module basic_5000_50000_5000_5_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xor U0 (N_0,In_4689,In_496);
xnor U1 (N_1,In_3829,In_2219);
nand U2 (N_2,In_464,In_4621);
and U3 (N_3,In_3310,In_4652);
or U4 (N_4,In_262,In_3231);
xor U5 (N_5,In_4396,In_1098);
nand U6 (N_6,In_1685,In_3352);
nand U7 (N_7,In_1339,In_638);
nand U8 (N_8,In_4196,In_4610);
nand U9 (N_9,In_377,In_4951);
xnor U10 (N_10,In_586,In_387);
or U11 (N_11,In_4439,In_4055);
or U12 (N_12,In_3712,In_4253);
or U13 (N_13,In_4500,In_4954);
nor U14 (N_14,In_769,In_1353);
and U15 (N_15,In_2069,In_1654);
or U16 (N_16,In_3279,In_766);
nor U17 (N_17,In_2142,In_548);
xor U18 (N_18,In_3610,In_42);
nand U19 (N_19,In_4090,In_3460);
nor U20 (N_20,In_3302,In_469);
xnor U21 (N_21,In_2736,In_4892);
xnor U22 (N_22,In_3463,In_3411);
xor U23 (N_23,In_1532,In_3818);
or U24 (N_24,In_314,In_1566);
and U25 (N_25,In_4879,In_4878);
xnor U26 (N_26,In_1198,In_2062);
nand U27 (N_27,In_4476,In_1838);
nand U28 (N_28,In_1483,In_4628);
nor U29 (N_29,In_514,In_3097);
or U30 (N_30,In_4542,In_1272);
or U31 (N_31,In_1173,In_4767);
and U32 (N_32,In_3237,In_3771);
nand U33 (N_33,In_765,In_3011);
nand U34 (N_34,In_352,In_1110);
xor U35 (N_35,In_575,In_679);
nor U36 (N_36,In_1722,In_2155);
nor U37 (N_37,In_3559,In_2930);
and U38 (N_38,In_4042,In_1292);
or U39 (N_39,In_2309,In_4522);
or U40 (N_40,In_1213,In_1236);
xor U41 (N_41,In_3933,In_4989);
and U42 (N_42,In_3077,In_2478);
nor U43 (N_43,In_3867,In_3092);
xnor U44 (N_44,In_4045,In_191);
nor U45 (N_45,In_58,In_3920);
and U46 (N_46,In_2541,In_1808);
and U47 (N_47,In_4785,In_748);
or U48 (N_48,In_2328,In_3700);
and U49 (N_49,In_1218,In_4204);
xnor U50 (N_50,In_1803,In_2368);
xor U51 (N_51,In_1958,In_2750);
xnor U52 (N_52,In_947,In_1644);
nand U53 (N_53,In_1643,In_4023);
nand U54 (N_54,In_1973,In_61);
or U55 (N_55,In_392,In_4386);
nand U56 (N_56,In_930,In_2709);
xor U57 (N_57,In_348,In_2582);
nand U58 (N_58,In_3655,In_3733);
and U59 (N_59,In_3013,In_310);
and U60 (N_60,In_1579,In_1814);
and U61 (N_61,In_862,In_3794);
or U62 (N_62,In_4289,In_4228);
nand U63 (N_63,In_3911,In_4885);
and U64 (N_64,In_1874,In_2792);
nor U65 (N_65,In_3975,In_4472);
or U66 (N_66,In_2795,In_3560);
nand U67 (N_67,In_1004,In_2801);
or U68 (N_68,In_3450,In_3654);
and U69 (N_69,In_1693,In_1165);
or U70 (N_70,In_825,In_509);
nor U71 (N_71,In_1488,In_1266);
nand U72 (N_72,In_2825,In_3935);
xor U73 (N_73,In_3034,In_863);
and U74 (N_74,In_357,In_3282);
nand U75 (N_75,In_751,In_3458);
nor U76 (N_76,In_4291,In_2776);
xor U77 (N_77,In_63,In_1791);
or U78 (N_78,In_64,In_2229);
nor U79 (N_79,In_2904,In_4708);
xnor U80 (N_80,In_4587,In_3909);
and U81 (N_81,In_3688,In_23);
or U82 (N_82,In_1856,In_4536);
xnor U83 (N_83,In_3495,In_1100);
xnor U84 (N_84,In_2338,In_3219);
nor U85 (N_85,In_3421,In_315);
xnor U86 (N_86,In_539,In_1556);
nor U87 (N_87,In_3455,In_3873);
nor U88 (N_88,In_270,In_396);
nor U89 (N_89,In_4457,In_15);
and U90 (N_90,In_2078,In_2608);
nand U91 (N_91,In_4188,In_1944);
and U92 (N_92,In_3950,In_2990);
nor U93 (N_93,In_3064,In_1438);
nand U94 (N_94,In_1805,In_2133);
xor U95 (N_95,In_794,In_2717);
xnor U96 (N_96,In_2244,In_4452);
xnor U97 (N_97,In_2361,In_3461);
or U98 (N_98,In_320,In_3457);
xor U99 (N_99,In_2479,In_4836);
xnor U100 (N_100,In_2282,In_4465);
or U101 (N_101,In_2176,In_4590);
xnor U102 (N_102,In_841,In_1385);
and U103 (N_103,In_3151,In_4846);
and U104 (N_104,In_4438,In_560);
nand U105 (N_105,In_275,In_4294);
and U106 (N_106,In_2392,In_532);
xor U107 (N_107,In_4506,In_1711);
and U108 (N_108,In_2198,In_2880);
nand U109 (N_109,In_1917,In_171);
nor U110 (N_110,In_3136,In_4533);
xor U111 (N_111,In_3965,In_3924);
and U112 (N_112,In_1321,In_478);
and U113 (N_113,In_2503,In_4895);
xnor U114 (N_114,In_790,In_4490);
and U115 (N_115,In_3084,In_4887);
xor U116 (N_116,In_1009,In_1696);
or U117 (N_117,In_699,In_594);
nand U118 (N_118,In_3387,In_434);
xnor U119 (N_119,In_604,In_4532);
nor U120 (N_120,In_3889,In_2033);
nand U121 (N_121,In_4557,In_2909);
and U122 (N_122,In_4283,In_374);
or U123 (N_123,In_2152,In_2914);
xor U124 (N_124,In_2651,In_4795);
nor U125 (N_125,In_3424,In_4877);
nor U126 (N_126,In_2784,In_292);
xor U127 (N_127,In_1204,In_3947);
xnor U128 (N_128,In_4526,In_2462);
or U129 (N_129,In_4872,In_3227);
nor U130 (N_130,In_4827,In_4300);
or U131 (N_131,In_1967,In_2046);
nor U132 (N_132,In_805,In_3747);
or U133 (N_133,In_2430,In_4194);
and U134 (N_134,In_1020,In_4241);
nand U135 (N_135,In_4029,In_2363);
nand U136 (N_136,In_4978,In_2094);
or U137 (N_137,In_1107,In_2639);
nand U138 (N_138,In_3540,In_1155);
nand U139 (N_139,In_4493,In_1143);
nand U140 (N_140,In_4984,In_569);
nand U141 (N_141,In_816,In_840);
nand U142 (N_142,In_1725,In_220);
nand U143 (N_143,In_1486,In_4317);
xnor U144 (N_144,In_4141,In_26);
xor U145 (N_145,In_2878,In_738);
or U146 (N_146,In_2369,In_3451);
or U147 (N_147,In_2104,In_2114);
nand U148 (N_148,In_1132,In_3659);
nor U149 (N_149,In_1773,In_1044);
nor U150 (N_150,In_2100,In_2339);
and U151 (N_151,In_940,In_1464);
nand U152 (N_152,In_3257,In_696);
and U153 (N_153,In_4786,In_4116);
or U154 (N_154,In_4694,In_3772);
nand U155 (N_155,In_1220,In_954);
or U156 (N_156,In_1749,In_1337);
nor U157 (N_157,In_2056,In_2386);
xnor U158 (N_158,In_2358,In_4809);
and U159 (N_159,In_824,In_4297);
nor U160 (N_160,In_1593,In_4709);
nor U161 (N_161,In_3614,In_4028);
nand U162 (N_162,In_4299,In_849);
and U163 (N_163,In_339,In_95);
nand U164 (N_164,In_1758,In_2247);
or U165 (N_165,In_4354,In_3472);
nor U166 (N_166,In_1855,In_3898);
or U167 (N_167,In_2236,In_4595);
and U168 (N_168,In_2168,In_3970);
and U169 (N_169,In_3521,In_729);
nand U170 (N_170,In_668,In_3797);
nor U171 (N_171,In_201,In_443);
nor U172 (N_172,In_4421,In_247);
or U173 (N_173,In_132,In_178);
and U174 (N_174,In_1957,In_3594);
nand U175 (N_175,In_2401,In_1407);
xor U176 (N_176,In_46,In_219);
and U177 (N_177,In_2970,In_1786);
or U178 (N_178,In_2992,In_926);
or U179 (N_179,In_2864,In_2558);
and U180 (N_180,In_1778,In_3531);
and U181 (N_181,In_2530,In_1502);
nand U182 (N_182,In_463,In_3022);
nand U183 (N_183,In_4169,In_3350);
nor U184 (N_184,In_4047,In_3895);
xor U185 (N_185,In_2972,In_1551);
and U186 (N_186,In_265,In_1179);
nand U187 (N_187,In_1421,In_1441);
xor U188 (N_188,In_3859,In_1028);
or U189 (N_189,In_4734,In_2111);
nor U190 (N_190,In_682,In_4470);
xnor U191 (N_191,In_284,In_4349);
or U192 (N_192,In_4560,In_268);
xor U193 (N_193,In_4637,In_1949);
and U194 (N_194,In_4927,In_2735);
nor U195 (N_195,In_2365,In_4365);
nor U196 (N_196,In_510,In_4655);
and U197 (N_197,In_3316,In_4469);
xnor U198 (N_198,In_3112,In_1365);
xor U199 (N_199,In_3108,In_2573);
nand U200 (N_200,In_4301,In_2492);
and U201 (N_201,In_3040,In_3364);
nor U202 (N_202,In_1592,In_924);
or U203 (N_203,In_4670,In_815);
nor U204 (N_204,In_2790,In_1095);
nor U205 (N_205,In_2256,In_3927);
and U206 (N_206,In_2669,In_2186);
nor U207 (N_207,In_3070,In_4935);
or U208 (N_208,In_3995,In_344);
and U209 (N_209,In_2729,In_1168);
nand U210 (N_210,In_2194,In_4458);
or U211 (N_211,In_2473,In_203);
or U212 (N_212,In_2683,In_163);
or U213 (N_213,In_1351,In_27);
xnor U214 (N_214,In_4504,In_237);
nand U215 (N_215,In_4156,In_1625);
and U216 (N_216,In_1982,In_2308);
nor U217 (N_217,In_1613,In_4074);
nor U218 (N_218,In_3519,In_4696);
or U219 (N_219,In_4171,In_752);
xor U220 (N_220,In_466,In_3726);
nand U221 (N_221,In_4960,In_231);
xnor U222 (N_222,In_801,In_508);
nand U223 (N_223,In_318,In_4048);
nand U224 (N_224,In_1058,In_4229);
nand U225 (N_225,In_3879,In_1118);
xnor U226 (N_226,In_3183,In_1871);
and U227 (N_227,In_880,In_4657);
nor U228 (N_228,In_1756,In_2918);
xnor U229 (N_229,In_1909,In_3695);
nor U230 (N_230,In_4890,In_2989);
nor U231 (N_231,In_4781,In_2635);
xor U232 (N_232,In_4161,In_4808);
nor U233 (N_233,In_2173,In_917);
nand U234 (N_234,In_932,In_2354);
xor U235 (N_235,In_2450,In_4408);
nand U236 (N_236,In_4736,In_4273);
nor U237 (N_237,In_4632,In_3915);
xor U238 (N_238,In_2845,In_762);
nor U239 (N_239,In_1907,In_2088);
nand U240 (N_240,In_4260,In_433);
and U241 (N_241,In_2484,In_1243);
or U242 (N_242,In_732,In_3557);
or U243 (N_243,In_3441,In_3131);
and U244 (N_244,In_2140,In_362);
nor U245 (N_245,In_2243,In_593);
nand U246 (N_246,In_2317,In_522);
or U247 (N_247,In_2756,In_4824);
nand U248 (N_248,In_2738,In_461);
or U249 (N_249,In_821,In_1499);
xor U250 (N_250,In_3994,In_4344);
nor U251 (N_251,In_553,In_931);
nand U252 (N_252,In_1210,In_717);
nor U253 (N_253,In_4605,In_167);
nor U254 (N_254,In_2642,In_1877);
and U255 (N_255,In_2894,In_235);
nor U256 (N_256,In_4036,In_1568);
nand U257 (N_257,In_2707,In_4946);
nand U258 (N_258,In_358,In_2858);
xor U259 (N_259,In_1211,In_115);
xor U260 (N_260,In_2252,In_4612);
or U261 (N_261,In_1661,In_3508);
nor U262 (N_262,In_3195,In_1624);
nor U263 (N_263,In_861,In_4309);
and U264 (N_264,In_436,In_3634);
and U265 (N_265,In_1746,In_492);
nand U266 (N_266,In_2139,In_4841);
or U267 (N_267,In_1987,In_3912);
xnor U268 (N_268,In_4661,In_3764);
xnor U269 (N_269,In_2287,In_3199);
or U270 (N_270,In_2120,In_4796);
nand U271 (N_271,In_3471,In_1699);
nor U272 (N_272,In_2004,In_4530);
or U273 (N_273,In_2819,In_1150);
or U274 (N_274,In_883,In_4627);
xor U275 (N_275,In_3033,In_2625);
or U276 (N_276,In_4963,In_4602);
nand U277 (N_277,In_3045,In_2267);
nand U278 (N_278,In_4281,In_2949);
xor U279 (N_279,In_3464,In_1806);
nand U280 (N_280,In_1854,In_2733);
nor U281 (N_281,In_2352,In_2440);
nand U282 (N_282,In_4370,In_4174);
or U283 (N_283,In_4412,In_4117);
nand U284 (N_284,In_4282,In_3256);
xnor U285 (N_285,In_1194,In_3869);
or U286 (N_286,In_4347,In_3354);
or U287 (N_287,In_2906,In_1999);
and U288 (N_288,In_4460,In_2629);
nor U289 (N_289,In_4712,In_2882);
nor U290 (N_290,In_2638,In_327);
nor U291 (N_291,In_3528,In_3565);
nor U292 (N_292,In_2432,In_2574);
or U293 (N_293,In_4749,In_1843);
xnor U294 (N_294,In_3403,In_3749);
nor U295 (N_295,In_2588,In_1043);
nand U296 (N_296,In_1373,In_481);
nor U297 (N_297,In_1347,In_2546);
xnor U298 (N_298,In_1108,In_19);
nor U299 (N_299,In_2178,In_2941);
xor U300 (N_300,In_4549,In_3174);
and U301 (N_301,In_1115,In_2675);
nand U302 (N_302,In_3903,In_2869);
and U303 (N_303,In_1175,In_991);
nor U304 (N_304,In_4553,In_335);
xor U305 (N_305,In_2065,In_2777);
nand U306 (N_306,In_3855,In_2705);
nor U307 (N_307,In_4276,In_1869);
or U308 (N_308,In_2595,In_3534);
or U309 (N_309,In_1775,In_1993);
and U310 (N_310,In_2911,In_3778);
or U311 (N_311,In_2877,In_1303);
xor U312 (N_312,In_2136,In_1608);
nor U313 (N_313,In_3459,In_2748);
xor U314 (N_314,In_457,In_874);
nor U315 (N_315,In_733,In_3505);
xnor U316 (N_316,In_1352,In_3288);
and U317 (N_317,In_3775,In_879);
or U318 (N_318,In_2859,In_2585);
xor U319 (N_319,In_2203,In_3117);
and U320 (N_320,In_3142,In_4513);
nor U321 (N_321,In_3916,In_1837);
and U322 (N_322,In_1338,In_1490);
nor U323 (N_323,In_4692,In_1586);
or U324 (N_324,In_4017,In_506);
or U325 (N_325,In_1291,In_1587);
nand U326 (N_326,In_1789,In_3913);
nand U327 (N_327,In_588,In_877);
and U328 (N_328,In_3544,In_4287);
nor U329 (N_329,In_383,In_3479);
xor U330 (N_330,In_1694,In_4288);
nand U331 (N_331,In_4883,In_1498);
nor U332 (N_332,In_1809,In_4999);
or U333 (N_333,In_4826,In_2150);
or U334 (N_334,In_2289,In_158);
nor U335 (N_335,In_4625,In_286);
nand U336 (N_336,In_1312,In_2596);
xor U337 (N_337,In_2232,In_1908);
or U338 (N_338,In_3653,In_937);
xor U339 (N_339,In_2307,In_1922);
xnor U340 (N_340,In_4973,In_2617);
or U341 (N_341,In_342,In_898);
and U342 (N_342,In_3500,In_1197);
and U343 (N_343,In_3574,In_2237);
nor U344 (N_344,In_1309,In_1757);
or U345 (N_345,In_1770,In_3577);
nor U346 (N_346,In_1406,In_4852);
and U347 (N_347,In_2161,In_332);
and U348 (N_348,In_304,In_533);
nand U349 (N_349,In_3320,In_4318);
nand U350 (N_350,In_995,In_3446);
nor U351 (N_351,In_126,In_3192);
nand U352 (N_352,In_1193,In_1015);
nor U353 (N_353,In_3334,In_2843);
nor U354 (N_354,In_2905,In_4710);
nor U355 (N_355,In_1,In_3906);
xor U356 (N_356,In_1578,In_4402);
xnor U357 (N_357,In_2362,In_4925);
xor U358 (N_358,In_2895,In_2632);
and U359 (N_359,In_4975,In_296);
nor U360 (N_360,In_345,In_970);
or U361 (N_361,In_4085,In_28);
and U362 (N_362,In_1129,In_886);
nor U363 (N_363,In_1708,In_1176);
or U364 (N_364,In_1620,In_3072);
xnor U365 (N_365,In_2476,In_4304);
xor U366 (N_366,In_1336,In_1430);
or U367 (N_367,In_2722,In_1847);
xnor U368 (N_368,In_3709,In_2245);
nor U369 (N_369,In_759,In_1230);
and U370 (N_370,In_31,In_1422);
or U371 (N_371,In_4364,In_3760);
xor U372 (N_372,In_2725,In_2066);
xnor U373 (N_373,In_3135,In_2223);
xnor U374 (N_374,In_254,In_1202);
nor U375 (N_375,In_3333,In_2189);
xor U376 (N_376,In_3941,In_3419);
nor U377 (N_377,In_2837,In_1027);
xor U378 (N_378,In_412,In_3746);
and U379 (N_379,In_3272,In_798);
xor U380 (N_380,In_1600,In_1637);
and U381 (N_381,In_667,In_4166);
nand U382 (N_382,In_3851,In_225);
xnor U383 (N_383,In_4389,In_1269);
nor U384 (N_384,In_4144,In_1879);
nand U385 (N_385,In_431,In_1133);
or U386 (N_386,In_1656,In_2019);
nand U387 (N_387,In_4818,In_2118);
nand U388 (N_388,In_1077,In_1641);
nand U389 (N_389,In_1961,In_2041);
nor U390 (N_390,In_4268,In_1583);
or U391 (N_391,In_2405,In_4149);
xnor U392 (N_392,In_3856,In_417);
nor U393 (N_393,In_118,In_1295);
nor U394 (N_394,In_1283,In_3285);
nand U395 (N_395,In_3510,In_2431);
nor U396 (N_396,In_1258,In_3787);
xor U397 (N_397,In_1889,In_1327);
nor U398 (N_398,In_3551,In_1041);
or U399 (N_399,In_2811,In_3809);
nor U400 (N_400,In_4782,In_2598);
xnor U401 (N_401,In_4740,In_705);
and U402 (N_402,In_1911,In_1942);
nor U403 (N_403,In_2985,In_3188);
or U404 (N_404,In_2318,In_1774);
nand U405 (N_405,In_1163,In_2716);
or U406 (N_406,In_105,In_1975);
nand U407 (N_407,In_274,In_4966);
and U408 (N_408,In_2402,In_3762);
or U409 (N_409,In_3669,In_370);
nand U410 (N_410,In_1687,In_4444);
xnor U411 (N_411,In_890,In_2006);
xor U412 (N_412,In_897,In_3862);
or U413 (N_413,In_4145,In_4053);
nand U414 (N_414,In_1609,In_606);
nor U415 (N_415,In_2517,In_4003);
xnor U416 (N_416,In_3175,In_4494);
or U417 (N_417,In_3093,In_1793);
nor U418 (N_418,In_2965,In_2994);
or U419 (N_419,In_2523,In_1867);
and U420 (N_420,In_3041,In_3098);
and U421 (N_421,In_4860,In_987);
or U422 (N_422,In_3946,In_4051);
nand U423 (N_423,In_4030,In_3109);
or U424 (N_424,In_4934,In_706);
nor U425 (N_425,In_159,In_2209);
nand U426 (N_426,In_662,In_317);
xor U427 (N_427,In_108,In_285);
and U428 (N_428,In_2991,In_1648);
or U429 (N_429,In_4216,In_3398);
xor U430 (N_430,In_3523,In_623);
xnor U431 (N_431,In_4721,In_3622);
and U432 (N_432,In_2800,In_4009);
or U433 (N_433,In_1745,In_4018);
and U434 (N_434,In_1304,In_3373);
nor U435 (N_435,In_360,In_2891);
or U436 (N_436,In_110,In_4377);
nand U437 (N_437,In_3966,In_3542);
and U438 (N_438,In_4013,In_3481);
or U439 (N_439,In_1263,In_1622);
or U440 (N_440,In_4608,In_1316);
xnor U441 (N_441,In_633,In_4983);
or U442 (N_442,In_4544,In_473);
xor U443 (N_443,In_3843,In_4947);
nand U444 (N_444,In_3005,In_800);
nor U445 (N_445,In_2141,In_1456);
or U446 (N_446,In_3020,In_107);
or U447 (N_447,In_4683,In_2148);
and U448 (N_448,In_1423,In_2132);
nor U449 (N_449,In_1315,In_480);
or U450 (N_450,In_3805,In_4578);
xor U451 (N_451,In_1461,In_1599);
nor U452 (N_452,In_1826,In_2332);
nor U453 (N_453,In_2958,In_2117);
or U454 (N_454,In_4168,In_2922);
nand U455 (N_455,In_845,In_4286);
or U456 (N_456,In_228,In_4005);
and U457 (N_457,In_2953,In_3454);
and U458 (N_458,In_1181,In_4611);
nor U459 (N_459,In_2760,In_2039);
and U460 (N_460,In_1083,In_4640);
or U461 (N_461,In_3368,In_249);
xnor U462 (N_462,In_3187,In_2907);
or U463 (N_463,In_3453,In_3325);
or U464 (N_464,In_3046,In_1933);
nor U465 (N_465,In_3917,In_18);
and U466 (N_466,In_3021,In_3800);
nor U467 (N_467,In_2863,In_3707);
or U468 (N_468,In_2516,In_1189);
and U469 (N_469,In_2359,In_213);
or U470 (N_470,In_3740,In_1081);
nor U471 (N_471,In_1192,In_1686);
nand U472 (N_472,In_1726,In_2269);
xor U473 (N_473,In_1507,In_299);
or U474 (N_474,In_4898,In_414);
xnor U475 (N_475,In_1974,In_1635);
nor U476 (N_476,In_4008,In_3821);
nor U477 (N_477,In_1362,In_3576);
nor U478 (N_478,In_3095,In_2197);
nor U479 (N_479,In_4772,In_151);
and U480 (N_480,In_40,In_9);
and U481 (N_481,In_2337,In_1816);
or U482 (N_482,In_2589,In_1396);
nor U483 (N_483,In_986,In_572);
nand U484 (N_484,In_649,In_635);
nand U485 (N_485,In_493,In_1207);
nor U486 (N_486,In_437,In_4487);
nand U487 (N_487,In_4019,In_1807);
nand U488 (N_488,In_226,In_3602);
nand U489 (N_489,In_1704,In_2013);
nand U490 (N_490,In_4964,In_441);
nand U491 (N_491,In_2242,In_20);
nand U492 (N_492,In_2902,In_3765);
or U493 (N_493,In_84,In_1302);
and U494 (N_494,In_723,In_3491);
and U495 (N_495,In_4134,In_1997);
nor U496 (N_496,In_4691,In_904);
and U497 (N_497,In_1506,In_279);
or U498 (N_498,In_3679,In_1576);
and U499 (N_499,In_74,In_4894);
and U500 (N_500,In_1567,In_2619);
nor U501 (N_501,In_967,In_1006);
and U502 (N_502,In_3284,In_4056);
or U503 (N_503,In_1349,In_372);
and U504 (N_504,In_4434,In_3864);
xnor U505 (N_505,In_3023,In_3832);
or U506 (N_506,In_3845,In_3944);
or U507 (N_507,In_2655,In_1674);
nor U508 (N_508,In_4523,In_1870);
nand U509 (N_509,In_1493,In_3330);
nand U510 (N_510,In_2439,In_2881);
xnor U511 (N_511,In_4131,In_2694);
and U512 (N_512,In_4150,In_2908);
nor U513 (N_513,In_922,In_1395);
and U514 (N_514,In_4725,In_3415);
nand U515 (N_515,In_4183,In_94);
nand U516 (N_516,In_1389,In_2520);
nor U517 (N_517,In_2979,In_4695);
and U518 (N_518,In_4077,In_1345);
and U519 (N_519,In_1581,In_3866);
xor U520 (N_520,In_4035,In_4);
nor U521 (N_521,In_2112,In_2633);
nand U522 (N_522,In_36,In_1765);
and U523 (N_523,In_3919,In_3595);
or U524 (N_524,In_3937,In_1671);
and U525 (N_525,In_465,In_2701);
or U526 (N_526,In_557,In_2171);
or U527 (N_527,In_287,In_3342);
xnor U528 (N_528,In_4121,In_1896);
nor U529 (N_529,In_2437,In_3969);
or U530 (N_530,In_3721,In_4034);
nor U531 (N_531,In_4011,In_4499);
xnor U532 (N_532,In_810,In_4345);
nor U533 (N_533,In_3308,In_1501);
and U534 (N_534,In_3128,In_354);
nor U535 (N_535,In_1597,In_2315);
nand U536 (N_536,In_1380,In_485);
nand U537 (N_537,In_536,In_3028);
xnor U538 (N_538,In_12,In_1307);
nand U539 (N_539,In_1753,In_1364);
nand U540 (N_540,In_3720,In_144);
and U541 (N_541,In_2248,In_757);
nor U542 (N_542,In_1730,In_4264);
nand U543 (N_543,In_497,In_8);
xnor U544 (N_544,In_2191,In_1036);
and U545 (N_545,In_2156,In_1102);
nand U546 (N_546,In_1392,In_1950);
nand U547 (N_547,In_4897,In_2326);
nand U548 (N_548,In_1741,In_4777);
nor U549 (N_549,In_3608,In_1184);
or U550 (N_550,In_3872,In_3477);
or U551 (N_551,In_3370,In_2531);
nor U552 (N_552,In_4323,In_1051);
nor U553 (N_553,In_1899,In_4832);
and U554 (N_554,In_470,In_4780);
nor U555 (N_555,In_2544,In_3616);
xor U556 (N_556,In_4060,In_1138);
nor U557 (N_557,In_3423,In_876);
nand U558 (N_558,In_3340,In_3759);
nor U559 (N_559,In_1090,In_1473);
xnor U560 (N_560,In_3893,In_634);
and U561 (N_561,In_3049,In_1085);
nor U562 (N_562,In_2600,In_3786);
nand U563 (N_563,In_4037,In_3179);
nor U564 (N_564,In_184,In_2592);
nor U565 (N_565,In_2491,In_56);
xnor U566 (N_566,In_4212,In_3561);
xnor U567 (N_567,In_4997,In_3074);
and U568 (N_568,In_4580,In_3734);
or U569 (N_569,In_3948,In_1744);
or U570 (N_570,In_4118,In_3428);
xor U571 (N_571,In_2715,In_121);
nand U572 (N_572,In_3611,In_4910);
nand U573 (N_573,In_4679,In_2389);
or U574 (N_574,In_2355,In_3305);
nand U575 (N_575,In_1013,In_685);
and U576 (N_576,In_4546,In_1640);
or U577 (N_577,In_1480,In_331);
or U578 (N_578,In_1690,In_3846);
nor U579 (N_579,In_1530,In_1172);
or U580 (N_580,In_665,In_2043);
xor U581 (N_581,In_1658,In_399);
nand U582 (N_582,In_4851,In_4098);
xnor U583 (N_583,In_888,In_1073);
nor U584 (N_584,In_2193,In_4848);
or U585 (N_585,In_600,In_3138);
or U586 (N_586,In_3071,In_4385);
xnor U587 (N_587,In_3629,In_4352);
nand U588 (N_588,In_1403,In_4728);
nor U589 (N_589,In_4329,In_3512);
nor U590 (N_590,In_1817,In_686);
nor U591 (N_591,In_1278,In_356);
nand U592 (N_592,In_170,In_517);
nor U593 (N_593,In_1802,In_3717);
and U594 (N_594,In_4496,In_1589);
and U595 (N_595,In_3804,In_2438);
nor U596 (N_596,In_2260,In_3784);
or U597 (N_597,In_2723,In_4341);
or U598 (N_598,In_4641,In_242);
nor U599 (N_599,In_3918,In_13);
nand U600 (N_600,In_1078,In_2003);
or U601 (N_601,In_2565,In_4160);
xor U602 (N_602,In_3957,In_3921);
xnor U603 (N_603,In_1662,In_3303);
or U604 (N_604,In_4124,In_3766);
nor U605 (N_605,In_81,In_3353);
or U606 (N_606,In_4337,In_3537);
nand U607 (N_607,In_2665,In_384);
xor U608 (N_608,In_2384,In_2350);
nand U609 (N_609,In_3991,In_197);
nand U610 (N_610,In_3413,In_647);
xnor U611 (N_611,In_3753,In_3696);
xor U612 (N_612,In_2645,In_428);
xnor U613 (N_613,In_4269,In_951);
nand U614 (N_614,In_1147,In_2929);
or U615 (N_615,In_2449,In_2844);
and U616 (N_616,In_725,In_91);
xnor U617 (N_617,In_646,In_4440);
xnor U618 (N_618,In_1117,In_1963);
nand U619 (N_619,In_2076,In_4103);
or U620 (N_620,In_1076,In_288);
and U621 (N_621,In_373,In_1019);
and U622 (N_622,In_2964,In_3882);
nand U623 (N_623,In_4609,In_2275);
nand U624 (N_624,In_519,In_3374);
nor U625 (N_625,In_3852,In_208);
or U626 (N_626,In_2628,In_277);
or U627 (N_627,In_2444,In_3545);
and U628 (N_628,In_1404,In_3067);
nor U629 (N_629,In_2578,In_2077);
or U630 (N_630,In_4367,In_4007);
and U631 (N_631,In_4516,In_985);
and U632 (N_632,In_2082,In_4682);
or U633 (N_633,In_3819,In_3587);
and U634 (N_634,In_3684,In_4662);
nand U635 (N_635,In_3026,In_3767);
nor U636 (N_636,In_1399,In_4073);
xor U637 (N_637,In_885,In_4020);
nand U638 (N_638,In_581,In_4825);
and U639 (N_639,In_1684,In_599);
and U640 (N_640,In_1617,In_1035);
or U641 (N_641,In_4217,In_1529);
or U642 (N_642,In_655,In_2433);
xor U643 (N_643,In_963,In_4479);
xor U644 (N_644,In_1925,In_1135);
nor U645 (N_645,In_4126,In_1196);
nand U646 (N_646,In_3184,In_784);
nor U647 (N_647,In_4847,In_2959);
nor U648 (N_648,In_4958,In_487);
nor U649 (N_649,In_4477,In_60);
nand U650 (N_650,In_2306,In_3376);
and U651 (N_651,In_1415,In_472);
and U652 (N_652,In_2455,In_4914);
or U653 (N_653,In_4733,In_1029);
xnor U654 (N_654,In_4266,In_4693);
nand U655 (N_655,In_1571,In_3152);
xor U656 (N_656,In_1458,In_4673);
or U657 (N_657,In_2657,In_1956);
xor U658 (N_658,In_113,In_2137);
and U659 (N_659,In_1737,In_826);
xor U660 (N_660,In_3914,In_3763);
or U661 (N_661,In_223,In_4940);
and U662 (N_662,In_3019,In_3748);
nor U663 (N_663,In_4697,In_3094);
or U664 (N_664,In_1522,In_4739);
and U665 (N_665,In_2413,In_395);
nand U666 (N_666,In_1951,In_4591);
xnor U667 (N_667,In_4766,In_3673);
and U668 (N_668,In_3632,In_4139);
nand U669 (N_669,In_4445,In_956);
nor U670 (N_670,In_3051,In_111);
nor U671 (N_671,In_1565,In_3892);
nor U672 (N_672,In_3548,In_4142);
or U673 (N_673,In_4091,In_2280);
nand U674 (N_674,In_516,In_524);
or U675 (N_675,In_1892,In_983);
nor U676 (N_676,In_2034,In_1820);
xnor U677 (N_677,In_591,In_4653);
or U678 (N_678,In_920,In_3004);
nand U679 (N_679,In_3671,In_799);
nor U680 (N_680,In_739,In_3546);
or U681 (N_681,In_2872,In_4856);
or U682 (N_682,In_537,In_1865);
or U683 (N_683,In_3171,In_2488);
or U684 (N_684,In_1279,In_3890);
and U685 (N_685,In_2264,In_3036);
nor U686 (N_686,In_1358,In_4775);
or U687 (N_687,In_1538,In_1411);
and U688 (N_688,In_4380,In_1825);
nor U689 (N_689,In_4012,In_2797);
nor U690 (N_690,In_3249,In_2862);
and U691 (N_691,In_2072,In_3384);
or U692 (N_692,In_2997,In_4569);
nor U693 (N_693,In_3939,In_4044);
nor U694 (N_694,In_294,In_1564);
and U695 (N_695,In_1828,In_1439);
or U696 (N_696,In_2680,In_2390);
nand U697 (N_697,In_3943,In_866);
nor U698 (N_698,In_4774,In_1893);
or U699 (N_699,In_4135,In_997);
and U700 (N_700,In_2765,In_333);
or U701 (N_701,In_871,In_4561);
nand U702 (N_702,In_1002,In_3828);
or U703 (N_703,In_101,In_153);
and U704 (N_704,In_1428,In_1325);
xor U705 (N_705,In_4950,In_2210);
nand U706 (N_706,In_571,In_4057);
and U707 (N_707,In_4737,In_4665);
nand U708 (N_708,In_4511,In_2090);
xor U709 (N_709,In_258,In_4398);
xnor U710 (N_710,In_4735,In_2299);
nor U711 (N_711,In_474,In_823);
nand U712 (N_712,In_1324,In_1733);
and U713 (N_713,In_4061,In_4251);
xnor U714 (N_714,In_2606,In_2936);
and U715 (N_715,In_4550,In_619);
nand U716 (N_716,In_4944,In_4218);
nor U717 (N_717,In_3292,In_71);
nor U718 (N_718,In_1187,In_1721);
or U719 (N_719,In_1985,In_2551);
and U720 (N_720,In_1229,In_637);
nand U721 (N_721,In_1039,In_4209);
nor U722 (N_722,In_2427,In_2157);
nand U723 (N_723,In_835,In_2831);
and U724 (N_724,In_2356,In_1299);
nor U725 (N_725,In_527,In_3147);
and U726 (N_726,In_2266,In_4065);
xor U727 (N_727,In_1882,In_906);
nor U728 (N_728,In_2696,In_2560);
and U729 (N_729,In_2559,In_4575);
nor U730 (N_730,In_1842,In_2278);
nand U731 (N_731,In_2621,In_4327);
and U732 (N_732,In_3811,In_3631);
nor U733 (N_733,In_1419,In_4998);
xnor U734 (N_734,In_1827,In_2028);
and U735 (N_735,In_2029,In_1429);
xor U736 (N_736,In_341,In_4762);
and U737 (N_737,In_4510,In_3822);
nand U738 (N_738,In_4994,In_4527);
nand U739 (N_739,In_4664,In_393);
or U740 (N_740,In_4443,In_298);
nand U741 (N_741,In_3048,In_4741);
nand U742 (N_742,In_1088,In_737);
nand U743 (N_743,In_4338,In_283);
xor U744 (N_744,In_2938,In_4384);
or U745 (N_745,In_4816,In_4159);
and U746 (N_746,In_4334,In_1841);
and U747 (N_747,In_3329,In_1573);
nand U748 (N_748,In_4348,In_1618);
nand U749 (N_749,In_2089,In_252);
or U750 (N_750,In_3953,In_3168);
xor U751 (N_751,In_839,In_351);
nand U752 (N_752,In_2841,In_1514);
and U753 (N_753,In_673,In_1251);
xnor U754 (N_754,In_185,In_4779);
nand U755 (N_755,In_1692,In_475);
and U756 (N_756,In_1768,In_3210);
and U757 (N_757,In_1367,In_654);
nor U758 (N_758,In_3444,In_4122);
xnor U759 (N_759,In_3897,In_2037);
and U760 (N_760,In_186,In_3752);
xnor U761 (N_761,In_1160,In_2480);
nand U762 (N_762,In_2641,In_32);
or U763 (N_763,In_2730,In_369);
xor U764 (N_764,In_3322,In_858);
or U765 (N_765,In_421,In_631);
nor U766 (N_766,In_4226,In_1798);
or U767 (N_767,In_102,In_3445);
nor U768 (N_768,In_2182,In_3000);
xnor U769 (N_769,In_3264,In_2091);
xnor U770 (N_770,In_1519,In_4456);
xnor U771 (N_771,In_1859,In_4538);
nand U772 (N_772,In_4190,In_2321);
and U773 (N_773,In_2216,In_2700);
and U774 (N_774,In_3990,In_1771);
nor U775 (N_775,In_1391,In_3888);
or U776 (N_776,In_119,In_4486);
nand U777 (N_777,In_1575,In_404);
nand U778 (N_778,In_3185,In_2017);
nand U779 (N_779,In_3620,In_774);
xnor U780 (N_780,In_3258,In_68);
or U781 (N_781,In_2257,In_3079);
nand U782 (N_782,In_1208,In_2461);
nand U783 (N_783,In_2703,In_4814);
or U784 (N_784,In_267,In_652);
nor U785 (N_785,In_4478,In_2008);
and U786 (N_786,In_3666,In_302);
nand U787 (N_787,In_3863,In_3774);
nand U788 (N_788,In_1886,In_3609);
xnor U789 (N_789,In_3420,In_4473);
and U790 (N_790,In_3357,In_1782);
and U791 (N_791,In_2031,In_397);
or U792 (N_792,In_4813,In_4639);
or U793 (N_793,In_914,In_2052);
xor U794 (N_794,In_1249,In_2061);
and U795 (N_795,In_3278,In_609);
xnor U796 (N_796,In_3416,In_1393);
nand U797 (N_797,In_744,In_3346);
nand U798 (N_798,In_2984,In_3960);
nand U799 (N_799,In_1082,In_238);
nand U800 (N_800,In_4913,In_2622);
nor U801 (N_801,In_4865,In_1544);
and U802 (N_802,In_1594,In_4604);
and U803 (N_803,In_232,In_3955);
or U804 (N_804,In_141,In_2235);
nor U805 (N_805,In_3377,In_848);
xor U806 (N_806,In_543,In_2372);
nor U807 (N_807,In_1158,In_1990);
or U808 (N_808,In_4672,In_127);
and U809 (N_809,In_2828,In_4422);
and U810 (N_810,In_4588,In_1813);
xor U811 (N_811,In_2806,In_2810);
or U812 (N_812,In_245,In_2131);
and U813 (N_813,In_155,In_2887);
nand U814 (N_814,In_1190,In_4724);
xnor U815 (N_815,In_1094,In_2227);
nor U816 (N_816,In_4936,In_2671);
or U817 (N_817,In_1446,In_2927);
and U818 (N_818,In_2233,In_2956);
or U819 (N_819,In_3932,In_3743);
nor U820 (N_820,In_2125,In_3473);
or U821 (N_821,In_4409,In_2714);
nand U822 (N_822,In_4497,In_3238);
nand U823 (N_823,In_1947,In_1785);
and U824 (N_824,In_881,In_1790);
nand U825 (N_825,In_1862,In_3641);
and U826 (N_826,In_608,In_2815);
or U827 (N_827,In_1885,In_2348);
nor U828 (N_828,In_4292,In_2153);
nor U829 (N_829,In_3002,In_1235);
xnor U830 (N_830,In_2102,In_1524);
xor U831 (N_831,In_2873,In_3299);
xnor U832 (N_832,In_812,In_1833);
xnor U833 (N_833,In_2202,In_2647);
nand U834 (N_834,In_3328,In_3209);
xnor U835 (N_835,In_114,In_3059);
and U836 (N_836,In_4539,In_2802);
xnor U837 (N_837,In_1319,In_2720);
xor U838 (N_838,In_584,In_3780);
nor U839 (N_839,In_656,In_453);
nand U840 (N_840,In_1462,In_2923);
and U841 (N_841,In_2961,In_4907);
xor U842 (N_842,In_1517,In_4981);
xnor U843 (N_843,In_1267,In_2283);
and U844 (N_844,In_3283,In_4761);
or U845 (N_845,In_313,In_544);
nor U846 (N_846,In_4649,In_4915);
nor U847 (N_847,In_1751,In_1167);
or U848 (N_848,In_4770,In_3114);
or U849 (N_849,In_518,In_2080);
xnor U850 (N_850,In_2940,In_4176);
nor U851 (N_851,In_4001,In_4830);
or U852 (N_852,In_2667,In_1559);
xor U853 (N_853,In_2279,In_2505);
nand U854 (N_854,In_1800,In_1830);
or U855 (N_855,In_2509,In_1151);
xor U856 (N_856,In_1646,In_4684);
nor U857 (N_857,In_546,In_1122);
xor U858 (N_858,In_2803,In_2086);
or U859 (N_859,In_2172,In_1436);
or U860 (N_860,In_1274,In_1125);
and U861 (N_861,In_243,In_1127);
nand U862 (N_862,In_282,In_780);
nor U863 (N_863,In_303,In_3844);
or U864 (N_864,In_194,In_2347);
and U865 (N_865,In_3986,In_952);
xnor U866 (N_866,In_3761,In_4718);
nand U867 (N_867,In_4675,In_929);
nor U868 (N_868,In_2495,In_3332);
nand U869 (N_869,In_4688,In_2251);
nor U870 (N_870,In_640,In_2977);
xnor U871 (N_871,In_2255,In_3567);
or U872 (N_872,In_3599,In_321);
or U873 (N_873,In_4336,In_411);
or U874 (N_874,In_378,In_1120);
nor U875 (N_875,In_2510,In_1543);
nand U876 (N_876,In_3,In_2698);
nor U877 (N_877,In_3738,In_1651);
nand U878 (N_878,In_4324,In_4622);
xor U879 (N_879,In_37,In_504);
xnor U880 (N_880,In_959,In_1679);
nor U881 (N_881,In_1159,In_830);
nor U882 (N_882,In_4014,In_4939);
nand U883 (N_883,In_4520,In_1141);
nand U884 (N_884,In_1943,In_795);
nor U885 (N_885,In_4659,In_375);
or U886 (N_886,In_2110,In_773);
xnor U887 (N_887,In_479,In_4298);
and U888 (N_888,In_664,In_2577);
and U889 (N_889,In_125,In_3372);
and U890 (N_890,In_2752,In_1705);
nand U891 (N_891,In_636,In_3490);
or U892 (N_892,In_4010,In_4491);
and U893 (N_893,In_1067,In_2407);
or U894 (N_894,In_2870,In_3160);
and U895 (N_895,In_1759,In_2420);
nor U896 (N_896,In_2555,In_3113);
nand U897 (N_897,In_2556,In_2853);
and U898 (N_898,In_2623,In_3216);
nand U899 (N_899,In_1901,In_4004);
nor U900 (N_900,In_2011,In_1418);
xor U901 (N_901,In_4249,In_4203);
nor U902 (N_902,In_1823,In_1959);
xor U903 (N_903,In_3690,In_887);
or U904 (N_904,In_4647,In_2597);
nor U905 (N_905,In_2519,In_2458);
nor U906 (N_906,In_70,In_2434);
and U907 (N_907,In_3392,In_3793);
or U908 (N_908,In_1045,In_3101);
or U909 (N_909,In_3744,In_3550);
nor U910 (N_910,In_989,In_1478);
and U911 (N_911,In_3563,In_3498);
nor U912 (N_912,In_1154,In_3198);
or U913 (N_913,In_3642,In_834);
nor U914 (N_914,In_2313,In_4650);
and U915 (N_915,In_3930,In_1669);
and U916 (N_916,In_3436,In_2409);
or U917 (N_917,In_945,In_3881);
nor U918 (N_918,In_2852,In_4731);
nor U919 (N_919,In_3482,In_666);
xnor U920 (N_920,In_1386,In_2687);
xor U921 (N_921,In_4503,In_893);
nor U922 (N_922,In_3166,In_2839);
nor U923 (N_923,In_3061,In_4238);
xor U924 (N_924,In_836,In_3493);
xnor U925 (N_925,In_1977,In_2045);
or U926 (N_926,In_580,In_1145);
and U927 (N_927,In_4797,In_3295);
and U928 (N_928,In_1284,In_2987);
or U929 (N_929,In_3723,In_1927);
nor U930 (N_930,In_1616,In_3589);
xnor U931 (N_931,In_4932,In_1216);
xor U932 (N_932,In_3725,In_2614);
xnor U933 (N_933,In_4558,In_842);
nand U934 (N_934,In_2016,In_329);
nand U935 (N_935,In_2471,In_680);
nand U936 (N_936,In_3596,In_1388);
nand U937 (N_937,In_2654,In_1465);
and U938 (N_938,In_971,In_540);
nor U939 (N_939,In_192,In_4058);
nor U940 (N_940,In_4075,In_3683);
xnor U941 (N_941,In_3399,In_1520);
and U942 (N_942,In_448,In_255);
or U943 (N_943,In_3541,In_530);
and U944 (N_944,In_3096,In_3139);
and U945 (N_945,In_3954,In_1032);
xor U946 (N_946,In_2653,In_701);
or U947 (N_947,In_1864,In_2526);
nand U948 (N_948,In_4889,In_642);
nor U949 (N_949,In_183,In_703);
or U950 (N_950,In_3039,In_4668);
or U951 (N_951,In_4943,In_1994);
and U952 (N_952,In_408,In_1719);
nor U953 (N_953,In_727,In_4867);
xor U954 (N_954,In_2821,In_1205);
nor U955 (N_955,In_2371,In_2221);
xnor U956 (N_956,In_4427,In_875);
nor U957 (N_957,In_2529,In_4070);
and U958 (N_958,In_236,In_1186);
nand U959 (N_959,In_2913,In_3027);
xor U960 (N_960,In_614,In_2496);
xnor U961 (N_961,In_4446,In_2166);
nand U962 (N_962,In_4311,In_4455);
nor U963 (N_963,In_4568,In_3504);
xor U964 (N_964,In_2415,In_338);
xor U965 (N_965,In_1981,In_561);
nand U966 (N_966,In_1308,In_982);
or U967 (N_967,In_3637,In_1334);
nand U968 (N_968,In_4577,In_2201);
and U969 (N_969,In_2485,In_3047);
or U970 (N_970,In_2366,In_4252);
nor U971 (N_971,In_2652,In_3452);
nand U972 (N_972,In_2793,In_214);
or U973 (N_973,In_1131,In_3830);
or U974 (N_974,In_2605,In_29);
and U975 (N_975,In_1162,In_164);
xnor U976 (N_976,In_1653,In_3757);
xnor U977 (N_977,In_4677,In_429);
nor U978 (N_978,In_2609,In_2751);
and U979 (N_979,In_3854,In_2636);
xor U980 (N_980,In_1743,In_4207);
nor U981 (N_981,In_4069,In_4346);
nor U982 (N_982,In_4801,In_3526);
and U983 (N_983,In_659,In_2380);
nand U984 (N_984,In_143,In_758);
or U985 (N_985,In_3358,In_793);
nand U986 (N_986,In_4049,In_3409);
xor U987 (N_987,In_1232,In_1096);
xor U988 (N_988,In_2002,In_3676);
nor U989 (N_989,In_1873,In_21);
and U990 (N_990,In_4080,In_3180);
nor U991 (N_991,In_1424,In_761);
and U992 (N_992,In_4246,In_502);
and U993 (N_993,In_4182,In_4078);
xnor U994 (N_994,In_4369,In_4988);
and U995 (N_995,In_4451,In_2001);
or U996 (N_996,In_4108,In_1063);
nand U997 (N_997,In_4991,In_4381);
nand U998 (N_998,In_2774,In_2593);
and U999 (N_999,In_2830,In_3014);
xnor U1000 (N_1000,In_894,In_711);
or U1001 (N_1001,In_583,In_3750);
or U1002 (N_1002,In_2188,In_3024);
and U1003 (N_1003,In_1093,In_3251);
and U1004 (N_1004,In_1881,In_4064);
xnor U1005 (N_1005,In_2789,In_1425);
or U1006 (N_1006,In_2950,In_1233);
xor U1007 (N_1007,In_3337,In_1534);
or U1008 (N_1008,In_4485,In_1432);
nor U1009 (N_1009,In_661,In_4133);
nor U1010 (N_1010,In_622,In_3886);
xor U1011 (N_1011,In_4063,In_2360);
and U1012 (N_1012,In_768,In_4900);
and U1013 (N_1013,In_2406,In_1289);
nand U1014 (N_1014,In_4153,In_4589);
xnor U1015 (N_1015,In_3682,In_4823);
or U1016 (N_1016,In_216,In_1760);
or U1017 (N_1017,In_4844,In_3971);
nand U1018 (N_1018,In_3215,In_6);
xor U1019 (N_1019,In_4919,In_3901);
and U1020 (N_1020,In_4886,In_4756);
or U1021 (N_1021,In_4198,In_3476);
nor U1022 (N_1022,In_4177,In_3137);
and U1023 (N_1023,In_4101,In_2754);
and U1024 (N_1024,In_2610,In_2504);
nor U1025 (N_1025,In_3974,In_4106);
nand U1026 (N_1026,In_1991,In_674);
or U1027 (N_1027,In_1742,In_3081);
or U1028 (N_1028,In_2986,In_4437);
nor U1029 (N_1029,In_4937,In_783);
nor U1030 (N_1030,In_1912,In_2115);
nor U1031 (N_1031,In_4104,In_2612);
nand U1032 (N_1032,In_3085,In_1557);
xor U1033 (N_1033,In_3525,In_4043);
nand U1034 (N_1034,In_2270,In_3520);
nor U1035 (N_1035,In_1598,In_3087);
nand U1036 (N_1036,In_554,In_980);
nand U1037 (N_1037,In_3391,In_3107);
and U1038 (N_1038,In_4850,In_3486);
xor U1039 (N_1039,In_2231,In_4272);
nor U1040 (N_1040,In_446,In_2866);
nand U1041 (N_1041,In_992,In_658);
and U1042 (N_1042,In_512,In_2381);
nor U1043 (N_1043,In_204,In_817);
nor U1044 (N_1044,In_4373,In_697);
nor U1045 (N_1045,In_4441,In_3985);
or U1046 (N_1046,In_4667,In_2749);
xor U1047 (N_1047,In_1071,In_2327);
xnor U1048 (N_1048,In_2304,In_1516);
nor U1049 (N_1049,In_4505,In_1915);
nand U1050 (N_1050,In_511,In_388);
nor U1051 (N_1051,In_2846,In_3153);
xor U1052 (N_1052,In_3701,In_1852);
or U1053 (N_1053,In_4219,In_4599);
nor U1054 (N_1054,In_882,In_2340);
or U1055 (N_1055,In_916,In_4332);
xor U1056 (N_1056,In_4243,In_2935);
nand U1057 (N_1057,In_273,In_422);
or U1058 (N_1058,In_3447,In_2027);
nor U1059 (N_1059,In_4214,In_909);
and U1060 (N_1060,In_1268,In_3043);
nand U1061 (N_1061,In_1306,In_2512);
nand U1062 (N_1062,In_1329,In_3796);
xnor U1063 (N_1063,In_847,In_2945);
nand U1064 (N_1064,In_3672,In_3578);
nor U1065 (N_1065,In_3467,In_3792);
or U1066 (N_1066,In_4303,In_2527);
and U1067 (N_1067,In_3324,In_53);
nor U1068 (N_1068,In_3782,In_2664);
and U1069 (N_1069,In_3449,In_4474);
nor U1070 (N_1070,In_3060,In_1966);
nor U1071 (N_1071,In_4861,In_1836);
nor U1072 (N_1072,In_4178,In_3773);
or U1073 (N_1073,In_3651,In_808);
and U1074 (N_1074,In_1037,In_1443);
xor U1075 (N_1075,In_363,In_2276);
xnor U1076 (N_1076,In_2330,In_612);
nor U1077 (N_1077,In_2058,In_195);
and U1078 (N_1078,In_3514,In_1796);
nand U1079 (N_1079,In_4170,In_4956);
and U1080 (N_1080,In_1320,In_4837);
nand U1081 (N_1081,In_3127,In_3066);
or U1082 (N_1082,In_1840,In_3439);
xor U1083 (N_1083,In_2855,In_3705);
nand U1084 (N_1084,In_1747,In_1156);
nor U1085 (N_1085,In_2497,In_439);
and U1086 (N_1086,In_4976,In_334);
xnor U1087 (N_1087,In_754,In_4880);
xnor U1088 (N_1088,In_1091,In_3306);
nand U1089 (N_1089,In_4969,In_2410);
nand U1090 (N_1090,In_4552,In_2886);
nand U1091 (N_1091,In_1849,In_1048);
nand U1092 (N_1092,In_181,In_2704);
xnor U1093 (N_1093,In_2343,In_4081);
nor U1094 (N_1094,In_3178,In_3618);
or U1095 (N_1095,In_3121,In_1463);
nor U1096 (N_1096,In_3088,In_3894);
xnor U1097 (N_1097,In_1698,In_460);
xnor U1098 (N_1098,In_2271,In_2742);
nand U1099 (N_1099,In_2408,In_1089);
nor U1100 (N_1100,In_366,In_928);
nand U1101 (N_1101,In_628,In_4387);
or U1102 (N_1102,In_3010,In_4436);
nor U1103 (N_1103,In_2097,In_3756);
nand U1104 (N_1104,In_3008,In_2934);
or U1105 (N_1105,In_2739,In_3711);
xnor U1106 (N_1106,In_2200,In_828);
nor U1107 (N_1107,In_490,In_3952);
or U1108 (N_1108,In_4462,In_4938);
or U1109 (N_1109,In_4586,In_3119);
and U1110 (N_1110,In_2051,In_1984);
xor U1111 (N_1111,In_1069,In_1469);
nor U1112 (N_1112,In_2357,In_1647);
xnor U1113 (N_1113,In_602,In_3348);
nand U1114 (N_1114,In_278,In_4062);
xnor U1115 (N_1115,In_3706,In_1128);
xnor U1116 (N_1116,In_2728,In_2412);
xor U1117 (N_1117,In_4518,In_3307);
nor U1118 (N_1118,In_3250,In_222);
and U1119 (N_1119,In_3543,In_2755);
or U1120 (N_1120,In_1979,In_3053);
xor U1121 (N_1121,In_3240,In_2912);
xnor U1122 (N_1122,In_1548,In_4459);
nor U1123 (N_1123,In_1259,In_4340);
or U1124 (N_1124,In_4084,In_3801);
xor U1125 (N_1125,In_3492,In_2699);
nor U1126 (N_1126,In_432,In_3976);
nor U1127 (N_1127,In_2014,In_3266);
xor U1128 (N_1128,In_4227,In_1652);
xnor U1129 (N_1129,In_2769,In_2333);
nor U1130 (N_1130,In_3964,In_80);
and U1131 (N_1131,In_3105,In_3404);
or U1132 (N_1132,In_1906,In_4200);
nand U1133 (N_1133,In_2620,In_2254);
or U1134 (N_1134,In_653,In_1675);
and U1135 (N_1135,In_1038,In_4181);
xnor U1136 (N_1136,In_1468,In_1153);
nor U1137 (N_1137,In_2637,In_3029);
nor U1138 (N_1138,In_4572,In_2955);
nand U1139 (N_1139,In_1426,In_3344);
and U1140 (N_1140,In_241,In_4820);
or U1141 (N_1141,In_4713,In_1761);
xor U1142 (N_1142,In_1512,In_1342);
or U1143 (N_1143,In_4360,In_1164);
and U1144 (N_1144,In_4410,In_250);
nand U1145 (N_1145,In_1604,In_4583);
nand U1146 (N_1146,In_452,In_2151);
and U1147 (N_1147,In_2295,In_2422);
or U1148 (N_1148,In_198,In_3326);
nor U1149 (N_1149,In_1180,In_570);
xor U1150 (N_1150,In_4751,In_1633);
or U1151 (N_1151,In_4040,In_4356);
and U1152 (N_1152,In_1343,In_745);
xor U1153 (N_1153,In_3091,In_3030);
or U1154 (N_1154,In_3877,In_4033);
and U1155 (N_1155,In_710,In_281);
xnor U1156 (N_1156,In_4221,In_1863);
or U1157 (N_1157,In_3849,In_2456);
nand U1158 (N_1158,In_763,In_3612);
and U1159 (N_1159,In_2329,In_3770);
nand U1160 (N_1160,In_3089,In_1513);
nor U1161 (N_1161,In_3390,In_833);
nor U1162 (N_1162,In_1030,In_2947);
nand U1163 (N_1163,In_3123,In_2465);
or U1164 (N_1164,In_4235,In_2921);
nor U1165 (N_1165,In_1471,In_3056);
nor U1166 (N_1166,In_4904,In_1664);
and U1167 (N_1167,In_47,In_2319);
nor U1168 (N_1168,In_4418,In_2053);
and U1169 (N_1169,In_2849,In_2579);
or U1170 (N_1170,In_3511,In_598);
nand U1171 (N_1171,In_2105,In_4343);
xnor U1172 (N_1172,In_1965,In_688);
xnor U1173 (N_1173,In_4374,In_4799);
xnor U1174 (N_1174,In_3769,In_3936);
nor U1175 (N_1175,In_856,In_2364);
nor U1176 (N_1176,In_3785,In_1348);
and U1177 (N_1177,In_1562,In_2116);
nor U1178 (N_1178,In_2757,In_1474);
or U1179 (N_1179,In_3281,In_4722);
xnor U1180 (N_1180,In_2180,In_3434);
xor U1181 (N_1181,In_2272,In_1318);
nor U1182 (N_1182,In_2542,In_979);
nand U1183 (N_1183,In_1505,In_1537);
nand U1184 (N_1184,In_1976,In_749);
xnor U1185 (N_1185,In_2387,In_2170);
or U1186 (N_1186,In_1286,In_142);
xor U1187 (N_1187,In_3923,In_4382);
nand U1188 (N_1188,In_2601,In_1255);
xnor U1189 (N_1189,In_3365,In_639);
and U1190 (N_1190,In_4400,In_644);
and U1191 (N_1191,In_4645,In_1923);
or U1192 (N_1192,In_4977,In_1080);
nor U1193 (N_1193,In_4974,In_641);
nor U1194 (N_1194,In_2475,In_2594);
xnor U1195 (N_1195,In_3646,In_1040);
nor U1196 (N_1196,In_1755,In_965);
nor U1197 (N_1197,In_4899,In_3860);
and U1198 (N_1198,In_4918,In_4791);
nor U1199 (N_1199,In_1023,In_3289);
nor U1200 (N_1200,In_4502,In_494);
nand U1201 (N_1201,In_78,In_4873);
or U1202 (N_1202,In_3478,In_4071);
or U1203 (N_1203,In_1811,In_1011);
xnor U1204 (N_1204,In_295,In_925);
nand U1205 (N_1205,In_3162,In_3336);
nand U1206 (N_1206,In_1509,In_3779);
nand U1207 (N_1207,In_2466,In_2662);
nand U1208 (N_1208,In_718,In_476);
xor U1209 (N_1209,In_1113,In_4355);
xnor U1210 (N_1210,In_3640,In_785);
xnor U1211 (N_1211,In_2018,In_2351);
nor U1212 (N_1212,In_4002,In_3475);
or U1213 (N_1213,In_1435,In_2367);
nor U1214 (N_1214,In_3798,In_2856);
and U1215 (N_1215,In_1402,In_4038);
xnor U1216 (N_1216,In_1238,In_1857);
and U1217 (N_1217,In_3621,In_3824);
nor U1218 (N_1218,In_4125,In_3681);
and U1219 (N_1219,In_2230,In_2419);
and U1220 (N_1220,In_789,In_1491);
or U1221 (N_1221,In_246,In_2673);
or U1222 (N_1222,In_3810,In_2535);
nand U1223 (N_1223,In_477,In_3200);
xnor U1224 (N_1224,In_4574,In_1630);
and U1225 (N_1225,In_4926,In_336);
nor U1226 (N_1226,In_1262,In_196);
and U1227 (N_1227,In_229,In_1379);
nor U1228 (N_1228,In_4368,In_3826);
or U1229 (N_1229,In_3680,In_1383);
or U1230 (N_1230,In_2382,In_3349);
nor U1231 (N_1231,In_4812,In_4871);
xor U1232 (N_1232,In_2971,In_2084);
and U1233 (N_1233,In_3737,In_4046);
nor U1234 (N_1234,In_3812,In_990);
nand U1235 (N_1235,In_82,In_2414);
and U1236 (N_1236,In_365,In_4726);
xnor U1237 (N_1237,In_4006,In_2817);
nand U1238 (N_1238,In_200,In_750);
nor U1239 (N_1239,In_1937,In_4993);
xor U1240 (N_1240,In_981,In_1355);
xor U1241 (N_1241,In_4633,In_3562);
nand U1242 (N_1242,In_573,In_79);
or U1243 (N_1243,In_915,In_4888);
and U1244 (N_1244,In_24,In_2676);
or U1245 (N_1245,In_2995,In_2539);
or U1246 (N_1246,In_974,In_3963);
xor U1247 (N_1247,In_1397,In_683);
nand U1248 (N_1248,In_2493,In_1007);
nand U1249 (N_1249,In_2303,In_4924);
or U1250 (N_1250,In_2284,In_3335);
nor U1251 (N_1251,In_4719,In_1482);
nor U1252 (N_1252,In_4644,In_1948);
nor U1253 (N_1253,In_1621,In_4715);
nand U1254 (N_1254,In_3120,In_1273);
or U1255 (N_1255,In_1253,In_1955);
xnor U1256 (N_1256,In_3448,In_1200);
or U1257 (N_1257,In_189,In_1689);
or U1258 (N_1258,In_4359,In_4275);
or U1259 (N_1259,In_1341,In_1542);
and U1260 (N_1260,In_1014,In_2211);
and U1261 (N_1261,In_3997,In_1225);
nand U1262 (N_1262,In_2379,In_33);
xnor U1263 (N_1263,In_1834,In_234);
nand U1264 (N_1264,In_1209,In_3062);
nor U1265 (N_1265,In_4835,In_2234);
nor U1266 (N_1266,In_4565,In_390);
nand U1267 (N_1267,In_1850,In_3236);
and U1268 (N_1268,In_4987,In_4744);
or U1269 (N_1269,In_386,In_969);
nand U1270 (N_1270,In_2206,In_2047);
nor U1271 (N_1271,In_3588,In_3708);
or U1272 (N_1272,In_3962,In_1804);
and U1273 (N_1273,In_1666,In_2660);
nor U1274 (N_1274,In_2868,In_2809);
and U1275 (N_1275,In_2726,In_2564);
and U1276 (N_1276,In_579,In_1701);
or U1277 (N_1277,In_4320,In_427);
or U1278 (N_1278,In_2024,In_3871);
nor U1279 (N_1279,In_955,In_385);
or U1280 (N_1280,In_3781,In_3012);
or U1281 (N_1281,In_1479,In_1619);
or U1282 (N_1282,In_1330,In_4985);
nand U1283 (N_1283,In_3715,In_3202);
xor U1284 (N_1284,In_3396,In_4270);
and U1285 (N_1285,In_1016,In_128);
or U1286 (N_1286,In_1293,In_3554);
nand U1287 (N_1287,In_2258,In_1185);
nand U1288 (N_1288,In_3838,In_4720);
xor U1289 (N_1289,In_89,In_4930);
xor U1290 (N_1290,In_692,In_4102);
or U1291 (N_1291,In_1612,In_4507);
nor U1292 (N_1292,In_1584,In_993);
xor U1293 (N_1293,In_3579,In_1390);
or U1294 (N_1294,In_1024,In_3662);
and U1295 (N_1295,In_398,In_4911);
nor U1296 (N_1296,In_3876,In_11);
and U1297 (N_1297,In_2993,In_961);
nand U1298 (N_1298,In_513,In_853);
nor U1299 (N_1299,In_3293,In_3580);
nor U1300 (N_1300,In_2199,In_3516);
nor U1301 (N_1301,In_850,In_1891);
or U1302 (N_1302,In_1697,In_3208);
nor U1303 (N_1303,In_1409,In_551);
nor U1304 (N_1304,In_1888,In_1064);
and U1305 (N_1305,In_361,In_2525);
or U1306 (N_1306,In_4663,In_3193);
or U1307 (N_1307,In_3790,In_2627);
nor U1308 (N_1308,In_3191,In_2184);
xor U1309 (N_1309,In_3624,In_597);
or U1310 (N_1310,In_2296,In_2602);
and U1311 (N_1311,In_873,In_2502);
xnor U1312 (N_1312,In_4403,In_4965);
or U1313 (N_1313,In_1437,In_3984);
and U1314 (N_1314,In_1549,In_2079);
nor U1315 (N_1315,In_1650,In_4115);
xor U1316 (N_1316,In_4833,In_2646);
xnor U1317 (N_1317,In_420,In_1265);
nor U1318 (N_1318,In_1777,In_3795);
and U1319 (N_1319,In_1356,In_3713);
nor U1320 (N_1320,In_4854,In_124);
nor U1321 (N_1321,In_4748,In_1724);
and U1322 (N_1322,In_3880,In_3878);
or U1323 (N_1323,In_3134,In_4379);
or U1324 (N_1324,In_1183,In_353);
and U1325 (N_1325,In_1894,In_1119);
or U1326 (N_1326,In_4723,In_435);
and U1327 (N_1327,In_651,In_3090);
nand U1328 (N_1328,In_4111,In_2135);
or U1329 (N_1329,In_2336,In_1580);
xor U1330 (N_1330,In_4032,In_3656);
or U1331 (N_1331,In_2160,In_3148);
or U1332 (N_1332,In_2834,In_4596);
nor U1333 (N_1333,In_2378,In_846);
nor U1334 (N_1334,In_2370,In_3730);
and U1335 (N_1335,In_4401,In_2036);
or U1336 (N_1336,In_1536,In_3345);
nor U1337 (N_1337,In_2215,In_721);
xnor U1338 (N_1338,In_3351,In_3233);
xor U1339 (N_1339,In_1234,In_3169);
or U1340 (N_1340,In_188,In_3116);
and U1341 (N_1341,In_4305,In_2106);
xnor U1342 (N_1342,In_3949,In_2778);
nor U1343 (N_1343,In_4097,In_2648);
xnor U1344 (N_1344,In_3728,In_735);
nand U1345 (N_1345,In_2867,In_4430);
nor U1346 (N_1346,In_4794,In_3025);
or U1347 (N_1347,In_10,In_2847);
or U1348 (N_1348,In_2468,In_1735);
nor U1349 (N_1349,In_3311,In_1494);
or U1350 (N_1350,In_4480,In_577);
xor U1351 (N_1351,In_3057,In_4600);
xnor U1352 (N_1352,In_960,In_3480);
and U1353 (N_1353,In_4096,In_2376);
nand U1354 (N_1354,In_3977,In_2499);
nand U1355 (N_1355,In_3229,In_2963);
nand U1356 (N_1356,In_772,In_100);
or U1357 (N_1357,In_41,In_741);
and U1358 (N_1358,In_538,In_1245);
and U1359 (N_1359,In_4559,In_1718);
nand U1360 (N_1360,In_4967,In_2195);
nand U1361 (N_1361,In_4702,In_206);
and U1362 (N_1362,In_104,In_994);
nand U1363 (N_1363,In_4624,In_2063);
or U1364 (N_1364,In_4788,In_2259);
nand U1365 (N_1365,In_1359,In_2666);
or U1366 (N_1366,In_2721,In_4773);
and U1367 (N_1367,In_2920,In_4262);
and U1368 (N_1368,In_615,In_51);
nand U1369 (N_1369,In_797,In_1022);
nand U1370 (N_1370,In_4630,In_169);
and U1371 (N_1371,In_2349,In_1250);
nor U1372 (N_1372,In_4256,In_1569);
or U1373 (N_1373,In_1060,In_1541);
or U1374 (N_1374,In_811,In_3273);
and U1375 (N_1375,In_3111,In_3983);
xnor U1376 (N_1376,In_3584,In_3430);
or U1377 (N_1377,In_1264,In_2126);
nand U1378 (N_1378,In_3564,In_1454);
xor U1379 (N_1379,In_663,In_2022);
and U1380 (N_1380,In_3825,In_2049);
xnor U1381 (N_1381,In_3277,In_1366);
xor U1382 (N_1382,In_3313,In_838);
or U1383 (N_1383,In_146,In_3758);
and U1384 (N_1384,In_3693,In_2967);
nor U1385 (N_1385,In_2239,In_4416);
xor U1386 (N_1386,In_4105,In_1485);
and U1387 (N_1387,In_3260,In_1056);
nand U1388 (N_1388,In_4488,In_4328);
nand U1389 (N_1389,In_2147,In_1795);
and U1390 (N_1390,In_1260,In_1195);
nor U1391 (N_1391,In_4534,In_4330);
xor U1392 (N_1392,In_4165,In_2590);
nand U1393 (N_1393,In_3331,In_1239);
nand U1394 (N_1394,In_1169,In_3104);
and U1395 (N_1395,In_4492,In_4839);
or U1396 (N_1396,In_2122,In_1731);
xnor U1397 (N_1397,In_419,In_4875);
and U1398 (N_1398,In_4151,In_1821);
or U1399 (N_1399,In_2040,In_1712);
nand U1400 (N_1400,In_1221,In_154);
xnor U1401 (N_1401,In_190,In_4371);
and U1402 (N_1402,In_620,In_3908);
xnor U1403 (N_1403,In_1606,In_3242);
xor U1404 (N_1404,In_1875,In_4187);
nor U1405 (N_1405,In_4942,In_1561);
nand U1406 (N_1406,In_1560,In_4202);
nor U1407 (N_1407,In_4566,In_813);
nand U1408 (N_1408,In_199,In_627);
nand U1409 (N_1409,In_4817,In_566);
or U1410 (N_1410,In_4335,In_2644);
xnor U1411 (N_1411,In_133,In_4107);
or U1412 (N_1412,In_2353,In_4893);
and U1413 (N_1413,In_1851,In_2334);
nand U1414 (N_1414,In_4411,In_775);
or U1415 (N_1415,In_4512,In_4798);
nand U1416 (N_1416,In_4619,In_1457);
or U1417 (N_1417,In_471,In_4405);
nor U1418 (N_1418,In_3408,In_948);
xnor U1419 (N_1419,In_4822,In_4792);
and U1420 (N_1420,In_3182,In_4086);
nand U1421 (N_1421,In_4129,In_3848);
or U1422 (N_1422,In_1378,In_3379);
nand U1423 (N_1423,In_4614,In_86);
nor U1424 (N_1424,In_4528,In_3731);
nor U1425 (N_1425,In_355,In_2087);
nor U1426 (N_1426,In_1097,In_695);
xor U1427 (N_1427,In_3417,In_4239);
nor U1428 (N_1428,In_2861,In_3466);
and U1429 (N_1429,In_3925,In_978);
or U1430 (N_1430,In_0,In_2567);
nand U1431 (N_1431,In_176,In_1919);
xnor U1432 (N_1432,In_2399,In_1787);
nand U1433 (N_1433,In_4923,In_4953);
nand U1434 (N_1434,In_2557,In_413);
xor U1435 (N_1435,In_4864,In_2832);
and U1436 (N_1436,In_3143,In_2768);
or U1437 (N_1437,In_843,In_1099);
and U1438 (N_1438,In_3702,In_687);
or U1439 (N_1439,In_131,In_2640);
xor U1440 (N_1440,In_2857,In_1555);
and U1441 (N_1441,In_367,In_1400);
xor U1442 (N_1442,In_1695,In_202);
nor U1443 (N_1443,In_1310,In_2919);
nor U1444 (N_1444,In_2903,In_4986);
nand U1445 (N_1445,In_1261,In_2973);
xnor U1446 (N_1446,In_4598,In_3870);
or U1447 (N_1447,In_613,In_3980);
and U1448 (N_1448,In_4350,In_507);
nand U1449 (N_1449,In_4962,In_2451);
nor U1450 (N_1450,In_4362,In_4920);
or U1451 (N_1451,In_4172,In_2121);
or U1452 (N_1452,In_174,In_3381);
xnor U1453 (N_1453,In_2071,In_984);
xor U1454 (N_1454,In_2634,In_2085);
or U1455 (N_1455,In_410,In_495);
and U1456 (N_1456,In_3149,In_177);
and U1457 (N_1457,In_2740,In_1627);
or U1458 (N_1458,In_3158,In_2375);
nor U1459 (N_1459,In_1116,In_3226);
or U1460 (N_1460,In_2827,In_1106);
nand U1461 (N_1461,In_3591,In_445);
or U1462 (N_1462,In_1628,In_2799);
xnor U1463 (N_1463,In_3083,In_1887);
nand U1464 (N_1464,In_4514,In_2772);
nor U1465 (N_1465,In_1962,In_4620);
nand U1466 (N_1466,In_3165,In_3934);
and U1467 (N_1467,In_2445,In_4576);
and U1468 (N_1468,In_93,In_1631);
nor U1469 (N_1469,In_1003,In_1766);
and U1470 (N_1470,In_3791,In_328);
xor U1471 (N_1471,In_1287,In_3710);
nand U1472 (N_1472,In_55,In_3214);
and U1473 (N_1473,In_4175,In_3902);
or U1474 (N_1474,In_1574,In_2584);
nand U1475 (N_1475,In_401,In_3429);
or U1476 (N_1476,In_4466,In_3405);
nand U1477 (N_1477,In_106,In_975);
xnor U1478 (N_1478,In_4916,In_1601);
nand U1479 (N_1479,In_77,In_1311);
nand U1480 (N_1480,In_227,In_562);
xor U1481 (N_1481,In_2944,In_2506);
or U1482 (N_1482,In_4351,In_444);
nand U1483 (N_1483,In_3907,In_1540);
xnor U1484 (N_1484,In_3176,In_4094);
and U1485 (N_1485,In_563,In_596);
nor U1486 (N_1486,In_2452,In_2143);
or U1487 (N_1487,In_3406,In_4755);
or U1488 (N_1488,In_3698,In_4831);
and U1489 (N_1489,In_2123,In_3751);
nor U1490 (N_1490,In_1074,In_4388);
nand U1491 (N_1491,In_796,In_2113);
xnor U1492 (N_1492,In_4279,In_1639);
and U1493 (N_1493,In_4315,In_483);
nor U1494 (N_1494,In_4671,In_3501);
or U1495 (N_1495,In_447,In_300);
nand U1496 (N_1496,In_4800,In_4277);
and U1497 (N_1497,In_3978,In_670);
nor U1498 (N_1498,In_4778,In_2672);
nand U1499 (N_1499,In_4482,In_4404);
nor U1500 (N_1500,In_2163,In_2630);
nor U1501 (N_1501,In_2798,In_4971);
nand U1502 (N_1502,In_4498,In_521);
xor U1503 (N_1503,In_3222,In_2119);
nand U1504 (N_1504,In_2968,In_3196);
xnor U1505 (N_1505,In_2547,In_4449);
or U1506 (N_1506,In_4603,In_2836);
or U1507 (N_1507,In_3205,In_2305);
and U1508 (N_1508,In_2098,In_3891);
and U1509 (N_1509,In_1878,In_2377);
xor U1510 (N_1510,In_4959,In_1980);
nor U1511 (N_1511,In_1492,In_4921);
nand U1512 (N_1512,In_4114,In_2889);
nand U1513 (N_1513,In_2568,In_359);
nand U1514 (N_1514,In_3999,In_1602);
nor U1515 (N_1515,In_340,In_1971);
nand U1516 (N_1516,In_4769,In_3228);
nor U1517 (N_1517,In_4278,In_3549);
and U1518 (N_1518,In_1521,In_4442);
xnor U1519 (N_1519,In_2346,In_4234);
nand U1520 (N_1520,In_3973,In_3951);
nand U1521 (N_1521,In_482,In_1528);
nor U1522 (N_1522,In_1780,In_1105);
nor U1523 (N_1523,In_1883,In_160);
nor U1524 (N_1524,In_1903,In_4426);
and U1525 (N_1525,In_1459,In_542);
nor U1526 (N_1526,In_4425,In_865);
or U1527 (N_1527,In_2624,In_3437);
or U1528 (N_1528,In_3945,In_2604);
nor U1529 (N_1529,In_2718,In_3015);
and U1530 (N_1530,In_2144,In_391);
and U1531 (N_1531,In_4615,In_3038);
nand U1532 (N_1532,In_2876,In_1703);
nor U1533 (N_1533,In_3401,In_3361);
nor U1534 (N_1534,In_3729,In_578);
nand U1535 (N_1535,In_1945,In_520);
nand U1536 (N_1536,In_4961,In_3253);
nor U1537 (N_1537,In_681,In_2498);
and U1538 (N_1538,In_1547,In_3426);
or U1539 (N_1539,In_69,In_829);
or U1540 (N_1540,In_1996,In_2423);
and U1541 (N_1541,In_3276,In_4274);
nor U1542 (N_1542,In_2268,In_4237);
nor U1543 (N_1543,In_3623,In_1144);
nand U1544 (N_1544,In_803,In_708);
nor U1545 (N_1545,In_312,In_4154);
nand U1546 (N_1546,In_4285,In_4447);
xor U1547 (N_1547,In_4531,In_2048);
and U1548 (N_1548,In_2459,In_776);
or U1549 (N_1549,In_381,In_1495);
and U1550 (N_1550,In_526,In_3626);
and U1551 (N_1551,In_3524,In_2583);
nor U1552 (N_1552,In_2813,In_2753);
nor U1553 (N_1553,In_4431,In_3050);
nor U1554 (N_1554,In_2312,In_498);
and U1555 (N_1555,In_1357,In_3298);
and U1556 (N_1556,In_781,In_3468);
nand U1557 (N_1557,In_4361,In_851);
and U1558 (N_1558,In_1408,In_1590);
or U1559 (N_1559,In_3603,In_988);
and U1560 (N_1560,In_2020,In_2074);
nand U1561 (N_1561,In_4067,In_3868);
and U1562 (N_1562,In_4284,In_3509);
nor U1563 (N_1563,In_4041,In_1372);
xor U1564 (N_1564,In_3073,In_3803);
and U1565 (N_1565,In_4109,In_3075);
or U1566 (N_1566,In_3555,In_4201);
nand U1567 (N_1567,In_3961,In_4746);
nor U1568 (N_1568,In_736,In_3221);
and U1569 (N_1569,In_1940,In_3440);
nand U1570 (N_1570,In_85,In_1752);
nand U1571 (N_1571,In_2508,In_3432);
and U1572 (N_1572,In_2766,In_3239);
and U1573 (N_1573,In_1018,In_1405);
and U1574 (N_1574,In_1824,In_3338);
nor U1575 (N_1575,In_4222,In_820);
nand U1576 (N_1576,In_1623,In_4271);
or U1577 (N_1577,In_3552,In_731);
nand U1578 (N_1578,In_4643,In_3035);
or U1579 (N_1579,In_1629,In_35);
nor U1580 (N_1580,In_3263,In_2342);
and U1581 (N_1581,In_1660,In_4529);
and U1582 (N_1582,In_760,In_322);
or U1583 (N_1583,In_2893,In_1769);
nand U1584 (N_1584,In_211,In_2658);
xor U1585 (N_1585,In_3037,In_3633);
and U1586 (N_1586,In_3371,In_4059);
nand U1587 (N_1587,In_4678,In_2744);
or U1588 (N_1588,In_630,In_589);
nand U1589 (N_1589,In_3268,In_964);
nand U1590 (N_1590,In_1477,In_3246);
or U1591 (N_1591,In_1764,In_2706);
or U1592 (N_1592,In_966,In_2686);
nand U1593 (N_1593,In_3427,In_2128);
nand U1594 (N_1594,In_3675,In_2708);
and U1595 (N_1595,In_2915,In_1992);
or U1596 (N_1596,In_1905,In_3513);
nand U1597 (N_1597,In_2015,In_4573);
nor U1598 (N_1598,In_4902,In_4302);
nor U1599 (N_1599,In_3687,In_3507);
and U1600 (N_1600,In_3356,In_1938);
or U1601 (N_1601,In_4376,In_3206);
xnor U1602 (N_1602,In_1526,In_2403);
xnor U1603 (N_1603,In_4232,In_528);
nor U1604 (N_1604,In_1139,In_4901);
or U1605 (N_1605,In_4236,In_468);
and U1606 (N_1606,In_2059,In_4592);
xnor U1607 (N_1607,In_1588,In_165);
nor U1608 (N_1608,In_4313,In_953);
and U1609 (N_1609,In_3628,In_87);
nand U1610 (N_1610,In_239,In_3186);
nor U1611 (N_1611,In_2472,In_3942);
nor U1612 (N_1612,In_3382,In_1256);
nor U1613 (N_1613,In_4760,In_2898);
nor U1614 (N_1614,In_409,In_3593);
and U1615 (N_1615,In_4509,In_2325);
or U1616 (N_1616,In_3359,In_756);
xnor U1617 (N_1617,In_1297,In_1033);
nand U1618 (N_1618,In_1611,In_4732);
xnor U1619 (N_1619,In_2747,In_998);
and U1620 (N_1620,In_3300,In_4180);
nand U1621 (N_1621,In_4146,In_4551);
or U1622 (N_1622,In_505,In_2960);
nor U1623 (N_1623,In_168,In_1815);
and U1624 (N_1624,In_416,In_256);
nand U1625 (N_1625,In_545,In_905);
nor U1626 (N_1626,In_4247,In_832);
nor U1627 (N_1627,In_1649,In_4100);
or U1628 (N_1628,In_4869,In_804);
nand U1629 (N_1629,In_2884,In_4099);
nand U1630 (N_1630,In_1452,In_2685);
nor U1631 (N_1631,In_632,In_2607);
nor U1632 (N_1632,In_2759,In_4157);
xor U1633 (N_1633,In_2917,In_4968);
nor U1634 (N_1634,In_2693,In_4990);
nand U1635 (N_1635,In_3989,In_4634);
nor U1636 (N_1636,In_2659,In_2226);
and U1637 (N_1637,In_4690,In_3674);
or U1638 (N_1638,In_1829,In_2124);
nor U1639 (N_1639,In_217,In_2314);
xnor U1640 (N_1640,In_4316,In_1866);
nor U1641 (N_1641,In_4753,In_700);
nand U1642 (N_1642,In_3547,In_852);
nand U1643 (N_1643,In_1750,In_1136);
nand U1644 (N_1644,In_4686,In_1596);
xnor U1645 (N_1645,In_1858,In_3380);
xnor U1646 (N_1646,In_306,In_2710);
and U1647 (N_1647,In_3644,In_3581);
and U1648 (N_1648,In_4855,In_918);
nor U1649 (N_1649,In_4681,In_65);
nand U1650 (N_1650,In_1872,In_4952);
and U1651 (N_1651,In_2534,In_4495);
nand U1652 (N_1652,In_3515,In_4419);
nor U1653 (N_1653,In_590,In_2814);
nand U1654 (N_1654,In_3301,In_2192);
nand U1655 (N_1655,In_884,In_3157);
nand U1656 (N_1656,In_2107,In_3201);
and U1657 (N_1657,In_4949,In_2951);
and U1658 (N_1658,In_4745,In_2900);
and U1659 (N_1659,In_459,In_4979);
and U1660 (N_1660,In_179,In_1012);
and U1661 (N_1661,In_1897,In_693);
nand U1662 (N_1662,In_1466,In_45);
or U1663 (N_1663,In_4541,In_1706);
or U1664 (N_1664,In_2816,In_4765);
xor U1665 (N_1665,In_230,In_2899);
xor U1666 (N_1666,In_3055,In_938);
nor U1667 (N_1667,In_4152,In_1448);
nor U1668 (N_1668,In_3979,In_2674);
and U1669 (N_1669,In_116,In_2713);
and U1670 (N_1670,In_901,In_1716);
or U1671 (N_1671,In_2791,In_4849);
nor U1672 (N_1672,In_193,In_2518);
xnor U1673 (N_1673,In_1005,In_4016);
xnor U1674 (N_1674,In_3736,In_423);
and U1675 (N_1675,In_595,In_908);
nor U1676 (N_1676,In_2481,In_166);
nor U1677 (N_1677,In_4803,In_2933);
nand U1678 (N_1678,In_2948,In_720);
and U1679 (N_1679,In_4420,In_2697);
xnor U1680 (N_1680,In_4257,In_3265);
xor U1681 (N_1681,In_4021,In_2411);
and U1682 (N_1682,In_2569,In_1792);
nand U1683 (N_1683,In_426,In_2070);
nor U1684 (N_1684,In_919,In_3742);
nand U1685 (N_1685,In_4905,In_555);
nor U1686 (N_1686,In_2263,In_3858);
or U1687 (N_1687,In_2783,In_2007);
nand U1688 (N_1688,In_1736,In_1475);
nor U1689 (N_1689,In_2838,In_2374);
nor U1690 (N_1690,In_1323,In_4876);
nor U1691 (N_1691,In_1904,In_2241);
nor U1692 (N_1692,In_2807,In_2311);
or U1693 (N_1693,In_1552,In_4821);
or U1694 (N_1694,In_574,In_2300);
nor U1695 (N_1695,In_99,In_2196);
nor U1696 (N_1696,In_1659,In_400);
nand U1697 (N_1697,In_324,In_2103);
xnor U1698 (N_1698,In_1363,In_4448);
nand U1699 (N_1699,In_407,In_3031);
xor U1700 (N_1700,In_1241,In_716);
nor U1701 (N_1701,In_2553,In_2885);
xnor U1702 (N_1702,In_4244,In_2599);
nand U1703 (N_1703,In_2785,In_4363);
xnor U1704 (N_1704,In_1460,In_3539);
xnor U1705 (N_1705,In_3529,In_1497);
xnor U1706 (N_1706,In_130,In_4050);
and U1707 (N_1707,In_958,In_2146);
nor U1708 (N_1708,In_1710,In_3958);
or U1709 (N_1709,In_4525,In_3776);
or U1710 (N_1710,In_3678,In_2575);
xnor U1711 (N_1711,In_4752,In_4392);
or U1712 (N_1712,In_4548,In_3100);
and U1713 (N_1713,In_1714,In_4211);
nor U1714 (N_1714,In_4128,In_4537);
or U1715 (N_1715,In_4186,In_1553);
nor U1716 (N_1716,In_1313,In_3339);
and U1717 (N_1717,In_1554,In_3267);
or U1718 (N_1718,In_3582,In_3535);
and U1719 (N_1719,In_3252,In_244);
and U1720 (N_1720,In_276,In_266);
nand U1721 (N_1721,In_3484,In_3274);
nand U1722 (N_1722,In_4524,In_3130);
and U1723 (N_1723,In_3489,In_4261);
and U1724 (N_1724,In_4399,In_672);
or U1725 (N_1725,In_2763,In_4093);
xor U1726 (N_1726,In_4859,In_814);
nor U1727 (N_1727,In_976,In_4375);
xnor U1728 (N_1728,In_891,In_1846);
nor U1729 (N_1729,In_3719,In_2794);
or U1730 (N_1730,In_4127,In_4123);
nor U1731 (N_1731,In_4660,In_4331);
or U1732 (N_1732,In_3689,In_2294);
and U1733 (N_1733,In_52,In_1171);
nor U1734 (N_1734,In_3910,In_1223);
and U1735 (N_1735,In_14,In_902);
or U1736 (N_1736,In_903,In_1839);
xnor U1737 (N_1737,In_4648,In_2571);
nand U1738 (N_1738,In_309,In_3823);
or U1739 (N_1739,In_1188,In_2463);
nand U1740 (N_1740,In_1518,In_3465);
xnor U1741 (N_1741,In_3309,In_648);
or U1742 (N_1742,In_911,In_607);
and U1743 (N_1743,In_1531,In_913);
xor U1744 (N_1744,In_1276,In_3590);
or U1745 (N_1745,In_2850,In_3808);
nand U1746 (N_1746,In_855,In_2416);
and U1747 (N_1747,In_3407,In_1832);
xnor U1748 (N_1748,In_1149,In_3244);
and U1749 (N_1749,In_4567,In_2293);
and U1750 (N_1750,In_2770,In_4545);
or U1751 (N_1751,In_4026,In_2026);
nor U1752 (N_1752,In_4868,In_4453);
nand U1753 (N_1753,In_1288,In_4413);
nand U1754 (N_1754,In_1065,In_1281);
or U1755 (N_1755,In_3718,In_4138);
nand U1756 (N_1756,In_43,In_3017);
and U1757 (N_1757,In_3788,In_4255);
nand U1758 (N_1758,In_4394,In_3314);
xnor U1759 (N_1759,In_67,In_3648);
and U1760 (N_1760,In_30,In_660);
xor U1761 (N_1761,In_2681,In_3558);
nand U1762 (N_1762,In_977,In_1614);
nand U1763 (N_1763,In_3412,In_403);
xnor U1764 (N_1764,In_1835,In_4933);
or U1765 (N_1765,In_3789,In_912);
nor U1766 (N_1766,In_3506,In_4024);
or U1767 (N_1767,In_1203,In_145);
nand U1768 (N_1768,In_4223,In_3807);
xor U1769 (N_1769,In_1550,In_2023);
nand U1770 (N_1770,In_271,In_4280);
and U1771 (N_1771,In_2781,In_4804);
nand U1772 (N_1772,In_2185,In_2297);
nor U1773 (N_1773,In_280,In_1322);
nand U1774 (N_1774,In_4267,In_152);
nor U1775 (N_1775,In_3496,In_4242);
nor U1776 (N_1776,In_1734,In_3319);
nor U1777 (N_1777,In_316,In_1092);
xnor U1778 (N_1778,In_2425,In_3571);
or U1779 (N_1779,In_418,In_3732);
and U1780 (N_1780,In_3375,In_1112);
xnor U1781 (N_1781,In_1707,In_3527);
or U1782 (N_1782,In_1215,In_2561);
or U1783 (N_1783,In_870,In_3494);
and U1784 (N_1784,In_1880,In_3294);
and U1785 (N_1785,In_2054,In_4395);
nand U1786 (N_1786,In_4088,In_1978);
nand U1787 (N_1787,In_2301,In_4119);
or U1788 (N_1788,In_618,In_972);
nand U1789 (N_1789,In_2572,In_1447);
and U1790 (N_1790,In_1290,In_4433);
or U1791 (N_1791,In_2682,In_1801);
or U1792 (N_1792,In_4858,In_4148);
xnor U1793 (N_1793,In_491,In_1427);
or U1794 (N_1794,In_1910,In_4185);
nand U1795 (N_1795,In_212,In_2);
nand U1796 (N_1796,In_872,In_1280);
nor U1797 (N_1797,In_2761,In_3630);
or U1798 (N_1798,In_1206,In_2344);
xor U1799 (N_1799,In_3745,In_2543);
xnor U1800 (N_1800,In_4321,In_1126);
nand U1801 (N_1801,In_4358,In_4783);
and U1802 (N_1802,In_379,In_2424);
nand U1803 (N_1803,In_3474,In_2127);
nor U1804 (N_1804,In_2323,In_1952);
and U1805 (N_1805,In_4092,In_3235);
xnor U1806 (N_1806,In_122,In_1017);
nor U1807 (N_1807,In_2661,In_2896);
and U1808 (N_1808,In_942,In_1876);
nor U1809 (N_1809,In_3488,In_2265);
nor U1810 (N_1810,In_3042,In_3570);
or U1811 (N_1811,In_4838,In_4570);
or U1812 (N_1812,In_3636,In_1394);
xnor U1813 (N_1813,In_2436,In_2083);
xnor U1814 (N_1814,In_1929,In_4703);
or U1815 (N_1815,In_2025,In_3386);
and U1816 (N_1816,In_4730,In_438);
nand U1817 (N_1817,In_4054,In_2692);
and U1818 (N_1818,In_4307,In_4922);
nand U1819 (N_1819,In_4254,In_3926);
nor U1820 (N_1820,In_1000,In_4082);
or U1821 (N_1821,In_4698,In_3568);
xor U1822 (N_1822,In_3755,In_2688);
and U1823 (N_1823,In_2073,In_34);
xor U1824 (N_1824,In_1895,In_103);
and U1825 (N_1825,In_3224,In_3605);
and U1826 (N_1826,In_1783,In_1585);
and U1827 (N_1827,In_2937,In_2974);
xnor U1828 (N_1828,In_3840,In_4191);
xnor U1829 (N_1829,In_3703,In_3900);
xor U1830 (N_1830,In_899,In_3967);
nor U1831 (N_1831,In_2983,In_4706);
or U1832 (N_1832,In_610,In_1723);
and U1833 (N_1833,In_4353,In_3317);
nand U1834 (N_1834,In_3132,In_2954);
xor U1835 (N_1835,In_2786,In_4461);
xor U1836 (N_1836,In_1217,In_719);
xnor U1837 (N_1837,In_3106,In_2044);
nand U1838 (N_1838,In_2513,In_3470);
nor U1839 (N_1839,In_2998,In_3223);
nand U1840 (N_1840,In_713,In_547);
xor U1841 (N_1841,In_2874,In_2871);
and U1842 (N_1842,In_291,In_1539);
xnor U1843 (N_1843,In_240,In_1788);
and U1844 (N_1844,In_3086,In_2208);
or U1845 (N_1845,In_1282,In_389);
nor U1846 (N_1846,In_3425,In_137);
nor U1847 (N_1847,In_1545,In_59);
and U1848 (N_1848,In_3931,In_1626);
or U1849 (N_1849,In_3280,In_4768);
or U1850 (N_1850,In_3243,In_1227);
xnor U1851 (N_1851,In_743,In_3834);
nand U1852 (N_1852,In_500,In_2820);
and U1853 (N_1853,In_3385,In_1417);
nor U1854 (N_1854,In_603,In_2848);
xor U1855 (N_1855,In_2695,In_617);
xor U1856 (N_1856,In_149,In_4428);
or U1857 (N_1857,In_3583,In_3082);
and U1858 (N_1858,In_3241,In_564);
or U1859 (N_1859,In_4543,In_3110);
or U1860 (N_1860,In_1884,In_944);
nand U1861 (N_1861,In_1157,In_1972);
xnor U1862 (N_1862,In_2159,In_2012);
nand U1863 (N_1863,In_2331,In_2888);
nand U1864 (N_1864,In_4727,In_1152);
and U1865 (N_1865,In_4874,In_4259);
and U1866 (N_1866,In_2400,In_694);
nand U1867 (N_1867,In_147,In_4208);
xnor U1868 (N_1868,In_4326,In_4230);
nor U1869 (N_1869,In_1049,In_503);
xor U1870 (N_1870,In_2711,In_1763);
or U1871 (N_1871,In_1920,In_3211);
or U1872 (N_1872,In_1968,In_2441);
xnor U1873 (N_1873,In_1021,In_3063);
or U1874 (N_1874,In_4884,In_406);
xor U1875 (N_1875,In_4828,In_1381);
xnor U1876 (N_1876,In_3841,In_450);
nand U1877 (N_1877,In_702,In_39);
nand U1878 (N_1878,In_4554,In_1591);
nand U1879 (N_1879,In_4066,In_3141);
nor U1880 (N_1880,In_3247,In_1989);
or U1881 (N_1881,In_2626,In_3369);
or U1882 (N_1882,In_1068,In_1898);
xnor U1883 (N_1883,In_4705,In_764);
nor U1884 (N_1884,In_2548,In_2453);
and U1885 (N_1885,In_3296,In_1527);
xnor U1886 (N_1886,In_3362,In_1387);
xor U1887 (N_1887,In_3573,In_3400);
or U1888 (N_1888,In_1109,In_1484);
xnor U1889 (N_1889,In_3118,In_4613);
and U1890 (N_1890,In_2385,In_1939);
and U1891 (N_1891,In_4757,In_2879);
or U1892 (N_1892,In_2875,In_2618);
nor U1893 (N_1893,In_3287,In_2298);
nand U1894 (N_1894,In_2129,In_605);
xor U1895 (N_1895,In_1921,In_4579);
xor U1896 (N_1896,In_2691,In_251);
nand U1897 (N_1897,In_92,In_3768);
or U1898 (N_1898,In_2840,In_2238);
or U1899 (N_1899,In_684,In_1034);
nand U1900 (N_1900,In_3418,In_4205);
xor U1901 (N_1901,In_2767,In_1572);
or U1902 (N_1902,In_3318,In_3261);
nand U1903 (N_1903,In_4955,In_4931);
nor U1904 (N_1904,In_4179,In_3291);
nand U1905 (N_1905,In_2952,In_4790);
nand U1906 (N_1906,In_4776,In_50);
nor U1907 (N_1907,In_4759,In_1361);
nand U1908 (N_1908,In_4454,In_2418);
and U1909 (N_1909,In_2521,In_4022);
or U1910 (N_1910,In_261,In_2591);
or U1911 (N_1911,In_1369,In_3839);
xnor U1912 (N_1912,In_895,In_778);
nor U1913 (N_1913,In_3397,In_629);
nor U1914 (N_1914,In_525,In_3275);
or U1915 (N_1915,In_4654,In_1496);
nor U1916 (N_1916,In_868,In_771);
nor U1917 (N_1917,In_2322,In_4912);
xor U1918 (N_1918,In_4970,In_818);
xor U1919 (N_1919,In_2448,In_2932);
nor U1920 (N_1920,In_4564,In_4928);
and U1921 (N_1921,In_1046,In_3218);
xor U1922 (N_1922,In_1374,In_1442);
xor U1923 (N_1923,In_3847,In_3677);
nor U1924 (N_1924,In_3722,In_2540);
nor U1925 (N_1925,In_2273,In_4714);
and U1926 (N_1926,In_3727,In_3343);
xnor U1927 (N_1927,In_4658,In_3783);
or U1928 (N_1928,In_550,In_1818);
nand U1929 (N_1929,In_1248,In_2099);
nand U1930 (N_1930,In_2302,In_2663);
or U1931 (N_1931,In_269,In_2670);
and U1932 (N_1932,In_4601,In_4306);
nor U1933 (N_1933,In_2925,In_837);
nand U1934 (N_1934,In_3204,In_809);
or U1935 (N_1935,In_3601,In_455);
and U1936 (N_1936,In_3928,In_864);
nor U1937 (N_1937,In_3433,In_4342);
xnor U1938 (N_1938,In_4517,In_3052);
or U1939 (N_1939,In_941,In_2570);
xor U1940 (N_1940,In_3438,In_690);
nor U1941 (N_1941,In_2943,In_1137);
nand U1942 (N_1942,In_730,In_724);
xor U1943 (N_1943,In_4424,In_3617);
nand U1944 (N_1944,In_4699,In_3254);
and U1945 (N_1945,In_2764,In_3032);
and U1946 (N_1946,In_698,In_1713);
xor U1947 (N_1947,In_1678,In_1645);
nand U1948 (N_1948,In_3883,In_2050);
nand U1949 (N_1949,In_1244,In_1822);
nor U1950 (N_1950,In_2833,In_1767);
nor U1951 (N_1951,In_1008,In_140);
nand U1952 (N_1952,In_2731,In_3647);
and U1953 (N_1953,In_3940,In_1998);
or U1954 (N_1954,In_4293,In_1246);
and U1955 (N_1955,In_1663,In_1191);
or U1956 (N_1956,In_3815,In_691);
nand U1957 (N_1957,In_1354,In_83);
nor U1958 (N_1958,In_3668,In_1222);
xnor U1959 (N_1959,In_3827,In_430);
or U1960 (N_1960,In_1558,In_2999);
and U1961 (N_1961,In_182,In_4747);
and U1962 (N_1962,In_4333,In_4471);
nor U1963 (N_1963,In_4072,In_260);
nor U1964 (N_1964,In_1375,In_4167);
xor U1965 (N_1965,In_2563,In_205);
and U1966 (N_1966,In_1848,In_1219);
nand U1967 (N_1967,In_2537,In_2324);
xor U1968 (N_1968,In_3850,In_962);
xnor U1969 (N_1969,In_4162,In_2656);
nor U1970 (N_1970,In_3664,In_187);
and U1971 (N_1971,In_3321,In_3735);
and U1972 (N_1972,In_2169,In_3395);
nor U1973 (N_1973,In_1271,In_2883);
nor U1974 (N_1974,In_2246,In_3003);
or U1975 (N_1975,In_1166,In_1794);
nor U1976 (N_1976,In_2982,In_1072);
nand U1977 (N_1977,In_425,In_2524);
nor U1978 (N_1978,In_746,In_4143);
nand U1979 (N_1979,In_2005,In_2190);
and U1980 (N_1980,In_4646,In_382);
and U1981 (N_1981,In_3833,In_1797);
or U1982 (N_1982,In_3469,In_2835);
nor U1983 (N_1983,In_2823,In_2426);
nand U1984 (N_1984,In_4213,In_2130);
xnor U1985 (N_1985,In_4220,In_4806);
and U1986 (N_1986,In_2780,In_2021);
nand U1987 (N_1987,In_1254,In_3248);
xor U1988 (N_1988,In_625,In_76);
nand U1989 (N_1989,In_1603,In_4258);
nand U1990 (N_1990,In_1570,In_3652);
or U1991 (N_1991,In_1332,In_4489);
xnor U1992 (N_1992,In_910,In_156);
or U1993 (N_1993,In_3799,In_3904);
and U1994 (N_1994,In_2075,In_1382);
nor U1995 (N_1995,In_2988,In_556);
nor U1996 (N_1996,In_4000,In_2787);
xnor U1997 (N_1997,In_645,In_1853);
and U1998 (N_1998,In_2771,In_1508);
xor U1999 (N_1999,In_25,In_209);
nand U2000 (N_2000,In_2892,In_3217);
xor U2001 (N_2001,In_157,In_4025);
nor U2002 (N_2002,In_567,In_2901);
or U2003 (N_2003,In_3660,In_782);
nand U2004 (N_2004,In_1340,In_2842);
or U2005 (N_2005,In_2447,In_2719);
and U2006 (N_2006,In_1970,In_4581);
xnor U2007 (N_2007,In_1025,In_4250);
and U2008 (N_2008,In_689,In_1449);
and U2009 (N_2009,In_1691,In_4319);
xor U2010 (N_2010,In_831,In_3181);
nor U2011 (N_2011,In_2631,In_807);
nor U2012 (N_2012,In_3837,In_290);
nand U2013 (N_2013,In_3155,In_854);
xnor U2014 (N_2014,In_3255,In_257);
or U2015 (N_2015,In_650,In_3998);
nor U2016 (N_2016,In_1720,In_1075);
nand U2017 (N_2017,In_1845,In_3522);
and U2018 (N_2018,In_4815,In_218);
nand U2019 (N_2019,In_4700,In_2812);
nor U2020 (N_2020,In_134,In_2536);
nor U2021 (N_2021,In_3956,In_2957);
nand U2022 (N_2022,In_3262,In_3363);
or U2023 (N_2023,In_3245,In_486);
or U2024 (N_2024,In_4391,In_2417);
and U2025 (N_2025,In_3009,In_2500);
or U2026 (N_2026,In_3530,In_1930);
or U2027 (N_2027,In_3663,In_3212);
or U2028 (N_2028,In_3173,In_1986);
xnor U2029 (N_2029,In_4215,In_3402);
xnor U2030 (N_2030,In_4597,In_1740);
nand U2031 (N_2031,In_394,In_66);
and U2032 (N_2032,In_2976,In_2533);
nand U2033 (N_2033,In_1523,In_3981);
or U2034 (N_2034,In_4771,In_4417);
nor U2035 (N_2035,In_4357,In_1683);
nor U2036 (N_2036,In_3658,In_3177);
nand U2037 (N_2037,In_4866,In_2038);
and U2038 (N_2038,In_892,In_4863);
nor U2039 (N_2039,In_788,In_2093);
nor U2040 (N_2040,In_4383,In_109);
nand U2041 (N_2041,In_4882,In_4501);
nand U2042 (N_2042,In_4231,In_4173);
or U2043 (N_2043,In_4039,In_2489);
nand U2044 (N_2044,In_4310,In_806);
nand U2045 (N_2045,In_4606,In_878);
or U2046 (N_2046,In_4423,In_1031);
or U2047 (N_2047,In_4519,In_3615);
or U2048 (N_2048,In_1054,In_1057);
and U2049 (N_2049,In_3816,In_1335);
or U2050 (N_2050,In_3146,In_349);
nor U2051 (N_2051,In_1052,In_1636);
xor U2052 (N_2052,In_3777,In_2395);
xor U2053 (N_2053,In_1103,In_1079);
or U2054 (N_2054,In_4842,In_2511);
and U2055 (N_2055,In_2055,In_2383);
or U2056 (N_2056,In_272,In_558);
nand U2057 (N_2057,In_2678,In_2745);
or U2058 (N_2058,In_4616,In_2732);
nor U2059 (N_2059,In_3144,In_2939);
xnor U2060 (N_2060,In_2980,In_4623);
nand U2061 (N_2061,In_2212,In_2566);
or U2062 (N_2062,In_4515,In_1605);
and U2063 (N_2063,In_3597,In_921);
xor U2064 (N_2064,In_1728,In_4929);
nand U2065 (N_2065,In_3714,In_3126);
or U2066 (N_2066,In_1368,In_715);
nor U2067 (N_2067,In_488,In_1954);
nor U2068 (N_2068,In_2035,In_3645);
or U2069 (N_2069,In_946,In_215);
and U2070 (N_2070,In_1615,In_1727);
nor U2071 (N_2071,In_4206,In_2854);
xor U2072 (N_2072,In_2064,In_2373);
and U2073 (N_2073,In_319,In_1739);
xnor U2074 (N_2074,In_1515,In_4903);
xnor U2075 (N_2075,In_582,In_3099);
and U2076 (N_2076,In_2690,In_1370);
nand U2077 (N_2077,In_1294,In_371);
nor U2078 (N_2078,In_1914,In_4819);
and U2079 (N_2079,In_4996,In_3355);
or U2080 (N_2080,In_4870,In_4891);
or U2081 (N_2081,In_2187,In_456);
nand U2082 (N_2082,In_4450,In_3670);
nor U2083 (N_2083,In_1066,In_1296);
nor U2084 (N_2084,In_135,In_4669);
xor U2085 (N_2085,In_3988,In_1511);
and U2086 (N_2086,In_1677,In_4110);
xnor U2087 (N_2087,In_4113,In_4407);
or U2088 (N_2088,In_3422,In_4290);
or U2089 (N_2089,In_549,In_4120);
nand U2090 (N_2090,In_860,In_1305);
and U2091 (N_2091,In_2796,In_4636);
xnor U2092 (N_2092,In_3341,In_1242);
xnor U2093 (N_2093,In_4393,In_4631);
nor U2094 (N_2094,In_4435,In_4390);
nand U2095 (N_2095,In_1384,In_2286);
xnor U2096 (N_2096,In_3462,In_1890);
or U2097 (N_2097,In_3394,In_1134);
xnor U2098 (N_2098,In_2613,In_1510);
and U2099 (N_2099,In_49,In_3145);
and U2100 (N_2100,In_1410,In_2095);
and U2101 (N_2101,In_2734,In_1328);
nor U2102 (N_2102,In_96,In_2443);
and U2103 (N_2103,In_1472,In_3414);
nor U2104 (N_2104,In_671,In_3835);
nor U2105 (N_2105,In_4265,In_139);
and U2106 (N_2106,In_3639,In_2218);
or U2107 (N_2107,In_90,In_2165);
xor U2108 (N_2108,In_2292,In_4562);
xor U2109 (N_2109,In_3556,In_2928);
and U2110 (N_2110,In_996,In_1161);
xor U2111 (N_2111,In_3080,In_1148);
or U2112 (N_2112,In_117,In_1928);
nand U2113 (N_2113,In_2213,In_1240);
xor U2114 (N_2114,In_559,In_368);
and U2115 (N_2115,In_2924,In_1142);
nand U2116 (N_2116,In_2824,In_1377);
nand U2117 (N_2117,In_2741,In_1285);
or U2118 (N_2118,In_3125,In_2274);
xor U2119 (N_2119,In_1781,In_753);
or U2120 (N_2120,In_3972,In_3194);
nor U2121 (N_2121,In_4711,In_4406);
nor U2122 (N_2122,In_4853,In_3378);
or U2123 (N_2123,In_585,In_311);
nand U2124 (N_2124,In_489,In_4136);
and U2125 (N_2125,In_1434,In_740);
or U2126 (N_2126,In_415,In_2477);
or U2127 (N_2127,In_120,In_297);
nand U2128 (N_2128,In_3704,In_3078);
xor U2129 (N_2129,In_4805,In_2483);
and U2130 (N_2130,In_3699,In_4701);
nand U2131 (N_2131,In_4585,In_364);
or U2132 (N_2132,In_4481,In_2981);
or U2133 (N_2133,In_1861,In_1582);
nand U2134 (N_2134,In_1868,In_531);
nor U2135 (N_2135,In_2996,In_2341);
nand U2136 (N_2136,In_2773,In_2865);
xnor U2137 (N_2137,In_3230,In_2454);
xnor U2138 (N_2138,In_4233,In_1247);
xnor U2139 (N_2139,In_22,In_2000);
xor U2140 (N_2140,In_1799,In_2712);
or U2141 (N_2141,In_3150,In_677);
xnor U2142 (N_2142,In_675,In_4484);
and U2143 (N_2143,In_2851,In_3312);
xnor U2144 (N_2144,In_1026,In_2457);
and U2145 (N_2145,In_2277,In_3054);
or U2146 (N_2146,In_3716,In_626);
or U2147 (N_2147,In_2158,In_2515);
nor U2148 (N_2148,In_3327,In_2446);
xnor U2149 (N_2149,In_3518,In_936);
and U2150 (N_2150,In_4906,In_2545);
or U2151 (N_2151,In_1467,In_1453);
or U2152 (N_2152,In_907,In_97);
nand U2153 (N_2153,In_1964,In_1226);
nor U2154 (N_2154,In_2942,In_3533);
and U2155 (N_2155,In_1350,In_3987);
and U2156 (N_2156,In_2482,In_2057);
nand U2157 (N_2157,In_4980,In_175);
nand U2158 (N_2158,In_1053,In_4845);
and U2159 (N_2159,In_2532,In_4676);
or U2160 (N_2160,In_1812,In_1414);
and U2161 (N_2161,In_1487,In_3625);
xnor U2162 (N_2162,In_4193,In_1546);
or U2163 (N_2163,In_3442,In_4295);
xor U2164 (N_2164,In_4163,In_4189);
xnor U2165 (N_2165,In_1481,In_1667);
nor U2166 (N_2166,In_2550,In_2207);
or U2167 (N_2167,In_3686,In_2224);
and U2168 (N_2168,In_2167,In_3315);
or U2169 (N_2169,In_1682,In_1754);
nand U2170 (N_2170,In_1831,In_4995);
or U2171 (N_2171,In_2032,In_307);
nor U2172 (N_2172,In_350,In_2222);
nor U2173 (N_2173,In_172,In_2470);
or U2174 (N_2174,In_3103,In_233);
xnor U2175 (N_2175,In_2580,In_458);
nand U2176 (N_2176,In_4556,In_1174);
or U2177 (N_2177,In_1346,In_2217);
and U2178 (N_2178,In_1688,In_2285);
or U2179 (N_2179,In_3566,In_3076);
nand U2180 (N_2180,In_1412,In_1595);
and U2181 (N_2181,In_973,In_1331);
nor U2182 (N_2182,In_2281,In_3234);
nor U2183 (N_2183,In_4463,In_1776);
xor U2184 (N_2184,In_3367,In_1257);
nor U2185 (N_2185,In_2603,In_950);
and U2186 (N_2186,In_501,In_3163);
xnor U2187 (N_2187,In_3007,In_3532);
nor U2188 (N_2188,In_1413,In_4843);
and U2189 (N_2189,In_1931,In_1170);
and U2190 (N_2190,In_2931,In_4957);
or U2191 (N_2191,In_1700,In_2762);
nor U2192 (N_2192,In_933,In_859);
or U2193 (N_2193,In_499,In_1772);
or U2194 (N_2194,In_1932,In_3203);
nand U2195 (N_2195,In_3167,In_330);
or U2196 (N_2196,In_1314,In_2615);
nor U2197 (N_2197,In_1445,In_2081);
nor U2198 (N_2198,In_4584,In_1114);
and U2199 (N_2199,In_4754,In_2250);
or U2200 (N_2200,In_4992,In_900);
xor U2201 (N_2201,In_4642,In_2969);
or U2202 (N_2202,In_3065,In_3297);
xnor U2203 (N_2203,In_4132,In_1610);
xor U2204 (N_2204,In_3813,In_259);
xnor U2205 (N_2205,In_1476,In_1450);
or U2206 (N_2206,In_2010,In_3485);
nor U2207 (N_2207,In_3569,In_2975);
nor U2208 (N_2208,In_3553,In_1681);
xor U2209 (N_2209,In_3269,In_57);
xnor U2210 (N_2210,In_1050,In_1199);
or U2211 (N_2211,In_2818,In_2650);
nand U2212 (N_2212,In_75,In_2149);
nand U2213 (N_2213,In_791,In_2679);
xor U2214 (N_2214,In_2962,In_3347);
or U2215 (N_2215,In_3600,In_3649);
xor U2216 (N_2216,In_1642,In_3159);
and U2217 (N_2217,In_2179,In_3836);
or U2218 (N_2218,In_3993,In_1969);
nand U2219 (N_2219,In_4339,In_1333);
or U2220 (N_2220,In_4397,In_4707);
and U2221 (N_2221,In_98,In_2145);
or U2222 (N_2222,In_4948,In_1010);
and U2223 (N_2223,In_1431,In_779);
or U2224 (N_2224,In_4052,In_3592);
or U2225 (N_2225,In_2464,In_657);
nor U2226 (N_2226,In_2096,In_2175);
nand U2227 (N_2227,In_2822,In_4563);
xor U2228 (N_2228,In_1953,In_3383);
or U2229 (N_2229,In_4638,In_337);
and U2230 (N_2230,In_2225,In_1638);
xor U2231 (N_2231,In_4972,In_405);
and U2232 (N_2232,In_3697,In_2181);
and U2233 (N_2233,In_3598,In_3286);
xnor U2234 (N_2234,In_3497,In_2214);
and U2235 (N_2235,In_3875,In_3661);
or U2236 (N_2236,In_4263,In_3635);
and U2237 (N_2237,In_3814,In_643);
or U2238 (N_2238,In_3443,In_3538);
or U2239 (N_2239,In_2689,In_1717);
nor U2240 (N_2240,In_4372,In_3685);
or U2241 (N_2241,In_1401,In_1665);
and U2242 (N_2242,In_4540,In_1059);
and U2243 (N_2243,In_1926,In_1634);
or U2244 (N_2244,In_2684,In_3018);
xor U2245 (N_2245,In_4015,In_4593);
or U2246 (N_2246,In_451,In_2562);
or U2247 (N_2247,In_4415,In_999);
nand U2248 (N_2248,In_3575,In_1632);
nand U2249 (N_2249,In_3156,In_3164);
nor U2250 (N_2250,In_714,In_844);
xor U2251 (N_2251,In_3124,In_4909);
nand U2252 (N_2252,In_1988,In_4789);
or U2253 (N_2253,In_2162,In_4941);
nor U2254 (N_2254,In_1277,In_148);
xor U2255 (N_2255,In_4432,In_1670);
nor U2256 (N_2256,In_1860,In_4464);
xnor U2257 (N_2257,In_4685,In_2486);
xor U2258 (N_2258,In_4027,In_3959);
or U2259 (N_2259,In_968,In_88);
and U2260 (N_2260,In_4680,In_1680);
nand U2261 (N_2261,In_777,In_424);
xnor U2262 (N_2262,In_709,In_2320);
xnor U2263 (N_2263,In_2335,In_4195);
nand U2264 (N_2264,In_207,In_3536);
nor U2265 (N_2265,In_1762,In_857);
nor U2266 (N_2266,In_1563,In_2316);
and U2267 (N_2267,In_1936,In_4076);
or U2268 (N_2268,In_869,In_3857);
xor U2269 (N_2269,In_4607,In_3586);
xor U2270 (N_2270,In_1983,In_728);
nor U2271 (N_2271,In_1416,In_4750);
nand U2272 (N_2272,In_347,In_2391);
and U2273 (N_2273,In_1729,In_161);
nand U2274 (N_2274,In_1503,In_2775);
nor U2275 (N_2275,In_3170,In_2397);
and U2276 (N_2276,In_4743,In_2154);
or U2277 (N_2277,In_1672,In_2177);
xnor U2278 (N_2278,In_515,In_2164);
or U2279 (N_2279,In_3724,In_2174);
xor U2280 (N_2280,In_3572,In_3502);
and U2281 (N_2281,In_1270,In_2926);
or U2282 (N_2282,In_5,In_4793);
and U2283 (N_2283,In_2067,In_1086);
or U2284 (N_2284,In_449,In_3483);
or U2285 (N_2285,In_1420,In_867);
nor U2286 (N_2286,In_2702,In_4192);
nor U2287 (N_2287,In_2421,In_264);
and U2288 (N_2288,In_1784,In_4742);
nor U2289 (N_2289,In_3650,In_3435);
or U2290 (N_2290,In_467,In_534);
nor U2291 (N_2291,In_4240,In_1360);
and U2292 (N_2292,In_4704,In_3388);
and U2293 (N_2293,In_2522,In_4508);
and U2294 (N_2294,In_1810,In_3517);
and U2295 (N_2295,In_2611,In_2109);
or U2296 (N_2296,In_1061,In_1371);
xor U2297 (N_2297,In_2030,In_3842);
xnor U2298 (N_2298,In_755,In_4158);
nand U2299 (N_2299,In_2398,In_621);
and U2300 (N_2300,In_2805,In_3992);
xor U2301 (N_2301,In_568,In_1070);
nor U2302 (N_2302,In_3393,In_1451);
nand U2303 (N_2303,In_2552,In_1228);
xnor U2304 (N_2304,In_2009,In_2435);
nor U2305 (N_2305,In_1275,In_819);
or U2306 (N_2306,In_770,In_1201);
nor U2307 (N_2307,In_2204,In_1535);
or U2308 (N_2308,In_1344,In_2253);
or U2309 (N_2309,In_4617,In_3643);
xnor U2310 (N_2310,In_2677,In_3044);
or U2311 (N_2311,In_2808,In_4857);
nor U2312 (N_2312,In_3982,In_1062);
or U2313 (N_2313,In_72,In_2467);
nor U2314 (N_2314,In_2514,In_2240);
and U2315 (N_2315,In_3259,In_2092);
nand U2316 (N_2316,In_4325,In_2946);
or U2317 (N_2317,In_3232,In_3739);
or U2318 (N_2318,In_726,In_2587);
or U2319 (N_2319,In_2978,In_4308);
and U2320 (N_2320,In_4571,In_3456);
or U2321 (N_2321,In_1657,In_3190);
and U2322 (N_2322,In_3865,In_1455);
nand U2323 (N_2323,In_747,In_4787);
xnor U2324 (N_2324,In_4717,In_248);
xor U2325 (N_2325,In_3899,In_4764);
or U2326 (N_2326,In_2428,In_454);
nand U2327 (N_2327,In_722,In_3885);
nor U2328 (N_2328,In_4656,In_221);
xnor U2329 (N_2329,In_162,In_2743);
or U2330 (N_2330,In_4802,In_1101);
or U2331 (N_2331,In_1301,In_1913);
xor U2332 (N_2332,In_624,In_3069);
nand U2333 (N_2333,In_2782,In_4729);
nor U2334 (N_2334,In_4475,In_2460);
or U2335 (N_2335,In_1748,In_669);
nand U2336 (N_2336,In_2829,In_1182);
or U2337 (N_2337,In_541,In_611);
nand U2338 (N_2338,In_3225,In_1525);
and U2339 (N_2339,In_939,In_2890);
nand U2340 (N_2340,In_54,In_2897);
and U2341 (N_2341,In_4666,In_323);
nor U2342 (N_2342,In_4810,In_4296);
nor U2343 (N_2343,In_3691,In_376);
and U2344 (N_2344,In_3627,In_1104);
and U2345 (N_2345,In_4155,In_2068);
and U2346 (N_2346,In_3410,In_3270);
or U2347 (N_2347,In_1732,In_3905);
nand U2348 (N_2348,In_1676,In_896);
nand U2349 (N_2349,In_4314,In_4917);
nand U2350 (N_2350,In_1709,In_4582);
or U2351 (N_2351,In_2228,In_402);
or U2352 (N_2352,In_2788,In_380);
and U2353 (N_2353,In_2388,In_346);
nor U2354 (N_2354,In_4908,In_4164);
and U2355 (N_2355,In_4079,In_1738);
nor U2356 (N_2356,In_592,In_4807);
nor U2357 (N_2357,In_529,In_1935);
xnor U2358 (N_2358,In_4535,In_4468);
or U2359 (N_2359,In_3006,In_4521);
nand U2360 (N_2360,In_4378,In_3817);
nor U2361 (N_2361,In_2290,In_4137);
or U2362 (N_2362,In_3968,In_1673);
xor U2363 (N_2363,In_3657,In_3806);
or U2364 (N_2364,In_1212,In_1504);
nand U2365 (N_2365,In_1433,In_1934);
nand U2366 (N_2366,In_4763,In_792);
nor U2367 (N_2367,In_2538,In_2487);
nand U2368 (N_2368,In_4635,In_2220);
or U2369 (N_2369,In_1042,In_3102);
or U2370 (N_2370,In_2860,In_767);
or U2371 (N_2371,In_2554,In_3360);
and U2372 (N_2372,In_4547,In_1715);
xnor U2373 (N_2373,In_4068,In_293);
nand U2374 (N_2374,In_484,In_4881);
and U2375 (N_2375,In_1470,In_308);
nor U2376 (N_2376,In_2586,In_2804);
and U2377 (N_2377,In_3887,In_4626);
or U2378 (N_2378,In_3207,In_535);
and U2379 (N_2379,In_3938,In_4130);
nand U2380 (N_2380,In_3619,In_827);
xor U2381 (N_2381,In_3068,In_3323);
or U2382 (N_2382,In_3140,In_2042);
nand U2383 (N_2383,In_3667,In_678);
and U2384 (N_2384,In_2101,In_1489);
and U2385 (N_2385,In_3638,In_3996);
and U2386 (N_2386,In_4834,In_210);
nand U2387 (N_2387,In_3220,In_2183);
nor U2388 (N_2388,In_150,In_1924);
and U2389 (N_2389,In_73,In_1844);
and U2390 (N_2390,In_1900,In_4366);
and U2391 (N_2391,In_1317,In_2916);
nand U2392 (N_2392,In_734,In_3133);
nor U2393 (N_2393,In_129,In_4083);
and U2394 (N_2394,In_1941,In_601);
nand U2395 (N_2395,In_138,In_2138);
nor U2396 (N_2396,In_3154,In_2249);
and U2397 (N_2397,In_2108,In_2581);
and U2398 (N_2398,In_3213,In_3607);
nand U2399 (N_2399,In_3606,In_343);
nor U2400 (N_2400,In_4896,In_44);
or U2401 (N_2401,In_1607,In_224);
and U2402 (N_2402,In_3189,In_3122);
nand U2403 (N_2403,In_712,In_4089);
xor U2404 (N_2404,In_934,In_4716);
or U2405 (N_2405,In_4862,In_2668);
and U2406 (N_2406,In_2727,In_4467);
xnor U2407 (N_2407,In_3922,In_3884);
or U2408 (N_2408,In_1055,In_4322);
nand U2409 (N_2409,In_1252,In_2429);
or U2410 (N_2410,In_4829,In_1946);
nor U2411 (N_2411,In_2737,In_4095);
or U2412 (N_2412,In_4758,In_1084);
xnor U2413 (N_2413,In_2393,In_889);
or U2414 (N_2414,In_1916,In_786);
nor U2415 (N_2415,In_1500,In_2576);
xor U2416 (N_2416,In_3172,In_3304);
or U2417 (N_2417,In_4414,In_2649);
xnor U2418 (N_2418,In_3802,In_326);
or U2419 (N_2419,In_3271,In_17);
xor U2420 (N_2420,In_4031,In_3613);
nand U2421 (N_2421,In_1146,In_4429);
nor U2422 (N_2422,In_3896,In_2310);
and U2423 (N_2423,In_3366,In_1111);
and U2424 (N_2424,In_305,In_1819);
nand U2425 (N_2425,In_136,In_2345);
xor U2426 (N_2426,In_576,In_2474);
xor U2427 (N_2427,In_2394,In_4224);
nor U2428 (N_2428,In_263,In_1214);
and U2429 (N_2429,In_2616,In_1577);
and U2430 (N_2430,In_587,In_4784);
or U2431 (N_2431,In_742,In_1398);
nand U2432 (N_2432,In_4225,In_3197);
or U2433 (N_2433,In_2134,In_1918);
or U2434 (N_2434,In_3129,In_4147);
and U2435 (N_2435,In_4674,In_4184);
nor U2436 (N_2436,In_1178,In_440);
and U2437 (N_2437,In_1123,In_4112);
nor U2438 (N_2438,In_3431,In_2501);
and U2439 (N_2439,In_1087,In_1995);
or U2440 (N_2440,In_2507,In_707);
xor U2441 (N_2441,In_676,In_565);
nor U2442 (N_2442,In_1124,In_3503);
nand U2443 (N_2443,In_1177,In_4982);
xnor U2444 (N_2444,In_3389,In_1444);
and U2445 (N_2445,In_957,In_523);
or U2446 (N_2446,In_2490,In_1231);
nand U2447 (N_2447,In_787,In_62);
nand U2448 (N_2448,In_2528,In_3161);
xnor U2449 (N_2449,In_38,In_1298);
nand U2450 (N_2450,In_935,In_3115);
nor U2451 (N_2451,In_4140,In_4199);
xnor U2452 (N_2452,In_3499,In_173);
xnor U2453 (N_2453,In_4483,In_2724);
nor U2454 (N_2454,In_1047,In_253);
nand U2455 (N_2455,In_2261,In_1655);
nor U2456 (N_2456,In_3016,In_3665);
or U2457 (N_2457,In_3853,In_3754);
nand U2458 (N_2458,In_3820,In_3058);
xor U2459 (N_2459,In_301,In_462);
nand U2460 (N_2460,In_3585,In_616);
nor U2461 (N_2461,In_2549,In_1130);
xnor U2462 (N_2462,In_1376,In_1224);
nand U2463 (N_2463,In_3929,In_2643);
xnor U2464 (N_2464,In_4811,In_2404);
and U2465 (N_2465,In_4594,In_1533);
and U2466 (N_2466,In_2442,In_3604);
or U2467 (N_2467,In_2060,In_822);
or U2468 (N_2468,In_1121,In_4312);
nor U2469 (N_2469,In_3001,In_4248);
nand U2470 (N_2470,In_2966,In_123);
and U2471 (N_2471,In_7,In_2288);
xor U2472 (N_2472,In_2291,In_289);
and U2473 (N_2473,In_3861,In_4840);
xnor U2474 (N_2474,In_3692,In_3874);
nand U2475 (N_2475,In_1902,In_442);
and U2476 (N_2476,In_112,In_4629);
or U2477 (N_2477,In_2910,In_1960);
and U2478 (N_2478,In_325,In_3741);
and U2479 (N_2479,In_1001,In_2746);
nor U2480 (N_2480,In_2826,In_4651);
nor U2481 (N_2481,In_2469,In_1300);
or U2482 (N_2482,In_2396,In_3487);
or U2483 (N_2483,In_923,In_943);
xor U2484 (N_2484,In_704,In_1702);
or U2485 (N_2485,In_4210,In_4555);
and U2486 (N_2486,In_1779,In_4618);
xnor U2487 (N_2487,In_180,In_3831);
xor U2488 (N_2488,In_2494,In_2205);
xor U2489 (N_2489,In_1668,In_552);
and U2490 (N_2490,In_1326,In_4738);
nand U2491 (N_2491,In_1440,In_4245);
nor U2492 (N_2492,In_2262,In_4945);
or U2493 (N_2493,In_4087,In_4197);
or U2494 (N_2494,In_949,In_1237);
nand U2495 (N_2495,In_802,In_3694);
or U2496 (N_2496,In_48,In_1140);
or U2497 (N_2497,In_2779,In_2758);
and U2498 (N_2498,In_3290,In_927);
xor U2499 (N_2499,In_4687,In_16);
and U2500 (N_2500,In_2767,In_922);
and U2501 (N_2501,In_4238,In_4027);
xnor U2502 (N_2502,In_2816,In_1596);
xor U2503 (N_2503,In_4575,In_72);
nand U2504 (N_2504,In_957,In_3306);
nand U2505 (N_2505,In_1022,In_2545);
xnor U2506 (N_2506,In_828,In_1366);
and U2507 (N_2507,In_1494,In_4732);
and U2508 (N_2508,In_3060,In_4305);
nand U2509 (N_2509,In_2121,In_2048);
xnor U2510 (N_2510,In_4598,In_1109);
or U2511 (N_2511,In_1794,In_1844);
nand U2512 (N_2512,In_476,In_3423);
xor U2513 (N_2513,In_3106,In_1917);
or U2514 (N_2514,In_1290,In_2120);
and U2515 (N_2515,In_401,In_3671);
or U2516 (N_2516,In_891,In_2276);
nand U2517 (N_2517,In_2052,In_141);
or U2518 (N_2518,In_2660,In_4318);
and U2519 (N_2519,In_11,In_2908);
and U2520 (N_2520,In_2948,In_1947);
and U2521 (N_2521,In_72,In_3607);
nand U2522 (N_2522,In_559,In_1640);
and U2523 (N_2523,In_3571,In_2616);
or U2524 (N_2524,In_2942,In_1620);
nand U2525 (N_2525,In_2137,In_119);
nor U2526 (N_2526,In_1828,In_392);
and U2527 (N_2527,In_3734,In_4228);
nor U2528 (N_2528,In_515,In_2187);
nand U2529 (N_2529,In_405,In_743);
xnor U2530 (N_2530,In_3681,In_2744);
or U2531 (N_2531,In_741,In_1929);
xor U2532 (N_2532,In_4438,In_1741);
xor U2533 (N_2533,In_4597,In_3194);
nand U2534 (N_2534,In_3344,In_1020);
xnor U2535 (N_2535,In_2733,In_2806);
xnor U2536 (N_2536,In_3468,In_2973);
or U2537 (N_2537,In_2760,In_778);
and U2538 (N_2538,In_987,In_157);
xnor U2539 (N_2539,In_3399,In_1991);
or U2540 (N_2540,In_4751,In_41);
and U2541 (N_2541,In_507,In_3109);
or U2542 (N_2542,In_4290,In_3396);
and U2543 (N_2543,In_189,In_3289);
xor U2544 (N_2544,In_3614,In_2923);
and U2545 (N_2545,In_3037,In_2901);
and U2546 (N_2546,In_529,In_1974);
xnor U2547 (N_2547,In_4178,In_981);
nand U2548 (N_2548,In_1941,In_233);
and U2549 (N_2549,In_3076,In_3243);
nand U2550 (N_2550,In_2425,In_4601);
or U2551 (N_2551,In_259,In_610);
nand U2552 (N_2552,In_1483,In_108);
nor U2553 (N_2553,In_2083,In_4975);
nor U2554 (N_2554,In_545,In_1545);
xnor U2555 (N_2555,In_1390,In_1264);
or U2556 (N_2556,In_3236,In_61);
xor U2557 (N_2557,In_2275,In_1318);
and U2558 (N_2558,In_3845,In_710);
and U2559 (N_2559,In_411,In_3568);
nor U2560 (N_2560,In_2655,In_1418);
or U2561 (N_2561,In_4998,In_1934);
xnor U2562 (N_2562,In_4104,In_2715);
xor U2563 (N_2563,In_3106,In_2656);
xor U2564 (N_2564,In_1251,In_4624);
nor U2565 (N_2565,In_2137,In_3548);
xnor U2566 (N_2566,In_4245,In_1233);
xor U2567 (N_2567,In_1159,In_2109);
or U2568 (N_2568,In_4286,In_4774);
nor U2569 (N_2569,In_4948,In_926);
nor U2570 (N_2570,In_3480,In_2722);
nor U2571 (N_2571,In_4073,In_474);
nand U2572 (N_2572,In_4897,In_2275);
nor U2573 (N_2573,In_2272,In_740);
nand U2574 (N_2574,In_3871,In_2458);
or U2575 (N_2575,In_3909,In_4969);
xor U2576 (N_2576,In_3035,In_1610);
xnor U2577 (N_2577,In_4355,In_3141);
nor U2578 (N_2578,In_4573,In_3128);
or U2579 (N_2579,In_4146,In_1628);
nor U2580 (N_2580,In_1227,In_2330);
xnor U2581 (N_2581,In_1250,In_21);
xnor U2582 (N_2582,In_1496,In_2249);
or U2583 (N_2583,In_4396,In_4446);
nor U2584 (N_2584,In_199,In_4528);
nand U2585 (N_2585,In_3116,In_4899);
and U2586 (N_2586,In_2698,In_4395);
or U2587 (N_2587,In_2579,In_2476);
and U2588 (N_2588,In_4135,In_1696);
and U2589 (N_2589,In_128,In_2826);
nor U2590 (N_2590,In_2514,In_761);
and U2591 (N_2591,In_2352,In_3484);
nor U2592 (N_2592,In_4744,In_2128);
nand U2593 (N_2593,In_2935,In_963);
or U2594 (N_2594,In_634,In_1148);
or U2595 (N_2595,In_0,In_2219);
or U2596 (N_2596,In_1291,In_4092);
or U2597 (N_2597,In_2168,In_4026);
nor U2598 (N_2598,In_1790,In_4500);
xor U2599 (N_2599,In_4850,In_2496);
nor U2600 (N_2600,In_2783,In_3123);
xor U2601 (N_2601,In_4853,In_82);
nor U2602 (N_2602,In_3551,In_4190);
xor U2603 (N_2603,In_2378,In_4795);
and U2604 (N_2604,In_1224,In_1022);
nor U2605 (N_2605,In_655,In_4930);
and U2606 (N_2606,In_562,In_4316);
or U2607 (N_2607,In_3697,In_4739);
or U2608 (N_2608,In_967,In_1261);
and U2609 (N_2609,In_2823,In_2067);
nor U2610 (N_2610,In_4268,In_3270);
or U2611 (N_2611,In_3124,In_1102);
xor U2612 (N_2612,In_3963,In_1354);
nand U2613 (N_2613,In_3134,In_921);
nor U2614 (N_2614,In_3215,In_910);
and U2615 (N_2615,In_4559,In_3827);
and U2616 (N_2616,In_1322,In_4487);
or U2617 (N_2617,In_3457,In_2605);
nor U2618 (N_2618,In_605,In_3526);
and U2619 (N_2619,In_2599,In_341);
nor U2620 (N_2620,In_2824,In_656);
or U2621 (N_2621,In_3396,In_85);
or U2622 (N_2622,In_3987,In_125);
nor U2623 (N_2623,In_2211,In_1592);
nand U2624 (N_2624,In_2713,In_3314);
xor U2625 (N_2625,In_1655,In_2762);
and U2626 (N_2626,In_1202,In_897);
xnor U2627 (N_2627,In_3404,In_2045);
nor U2628 (N_2628,In_1927,In_4812);
and U2629 (N_2629,In_3374,In_3231);
or U2630 (N_2630,In_3585,In_280);
nor U2631 (N_2631,In_2177,In_4328);
nand U2632 (N_2632,In_2918,In_1396);
nand U2633 (N_2633,In_1576,In_1069);
and U2634 (N_2634,In_538,In_3439);
and U2635 (N_2635,In_265,In_3464);
nor U2636 (N_2636,In_656,In_2443);
xnor U2637 (N_2637,In_1445,In_1647);
or U2638 (N_2638,In_2964,In_89);
nor U2639 (N_2639,In_2468,In_3503);
nand U2640 (N_2640,In_1609,In_3962);
or U2641 (N_2641,In_1807,In_2536);
and U2642 (N_2642,In_3262,In_4485);
nand U2643 (N_2643,In_1091,In_4287);
and U2644 (N_2644,In_4208,In_3237);
and U2645 (N_2645,In_3758,In_1692);
xnor U2646 (N_2646,In_2054,In_4804);
and U2647 (N_2647,In_3962,In_1514);
xor U2648 (N_2648,In_4311,In_3338);
or U2649 (N_2649,In_1149,In_1098);
or U2650 (N_2650,In_2594,In_3262);
and U2651 (N_2651,In_646,In_3647);
and U2652 (N_2652,In_1658,In_4624);
nor U2653 (N_2653,In_3983,In_4366);
nand U2654 (N_2654,In_251,In_1392);
nor U2655 (N_2655,In_2639,In_3273);
nand U2656 (N_2656,In_3235,In_4100);
nor U2657 (N_2657,In_2960,In_2099);
nand U2658 (N_2658,In_145,In_960);
or U2659 (N_2659,In_4044,In_4365);
and U2660 (N_2660,In_3319,In_1858);
and U2661 (N_2661,In_3445,In_2016);
xor U2662 (N_2662,In_1796,In_3004);
nor U2663 (N_2663,In_4067,In_2273);
or U2664 (N_2664,In_4442,In_3598);
nor U2665 (N_2665,In_1954,In_4354);
xor U2666 (N_2666,In_3939,In_4914);
nor U2667 (N_2667,In_243,In_4445);
or U2668 (N_2668,In_4944,In_3617);
nand U2669 (N_2669,In_555,In_78);
or U2670 (N_2670,In_314,In_4693);
and U2671 (N_2671,In_436,In_2074);
and U2672 (N_2672,In_807,In_1125);
nor U2673 (N_2673,In_4894,In_3038);
or U2674 (N_2674,In_3733,In_1626);
or U2675 (N_2675,In_695,In_4637);
nand U2676 (N_2676,In_4880,In_543);
and U2677 (N_2677,In_4197,In_1473);
nand U2678 (N_2678,In_4783,In_1137);
nor U2679 (N_2679,In_2223,In_2320);
nand U2680 (N_2680,In_3130,In_3619);
and U2681 (N_2681,In_1557,In_618);
and U2682 (N_2682,In_4043,In_604);
and U2683 (N_2683,In_1465,In_756);
nor U2684 (N_2684,In_1713,In_4922);
nand U2685 (N_2685,In_2899,In_4345);
nand U2686 (N_2686,In_4417,In_758);
nor U2687 (N_2687,In_4016,In_2838);
nor U2688 (N_2688,In_108,In_3481);
xor U2689 (N_2689,In_602,In_1512);
or U2690 (N_2690,In_3570,In_2677);
nor U2691 (N_2691,In_4613,In_2189);
or U2692 (N_2692,In_1859,In_1266);
xnor U2693 (N_2693,In_2055,In_110);
and U2694 (N_2694,In_3354,In_2182);
or U2695 (N_2695,In_4034,In_3107);
or U2696 (N_2696,In_3413,In_2743);
nand U2697 (N_2697,In_1313,In_68);
and U2698 (N_2698,In_2612,In_3231);
nand U2699 (N_2699,In_3300,In_4827);
or U2700 (N_2700,In_1763,In_789);
or U2701 (N_2701,In_3282,In_4521);
and U2702 (N_2702,In_1208,In_2709);
nand U2703 (N_2703,In_2478,In_2718);
or U2704 (N_2704,In_4040,In_3931);
nor U2705 (N_2705,In_1460,In_1290);
nor U2706 (N_2706,In_3013,In_4970);
xnor U2707 (N_2707,In_4248,In_1371);
xor U2708 (N_2708,In_4325,In_2280);
and U2709 (N_2709,In_719,In_2892);
or U2710 (N_2710,In_2032,In_4684);
nand U2711 (N_2711,In_1098,In_4825);
and U2712 (N_2712,In_1332,In_3669);
or U2713 (N_2713,In_3877,In_4299);
or U2714 (N_2714,In_4770,In_4827);
or U2715 (N_2715,In_4936,In_282);
and U2716 (N_2716,In_1995,In_1531);
and U2717 (N_2717,In_1674,In_2601);
nand U2718 (N_2718,In_779,In_929);
and U2719 (N_2719,In_1597,In_2898);
or U2720 (N_2720,In_2307,In_1128);
nand U2721 (N_2721,In_4589,In_2307);
nand U2722 (N_2722,In_3180,In_3270);
or U2723 (N_2723,In_3963,In_4138);
nor U2724 (N_2724,In_842,In_1795);
nand U2725 (N_2725,In_1038,In_665);
or U2726 (N_2726,In_2078,In_1474);
nand U2727 (N_2727,In_2792,In_2017);
and U2728 (N_2728,In_667,In_3655);
and U2729 (N_2729,In_2890,In_3054);
xnor U2730 (N_2730,In_3786,In_1104);
nor U2731 (N_2731,In_375,In_249);
nand U2732 (N_2732,In_4916,In_2207);
xor U2733 (N_2733,In_3839,In_4987);
xor U2734 (N_2734,In_491,In_2193);
nand U2735 (N_2735,In_3776,In_633);
or U2736 (N_2736,In_3020,In_3236);
nand U2737 (N_2737,In_1648,In_4024);
nand U2738 (N_2738,In_2135,In_4320);
or U2739 (N_2739,In_2151,In_960);
or U2740 (N_2740,In_516,In_2371);
or U2741 (N_2741,In_2090,In_3745);
xnor U2742 (N_2742,In_4050,In_3473);
nor U2743 (N_2743,In_1411,In_3820);
xnor U2744 (N_2744,In_87,In_1652);
xor U2745 (N_2745,In_156,In_2120);
or U2746 (N_2746,In_2880,In_1652);
and U2747 (N_2747,In_73,In_507);
or U2748 (N_2748,In_1471,In_1858);
nand U2749 (N_2749,In_1853,In_4942);
xor U2750 (N_2750,In_4898,In_310);
or U2751 (N_2751,In_4804,In_2179);
xor U2752 (N_2752,In_1184,In_4494);
or U2753 (N_2753,In_164,In_2035);
or U2754 (N_2754,In_170,In_2518);
or U2755 (N_2755,In_4616,In_4963);
nand U2756 (N_2756,In_409,In_1426);
and U2757 (N_2757,In_4536,In_379);
and U2758 (N_2758,In_1375,In_3346);
and U2759 (N_2759,In_2847,In_3246);
nor U2760 (N_2760,In_2208,In_2086);
nor U2761 (N_2761,In_1961,In_181);
nand U2762 (N_2762,In_2904,In_1910);
nand U2763 (N_2763,In_3992,In_957);
nand U2764 (N_2764,In_882,In_3224);
nor U2765 (N_2765,In_10,In_1138);
xor U2766 (N_2766,In_4231,In_2917);
xor U2767 (N_2767,In_4112,In_1593);
nand U2768 (N_2768,In_204,In_3611);
xnor U2769 (N_2769,In_658,In_468);
nor U2770 (N_2770,In_1899,In_2698);
nand U2771 (N_2771,In_3283,In_3359);
nand U2772 (N_2772,In_523,In_2013);
nor U2773 (N_2773,In_1298,In_2181);
xor U2774 (N_2774,In_4419,In_887);
and U2775 (N_2775,In_2111,In_4529);
nand U2776 (N_2776,In_2397,In_2691);
nand U2777 (N_2777,In_3022,In_4696);
and U2778 (N_2778,In_3727,In_2741);
xnor U2779 (N_2779,In_2131,In_760);
nand U2780 (N_2780,In_2256,In_4405);
xnor U2781 (N_2781,In_2263,In_4395);
and U2782 (N_2782,In_3854,In_1273);
or U2783 (N_2783,In_3088,In_4916);
or U2784 (N_2784,In_4071,In_380);
nor U2785 (N_2785,In_3132,In_171);
nand U2786 (N_2786,In_549,In_265);
nand U2787 (N_2787,In_123,In_3878);
nand U2788 (N_2788,In_2707,In_1073);
xnor U2789 (N_2789,In_428,In_1148);
or U2790 (N_2790,In_4839,In_477);
and U2791 (N_2791,In_4161,In_4053);
or U2792 (N_2792,In_1313,In_1998);
xor U2793 (N_2793,In_991,In_3189);
xor U2794 (N_2794,In_2620,In_3824);
nand U2795 (N_2795,In_4551,In_1251);
xnor U2796 (N_2796,In_332,In_1175);
nor U2797 (N_2797,In_3851,In_3064);
nor U2798 (N_2798,In_3805,In_1369);
or U2799 (N_2799,In_1988,In_439);
or U2800 (N_2800,In_1840,In_167);
or U2801 (N_2801,In_1151,In_3231);
nor U2802 (N_2802,In_316,In_65);
or U2803 (N_2803,In_2871,In_585);
xor U2804 (N_2804,In_720,In_3631);
nor U2805 (N_2805,In_3371,In_2802);
nor U2806 (N_2806,In_2798,In_4164);
nand U2807 (N_2807,In_765,In_1820);
nor U2808 (N_2808,In_4660,In_1102);
nand U2809 (N_2809,In_534,In_1178);
and U2810 (N_2810,In_2300,In_1115);
and U2811 (N_2811,In_3810,In_884);
nor U2812 (N_2812,In_4488,In_2827);
and U2813 (N_2813,In_3213,In_2912);
nor U2814 (N_2814,In_4335,In_4261);
xor U2815 (N_2815,In_2071,In_4042);
or U2816 (N_2816,In_4151,In_3285);
nor U2817 (N_2817,In_4201,In_2301);
xnor U2818 (N_2818,In_4365,In_4019);
nor U2819 (N_2819,In_3579,In_813);
nor U2820 (N_2820,In_2308,In_31);
xnor U2821 (N_2821,In_952,In_4012);
nand U2822 (N_2822,In_4396,In_2516);
nand U2823 (N_2823,In_2034,In_3645);
and U2824 (N_2824,In_4467,In_3967);
xor U2825 (N_2825,In_1702,In_1831);
and U2826 (N_2826,In_4997,In_2925);
and U2827 (N_2827,In_4122,In_4098);
or U2828 (N_2828,In_569,In_3366);
nor U2829 (N_2829,In_1510,In_2167);
and U2830 (N_2830,In_2754,In_231);
and U2831 (N_2831,In_820,In_2038);
and U2832 (N_2832,In_4343,In_88);
nand U2833 (N_2833,In_3594,In_1084);
nand U2834 (N_2834,In_1405,In_723);
and U2835 (N_2835,In_1303,In_4425);
nor U2836 (N_2836,In_2800,In_4687);
nand U2837 (N_2837,In_3896,In_685);
nand U2838 (N_2838,In_1579,In_4595);
or U2839 (N_2839,In_3960,In_2511);
or U2840 (N_2840,In_1198,In_3247);
nor U2841 (N_2841,In_4117,In_4506);
nor U2842 (N_2842,In_3786,In_2768);
and U2843 (N_2843,In_1242,In_3797);
nor U2844 (N_2844,In_4689,In_2074);
and U2845 (N_2845,In_1769,In_1679);
and U2846 (N_2846,In_254,In_4973);
nor U2847 (N_2847,In_4510,In_2011);
nand U2848 (N_2848,In_25,In_610);
xor U2849 (N_2849,In_1206,In_4302);
and U2850 (N_2850,In_4394,In_1304);
and U2851 (N_2851,In_4095,In_1896);
or U2852 (N_2852,In_4446,In_2044);
or U2853 (N_2853,In_1325,In_795);
xnor U2854 (N_2854,In_2057,In_4799);
or U2855 (N_2855,In_4329,In_1754);
or U2856 (N_2856,In_840,In_4890);
nand U2857 (N_2857,In_136,In_2039);
nor U2858 (N_2858,In_1193,In_3507);
or U2859 (N_2859,In_3185,In_61);
nand U2860 (N_2860,In_4185,In_4013);
or U2861 (N_2861,In_3636,In_596);
nand U2862 (N_2862,In_1500,In_481);
or U2863 (N_2863,In_1897,In_1076);
and U2864 (N_2864,In_643,In_4950);
and U2865 (N_2865,In_3654,In_3691);
and U2866 (N_2866,In_4513,In_4369);
nand U2867 (N_2867,In_876,In_4060);
and U2868 (N_2868,In_3876,In_3831);
or U2869 (N_2869,In_375,In_3386);
or U2870 (N_2870,In_2598,In_22);
xor U2871 (N_2871,In_2532,In_1142);
nand U2872 (N_2872,In_2257,In_1022);
or U2873 (N_2873,In_490,In_1245);
nand U2874 (N_2874,In_162,In_3834);
nor U2875 (N_2875,In_2963,In_481);
nand U2876 (N_2876,In_2772,In_3124);
nand U2877 (N_2877,In_3785,In_4511);
nor U2878 (N_2878,In_1568,In_4944);
nand U2879 (N_2879,In_924,In_233);
and U2880 (N_2880,In_122,In_2934);
nand U2881 (N_2881,In_3875,In_4548);
nor U2882 (N_2882,In_1652,In_2105);
or U2883 (N_2883,In_707,In_143);
nand U2884 (N_2884,In_738,In_4661);
nor U2885 (N_2885,In_1091,In_2300);
and U2886 (N_2886,In_1404,In_2157);
nand U2887 (N_2887,In_3452,In_3290);
nand U2888 (N_2888,In_1999,In_1404);
and U2889 (N_2889,In_1584,In_872);
or U2890 (N_2890,In_1785,In_824);
or U2891 (N_2891,In_2578,In_3575);
nand U2892 (N_2892,In_459,In_3451);
nand U2893 (N_2893,In_4598,In_3661);
xnor U2894 (N_2894,In_3919,In_2315);
and U2895 (N_2895,In_4199,In_2843);
and U2896 (N_2896,In_4213,In_1943);
and U2897 (N_2897,In_1371,In_2448);
nor U2898 (N_2898,In_167,In_142);
xnor U2899 (N_2899,In_3116,In_4549);
xnor U2900 (N_2900,In_769,In_598);
xor U2901 (N_2901,In_4035,In_1864);
or U2902 (N_2902,In_3455,In_688);
nand U2903 (N_2903,In_1469,In_264);
or U2904 (N_2904,In_1594,In_2011);
nand U2905 (N_2905,In_3676,In_3696);
xnor U2906 (N_2906,In_1146,In_810);
and U2907 (N_2907,In_4614,In_4373);
xor U2908 (N_2908,In_2921,In_708);
nand U2909 (N_2909,In_998,In_2970);
nand U2910 (N_2910,In_664,In_1714);
and U2911 (N_2911,In_2329,In_973);
or U2912 (N_2912,In_1904,In_47);
nor U2913 (N_2913,In_1796,In_2439);
and U2914 (N_2914,In_1208,In_4825);
and U2915 (N_2915,In_868,In_12);
nor U2916 (N_2916,In_3752,In_1320);
or U2917 (N_2917,In_908,In_4594);
and U2918 (N_2918,In_2572,In_1348);
and U2919 (N_2919,In_1508,In_2281);
nand U2920 (N_2920,In_4016,In_4384);
xor U2921 (N_2921,In_783,In_719);
xnor U2922 (N_2922,In_120,In_1429);
and U2923 (N_2923,In_1322,In_3119);
xor U2924 (N_2924,In_2272,In_1006);
and U2925 (N_2925,In_2426,In_59);
xor U2926 (N_2926,In_3875,In_4368);
or U2927 (N_2927,In_598,In_3922);
or U2928 (N_2928,In_3525,In_4485);
xor U2929 (N_2929,In_400,In_404);
or U2930 (N_2930,In_4680,In_1958);
nor U2931 (N_2931,In_2795,In_4954);
and U2932 (N_2932,In_2595,In_4963);
xor U2933 (N_2933,In_2396,In_4023);
or U2934 (N_2934,In_226,In_3903);
nor U2935 (N_2935,In_2255,In_4736);
nand U2936 (N_2936,In_2844,In_261);
nor U2937 (N_2937,In_2402,In_1850);
and U2938 (N_2938,In_4279,In_348);
nand U2939 (N_2939,In_701,In_181);
nand U2940 (N_2940,In_993,In_948);
and U2941 (N_2941,In_342,In_217);
and U2942 (N_2942,In_197,In_661);
and U2943 (N_2943,In_2132,In_2834);
nand U2944 (N_2944,In_368,In_4659);
and U2945 (N_2945,In_898,In_784);
nor U2946 (N_2946,In_606,In_1293);
or U2947 (N_2947,In_2550,In_178);
xor U2948 (N_2948,In_2863,In_3911);
xor U2949 (N_2949,In_4211,In_3033);
nand U2950 (N_2950,In_285,In_4727);
and U2951 (N_2951,In_1166,In_1311);
or U2952 (N_2952,In_4224,In_414);
and U2953 (N_2953,In_3038,In_348);
xor U2954 (N_2954,In_1945,In_4806);
nor U2955 (N_2955,In_148,In_1123);
nand U2956 (N_2956,In_1170,In_3680);
xor U2957 (N_2957,In_3799,In_2696);
xor U2958 (N_2958,In_1495,In_3902);
nand U2959 (N_2959,In_4853,In_4920);
and U2960 (N_2960,In_2858,In_2674);
nand U2961 (N_2961,In_971,In_149);
and U2962 (N_2962,In_3107,In_4579);
nand U2963 (N_2963,In_3439,In_646);
nor U2964 (N_2964,In_4788,In_2992);
and U2965 (N_2965,In_4496,In_1410);
and U2966 (N_2966,In_193,In_4172);
xnor U2967 (N_2967,In_1266,In_1165);
nand U2968 (N_2968,In_561,In_4787);
and U2969 (N_2969,In_370,In_1719);
nand U2970 (N_2970,In_1882,In_1260);
or U2971 (N_2971,In_1189,In_1821);
and U2972 (N_2972,In_1058,In_4372);
nand U2973 (N_2973,In_326,In_121);
or U2974 (N_2974,In_1885,In_389);
nand U2975 (N_2975,In_3031,In_1719);
nand U2976 (N_2976,In_1860,In_1457);
or U2977 (N_2977,In_3911,In_2783);
or U2978 (N_2978,In_1967,In_2919);
and U2979 (N_2979,In_288,In_925);
nand U2980 (N_2980,In_4551,In_750);
nor U2981 (N_2981,In_2912,In_4633);
nand U2982 (N_2982,In_3809,In_1581);
nand U2983 (N_2983,In_18,In_2209);
or U2984 (N_2984,In_4964,In_2173);
and U2985 (N_2985,In_1723,In_1238);
nand U2986 (N_2986,In_3339,In_2464);
nor U2987 (N_2987,In_4478,In_1059);
or U2988 (N_2988,In_119,In_3849);
xnor U2989 (N_2989,In_4435,In_4980);
nand U2990 (N_2990,In_2259,In_932);
xnor U2991 (N_2991,In_540,In_331);
nor U2992 (N_2992,In_3973,In_1018);
xor U2993 (N_2993,In_2684,In_3962);
nor U2994 (N_2994,In_3317,In_4463);
and U2995 (N_2995,In_1781,In_3933);
nor U2996 (N_2996,In_1545,In_1610);
or U2997 (N_2997,In_2034,In_3815);
and U2998 (N_2998,In_764,In_3785);
xor U2999 (N_2999,In_4139,In_2993);
or U3000 (N_3000,In_879,In_2949);
xnor U3001 (N_3001,In_2304,In_180);
xor U3002 (N_3002,In_2815,In_3095);
or U3003 (N_3003,In_2362,In_4932);
or U3004 (N_3004,In_1871,In_4291);
nor U3005 (N_3005,In_4510,In_1763);
nor U3006 (N_3006,In_3109,In_648);
or U3007 (N_3007,In_3829,In_2363);
or U3008 (N_3008,In_1401,In_3928);
nor U3009 (N_3009,In_901,In_886);
nand U3010 (N_3010,In_1088,In_855);
xnor U3011 (N_3011,In_1794,In_1127);
nor U3012 (N_3012,In_2579,In_2441);
nor U3013 (N_3013,In_2540,In_3212);
or U3014 (N_3014,In_852,In_1757);
xnor U3015 (N_3015,In_4694,In_984);
nor U3016 (N_3016,In_3162,In_3804);
or U3017 (N_3017,In_148,In_663);
nand U3018 (N_3018,In_3148,In_774);
and U3019 (N_3019,In_3077,In_4914);
nand U3020 (N_3020,In_1624,In_283);
nor U3021 (N_3021,In_3171,In_4412);
and U3022 (N_3022,In_3033,In_3802);
or U3023 (N_3023,In_4966,In_3147);
or U3024 (N_3024,In_847,In_1582);
xor U3025 (N_3025,In_2514,In_641);
and U3026 (N_3026,In_3916,In_4666);
nor U3027 (N_3027,In_3576,In_3516);
nor U3028 (N_3028,In_3481,In_4222);
nor U3029 (N_3029,In_1993,In_2046);
or U3030 (N_3030,In_4719,In_3601);
xnor U3031 (N_3031,In_1362,In_1559);
or U3032 (N_3032,In_3871,In_1778);
nand U3033 (N_3033,In_2160,In_3555);
xnor U3034 (N_3034,In_4160,In_2955);
nand U3035 (N_3035,In_2624,In_4431);
or U3036 (N_3036,In_2458,In_2372);
and U3037 (N_3037,In_2800,In_814);
nand U3038 (N_3038,In_4686,In_994);
or U3039 (N_3039,In_1866,In_3446);
or U3040 (N_3040,In_4002,In_1285);
and U3041 (N_3041,In_2955,In_691);
or U3042 (N_3042,In_3098,In_3227);
nand U3043 (N_3043,In_3173,In_4692);
and U3044 (N_3044,In_4723,In_2370);
nand U3045 (N_3045,In_125,In_4841);
xnor U3046 (N_3046,In_2125,In_479);
and U3047 (N_3047,In_2259,In_3880);
nand U3048 (N_3048,In_2721,In_3675);
nand U3049 (N_3049,In_1223,In_1743);
nor U3050 (N_3050,In_4820,In_922);
or U3051 (N_3051,In_1143,In_168);
or U3052 (N_3052,In_502,In_1871);
xnor U3053 (N_3053,In_2852,In_2331);
and U3054 (N_3054,In_73,In_3974);
nor U3055 (N_3055,In_2234,In_3435);
xor U3056 (N_3056,In_569,In_2040);
nand U3057 (N_3057,In_2000,In_3080);
or U3058 (N_3058,In_4246,In_2762);
nor U3059 (N_3059,In_2603,In_3820);
nor U3060 (N_3060,In_816,In_1826);
or U3061 (N_3061,In_622,In_4872);
or U3062 (N_3062,In_1316,In_4729);
nor U3063 (N_3063,In_3831,In_3646);
and U3064 (N_3064,In_1755,In_477);
or U3065 (N_3065,In_259,In_3256);
nand U3066 (N_3066,In_217,In_1854);
nor U3067 (N_3067,In_4471,In_2030);
xnor U3068 (N_3068,In_1172,In_4375);
xnor U3069 (N_3069,In_4704,In_4619);
nand U3070 (N_3070,In_2917,In_2033);
xor U3071 (N_3071,In_4405,In_1244);
xnor U3072 (N_3072,In_2887,In_3998);
and U3073 (N_3073,In_2436,In_2426);
and U3074 (N_3074,In_4171,In_2963);
or U3075 (N_3075,In_2530,In_3387);
nand U3076 (N_3076,In_4086,In_2464);
or U3077 (N_3077,In_1353,In_4000);
nand U3078 (N_3078,In_4571,In_3069);
nand U3079 (N_3079,In_1345,In_2180);
nor U3080 (N_3080,In_4940,In_2071);
xor U3081 (N_3081,In_486,In_1747);
nor U3082 (N_3082,In_1584,In_2620);
and U3083 (N_3083,In_2549,In_4349);
or U3084 (N_3084,In_457,In_4694);
or U3085 (N_3085,In_3460,In_3988);
nor U3086 (N_3086,In_2073,In_587);
and U3087 (N_3087,In_1084,In_2596);
nand U3088 (N_3088,In_33,In_1047);
nor U3089 (N_3089,In_1277,In_2218);
nor U3090 (N_3090,In_4100,In_2765);
nand U3091 (N_3091,In_1883,In_2442);
or U3092 (N_3092,In_3250,In_4893);
nand U3093 (N_3093,In_2823,In_4455);
xor U3094 (N_3094,In_2923,In_4937);
nand U3095 (N_3095,In_3533,In_4136);
and U3096 (N_3096,In_675,In_3978);
nand U3097 (N_3097,In_2710,In_3171);
nor U3098 (N_3098,In_2730,In_4785);
xor U3099 (N_3099,In_3975,In_3146);
and U3100 (N_3100,In_4381,In_4667);
or U3101 (N_3101,In_3324,In_1968);
or U3102 (N_3102,In_1652,In_1950);
and U3103 (N_3103,In_2321,In_662);
or U3104 (N_3104,In_2282,In_4091);
and U3105 (N_3105,In_2160,In_737);
or U3106 (N_3106,In_2021,In_2462);
nand U3107 (N_3107,In_4965,In_2988);
nor U3108 (N_3108,In_1809,In_1217);
and U3109 (N_3109,In_4927,In_170);
or U3110 (N_3110,In_716,In_3123);
nand U3111 (N_3111,In_968,In_1815);
xor U3112 (N_3112,In_752,In_25);
and U3113 (N_3113,In_1640,In_1838);
and U3114 (N_3114,In_4940,In_1252);
nand U3115 (N_3115,In_2094,In_2136);
or U3116 (N_3116,In_3005,In_2219);
xnor U3117 (N_3117,In_3849,In_4734);
or U3118 (N_3118,In_3600,In_442);
and U3119 (N_3119,In_1612,In_1259);
and U3120 (N_3120,In_3259,In_2162);
or U3121 (N_3121,In_4764,In_566);
nand U3122 (N_3122,In_3150,In_3994);
and U3123 (N_3123,In_1885,In_3734);
nor U3124 (N_3124,In_2673,In_1578);
or U3125 (N_3125,In_2789,In_1160);
nand U3126 (N_3126,In_569,In_2556);
or U3127 (N_3127,In_4866,In_2023);
and U3128 (N_3128,In_906,In_1926);
nand U3129 (N_3129,In_4486,In_1973);
and U3130 (N_3130,In_4773,In_3017);
xor U3131 (N_3131,In_4365,In_2263);
and U3132 (N_3132,In_269,In_4780);
nand U3133 (N_3133,In_2143,In_4299);
nand U3134 (N_3134,In_2752,In_980);
nor U3135 (N_3135,In_2288,In_2684);
xnor U3136 (N_3136,In_4250,In_579);
nand U3137 (N_3137,In_2573,In_3442);
and U3138 (N_3138,In_718,In_1235);
xor U3139 (N_3139,In_295,In_2183);
or U3140 (N_3140,In_2155,In_643);
or U3141 (N_3141,In_217,In_3299);
or U3142 (N_3142,In_1232,In_1344);
or U3143 (N_3143,In_2714,In_325);
and U3144 (N_3144,In_3136,In_3708);
and U3145 (N_3145,In_2216,In_4929);
nand U3146 (N_3146,In_2739,In_2845);
and U3147 (N_3147,In_3820,In_262);
xnor U3148 (N_3148,In_4989,In_2579);
nand U3149 (N_3149,In_4089,In_2049);
or U3150 (N_3150,In_1049,In_3635);
xor U3151 (N_3151,In_13,In_4803);
nor U3152 (N_3152,In_2141,In_4728);
or U3153 (N_3153,In_1672,In_512);
nor U3154 (N_3154,In_3671,In_2122);
xor U3155 (N_3155,In_4749,In_3848);
xor U3156 (N_3156,In_2766,In_2491);
nor U3157 (N_3157,In_451,In_200);
xor U3158 (N_3158,In_1049,In_1746);
and U3159 (N_3159,In_323,In_3966);
xor U3160 (N_3160,In_3121,In_1179);
nor U3161 (N_3161,In_3722,In_4570);
or U3162 (N_3162,In_4149,In_2524);
nor U3163 (N_3163,In_23,In_2526);
xnor U3164 (N_3164,In_2046,In_4883);
nor U3165 (N_3165,In_274,In_2291);
nand U3166 (N_3166,In_2265,In_2789);
nand U3167 (N_3167,In_3685,In_4285);
or U3168 (N_3168,In_3260,In_4557);
nand U3169 (N_3169,In_582,In_2437);
and U3170 (N_3170,In_1967,In_62);
and U3171 (N_3171,In_1547,In_1922);
nor U3172 (N_3172,In_941,In_511);
and U3173 (N_3173,In_4035,In_2299);
nand U3174 (N_3174,In_1729,In_3324);
nor U3175 (N_3175,In_3101,In_579);
nor U3176 (N_3176,In_734,In_2138);
nand U3177 (N_3177,In_1141,In_3613);
nor U3178 (N_3178,In_3370,In_2640);
and U3179 (N_3179,In_1426,In_2840);
or U3180 (N_3180,In_4357,In_642);
nor U3181 (N_3181,In_4096,In_1438);
nand U3182 (N_3182,In_2288,In_586);
or U3183 (N_3183,In_2998,In_1606);
or U3184 (N_3184,In_338,In_1073);
or U3185 (N_3185,In_3723,In_4876);
xnor U3186 (N_3186,In_3614,In_3958);
xnor U3187 (N_3187,In_4717,In_2588);
nor U3188 (N_3188,In_813,In_525);
xor U3189 (N_3189,In_4247,In_3276);
and U3190 (N_3190,In_2011,In_1603);
and U3191 (N_3191,In_4727,In_330);
nand U3192 (N_3192,In_2880,In_2520);
xnor U3193 (N_3193,In_4603,In_1115);
or U3194 (N_3194,In_2221,In_4247);
nor U3195 (N_3195,In_4040,In_816);
xnor U3196 (N_3196,In_806,In_4290);
nor U3197 (N_3197,In_1866,In_4172);
nor U3198 (N_3198,In_1808,In_933);
or U3199 (N_3199,In_4191,In_4770);
nor U3200 (N_3200,In_2094,In_2591);
or U3201 (N_3201,In_470,In_1526);
nor U3202 (N_3202,In_1753,In_1905);
nor U3203 (N_3203,In_895,In_3040);
nand U3204 (N_3204,In_1218,In_2063);
or U3205 (N_3205,In_1425,In_1726);
or U3206 (N_3206,In_1816,In_1612);
xor U3207 (N_3207,In_830,In_4468);
and U3208 (N_3208,In_1682,In_3708);
and U3209 (N_3209,In_2233,In_2674);
nand U3210 (N_3210,In_4277,In_1290);
and U3211 (N_3211,In_4087,In_2266);
nor U3212 (N_3212,In_1330,In_4285);
or U3213 (N_3213,In_1012,In_3900);
nor U3214 (N_3214,In_232,In_470);
or U3215 (N_3215,In_1978,In_951);
and U3216 (N_3216,In_68,In_3082);
xor U3217 (N_3217,In_1343,In_1362);
and U3218 (N_3218,In_3785,In_881);
nand U3219 (N_3219,In_4824,In_1130);
nand U3220 (N_3220,In_3691,In_2906);
nand U3221 (N_3221,In_4055,In_3211);
xnor U3222 (N_3222,In_4148,In_3886);
nor U3223 (N_3223,In_2597,In_2169);
or U3224 (N_3224,In_1399,In_2969);
nand U3225 (N_3225,In_1214,In_1748);
xor U3226 (N_3226,In_3847,In_2469);
or U3227 (N_3227,In_3121,In_3584);
xnor U3228 (N_3228,In_502,In_1910);
nor U3229 (N_3229,In_1345,In_4772);
and U3230 (N_3230,In_2301,In_1025);
or U3231 (N_3231,In_4336,In_1355);
xor U3232 (N_3232,In_3999,In_4170);
nand U3233 (N_3233,In_4630,In_1667);
xnor U3234 (N_3234,In_1545,In_4080);
nor U3235 (N_3235,In_1750,In_2415);
xor U3236 (N_3236,In_4286,In_2681);
xor U3237 (N_3237,In_3097,In_4934);
nor U3238 (N_3238,In_906,In_4327);
and U3239 (N_3239,In_3561,In_2450);
or U3240 (N_3240,In_2998,In_1586);
or U3241 (N_3241,In_1402,In_1589);
and U3242 (N_3242,In_2132,In_3120);
nor U3243 (N_3243,In_195,In_4887);
nor U3244 (N_3244,In_4523,In_4461);
nor U3245 (N_3245,In_1225,In_3243);
and U3246 (N_3246,In_1580,In_3288);
nor U3247 (N_3247,In_3116,In_1274);
nor U3248 (N_3248,In_1315,In_2345);
xnor U3249 (N_3249,In_2332,In_4150);
nor U3250 (N_3250,In_4530,In_1925);
or U3251 (N_3251,In_4369,In_3156);
or U3252 (N_3252,In_1924,In_215);
and U3253 (N_3253,In_1623,In_2472);
and U3254 (N_3254,In_4544,In_4126);
and U3255 (N_3255,In_94,In_1997);
xor U3256 (N_3256,In_3387,In_2557);
nand U3257 (N_3257,In_3626,In_433);
nor U3258 (N_3258,In_3030,In_2968);
nor U3259 (N_3259,In_4519,In_247);
xnor U3260 (N_3260,In_2171,In_3551);
and U3261 (N_3261,In_3642,In_4714);
or U3262 (N_3262,In_2949,In_2651);
and U3263 (N_3263,In_1275,In_2924);
nand U3264 (N_3264,In_736,In_1102);
nor U3265 (N_3265,In_2727,In_979);
or U3266 (N_3266,In_2362,In_1340);
or U3267 (N_3267,In_1216,In_2310);
nor U3268 (N_3268,In_4707,In_970);
xor U3269 (N_3269,In_1255,In_4609);
and U3270 (N_3270,In_2643,In_535);
nor U3271 (N_3271,In_1730,In_4914);
xor U3272 (N_3272,In_3497,In_1447);
or U3273 (N_3273,In_4739,In_1445);
and U3274 (N_3274,In_1198,In_1146);
xor U3275 (N_3275,In_1742,In_3647);
and U3276 (N_3276,In_2188,In_3003);
nor U3277 (N_3277,In_422,In_1066);
xnor U3278 (N_3278,In_4968,In_2163);
nand U3279 (N_3279,In_587,In_3693);
and U3280 (N_3280,In_2354,In_1261);
and U3281 (N_3281,In_1470,In_1281);
nor U3282 (N_3282,In_1143,In_2206);
nand U3283 (N_3283,In_4075,In_2352);
nor U3284 (N_3284,In_3544,In_1555);
nor U3285 (N_3285,In_4382,In_2121);
xnor U3286 (N_3286,In_2494,In_2364);
nand U3287 (N_3287,In_2570,In_4708);
nor U3288 (N_3288,In_2641,In_1342);
and U3289 (N_3289,In_2230,In_1205);
and U3290 (N_3290,In_859,In_4326);
nand U3291 (N_3291,In_4085,In_2165);
nand U3292 (N_3292,In_1691,In_303);
and U3293 (N_3293,In_1436,In_2319);
and U3294 (N_3294,In_4994,In_4891);
xnor U3295 (N_3295,In_2086,In_618);
and U3296 (N_3296,In_597,In_3861);
xnor U3297 (N_3297,In_1611,In_2064);
and U3298 (N_3298,In_1670,In_4618);
nor U3299 (N_3299,In_2484,In_1355);
or U3300 (N_3300,In_2924,In_2383);
or U3301 (N_3301,In_3735,In_63);
or U3302 (N_3302,In_4158,In_4439);
or U3303 (N_3303,In_4094,In_2992);
xnor U3304 (N_3304,In_258,In_428);
xnor U3305 (N_3305,In_3708,In_2396);
nand U3306 (N_3306,In_2840,In_1410);
or U3307 (N_3307,In_2320,In_3633);
and U3308 (N_3308,In_3302,In_687);
and U3309 (N_3309,In_2117,In_3816);
nand U3310 (N_3310,In_4219,In_823);
and U3311 (N_3311,In_319,In_2338);
xnor U3312 (N_3312,In_4762,In_1198);
xor U3313 (N_3313,In_3818,In_1479);
nor U3314 (N_3314,In_4155,In_3880);
or U3315 (N_3315,In_3145,In_4703);
or U3316 (N_3316,In_105,In_2776);
nand U3317 (N_3317,In_3796,In_1691);
nor U3318 (N_3318,In_2145,In_2131);
or U3319 (N_3319,In_237,In_4037);
nor U3320 (N_3320,In_3827,In_1456);
nor U3321 (N_3321,In_658,In_2371);
nand U3322 (N_3322,In_1053,In_765);
or U3323 (N_3323,In_289,In_4859);
or U3324 (N_3324,In_3968,In_459);
or U3325 (N_3325,In_4173,In_1325);
or U3326 (N_3326,In_4113,In_1730);
or U3327 (N_3327,In_4500,In_1016);
nand U3328 (N_3328,In_4325,In_2513);
and U3329 (N_3329,In_2234,In_2036);
nor U3330 (N_3330,In_658,In_2374);
and U3331 (N_3331,In_1329,In_3717);
nor U3332 (N_3332,In_4852,In_362);
nand U3333 (N_3333,In_3633,In_4643);
nor U3334 (N_3334,In_3340,In_2619);
and U3335 (N_3335,In_825,In_308);
nand U3336 (N_3336,In_4436,In_1076);
xnor U3337 (N_3337,In_3919,In_4799);
xnor U3338 (N_3338,In_1089,In_534);
and U3339 (N_3339,In_2425,In_3077);
xnor U3340 (N_3340,In_192,In_2458);
nor U3341 (N_3341,In_64,In_3039);
nor U3342 (N_3342,In_2083,In_1152);
xor U3343 (N_3343,In_141,In_576);
nand U3344 (N_3344,In_3786,In_3061);
nor U3345 (N_3345,In_247,In_4324);
nor U3346 (N_3346,In_4192,In_3438);
and U3347 (N_3347,In_1334,In_3098);
nand U3348 (N_3348,In_2525,In_2042);
nand U3349 (N_3349,In_493,In_4818);
and U3350 (N_3350,In_4453,In_1897);
or U3351 (N_3351,In_1625,In_4162);
and U3352 (N_3352,In_3986,In_2163);
xor U3353 (N_3353,In_3851,In_3222);
nand U3354 (N_3354,In_767,In_1311);
xor U3355 (N_3355,In_4954,In_3974);
nor U3356 (N_3356,In_4488,In_2771);
nor U3357 (N_3357,In_2650,In_2532);
and U3358 (N_3358,In_2379,In_688);
and U3359 (N_3359,In_2138,In_2634);
nand U3360 (N_3360,In_3437,In_4145);
or U3361 (N_3361,In_1131,In_3661);
or U3362 (N_3362,In_268,In_3665);
or U3363 (N_3363,In_4512,In_2417);
nand U3364 (N_3364,In_3677,In_2692);
xnor U3365 (N_3365,In_1074,In_834);
nand U3366 (N_3366,In_3551,In_273);
nor U3367 (N_3367,In_3380,In_553);
or U3368 (N_3368,In_208,In_4982);
nand U3369 (N_3369,In_490,In_4504);
xor U3370 (N_3370,In_3866,In_3657);
nor U3371 (N_3371,In_2902,In_578);
and U3372 (N_3372,In_1007,In_4688);
and U3373 (N_3373,In_2721,In_695);
nand U3374 (N_3374,In_4509,In_4047);
and U3375 (N_3375,In_4263,In_2753);
nand U3376 (N_3376,In_3418,In_278);
nor U3377 (N_3377,In_4870,In_350);
or U3378 (N_3378,In_1091,In_4887);
and U3379 (N_3379,In_171,In_2659);
nand U3380 (N_3380,In_3304,In_165);
nand U3381 (N_3381,In_3158,In_1848);
nand U3382 (N_3382,In_92,In_4509);
nor U3383 (N_3383,In_666,In_736);
or U3384 (N_3384,In_892,In_681);
or U3385 (N_3385,In_381,In_3849);
nor U3386 (N_3386,In_81,In_3227);
xor U3387 (N_3387,In_145,In_1294);
xnor U3388 (N_3388,In_3497,In_4220);
xnor U3389 (N_3389,In_3137,In_376);
and U3390 (N_3390,In_2853,In_4576);
and U3391 (N_3391,In_1740,In_2907);
or U3392 (N_3392,In_2200,In_4507);
nand U3393 (N_3393,In_3971,In_3);
xnor U3394 (N_3394,In_760,In_4290);
xor U3395 (N_3395,In_279,In_3989);
nor U3396 (N_3396,In_2165,In_3474);
xor U3397 (N_3397,In_2736,In_4839);
and U3398 (N_3398,In_996,In_2392);
nor U3399 (N_3399,In_3181,In_477);
and U3400 (N_3400,In_624,In_3716);
and U3401 (N_3401,In_2675,In_351);
and U3402 (N_3402,In_675,In_1380);
nor U3403 (N_3403,In_2912,In_4354);
or U3404 (N_3404,In_1046,In_831);
and U3405 (N_3405,In_3279,In_660);
and U3406 (N_3406,In_3786,In_1824);
or U3407 (N_3407,In_2382,In_3388);
xnor U3408 (N_3408,In_735,In_3676);
nor U3409 (N_3409,In_3784,In_2708);
xor U3410 (N_3410,In_2836,In_451);
and U3411 (N_3411,In_2340,In_2386);
nand U3412 (N_3412,In_1834,In_4377);
xor U3413 (N_3413,In_2035,In_3467);
nand U3414 (N_3414,In_1235,In_4050);
xor U3415 (N_3415,In_1372,In_2280);
nor U3416 (N_3416,In_949,In_2343);
xor U3417 (N_3417,In_646,In_3136);
or U3418 (N_3418,In_2242,In_1118);
xnor U3419 (N_3419,In_131,In_1088);
nand U3420 (N_3420,In_1143,In_1111);
and U3421 (N_3421,In_3379,In_2987);
or U3422 (N_3422,In_2308,In_4264);
or U3423 (N_3423,In_4523,In_4083);
and U3424 (N_3424,In_861,In_3737);
nor U3425 (N_3425,In_2583,In_2887);
and U3426 (N_3426,In_2810,In_2964);
nor U3427 (N_3427,In_3567,In_1207);
nand U3428 (N_3428,In_2794,In_3381);
nor U3429 (N_3429,In_3173,In_4809);
or U3430 (N_3430,In_1359,In_2306);
xnor U3431 (N_3431,In_42,In_3680);
nand U3432 (N_3432,In_2423,In_3879);
nor U3433 (N_3433,In_4212,In_3663);
and U3434 (N_3434,In_4667,In_571);
nand U3435 (N_3435,In_2829,In_1274);
xnor U3436 (N_3436,In_2687,In_4552);
nor U3437 (N_3437,In_4195,In_279);
xnor U3438 (N_3438,In_1761,In_3622);
or U3439 (N_3439,In_3200,In_1729);
nor U3440 (N_3440,In_3189,In_319);
or U3441 (N_3441,In_1007,In_4835);
nor U3442 (N_3442,In_3368,In_4179);
nand U3443 (N_3443,In_4804,In_2408);
nor U3444 (N_3444,In_3635,In_3682);
or U3445 (N_3445,In_4028,In_3346);
and U3446 (N_3446,In_2070,In_2895);
or U3447 (N_3447,In_1994,In_4602);
xnor U3448 (N_3448,In_553,In_1799);
xor U3449 (N_3449,In_3875,In_2417);
nor U3450 (N_3450,In_1797,In_665);
nand U3451 (N_3451,In_2225,In_657);
xnor U3452 (N_3452,In_3865,In_4004);
xor U3453 (N_3453,In_3637,In_1853);
and U3454 (N_3454,In_3260,In_3568);
nand U3455 (N_3455,In_4718,In_2145);
and U3456 (N_3456,In_4350,In_1298);
and U3457 (N_3457,In_526,In_2594);
xnor U3458 (N_3458,In_918,In_3659);
xor U3459 (N_3459,In_3553,In_4968);
nand U3460 (N_3460,In_3353,In_4104);
nand U3461 (N_3461,In_293,In_1331);
xnor U3462 (N_3462,In_929,In_43);
or U3463 (N_3463,In_2532,In_1402);
and U3464 (N_3464,In_4767,In_504);
nand U3465 (N_3465,In_4586,In_783);
and U3466 (N_3466,In_4551,In_267);
nor U3467 (N_3467,In_1348,In_1366);
xor U3468 (N_3468,In_2920,In_1637);
nand U3469 (N_3469,In_4177,In_1121);
xor U3470 (N_3470,In_3310,In_2713);
nor U3471 (N_3471,In_263,In_4079);
xor U3472 (N_3472,In_1741,In_415);
nor U3473 (N_3473,In_4407,In_3087);
and U3474 (N_3474,In_2413,In_3705);
nand U3475 (N_3475,In_2167,In_890);
and U3476 (N_3476,In_894,In_4524);
and U3477 (N_3477,In_1294,In_2895);
or U3478 (N_3478,In_1505,In_1856);
xnor U3479 (N_3479,In_2031,In_1668);
nor U3480 (N_3480,In_1096,In_3274);
xor U3481 (N_3481,In_4439,In_3365);
nand U3482 (N_3482,In_4043,In_2915);
or U3483 (N_3483,In_444,In_3355);
or U3484 (N_3484,In_3323,In_2459);
nand U3485 (N_3485,In_869,In_2153);
nor U3486 (N_3486,In_542,In_3251);
nor U3487 (N_3487,In_3318,In_1287);
or U3488 (N_3488,In_4363,In_998);
nor U3489 (N_3489,In_2188,In_3112);
xor U3490 (N_3490,In_3367,In_2337);
and U3491 (N_3491,In_3723,In_254);
xnor U3492 (N_3492,In_3011,In_2429);
nand U3493 (N_3493,In_2515,In_1332);
or U3494 (N_3494,In_4468,In_1711);
and U3495 (N_3495,In_1902,In_3126);
xor U3496 (N_3496,In_2354,In_3708);
xnor U3497 (N_3497,In_1734,In_2150);
nand U3498 (N_3498,In_4479,In_433);
or U3499 (N_3499,In_4741,In_1813);
xnor U3500 (N_3500,In_4588,In_3909);
or U3501 (N_3501,In_3343,In_1099);
nor U3502 (N_3502,In_2556,In_2619);
xor U3503 (N_3503,In_3989,In_2503);
nand U3504 (N_3504,In_4828,In_4476);
or U3505 (N_3505,In_4502,In_1596);
xnor U3506 (N_3506,In_991,In_4899);
and U3507 (N_3507,In_212,In_3585);
or U3508 (N_3508,In_430,In_4220);
xnor U3509 (N_3509,In_1929,In_1284);
nand U3510 (N_3510,In_4918,In_3616);
nor U3511 (N_3511,In_1401,In_1579);
nand U3512 (N_3512,In_2492,In_4104);
xor U3513 (N_3513,In_4136,In_3444);
and U3514 (N_3514,In_1885,In_4480);
xor U3515 (N_3515,In_2974,In_4405);
nor U3516 (N_3516,In_897,In_2546);
or U3517 (N_3517,In_1314,In_2025);
xor U3518 (N_3518,In_4352,In_632);
and U3519 (N_3519,In_1867,In_1044);
or U3520 (N_3520,In_1831,In_848);
or U3521 (N_3521,In_511,In_705);
xnor U3522 (N_3522,In_3759,In_4674);
xor U3523 (N_3523,In_4949,In_2022);
nor U3524 (N_3524,In_3919,In_784);
nand U3525 (N_3525,In_3217,In_3150);
and U3526 (N_3526,In_1134,In_3193);
nor U3527 (N_3527,In_4436,In_1068);
nand U3528 (N_3528,In_1433,In_1695);
nor U3529 (N_3529,In_4978,In_1734);
xnor U3530 (N_3530,In_689,In_3511);
or U3531 (N_3531,In_2772,In_2281);
nor U3532 (N_3532,In_2795,In_2245);
and U3533 (N_3533,In_1002,In_2530);
or U3534 (N_3534,In_2276,In_4029);
nor U3535 (N_3535,In_1142,In_2628);
nor U3536 (N_3536,In_1069,In_185);
nor U3537 (N_3537,In_4826,In_818);
nor U3538 (N_3538,In_89,In_1585);
nand U3539 (N_3539,In_2305,In_3187);
nand U3540 (N_3540,In_2668,In_3900);
nand U3541 (N_3541,In_763,In_785);
xnor U3542 (N_3542,In_2808,In_768);
nor U3543 (N_3543,In_4713,In_2990);
or U3544 (N_3544,In_2891,In_4739);
and U3545 (N_3545,In_71,In_1112);
nor U3546 (N_3546,In_3160,In_2150);
nor U3547 (N_3547,In_2615,In_3491);
or U3548 (N_3548,In_706,In_2049);
and U3549 (N_3549,In_4596,In_4211);
xnor U3550 (N_3550,In_4086,In_4537);
nand U3551 (N_3551,In_2731,In_1771);
nor U3552 (N_3552,In_2416,In_3090);
xnor U3553 (N_3553,In_4952,In_217);
or U3554 (N_3554,In_2608,In_3985);
or U3555 (N_3555,In_2858,In_2363);
and U3556 (N_3556,In_307,In_1319);
or U3557 (N_3557,In_2754,In_1692);
xor U3558 (N_3558,In_3359,In_3932);
or U3559 (N_3559,In_1435,In_3567);
and U3560 (N_3560,In_3520,In_4254);
or U3561 (N_3561,In_996,In_4143);
nor U3562 (N_3562,In_1742,In_4226);
nor U3563 (N_3563,In_2104,In_89);
nor U3564 (N_3564,In_323,In_4481);
and U3565 (N_3565,In_4054,In_4633);
nor U3566 (N_3566,In_1004,In_3856);
or U3567 (N_3567,In_341,In_679);
nand U3568 (N_3568,In_4486,In_4638);
xor U3569 (N_3569,In_4957,In_2996);
and U3570 (N_3570,In_4193,In_1618);
nand U3571 (N_3571,In_3563,In_4884);
and U3572 (N_3572,In_4052,In_1917);
or U3573 (N_3573,In_4880,In_2822);
and U3574 (N_3574,In_1433,In_2057);
xnor U3575 (N_3575,In_126,In_3754);
xor U3576 (N_3576,In_2526,In_4310);
nor U3577 (N_3577,In_2684,In_1725);
or U3578 (N_3578,In_2966,In_2008);
nand U3579 (N_3579,In_1812,In_2459);
nor U3580 (N_3580,In_3083,In_4590);
nand U3581 (N_3581,In_1085,In_3501);
and U3582 (N_3582,In_2138,In_4347);
nor U3583 (N_3583,In_2645,In_4738);
or U3584 (N_3584,In_3657,In_537);
or U3585 (N_3585,In_2684,In_1499);
or U3586 (N_3586,In_4453,In_1654);
and U3587 (N_3587,In_4164,In_1452);
nand U3588 (N_3588,In_1494,In_2732);
and U3589 (N_3589,In_1526,In_4528);
or U3590 (N_3590,In_3323,In_2201);
nand U3591 (N_3591,In_1576,In_609);
nand U3592 (N_3592,In_2773,In_2038);
or U3593 (N_3593,In_4473,In_1595);
nand U3594 (N_3594,In_1661,In_1428);
and U3595 (N_3595,In_2384,In_1127);
nor U3596 (N_3596,In_4937,In_4842);
xnor U3597 (N_3597,In_2782,In_2885);
nor U3598 (N_3598,In_2556,In_1988);
xor U3599 (N_3599,In_2442,In_621);
xor U3600 (N_3600,In_2049,In_4853);
or U3601 (N_3601,In_4787,In_606);
nor U3602 (N_3602,In_4073,In_992);
or U3603 (N_3603,In_1710,In_2833);
or U3604 (N_3604,In_1588,In_1768);
nand U3605 (N_3605,In_4621,In_778);
nor U3606 (N_3606,In_2931,In_1181);
or U3607 (N_3607,In_296,In_1900);
xnor U3608 (N_3608,In_4876,In_4465);
and U3609 (N_3609,In_4967,In_2724);
nand U3610 (N_3610,In_2270,In_3481);
and U3611 (N_3611,In_3082,In_2646);
nor U3612 (N_3612,In_4711,In_3956);
or U3613 (N_3613,In_1505,In_1025);
nand U3614 (N_3614,In_4050,In_1477);
or U3615 (N_3615,In_4474,In_1273);
nor U3616 (N_3616,In_3380,In_2157);
nor U3617 (N_3617,In_658,In_3988);
nor U3618 (N_3618,In_4746,In_4222);
xor U3619 (N_3619,In_4931,In_4312);
and U3620 (N_3620,In_1130,In_3376);
and U3621 (N_3621,In_1096,In_4222);
or U3622 (N_3622,In_1002,In_2236);
nor U3623 (N_3623,In_3071,In_1367);
xnor U3624 (N_3624,In_247,In_4853);
xor U3625 (N_3625,In_4252,In_382);
nor U3626 (N_3626,In_1347,In_241);
or U3627 (N_3627,In_2211,In_1399);
and U3628 (N_3628,In_3433,In_4090);
or U3629 (N_3629,In_4802,In_1353);
nand U3630 (N_3630,In_1440,In_1690);
nand U3631 (N_3631,In_3547,In_1271);
nor U3632 (N_3632,In_2088,In_1817);
nand U3633 (N_3633,In_4992,In_2068);
nor U3634 (N_3634,In_946,In_2780);
or U3635 (N_3635,In_2477,In_1514);
xor U3636 (N_3636,In_4090,In_1096);
xnor U3637 (N_3637,In_1410,In_2004);
xor U3638 (N_3638,In_1985,In_3960);
nand U3639 (N_3639,In_1523,In_1443);
nand U3640 (N_3640,In_3619,In_1976);
or U3641 (N_3641,In_2320,In_4120);
and U3642 (N_3642,In_210,In_3912);
or U3643 (N_3643,In_3939,In_1917);
and U3644 (N_3644,In_1873,In_1968);
nand U3645 (N_3645,In_3589,In_2926);
and U3646 (N_3646,In_3970,In_568);
and U3647 (N_3647,In_480,In_2106);
xnor U3648 (N_3648,In_1854,In_4626);
and U3649 (N_3649,In_4465,In_724);
xnor U3650 (N_3650,In_2718,In_3908);
or U3651 (N_3651,In_2907,In_3733);
nand U3652 (N_3652,In_235,In_4779);
nor U3653 (N_3653,In_3565,In_4510);
nor U3654 (N_3654,In_1533,In_1175);
nand U3655 (N_3655,In_3132,In_4806);
and U3656 (N_3656,In_4878,In_4985);
xnor U3657 (N_3657,In_4287,In_2589);
and U3658 (N_3658,In_4106,In_4303);
nand U3659 (N_3659,In_1228,In_4246);
or U3660 (N_3660,In_2485,In_157);
nor U3661 (N_3661,In_3372,In_4328);
nor U3662 (N_3662,In_1563,In_720);
or U3663 (N_3663,In_3710,In_2826);
and U3664 (N_3664,In_2645,In_1739);
xor U3665 (N_3665,In_1502,In_3277);
and U3666 (N_3666,In_1018,In_2042);
or U3667 (N_3667,In_1076,In_625);
nor U3668 (N_3668,In_2990,In_2503);
or U3669 (N_3669,In_1890,In_3853);
and U3670 (N_3670,In_2181,In_2702);
nor U3671 (N_3671,In_489,In_125);
or U3672 (N_3672,In_4085,In_2643);
xor U3673 (N_3673,In_2056,In_3039);
and U3674 (N_3674,In_996,In_2918);
nand U3675 (N_3675,In_3688,In_85);
or U3676 (N_3676,In_2873,In_1401);
nor U3677 (N_3677,In_4983,In_2386);
xor U3678 (N_3678,In_4187,In_1270);
xor U3679 (N_3679,In_416,In_3591);
nor U3680 (N_3680,In_1319,In_3764);
xnor U3681 (N_3681,In_1007,In_1662);
nand U3682 (N_3682,In_4401,In_1873);
nand U3683 (N_3683,In_903,In_2559);
and U3684 (N_3684,In_3513,In_1829);
and U3685 (N_3685,In_696,In_1993);
and U3686 (N_3686,In_1248,In_4013);
xnor U3687 (N_3687,In_3979,In_3311);
nand U3688 (N_3688,In_4436,In_1110);
xor U3689 (N_3689,In_4031,In_1931);
or U3690 (N_3690,In_3957,In_1916);
or U3691 (N_3691,In_1525,In_791);
nand U3692 (N_3692,In_2883,In_1039);
or U3693 (N_3693,In_2045,In_1408);
nor U3694 (N_3694,In_1633,In_3589);
nor U3695 (N_3695,In_2061,In_2758);
or U3696 (N_3696,In_2787,In_2818);
nor U3697 (N_3697,In_3282,In_4354);
or U3698 (N_3698,In_2690,In_4430);
xnor U3699 (N_3699,In_2840,In_534);
or U3700 (N_3700,In_4464,In_2818);
and U3701 (N_3701,In_4212,In_641);
nand U3702 (N_3702,In_1816,In_2389);
or U3703 (N_3703,In_2946,In_1574);
or U3704 (N_3704,In_3884,In_3358);
nand U3705 (N_3705,In_523,In_1229);
xor U3706 (N_3706,In_83,In_3613);
nand U3707 (N_3707,In_1430,In_3776);
nand U3708 (N_3708,In_3600,In_3088);
or U3709 (N_3709,In_4226,In_4679);
or U3710 (N_3710,In_4503,In_2450);
xor U3711 (N_3711,In_2644,In_364);
xor U3712 (N_3712,In_1006,In_3287);
nor U3713 (N_3713,In_1480,In_1065);
nor U3714 (N_3714,In_2401,In_1546);
nor U3715 (N_3715,In_4886,In_4444);
xnor U3716 (N_3716,In_1792,In_4906);
or U3717 (N_3717,In_63,In_4528);
or U3718 (N_3718,In_3679,In_4922);
nand U3719 (N_3719,In_576,In_2510);
or U3720 (N_3720,In_3685,In_2238);
xnor U3721 (N_3721,In_85,In_3198);
xor U3722 (N_3722,In_3631,In_4096);
nor U3723 (N_3723,In_615,In_1241);
xor U3724 (N_3724,In_2598,In_2132);
xor U3725 (N_3725,In_4444,In_3090);
and U3726 (N_3726,In_2541,In_451);
xor U3727 (N_3727,In_1200,In_4059);
or U3728 (N_3728,In_4098,In_4062);
nand U3729 (N_3729,In_3974,In_2247);
nor U3730 (N_3730,In_2238,In_1373);
nor U3731 (N_3731,In_1557,In_4169);
xnor U3732 (N_3732,In_120,In_1076);
and U3733 (N_3733,In_659,In_1130);
xor U3734 (N_3734,In_3859,In_3661);
nor U3735 (N_3735,In_3860,In_1136);
and U3736 (N_3736,In_2305,In_687);
or U3737 (N_3737,In_1698,In_471);
nand U3738 (N_3738,In_1818,In_4962);
nand U3739 (N_3739,In_1006,In_4948);
and U3740 (N_3740,In_2049,In_36);
xnor U3741 (N_3741,In_84,In_937);
xor U3742 (N_3742,In_935,In_3387);
or U3743 (N_3743,In_4384,In_788);
and U3744 (N_3744,In_3341,In_2758);
xnor U3745 (N_3745,In_4300,In_1902);
xnor U3746 (N_3746,In_3136,In_571);
or U3747 (N_3747,In_2277,In_1275);
xnor U3748 (N_3748,In_3439,In_3115);
xor U3749 (N_3749,In_3273,In_2649);
nor U3750 (N_3750,In_3559,In_2858);
xor U3751 (N_3751,In_1289,In_4016);
nand U3752 (N_3752,In_736,In_2420);
or U3753 (N_3753,In_17,In_3293);
xor U3754 (N_3754,In_4348,In_2413);
xnor U3755 (N_3755,In_2987,In_708);
and U3756 (N_3756,In_1719,In_2959);
xnor U3757 (N_3757,In_3441,In_4899);
xnor U3758 (N_3758,In_4267,In_3916);
nor U3759 (N_3759,In_4904,In_2860);
xor U3760 (N_3760,In_163,In_2486);
and U3761 (N_3761,In_4090,In_1352);
and U3762 (N_3762,In_982,In_1875);
nor U3763 (N_3763,In_3564,In_3313);
and U3764 (N_3764,In_1735,In_3212);
nand U3765 (N_3765,In_2587,In_1624);
or U3766 (N_3766,In_1635,In_2112);
or U3767 (N_3767,In_4519,In_2338);
xnor U3768 (N_3768,In_186,In_2386);
and U3769 (N_3769,In_3296,In_4726);
xnor U3770 (N_3770,In_4615,In_4739);
nor U3771 (N_3771,In_4209,In_2468);
and U3772 (N_3772,In_2040,In_2036);
xnor U3773 (N_3773,In_3921,In_2815);
or U3774 (N_3774,In_1998,In_4978);
nand U3775 (N_3775,In_1585,In_1175);
or U3776 (N_3776,In_2259,In_1838);
xor U3777 (N_3777,In_2618,In_3459);
xor U3778 (N_3778,In_518,In_4485);
nor U3779 (N_3779,In_1632,In_1813);
or U3780 (N_3780,In_3084,In_4501);
nand U3781 (N_3781,In_4639,In_2818);
and U3782 (N_3782,In_2682,In_4930);
nor U3783 (N_3783,In_4309,In_3743);
or U3784 (N_3784,In_3604,In_4469);
and U3785 (N_3785,In_4268,In_3196);
xnor U3786 (N_3786,In_2285,In_2970);
and U3787 (N_3787,In_3086,In_4423);
nand U3788 (N_3788,In_4367,In_583);
nor U3789 (N_3789,In_2800,In_3063);
or U3790 (N_3790,In_1077,In_119);
xnor U3791 (N_3791,In_2543,In_1128);
and U3792 (N_3792,In_1593,In_2837);
nand U3793 (N_3793,In_4689,In_2854);
nor U3794 (N_3794,In_4076,In_3428);
or U3795 (N_3795,In_3269,In_49);
nor U3796 (N_3796,In_189,In_150);
and U3797 (N_3797,In_807,In_4448);
or U3798 (N_3798,In_895,In_3238);
and U3799 (N_3799,In_1453,In_2057);
nor U3800 (N_3800,In_2693,In_3023);
and U3801 (N_3801,In_1307,In_4191);
or U3802 (N_3802,In_1819,In_4057);
or U3803 (N_3803,In_1484,In_1340);
nand U3804 (N_3804,In_3945,In_2244);
nand U3805 (N_3805,In_2459,In_4947);
xnor U3806 (N_3806,In_2884,In_4351);
nor U3807 (N_3807,In_1484,In_4455);
xor U3808 (N_3808,In_1182,In_1550);
or U3809 (N_3809,In_3906,In_1681);
or U3810 (N_3810,In_4302,In_2845);
nand U3811 (N_3811,In_3099,In_3608);
nor U3812 (N_3812,In_2666,In_4394);
nand U3813 (N_3813,In_3945,In_2268);
and U3814 (N_3814,In_1658,In_2107);
nor U3815 (N_3815,In_2836,In_2745);
or U3816 (N_3816,In_3217,In_2199);
or U3817 (N_3817,In_564,In_122);
and U3818 (N_3818,In_4617,In_4129);
and U3819 (N_3819,In_840,In_2549);
and U3820 (N_3820,In_4992,In_3585);
or U3821 (N_3821,In_2585,In_2271);
and U3822 (N_3822,In_1994,In_1424);
nor U3823 (N_3823,In_61,In_701);
and U3824 (N_3824,In_4153,In_3708);
nor U3825 (N_3825,In_439,In_1696);
nand U3826 (N_3826,In_4480,In_3019);
or U3827 (N_3827,In_2402,In_3076);
nand U3828 (N_3828,In_1508,In_4266);
xor U3829 (N_3829,In_288,In_68);
and U3830 (N_3830,In_1264,In_1401);
nor U3831 (N_3831,In_1125,In_2349);
nand U3832 (N_3832,In_1200,In_426);
nor U3833 (N_3833,In_4885,In_2956);
xor U3834 (N_3834,In_3610,In_1199);
or U3835 (N_3835,In_90,In_2524);
nor U3836 (N_3836,In_587,In_806);
and U3837 (N_3837,In_2316,In_279);
nand U3838 (N_3838,In_3350,In_6);
or U3839 (N_3839,In_4351,In_3501);
nor U3840 (N_3840,In_3894,In_216);
or U3841 (N_3841,In_413,In_4032);
and U3842 (N_3842,In_4738,In_2913);
or U3843 (N_3843,In_4778,In_2078);
nand U3844 (N_3844,In_1890,In_403);
nand U3845 (N_3845,In_2953,In_4745);
and U3846 (N_3846,In_817,In_602);
and U3847 (N_3847,In_310,In_4172);
xnor U3848 (N_3848,In_362,In_4617);
xor U3849 (N_3849,In_913,In_3416);
nor U3850 (N_3850,In_3726,In_3356);
nor U3851 (N_3851,In_4761,In_3073);
nor U3852 (N_3852,In_3219,In_3743);
nor U3853 (N_3853,In_3875,In_2540);
nor U3854 (N_3854,In_2333,In_1675);
and U3855 (N_3855,In_3540,In_933);
xor U3856 (N_3856,In_2601,In_4499);
and U3857 (N_3857,In_2713,In_3674);
and U3858 (N_3858,In_3196,In_507);
nor U3859 (N_3859,In_3207,In_447);
nand U3860 (N_3860,In_2674,In_1968);
or U3861 (N_3861,In_589,In_852);
nor U3862 (N_3862,In_1982,In_4931);
and U3863 (N_3863,In_1275,In_494);
nor U3864 (N_3864,In_2996,In_3265);
nand U3865 (N_3865,In_1945,In_631);
xnor U3866 (N_3866,In_2349,In_3843);
and U3867 (N_3867,In_1458,In_658);
xor U3868 (N_3868,In_2686,In_2997);
xnor U3869 (N_3869,In_4653,In_1907);
and U3870 (N_3870,In_1946,In_3550);
nor U3871 (N_3871,In_911,In_2193);
nand U3872 (N_3872,In_4587,In_711);
and U3873 (N_3873,In_1748,In_1144);
nor U3874 (N_3874,In_3847,In_2632);
nand U3875 (N_3875,In_4739,In_1096);
nor U3876 (N_3876,In_4951,In_575);
nor U3877 (N_3877,In_4874,In_4842);
nand U3878 (N_3878,In_395,In_4621);
nor U3879 (N_3879,In_1360,In_2810);
xor U3880 (N_3880,In_1137,In_4883);
and U3881 (N_3881,In_3534,In_2419);
and U3882 (N_3882,In_1946,In_1515);
or U3883 (N_3883,In_901,In_4230);
nor U3884 (N_3884,In_1147,In_1184);
nand U3885 (N_3885,In_1802,In_2782);
xnor U3886 (N_3886,In_4003,In_2267);
nand U3887 (N_3887,In_1191,In_631);
or U3888 (N_3888,In_3851,In_1262);
xor U3889 (N_3889,In_3786,In_2122);
xnor U3890 (N_3890,In_4126,In_1561);
nand U3891 (N_3891,In_2538,In_3339);
or U3892 (N_3892,In_3011,In_3915);
and U3893 (N_3893,In_2543,In_3614);
or U3894 (N_3894,In_556,In_3655);
nor U3895 (N_3895,In_4878,In_1441);
nand U3896 (N_3896,In_3780,In_3486);
or U3897 (N_3897,In_2902,In_1047);
nand U3898 (N_3898,In_2025,In_3353);
or U3899 (N_3899,In_1661,In_62);
xnor U3900 (N_3900,In_2646,In_1418);
nor U3901 (N_3901,In_2394,In_1782);
nor U3902 (N_3902,In_4811,In_2763);
and U3903 (N_3903,In_1010,In_2505);
nor U3904 (N_3904,In_1502,In_2871);
nor U3905 (N_3905,In_634,In_479);
nor U3906 (N_3906,In_716,In_795);
and U3907 (N_3907,In_2036,In_2515);
and U3908 (N_3908,In_1239,In_3252);
and U3909 (N_3909,In_190,In_3307);
and U3910 (N_3910,In_1513,In_4528);
or U3911 (N_3911,In_1607,In_1718);
nor U3912 (N_3912,In_4217,In_1679);
nand U3913 (N_3913,In_3589,In_3478);
or U3914 (N_3914,In_3006,In_38);
nor U3915 (N_3915,In_1765,In_4830);
nor U3916 (N_3916,In_2742,In_1451);
and U3917 (N_3917,In_3824,In_1519);
nand U3918 (N_3918,In_4491,In_1465);
nor U3919 (N_3919,In_1295,In_1781);
nor U3920 (N_3920,In_4202,In_1572);
xor U3921 (N_3921,In_1858,In_4605);
nor U3922 (N_3922,In_4969,In_3708);
or U3923 (N_3923,In_1121,In_4139);
or U3924 (N_3924,In_2919,In_4125);
or U3925 (N_3925,In_1534,In_3676);
nand U3926 (N_3926,In_1899,In_1500);
or U3927 (N_3927,In_4518,In_4222);
nand U3928 (N_3928,In_1532,In_1153);
xnor U3929 (N_3929,In_1697,In_4170);
and U3930 (N_3930,In_4459,In_2590);
or U3931 (N_3931,In_4897,In_4638);
xor U3932 (N_3932,In_4355,In_2315);
and U3933 (N_3933,In_3567,In_1411);
nor U3934 (N_3934,In_2787,In_2761);
and U3935 (N_3935,In_1322,In_2584);
and U3936 (N_3936,In_3348,In_2743);
or U3937 (N_3937,In_2548,In_895);
xnor U3938 (N_3938,In_3821,In_1474);
nand U3939 (N_3939,In_2349,In_753);
nor U3940 (N_3940,In_4133,In_3434);
nor U3941 (N_3941,In_1911,In_1325);
nand U3942 (N_3942,In_3395,In_10);
nor U3943 (N_3943,In_523,In_974);
nor U3944 (N_3944,In_2031,In_105);
or U3945 (N_3945,In_18,In_2585);
nand U3946 (N_3946,In_4272,In_90);
xor U3947 (N_3947,In_801,In_2278);
or U3948 (N_3948,In_2377,In_2429);
or U3949 (N_3949,In_2889,In_1567);
nand U3950 (N_3950,In_1211,In_850);
xor U3951 (N_3951,In_3480,In_4368);
or U3952 (N_3952,In_1116,In_1502);
nor U3953 (N_3953,In_3124,In_2986);
nand U3954 (N_3954,In_2340,In_4940);
nand U3955 (N_3955,In_4106,In_4651);
nand U3956 (N_3956,In_4474,In_3507);
and U3957 (N_3957,In_323,In_1038);
and U3958 (N_3958,In_4884,In_3615);
and U3959 (N_3959,In_4765,In_2984);
nor U3960 (N_3960,In_871,In_4438);
nand U3961 (N_3961,In_1093,In_3334);
and U3962 (N_3962,In_1167,In_4435);
xor U3963 (N_3963,In_166,In_2378);
xnor U3964 (N_3964,In_2556,In_2578);
or U3965 (N_3965,In_1292,In_971);
and U3966 (N_3966,In_4178,In_4632);
xor U3967 (N_3967,In_3791,In_2835);
and U3968 (N_3968,In_1465,In_612);
xnor U3969 (N_3969,In_3405,In_3623);
xor U3970 (N_3970,In_717,In_405);
and U3971 (N_3971,In_4066,In_3667);
nor U3972 (N_3972,In_2640,In_2802);
or U3973 (N_3973,In_2065,In_382);
nand U3974 (N_3974,In_2348,In_646);
or U3975 (N_3975,In_3139,In_4442);
and U3976 (N_3976,In_2965,In_4463);
and U3977 (N_3977,In_1161,In_4032);
nor U3978 (N_3978,In_891,In_4441);
xnor U3979 (N_3979,In_4862,In_626);
nand U3980 (N_3980,In_3821,In_4904);
nor U3981 (N_3981,In_3723,In_2711);
or U3982 (N_3982,In_4879,In_1418);
or U3983 (N_3983,In_3499,In_4318);
nand U3984 (N_3984,In_3273,In_3865);
and U3985 (N_3985,In_2640,In_1536);
nand U3986 (N_3986,In_4180,In_575);
nor U3987 (N_3987,In_1735,In_2532);
and U3988 (N_3988,In_2881,In_4639);
nor U3989 (N_3989,In_1226,In_881);
nor U3990 (N_3990,In_1064,In_4067);
and U3991 (N_3991,In_2947,In_77);
or U3992 (N_3992,In_772,In_2025);
xnor U3993 (N_3993,In_3534,In_726);
and U3994 (N_3994,In_162,In_1594);
nand U3995 (N_3995,In_4600,In_2683);
nand U3996 (N_3996,In_960,In_4158);
xor U3997 (N_3997,In_596,In_4429);
nor U3998 (N_3998,In_1390,In_4046);
nor U3999 (N_3999,In_4664,In_3788);
xor U4000 (N_4000,In_1060,In_3627);
or U4001 (N_4001,In_1452,In_2671);
and U4002 (N_4002,In_2565,In_4905);
or U4003 (N_4003,In_1918,In_819);
and U4004 (N_4004,In_4523,In_662);
nor U4005 (N_4005,In_770,In_1209);
nor U4006 (N_4006,In_2865,In_2143);
and U4007 (N_4007,In_4943,In_245);
and U4008 (N_4008,In_227,In_1580);
and U4009 (N_4009,In_1128,In_2135);
xor U4010 (N_4010,In_2651,In_1870);
nand U4011 (N_4011,In_2374,In_3438);
nor U4012 (N_4012,In_1035,In_4989);
nor U4013 (N_4013,In_3160,In_2955);
xor U4014 (N_4014,In_48,In_1804);
nor U4015 (N_4015,In_4634,In_4368);
xnor U4016 (N_4016,In_3713,In_3278);
or U4017 (N_4017,In_3786,In_1221);
and U4018 (N_4018,In_1860,In_4728);
xnor U4019 (N_4019,In_433,In_1754);
and U4020 (N_4020,In_4786,In_3565);
xor U4021 (N_4021,In_4600,In_1792);
or U4022 (N_4022,In_3965,In_1410);
or U4023 (N_4023,In_2622,In_3018);
xnor U4024 (N_4024,In_4199,In_4985);
nor U4025 (N_4025,In_2219,In_4215);
xor U4026 (N_4026,In_4132,In_2343);
xor U4027 (N_4027,In_4349,In_3390);
nor U4028 (N_4028,In_2841,In_2412);
or U4029 (N_4029,In_359,In_4718);
xnor U4030 (N_4030,In_4260,In_4671);
nor U4031 (N_4031,In_3301,In_3107);
nor U4032 (N_4032,In_2589,In_793);
nand U4033 (N_4033,In_2934,In_2834);
nor U4034 (N_4034,In_1202,In_2669);
or U4035 (N_4035,In_1088,In_3174);
and U4036 (N_4036,In_711,In_4690);
nor U4037 (N_4037,In_2172,In_3033);
xor U4038 (N_4038,In_2587,In_655);
nor U4039 (N_4039,In_1792,In_2419);
nor U4040 (N_4040,In_2970,In_586);
xor U4041 (N_4041,In_2594,In_2914);
nand U4042 (N_4042,In_2021,In_2094);
nand U4043 (N_4043,In_1187,In_3848);
nand U4044 (N_4044,In_2686,In_1507);
or U4045 (N_4045,In_4353,In_3868);
nand U4046 (N_4046,In_4993,In_3804);
xor U4047 (N_4047,In_1824,In_418);
and U4048 (N_4048,In_3954,In_72);
xor U4049 (N_4049,In_4832,In_1887);
and U4050 (N_4050,In_1655,In_4222);
nor U4051 (N_4051,In_3020,In_1125);
xor U4052 (N_4052,In_4593,In_1584);
xnor U4053 (N_4053,In_3474,In_3473);
nand U4054 (N_4054,In_1656,In_351);
nand U4055 (N_4055,In_1597,In_463);
nand U4056 (N_4056,In_502,In_4314);
nand U4057 (N_4057,In_865,In_1402);
nand U4058 (N_4058,In_822,In_3035);
or U4059 (N_4059,In_1564,In_3196);
or U4060 (N_4060,In_2554,In_2905);
xor U4061 (N_4061,In_2093,In_2191);
or U4062 (N_4062,In_2241,In_4351);
nor U4063 (N_4063,In_392,In_548);
xor U4064 (N_4064,In_723,In_2326);
nand U4065 (N_4065,In_1006,In_2863);
nand U4066 (N_4066,In_1436,In_383);
or U4067 (N_4067,In_3006,In_650);
xnor U4068 (N_4068,In_221,In_4949);
and U4069 (N_4069,In_4432,In_4176);
or U4070 (N_4070,In_3756,In_1955);
or U4071 (N_4071,In_4325,In_3477);
or U4072 (N_4072,In_2728,In_1963);
nand U4073 (N_4073,In_1025,In_2667);
and U4074 (N_4074,In_1416,In_290);
and U4075 (N_4075,In_4801,In_2090);
or U4076 (N_4076,In_3545,In_268);
or U4077 (N_4077,In_2343,In_389);
nand U4078 (N_4078,In_4963,In_4692);
nor U4079 (N_4079,In_1575,In_3095);
nand U4080 (N_4080,In_1602,In_1233);
nor U4081 (N_4081,In_402,In_1277);
and U4082 (N_4082,In_4168,In_2805);
nand U4083 (N_4083,In_4687,In_76);
or U4084 (N_4084,In_1086,In_4221);
xnor U4085 (N_4085,In_3435,In_791);
xor U4086 (N_4086,In_3757,In_4047);
and U4087 (N_4087,In_1933,In_3487);
xor U4088 (N_4088,In_533,In_2053);
or U4089 (N_4089,In_3363,In_1251);
or U4090 (N_4090,In_741,In_3276);
nand U4091 (N_4091,In_2966,In_3125);
and U4092 (N_4092,In_2442,In_120);
xnor U4093 (N_4093,In_4074,In_4462);
nor U4094 (N_4094,In_4023,In_234);
or U4095 (N_4095,In_4100,In_1743);
nand U4096 (N_4096,In_4511,In_1052);
and U4097 (N_4097,In_1734,In_1453);
nor U4098 (N_4098,In_10,In_2072);
nand U4099 (N_4099,In_242,In_3837);
and U4100 (N_4100,In_927,In_4056);
or U4101 (N_4101,In_61,In_472);
and U4102 (N_4102,In_1216,In_353);
and U4103 (N_4103,In_4153,In_2602);
xnor U4104 (N_4104,In_4628,In_2790);
or U4105 (N_4105,In_707,In_641);
nand U4106 (N_4106,In_903,In_4533);
and U4107 (N_4107,In_2517,In_4427);
and U4108 (N_4108,In_2074,In_223);
or U4109 (N_4109,In_2079,In_274);
nor U4110 (N_4110,In_2314,In_576);
xor U4111 (N_4111,In_4798,In_4137);
xnor U4112 (N_4112,In_2594,In_3089);
xor U4113 (N_4113,In_2783,In_1618);
xnor U4114 (N_4114,In_422,In_1975);
nor U4115 (N_4115,In_2215,In_604);
and U4116 (N_4116,In_577,In_934);
xnor U4117 (N_4117,In_506,In_1297);
xnor U4118 (N_4118,In_44,In_3687);
and U4119 (N_4119,In_3036,In_3880);
and U4120 (N_4120,In_2871,In_3000);
nand U4121 (N_4121,In_259,In_2674);
xor U4122 (N_4122,In_2852,In_3067);
nand U4123 (N_4123,In_980,In_4202);
nand U4124 (N_4124,In_142,In_2006);
nor U4125 (N_4125,In_4377,In_1875);
and U4126 (N_4126,In_1947,In_865);
xor U4127 (N_4127,In_4072,In_2572);
or U4128 (N_4128,In_2948,In_1935);
nor U4129 (N_4129,In_2759,In_4132);
xnor U4130 (N_4130,In_565,In_1813);
nor U4131 (N_4131,In_2781,In_957);
or U4132 (N_4132,In_1932,In_1268);
xnor U4133 (N_4133,In_2677,In_1664);
or U4134 (N_4134,In_201,In_3168);
nor U4135 (N_4135,In_2859,In_1507);
nand U4136 (N_4136,In_1600,In_1269);
or U4137 (N_4137,In_2638,In_1984);
and U4138 (N_4138,In_1018,In_2872);
nor U4139 (N_4139,In_527,In_3115);
xor U4140 (N_4140,In_731,In_4722);
xor U4141 (N_4141,In_4834,In_3798);
or U4142 (N_4142,In_1446,In_1676);
or U4143 (N_4143,In_4500,In_3645);
nor U4144 (N_4144,In_830,In_2290);
nor U4145 (N_4145,In_3325,In_2180);
and U4146 (N_4146,In_3283,In_4093);
xor U4147 (N_4147,In_4561,In_103);
or U4148 (N_4148,In_1250,In_403);
and U4149 (N_4149,In_4039,In_84);
and U4150 (N_4150,In_2794,In_3843);
nand U4151 (N_4151,In_962,In_1251);
or U4152 (N_4152,In_2574,In_4530);
and U4153 (N_4153,In_47,In_3554);
xor U4154 (N_4154,In_3326,In_15);
nand U4155 (N_4155,In_4255,In_409);
or U4156 (N_4156,In_1284,In_4517);
and U4157 (N_4157,In_4612,In_4482);
nor U4158 (N_4158,In_1088,In_4711);
or U4159 (N_4159,In_1810,In_581);
and U4160 (N_4160,In_1468,In_1522);
and U4161 (N_4161,In_822,In_3667);
or U4162 (N_4162,In_2733,In_4723);
nor U4163 (N_4163,In_1348,In_4630);
nand U4164 (N_4164,In_3490,In_4910);
and U4165 (N_4165,In_2865,In_1763);
or U4166 (N_4166,In_4609,In_4570);
nand U4167 (N_4167,In_571,In_1911);
and U4168 (N_4168,In_3333,In_1682);
or U4169 (N_4169,In_681,In_3507);
and U4170 (N_4170,In_803,In_3147);
or U4171 (N_4171,In_531,In_214);
nor U4172 (N_4172,In_1722,In_1558);
xor U4173 (N_4173,In_169,In_1701);
xor U4174 (N_4174,In_2205,In_4481);
and U4175 (N_4175,In_3697,In_4861);
nor U4176 (N_4176,In_4247,In_3957);
nand U4177 (N_4177,In_410,In_4696);
nor U4178 (N_4178,In_1750,In_4759);
and U4179 (N_4179,In_4675,In_26);
nand U4180 (N_4180,In_2961,In_2054);
or U4181 (N_4181,In_1272,In_3105);
nor U4182 (N_4182,In_1323,In_2442);
xor U4183 (N_4183,In_642,In_1472);
xor U4184 (N_4184,In_1916,In_4584);
nand U4185 (N_4185,In_2034,In_3211);
xnor U4186 (N_4186,In_3518,In_3549);
and U4187 (N_4187,In_4301,In_1684);
nor U4188 (N_4188,In_2458,In_1764);
or U4189 (N_4189,In_1353,In_3181);
nand U4190 (N_4190,In_2549,In_1664);
or U4191 (N_4191,In_946,In_4544);
nor U4192 (N_4192,In_1022,In_719);
or U4193 (N_4193,In_4009,In_775);
xnor U4194 (N_4194,In_4956,In_1972);
nor U4195 (N_4195,In_1993,In_2256);
xor U4196 (N_4196,In_3882,In_3690);
and U4197 (N_4197,In_1164,In_4135);
and U4198 (N_4198,In_3367,In_2583);
nand U4199 (N_4199,In_4399,In_2543);
and U4200 (N_4200,In_4260,In_2399);
nor U4201 (N_4201,In_4909,In_639);
nor U4202 (N_4202,In_1853,In_1551);
or U4203 (N_4203,In_2884,In_1967);
xnor U4204 (N_4204,In_4434,In_3884);
and U4205 (N_4205,In_3638,In_969);
and U4206 (N_4206,In_3685,In_550);
nor U4207 (N_4207,In_676,In_3676);
and U4208 (N_4208,In_4352,In_4976);
or U4209 (N_4209,In_1474,In_2286);
nand U4210 (N_4210,In_4479,In_845);
xnor U4211 (N_4211,In_4210,In_4461);
nand U4212 (N_4212,In_33,In_1767);
xnor U4213 (N_4213,In_4575,In_2897);
or U4214 (N_4214,In_2204,In_3431);
nor U4215 (N_4215,In_1007,In_2016);
and U4216 (N_4216,In_2776,In_97);
or U4217 (N_4217,In_711,In_4769);
nand U4218 (N_4218,In_4598,In_3595);
xnor U4219 (N_4219,In_4356,In_2611);
and U4220 (N_4220,In_4905,In_4474);
nand U4221 (N_4221,In_4941,In_144);
nor U4222 (N_4222,In_636,In_759);
nand U4223 (N_4223,In_4326,In_4178);
and U4224 (N_4224,In_4757,In_2147);
nand U4225 (N_4225,In_1667,In_2291);
xnor U4226 (N_4226,In_3360,In_4265);
nor U4227 (N_4227,In_4775,In_1072);
nand U4228 (N_4228,In_1714,In_3964);
nor U4229 (N_4229,In_3527,In_1458);
xnor U4230 (N_4230,In_640,In_3835);
nor U4231 (N_4231,In_1840,In_2476);
or U4232 (N_4232,In_4968,In_2546);
and U4233 (N_4233,In_3808,In_1620);
and U4234 (N_4234,In_2706,In_3831);
nand U4235 (N_4235,In_3795,In_4364);
nor U4236 (N_4236,In_3273,In_1330);
nor U4237 (N_4237,In_2683,In_932);
nor U4238 (N_4238,In_1196,In_3713);
and U4239 (N_4239,In_1212,In_4339);
nor U4240 (N_4240,In_485,In_1284);
nand U4241 (N_4241,In_2676,In_3043);
or U4242 (N_4242,In_469,In_4945);
xor U4243 (N_4243,In_691,In_2918);
or U4244 (N_4244,In_3146,In_1171);
nand U4245 (N_4245,In_2227,In_3099);
and U4246 (N_4246,In_1315,In_4291);
nor U4247 (N_4247,In_4154,In_3482);
and U4248 (N_4248,In_899,In_2667);
nor U4249 (N_4249,In_1435,In_4251);
nor U4250 (N_4250,In_4862,In_2734);
and U4251 (N_4251,In_3179,In_1978);
and U4252 (N_4252,In_2745,In_1864);
or U4253 (N_4253,In_3321,In_3073);
and U4254 (N_4254,In_1239,In_661);
xnor U4255 (N_4255,In_3012,In_4027);
nand U4256 (N_4256,In_1937,In_1036);
nor U4257 (N_4257,In_4476,In_4833);
or U4258 (N_4258,In_2515,In_3214);
xor U4259 (N_4259,In_536,In_1516);
and U4260 (N_4260,In_3303,In_2616);
and U4261 (N_4261,In_1500,In_2508);
or U4262 (N_4262,In_3298,In_2669);
nor U4263 (N_4263,In_3176,In_1625);
nand U4264 (N_4264,In_4918,In_2812);
and U4265 (N_4265,In_1109,In_993);
nand U4266 (N_4266,In_2247,In_4955);
xnor U4267 (N_4267,In_1092,In_1759);
or U4268 (N_4268,In_2054,In_4552);
xnor U4269 (N_4269,In_3826,In_4354);
or U4270 (N_4270,In_4873,In_3622);
nor U4271 (N_4271,In_4313,In_88);
nand U4272 (N_4272,In_103,In_108);
nor U4273 (N_4273,In_560,In_4352);
or U4274 (N_4274,In_3544,In_3206);
nor U4275 (N_4275,In_3841,In_1568);
nand U4276 (N_4276,In_181,In_3167);
and U4277 (N_4277,In_2176,In_4814);
and U4278 (N_4278,In_3305,In_641);
or U4279 (N_4279,In_120,In_2952);
nor U4280 (N_4280,In_2995,In_4123);
nand U4281 (N_4281,In_760,In_1811);
xor U4282 (N_4282,In_2140,In_1212);
nor U4283 (N_4283,In_4378,In_2786);
xnor U4284 (N_4284,In_428,In_4985);
nand U4285 (N_4285,In_877,In_87);
nor U4286 (N_4286,In_4906,In_1562);
xnor U4287 (N_4287,In_4155,In_50);
nor U4288 (N_4288,In_1369,In_3341);
xor U4289 (N_4289,In_3171,In_1568);
nor U4290 (N_4290,In_4205,In_1847);
and U4291 (N_4291,In_1180,In_1829);
and U4292 (N_4292,In_2267,In_4797);
nor U4293 (N_4293,In_451,In_559);
nor U4294 (N_4294,In_4474,In_1246);
nor U4295 (N_4295,In_3529,In_4397);
and U4296 (N_4296,In_511,In_243);
nand U4297 (N_4297,In_4172,In_1312);
nor U4298 (N_4298,In_541,In_3391);
and U4299 (N_4299,In_3223,In_110);
or U4300 (N_4300,In_2062,In_2894);
xnor U4301 (N_4301,In_3840,In_4886);
and U4302 (N_4302,In_2923,In_4837);
or U4303 (N_4303,In_4476,In_4384);
nand U4304 (N_4304,In_1232,In_2044);
nand U4305 (N_4305,In_3393,In_3163);
nand U4306 (N_4306,In_3544,In_248);
nor U4307 (N_4307,In_1083,In_1585);
nor U4308 (N_4308,In_895,In_2011);
nor U4309 (N_4309,In_2214,In_3862);
and U4310 (N_4310,In_3196,In_3922);
nand U4311 (N_4311,In_237,In_4270);
and U4312 (N_4312,In_1150,In_4615);
or U4313 (N_4313,In_3410,In_59);
xnor U4314 (N_4314,In_4605,In_1198);
or U4315 (N_4315,In_2754,In_2646);
xnor U4316 (N_4316,In_3005,In_2562);
nand U4317 (N_4317,In_4289,In_4330);
and U4318 (N_4318,In_3086,In_1379);
nand U4319 (N_4319,In_875,In_2183);
or U4320 (N_4320,In_1776,In_3115);
nor U4321 (N_4321,In_4510,In_2414);
xnor U4322 (N_4322,In_4381,In_3482);
nor U4323 (N_4323,In_1400,In_2503);
and U4324 (N_4324,In_2176,In_1006);
nor U4325 (N_4325,In_4195,In_3433);
xnor U4326 (N_4326,In_4468,In_885);
or U4327 (N_4327,In_2924,In_3517);
or U4328 (N_4328,In_804,In_611);
nand U4329 (N_4329,In_3511,In_3853);
or U4330 (N_4330,In_2265,In_4948);
or U4331 (N_4331,In_305,In_216);
or U4332 (N_4332,In_3905,In_4589);
nor U4333 (N_4333,In_2076,In_1642);
xnor U4334 (N_4334,In_1369,In_2303);
nor U4335 (N_4335,In_1653,In_2041);
xnor U4336 (N_4336,In_2845,In_2067);
nor U4337 (N_4337,In_4759,In_4172);
nand U4338 (N_4338,In_2863,In_3652);
nand U4339 (N_4339,In_4158,In_3653);
or U4340 (N_4340,In_2406,In_4361);
xor U4341 (N_4341,In_771,In_3408);
xnor U4342 (N_4342,In_2162,In_2387);
xnor U4343 (N_4343,In_284,In_451);
xnor U4344 (N_4344,In_1249,In_867);
or U4345 (N_4345,In_3612,In_4471);
nand U4346 (N_4346,In_399,In_2064);
nand U4347 (N_4347,In_2177,In_2691);
nor U4348 (N_4348,In_2705,In_624);
xnor U4349 (N_4349,In_4406,In_1088);
xnor U4350 (N_4350,In_3919,In_2513);
nand U4351 (N_4351,In_853,In_156);
or U4352 (N_4352,In_1141,In_2685);
or U4353 (N_4353,In_4043,In_3766);
xor U4354 (N_4354,In_1578,In_2392);
xnor U4355 (N_4355,In_1217,In_845);
or U4356 (N_4356,In_2654,In_1444);
nor U4357 (N_4357,In_1365,In_3924);
and U4358 (N_4358,In_1307,In_1117);
xnor U4359 (N_4359,In_4704,In_921);
or U4360 (N_4360,In_1358,In_3737);
nand U4361 (N_4361,In_3189,In_380);
and U4362 (N_4362,In_1616,In_1628);
and U4363 (N_4363,In_3932,In_3392);
xnor U4364 (N_4364,In_3351,In_3881);
or U4365 (N_4365,In_2393,In_2507);
xnor U4366 (N_4366,In_1532,In_2498);
xnor U4367 (N_4367,In_4550,In_4190);
or U4368 (N_4368,In_327,In_4687);
nand U4369 (N_4369,In_1005,In_307);
nor U4370 (N_4370,In_1911,In_2713);
nand U4371 (N_4371,In_4165,In_1967);
nand U4372 (N_4372,In_1349,In_4023);
or U4373 (N_4373,In_4731,In_2618);
nor U4374 (N_4374,In_4942,In_3717);
xnor U4375 (N_4375,In_361,In_4667);
xnor U4376 (N_4376,In_3530,In_4360);
xnor U4377 (N_4377,In_3214,In_2492);
or U4378 (N_4378,In_2741,In_530);
xnor U4379 (N_4379,In_2455,In_2679);
and U4380 (N_4380,In_1055,In_4650);
nand U4381 (N_4381,In_568,In_2887);
nor U4382 (N_4382,In_1114,In_3605);
xnor U4383 (N_4383,In_1432,In_3658);
and U4384 (N_4384,In_973,In_3382);
nor U4385 (N_4385,In_182,In_3622);
nand U4386 (N_4386,In_91,In_1836);
and U4387 (N_4387,In_2196,In_1247);
or U4388 (N_4388,In_57,In_2865);
nand U4389 (N_4389,In_1321,In_2709);
nor U4390 (N_4390,In_3519,In_4861);
or U4391 (N_4391,In_3136,In_1584);
and U4392 (N_4392,In_1755,In_3337);
and U4393 (N_4393,In_4887,In_3849);
xor U4394 (N_4394,In_45,In_4234);
xnor U4395 (N_4395,In_183,In_3003);
or U4396 (N_4396,In_35,In_4659);
xor U4397 (N_4397,In_4426,In_3806);
nor U4398 (N_4398,In_1901,In_983);
xor U4399 (N_4399,In_4545,In_59);
nand U4400 (N_4400,In_697,In_1201);
and U4401 (N_4401,In_3047,In_462);
and U4402 (N_4402,In_2870,In_4568);
nand U4403 (N_4403,In_4770,In_4916);
or U4404 (N_4404,In_3264,In_163);
nand U4405 (N_4405,In_4746,In_3271);
xor U4406 (N_4406,In_157,In_4191);
and U4407 (N_4407,In_274,In_3489);
xnor U4408 (N_4408,In_871,In_4913);
nand U4409 (N_4409,In_4911,In_67);
xnor U4410 (N_4410,In_465,In_4715);
and U4411 (N_4411,In_1678,In_1303);
nor U4412 (N_4412,In_3291,In_4814);
and U4413 (N_4413,In_1193,In_2988);
nand U4414 (N_4414,In_585,In_2063);
nor U4415 (N_4415,In_1235,In_2404);
nand U4416 (N_4416,In_2261,In_2227);
nor U4417 (N_4417,In_1905,In_988);
xor U4418 (N_4418,In_33,In_2502);
nand U4419 (N_4419,In_1994,In_1380);
nor U4420 (N_4420,In_3380,In_1959);
or U4421 (N_4421,In_1857,In_2318);
xor U4422 (N_4422,In_1958,In_1518);
xnor U4423 (N_4423,In_100,In_1825);
xor U4424 (N_4424,In_2631,In_4137);
or U4425 (N_4425,In_3197,In_3795);
nand U4426 (N_4426,In_2065,In_2834);
xor U4427 (N_4427,In_964,In_1509);
xnor U4428 (N_4428,In_3576,In_2650);
or U4429 (N_4429,In_837,In_3837);
and U4430 (N_4430,In_4754,In_1447);
or U4431 (N_4431,In_1246,In_3576);
xor U4432 (N_4432,In_4942,In_2006);
xor U4433 (N_4433,In_1079,In_3161);
or U4434 (N_4434,In_3272,In_2671);
and U4435 (N_4435,In_174,In_1320);
and U4436 (N_4436,In_118,In_3913);
or U4437 (N_4437,In_717,In_4878);
nor U4438 (N_4438,In_232,In_2214);
nand U4439 (N_4439,In_1186,In_1375);
nand U4440 (N_4440,In_864,In_4388);
or U4441 (N_4441,In_1356,In_1999);
or U4442 (N_4442,In_579,In_4896);
or U4443 (N_4443,In_2125,In_3703);
nor U4444 (N_4444,In_4799,In_2353);
or U4445 (N_4445,In_2087,In_3495);
xnor U4446 (N_4446,In_4541,In_3948);
or U4447 (N_4447,In_2872,In_314);
xor U4448 (N_4448,In_4845,In_4650);
nand U4449 (N_4449,In_411,In_2057);
and U4450 (N_4450,In_3615,In_4910);
or U4451 (N_4451,In_1027,In_3654);
xor U4452 (N_4452,In_1143,In_166);
nand U4453 (N_4453,In_867,In_1247);
xor U4454 (N_4454,In_155,In_2590);
or U4455 (N_4455,In_2572,In_2529);
nor U4456 (N_4456,In_2194,In_2748);
and U4457 (N_4457,In_2321,In_2204);
and U4458 (N_4458,In_1994,In_3740);
or U4459 (N_4459,In_2884,In_3681);
nor U4460 (N_4460,In_3597,In_1889);
or U4461 (N_4461,In_2940,In_1164);
xor U4462 (N_4462,In_3050,In_129);
xnor U4463 (N_4463,In_1187,In_4782);
nor U4464 (N_4464,In_1014,In_3799);
nand U4465 (N_4465,In_2066,In_4121);
nor U4466 (N_4466,In_4059,In_3141);
or U4467 (N_4467,In_678,In_2892);
xor U4468 (N_4468,In_1787,In_2279);
nor U4469 (N_4469,In_657,In_4927);
nor U4470 (N_4470,In_1500,In_1515);
xor U4471 (N_4471,In_2027,In_3610);
or U4472 (N_4472,In_1977,In_3108);
and U4473 (N_4473,In_3322,In_2062);
or U4474 (N_4474,In_3386,In_4372);
and U4475 (N_4475,In_3142,In_3662);
nand U4476 (N_4476,In_564,In_1292);
or U4477 (N_4477,In_174,In_4176);
nand U4478 (N_4478,In_2600,In_2749);
nand U4479 (N_4479,In_4738,In_818);
nand U4480 (N_4480,In_474,In_4120);
nor U4481 (N_4481,In_2833,In_2068);
and U4482 (N_4482,In_1840,In_439);
xor U4483 (N_4483,In_423,In_330);
xor U4484 (N_4484,In_2586,In_1424);
and U4485 (N_4485,In_12,In_2339);
or U4486 (N_4486,In_2010,In_399);
xnor U4487 (N_4487,In_1697,In_1821);
and U4488 (N_4488,In_1542,In_4905);
nand U4489 (N_4489,In_3936,In_892);
or U4490 (N_4490,In_2285,In_795);
or U4491 (N_4491,In_3705,In_1130);
and U4492 (N_4492,In_2595,In_1928);
nand U4493 (N_4493,In_466,In_4287);
xor U4494 (N_4494,In_4111,In_3323);
xor U4495 (N_4495,In_2740,In_2950);
nor U4496 (N_4496,In_261,In_2891);
xor U4497 (N_4497,In_189,In_4022);
nand U4498 (N_4498,In_914,In_696);
or U4499 (N_4499,In_2116,In_2547);
and U4500 (N_4500,In_3999,In_2488);
nor U4501 (N_4501,In_3476,In_701);
xor U4502 (N_4502,In_4768,In_1169);
and U4503 (N_4503,In_4084,In_2205);
or U4504 (N_4504,In_1842,In_4012);
and U4505 (N_4505,In_1177,In_876);
or U4506 (N_4506,In_589,In_49);
nand U4507 (N_4507,In_2796,In_2265);
nand U4508 (N_4508,In_3614,In_2386);
nand U4509 (N_4509,In_1121,In_4152);
nand U4510 (N_4510,In_469,In_3385);
nand U4511 (N_4511,In_4542,In_3047);
and U4512 (N_4512,In_9,In_2922);
nor U4513 (N_4513,In_1120,In_1710);
and U4514 (N_4514,In_2386,In_3443);
nor U4515 (N_4515,In_3647,In_4209);
xnor U4516 (N_4516,In_3551,In_1613);
nand U4517 (N_4517,In_126,In_2420);
nand U4518 (N_4518,In_827,In_4280);
xor U4519 (N_4519,In_2856,In_3766);
nand U4520 (N_4520,In_2576,In_1984);
or U4521 (N_4521,In_2634,In_2175);
xnor U4522 (N_4522,In_2184,In_461);
nand U4523 (N_4523,In_3555,In_788);
nand U4524 (N_4524,In_3348,In_3961);
xor U4525 (N_4525,In_2648,In_4638);
or U4526 (N_4526,In_3650,In_1000);
xnor U4527 (N_4527,In_4245,In_583);
xor U4528 (N_4528,In_4314,In_1574);
nor U4529 (N_4529,In_2093,In_2931);
or U4530 (N_4530,In_2052,In_804);
nand U4531 (N_4531,In_1972,In_4623);
nand U4532 (N_4532,In_3724,In_1667);
and U4533 (N_4533,In_3942,In_741);
or U4534 (N_4534,In_3157,In_2431);
nand U4535 (N_4535,In_1950,In_2287);
xor U4536 (N_4536,In_4772,In_4072);
nand U4537 (N_4537,In_4198,In_2450);
and U4538 (N_4538,In_1623,In_4220);
xor U4539 (N_4539,In_4225,In_3611);
xor U4540 (N_4540,In_3014,In_4673);
xor U4541 (N_4541,In_4825,In_2396);
nor U4542 (N_4542,In_1986,In_103);
xor U4543 (N_4543,In_4760,In_4336);
nor U4544 (N_4544,In_248,In_4141);
nand U4545 (N_4545,In_3655,In_1038);
xor U4546 (N_4546,In_1446,In_575);
nor U4547 (N_4547,In_3315,In_607);
or U4548 (N_4548,In_1402,In_4557);
nor U4549 (N_4549,In_2126,In_3313);
nand U4550 (N_4550,In_648,In_4148);
and U4551 (N_4551,In_2498,In_3581);
nand U4552 (N_4552,In_3927,In_3541);
xnor U4553 (N_4553,In_2951,In_1378);
xnor U4554 (N_4554,In_4817,In_238);
and U4555 (N_4555,In_4626,In_2225);
nor U4556 (N_4556,In_1150,In_4103);
and U4557 (N_4557,In_1401,In_4936);
and U4558 (N_4558,In_4744,In_1206);
or U4559 (N_4559,In_2137,In_4543);
and U4560 (N_4560,In_2855,In_4624);
nand U4561 (N_4561,In_2112,In_949);
and U4562 (N_4562,In_2706,In_1175);
xor U4563 (N_4563,In_574,In_1975);
or U4564 (N_4564,In_3532,In_148);
nand U4565 (N_4565,In_4330,In_4261);
xor U4566 (N_4566,In_977,In_4789);
xnor U4567 (N_4567,In_4330,In_853);
nor U4568 (N_4568,In_1108,In_4826);
nor U4569 (N_4569,In_4047,In_3690);
xor U4570 (N_4570,In_1539,In_2719);
or U4571 (N_4571,In_2752,In_2263);
xor U4572 (N_4572,In_2858,In_614);
nand U4573 (N_4573,In_3460,In_3148);
nor U4574 (N_4574,In_3144,In_4008);
nand U4575 (N_4575,In_4661,In_4823);
xnor U4576 (N_4576,In_608,In_1835);
and U4577 (N_4577,In_3428,In_3239);
xnor U4578 (N_4578,In_2221,In_3703);
nor U4579 (N_4579,In_638,In_4236);
or U4580 (N_4580,In_644,In_4450);
xnor U4581 (N_4581,In_2185,In_2961);
and U4582 (N_4582,In_3760,In_3203);
xor U4583 (N_4583,In_4086,In_474);
and U4584 (N_4584,In_342,In_3608);
or U4585 (N_4585,In_3021,In_545);
nand U4586 (N_4586,In_144,In_1692);
nand U4587 (N_4587,In_147,In_4886);
or U4588 (N_4588,In_3010,In_2324);
nor U4589 (N_4589,In_1224,In_4189);
or U4590 (N_4590,In_1406,In_976);
xnor U4591 (N_4591,In_3979,In_2283);
or U4592 (N_4592,In_3043,In_2266);
and U4593 (N_4593,In_3032,In_4618);
and U4594 (N_4594,In_1624,In_3753);
and U4595 (N_4595,In_645,In_4226);
nand U4596 (N_4596,In_1455,In_2209);
or U4597 (N_4597,In_381,In_4465);
nand U4598 (N_4598,In_482,In_342);
nor U4599 (N_4599,In_2794,In_228);
xnor U4600 (N_4600,In_4065,In_1044);
xor U4601 (N_4601,In_4724,In_3105);
xor U4602 (N_4602,In_2198,In_2067);
or U4603 (N_4603,In_1203,In_42);
nand U4604 (N_4604,In_2049,In_1766);
nor U4605 (N_4605,In_1062,In_4993);
nor U4606 (N_4606,In_3217,In_1315);
or U4607 (N_4607,In_221,In_2689);
nand U4608 (N_4608,In_2323,In_2398);
xor U4609 (N_4609,In_599,In_1392);
or U4610 (N_4610,In_2684,In_818);
xnor U4611 (N_4611,In_4140,In_3033);
nand U4612 (N_4612,In_1431,In_3530);
or U4613 (N_4613,In_2590,In_827);
and U4614 (N_4614,In_3971,In_1872);
nor U4615 (N_4615,In_977,In_846);
nand U4616 (N_4616,In_2748,In_1759);
nand U4617 (N_4617,In_2259,In_188);
or U4618 (N_4618,In_3590,In_2975);
nor U4619 (N_4619,In_1768,In_1349);
nand U4620 (N_4620,In_4660,In_943);
or U4621 (N_4621,In_1248,In_1346);
nor U4622 (N_4622,In_503,In_3495);
or U4623 (N_4623,In_2223,In_2920);
nand U4624 (N_4624,In_4977,In_4974);
and U4625 (N_4625,In_4033,In_2354);
and U4626 (N_4626,In_1404,In_1401);
nand U4627 (N_4627,In_3386,In_2923);
or U4628 (N_4628,In_1568,In_3037);
and U4629 (N_4629,In_4625,In_2950);
or U4630 (N_4630,In_1841,In_694);
xnor U4631 (N_4631,In_3061,In_492);
nor U4632 (N_4632,In_3618,In_399);
xnor U4633 (N_4633,In_3630,In_1269);
nor U4634 (N_4634,In_937,In_303);
xor U4635 (N_4635,In_2998,In_3180);
and U4636 (N_4636,In_99,In_2170);
and U4637 (N_4637,In_1234,In_2306);
and U4638 (N_4638,In_4656,In_2188);
and U4639 (N_4639,In_4317,In_4390);
and U4640 (N_4640,In_4195,In_1964);
or U4641 (N_4641,In_4237,In_4112);
or U4642 (N_4642,In_2533,In_2331);
and U4643 (N_4643,In_1878,In_996);
or U4644 (N_4644,In_2667,In_4965);
and U4645 (N_4645,In_3058,In_993);
or U4646 (N_4646,In_2339,In_4962);
and U4647 (N_4647,In_972,In_4159);
and U4648 (N_4648,In_1409,In_3422);
or U4649 (N_4649,In_3743,In_3194);
and U4650 (N_4650,In_4379,In_4142);
xnor U4651 (N_4651,In_506,In_2547);
nand U4652 (N_4652,In_3644,In_2989);
xor U4653 (N_4653,In_1075,In_4238);
xnor U4654 (N_4654,In_1658,In_1007);
nand U4655 (N_4655,In_4600,In_2454);
nand U4656 (N_4656,In_3246,In_3714);
and U4657 (N_4657,In_549,In_32);
and U4658 (N_4658,In_4377,In_213);
xor U4659 (N_4659,In_1380,In_3078);
and U4660 (N_4660,In_3292,In_1279);
nand U4661 (N_4661,In_99,In_4680);
or U4662 (N_4662,In_824,In_2960);
nor U4663 (N_4663,In_2260,In_1298);
xor U4664 (N_4664,In_2957,In_3948);
nand U4665 (N_4665,In_1785,In_2367);
nand U4666 (N_4666,In_4155,In_685);
and U4667 (N_4667,In_1493,In_2118);
and U4668 (N_4668,In_3968,In_4255);
nor U4669 (N_4669,In_4510,In_4448);
or U4670 (N_4670,In_2337,In_1777);
xor U4671 (N_4671,In_1746,In_3800);
or U4672 (N_4672,In_969,In_1499);
nor U4673 (N_4673,In_2251,In_186);
xor U4674 (N_4674,In_1414,In_306);
and U4675 (N_4675,In_4209,In_991);
and U4676 (N_4676,In_179,In_730);
or U4677 (N_4677,In_4633,In_2349);
nor U4678 (N_4678,In_1376,In_932);
nor U4679 (N_4679,In_2029,In_2733);
nand U4680 (N_4680,In_2096,In_1942);
nor U4681 (N_4681,In_420,In_377);
nand U4682 (N_4682,In_1091,In_450);
nor U4683 (N_4683,In_2464,In_1593);
nand U4684 (N_4684,In_1009,In_2975);
nor U4685 (N_4685,In_742,In_226);
xor U4686 (N_4686,In_1467,In_1767);
or U4687 (N_4687,In_630,In_3280);
or U4688 (N_4688,In_4741,In_1281);
xnor U4689 (N_4689,In_1010,In_397);
or U4690 (N_4690,In_4193,In_492);
and U4691 (N_4691,In_3224,In_4638);
or U4692 (N_4692,In_3499,In_1911);
nand U4693 (N_4693,In_2405,In_1060);
nor U4694 (N_4694,In_4589,In_622);
nand U4695 (N_4695,In_128,In_4231);
and U4696 (N_4696,In_4776,In_3465);
nand U4697 (N_4697,In_1525,In_1515);
and U4698 (N_4698,In_1097,In_1956);
or U4699 (N_4699,In_3152,In_223);
nand U4700 (N_4700,In_4996,In_4979);
nand U4701 (N_4701,In_4122,In_3134);
or U4702 (N_4702,In_4489,In_1584);
and U4703 (N_4703,In_4667,In_4391);
xor U4704 (N_4704,In_3001,In_3039);
and U4705 (N_4705,In_1786,In_3470);
or U4706 (N_4706,In_3907,In_4907);
xor U4707 (N_4707,In_4131,In_461);
nor U4708 (N_4708,In_1729,In_1498);
nor U4709 (N_4709,In_1971,In_4497);
xor U4710 (N_4710,In_1552,In_3207);
or U4711 (N_4711,In_1157,In_935);
xor U4712 (N_4712,In_2348,In_1987);
or U4713 (N_4713,In_831,In_4054);
and U4714 (N_4714,In_2833,In_1016);
and U4715 (N_4715,In_4391,In_3584);
or U4716 (N_4716,In_4326,In_95);
xor U4717 (N_4717,In_904,In_1325);
or U4718 (N_4718,In_1859,In_4091);
or U4719 (N_4719,In_3990,In_2832);
or U4720 (N_4720,In_132,In_4293);
xnor U4721 (N_4721,In_863,In_2330);
nor U4722 (N_4722,In_1943,In_4303);
or U4723 (N_4723,In_3398,In_4715);
and U4724 (N_4724,In_624,In_3526);
nand U4725 (N_4725,In_291,In_4276);
nand U4726 (N_4726,In_2615,In_4978);
and U4727 (N_4727,In_3747,In_1438);
and U4728 (N_4728,In_4689,In_2106);
xor U4729 (N_4729,In_742,In_4987);
nor U4730 (N_4730,In_597,In_4815);
and U4731 (N_4731,In_4973,In_2505);
or U4732 (N_4732,In_1263,In_3876);
xor U4733 (N_4733,In_526,In_287);
nand U4734 (N_4734,In_1589,In_4248);
nand U4735 (N_4735,In_1863,In_854);
nor U4736 (N_4736,In_176,In_4559);
nor U4737 (N_4737,In_4096,In_3034);
and U4738 (N_4738,In_2775,In_2055);
and U4739 (N_4739,In_4803,In_4898);
xor U4740 (N_4740,In_992,In_696);
or U4741 (N_4741,In_2277,In_2411);
and U4742 (N_4742,In_3238,In_3824);
xnor U4743 (N_4743,In_2231,In_248);
xnor U4744 (N_4744,In_4624,In_2461);
and U4745 (N_4745,In_2965,In_1727);
or U4746 (N_4746,In_3219,In_2635);
xnor U4747 (N_4747,In_126,In_2445);
nor U4748 (N_4748,In_518,In_1452);
or U4749 (N_4749,In_3199,In_1698);
nor U4750 (N_4750,In_1826,In_1656);
nor U4751 (N_4751,In_4883,In_2237);
xnor U4752 (N_4752,In_208,In_3081);
xnor U4753 (N_4753,In_2919,In_4622);
and U4754 (N_4754,In_856,In_3331);
and U4755 (N_4755,In_407,In_1377);
xor U4756 (N_4756,In_4686,In_1562);
xnor U4757 (N_4757,In_778,In_4962);
or U4758 (N_4758,In_4567,In_292);
xnor U4759 (N_4759,In_1133,In_1879);
or U4760 (N_4760,In_1637,In_1638);
nor U4761 (N_4761,In_4141,In_698);
or U4762 (N_4762,In_2543,In_549);
nor U4763 (N_4763,In_3956,In_952);
and U4764 (N_4764,In_862,In_3528);
and U4765 (N_4765,In_4001,In_4908);
or U4766 (N_4766,In_1921,In_2957);
nor U4767 (N_4767,In_2015,In_36);
and U4768 (N_4768,In_3903,In_663);
xor U4769 (N_4769,In_2587,In_4821);
nand U4770 (N_4770,In_1992,In_4304);
and U4771 (N_4771,In_1879,In_4605);
or U4772 (N_4772,In_692,In_1805);
or U4773 (N_4773,In_4072,In_2881);
and U4774 (N_4774,In_2693,In_767);
and U4775 (N_4775,In_149,In_357);
or U4776 (N_4776,In_1546,In_2733);
xor U4777 (N_4777,In_1585,In_2276);
or U4778 (N_4778,In_1875,In_3531);
nand U4779 (N_4779,In_1359,In_3255);
xnor U4780 (N_4780,In_4965,In_4851);
nand U4781 (N_4781,In_4632,In_3314);
nor U4782 (N_4782,In_4725,In_2134);
nor U4783 (N_4783,In_1368,In_2042);
nor U4784 (N_4784,In_3058,In_1569);
nor U4785 (N_4785,In_2890,In_4519);
nand U4786 (N_4786,In_3315,In_1784);
nand U4787 (N_4787,In_1593,In_4507);
nor U4788 (N_4788,In_2655,In_436);
or U4789 (N_4789,In_1360,In_788);
and U4790 (N_4790,In_4449,In_1863);
xnor U4791 (N_4791,In_4425,In_2761);
or U4792 (N_4792,In_2983,In_4764);
nor U4793 (N_4793,In_1034,In_2973);
xnor U4794 (N_4794,In_1849,In_4294);
and U4795 (N_4795,In_1634,In_1675);
or U4796 (N_4796,In_122,In_1875);
nor U4797 (N_4797,In_949,In_1493);
xnor U4798 (N_4798,In_3858,In_1094);
nor U4799 (N_4799,In_3664,In_3302);
and U4800 (N_4800,In_831,In_2227);
or U4801 (N_4801,In_2216,In_4355);
xnor U4802 (N_4802,In_3148,In_1575);
or U4803 (N_4803,In_4886,In_3699);
nor U4804 (N_4804,In_3260,In_1058);
or U4805 (N_4805,In_4795,In_4304);
or U4806 (N_4806,In_4897,In_2315);
and U4807 (N_4807,In_3936,In_588);
nor U4808 (N_4808,In_3935,In_2644);
xnor U4809 (N_4809,In_4829,In_3287);
xor U4810 (N_4810,In_1990,In_521);
and U4811 (N_4811,In_2559,In_4043);
xnor U4812 (N_4812,In_3018,In_2996);
or U4813 (N_4813,In_3463,In_2727);
xor U4814 (N_4814,In_3315,In_3346);
nand U4815 (N_4815,In_2100,In_611);
nor U4816 (N_4816,In_1572,In_2864);
and U4817 (N_4817,In_550,In_2583);
nor U4818 (N_4818,In_2903,In_2095);
nand U4819 (N_4819,In_336,In_2088);
nor U4820 (N_4820,In_1264,In_4310);
nand U4821 (N_4821,In_3505,In_4209);
nand U4822 (N_4822,In_1579,In_4713);
xnor U4823 (N_4823,In_2599,In_3149);
and U4824 (N_4824,In_205,In_2874);
nand U4825 (N_4825,In_2375,In_741);
and U4826 (N_4826,In_3004,In_2657);
or U4827 (N_4827,In_1124,In_1276);
nand U4828 (N_4828,In_3896,In_4563);
xnor U4829 (N_4829,In_3382,In_3696);
xnor U4830 (N_4830,In_3549,In_1351);
xnor U4831 (N_4831,In_2060,In_170);
xor U4832 (N_4832,In_2719,In_3593);
and U4833 (N_4833,In_3180,In_1526);
xor U4834 (N_4834,In_3341,In_1509);
nor U4835 (N_4835,In_3789,In_1548);
nor U4836 (N_4836,In_1095,In_4117);
or U4837 (N_4837,In_2753,In_4556);
or U4838 (N_4838,In_4017,In_3197);
xor U4839 (N_4839,In_1369,In_2491);
nor U4840 (N_4840,In_476,In_4006);
xor U4841 (N_4841,In_2490,In_2588);
or U4842 (N_4842,In_4184,In_2871);
and U4843 (N_4843,In_1572,In_4568);
nand U4844 (N_4844,In_4311,In_4012);
and U4845 (N_4845,In_3609,In_1755);
xnor U4846 (N_4846,In_4258,In_3852);
or U4847 (N_4847,In_2973,In_1118);
xnor U4848 (N_4848,In_177,In_4809);
xnor U4849 (N_4849,In_356,In_2765);
nor U4850 (N_4850,In_3489,In_388);
nand U4851 (N_4851,In_3197,In_3784);
nor U4852 (N_4852,In_1982,In_2450);
nor U4853 (N_4853,In_2647,In_3371);
and U4854 (N_4854,In_3321,In_4289);
and U4855 (N_4855,In_2705,In_181);
nor U4856 (N_4856,In_811,In_4516);
and U4857 (N_4857,In_4515,In_374);
nor U4858 (N_4858,In_1816,In_490);
or U4859 (N_4859,In_1831,In_323);
and U4860 (N_4860,In_4880,In_39);
and U4861 (N_4861,In_4323,In_3913);
xor U4862 (N_4862,In_3425,In_397);
xnor U4863 (N_4863,In_529,In_741);
nand U4864 (N_4864,In_261,In_1712);
nand U4865 (N_4865,In_518,In_291);
nor U4866 (N_4866,In_4190,In_3197);
or U4867 (N_4867,In_4312,In_486);
xnor U4868 (N_4868,In_3362,In_898);
nand U4869 (N_4869,In_2626,In_29);
or U4870 (N_4870,In_988,In_4930);
xnor U4871 (N_4871,In_813,In_4587);
and U4872 (N_4872,In_759,In_4304);
nand U4873 (N_4873,In_4343,In_2467);
nand U4874 (N_4874,In_4930,In_2413);
and U4875 (N_4875,In_3901,In_1144);
nand U4876 (N_4876,In_42,In_536);
nand U4877 (N_4877,In_173,In_1836);
nand U4878 (N_4878,In_1962,In_1638);
nand U4879 (N_4879,In_1216,In_716);
or U4880 (N_4880,In_4625,In_537);
xor U4881 (N_4881,In_1632,In_2516);
xor U4882 (N_4882,In_1281,In_2927);
xor U4883 (N_4883,In_27,In_1205);
nand U4884 (N_4884,In_4233,In_3762);
and U4885 (N_4885,In_3009,In_2730);
or U4886 (N_4886,In_2899,In_1772);
nor U4887 (N_4887,In_2980,In_4883);
nor U4888 (N_4888,In_2563,In_3710);
and U4889 (N_4889,In_704,In_528);
nand U4890 (N_4890,In_1498,In_4222);
and U4891 (N_4891,In_1319,In_3108);
xor U4892 (N_4892,In_54,In_4635);
or U4893 (N_4893,In_2818,In_84);
nand U4894 (N_4894,In_1274,In_1559);
nand U4895 (N_4895,In_330,In_2854);
or U4896 (N_4896,In_629,In_2088);
or U4897 (N_4897,In_1234,In_1379);
or U4898 (N_4898,In_4175,In_2720);
and U4899 (N_4899,In_3188,In_1397);
or U4900 (N_4900,In_4144,In_4799);
nand U4901 (N_4901,In_1031,In_3362);
nor U4902 (N_4902,In_3097,In_3575);
and U4903 (N_4903,In_3545,In_814);
or U4904 (N_4904,In_2455,In_4029);
nor U4905 (N_4905,In_2060,In_1507);
and U4906 (N_4906,In_832,In_1855);
or U4907 (N_4907,In_2535,In_3201);
xor U4908 (N_4908,In_939,In_1338);
and U4909 (N_4909,In_4075,In_2529);
nor U4910 (N_4910,In_715,In_3450);
nor U4911 (N_4911,In_4479,In_2967);
xor U4912 (N_4912,In_4344,In_2898);
and U4913 (N_4913,In_4218,In_3879);
xor U4914 (N_4914,In_3153,In_3591);
xor U4915 (N_4915,In_2051,In_2967);
and U4916 (N_4916,In_1462,In_1648);
and U4917 (N_4917,In_109,In_2481);
nor U4918 (N_4918,In_4174,In_3694);
and U4919 (N_4919,In_4793,In_3687);
and U4920 (N_4920,In_922,In_3433);
nor U4921 (N_4921,In_2982,In_1170);
or U4922 (N_4922,In_1517,In_2775);
nor U4923 (N_4923,In_1394,In_1253);
nand U4924 (N_4924,In_2457,In_1156);
nor U4925 (N_4925,In_3074,In_168);
nor U4926 (N_4926,In_691,In_4980);
and U4927 (N_4927,In_3819,In_2819);
xnor U4928 (N_4928,In_2780,In_4202);
nor U4929 (N_4929,In_946,In_4790);
and U4930 (N_4930,In_3929,In_599);
xor U4931 (N_4931,In_3611,In_3514);
and U4932 (N_4932,In_3778,In_2568);
nor U4933 (N_4933,In_3257,In_3362);
or U4934 (N_4934,In_694,In_2825);
and U4935 (N_4935,In_4844,In_2199);
nor U4936 (N_4936,In_923,In_3647);
or U4937 (N_4937,In_4648,In_2404);
and U4938 (N_4938,In_2475,In_3659);
nor U4939 (N_4939,In_4794,In_3045);
and U4940 (N_4940,In_4425,In_4514);
and U4941 (N_4941,In_3178,In_2466);
nor U4942 (N_4942,In_4954,In_3283);
nand U4943 (N_4943,In_1126,In_2985);
nor U4944 (N_4944,In_4714,In_1336);
and U4945 (N_4945,In_1848,In_2563);
xor U4946 (N_4946,In_4365,In_4554);
xnor U4947 (N_4947,In_1674,In_4569);
xnor U4948 (N_4948,In_2408,In_3805);
xor U4949 (N_4949,In_4073,In_3366);
or U4950 (N_4950,In_1745,In_388);
and U4951 (N_4951,In_2662,In_1113);
nor U4952 (N_4952,In_456,In_2398);
and U4953 (N_4953,In_4557,In_151);
nor U4954 (N_4954,In_2003,In_820);
and U4955 (N_4955,In_1727,In_1698);
xnor U4956 (N_4956,In_2413,In_95);
nand U4957 (N_4957,In_2551,In_851);
or U4958 (N_4958,In_2290,In_4710);
xnor U4959 (N_4959,In_4083,In_2629);
or U4960 (N_4960,In_4410,In_2172);
xnor U4961 (N_4961,In_4708,In_1217);
or U4962 (N_4962,In_469,In_1063);
or U4963 (N_4963,In_4027,In_1140);
and U4964 (N_4964,In_4629,In_4530);
or U4965 (N_4965,In_1664,In_1819);
or U4966 (N_4966,In_4987,In_1706);
nand U4967 (N_4967,In_923,In_1493);
xnor U4968 (N_4968,In_382,In_4197);
or U4969 (N_4969,In_2946,In_3590);
nor U4970 (N_4970,In_1413,In_3767);
and U4971 (N_4971,In_1735,In_3674);
nor U4972 (N_4972,In_332,In_2775);
or U4973 (N_4973,In_3363,In_449);
or U4974 (N_4974,In_1854,In_4109);
and U4975 (N_4975,In_3951,In_1651);
and U4976 (N_4976,In_1559,In_1147);
nor U4977 (N_4977,In_799,In_584);
and U4978 (N_4978,In_3078,In_4578);
and U4979 (N_4979,In_4289,In_4079);
nand U4980 (N_4980,In_1001,In_3549);
xnor U4981 (N_4981,In_3637,In_2491);
nand U4982 (N_4982,In_4524,In_3674);
and U4983 (N_4983,In_3920,In_4925);
nand U4984 (N_4984,In_999,In_1393);
and U4985 (N_4985,In_4451,In_2007);
nor U4986 (N_4986,In_1563,In_1731);
or U4987 (N_4987,In_1546,In_1938);
or U4988 (N_4988,In_4647,In_3267);
nand U4989 (N_4989,In_316,In_3594);
nor U4990 (N_4990,In_3981,In_2101);
or U4991 (N_4991,In_283,In_215);
and U4992 (N_4992,In_4230,In_4196);
and U4993 (N_4993,In_2858,In_1261);
nand U4994 (N_4994,In_607,In_1031);
nand U4995 (N_4995,In_2866,In_3894);
or U4996 (N_4996,In_4024,In_1284);
xor U4997 (N_4997,In_1173,In_656);
xnor U4998 (N_4998,In_1602,In_3413);
nor U4999 (N_4999,In_4890,In_1919);
nor U5000 (N_5000,In_2408,In_352);
and U5001 (N_5001,In_2516,In_2340);
nor U5002 (N_5002,In_2337,In_4500);
nor U5003 (N_5003,In_3310,In_3084);
nor U5004 (N_5004,In_292,In_354);
xnor U5005 (N_5005,In_4726,In_299);
nor U5006 (N_5006,In_2300,In_1158);
nand U5007 (N_5007,In_1028,In_4483);
nor U5008 (N_5008,In_4369,In_3847);
or U5009 (N_5009,In_4260,In_2082);
nand U5010 (N_5010,In_2787,In_56);
nand U5011 (N_5011,In_3352,In_2660);
nand U5012 (N_5012,In_4410,In_3554);
nor U5013 (N_5013,In_3643,In_1707);
or U5014 (N_5014,In_3387,In_3975);
nor U5015 (N_5015,In_3670,In_2840);
xnor U5016 (N_5016,In_4546,In_3504);
xnor U5017 (N_5017,In_2446,In_4357);
nor U5018 (N_5018,In_3460,In_3203);
or U5019 (N_5019,In_170,In_2921);
nor U5020 (N_5020,In_3610,In_1916);
or U5021 (N_5021,In_3406,In_3789);
nand U5022 (N_5022,In_3645,In_4629);
nor U5023 (N_5023,In_409,In_2348);
or U5024 (N_5024,In_1301,In_4693);
or U5025 (N_5025,In_378,In_2219);
xnor U5026 (N_5026,In_1538,In_4651);
nand U5027 (N_5027,In_4464,In_1992);
or U5028 (N_5028,In_2888,In_3941);
and U5029 (N_5029,In_2795,In_4334);
nor U5030 (N_5030,In_2339,In_4797);
nor U5031 (N_5031,In_4171,In_3278);
and U5032 (N_5032,In_3464,In_4292);
nor U5033 (N_5033,In_2215,In_3076);
xor U5034 (N_5034,In_548,In_1561);
or U5035 (N_5035,In_324,In_2341);
nor U5036 (N_5036,In_2207,In_4344);
or U5037 (N_5037,In_4663,In_4044);
nor U5038 (N_5038,In_2932,In_2285);
xnor U5039 (N_5039,In_2567,In_2439);
or U5040 (N_5040,In_950,In_429);
nand U5041 (N_5041,In_4977,In_1903);
and U5042 (N_5042,In_2883,In_864);
xor U5043 (N_5043,In_4836,In_4109);
and U5044 (N_5044,In_84,In_2641);
and U5045 (N_5045,In_4166,In_3221);
or U5046 (N_5046,In_2417,In_945);
and U5047 (N_5047,In_1432,In_3945);
and U5048 (N_5048,In_2758,In_129);
nor U5049 (N_5049,In_567,In_1346);
or U5050 (N_5050,In_2894,In_555);
and U5051 (N_5051,In_2158,In_3040);
or U5052 (N_5052,In_1727,In_4814);
or U5053 (N_5053,In_361,In_2515);
nand U5054 (N_5054,In_1585,In_183);
xor U5055 (N_5055,In_1987,In_4425);
and U5056 (N_5056,In_1777,In_1655);
nand U5057 (N_5057,In_212,In_1577);
xor U5058 (N_5058,In_3594,In_817);
nor U5059 (N_5059,In_4090,In_399);
xnor U5060 (N_5060,In_1739,In_1461);
nand U5061 (N_5061,In_576,In_397);
or U5062 (N_5062,In_4059,In_2832);
nor U5063 (N_5063,In_1181,In_1122);
and U5064 (N_5064,In_3260,In_4455);
or U5065 (N_5065,In_2899,In_2253);
nand U5066 (N_5066,In_3022,In_2108);
xor U5067 (N_5067,In_4603,In_1837);
xor U5068 (N_5068,In_2994,In_4832);
nor U5069 (N_5069,In_2671,In_2779);
and U5070 (N_5070,In_2556,In_2585);
xnor U5071 (N_5071,In_47,In_1857);
nor U5072 (N_5072,In_2788,In_4368);
nor U5073 (N_5073,In_70,In_4970);
nor U5074 (N_5074,In_4506,In_4037);
and U5075 (N_5075,In_2088,In_4310);
nor U5076 (N_5076,In_216,In_4735);
and U5077 (N_5077,In_1558,In_4675);
nor U5078 (N_5078,In_2575,In_2237);
or U5079 (N_5079,In_221,In_3215);
and U5080 (N_5080,In_1737,In_3391);
and U5081 (N_5081,In_95,In_4928);
nor U5082 (N_5082,In_460,In_1677);
or U5083 (N_5083,In_1805,In_4399);
xor U5084 (N_5084,In_1830,In_352);
nor U5085 (N_5085,In_1845,In_4338);
xnor U5086 (N_5086,In_3754,In_289);
and U5087 (N_5087,In_1965,In_4998);
nand U5088 (N_5088,In_3604,In_1483);
or U5089 (N_5089,In_918,In_743);
xnor U5090 (N_5090,In_4064,In_2807);
and U5091 (N_5091,In_4179,In_3480);
nand U5092 (N_5092,In_4220,In_1086);
nor U5093 (N_5093,In_1996,In_1238);
or U5094 (N_5094,In_1402,In_3628);
and U5095 (N_5095,In_2753,In_4037);
or U5096 (N_5096,In_4170,In_449);
nand U5097 (N_5097,In_2912,In_673);
or U5098 (N_5098,In_2946,In_3422);
nand U5099 (N_5099,In_1925,In_4908);
nand U5100 (N_5100,In_4900,In_1058);
nor U5101 (N_5101,In_3885,In_3499);
or U5102 (N_5102,In_1567,In_2012);
xnor U5103 (N_5103,In_335,In_3295);
nand U5104 (N_5104,In_3735,In_4758);
xnor U5105 (N_5105,In_4826,In_754);
xnor U5106 (N_5106,In_939,In_1400);
or U5107 (N_5107,In_434,In_3263);
or U5108 (N_5108,In_474,In_1897);
xor U5109 (N_5109,In_4896,In_4920);
or U5110 (N_5110,In_2518,In_2090);
and U5111 (N_5111,In_1280,In_1476);
nor U5112 (N_5112,In_3953,In_1045);
xnor U5113 (N_5113,In_3304,In_3242);
xnor U5114 (N_5114,In_597,In_1040);
xor U5115 (N_5115,In_509,In_1921);
or U5116 (N_5116,In_2107,In_4362);
nand U5117 (N_5117,In_4964,In_655);
nand U5118 (N_5118,In_3461,In_1863);
nor U5119 (N_5119,In_4062,In_165);
and U5120 (N_5120,In_2127,In_2624);
or U5121 (N_5121,In_2090,In_158);
nand U5122 (N_5122,In_2141,In_3549);
nor U5123 (N_5123,In_3270,In_2339);
or U5124 (N_5124,In_322,In_3365);
nor U5125 (N_5125,In_4325,In_3211);
xnor U5126 (N_5126,In_3269,In_3801);
and U5127 (N_5127,In_2694,In_549);
nand U5128 (N_5128,In_3774,In_4654);
and U5129 (N_5129,In_3201,In_4705);
xor U5130 (N_5130,In_591,In_4516);
xnor U5131 (N_5131,In_595,In_3781);
nor U5132 (N_5132,In_2342,In_532);
nor U5133 (N_5133,In_1118,In_2460);
xor U5134 (N_5134,In_3184,In_14);
xor U5135 (N_5135,In_2971,In_2001);
nor U5136 (N_5136,In_894,In_1970);
and U5137 (N_5137,In_2142,In_1973);
or U5138 (N_5138,In_4859,In_195);
nand U5139 (N_5139,In_2035,In_2203);
xor U5140 (N_5140,In_3508,In_1457);
or U5141 (N_5141,In_2803,In_3921);
or U5142 (N_5142,In_4785,In_403);
and U5143 (N_5143,In_3219,In_3886);
nand U5144 (N_5144,In_632,In_2623);
xor U5145 (N_5145,In_4101,In_2684);
nor U5146 (N_5146,In_1271,In_4602);
nor U5147 (N_5147,In_2495,In_3660);
nand U5148 (N_5148,In_1193,In_4952);
xnor U5149 (N_5149,In_2628,In_280);
or U5150 (N_5150,In_2366,In_1770);
or U5151 (N_5151,In_2981,In_698);
or U5152 (N_5152,In_3981,In_4714);
xor U5153 (N_5153,In_3623,In_3415);
xnor U5154 (N_5154,In_1180,In_3380);
or U5155 (N_5155,In_1992,In_1210);
nor U5156 (N_5156,In_2235,In_33);
or U5157 (N_5157,In_3577,In_3766);
nor U5158 (N_5158,In_3959,In_1822);
or U5159 (N_5159,In_2082,In_1915);
nor U5160 (N_5160,In_3108,In_4547);
nor U5161 (N_5161,In_1509,In_4470);
or U5162 (N_5162,In_4986,In_3949);
xor U5163 (N_5163,In_1663,In_3391);
or U5164 (N_5164,In_1242,In_3057);
nand U5165 (N_5165,In_1834,In_3266);
nand U5166 (N_5166,In_3250,In_4295);
xor U5167 (N_5167,In_1091,In_2402);
nor U5168 (N_5168,In_3607,In_3086);
nor U5169 (N_5169,In_3129,In_2964);
and U5170 (N_5170,In_2418,In_3349);
and U5171 (N_5171,In_4903,In_2234);
nand U5172 (N_5172,In_3107,In_2603);
xnor U5173 (N_5173,In_4159,In_3884);
xor U5174 (N_5174,In_4335,In_3369);
nand U5175 (N_5175,In_3309,In_2522);
xor U5176 (N_5176,In_4562,In_1915);
and U5177 (N_5177,In_4684,In_540);
or U5178 (N_5178,In_602,In_1231);
xnor U5179 (N_5179,In_4379,In_4040);
nand U5180 (N_5180,In_989,In_4099);
nor U5181 (N_5181,In_3839,In_2340);
and U5182 (N_5182,In_830,In_3917);
and U5183 (N_5183,In_4509,In_4403);
nand U5184 (N_5184,In_3538,In_2507);
xor U5185 (N_5185,In_1751,In_1342);
xor U5186 (N_5186,In_3271,In_1752);
and U5187 (N_5187,In_4748,In_980);
nor U5188 (N_5188,In_771,In_363);
and U5189 (N_5189,In_90,In_1280);
nor U5190 (N_5190,In_2459,In_1520);
nor U5191 (N_5191,In_158,In_2387);
nor U5192 (N_5192,In_4172,In_1946);
and U5193 (N_5193,In_1191,In_3233);
xnor U5194 (N_5194,In_1700,In_2523);
nor U5195 (N_5195,In_973,In_1782);
nor U5196 (N_5196,In_2401,In_4733);
nor U5197 (N_5197,In_3480,In_2261);
or U5198 (N_5198,In_49,In_1290);
xor U5199 (N_5199,In_4386,In_2617);
nand U5200 (N_5200,In_4277,In_131);
nor U5201 (N_5201,In_3598,In_4898);
nand U5202 (N_5202,In_1280,In_4548);
xnor U5203 (N_5203,In_369,In_3911);
nand U5204 (N_5204,In_4943,In_4191);
nor U5205 (N_5205,In_4282,In_708);
nor U5206 (N_5206,In_967,In_3812);
and U5207 (N_5207,In_1029,In_883);
nand U5208 (N_5208,In_27,In_4510);
nor U5209 (N_5209,In_3751,In_2385);
xor U5210 (N_5210,In_2935,In_1621);
or U5211 (N_5211,In_4590,In_486);
nor U5212 (N_5212,In_2454,In_1126);
or U5213 (N_5213,In_2085,In_3493);
xnor U5214 (N_5214,In_3385,In_1314);
nor U5215 (N_5215,In_3965,In_698);
or U5216 (N_5216,In_1236,In_3707);
nor U5217 (N_5217,In_2246,In_4527);
or U5218 (N_5218,In_1579,In_4651);
xnor U5219 (N_5219,In_1703,In_1536);
or U5220 (N_5220,In_4647,In_2034);
nand U5221 (N_5221,In_3316,In_4982);
nor U5222 (N_5222,In_4440,In_196);
or U5223 (N_5223,In_93,In_1443);
or U5224 (N_5224,In_2501,In_2267);
nand U5225 (N_5225,In_2108,In_2732);
nand U5226 (N_5226,In_3606,In_3454);
or U5227 (N_5227,In_2680,In_2835);
or U5228 (N_5228,In_3033,In_713);
and U5229 (N_5229,In_2732,In_4851);
or U5230 (N_5230,In_2244,In_2622);
nor U5231 (N_5231,In_504,In_3343);
xnor U5232 (N_5232,In_1755,In_4375);
and U5233 (N_5233,In_4703,In_4981);
nand U5234 (N_5234,In_2747,In_4518);
or U5235 (N_5235,In_2747,In_3152);
or U5236 (N_5236,In_4213,In_1452);
nor U5237 (N_5237,In_1175,In_4092);
nor U5238 (N_5238,In_3192,In_233);
nand U5239 (N_5239,In_552,In_1006);
and U5240 (N_5240,In_1147,In_4541);
and U5241 (N_5241,In_1662,In_3628);
nand U5242 (N_5242,In_2776,In_2023);
xnor U5243 (N_5243,In_615,In_2867);
and U5244 (N_5244,In_3134,In_1140);
nand U5245 (N_5245,In_3784,In_4864);
xor U5246 (N_5246,In_3916,In_2620);
nor U5247 (N_5247,In_3337,In_2308);
nand U5248 (N_5248,In_836,In_139);
nand U5249 (N_5249,In_4554,In_792);
nor U5250 (N_5250,In_3891,In_4029);
xnor U5251 (N_5251,In_4111,In_1043);
nor U5252 (N_5252,In_4992,In_3215);
nor U5253 (N_5253,In_224,In_871);
nor U5254 (N_5254,In_1905,In_1614);
nand U5255 (N_5255,In_539,In_70);
nor U5256 (N_5256,In_3288,In_2476);
nand U5257 (N_5257,In_1769,In_4094);
nand U5258 (N_5258,In_3079,In_2582);
and U5259 (N_5259,In_3343,In_4028);
and U5260 (N_5260,In_4801,In_2347);
nor U5261 (N_5261,In_895,In_2852);
nand U5262 (N_5262,In_3061,In_893);
and U5263 (N_5263,In_758,In_3561);
nand U5264 (N_5264,In_3597,In_172);
or U5265 (N_5265,In_1279,In_4661);
and U5266 (N_5266,In_2653,In_1233);
nand U5267 (N_5267,In_1255,In_1607);
nor U5268 (N_5268,In_1146,In_672);
nor U5269 (N_5269,In_4694,In_219);
nor U5270 (N_5270,In_2888,In_4537);
nor U5271 (N_5271,In_3187,In_1249);
or U5272 (N_5272,In_2307,In_3928);
nand U5273 (N_5273,In_4052,In_4671);
nand U5274 (N_5274,In_4605,In_3629);
and U5275 (N_5275,In_4374,In_1484);
nor U5276 (N_5276,In_1765,In_4945);
or U5277 (N_5277,In_3873,In_1573);
nand U5278 (N_5278,In_2121,In_3481);
nand U5279 (N_5279,In_3657,In_2642);
and U5280 (N_5280,In_2208,In_1471);
or U5281 (N_5281,In_488,In_177);
xnor U5282 (N_5282,In_4442,In_1061);
xnor U5283 (N_5283,In_2609,In_0);
nor U5284 (N_5284,In_2170,In_697);
nor U5285 (N_5285,In_970,In_2901);
nor U5286 (N_5286,In_1078,In_1645);
and U5287 (N_5287,In_3250,In_2421);
xor U5288 (N_5288,In_1670,In_4851);
xor U5289 (N_5289,In_312,In_2820);
or U5290 (N_5290,In_390,In_4647);
or U5291 (N_5291,In_4221,In_2146);
xor U5292 (N_5292,In_3044,In_1700);
and U5293 (N_5293,In_992,In_622);
or U5294 (N_5294,In_547,In_912);
or U5295 (N_5295,In_2152,In_2714);
xor U5296 (N_5296,In_1394,In_4704);
and U5297 (N_5297,In_2452,In_1762);
and U5298 (N_5298,In_2391,In_986);
xnor U5299 (N_5299,In_3553,In_2669);
and U5300 (N_5300,In_1320,In_749);
or U5301 (N_5301,In_4887,In_1050);
xor U5302 (N_5302,In_3794,In_3851);
and U5303 (N_5303,In_4366,In_4079);
or U5304 (N_5304,In_2130,In_3187);
nor U5305 (N_5305,In_1922,In_3123);
or U5306 (N_5306,In_4900,In_2351);
xnor U5307 (N_5307,In_199,In_4863);
xnor U5308 (N_5308,In_207,In_2729);
and U5309 (N_5309,In_4050,In_264);
xor U5310 (N_5310,In_722,In_523);
or U5311 (N_5311,In_1301,In_2526);
or U5312 (N_5312,In_1995,In_3982);
xnor U5313 (N_5313,In_4324,In_809);
nor U5314 (N_5314,In_1427,In_2275);
xnor U5315 (N_5315,In_1718,In_2932);
xor U5316 (N_5316,In_4305,In_2354);
or U5317 (N_5317,In_1317,In_1536);
nor U5318 (N_5318,In_2622,In_2508);
nand U5319 (N_5319,In_739,In_2510);
xnor U5320 (N_5320,In_1741,In_1030);
nand U5321 (N_5321,In_908,In_2413);
or U5322 (N_5322,In_3299,In_2153);
or U5323 (N_5323,In_452,In_2434);
and U5324 (N_5324,In_4844,In_3615);
xor U5325 (N_5325,In_2751,In_4933);
nand U5326 (N_5326,In_4601,In_4247);
and U5327 (N_5327,In_2666,In_3761);
nand U5328 (N_5328,In_178,In_3533);
nor U5329 (N_5329,In_2936,In_2831);
nor U5330 (N_5330,In_104,In_1325);
or U5331 (N_5331,In_3085,In_1188);
nand U5332 (N_5332,In_647,In_4785);
nand U5333 (N_5333,In_4602,In_3024);
xor U5334 (N_5334,In_3516,In_3391);
xor U5335 (N_5335,In_3619,In_3129);
nand U5336 (N_5336,In_1315,In_1286);
xor U5337 (N_5337,In_960,In_2442);
nor U5338 (N_5338,In_1248,In_1545);
or U5339 (N_5339,In_856,In_1729);
nand U5340 (N_5340,In_1342,In_854);
xor U5341 (N_5341,In_2455,In_3585);
nor U5342 (N_5342,In_3510,In_3972);
and U5343 (N_5343,In_2035,In_998);
xor U5344 (N_5344,In_1563,In_50);
and U5345 (N_5345,In_2961,In_967);
nand U5346 (N_5346,In_3587,In_4378);
xnor U5347 (N_5347,In_3099,In_3988);
nand U5348 (N_5348,In_3325,In_1840);
nor U5349 (N_5349,In_1413,In_1009);
and U5350 (N_5350,In_2385,In_4377);
xnor U5351 (N_5351,In_923,In_4924);
xnor U5352 (N_5352,In_1694,In_2562);
nand U5353 (N_5353,In_2063,In_4679);
nand U5354 (N_5354,In_316,In_2687);
xnor U5355 (N_5355,In_2371,In_334);
nand U5356 (N_5356,In_1994,In_2463);
xnor U5357 (N_5357,In_1065,In_3240);
nand U5358 (N_5358,In_286,In_253);
nor U5359 (N_5359,In_2388,In_4551);
nand U5360 (N_5360,In_4099,In_4440);
nand U5361 (N_5361,In_289,In_4803);
nand U5362 (N_5362,In_4165,In_133);
xor U5363 (N_5363,In_2564,In_1618);
or U5364 (N_5364,In_3956,In_1065);
nand U5365 (N_5365,In_2489,In_3417);
xor U5366 (N_5366,In_4223,In_3580);
nand U5367 (N_5367,In_4931,In_4043);
nor U5368 (N_5368,In_3707,In_4081);
xor U5369 (N_5369,In_3267,In_1192);
xnor U5370 (N_5370,In_423,In_4955);
nand U5371 (N_5371,In_1109,In_4529);
nand U5372 (N_5372,In_3790,In_1745);
xor U5373 (N_5373,In_2932,In_1961);
xnor U5374 (N_5374,In_4587,In_493);
nand U5375 (N_5375,In_277,In_2475);
xnor U5376 (N_5376,In_2518,In_1182);
xnor U5377 (N_5377,In_580,In_3364);
xnor U5378 (N_5378,In_4719,In_2380);
nand U5379 (N_5379,In_4339,In_339);
nand U5380 (N_5380,In_762,In_3732);
nor U5381 (N_5381,In_4700,In_1478);
or U5382 (N_5382,In_4601,In_1625);
or U5383 (N_5383,In_3223,In_2847);
and U5384 (N_5384,In_2640,In_687);
or U5385 (N_5385,In_4193,In_1972);
and U5386 (N_5386,In_411,In_2303);
nand U5387 (N_5387,In_1794,In_2488);
or U5388 (N_5388,In_3130,In_1008);
nand U5389 (N_5389,In_2399,In_140);
nor U5390 (N_5390,In_4243,In_2897);
nor U5391 (N_5391,In_2741,In_4551);
or U5392 (N_5392,In_4285,In_2675);
and U5393 (N_5393,In_605,In_1106);
or U5394 (N_5394,In_279,In_2772);
and U5395 (N_5395,In_2166,In_4779);
nand U5396 (N_5396,In_4520,In_864);
or U5397 (N_5397,In_1481,In_1690);
xnor U5398 (N_5398,In_2299,In_3280);
and U5399 (N_5399,In_1925,In_1038);
xnor U5400 (N_5400,In_417,In_4391);
nand U5401 (N_5401,In_522,In_110);
xnor U5402 (N_5402,In_216,In_2775);
nor U5403 (N_5403,In_46,In_126);
and U5404 (N_5404,In_4130,In_3787);
or U5405 (N_5405,In_760,In_2293);
or U5406 (N_5406,In_1157,In_346);
or U5407 (N_5407,In_3163,In_570);
and U5408 (N_5408,In_2767,In_194);
xor U5409 (N_5409,In_557,In_307);
and U5410 (N_5410,In_642,In_2156);
or U5411 (N_5411,In_1987,In_1679);
nor U5412 (N_5412,In_1,In_2552);
and U5413 (N_5413,In_947,In_2031);
nor U5414 (N_5414,In_2165,In_4141);
xnor U5415 (N_5415,In_3249,In_4672);
nand U5416 (N_5416,In_90,In_3331);
and U5417 (N_5417,In_3447,In_3873);
or U5418 (N_5418,In_4391,In_3882);
and U5419 (N_5419,In_4001,In_3808);
and U5420 (N_5420,In_4214,In_3044);
and U5421 (N_5421,In_1126,In_3710);
nand U5422 (N_5422,In_1,In_1905);
nor U5423 (N_5423,In_2477,In_246);
xor U5424 (N_5424,In_811,In_248);
nor U5425 (N_5425,In_3082,In_925);
nand U5426 (N_5426,In_945,In_2688);
and U5427 (N_5427,In_4873,In_4251);
nor U5428 (N_5428,In_4329,In_3402);
nand U5429 (N_5429,In_2701,In_4301);
xor U5430 (N_5430,In_2058,In_1474);
nand U5431 (N_5431,In_4575,In_864);
xor U5432 (N_5432,In_4876,In_3884);
or U5433 (N_5433,In_3010,In_960);
xor U5434 (N_5434,In_0,In_1798);
xor U5435 (N_5435,In_2127,In_3964);
nand U5436 (N_5436,In_3159,In_3826);
or U5437 (N_5437,In_1813,In_1965);
xor U5438 (N_5438,In_1277,In_52);
nand U5439 (N_5439,In_4549,In_1013);
xor U5440 (N_5440,In_1960,In_3538);
and U5441 (N_5441,In_4507,In_1020);
nor U5442 (N_5442,In_3005,In_1523);
or U5443 (N_5443,In_4048,In_999);
nand U5444 (N_5444,In_1287,In_1615);
and U5445 (N_5445,In_3733,In_2153);
or U5446 (N_5446,In_4834,In_1901);
or U5447 (N_5447,In_3905,In_2646);
xnor U5448 (N_5448,In_3887,In_209);
and U5449 (N_5449,In_3056,In_367);
and U5450 (N_5450,In_3383,In_2641);
and U5451 (N_5451,In_2706,In_4523);
and U5452 (N_5452,In_933,In_368);
nor U5453 (N_5453,In_503,In_1657);
or U5454 (N_5454,In_628,In_4416);
nand U5455 (N_5455,In_2471,In_3370);
nand U5456 (N_5456,In_2761,In_3022);
nor U5457 (N_5457,In_4798,In_2438);
nand U5458 (N_5458,In_587,In_1428);
nand U5459 (N_5459,In_626,In_4498);
or U5460 (N_5460,In_4755,In_2302);
nor U5461 (N_5461,In_1124,In_1026);
nand U5462 (N_5462,In_3501,In_562);
nor U5463 (N_5463,In_450,In_2201);
and U5464 (N_5464,In_3289,In_3821);
nand U5465 (N_5465,In_4787,In_3298);
or U5466 (N_5466,In_1566,In_1147);
and U5467 (N_5467,In_1586,In_68);
xor U5468 (N_5468,In_1016,In_464);
nor U5469 (N_5469,In_2889,In_3812);
xor U5470 (N_5470,In_4562,In_1666);
or U5471 (N_5471,In_956,In_208);
xnor U5472 (N_5472,In_4224,In_1566);
nor U5473 (N_5473,In_3496,In_1940);
and U5474 (N_5474,In_731,In_4846);
xnor U5475 (N_5475,In_2807,In_4856);
or U5476 (N_5476,In_2417,In_3669);
nor U5477 (N_5477,In_3269,In_224);
nor U5478 (N_5478,In_599,In_1923);
and U5479 (N_5479,In_2724,In_3186);
or U5480 (N_5480,In_3268,In_1361);
nor U5481 (N_5481,In_1635,In_3483);
xnor U5482 (N_5482,In_1747,In_2703);
or U5483 (N_5483,In_37,In_838);
xnor U5484 (N_5484,In_1081,In_787);
and U5485 (N_5485,In_231,In_3448);
and U5486 (N_5486,In_4336,In_4052);
and U5487 (N_5487,In_3098,In_2632);
and U5488 (N_5488,In_2654,In_58);
xor U5489 (N_5489,In_655,In_1778);
and U5490 (N_5490,In_4553,In_1443);
xnor U5491 (N_5491,In_3727,In_1399);
xor U5492 (N_5492,In_1550,In_2415);
or U5493 (N_5493,In_4145,In_251);
and U5494 (N_5494,In_4195,In_910);
nor U5495 (N_5495,In_2371,In_172);
xor U5496 (N_5496,In_1718,In_900);
and U5497 (N_5497,In_2234,In_3858);
nand U5498 (N_5498,In_1853,In_2066);
and U5499 (N_5499,In_4768,In_851);
xnor U5500 (N_5500,In_2808,In_3096);
nand U5501 (N_5501,In_3076,In_3487);
nor U5502 (N_5502,In_1803,In_1257);
xnor U5503 (N_5503,In_3661,In_4942);
and U5504 (N_5504,In_1045,In_856);
and U5505 (N_5505,In_3353,In_2730);
or U5506 (N_5506,In_4045,In_1690);
xnor U5507 (N_5507,In_358,In_2577);
and U5508 (N_5508,In_2846,In_1076);
xnor U5509 (N_5509,In_1636,In_3115);
and U5510 (N_5510,In_2650,In_2023);
or U5511 (N_5511,In_691,In_608);
and U5512 (N_5512,In_4536,In_2200);
nor U5513 (N_5513,In_3354,In_1802);
xnor U5514 (N_5514,In_3582,In_4019);
xnor U5515 (N_5515,In_340,In_691);
xnor U5516 (N_5516,In_2110,In_2798);
and U5517 (N_5517,In_2153,In_3467);
nor U5518 (N_5518,In_3904,In_2800);
or U5519 (N_5519,In_3918,In_4496);
nand U5520 (N_5520,In_2610,In_3229);
and U5521 (N_5521,In_4829,In_97);
and U5522 (N_5522,In_2641,In_1680);
nor U5523 (N_5523,In_1173,In_2803);
nor U5524 (N_5524,In_4953,In_909);
or U5525 (N_5525,In_3525,In_4156);
nor U5526 (N_5526,In_4918,In_733);
nand U5527 (N_5527,In_410,In_4698);
and U5528 (N_5528,In_1932,In_1855);
and U5529 (N_5529,In_440,In_585);
nor U5530 (N_5530,In_3999,In_4715);
xnor U5531 (N_5531,In_2557,In_4364);
and U5532 (N_5532,In_1209,In_424);
nand U5533 (N_5533,In_3380,In_1940);
or U5534 (N_5534,In_1140,In_1671);
nor U5535 (N_5535,In_3944,In_4447);
nand U5536 (N_5536,In_2114,In_3224);
nor U5537 (N_5537,In_4675,In_3528);
xor U5538 (N_5538,In_1305,In_71);
xor U5539 (N_5539,In_998,In_4544);
nor U5540 (N_5540,In_1048,In_4964);
nor U5541 (N_5541,In_3140,In_3104);
or U5542 (N_5542,In_3172,In_2277);
xor U5543 (N_5543,In_1873,In_589);
xor U5544 (N_5544,In_18,In_2010);
or U5545 (N_5545,In_4992,In_4168);
nor U5546 (N_5546,In_438,In_4155);
and U5547 (N_5547,In_2882,In_4662);
and U5548 (N_5548,In_1634,In_3971);
or U5549 (N_5549,In_641,In_699);
nand U5550 (N_5550,In_488,In_206);
xor U5551 (N_5551,In_153,In_4975);
nand U5552 (N_5552,In_2751,In_3465);
nor U5553 (N_5553,In_4016,In_3965);
xor U5554 (N_5554,In_2309,In_1473);
or U5555 (N_5555,In_3606,In_2718);
nand U5556 (N_5556,In_1525,In_731);
xor U5557 (N_5557,In_3890,In_4145);
xor U5558 (N_5558,In_1009,In_3767);
nand U5559 (N_5559,In_4450,In_2868);
nor U5560 (N_5560,In_817,In_4802);
nor U5561 (N_5561,In_4230,In_1611);
xnor U5562 (N_5562,In_2503,In_573);
nor U5563 (N_5563,In_120,In_2974);
nand U5564 (N_5564,In_789,In_3612);
nand U5565 (N_5565,In_1601,In_2165);
xnor U5566 (N_5566,In_4502,In_2653);
xnor U5567 (N_5567,In_2881,In_2231);
nand U5568 (N_5568,In_185,In_4762);
nand U5569 (N_5569,In_734,In_4434);
nor U5570 (N_5570,In_3090,In_4310);
or U5571 (N_5571,In_4776,In_2369);
nor U5572 (N_5572,In_4962,In_3574);
xor U5573 (N_5573,In_813,In_1652);
nand U5574 (N_5574,In_4818,In_2717);
and U5575 (N_5575,In_3776,In_1113);
nand U5576 (N_5576,In_317,In_4033);
and U5577 (N_5577,In_1329,In_2594);
or U5578 (N_5578,In_406,In_947);
nand U5579 (N_5579,In_1546,In_248);
nand U5580 (N_5580,In_4934,In_1119);
nor U5581 (N_5581,In_3798,In_1582);
nand U5582 (N_5582,In_778,In_236);
and U5583 (N_5583,In_718,In_3006);
nand U5584 (N_5584,In_4036,In_90);
nand U5585 (N_5585,In_2837,In_1247);
xnor U5586 (N_5586,In_2711,In_1740);
and U5587 (N_5587,In_3997,In_4718);
and U5588 (N_5588,In_2520,In_4546);
xor U5589 (N_5589,In_4373,In_4061);
xor U5590 (N_5590,In_2276,In_3711);
nand U5591 (N_5591,In_4534,In_2958);
or U5592 (N_5592,In_1283,In_3202);
xnor U5593 (N_5593,In_4426,In_4520);
or U5594 (N_5594,In_3026,In_4116);
nor U5595 (N_5595,In_3721,In_2565);
nand U5596 (N_5596,In_2869,In_4212);
xor U5597 (N_5597,In_3249,In_431);
nand U5598 (N_5598,In_1501,In_2323);
or U5599 (N_5599,In_3459,In_1276);
nand U5600 (N_5600,In_330,In_2191);
and U5601 (N_5601,In_1572,In_1737);
xor U5602 (N_5602,In_1882,In_1489);
nand U5603 (N_5603,In_3962,In_657);
and U5604 (N_5604,In_4476,In_143);
nor U5605 (N_5605,In_3177,In_284);
nand U5606 (N_5606,In_4691,In_2989);
xnor U5607 (N_5607,In_695,In_4451);
nand U5608 (N_5608,In_2758,In_3186);
or U5609 (N_5609,In_1269,In_2165);
xor U5610 (N_5610,In_1770,In_3842);
and U5611 (N_5611,In_2463,In_2326);
or U5612 (N_5612,In_133,In_417);
and U5613 (N_5613,In_2051,In_3575);
nor U5614 (N_5614,In_4890,In_4838);
and U5615 (N_5615,In_2628,In_3876);
nand U5616 (N_5616,In_4507,In_271);
and U5617 (N_5617,In_2447,In_4827);
and U5618 (N_5618,In_3246,In_1496);
or U5619 (N_5619,In_2004,In_286);
nor U5620 (N_5620,In_3632,In_4172);
nor U5621 (N_5621,In_3638,In_4807);
or U5622 (N_5622,In_2190,In_4492);
and U5623 (N_5623,In_4195,In_4409);
xnor U5624 (N_5624,In_1027,In_328);
xor U5625 (N_5625,In_670,In_731);
and U5626 (N_5626,In_4536,In_4006);
nand U5627 (N_5627,In_383,In_3915);
or U5628 (N_5628,In_1720,In_3274);
nand U5629 (N_5629,In_3409,In_1392);
nor U5630 (N_5630,In_1092,In_4881);
xor U5631 (N_5631,In_4979,In_3727);
or U5632 (N_5632,In_2280,In_2689);
and U5633 (N_5633,In_2767,In_3717);
nor U5634 (N_5634,In_4013,In_2802);
nand U5635 (N_5635,In_1207,In_4046);
or U5636 (N_5636,In_3040,In_315);
and U5637 (N_5637,In_1117,In_3133);
and U5638 (N_5638,In_2486,In_1357);
or U5639 (N_5639,In_3847,In_2363);
or U5640 (N_5640,In_445,In_4354);
nand U5641 (N_5641,In_2505,In_4622);
nor U5642 (N_5642,In_1626,In_4485);
nand U5643 (N_5643,In_179,In_2074);
nor U5644 (N_5644,In_672,In_342);
or U5645 (N_5645,In_3749,In_2799);
and U5646 (N_5646,In_3569,In_223);
nor U5647 (N_5647,In_4402,In_3153);
xor U5648 (N_5648,In_3463,In_975);
nor U5649 (N_5649,In_4465,In_4954);
or U5650 (N_5650,In_2449,In_2041);
nor U5651 (N_5651,In_2962,In_236);
or U5652 (N_5652,In_4464,In_86);
or U5653 (N_5653,In_1901,In_2124);
and U5654 (N_5654,In_4605,In_3503);
xor U5655 (N_5655,In_2587,In_1678);
nor U5656 (N_5656,In_2275,In_2105);
or U5657 (N_5657,In_3237,In_4457);
or U5658 (N_5658,In_695,In_1636);
xnor U5659 (N_5659,In_2382,In_4138);
and U5660 (N_5660,In_706,In_321);
and U5661 (N_5661,In_715,In_4026);
or U5662 (N_5662,In_2993,In_3105);
nor U5663 (N_5663,In_374,In_2027);
nor U5664 (N_5664,In_3373,In_1171);
nor U5665 (N_5665,In_3434,In_3917);
nor U5666 (N_5666,In_3727,In_3491);
xor U5667 (N_5667,In_584,In_957);
xor U5668 (N_5668,In_1211,In_774);
or U5669 (N_5669,In_4609,In_1932);
and U5670 (N_5670,In_4205,In_1277);
xnor U5671 (N_5671,In_2289,In_3025);
nor U5672 (N_5672,In_1157,In_671);
or U5673 (N_5673,In_226,In_758);
nand U5674 (N_5674,In_2059,In_2733);
xnor U5675 (N_5675,In_2547,In_2086);
and U5676 (N_5676,In_1693,In_1871);
nor U5677 (N_5677,In_2119,In_2184);
xor U5678 (N_5678,In_4607,In_973);
nand U5679 (N_5679,In_3719,In_1403);
nor U5680 (N_5680,In_2058,In_1765);
xnor U5681 (N_5681,In_614,In_2302);
or U5682 (N_5682,In_2140,In_2082);
xor U5683 (N_5683,In_681,In_3044);
nand U5684 (N_5684,In_2797,In_2871);
nor U5685 (N_5685,In_3124,In_2801);
nand U5686 (N_5686,In_3235,In_4337);
nor U5687 (N_5687,In_793,In_980);
and U5688 (N_5688,In_1902,In_3116);
nor U5689 (N_5689,In_4394,In_472);
and U5690 (N_5690,In_4887,In_876);
nand U5691 (N_5691,In_2492,In_4171);
nor U5692 (N_5692,In_895,In_866);
nand U5693 (N_5693,In_3073,In_3772);
nor U5694 (N_5694,In_4547,In_2710);
nor U5695 (N_5695,In_1376,In_3194);
xor U5696 (N_5696,In_115,In_3745);
nor U5697 (N_5697,In_3506,In_2608);
nand U5698 (N_5698,In_3250,In_3150);
nand U5699 (N_5699,In_237,In_861);
nor U5700 (N_5700,In_1745,In_4853);
nor U5701 (N_5701,In_1474,In_529);
xor U5702 (N_5702,In_2948,In_2181);
nand U5703 (N_5703,In_4435,In_3357);
or U5704 (N_5704,In_4876,In_2437);
nor U5705 (N_5705,In_4633,In_1014);
nand U5706 (N_5706,In_274,In_4231);
nand U5707 (N_5707,In_2729,In_4563);
nand U5708 (N_5708,In_3871,In_1580);
or U5709 (N_5709,In_4080,In_3360);
nand U5710 (N_5710,In_4455,In_4586);
and U5711 (N_5711,In_2057,In_612);
xnor U5712 (N_5712,In_4716,In_66);
nand U5713 (N_5713,In_899,In_819);
and U5714 (N_5714,In_686,In_1538);
nand U5715 (N_5715,In_2274,In_2079);
or U5716 (N_5716,In_2437,In_967);
nand U5717 (N_5717,In_605,In_724);
nor U5718 (N_5718,In_2153,In_1053);
or U5719 (N_5719,In_1243,In_1930);
or U5720 (N_5720,In_3762,In_804);
nand U5721 (N_5721,In_2032,In_4397);
xnor U5722 (N_5722,In_1237,In_3270);
nor U5723 (N_5723,In_4878,In_2359);
and U5724 (N_5724,In_1147,In_2558);
nor U5725 (N_5725,In_3451,In_4438);
nor U5726 (N_5726,In_2835,In_2356);
nand U5727 (N_5727,In_2207,In_2970);
xor U5728 (N_5728,In_3488,In_2127);
and U5729 (N_5729,In_4683,In_955);
or U5730 (N_5730,In_3000,In_4304);
nor U5731 (N_5731,In_3686,In_297);
nor U5732 (N_5732,In_829,In_910);
and U5733 (N_5733,In_735,In_4339);
xor U5734 (N_5734,In_4024,In_4530);
nor U5735 (N_5735,In_4630,In_1622);
and U5736 (N_5736,In_2253,In_4970);
nor U5737 (N_5737,In_905,In_2282);
xor U5738 (N_5738,In_2708,In_1548);
nor U5739 (N_5739,In_2205,In_2153);
or U5740 (N_5740,In_2908,In_1726);
xor U5741 (N_5741,In_3743,In_2926);
and U5742 (N_5742,In_799,In_804);
nor U5743 (N_5743,In_939,In_4541);
nand U5744 (N_5744,In_4341,In_2015);
nor U5745 (N_5745,In_2293,In_2870);
xor U5746 (N_5746,In_4927,In_4009);
xnor U5747 (N_5747,In_1646,In_3004);
xor U5748 (N_5748,In_762,In_1002);
and U5749 (N_5749,In_2462,In_3086);
and U5750 (N_5750,In_2952,In_153);
or U5751 (N_5751,In_2397,In_2859);
and U5752 (N_5752,In_3741,In_4044);
nor U5753 (N_5753,In_856,In_1941);
nor U5754 (N_5754,In_432,In_4923);
nor U5755 (N_5755,In_3899,In_1137);
xor U5756 (N_5756,In_4771,In_3683);
xnor U5757 (N_5757,In_4779,In_4980);
nand U5758 (N_5758,In_4027,In_2079);
nand U5759 (N_5759,In_4287,In_2385);
nor U5760 (N_5760,In_3874,In_3877);
nand U5761 (N_5761,In_4229,In_4984);
nor U5762 (N_5762,In_3251,In_3719);
nor U5763 (N_5763,In_3992,In_4589);
nor U5764 (N_5764,In_4685,In_1166);
nand U5765 (N_5765,In_1654,In_2057);
and U5766 (N_5766,In_4916,In_2514);
or U5767 (N_5767,In_1689,In_2719);
nor U5768 (N_5768,In_1942,In_483);
xor U5769 (N_5769,In_3042,In_3482);
nor U5770 (N_5770,In_1250,In_582);
nand U5771 (N_5771,In_3999,In_1172);
or U5772 (N_5772,In_4489,In_3825);
and U5773 (N_5773,In_2926,In_4086);
nor U5774 (N_5774,In_3741,In_58);
and U5775 (N_5775,In_2832,In_468);
and U5776 (N_5776,In_1993,In_158);
nor U5777 (N_5777,In_2068,In_3514);
nand U5778 (N_5778,In_134,In_4280);
nor U5779 (N_5779,In_3442,In_2519);
nand U5780 (N_5780,In_3538,In_1415);
xnor U5781 (N_5781,In_2355,In_1869);
and U5782 (N_5782,In_1821,In_458);
xor U5783 (N_5783,In_4702,In_2842);
or U5784 (N_5784,In_957,In_3426);
nand U5785 (N_5785,In_1123,In_3744);
and U5786 (N_5786,In_999,In_3428);
or U5787 (N_5787,In_2119,In_539);
nor U5788 (N_5788,In_4985,In_3682);
xnor U5789 (N_5789,In_396,In_2467);
nand U5790 (N_5790,In_4198,In_1624);
nand U5791 (N_5791,In_763,In_243);
and U5792 (N_5792,In_1749,In_837);
or U5793 (N_5793,In_3386,In_2169);
and U5794 (N_5794,In_3679,In_4805);
and U5795 (N_5795,In_3177,In_4972);
xor U5796 (N_5796,In_4501,In_4538);
or U5797 (N_5797,In_2482,In_4774);
nor U5798 (N_5798,In_1494,In_2164);
or U5799 (N_5799,In_4648,In_3826);
nor U5800 (N_5800,In_1473,In_2946);
or U5801 (N_5801,In_2723,In_4297);
nand U5802 (N_5802,In_1853,In_838);
and U5803 (N_5803,In_4331,In_3398);
and U5804 (N_5804,In_2522,In_3744);
xor U5805 (N_5805,In_4545,In_4809);
and U5806 (N_5806,In_3932,In_1683);
or U5807 (N_5807,In_1197,In_1376);
nand U5808 (N_5808,In_3010,In_2766);
or U5809 (N_5809,In_1884,In_1829);
nand U5810 (N_5810,In_2276,In_1227);
nor U5811 (N_5811,In_1865,In_434);
nand U5812 (N_5812,In_4284,In_1075);
and U5813 (N_5813,In_3484,In_3429);
and U5814 (N_5814,In_1639,In_3540);
nor U5815 (N_5815,In_817,In_3363);
nand U5816 (N_5816,In_1721,In_377);
nand U5817 (N_5817,In_4509,In_3968);
xor U5818 (N_5818,In_3741,In_4796);
or U5819 (N_5819,In_674,In_1269);
nand U5820 (N_5820,In_2836,In_4370);
and U5821 (N_5821,In_1316,In_1754);
xor U5822 (N_5822,In_3200,In_2272);
or U5823 (N_5823,In_1570,In_4026);
nand U5824 (N_5824,In_2534,In_3606);
nor U5825 (N_5825,In_1304,In_2860);
or U5826 (N_5826,In_2124,In_512);
xor U5827 (N_5827,In_3736,In_4888);
nand U5828 (N_5828,In_4320,In_4164);
and U5829 (N_5829,In_2227,In_1623);
or U5830 (N_5830,In_4566,In_870);
and U5831 (N_5831,In_3659,In_3083);
nor U5832 (N_5832,In_4660,In_1669);
nor U5833 (N_5833,In_4316,In_4808);
and U5834 (N_5834,In_700,In_1539);
nor U5835 (N_5835,In_4090,In_1479);
nand U5836 (N_5836,In_2373,In_1864);
xnor U5837 (N_5837,In_4696,In_2846);
nor U5838 (N_5838,In_3002,In_2590);
xnor U5839 (N_5839,In_3841,In_4785);
and U5840 (N_5840,In_64,In_3029);
or U5841 (N_5841,In_3182,In_1715);
nand U5842 (N_5842,In_3205,In_1655);
xnor U5843 (N_5843,In_367,In_1720);
nor U5844 (N_5844,In_287,In_2013);
nand U5845 (N_5845,In_3436,In_4449);
nand U5846 (N_5846,In_35,In_2913);
nand U5847 (N_5847,In_1453,In_3500);
xnor U5848 (N_5848,In_3237,In_63);
nand U5849 (N_5849,In_2543,In_185);
nor U5850 (N_5850,In_1209,In_3207);
xnor U5851 (N_5851,In_1880,In_725);
nor U5852 (N_5852,In_3148,In_4585);
nor U5853 (N_5853,In_802,In_3903);
nor U5854 (N_5854,In_192,In_4431);
nand U5855 (N_5855,In_1063,In_744);
xnor U5856 (N_5856,In_4389,In_3911);
or U5857 (N_5857,In_3625,In_1613);
nor U5858 (N_5858,In_3025,In_1237);
xor U5859 (N_5859,In_293,In_3589);
nand U5860 (N_5860,In_638,In_4879);
or U5861 (N_5861,In_4243,In_2915);
xor U5862 (N_5862,In_2794,In_4894);
and U5863 (N_5863,In_282,In_2741);
nor U5864 (N_5864,In_4260,In_2060);
nor U5865 (N_5865,In_268,In_2596);
nor U5866 (N_5866,In_3739,In_2459);
or U5867 (N_5867,In_3952,In_1717);
nand U5868 (N_5868,In_610,In_227);
and U5869 (N_5869,In_3488,In_955);
or U5870 (N_5870,In_3944,In_1855);
or U5871 (N_5871,In_2148,In_1149);
nand U5872 (N_5872,In_3096,In_1409);
nand U5873 (N_5873,In_3029,In_533);
or U5874 (N_5874,In_253,In_83);
xor U5875 (N_5875,In_4612,In_1120);
and U5876 (N_5876,In_63,In_1379);
nand U5877 (N_5877,In_4776,In_3236);
or U5878 (N_5878,In_3790,In_501);
xnor U5879 (N_5879,In_4206,In_4768);
xnor U5880 (N_5880,In_2835,In_268);
xor U5881 (N_5881,In_2414,In_1643);
or U5882 (N_5882,In_2239,In_1382);
xnor U5883 (N_5883,In_2748,In_2346);
xor U5884 (N_5884,In_3501,In_2830);
or U5885 (N_5885,In_254,In_1930);
or U5886 (N_5886,In_4710,In_1724);
nand U5887 (N_5887,In_763,In_534);
xor U5888 (N_5888,In_3360,In_870);
nand U5889 (N_5889,In_3547,In_949);
xnor U5890 (N_5890,In_2113,In_3614);
nand U5891 (N_5891,In_2655,In_2660);
nand U5892 (N_5892,In_4078,In_2056);
and U5893 (N_5893,In_4693,In_4655);
or U5894 (N_5894,In_3004,In_342);
nand U5895 (N_5895,In_1796,In_2724);
or U5896 (N_5896,In_401,In_1574);
nor U5897 (N_5897,In_4599,In_2847);
nor U5898 (N_5898,In_4791,In_2434);
or U5899 (N_5899,In_3064,In_1258);
nor U5900 (N_5900,In_3173,In_2884);
nor U5901 (N_5901,In_1750,In_3231);
nand U5902 (N_5902,In_2015,In_3122);
nor U5903 (N_5903,In_4201,In_1212);
nor U5904 (N_5904,In_1579,In_1192);
xor U5905 (N_5905,In_972,In_2388);
nand U5906 (N_5906,In_1957,In_2643);
or U5907 (N_5907,In_3540,In_1408);
and U5908 (N_5908,In_2228,In_1874);
or U5909 (N_5909,In_2335,In_4603);
nor U5910 (N_5910,In_793,In_3896);
nand U5911 (N_5911,In_651,In_1128);
xnor U5912 (N_5912,In_3637,In_1568);
nand U5913 (N_5913,In_327,In_4677);
and U5914 (N_5914,In_575,In_211);
nor U5915 (N_5915,In_3076,In_4407);
and U5916 (N_5916,In_4371,In_2500);
or U5917 (N_5917,In_3497,In_4348);
or U5918 (N_5918,In_303,In_3219);
xnor U5919 (N_5919,In_3523,In_1616);
nor U5920 (N_5920,In_2577,In_3132);
or U5921 (N_5921,In_3288,In_2357);
nor U5922 (N_5922,In_4006,In_1586);
xnor U5923 (N_5923,In_4454,In_3689);
nand U5924 (N_5924,In_3066,In_3593);
and U5925 (N_5925,In_2955,In_2561);
nand U5926 (N_5926,In_372,In_1715);
or U5927 (N_5927,In_4952,In_3971);
nor U5928 (N_5928,In_3989,In_1569);
and U5929 (N_5929,In_1222,In_912);
and U5930 (N_5930,In_4777,In_3930);
xor U5931 (N_5931,In_1849,In_3744);
xnor U5932 (N_5932,In_4840,In_2528);
nand U5933 (N_5933,In_1303,In_3707);
nor U5934 (N_5934,In_4796,In_3116);
nand U5935 (N_5935,In_4075,In_1323);
and U5936 (N_5936,In_711,In_4500);
nor U5937 (N_5937,In_688,In_580);
xor U5938 (N_5938,In_4076,In_3322);
or U5939 (N_5939,In_3151,In_4119);
and U5940 (N_5940,In_2954,In_1613);
and U5941 (N_5941,In_1139,In_854);
xnor U5942 (N_5942,In_1137,In_3903);
xnor U5943 (N_5943,In_1177,In_3723);
and U5944 (N_5944,In_2665,In_1568);
xnor U5945 (N_5945,In_1291,In_4073);
or U5946 (N_5946,In_3770,In_921);
nor U5947 (N_5947,In_2039,In_4635);
or U5948 (N_5948,In_1141,In_2054);
nor U5949 (N_5949,In_4304,In_1967);
nand U5950 (N_5950,In_1225,In_3432);
nor U5951 (N_5951,In_4804,In_4326);
nand U5952 (N_5952,In_3827,In_4163);
nand U5953 (N_5953,In_1145,In_1175);
or U5954 (N_5954,In_2931,In_3577);
nor U5955 (N_5955,In_2441,In_4545);
xor U5956 (N_5956,In_4291,In_0);
or U5957 (N_5957,In_652,In_333);
nor U5958 (N_5958,In_241,In_1987);
and U5959 (N_5959,In_4852,In_1181);
nand U5960 (N_5960,In_4764,In_4965);
nor U5961 (N_5961,In_914,In_1135);
nor U5962 (N_5962,In_747,In_413);
xnor U5963 (N_5963,In_977,In_3614);
or U5964 (N_5964,In_1641,In_687);
xor U5965 (N_5965,In_1952,In_963);
xor U5966 (N_5966,In_896,In_2853);
or U5967 (N_5967,In_201,In_4915);
or U5968 (N_5968,In_4344,In_1896);
nand U5969 (N_5969,In_3499,In_816);
or U5970 (N_5970,In_2971,In_168);
nor U5971 (N_5971,In_1681,In_2939);
xor U5972 (N_5972,In_4485,In_2602);
nand U5973 (N_5973,In_1590,In_3024);
or U5974 (N_5974,In_4238,In_3542);
xor U5975 (N_5975,In_2936,In_1131);
or U5976 (N_5976,In_2549,In_4531);
nor U5977 (N_5977,In_754,In_469);
nand U5978 (N_5978,In_3561,In_3391);
and U5979 (N_5979,In_2835,In_3101);
xnor U5980 (N_5980,In_971,In_1563);
xor U5981 (N_5981,In_3579,In_1077);
xor U5982 (N_5982,In_1698,In_439);
xor U5983 (N_5983,In_3706,In_1217);
and U5984 (N_5984,In_4671,In_592);
nand U5985 (N_5985,In_846,In_3833);
or U5986 (N_5986,In_2835,In_1486);
nand U5987 (N_5987,In_4784,In_933);
nor U5988 (N_5988,In_210,In_1712);
xnor U5989 (N_5989,In_1557,In_4428);
xor U5990 (N_5990,In_2864,In_916);
and U5991 (N_5991,In_1390,In_2509);
nand U5992 (N_5992,In_2044,In_769);
nor U5993 (N_5993,In_2152,In_2303);
and U5994 (N_5994,In_1480,In_4495);
or U5995 (N_5995,In_4205,In_4552);
or U5996 (N_5996,In_755,In_3170);
or U5997 (N_5997,In_3676,In_3435);
nand U5998 (N_5998,In_4465,In_3877);
or U5999 (N_5999,In_1266,In_1196);
and U6000 (N_6000,In_1302,In_638);
xor U6001 (N_6001,In_3998,In_663);
xnor U6002 (N_6002,In_463,In_3635);
and U6003 (N_6003,In_1900,In_889);
nand U6004 (N_6004,In_2458,In_2640);
xor U6005 (N_6005,In_1430,In_1995);
xnor U6006 (N_6006,In_3059,In_4348);
nor U6007 (N_6007,In_3041,In_4156);
nor U6008 (N_6008,In_1298,In_4479);
xnor U6009 (N_6009,In_2799,In_146);
nand U6010 (N_6010,In_627,In_545);
nor U6011 (N_6011,In_4004,In_3708);
nand U6012 (N_6012,In_1697,In_3863);
nand U6013 (N_6013,In_460,In_2719);
and U6014 (N_6014,In_2047,In_591);
or U6015 (N_6015,In_3865,In_4609);
xor U6016 (N_6016,In_3409,In_4736);
nor U6017 (N_6017,In_2769,In_3495);
nand U6018 (N_6018,In_3326,In_3580);
or U6019 (N_6019,In_1577,In_3886);
nor U6020 (N_6020,In_2919,In_1197);
xor U6021 (N_6021,In_1954,In_1260);
and U6022 (N_6022,In_3680,In_834);
nand U6023 (N_6023,In_4734,In_1344);
and U6024 (N_6024,In_489,In_3678);
and U6025 (N_6025,In_1304,In_1359);
or U6026 (N_6026,In_386,In_567);
or U6027 (N_6027,In_1716,In_3734);
and U6028 (N_6028,In_3751,In_1433);
and U6029 (N_6029,In_4837,In_1518);
nor U6030 (N_6030,In_4199,In_2697);
or U6031 (N_6031,In_3671,In_3896);
or U6032 (N_6032,In_105,In_3669);
nand U6033 (N_6033,In_3638,In_2143);
nand U6034 (N_6034,In_937,In_2391);
or U6035 (N_6035,In_508,In_4573);
or U6036 (N_6036,In_4213,In_268);
or U6037 (N_6037,In_3609,In_13);
nand U6038 (N_6038,In_3647,In_2631);
xnor U6039 (N_6039,In_3758,In_2326);
nand U6040 (N_6040,In_514,In_2525);
xor U6041 (N_6041,In_1314,In_1013);
and U6042 (N_6042,In_3190,In_1455);
and U6043 (N_6043,In_170,In_770);
and U6044 (N_6044,In_1768,In_2826);
xnor U6045 (N_6045,In_1072,In_4237);
or U6046 (N_6046,In_4971,In_2112);
nand U6047 (N_6047,In_2901,In_2040);
or U6048 (N_6048,In_934,In_4498);
xor U6049 (N_6049,In_2519,In_3631);
nor U6050 (N_6050,In_1698,In_2728);
or U6051 (N_6051,In_1176,In_3657);
or U6052 (N_6052,In_286,In_3005);
and U6053 (N_6053,In_1481,In_3682);
nor U6054 (N_6054,In_3334,In_440);
or U6055 (N_6055,In_154,In_1961);
or U6056 (N_6056,In_2409,In_3506);
or U6057 (N_6057,In_1029,In_2587);
nor U6058 (N_6058,In_4635,In_790);
nand U6059 (N_6059,In_1986,In_1379);
nor U6060 (N_6060,In_2460,In_4025);
nor U6061 (N_6061,In_2637,In_784);
and U6062 (N_6062,In_2881,In_1557);
xnor U6063 (N_6063,In_4224,In_2108);
or U6064 (N_6064,In_3064,In_2533);
and U6065 (N_6065,In_4538,In_1213);
nand U6066 (N_6066,In_443,In_62);
nand U6067 (N_6067,In_863,In_2224);
xor U6068 (N_6068,In_891,In_1781);
nand U6069 (N_6069,In_3731,In_1292);
and U6070 (N_6070,In_3822,In_2595);
xor U6071 (N_6071,In_1801,In_4051);
xnor U6072 (N_6072,In_4239,In_2563);
nor U6073 (N_6073,In_1853,In_4457);
or U6074 (N_6074,In_4831,In_1085);
or U6075 (N_6075,In_2715,In_842);
xnor U6076 (N_6076,In_1186,In_4057);
and U6077 (N_6077,In_2146,In_584);
or U6078 (N_6078,In_2023,In_4041);
and U6079 (N_6079,In_4988,In_1880);
xnor U6080 (N_6080,In_4886,In_2892);
or U6081 (N_6081,In_2596,In_2420);
nand U6082 (N_6082,In_1925,In_616);
and U6083 (N_6083,In_4495,In_979);
or U6084 (N_6084,In_3507,In_3965);
nor U6085 (N_6085,In_2701,In_1438);
and U6086 (N_6086,In_2831,In_4549);
nor U6087 (N_6087,In_3569,In_2721);
xor U6088 (N_6088,In_3674,In_252);
and U6089 (N_6089,In_782,In_3084);
nor U6090 (N_6090,In_1103,In_3459);
and U6091 (N_6091,In_3675,In_52);
or U6092 (N_6092,In_2776,In_1167);
nor U6093 (N_6093,In_3364,In_2562);
nand U6094 (N_6094,In_2616,In_4053);
xor U6095 (N_6095,In_2366,In_2944);
xnor U6096 (N_6096,In_4731,In_2492);
nand U6097 (N_6097,In_1385,In_3346);
nand U6098 (N_6098,In_2538,In_3432);
and U6099 (N_6099,In_3471,In_3706);
and U6100 (N_6100,In_104,In_4573);
xnor U6101 (N_6101,In_369,In_1364);
nor U6102 (N_6102,In_1590,In_230);
nand U6103 (N_6103,In_3904,In_4461);
xnor U6104 (N_6104,In_4190,In_3176);
or U6105 (N_6105,In_2704,In_659);
xor U6106 (N_6106,In_2882,In_3420);
nand U6107 (N_6107,In_4416,In_4399);
and U6108 (N_6108,In_161,In_3517);
and U6109 (N_6109,In_2274,In_2505);
and U6110 (N_6110,In_3341,In_3719);
nand U6111 (N_6111,In_1403,In_4234);
or U6112 (N_6112,In_612,In_4988);
and U6113 (N_6113,In_2503,In_3523);
xor U6114 (N_6114,In_4858,In_3332);
xor U6115 (N_6115,In_4389,In_4530);
xor U6116 (N_6116,In_4214,In_383);
nor U6117 (N_6117,In_1115,In_3686);
xnor U6118 (N_6118,In_628,In_4276);
nand U6119 (N_6119,In_2884,In_663);
xor U6120 (N_6120,In_1693,In_3066);
nand U6121 (N_6121,In_1284,In_4852);
nor U6122 (N_6122,In_4952,In_4480);
nor U6123 (N_6123,In_2814,In_3557);
xnor U6124 (N_6124,In_2945,In_3177);
and U6125 (N_6125,In_1500,In_3809);
nand U6126 (N_6126,In_3663,In_1898);
nand U6127 (N_6127,In_1040,In_1633);
and U6128 (N_6128,In_2122,In_2993);
nor U6129 (N_6129,In_3823,In_1079);
or U6130 (N_6130,In_431,In_2822);
nand U6131 (N_6131,In_1526,In_3505);
nor U6132 (N_6132,In_4727,In_2649);
nand U6133 (N_6133,In_2276,In_2682);
or U6134 (N_6134,In_1861,In_3800);
and U6135 (N_6135,In_2813,In_4312);
or U6136 (N_6136,In_3120,In_3846);
nor U6137 (N_6137,In_2166,In_1085);
and U6138 (N_6138,In_270,In_1189);
nand U6139 (N_6139,In_2644,In_2842);
or U6140 (N_6140,In_4280,In_2313);
and U6141 (N_6141,In_1792,In_1833);
nor U6142 (N_6142,In_1067,In_2845);
nand U6143 (N_6143,In_3057,In_3910);
or U6144 (N_6144,In_1968,In_672);
and U6145 (N_6145,In_4133,In_3645);
nor U6146 (N_6146,In_3967,In_3216);
or U6147 (N_6147,In_2881,In_2409);
nand U6148 (N_6148,In_58,In_3269);
xnor U6149 (N_6149,In_1952,In_4211);
xnor U6150 (N_6150,In_611,In_3725);
or U6151 (N_6151,In_4387,In_349);
xor U6152 (N_6152,In_1888,In_3515);
nand U6153 (N_6153,In_1033,In_2972);
xnor U6154 (N_6154,In_1526,In_3300);
xnor U6155 (N_6155,In_1165,In_2666);
nor U6156 (N_6156,In_3683,In_1822);
nor U6157 (N_6157,In_1041,In_2058);
and U6158 (N_6158,In_3379,In_2106);
and U6159 (N_6159,In_1469,In_2808);
xnor U6160 (N_6160,In_334,In_3938);
or U6161 (N_6161,In_2097,In_1986);
xor U6162 (N_6162,In_548,In_4565);
and U6163 (N_6163,In_1152,In_2035);
nor U6164 (N_6164,In_4356,In_1639);
and U6165 (N_6165,In_3645,In_2741);
nor U6166 (N_6166,In_1544,In_3512);
xor U6167 (N_6167,In_4298,In_4624);
xnor U6168 (N_6168,In_2585,In_889);
nand U6169 (N_6169,In_3109,In_3322);
and U6170 (N_6170,In_4001,In_1862);
or U6171 (N_6171,In_967,In_1535);
nand U6172 (N_6172,In_1613,In_2656);
nor U6173 (N_6173,In_22,In_3073);
and U6174 (N_6174,In_772,In_3790);
xor U6175 (N_6175,In_34,In_764);
or U6176 (N_6176,In_2316,In_4998);
xnor U6177 (N_6177,In_4451,In_4264);
nand U6178 (N_6178,In_1359,In_4894);
nor U6179 (N_6179,In_4024,In_1034);
and U6180 (N_6180,In_4348,In_1952);
or U6181 (N_6181,In_1509,In_3965);
or U6182 (N_6182,In_1951,In_1832);
or U6183 (N_6183,In_608,In_2474);
xnor U6184 (N_6184,In_4355,In_3860);
or U6185 (N_6185,In_13,In_4543);
or U6186 (N_6186,In_2412,In_2137);
and U6187 (N_6187,In_2170,In_1986);
xor U6188 (N_6188,In_1313,In_1587);
and U6189 (N_6189,In_3200,In_675);
xnor U6190 (N_6190,In_31,In_2144);
xor U6191 (N_6191,In_3381,In_3804);
xnor U6192 (N_6192,In_2652,In_942);
xnor U6193 (N_6193,In_1786,In_1468);
or U6194 (N_6194,In_1894,In_661);
nand U6195 (N_6195,In_1737,In_585);
nand U6196 (N_6196,In_2007,In_3021);
xnor U6197 (N_6197,In_3766,In_1255);
xor U6198 (N_6198,In_887,In_1069);
or U6199 (N_6199,In_925,In_3939);
and U6200 (N_6200,In_3335,In_3868);
and U6201 (N_6201,In_3071,In_229);
xor U6202 (N_6202,In_3512,In_447);
nor U6203 (N_6203,In_2801,In_2808);
or U6204 (N_6204,In_847,In_3014);
nand U6205 (N_6205,In_1593,In_4956);
nor U6206 (N_6206,In_1993,In_3284);
nand U6207 (N_6207,In_1639,In_1137);
or U6208 (N_6208,In_3453,In_785);
or U6209 (N_6209,In_4269,In_874);
or U6210 (N_6210,In_1120,In_4188);
xor U6211 (N_6211,In_1208,In_2610);
nand U6212 (N_6212,In_3021,In_2709);
nor U6213 (N_6213,In_2221,In_4040);
xnor U6214 (N_6214,In_4639,In_1040);
or U6215 (N_6215,In_4903,In_1115);
and U6216 (N_6216,In_1769,In_2245);
and U6217 (N_6217,In_4171,In_273);
nand U6218 (N_6218,In_2467,In_803);
xnor U6219 (N_6219,In_4710,In_1277);
xor U6220 (N_6220,In_1846,In_2401);
or U6221 (N_6221,In_2337,In_2612);
nand U6222 (N_6222,In_626,In_916);
nand U6223 (N_6223,In_4161,In_3519);
nor U6224 (N_6224,In_3259,In_1729);
nor U6225 (N_6225,In_1975,In_2347);
nor U6226 (N_6226,In_3957,In_4534);
xnor U6227 (N_6227,In_4275,In_333);
and U6228 (N_6228,In_3452,In_2398);
nand U6229 (N_6229,In_4503,In_1237);
or U6230 (N_6230,In_1296,In_4035);
and U6231 (N_6231,In_4706,In_4193);
nand U6232 (N_6232,In_3429,In_1637);
or U6233 (N_6233,In_4495,In_3251);
nor U6234 (N_6234,In_2422,In_4384);
and U6235 (N_6235,In_682,In_1902);
or U6236 (N_6236,In_3883,In_1836);
nor U6237 (N_6237,In_3989,In_4168);
nand U6238 (N_6238,In_3278,In_1538);
and U6239 (N_6239,In_4948,In_2937);
nand U6240 (N_6240,In_1927,In_4060);
or U6241 (N_6241,In_356,In_3910);
xor U6242 (N_6242,In_4248,In_4550);
or U6243 (N_6243,In_148,In_136);
nor U6244 (N_6244,In_524,In_453);
or U6245 (N_6245,In_3493,In_2779);
and U6246 (N_6246,In_3152,In_1310);
or U6247 (N_6247,In_4222,In_146);
and U6248 (N_6248,In_3285,In_1901);
xnor U6249 (N_6249,In_1923,In_3662);
and U6250 (N_6250,In_2046,In_3601);
xnor U6251 (N_6251,In_3309,In_1926);
xor U6252 (N_6252,In_1502,In_4585);
and U6253 (N_6253,In_2492,In_2138);
and U6254 (N_6254,In_4501,In_2696);
and U6255 (N_6255,In_4184,In_4332);
xnor U6256 (N_6256,In_3038,In_1123);
xor U6257 (N_6257,In_2035,In_3775);
nor U6258 (N_6258,In_155,In_2797);
xnor U6259 (N_6259,In_90,In_1781);
xor U6260 (N_6260,In_1922,In_3799);
xor U6261 (N_6261,In_3339,In_751);
or U6262 (N_6262,In_4823,In_1031);
or U6263 (N_6263,In_3209,In_2691);
and U6264 (N_6264,In_1415,In_1812);
or U6265 (N_6265,In_215,In_4767);
nor U6266 (N_6266,In_2120,In_3536);
nor U6267 (N_6267,In_3989,In_1905);
nand U6268 (N_6268,In_1243,In_1980);
nand U6269 (N_6269,In_1021,In_2369);
nand U6270 (N_6270,In_1809,In_84);
or U6271 (N_6271,In_4116,In_3499);
or U6272 (N_6272,In_613,In_1287);
xor U6273 (N_6273,In_599,In_1020);
or U6274 (N_6274,In_1044,In_2919);
and U6275 (N_6275,In_4049,In_3205);
xor U6276 (N_6276,In_3286,In_3215);
nand U6277 (N_6277,In_982,In_3846);
nor U6278 (N_6278,In_2202,In_3126);
nand U6279 (N_6279,In_4968,In_548);
and U6280 (N_6280,In_2925,In_1974);
or U6281 (N_6281,In_1709,In_2923);
nor U6282 (N_6282,In_3276,In_1163);
xnor U6283 (N_6283,In_1363,In_1362);
xor U6284 (N_6284,In_4155,In_4030);
xnor U6285 (N_6285,In_3890,In_4398);
xnor U6286 (N_6286,In_706,In_705);
nor U6287 (N_6287,In_3945,In_2041);
nand U6288 (N_6288,In_468,In_3799);
xnor U6289 (N_6289,In_2002,In_922);
and U6290 (N_6290,In_2492,In_3564);
nand U6291 (N_6291,In_885,In_1501);
nor U6292 (N_6292,In_2613,In_1904);
nor U6293 (N_6293,In_516,In_4745);
nor U6294 (N_6294,In_4784,In_2308);
nand U6295 (N_6295,In_1835,In_4842);
nor U6296 (N_6296,In_465,In_3762);
and U6297 (N_6297,In_4508,In_4380);
nor U6298 (N_6298,In_3567,In_133);
or U6299 (N_6299,In_858,In_3092);
or U6300 (N_6300,In_3110,In_1861);
and U6301 (N_6301,In_3353,In_4955);
or U6302 (N_6302,In_2866,In_2874);
nand U6303 (N_6303,In_4214,In_4538);
xor U6304 (N_6304,In_3550,In_494);
xnor U6305 (N_6305,In_3120,In_895);
nand U6306 (N_6306,In_2242,In_457);
and U6307 (N_6307,In_3230,In_2979);
nor U6308 (N_6308,In_3470,In_1620);
and U6309 (N_6309,In_3789,In_1146);
or U6310 (N_6310,In_2361,In_2858);
and U6311 (N_6311,In_4307,In_729);
and U6312 (N_6312,In_3414,In_4575);
and U6313 (N_6313,In_1154,In_1350);
nand U6314 (N_6314,In_4405,In_1692);
and U6315 (N_6315,In_142,In_3986);
or U6316 (N_6316,In_932,In_2415);
nor U6317 (N_6317,In_3290,In_2926);
xnor U6318 (N_6318,In_303,In_3013);
nor U6319 (N_6319,In_747,In_4610);
and U6320 (N_6320,In_2618,In_4535);
nand U6321 (N_6321,In_440,In_3457);
nor U6322 (N_6322,In_3784,In_699);
xor U6323 (N_6323,In_2252,In_221);
nand U6324 (N_6324,In_396,In_2620);
nor U6325 (N_6325,In_4165,In_4615);
nor U6326 (N_6326,In_3646,In_1870);
nand U6327 (N_6327,In_75,In_2437);
nand U6328 (N_6328,In_2877,In_4289);
xor U6329 (N_6329,In_914,In_1930);
nor U6330 (N_6330,In_1401,In_4529);
nand U6331 (N_6331,In_4884,In_61);
nand U6332 (N_6332,In_1028,In_4222);
nand U6333 (N_6333,In_4385,In_969);
xnor U6334 (N_6334,In_4256,In_412);
and U6335 (N_6335,In_2446,In_1848);
nand U6336 (N_6336,In_3953,In_1292);
nor U6337 (N_6337,In_1910,In_4781);
or U6338 (N_6338,In_3258,In_3673);
and U6339 (N_6339,In_1536,In_2757);
or U6340 (N_6340,In_2604,In_937);
or U6341 (N_6341,In_4251,In_318);
nand U6342 (N_6342,In_2721,In_351);
or U6343 (N_6343,In_2595,In_969);
xor U6344 (N_6344,In_4020,In_1865);
xor U6345 (N_6345,In_3216,In_772);
xor U6346 (N_6346,In_2529,In_4267);
xor U6347 (N_6347,In_4331,In_2791);
nand U6348 (N_6348,In_1394,In_4124);
or U6349 (N_6349,In_3900,In_1623);
nor U6350 (N_6350,In_3278,In_4621);
xnor U6351 (N_6351,In_4038,In_4441);
or U6352 (N_6352,In_3289,In_3125);
xor U6353 (N_6353,In_1266,In_2702);
or U6354 (N_6354,In_214,In_4499);
nand U6355 (N_6355,In_1004,In_562);
nand U6356 (N_6356,In_3450,In_2727);
xnor U6357 (N_6357,In_4758,In_2510);
and U6358 (N_6358,In_3767,In_3980);
and U6359 (N_6359,In_4041,In_3572);
nor U6360 (N_6360,In_3549,In_2399);
nor U6361 (N_6361,In_1962,In_430);
xor U6362 (N_6362,In_54,In_850);
nor U6363 (N_6363,In_2327,In_1278);
nor U6364 (N_6364,In_908,In_1114);
nand U6365 (N_6365,In_494,In_26);
and U6366 (N_6366,In_3301,In_3208);
xnor U6367 (N_6367,In_3943,In_829);
or U6368 (N_6368,In_4810,In_4128);
and U6369 (N_6369,In_3062,In_3010);
nor U6370 (N_6370,In_2236,In_4359);
and U6371 (N_6371,In_3812,In_4703);
and U6372 (N_6372,In_1703,In_2997);
xor U6373 (N_6373,In_1754,In_1025);
xor U6374 (N_6374,In_1430,In_326);
or U6375 (N_6375,In_1591,In_3514);
nand U6376 (N_6376,In_4995,In_2040);
or U6377 (N_6377,In_889,In_3574);
xnor U6378 (N_6378,In_4155,In_4218);
xor U6379 (N_6379,In_3337,In_2395);
and U6380 (N_6380,In_4292,In_2560);
or U6381 (N_6381,In_3562,In_2978);
or U6382 (N_6382,In_4524,In_4042);
nand U6383 (N_6383,In_1612,In_2172);
nand U6384 (N_6384,In_2356,In_1612);
nand U6385 (N_6385,In_1567,In_3075);
and U6386 (N_6386,In_2936,In_447);
or U6387 (N_6387,In_298,In_3761);
nand U6388 (N_6388,In_2145,In_2532);
and U6389 (N_6389,In_3370,In_2852);
nor U6390 (N_6390,In_3054,In_1571);
nand U6391 (N_6391,In_4157,In_460);
xor U6392 (N_6392,In_4009,In_329);
xnor U6393 (N_6393,In_617,In_3694);
and U6394 (N_6394,In_2510,In_2546);
xnor U6395 (N_6395,In_1600,In_3279);
or U6396 (N_6396,In_1820,In_2671);
xnor U6397 (N_6397,In_3352,In_774);
xor U6398 (N_6398,In_1400,In_1740);
nand U6399 (N_6399,In_2770,In_1934);
nor U6400 (N_6400,In_3990,In_3);
xor U6401 (N_6401,In_1029,In_4048);
or U6402 (N_6402,In_1367,In_4542);
or U6403 (N_6403,In_2643,In_2613);
and U6404 (N_6404,In_452,In_764);
and U6405 (N_6405,In_2133,In_1540);
nor U6406 (N_6406,In_2668,In_1712);
xor U6407 (N_6407,In_1729,In_4301);
nor U6408 (N_6408,In_2822,In_2869);
or U6409 (N_6409,In_1189,In_267);
nand U6410 (N_6410,In_821,In_551);
xnor U6411 (N_6411,In_17,In_2081);
nand U6412 (N_6412,In_285,In_3531);
and U6413 (N_6413,In_4273,In_1587);
or U6414 (N_6414,In_3766,In_4316);
xor U6415 (N_6415,In_4699,In_1543);
nor U6416 (N_6416,In_2757,In_4003);
or U6417 (N_6417,In_393,In_3652);
nand U6418 (N_6418,In_2876,In_109);
nor U6419 (N_6419,In_4924,In_1198);
or U6420 (N_6420,In_2920,In_3224);
or U6421 (N_6421,In_1500,In_521);
or U6422 (N_6422,In_2351,In_2371);
or U6423 (N_6423,In_3421,In_1583);
xnor U6424 (N_6424,In_3807,In_4888);
nand U6425 (N_6425,In_1783,In_2886);
nand U6426 (N_6426,In_4547,In_1265);
xnor U6427 (N_6427,In_878,In_4353);
and U6428 (N_6428,In_3812,In_552);
nor U6429 (N_6429,In_4589,In_1392);
and U6430 (N_6430,In_1162,In_9);
nand U6431 (N_6431,In_2335,In_1613);
xnor U6432 (N_6432,In_4273,In_744);
and U6433 (N_6433,In_2950,In_1873);
nand U6434 (N_6434,In_2606,In_544);
or U6435 (N_6435,In_2698,In_1717);
nor U6436 (N_6436,In_462,In_4589);
nand U6437 (N_6437,In_3827,In_545);
and U6438 (N_6438,In_964,In_3585);
nor U6439 (N_6439,In_1712,In_860);
and U6440 (N_6440,In_3992,In_2656);
xor U6441 (N_6441,In_4233,In_1403);
xnor U6442 (N_6442,In_1159,In_1315);
xor U6443 (N_6443,In_4216,In_2322);
xor U6444 (N_6444,In_1252,In_2524);
xnor U6445 (N_6445,In_4493,In_4100);
nand U6446 (N_6446,In_2065,In_1973);
nor U6447 (N_6447,In_2630,In_4241);
and U6448 (N_6448,In_4948,In_4027);
or U6449 (N_6449,In_1624,In_3636);
or U6450 (N_6450,In_2537,In_1395);
nor U6451 (N_6451,In_2026,In_2132);
xnor U6452 (N_6452,In_4488,In_1227);
and U6453 (N_6453,In_4669,In_3638);
or U6454 (N_6454,In_4870,In_2615);
xnor U6455 (N_6455,In_3530,In_2679);
or U6456 (N_6456,In_4872,In_3077);
and U6457 (N_6457,In_310,In_3184);
and U6458 (N_6458,In_4225,In_2787);
nor U6459 (N_6459,In_33,In_4533);
xnor U6460 (N_6460,In_4753,In_3186);
xnor U6461 (N_6461,In_2943,In_4644);
xor U6462 (N_6462,In_1907,In_3896);
and U6463 (N_6463,In_984,In_749);
or U6464 (N_6464,In_328,In_1772);
and U6465 (N_6465,In_871,In_2251);
nand U6466 (N_6466,In_1523,In_2155);
or U6467 (N_6467,In_371,In_3297);
xor U6468 (N_6468,In_4839,In_4394);
nor U6469 (N_6469,In_578,In_312);
nor U6470 (N_6470,In_2768,In_993);
xnor U6471 (N_6471,In_2037,In_1548);
nand U6472 (N_6472,In_1893,In_2804);
nor U6473 (N_6473,In_2396,In_511);
nor U6474 (N_6474,In_2188,In_4691);
and U6475 (N_6475,In_903,In_3798);
and U6476 (N_6476,In_833,In_277);
nand U6477 (N_6477,In_2678,In_2151);
and U6478 (N_6478,In_4117,In_2584);
and U6479 (N_6479,In_1377,In_1569);
nand U6480 (N_6480,In_791,In_2221);
or U6481 (N_6481,In_267,In_1982);
or U6482 (N_6482,In_3267,In_4834);
nor U6483 (N_6483,In_3366,In_3012);
xor U6484 (N_6484,In_4850,In_75);
xnor U6485 (N_6485,In_4850,In_155);
and U6486 (N_6486,In_3234,In_4553);
or U6487 (N_6487,In_680,In_4413);
or U6488 (N_6488,In_2732,In_938);
nand U6489 (N_6489,In_2152,In_2262);
xor U6490 (N_6490,In_1319,In_3236);
and U6491 (N_6491,In_2668,In_3949);
nor U6492 (N_6492,In_2218,In_204);
nor U6493 (N_6493,In_2931,In_2552);
and U6494 (N_6494,In_3695,In_4680);
nor U6495 (N_6495,In_2614,In_1410);
nand U6496 (N_6496,In_3950,In_3348);
nand U6497 (N_6497,In_4801,In_253);
nor U6498 (N_6498,In_4588,In_4943);
nor U6499 (N_6499,In_2372,In_3807);
xnor U6500 (N_6500,In_4143,In_957);
xnor U6501 (N_6501,In_779,In_2219);
or U6502 (N_6502,In_2128,In_330);
nor U6503 (N_6503,In_1635,In_1617);
nor U6504 (N_6504,In_1484,In_1971);
xnor U6505 (N_6505,In_115,In_3785);
xor U6506 (N_6506,In_3168,In_3293);
xnor U6507 (N_6507,In_1964,In_4655);
nand U6508 (N_6508,In_3233,In_1336);
xor U6509 (N_6509,In_2943,In_2744);
nand U6510 (N_6510,In_2315,In_289);
and U6511 (N_6511,In_4480,In_2061);
xnor U6512 (N_6512,In_1345,In_1913);
xnor U6513 (N_6513,In_2172,In_2640);
nand U6514 (N_6514,In_3172,In_4552);
or U6515 (N_6515,In_3168,In_1508);
nand U6516 (N_6516,In_4590,In_2317);
nand U6517 (N_6517,In_1665,In_3919);
nor U6518 (N_6518,In_4371,In_1616);
and U6519 (N_6519,In_2345,In_591);
or U6520 (N_6520,In_1264,In_3363);
and U6521 (N_6521,In_3443,In_741);
and U6522 (N_6522,In_3824,In_3960);
nor U6523 (N_6523,In_3523,In_3324);
xnor U6524 (N_6524,In_3969,In_658);
and U6525 (N_6525,In_2313,In_248);
xnor U6526 (N_6526,In_4498,In_747);
and U6527 (N_6527,In_3149,In_1378);
and U6528 (N_6528,In_3403,In_3469);
xor U6529 (N_6529,In_3288,In_564);
nor U6530 (N_6530,In_30,In_263);
xnor U6531 (N_6531,In_1798,In_3919);
and U6532 (N_6532,In_731,In_4067);
nand U6533 (N_6533,In_162,In_4274);
or U6534 (N_6534,In_2455,In_2720);
nor U6535 (N_6535,In_1881,In_86);
and U6536 (N_6536,In_53,In_3567);
xnor U6537 (N_6537,In_2850,In_69);
nor U6538 (N_6538,In_3406,In_4661);
xor U6539 (N_6539,In_2452,In_3314);
nand U6540 (N_6540,In_2205,In_1663);
nor U6541 (N_6541,In_4627,In_2355);
nor U6542 (N_6542,In_3327,In_148);
or U6543 (N_6543,In_4732,In_2279);
nand U6544 (N_6544,In_1991,In_1672);
nand U6545 (N_6545,In_4274,In_3817);
nand U6546 (N_6546,In_1888,In_4003);
and U6547 (N_6547,In_3986,In_520);
and U6548 (N_6548,In_1887,In_4839);
xnor U6549 (N_6549,In_4586,In_637);
nor U6550 (N_6550,In_2567,In_4984);
xnor U6551 (N_6551,In_4843,In_192);
or U6552 (N_6552,In_1000,In_4562);
nor U6553 (N_6553,In_3402,In_3566);
xnor U6554 (N_6554,In_3588,In_2355);
and U6555 (N_6555,In_1589,In_793);
and U6556 (N_6556,In_594,In_3712);
and U6557 (N_6557,In_464,In_1496);
xor U6558 (N_6558,In_1492,In_4730);
xor U6559 (N_6559,In_50,In_2938);
or U6560 (N_6560,In_140,In_1918);
nor U6561 (N_6561,In_4199,In_1507);
xnor U6562 (N_6562,In_3595,In_1326);
xnor U6563 (N_6563,In_1360,In_1753);
and U6564 (N_6564,In_4576,In_4255);
or U6565 (N_6565,In_4464,In_3731);
nor U6566 (N_6566,In_3166,In_320);
or U6567 (N_6567,In_3751,In_1649);
and U6568 (N_6568,In_3327,In_491);
nor U6569 (N_6569,In_4584,In_3589);
xor U6570 (N_6570,In_2729,In_54);
xnor U6571 (N_6571,In_3896,In_370);
and U6572 (N_6572,In_3106,In_1651);
nor U6573 (N_6573,In_4190,In_4505);
nor U6574 (N_6574,In_2417,In_385);
nand U6575 (N_6575,In_1311,In_3245);
or U6576 (N_6576,In_1402,In_212);
or U6577 (N_6577,In_1380,In_3724);
nand U6578 (N_6578,In_1028,In_4756);
or U6579 (N_6579,In_4782,In_778);
nor U6580 (N_6580,In_4366,In_4736);
nor U6581 (N_6581,In_493,In_764);
and U6582 (N_6582,In_1279,In_1627);
or U6583 (N_6583,In_393,In_1883);
nand U6584 (N_6584,In_4709,In_3564);
nor U6585 (N_6585,In_3611,In_2436);
nand U6586 (N_6586,In_4162,In_447);
and U6587 (N_6587,In_416,In_2888);
or U6588 (N_6588,In_1111,In_3583);
and U6589 (N_6589,In_597,In_216);
xor U6590 (N_6590,In_4015,In_3137);
and U6591 (N_6591,In_2019,In_479);
xnor U6592 (N_6592,In_1785,In_1992);
nor U6593 (N_6593,In_2835,In_2269);
nand U6594 (N_6594,In_2250,In_267);
nand U6595 (N_6595,In_573,In_1657);
and U6596 (N_6596,In_535,In_1454);
nor U6597 (N_6597,In_4728,In_1384);
or U6598 (N_6598,In_1414,In_1725);
and U6599 (N_6599,In_3153,In_1365);
nor U6600 (N_6600,In_333,In_3067);
xor U6601 (N_6601,In_8,In_4675);
and U6602 (N_6602,In_1907,In_1339);
nor U6603 (N_6603,In_3290,In_4169);
or U6604 (N_6604,In_1025,In_3620);
nand U6605 (N_6605,In_4534,In_2347);
nand U6606 (N_6606,In_4038,In_1819);
nand U6607 (N_6607,In_2098,In_3905);
and U6608 (N_6608,In_2895,In_1557);
nor U6609 (N_6609,In_3045,In_848);
and U6610 (N_6610,In_2388,In_3630);
nand U6611 (N_6611,In_3779,In_4288);
and U6612 (N_6612,In_4204,In_173);
and U6613 (N_6613,In_518,In_3559);
or U6614 (N_6614,In_1068,In_4359);
nand U6615 (N_6615,In_3658,In_1431);
or U6616 (N_6616,In_4677,In_1202);
nor U6617 (N_6617,In_3537,In_4192);
nand U6618 (N_6618,In_3687,In_4465);
or U6619 (N_6619,In_1347,In_4451);
or U6620 (N_6620,In_2253,In_567);
and U6621 (N_6621,In_1666,In_2955);
nor U6622 (N_6622,In_980,In_18);
nand U6623 (N_6623,In_1589,In_4660);
or U6624 (N_6624,In_3304,In_4833);
nor U6625 (N_6625,In_3040,In_3971);
and U6626 (N_6626,In_4784,In_1013);
xnor U6627 (N_6627,In_2550,In_1167);
xnor U6628 (N_6628,In_515,In_642);
xor U6629 (N_6629,In_4342,In_4606);
nor U6630 (N_6630,In_2917,In_150);
xor U6631 (N_6631,In_3513,In_1482);
xnor U6632 (N_6632,In_1225,In_550);
or U6633 (N_6633,In_4775,In_4678);
or U6634 (N_6634,In_3096,In_3277);
nor U6635 (N_6635,In_3650,In_2811);
xnor U6636 (N_6636,In_4493,In_1114);
or U6637 (N_6637,In_2717,In_4750);
and U6638 (N_6638,In_848,In_2582);
nor U6639 (N_6639,In_1256,In_311);
nor U6640 (N_6640,In_4571,In_2827);
xor U6641 (N_6641,In_2748,In_4534);
nand U6642 (N_6642,In_4373,In_2225);
nor U6643 (N_6643,In_2422,In_3432);
or U6644 (N_6644,In_1488,In_3133);
nor U6645 (N_6645,In_2261,In_3074);
and U6646 (N_6646,In_4187,In_2339);
nor U6647 (N_6647,In_3814,In_3404);
xor U6648 (N_6648,In_3526,In_718);
and U6649 (N_6649,In_1167,In_199);
nor U6650 (N_6650,In_3270,In_8);
or U6651 (N_6651,In_697,In_2078);
xor U6652 (N_6652,In_541,In_631);
nand U6653 (N_6653,In_2956,In_719);
and U6654 (N_6654,In_4453,In_806);
nor U6655 (N_6655,In_307,In_55);
xor U6656 (N_6656,In_1972,In_1408);
and U6657 (N_6657,In_4291,In_4231);
or U6658 (N_6658,In_221,In_3476);
or U6659 (N_6659,In_1561,In_3877);
nand U6660 (N_6660,In_3116,In_3331);
nor U6661 (N_6661,In_2452,In_3277);
and U6662 (N_6662,In_2006,In_1154);
nor U6663 (N_6663,In_2366,In_2338);
xor U6664 (N_6664,In_2781,In_2181);
xnor U6665 (N_6665,In_4867,In_2176);
nand U6666 (N_6666,In_2031,In_286);
and U6667 (N_6667,In_1533,In_2342);
nor U6668 (N_6668,In_3584,In_2072);
nand U6669 (N_6669,In_4541,In_1930);
or U6670 (N_6670,In_3852,In_605);
and U6671 (N_6671,In_1124,In_355);
and U6672 (N_6672,In_2002,In_3700);
nand U6673 (N_6673,In_4961,In_4838);
or U6674 (N_6674,In_2455,In_3930);
nand U6675 (N_6675,In_1822,In_3005);
nor U6676 (N_6676,In_2133,In_2032);
or U6677 (N_6677,In_2986,In_4903);
and U6678 (N_6678,In_4149,In_990);
or U6679 (N_6679,In_883,In_2330);
or U6680 (N_6680,In_3582,In_4267);
and U6681 (N_6681,In_333,In_545);
nand U6682 (N_6682,In_1051,In_1694);
nand U6683 (N_6683,In_4762,In_3339);
xor U6684 (N_6684,In_3710,In_3063);
and U6685 (N_6685,In_701,In_1645);
and U6686 (N_6686,In_1552,In_4453);
nor U6687 (N_6687,In_1111,In_1258);
nor U6688 (N_6688,In_57,In_3051);
nand U6689 (N_6689,In_3906,In_3335);
nand U6690 (N_6690,In_4809,In_4135);
nand U6691 (N_6691,In_1108,In_1435);
xor U6692 (N_6692,In_1142,In_4095);
nand U6693 (N_6693,In_308,In_2505);
xor U6694 (N_6694,In_1607,In_2138);
or U6695 (N_6695,In_1685,In_1303);
nor U6696 (N_6696,In_822,In_1813);
and U6697 (N_6697,In_234,In_2506);
or U6698 (N_6698,In_1578,In_654);
nor U6699 (N_6699,In_4335,In_1507);
and U6700 (N_6700,In_170,In_32);
nand U6701 (N_6701,In_3255,In_2434);
or U6702 (N_6702,In_3353,In_3208);
and U6703 (N_6703,In_2738,In_3358);
nor U6704 (N_6704,In_2271,In_1953);
and U6705 (N_6705,In_3863,In_3367);
nor U6706 (N_6706,In_326,In_2835);
xnor U6707 (N_6707,In_2202,In_100);
and U6708 (N_6708,In_527,In_2719);
or U6709 (N_6709,In_357,In_761);
and U6710 (N_6710,In_2423,In_348);
nor U6711 (N_6711,In_143,In_4215);
and U6712 (N_6712,In_1488,In_3605);
nand U6713 (N_6713,In_4880,In_1207);
and U6714 (N_6714,In_2110,In_2549);
nor U6715 (N_6715,In_3637,In_3753);
and U6716 (N_6716,In_4579,In_2107);
nor U6717 (N_6717,In_3720,In_722);
xnor U6718 (N_6718,In_1966,In_1395);
and U6719 (N_6719,In_124,In_4731);
nand U6720 (N_6720,In_1957,In_2087);
or U6721 (N_6721,In_1431,In_1304);
nor U6722 (N_6722,In_853,In_3208);
nor U6723 (N_6723,In_770,In_2501);
or U6724 (N_6724,In_4242,In_3724);
xnor U6725 (N_6725,In_3801,In_3257);
nor U6726 (N_6726,In_3141,In_622);
or U6727 (N_6727,In_1288,In_4048);
xnor U6728 (N_6728,In_2421,In_4839);
and U6729 (N_6729,In_1028,In_134);
nor U6730 (N_6730,In_2695,In_3754);
and U6731 (N_6731,In_621,In_1646);
nor U6732 (N_6732,In_3784,In_4517);
nand U6733 (N_6733,In_4289,In_1393);
xnor U6734 (N_6734,In_2839,In_4981);
nor U6735 (N_6735,In_2991,In_3289);
nand U6736 (N_6736,In_37,In_3371);
nor U6737 (N_6737,In_3429,In_4682);
nor U6738 (N_6738,In_3502,In_4453);
nand U6739 (N_6739,In_422,In_3428);
and U6740 (N_6740,In_1997,In_2682);
or U6741 (N_6741,In_2114,In_10);
nor U6742 (N_6742,In_1491,In_2063);
nand U6743 (N_6743,In_148,In_1571);
nor U6744 (N_6744,In_4832,In_2581);
or U6745 (N_6745,In_4263,In_2435);
or U6746 (N_6746,In_3070,In_167);
and U6747 (N_6747,In_627,In_1247);
nand U6748 (N_6748,In_4084,In_1414);
nor U6749 (N_6749,In_4446,In_4456);
xnor U6750 (N_6750,In_1211,In_1376);
xor U6751 (N_6751,In_1424,In_1286);
nand U6752 (N_6752,In_1531,In_1090);
xor U6753 (N_6753,In_3594,In_4706);
nand U6754 (N_6754,In_4461,In_1556);
or U6755 (N_6755,In_2220,In_3601);
nand U6756 (N_6756,In_4600,In_531);
xnor U6757 (N_6757,In_484,In_1276);
or U6758 (N_6758,In_943,In_284);
xor U6759 (N_6759,In_2695,In_1046);
and U6760 (N_6760,In_1023,In_2922);
nor U6761 (N_6761,In_1836,In_2061);
and U6762 (N_6762,In_137,In_1363);
or U6763 (N_6763,In_3875,In_4577);
nand U6764 (N_6764,In_2744,In_4621);
nor U6765 (N_6765,In_3471,In_421);
xor U6766 (N_6766,In_1114,In_3189);
xor U6767 (N_6767,In_3042,In_3571);
and U6768 (N_6768,In_3616,In_4081);
nor U6769 (N_6769,In_338,In_3061);
and U6770 (N_6770,In_1411,In_1592);
or U6771 (N_6771,In_3592,In_1736);
nor U6772 (N_6772,In_310,In_4505);
or U6773 (N_6773,In_3068,In_4932);
or U6774 (N_6774,In_845,In_4061);
xnor U6775 (N_6775,In_4172,In_1855);
nand U6776 (N_6776,In_206,In_54);
xor U6777 (N_6777,In_588,In_29);
nand U6778 (N_6778,In_4245,In_3147);
and U6779 (N_6779,In_344,In_4577);
xor U6780 (N_6780,In_385,In_2814);
and U6781 (N_6781,In_4458,In_1854);
nand U6782 (N_6782,In_2371,In_1986);
nand U6783 (N_6783,In_138,In_3061);
nor U6784 (N_6784,In_2266,In_1869);
or U6785 (N_6785,In_1821,In_3423);
or U6786 (N_6786,In_605,In_1624);
nor U6787 (N_6787,In_3150,In_4309);
xnor U6788 (N_6788,In_94,In_3970);
nor U6789 (N_6789,In_1791,In_3410);
or U6790 (N_6790,In_4734,In_4528);
and U6791 (N_6791,In_4501,In_1655);
xor U6792 (N_6792,In_2074,In_599);
nand U6793 (N_6793,In_3962,In_2168);
and U6794 (N_6794,In_3446,In_4708);
nor U6795 (N_6795,In_4605,In_3569);
and U6796 (N_6796,In_654,In_2035);
nor U6797 (N_6797,In_1404,In_2051);
nand U6798 (N_6798,In_3561,In_228);
or U6799 (N_6799,In_4751,In_2837);
or U6800 (N_6800,In_2759,In_2881);
and U6801 (N_6801,In_4993,In_868);
nand U6802 (N_6802,In_3296,In_1379);
nor U6803 (N_6803,In_4749,In_1840);
xor U6804 (N_6804,In_3333,In_351);
nand U6805 (N_6805,In_4660,In_3515);
nor U6806 (N_6806,In_4726,In_768);
or U6807 (N_6807,In_4201,In_3415);
xnor U6808 (N_6808,In_4551,In_4419);
xor U6809 (N_6809,In_3495,In_2364);
and U6810 (N_6810,In_3441,In_1767);
nor U6811 (N_6811,In_4570,In_3487);
xnor U6812 (N_6812,In_3547,In_892);
nor U6813 (N_6813,In_1273,In_2146);
nand U6814 (N_6814,In_3087,In_3074);
or U6815 (N_6815,In_978,In_990);
nand U6816 (N_6816,In_1332,In_2546);
nor U6817 (N_6817,In_4277,In_1734);
nor U6818 (N_6818,In_2030,In_2902);
nand U6819 (N_6819,In_340,In_3747);
and U6820 (N_6820,In_4717,In_3336);
and U6821 (N_6821,In_4311,In_1826);
or U6822 (N_6822,In_489,In_3280);
xnor U6823 (N_6823,In_2118,In_2928);
or U6824 (N_6824,In_4847,In_2595);
nor U6825 (N_6825,In_4384,In_1393);
and U6826 (N_6826,In_2348,In_3556);
nor U6827 (N_6827,In_2035,In_2254);
nand U6828 (N_6828,In_163,In_599);
nand U6829 (N_6829,In_2399,In_4296);
or U6830 (N_6830,In_1320,In_3970);
xnor U6831 (N_6831,In_1971,In_245);
and U6832 (N_6832,In_129,In_4383);
nor U6833 (N_6833,In_2818,In_1330);
xor U6834 (N_6834,In_342,In_1754);
or U6835 (N_6835,In_109,In_1720);
and U6836 (N_6836,In_1088,In_3063);
nor U6837 (N_6837,In_904,In_1445);
nor U6838 (N_6838,In_746,In_3266);
and U6839 (N_6839,In_864,In_3996);
nand U6840 (N_6840,In_1198,In_3358);
nand U6841 (N_6841,In_3185,In_1783);
or U6842 (N_6842,In_4424,In_1951);
xnor U6843 (N_6843,In_4759,In_2976);
or U6844 (N_6844,In_3013,In_1868);
nor U6845 (N_6845,In_2667,In_72);
xor U6846 (N_6846,In_3197,In_3896);
or U6847 (N_6847,In_2173,In_2517);
nand U6848 (N_6848,In_2248,In_760);
nand U6849 (N_6849,In_4716,In_1423);
nor U6850 (N_6850,In_4076,In_373);
nand U6851 (N_6851,In_1605,In_1735);
or U6852 (N_6852,In_466,In_2708);
nand U6853 (N_6853,In_3840,In_4368);
nor U6854 (N_6854,In_1047,In_3133);
or U6855 (N_6855,In_2923,In_4222);
xnor U6856 (N_6856,In_1608,In_1447);
and U6857 (N_6857,In_740,In_3814);
or U6858 (N_6858,In_672,In_4685);
nor U6859 (N_6859,In_1357,In_4580);
or U6860 (N_6860,In_2683,In_3176);
nor U6861 (N_6861,In_518,In_1980);
and U6862 (N_6862,In_4150,In_680);
and U6863 (N_6863,In_1006,In_2769);
nor U6864 (N_6864,In_3351,In_1177);
or U6865 (N_6865,In_1587,In_3802);
or U6866 (N_6866,In_1572,In_9);
nand U6867 (N_6867,In_1129,In_199);
or U6868 (N_6868,In_4300,In_2492);
nand U6869 (N_6869,In_2127,In_3136);
nand U6870 (N_6870,In_3342,In_3076);
nor U6871 (N_6871,In_3952,In_4636);
and U6872 (N_6872,In_2288,In_1683);
nand U6873 (N_6873,In_714,In_3377);
xnor U6874 (N_6874,In_1544,In_2838);
and U6875 (N_6875,In_3985,In_1451);
xor U6876 (N_6876,In_97,In_4342);
xor U6877 (N_6877,In_549,In_4279);
xor U6878 (N_6878,In_1281,In_2905);
or U6879 (N_6879,In_915,In_1594);
nand U6880 (N_6880,In_825,In_3767);
xnor U6881 (N_6881,In_1735,In_1496);
or U6882 (N_6882,In_3688,In_4797);
xnor U6883 (N_6883,In_3177,In_2953);
and U6884 (N_6884,In_4328,In_1656);
and U6885 (N_6885,In_1220,In_346);
nand U6886 (N_6886,In_2899,In_1618);
and U6887 (N_6887,In_1621,In_1351);
or U6888 (N_6888,In_4428,In_523);
nor U6889 (N_6889,In_1570,In_1290);
xor U6890 (N_6890,In_1024,In_1433);
and U6891 (N_6891,In_2787,In_3615);
or U6892 (N_6892,In_3706,In_2685);
nor U6893 (N_6893,In_2233,In_3395);
nand U6894 (N_6894,In_1544,In_3210);
nor U6895 (N_6895,In_1676,In_4732);
xor U6896 (N_6896,In_1268,In_2074);
xnor U6897 (N_6897,In_2198,In_614);
nor U6898 (N_6898,In_1522,In_4218);
and U6899 (N_6899,In_3219,In_553);
nand U6900 (N_6900,In_455,In_2737);
or U6901 (N_6901,In_4280,In_4636);
nor U6902 (N_6902,In_2074,In_4754);
xnor U6903 (N_6903,In_2291,In_4707);
and U6904 (N_6904,In_2811,In_4605);
and U6905 (N_6905,In_1529,In_1721);
xor U6906 (N_6906,In_3230,In_2448);
or U6907 (N_6907,In_3413,In_1900);
nand U6908 (N_6908,In_3173,In_3744);
and U6909 (N_6909,In_315,In_2623);
or U6910 (N_6910,In_2627,In_2577);
and U6911 (N_6911,In_2338,In_1962);
xnor U6912 (N_6912,In_385,In_4652);
and U6913 (N_6913,In_4878,In_1134);
nor U6914 (N_6914,In_718,In_2159);
nand U6915 (N_6915,In_472,In_2507);
or U6916 (N_6916,In_3259,In_4008);
nand U6917 (N_6917,In_2419,In_2386);
and U6918 (N_6918,In_605,In_2917);
nor U6919 (N_6919,In_3500,In_646);
nor U6920 (N_6920,In_3265,In_4839);
and U6921 (N_6921,In_2624,In_1840);
or U6922 (N_6922,In_2038,In_1625);
or U6923 (N_6923,In_536,In_3631);
nor U6924 (N_6924,In_507,In_852);
nand U6925 (N_6925,In_3216,In_1266);
xor U6926 (N_6926,In_1398,In_1035);
nor U6927 (N_6927,In_2152,In_1270);
xor U6928 (N_6928,In_2424,In_2568);
nand U6929 (N_6929,In_3832,In_20);
or U6930 (N_6930,In_1831,In_4764);
xor U6931 (N_6931,In_986,In_4858);
or U6932 (N_6932,In_2348,In_2896);
xnor U6933 (N_6933,In_1224,In_3651);
and U6934 (N_6934,In_3044,In_3973);
and U6935 (N_6935,In_1095,In_4786);
and U6936 (N_6936,In_1091,In_2172);
xor U6937 (N_6937,In_2894,In_3832);
or U6938 (N_6938,In_530,In_4246);
and U6939 (N_6939,In_428,In_1274);
nand U6940 (N_6940,In_752,In_3720);
nand U6941 (N_6941,In_195,In_3430);
and U6942 (N_6942,In_71,In_1981);
and U6943 (N_6943,In_1594,In_2278);
or U6944 (N_6944,In_100,In_2737);
nor U6945 (N_6945,In_3529,In_2944);
nand U6946 (N_6946,In_3357,In_4583);
or U6947 (N_6947,In_3516,In_4162);
or U6948 (N_6948,In_1622,In_4055);
nor U6949 (N_6949,In_2606,In_3555);
xnor U6950 (N_6950,In_4921,In_3580);
nor U6951 (N_6951,In_749,In_2837);
and U6952 (N_6952,In_726,In_3187);
xor U6953 (N_6953,In_1790,In_2931);
nor U6954 (N_6954,In_4472,In_352);
or U6955 (N_6955,In_2938,In_4953);
nor U6956 (N_6956,In_1906,In_744);
xnor U6957 (N_6957,In_624,In_479);
xnor U6958 (N_6958,In_4802,In_376);
nor U6959 (N_6959,In_602,In_1493);
or U6960 (N_6960,In_4822,In_381);
nand U6961 (N_6961,In_4221,In_4632);
or U6962 (N_6962,In_3376,In_3195);
nand U6963 (N_6963,In_4666,In_1545);
xor U6964 (N_6964,In_3039,In_2112);
xor U6965 (N_6965,In_2736,In_3387);
nor U6966 (N_6966,In_1035,In_2581);
xnor U6967 (N_6967,In_3729,In_3556);
xnor U6968 (N_6968,In_3569,In_1620);
or U6969 (N_6969,In_1623,In_135);
xnor U6970 (N_6970,In_2003,In_1544);
xor U6971 (N_6971,In_2076,In_179);
or U6972 (N_6972,In_2224,In_3307);
and U6973 (N_6973,In_3707,In_4578);
or U6974 (N_6974,In_232,In_774);
nor U6975 (N_6975,In_2952,In_1189);
or U6976 (N_6976,In_3997,In_126);
xor U6977 (N_6977,In_1863,In_3818);
nand U6978 (N_6978,In_2058,In_881);
and U6979 (N_6979,In_54,In_889);
xor U6980 (N_6980,In_2907,In_1929);
nor U6981 (N_6981,In_2677,In_2268);
xor U6982 (N_6982,In_3466,In_2739);
xor U6983 (N_6983,In_2154,In_1248);
and U6984 (N_6984,In_2354,In_1260);
or U6985 (N_6985,In_3906,In_3343);
or U6986 (N_6986,In_382,In_2838);
nand U6987 (N_6987,In_4514,In_2744);
nor U6988 (N_6988,In_2856,In_4468);
nor U6989 (N_6989,In_4905,In_3235);
xnor U6990 (N_6990,In_4072,In_1069);
xnor U6991 (N_6991,In_611,In_4300);
nand U6992 (N_6992,In_1385,In_768);
and U6993 (N_6993,In_3112,In_2287);
nor U6994 (N_6994,In_2751,In_3494);
nand U6995 (N_6995,In_4648,In_1256);
xor U6996 (N_6996,In_1177,In_452);
nor U6997 (N_6997,In_140,In_3067);
and U6998 (N_6998,In_4609,In_2581);
nor U6999 (N_6999,In_3829,In_3203);
nor U7000 (N_7000,In_2278,In_4322);
nand U7001 (N_7001,In_2363,In_1128);
xor U7002 (N_7002,In_4856,In_3119);
nand U7003 (N_7003,In_507,In_3130);
xor U7004 (N_7004,In_1112,In_4670);
and U7005 (N_7005,In_4596,In_4781);
nor U7006 (N_7006,In_2195,In_53);
nand U7007 (N_7007,In_3855,In_2104);
nand U7008 (N_7008,In_4838,In_3942);
and U7009 (N_7009,In_900,In_4424);
nor U7010 (N_7010,In_4719,In_3797);
and U7011 (N_7011,In_2103,In_1749);
xor U7012 (N_7012,In_1766,In_3379);
nand U7013 (N_7013,In_900,In_3190);
nor U7014 (N_7014,In_1368,In_4234);
or U7015 (N_7015,In_4621,In_2369);
or U7016 (N_7016,In_2237,In_2438);
xnor U7017 (N_7017,In_517,In_2791);
xnor U7018 (N_7018,In_88,In_1318);
nor U7019 (N_7019,In_4552,In_3149);
nand U7020 (N_7020,In_4901,In_3303);
nor U7021 (N_7021,In_1619,In_2937);
and U7022 (N_7022,In_4424,In_4024);
and U7023 (N_7023,In_177,In_2489);
or U7024 (N_7024,In_1304,In_1222);
or U7025 (N_7025,In_2345,In_1593);
nor U7026 (N_7026,In_1037,In_2124);
xor U7027 (N_7027,In_2415,In_1418);
nor U7028 (N_7028,In_4049,In_1516);
xnor U7029 (N_7029,In_927,In_13);
and U7030 (N_7030,In_1151,In_741);
nor U7031 (N_7031,In_2,In_3897);
and U7032 (N_7032,In_458,In_3147);
nand U7033 (N_7033,In_3433,In_2727);
nand U7034 (N_7034,In_2706,In_3007);
nand U7035 (N_7035,In_3380,In_1236);
nand U7036 (N_7036,In_2221,In_524);
or U7037 (N_7037,In_2446,In_447);
and U7038 (N_7038,In_414,In_4972);
or U7039 (N_7039,In_1814,In_3113);
nor U7040 (N_7040,In_1574,In_488);
or U7041 (N_7041,In_799,In_2344);
and U7042 (N_7042,In_2919,In_1264);
or U7043 (N_7043,In_4195,In_4689);
nand U7044 (N_7044,In_4653,In_1481);
or U7045 (N_7045,In_4465,In_1183);
nor U7046 (N_7046,In_2416,In_1018);
xnor U7047 (N_7047,In_1857,In_651);
xor U7048 (N_7048,In_472,In_2625);
or U7049 (N_7049,In_2929,In_4500);
and U7050 (N_7050,In_1641,In_2730);
nand U7051 (N_7051,In_2857,In_2741);
nor U7052 (N_7052,In_4086,In_1972);
xnor U7053 (N_7053,In_2875,In_568);
nand U7054 (N_7054,In_3726,In_1756);
xor U7055 (N_7055,In_4591,In_1936);
xnor U7056 (N_7056,In_3410,In_1169);
xor U7057 (N_7057,In_4762,In_233);
nor U7058 (N_7058,In_2141,In_2630);
xnor U7059 (N_7059,In_3540,In_471);
nor U7060 (N_7060,In_2356,In_166);
nor U7061 (N_7061,In_4969,In_344);
or U7062 (N_7062,In_2428,In_782);
nor U7063 (N_7063,In_4927,In_32);
xnor U7064 (N_7064,In_3070,In_2314);
and U7065 (N_7065,In_440,In_630);
nand U7066 (N_7066,In_2920,In_837);
xor U7067 (N_7067,In_4517,In_4522);
nor U7068 (N_7068,In_1668,In_3757);
and U7069 (N_7069,In_196,In_4115);
xnor U7070 (N_7070,In_4421,In_333);
or U7071 (N_7071,In_3783,In_30);
xnor U7072 (N_7072,In_1871,In_892);
xor U7073 (N_7073,In_2388,In_2236);
nor U7074 (N_7074,In_942,In_946);
or U7075 (N_7075,In_828,In_3546);
and U7076 (N_7076,In_3707,In_128);
and U7077 (N_7077,In_4079,In_2201);
xor U7078 (N_7078,In_3717,In_4993);
or U7079 (N_7079,In_2497,In_1271);
and U7080 (N_7080,In_148,In_3710);
nand U7081 (N_7081,In_4105,In_814);
nor U7082 (N_7082,In_3249,In_3222);
xnor U7083 (N_7083,In_3895,In_1778);
nand U7084 (N_7084,In_4813,In_4054);
xnor U7085 (N_7085,In_529,In_2072);
nor U7086 (N_7086,In_1597,In_668);
nand U7087 (N_7087,In_4611,In_831);
or U7088 (N_7088,In_184,In_2456);
and U7089 (N_7089,In_3041,In_722);
or U7090 (N_7090,In_507,In_3183);
nor U7091 (N_7091,In_419,In_4257);
nand U7092 (N_7092,In_834,In_911);
xnor U7093 (N_7093,In_3731,In_4353);
and U7094 (N_7094,In_4695,In_4718);
nor U7095 (N_7095,In_2292,In_189);
and U7096 (N_7096,In_694,In_2954);
xor U7097 (N_7097,In_871,In_1358);
and U7098 (N_7098,In_3512,In_4491);
nor U7099 (N_7099,In_4337,In_3795);
or U7100 (N_7100,In_735,In_1964);
xor U7101 (N_7101,In_2330,In_3884);
xnor U7102 (N_7102,In_4490,In_2626);
xor U7103 (N_7103,In_2929,In_2291);
and U7104 (N_7104,In_967,In_2168);
nor U7105 (N_7105,In_3675,In_2292);
xnor U7106 (N_7106,In_4525,In_3763);
or U7107 (N_7107,In_1431,In_4283);
and U7108 (N_7108,In_372,In_1260);
and U7109 (N_7109,In_4194,In_1120);
xor U7110 (N_7110,In_4612,In_1591);
nand U7111 (N_7111,In_4620,In_2255);
xnor U7112 (N_7112,In_1621,In_949);
nand U7113 (N_7113,In_4654,In_3982);
and U7114 (N_7114,In_1068,In_4473);
nor U7115 (N_7115,In_428,In_810);
nor U7116 (N_7116,In_1121,In_1680);
and U7117 (N_7117,In_2039,In_153);
and U7118 (N_7118,In_3899,In_2890);
nor U7119 (N_7119,In_1123,In_491);
and U7120 (N_7120,In_1177,In_3677);
and U7121 (N_7121,In_4937,In_1854);
or U7122 (N_7122,In_2515,In_4298);
nor U7123 (N_7123,In_2967,In_4076);
nand U7124 (N_7124,In_1316,In_1389);
xor U7125 (N_7125,In_2673,In_4295);
nor U7126 (N_7126,In_4304,In_970);
or U7127 (N_7127,In_3220,In_1);
and U7128 (N_7128,In_3038,In_21);
xnor U7129 (N_7129,In_4641,In_3816);
nor U7130 (N_7130,In_2936,In_3134);
or U7131 (N_7131,In_764,In_2379);
nor U7132 (N_7132,In_4461,In_2720);
nand U7133 (N_7133,In_1846,In_3711);
nand U7134 (N_7134,In_2014,In_2447);
and U7135 (N_7135,In_1367,In_1944);
or U7136 (N_7136,In_241,In_3706);
xnor U7137 (N_7137,In_520,In_2925);
nand U7138 (N_7138,In_376,In_1063);
xor U7139 (N_7139,In_35,In_1381);
or U7140 (N_7140,In_1765,In_1294);
or U7141 (N_7141,In_3918,In_3597);
or U7142 (N_7142,In_3516,In_3942);
nand U7143 (N_7143,In_892,In_2263);
or U7144 (N_7144,In_3701,In_3430);
nor U7145 (N_7145,In_1786,In_2305);
and U7146 (N_7146,In_1609,In_978);
xnor U7147 (N_7147,In_3901,In_441);
nand U7148 (N_7148,In_40,In_4575);
or U7149 (N_7149,In_728,In_2665);
and U7150 (N_7150,In_3103,In_2692);
and U7151 (N_7151,In_526,In_1372);
or U7152 (N_7152,In_1787,In_3220);
or U7153 (N_7153,In_4370,In_3797);
xnor U7154 (N_7154,In_4428,In_3625);
nor U7155 (N_7155,In_2577,In_3971);
and U7156 (N_7156,In_1842,In_148);
nor U7157 (N_7157,In_4619,In_1779);
nand U7158 (N_7158,In_1567,In_3989);
or U7159 (N_7159,In_4362,In_3597);
and U7160 (N_7160,In_4359,In_2244);
nand U7161 (N_7161,In_766,In_2343);
nor U7162 (N_7162,In_4703,In_514);
and U7163 (N_7163,In_3641,In_1380);
nor U7164 (N_7164,In_4494,In_3131);
xor U7165 (N_7165,In_4875,In_1681);
or U7166 (N_7166,In_3541,In_2445);
and U7167 (N_7167,In_768,In_1188);
nor U7168 (N_7168,In_591,In_222);
nor U7169 (N_7169,In_3630,In_4176);
xor U7170 (N_7170,In_3774,In_3453);
or U7171 (N_7171,In_4180,In_3280);
nand U7172 (N_7172,In_1657,In_2368);
xnor U7173 (N_7173,In_2925,In_4897);
nand U7174 (N_7174,In_3015,In_4606);
or U7175 (N_7175,In_4227,In_1747);
xnor U7176 (N_7176,In_712,In_73);
nor U7177 (N_7177,In_2741,In_3735);
nor U7178 (N_7178,In_1499,In_4004);
nor U7179 (N_7179,In_2698,In_2902);
nand U7180 (N_7180,In_781,In_2115);
or U7181 (N_7181,In_704,In_4909);
xor U7182 (N_7182,In_4655,In_1017);
nand U7183 (N_7183,In_4342,In_1822);
or U7184 (N_7184,In_1184,In_4448);
or U7185 (N_7185,In_52,In_2663);
nor U7186 (N_7186,In_740,In_1400);
and U7187 (N_7187,In_4341,In_663);
and U7188 (N_7188,In_794,In_3720);
nand U7189 (N_7189,In_2087,In_1159);
nor U7190 (N_7190,In_886,In_2474);
nand U7191 (N_7191,In_4772,In_3941);
or U7192 (N_7192,In_371,In_2625);
xnor U7193 (N_7193,In_4820,In_188);
and U7194 (N_7194,In_4717,In_883);
or U7195 (N_7195,In_2630,In_2131);
nor U7196 (N_7196,In_4907,In_1409);
xnor U7197 (N_7197,In_1309,In_2239);
nand U7198 (N_7198,In_32,In_4323);
or U7199 (N_7199,In_2413,In_469);
nor U7200 (N_7200,In_717,In_2674);
and U7201 (N_7201,In_4740,In_3243);
and U7202 (N_7202,In_3055,In_1177);
nand U7203 (N_7203,In_3450,In_1803);
nor U7204 (N_7204,In_2675,In_3027);
and U7205 (N_7205,In_2012,In_163);
nor U7206 (N_7206,In_4210,In_4114);
nand U7207 (N_7207,In_2702,In_1082);
or U7208 (N_7208,In_872,In_4773);
xnor U7209 (N_7209,In_1096,In_322);
xnor U7210 (N_7210,In_1370,In_3090);
or U7211 (N_7211,In_3777,In_4091);
or U7212 (N_7212,In_272,In_389);
nor U7213 (N_7213,In_3457,In_2586);
or U7214 (N_7214,In_885,In_297);
nor U7215 (N_7215,In_3142,In_3696);
nand U7216 (N_7216,In_3046,In_3794);
or U7217 (N_7217,In_472,In_2764);
and U7218 (N_7218,In_1023,In_2070);
and U7219 (N_7219,In_24,In_4825);
and U7220 (N_7220,In_2893,In_3647);
nand U7221 (N_7221,In_3675,In_3438);
and U7222 (N_7222,In_401,In_4004);
or U7223 (N_7223,In_477,In_1849);
nor U7224 (N_7224,In_3327,In_1198);
or U7225 (N_7225,In_394,In_4188);
xor U7226 (N_7226,In_3040,In_3981);
nand U7227 (N_7227,In_696,In_3783);
or U7228 (N_7228,In_1277,In_412);
nor U7229 (N_7229,In_3771,In_1493);
nand U7230 (N_7230,In_85,In_4128);
xnor U7231 (N_7231,In_110,In_186);
and U7232 (N_7232,In_4616,In_2870);
and U7233 (N_7233,In_1671,In_308);
or U7234 (N_7234,In_2040,In_1000);
nor U7235 (N_7235,In_2415,In_247);
or U7236 (N_7236,In_341,In_1621);
and U7237 (N_7237,In_3187,In_4412);
nor U7238 (N_7238,In_1528,In_4462);
or U7239 (N_7239,In_4686,In_4491);
xor U7240 (N_7240,In_604,In_4000);
or U7241 (N_7241,In_1710,In_4279);
or U7242 (N_7242,In_4297,In_478);
nand U7243 (N_7243,In_3016,In_130);
nand U7244 (N_7244,In_4553,In_1642);
nand U7245 (N_7245,In_4457,In_2431);
xnor U7246 (N_7246,In_2006,In_760);
and U7247 (N_7247,In_1136,In_3429);
xnor U7248 (N_7248,In_2821,In_2999);
nor U7249 (N_7249,In_1768,In_2927);
or U7250 (N_7250,In_1985,In_1846);
xor U7251 (N_7251,In_416,In_3487);
and U7252 (N_7252,In_3048,In_4750);
xnor U7253 (N_7253,In_797,In_522);
nor U7254 (N_7254,In_3436,In_1565);
nand U7255 (N_7255,In_3165,In_3483);
or U7256 (N_7256,In_1176,In_3873);
xor U7257 (N_7257,In_3375,In_4836);
nand U7258 (N_7258,In_2885,In_601);
xor U7259 (N_7259,In_1435,In_4727);
nand U7260 (N_7260,In_2517,In_2811);
xnor U7261 (N_7261,In_2626,In_1326);
xor U7262 (N_7262,In_4375,In_4602);
nor U7263 (N_7263,In_141,In_991);
xor U7264 (N_7264,In_969,In_3550);
or U7265 (N_7265,In_4548,In_749);
nor U7266 (N_7266,In_295,In_2927);
and U7267 (N_7267,In_432,In_2058);
or U7268 (N_7268,In_1195,In_2876);
xor U7269 (N_7269,In_838,In_2465);
nand U7270 (N_7270,In_2599,In_533);
and U7271 (N_7271,In_3354,In_2463);
and U7272 (N_7272,In_4611,In_2474);
nand U7273 (N_7273,In_4787,In_2576);
nor U7274 (N_7274,In_959,In_2456);
xnor U7275 (N_7275,In_2458,In_440);
and U7276 (N_7276,In_966,In_4423);
nor U7277 (N_7277,In_3007,In_1799);
nor U7278 (N_7278,In_1912,In_1118);
nor U7279 (N_7279,In_1713,In_1408);
or U7280 (N_7280,In_3942,In_4406);
xor U7281 (N_7281,In_2847,In_2084);
xor U7282 (N_7282,In_2986,In_417);
xor U7283 (N_7283,In_4091,In_1449);
nor U7284 (N_7284,In_4901,In_3410);
and U7285 (N_7285,In_1705,In_3941);
nor U7286 (N_7286,In_3506,In_4858);
and U7287 (N_7287,In_619,In_3075);
or U7288 (N_7288,In_1662,In_3923);
and U7289 (N_7289,In_3013,In_2787);
xor U7290 (N_7290,In_879,In_2305);
xor U7291 (N_7291,In_4334,In_2732);
nand U7292 (N_7292,In_1473,In_4572);
and U7293 (N_7293,In_1836,In_3770);
xor U7294 (N_7294,In_1819,In_1808);
xnor U7295 (N_7295,In_4854,In_3518);
or U7296 (N_7296,In_4323,In_1846);
nand U7297 (N_7297,In_4744,In_1341);
and U7298 (N_7298,In_133,In_2735);
nand U7299 (N_7299,In_448,In_4784);
xnor U7300 (N_7300,In_3457,In_3706);
or U7301 (N_7301,In_2817,In_569);
or U7302 (N_7302,In_1801,In_2769);
xor U7303 (N_7303,In_2282,In_1152);
nand U7304 (N_7304,In_3721,In_3679);
and U7305 (N_7305,In_2369,In_3551);
nor U7306 (N_7306,In_1319,In_1519);
nor U7307 (N_7307,In_586,In_239);
and U7308 (N_7308,In_1498,In_2582);
nor U7309 (N_7309,In_996,In_3389);
xnor U7310 (N_7310,In_3360,In_4955);
nor U7311 (N_7311,In_1670,In_3726);
nor U7312 (N_7312,In_1170,In_1435);
and U7313 (N_7313,In_305,In_1085);
or U7314 (N_7314,In_1639,In_4382);
xor U7315 (N_7315,In_2357,In_2038);
or U7316 (N_7316,In_2755,In_1891);
xnor U7317 (N_7317,In_780,In_1100);
and U7318 (N_7318,In_1526,In_297);
xor U7319 (N_7319,In_4573,In_3923);
xnor U7320 (N_7320,In_2716,In_344);
and U7321 (N_7321,In_3217,In_1435);
nor U7322 (N_7322,In_4075,In_95);
xnor U7323 (N_7323,In_1590,In_292);
or U7324 (N_7324,In_3422,In_2209);
xor U7325 (N_7325,In_4934,In_4010);
or U7326 (N_7326,In_2335,In_1921);
and U7327 (N_7327,In_4474,In_1616);
nor U7328 (N_7328,In_4066,In_1265);
nor U7329 (N_7329,In_2139,In_817);
or U7330 (N_7330,In_4778,In_3035);
nor U7331 (N_7331,In_4805,In_291);
nor U7332 (N_7332,In_1630,In_1354);
nor U7333 (N_7333,In_611,In_4571);
nor U7334 (N_7334,In_39,In_2547);
nand U7335 (N_7335,In_1560,In_3084);
xor U7336 (N_7336,In_2520,In_4418);
nand U7337 (N_7337,In_2512,In_4531);
nand U7338 (N_7338,In_721,In_3446);
or U7339 (N_7339,In_4842,In_3062);
nor U7340 (N_7340,In_229,In_4744);
or U7341 (N_7341,In_3099,In_4624);
or U7342 (N_7342,In_1435,In_3392);
and U7343 (N_7343,In_149,In_1053);
nor U7344 (N_7344,In_370,In_714);
nor U7345 (N_7345,In_2418,In_3871);
and U7346 (N_7346,In_1254,In_4738);
or U7347 (N_7347,In_1624,In_835);
nor U7348 (N_7348,In_3641,In_3103);
xnor U7349 (N_7349,In_2631,In_65);
and U7350 (N_7350,In_1344,In_3025);
nand U7351 (N_7351,In_1728,In_2625);
and U7352 (N_7352,In_1152,In_2705);
or U7353 (N_7353,In_2019,In_2163);
nor U7354 (N_7354,In_2778,In_1871);
xor U7355 (N_7355,In_3371,In_3392);
nor U7356 (N_7356,In_1609,In_1474);
nand U7357 (N_7357,In_4228,In_1353);
and U7358 (N_7358,In_699,In_2965);
nand U7359 (N_7359,In_2091,In_761);
nand U7360 (N_7360,In_4388,In_4781);
nand U7361 (N_7361,In_2110,In_828);
or U7362 (N_7362,In_4192,In_2550);
or U7363 (N_7363,In_2784,In_4045);
nor U7364 (N_7364,In_3132,In_1397);
or U7365 (N_7365,In_3856,In_1356);
and U7366 (N_7366,In_4673,In_598);
xor U7367 (N_7367,In_1769,In_4797);
or U7368 (N_7368,In_2211,In_3333);
xnor U7369 (N_7369,In_4886,In_817);
and U7370 (N_7370,In_3079,In_1056);
xor U7371 (N_7371,In_860,In_4315);
xnor U7372 (N_7372,In_2295,In_1307);
and U7373 (N_7373,In_2373,In_1731);
nand U7374 (N_7374,In_239,In_3547);
or U7375 (N_7375,In_2217,In_3812);
nor U7376 (N_7376,In_170,In_3765);
nor U7377 (N_7377,In_4338,In_4945);
nand U7378 (N_7378,In_2943,In_2271);
xnor U7379 (N_7379,In_1123,In_2166);
and U7380 (N_7380,In_1627,In_1950);
or U7381 (N_7381,In_988,In_1445);
nor U7382 (N_7382,In_4613,In_85);
nand U7383 (N_7383,In_688,In_2449);
nor U7384 (N_7384,In_3606,In_1959);
nand U7385 (N_7385,In_1103,In_582);
nor U7386 (N_7386,In_3492,In_3221);
nand U7387 (N_7387,In_4006,In_1256);
nor U7388 (N_7388,In_1162,In_312);
and U7389 (N_7389,In_874,In_4104);
and U7390 (N_7390,In_408,In_2259);
nand U7391 (N_7391,In_2960,In_1338);
nor U7392 (N_7392,In_2169,In_1279);
or U7393 (N_7393,In_4367,In_2564);
xnor U7394 (N_7394,In_518,In_3831);
and U7395 (N_7395,In_4247,In_202);
or U7396 (N_7396,In_1747,In_3954);
and U7397 (N_7397,In_600,In_2913);
nand U7398 (N_7398,In_4266,In_1070);
nor U7399 (N_7399,In_2668,In_4786);
xor U7400 (N_7400,In_1845,In_4354);
nor U7401 (N_7401,In_2560,In_4910);
xor U7402 (N_7402,In_770,In_4848);
and U7403 (N_7403,In_2293,In_66);
nand U7404 (N_7404,In_1322,In_3448);
or U7405 (N_7405,In_2788,In_3862);
nand U7406 (N_7406,In_2789,In_4717);
nor U7407 (N_7407,In_3932,In_2476);
nor U7408 (N_7408,In_1522,In_825);
or U7409 (N_7409,In_424,In_758);
nand U7410 (N_7410,In_830,In_3496);
nor U7411 (N_7411,In_2349,In_499);
and U7412 (N_7412,In_77,In_2058);
and U7413 (N_7413,In_4221,In_1630);
xor U7414 (N_7414,In_1685,In_2700);
and U7415 (N_7415,In_1685,In_4365);
and U7416 (N_7416,In_4144,In_2046);
xor U7417 (N_7417,In_4162,In_1273);
nand U7418 (N_7418,In_1598,In_1027);
and U7419 (N_7419,In_1832,In_3886);
and U7420 (N_7420,In_1521,In_1136);
nor U7421 (N_7421,In_3593,In_52);
nor U7422 (N_7422,In_205,In_2639);
and U7423 (N_7423,In_4967,In_3422);
nand U7424 (N_7424,In_3483,In_2213);
nor U7425 (N_7425,In_4137,In_2889);
nand U7426 (N_7426,In_739,In_551);
or U7427 (N_7427,In_2728,In_1752);
xor U7428 (N_7428,In_3269,In_215);
nor U7429 (N_7429,In_2180,In_4325);
nor U7430 (N_7430,In_2266,In_659);
and U7431 (N_7431,In_322,In_2999);
and U7432 (N_7432,In_2269,In_3710);
or U7433 (N_7433,In_4607,In_3724);
nor U7434 (N_7434,In_2940,In_3711);
nand U7435 (N_7435,In_2854,In_4598);
nand U7436 (N_7436,In_3222,In_34);
xnor U7437 (N_7437,In_2796,In_2335);
nor U7438 (N_7438,In_979,In_1065);
and U7439 (N_7439,In_1471,In_3720);
or U7440 (N_7440,In_1576,In_2433);
and U7441 (N_7441,In_4201,In_4536);
xor U7442 (N_7442,In_4626,In_207);
or U7443 (N_7443,In_744,In_4956);
nor U7444 (N_7444,In_660,In_4693);
and U7445 (N_7445,In_1725,In_285);
and U7446 (N_7446,In_713,In_1053);
nand U7447 (N_7447,In_1309,In_1251);
and U7448 (N_7448,In_2309,In_1514);
and U7449 (N_7449,In_2798,In_1043);
nand U7450 (N_7450,In_3277,In_3432);
xor U7451 (N_7451,In_1773,In_3968);
xor U7452 (N_7452,In_3337,In_3914);
and U7453 (N_7453,In_4417,In_2557);
xor U7454 (N_7454,In_298,In_4947);
or U7455 (N_7455,In_1798,In_1616);
xnor U7456 (N_7456,In_2273,In_3814);
xnor U7457 (N_7457,In_2345,In_4234);
nand U7458 (N_7458,In_593,In_2577);
nand U7459 (N_7459,In_3214,In_3888);
nand U7460 (N_7460,In_3867,In_4452);
nand U7461 (N_7461,In_489,In_289);
nor U7462 (N_7462,In_2018,In_96);
xor U7463 (N_7463,In_4523,In_249);
nand U7464 (N_7464,In_3734,In_3664);
nand U7465 (N_7465,In_459,In_2360);
xor U7466 (N_7466,In_163,In_4717);
or U7467 (N_7467,In_4842,In_3312);
and U7468 (N_7468,In_1572,In_3011);
and U7469 (N_7469,In_4682,In_2780);
nor U7470 (N_7470,In_4478,In_4982);
and U7471 (N_7471,In_4605,In_4480);
xor U7472 (N_7472,In_1037,In_3657);
or U7473 (N_7473,In_3187,In_2166);
xor U7474 (N_7474,In_830,In_1082);
nand U7475 (N_7475,In_217,In_4282);
or U7476 (N_7476,In_253,In_365);
and U7477 (N_7477,In_2310,In_3069);
nand U7478 (N_7478,In_4075,In_4786);
or U7479 (N_7479,In_3460,In_2674);
nor U7480 (N_7480,In_2465,In_4732);
nand U7481 (N_7481,In_903,In_2969);
nor U7482 (N_7482,In_3402,In_3326);
xnor U7483 (N_7483,In_3497,In_291);
or U7484 (N_7484,In_2630,In_527);
and U7485 (N_7485,In_554,In_262);
or U7486 (N_7486,In_4329,In_3594);
nand U7487 (N_7487,In_4384,In_1408);
and U7488 (N_7488,In_1042,In_931);
nand U7489 (N_7489,In_1135,In_3976);
xor U7490 (N_7490,In_1466,In_4680);
and U7491 (N_7491,In_1587,In_2209);
xor U7492 (N_7492,In_2968,In_621);
nand U7493 (N_7493,In_2069,In_3749);
nand U7494 (N_7494,In_1811,In_3596);
or U7495 (N_7495,In_4400,In_2938);
nand U7496 (N_7496,In_4725,In_3283);
nor U7497 (N_7497,In_1861,In_2963);
nand U7498 (N_7498,In_3192,In_1749);
or U7499 (N_7499,In_3287,In_334);
nand U7500 (N_7500,In_1406,In_546);
nand U7501 (N_7501,In_977,In_2086);
and U7502 (N_7502,In_99,In_2007);
or U7503 (N_7503,In_3130,In_2729);
and U7504 (N_7504,In_1263,In_3206);
nand U7505 (N_7505,In_3429,In_1152);
nand U7506 (N_7506,In_327,In_3440);
or U7507 (N_7507,In_1413,In_394);
nand U7508 (N_7508,In_2135,In_2150);
nor U7509 (N_7509,In_4223,In_3312);
and U7510 (N_7510,In_912,In_3679);
or U7511 (N_7511,In_982,In_662);
or U7512 (N_7512,In_2407,In_2733);
or U7513 (N_7513,In_913,In_1819);
xnor U7514 (N_7514,In_1634,In_3922);
and U7515 (N_7515,In_76,In_897);
xnor U7516 (N_7516,In_2666,In_1455);
or U7517 (N_7517,In_2668,In_4371);
nand U7518 (N_7518,In_2741,In_394);
nand U7519 (N_7519,In_4355,In_3260);
xnor U7520 (N_7520,In_2238,In_690);
xor U7521 (N_7521,In_407,In_292);
and U7522 (N_7522,In_3369,In_2738);
and U7523 (N_7523,In_3018,In_1756);
and U7524 (N_7524,In_3828,In_2954);
nor U7525 (N_7525,In_3454,In_3789);
or U7526 (N_7526,In_2851,In_1875);
nand U7527 (N_7527,In_2832,In_508);
nor U7528 (N_7528,In_3908,In_4092);
or U7529 (N_7529,In_2092,In_1509);
and U7530 (N_7530,In_3260,In_2023);
or U7531 (N_7531,In_2405,In_2569);
nor U7532 (N_7532,In_235,In_3213);
or U7533 (N_7533,In_704,In_4078);
nand U7534 (N_7534,In_1029,In_855);
and U7535 (N_7535,In_1615,In_3799);
nand U7536 (N_7536,In_787,In_1575);
or U7537 (N_7537,In_125,In_963);
and U7538 (N_7538,In_3859,In_4780);
and U7539 (N_7539,In_2529,In_3296);
xor U7540 (N_7540,In_214,In_3039);
nor U7541 (N_7541,In_4760,In_4088);
nand U7542 (N_7542,In_1617,In_2764);
nand U7543 (N_7543,In_44,In_1806);
nand U7544 (N_7544,In_3864,In_4005);
or U7545 (N_7545,In_3908,In_255);
nor U7546 (N_7546,In_4479,In_1982);
and U7547 (N_7547,In_4529,In_3142);
nor U7548 (N_7548,In_1053,In_668);
and U7549 (N_7549,In_1443,In_2659);
xor U7550 (N_7550,In_3393,In_4625);
nor U7551 (N_7551,In_194,In_1720);
or U7552 (N_7552,In_1452,In_2484);
xnor U7553 (N_7553,In_3677,In_4631);
and U7554 (N_7554,In_260,In_3268);
nor U7555 (N_7555,In_3970,In_178);
and U7556 (N_7556,In_4417,In_4841);
and U7557 (N_7557,In_248,In_432);
or U7558 (N_7558,In_1930,In_3253);
or U7559 (N_7559,In_771,In_3648);
nor U7560 (N_7560,In_4017,In_3879);
nor U7561 (N_7561,In_295,In_2285);
nor U7562 (N_7562,In_3345,In_4358);
and U7563 (N_7563,In_1216,In_1975);
and U7564 (N_7564,In_3171,In_1602);
xor U7565 (N_7565,In_4598,In_1595);
xnor U7566 (N_7566,In_2536,In_3996);
xor U7567 (N_7567,In_2050,In_4279);
nor U7568 (N_7568,In_4777,In_2373);
and U7569 (N_7569,In_4826,In_3460);
and U7570 (N_7570,In_1299,In_834);
nor U7571 (N_7571,In_3884,In_2898);
and U7572 (N_7572,In_695,In_1479);
nand U7573 (N_7573,In_4944,In_2174);
xnor U7574 (N_7574,In_1909,In_1820);
nand U7575 (N_7575,In_1347,In_4352);
or U7576 (N_7576,In_4593,In_507);
and U7577 (N_7577,In_3784,In_4717);
xnor U7578 (N_7578,In_611,In_4792);
and U7579 (N_7579,In_3909,In_4433);
and U7580 (N_7580,In_2334,In_709);
and U7581 (N_7581,In_1635,In_570);
or U7582 (N_7582,In_3344,In_271);
or U7583 (N_7583,In_4063,In_1581);
nand U7584 (N_7584,In_41,In_4441);
and U7585 (N_7585,In_418,In_1612);
and U7586 (N_7586,In_4330,In_4986);
and U7587 (N_7587,In_3935,In_3393);
and U7588 (N_7588,In_3551,In_3662);
or U7589 (N_7589,In_1930,In_2383);
and U7590 (N_7590,In_4417,In_2317);
nor U7591 (N_7591,In_4081,In_2867);
and U7592 (N_7592,In_597,In_4352);
nand U7593 (N_7593,In_531,In_2008);
and U7594 (N_7594,In_4076,In_3753);
xnor U7595 (N_7595,In_4251,In_1191);
xor U7596 (N_7596,In_517,In_4155);
nor U7597 (N_7597,In_1794,In_1345);
nand U7598 (N_7598,In_4274,In_2349);
or U7599 (N_7599,In_4141,In_3338);
nand U7600 (N_7600,In_3382,In_3151);
nor U7601 (N_7601,In_1798,In_1979);
nor U7602 (N_7602,In_2631,In_1896);
xnor U7603 (N_7603,In_390,In_1331);
nand U7604 (N_7604,In_110,In_4702);
nand U7605 (N_7605,In_3012,In_1596);
or U7606 (N_7606,In_2675,In_2023);
nor U7607 (N_7607,In_4130,In_796);
nor U7608 (N_7608,In_3166,In_3189);
xnor U7609 (N_7609,In_254,In_3968);
and U7610 (N_7610,In_152,In_2233);
nor U7611 (N_7611,In_1109,In_2883);
nand U7612 (N_7612,In_3391,In_4357);
and U7613 (N_7613,In_2405,In_2348);
or U7614 (N_7614,In_2406,In_2899);
or U7615 (N_7615,In_3008,In_422);
nand U7616 (N_7616,In_2240,In_249);
xor U7617 (N_7617,In_1121,In_3947);
or U7618 (N_7618,In_1142,In_660);
nand U7619 (N_7619,In_2961,In_4980);
and U7620 (N_7620,In_4999,In_3370);
or U7621 (N_7621,In_2628,In_702);
nand U7622 (N_7622,In_1674,In_4738);
and U7623 (N_7623,In_3265,In_2281);
nor U7624 (N_7624,In_1444,In_671);
nand U7625 (N_7625,In_421,In_1722);
and U7626 (N_7626,In_2728,In_1609);
nor U7627 (N_7627,In_1820,In_1160);
xor U7628 (N_7628,In_4610,In_4791);
xnor U7629 (N_7629,In_1932,In_2503);
and U7630 (N_7630,In_2446,In_1162);
or U7631 (N_7631,In_1514,In_1389);
or U7632 (N_7632,In_1696,In_2265);
and U7633 (N_7633,In_1561,In_3488);
and U7634 (N_7634,In_1389,In_3166);
nor U7635 (N_7635,In_1611,In_4526);
nand U7636 (N_7636,In_3074,In_3169);
nand U7637 (N_7637,In_82,In_3384);
and U7638 (N_7638,In_4702,In_1182);
xor U7639 (N_7639,In_876,In_2315);
xnor U7640 (N_7640,In_3240,In_2366);
and U7641 (N_7641,In_1589,In_1373);
and U7642 (N_7642,In_681,In_1182);
nand U7643 (N_7643,In_102,In_3395);
xor U7644 (N_7644,In_3191,In_2536);
xor U7645 (N_7645,In_1010,In_4464);
and U7646 (N_7646,In_3794,In_3906);
and U7647 (N_7647,In_3362,In_999);
or U7648 (N_7648,In_549,In_298);
and U7649 (N_7649,In_296,In_3885);
nand U7650 (N_7650,In_2574,In_3353);
and U7651 (N_7651,In_603,In_4237);
and U7652 (N_7652,In_4125,In_2772);
nand U7653 (N_7653,In_2920,In_3102);
or U7654 (N_7654,In_4372,In_1401);
and U7655 (N_7655,In_2691,In_2464);
and U7656 (N_7656,In_1827,In_370);
and U7657 (N_7657,In_4094,In_762);
and U7658 (N_7658,In_1622,In_898);
xnor U7659 (N_7659,In_48,In_1303);
and U7660 (N_7660,In_272,In_1329);
and U7661 (N_7661,In_3452,In_1743);
or U7662 (N_7662,In_4277,In_4851);
nor U7663 (N_7663,In_3318,In_1382);
and U7664 (N_7664,In_1036,In_3069);
nand U7665 (N_7665,In_4637,In_371);
nand U7666 (N_7666,In_4490,In_4957);
xnor U7667 (N_7667,In_2768,In_3511);
nand U7668 (N_7668,In_2004,In_197);
and U7669 (N_7669,In_1493,In_3921);
nor U7670 (N_7670,In_1854,In_3001);
nor U7671 (N_7671,In_4639,In_3520);
xor U7672 (N_7672,In_3496,In_4414);
xor U7673 (N_7673,In_57,In_3547);
and U7674 (N_7674,In_275,In_3063);
and U7675 (N_7675,In_4692,In_1612);
nand U7676 (N_7676,In_3493,In_3955);
xor U7677 (N_7677,In_2140,In_1745);
and U7678 (N_7678,In_2660,In_4846);
and U7679 (N_7679,In_3573,In_3462);
nor U7680 (N_7680,In_2510,In_3449);
xnor U7681 (N_7681,In_1918,In_1677);
xnor U7682 (N_7682,In_1135,In_3610);
nand U7683 (N_7683,In_3739,In_4491);
and U7684 (N_7684,In_1572,In_4137);
nor U7685 (N_7685,In_782,In_2053);
nor U7686 (N_7686,In_3801,In_870);
nor U7687 (N_7687,In_2414,In_1417);
xor U7688 (N_7688,In_2762,In_2207);
and U7689 (N_7689,In_4448,In_2413);
nor U7690 (N_7690,In_3630,In_2491);
xor U7691 (N_7691,In_3631,In_2284);
and U7692 (N_7692,In_1430,In_4150);
nor U7693 (N_7693,In_4261,In_3884);
nand U7694 (N_7694,In_809,In_2010);
and U7695 (N_7695,In_2501,In_616);
or U7696 (N_7696,In_1734,In_938);
nor U7697 (N_7697,In_4779,In_2401);
nand U7698 (N_7698,In_826,In_2467);
nand U7699 (N_7699,In_4678,In_763);
nand U7700 (N_7700,In_3467,In_716);
and U7701 (N_7701,In_3681,In_3134);
xor U7702 (N_7702,In_1062,In_2754);
nand U7703 (N_7703,In_3342,In_3654);
xor U7704 (N_7704,In_2198,In_3096);
or U7705 (N_7705,In_2510,In_1210);
and U7706 (N_7706,In_558,In_2602);
or U7707 (N_7707,In_3711,In_2861);
or U7708 (N_7708,In_2114,In_3129);
or U7709 (N_7709,In_1553,In_3877);
xor U7710 (N_7710,In_2955,In_1291);
or U7711 (N_7711,In_1554,In_4923);
or U7712 (N_7712,In_3561,In_2150);
xor U7713 (N_7713,In_1403,In_30);
or U7714 (N_7714,In_161,In_1189);
xnor U7715 (N_7715,In_3054,In_555);
and U7716 (N_7716,In_4810,In_3656);
nor U7717 (N_7717,In_2758,In_1508);
and U7718 (N_7718,In_3448,In_2736);
nor U7719 (N_7719,In_2177,In_4318);
nor U7720 (N_7720,In_512,In_4561);
nor U7721 (N_7721,In_4237,In_4725);
nor U7722 (N_7722,In_4685,In_4382);
or U7723 (N_7723,In_4043,In_752);
nor U7724 (N_7724,In_4744,In_1581);
and U7725 (N_7725,In_1534,In_1378);
xnor U7726 (N_7726,In_2460,In_1722);
and U7727 (N_7727,In_1877,In_3126);
or U7728 (N_7728,In_4209,In_2611);
nor U7729 (N_7729,In_945,In_1157);
nand U7730 (N_7730,In_669,In_4501);
or U7731 (N_7731,In_1753,In_2692);
nor U7732 (N_7732,In_2843,In_335);
or U7733 (N_7733,In_4296,In_3785);
nand U7734 (N_7734,In_3332,In_4332);
or U7735 (N_7735,In_337,In_811);
xnor U7736 (N_7736,In_280,In_2409);
nand U7737 (N_7737,In_1370,In_2996);
or U7738 (N_7738,In_3044,In_434);
xnor U7739 (N_7739,In_4518,In_4223);
xnor U7740 (N_7740,In_4690,In_171);
nor U7741 (N_7741,In_3992,In_764);
nor U7742 (N_7742,In_4524,In_84);
xor U7743 (N_7743,In_116,In_2972);
nor U7744 (N_7744,In_3528,In_2499);
nand U7745 (N_7745,In_1652,In_4174);
nand U7746 (N_7746,In_2460,In_84);
and U7747 (N_7747,In_4748,In_3669);
xor U7748 (N_7748,In_1037,In_1767);
and U7749 (N_7749,In_1906,In_4299);
nand U7750 (N_7750,In_1378,In_1031);
or U7751 (N_7751,In_1217,In_569);
and U7752 (N_7752,In_4061,In_2329);
nor U7753 (N_7753,In_3277,In_3928);
nor U7754 (N_7754,In_2873,In_2031);
xor U7755 (N_7755,In_672,In_494);
xor U7756 (N_7756,In_4918,In_82);
nor U7757 (N_7757,In_4679,In_510);
nor U7758 (N_7758,In_3019,In_4715);
and U7759 (N_7759,In_4944,In_348);
or U7760 (N_7760,In_3881,In_677);
or U7761 (N_7761,In_2135,In_981);
xor U7762 (N_7762,In_3929,In_3376);
and U7763 (N_7763,In_3625,In_1852);
nand U7764 (N_7764,In_4213,In_250);
nand U7765 (N_7765,In_3503,In_4248);
or U7766 (N_7766,In_3702,In_4700);
nor U7767 (N_7767,In_1574,In_1524);
and U7768 (N_7768,In_2443,In_3491);
nor U7769 (N_7769,In_45,In_231);
and U7770 (N_7770,In_987,In_1814);
nand U7771 (N_7771,In_201,In_992);
and U7772 (N_7772,In_3311,In_4863);
or U7773 (N_7773,In_2221,In_4469);
and U7774 (N_7774,In_1055,In_4732);
nand U7775 (N_7775,In_2417,In_2135);
nand U7776 (N_7776,In_2701,In_1966);
nor U7777 (N_7777,In_4088,In_1861);
or U7778 (N_7778,In_3968,In_841);
nor U7779 (N_7779,In_4633,In_790);
xnor U7780 (N_7780,In_3802,In_1303);
xnor U7781 (N_7781,In_4167,In_2229);
or U7782 (N_7782,In_863,In_1763);
nand U7783 (N_7783,In_2832,In_4711);
nand U7784 (N_7784,In_1343,In_2542);
xnor U7785 (N_7785,In_2778,In_19);
nor U7786 (N_7786,In_108,In_901);
nor U7787 (N_7787,In_1351,In_1190);
xor U7788 (N_7788,In_4281,In_3120);
or U7789 (N_7789,In_134,In_1010);
xnor U7790 (N_7790,In_189,In_3532);
and U7791 (N_7791,In_2639,In_4393);
nand U7792 (N_7792,In_3339,In_2309);
or U7793 (N_7793,In_4054,In_2360);
and U7794 (N_7794,In_4097,In_2000);
nor U7795 (N_7795,In_2125,In_269);
or U7796 (N_7796,In_1740,In_3533);
nand U7797 (N_7797,In_2793,In_4106);
and U7798 (N_7798,In_4070,In_2289);
xor U7799 (N_7799,In_4522,In_1556);
xor U7800 (N_7800,In_298,In_3016);
xnor U7801 (N_7801,In_3664,In_508);
or U7802 (N_7802,In_1206,In_3419);
xnor U7803 (N_7803,In_419,In_4780);
nor U7804 (N_7804,In_913,In_3720);
xor U7805 (N_7805,In_3271,In_1142);
or U7806 (N_7806,In_753,In_2186);
and U7807 (N_7807,In_714,In_3768);
nor U7808 (N_7808,In_3511,In_1760);
xnor U7809 (N_7809,In_2552,In_906);
nor U7810 (N_7810,In_4289,In_4765);
nor U7811 (N_7811,In_634,In_272);
or U7812 (N_7812,In_1049,In_927);
or U7813 (N_7813,In_2549,In_2475);
or U7814 (N_7814,In_1740,In_3034);
nand U7815 (N_7815,In_1426,In_1356);
and U7816 (N_7816,In_3787,In_2007);
nand U7817 (N_7817,In_2812,In_4824);
and U7818 (N_7818,In_3919,In_3193);
and U7819 (N_7819,In_3538,In_2246);
nor U7820 (N_7820,In_2051,In_648);
or U7821 (N_7821,In_4514,In_4880);
xnor U7822 (N_7822,In_2009,In_1556);
nand U7823 (N_7823,In_2223,In_4720);
and U7824 (N_7824,In_2109,In_2254);
xor U7825 (N_7825,In_112,In_1320);
nor U7826 (N_7826,In_199,In_4829);
or U7827 (N_7827,In_4179,In_3194);
xnor U7828 (N_7828,In_3244,In_1862);
or U7829 (N_7829,In_716,In_2512);
xor U7830 (N_7830,In_2879,In_4321);
and U7831 (N_7831,In_3044,In_2438);
nand U7832 (N_7832,In_2094,In_480);
and U7833 (N_7833,In_30,In_959);
nor U7834 (N_7834,In_246,In_984);
and U7835 (N_7835,In_4220,In_4861);
xnor U7836 (N_7836,In_1849,In_3072);
xnor U7837 (N_7837,In_2780,In_4896);
nor U7838 (N_7838,In_2992,In_4421);
nand U7839 (N_7839,In_2936,In_4111);
xnor U7840 (N_7840,In_462,In_3848);
nor U7841 (N_7841,In_3927,In_3271);
or U7842 (N_7842,In_3036,In_1024);
xnor U7843 (N_7843,In_3170,In_748);
xor U7844 (N_7844,In_4443,In_2288);
nor U7845 (N_7845,In_3744,In_1709);
nor U7846 (N_7846,In_3081,In_2086);
and U7847 (N_7847,In_815,In_4928);
or U7848 (N_7848,In_730,In_767);
nand U7849 (N_7849,In_3817,In_605);
xor U7850 (N_7850,In_3442,In_2968);
nand U7851 (N_7851,In_2448,In_829);
nor U7852 (N_7852,In_4890,In_2484);
xnor U7853 (N_7853,In_2087,In_2554);
and U7854 (N_7854,In_1295,In_3616);
and U7855 (N_7855,In_3910,In_2617);
nor U7856 (N_7856,In_175,In_3037);
or U7857 (N_7857,In_3258,In_3861);
xor U7858 (N_7858,In_2953,In_2820);
or U7859 (N_7859,In_4380,In_1986);
or U7860 (N_7860,In_3059,In_49);
nor U7861 (N_7861,In_942,In_714);
nor U7862 (N_7862,In_1920,In_151);
or U7863 (N_7863,In_3346,In_3365);
or U7864 (N_7864,In_4800,In_336);
xor U7865 (N_7865,In_4592,In_624);
nor U7866 (N_7866,In_1012,In_2335);
or U7867 (N_7867,In_2521,In_2627);
or U7868 (N_7868,In_4065,In_1191);
nand U7869 (N_7869,In_2346,In_3095);
xnor U7870 (N_7870,In_2835,In_4590);
nor U7871 (N_7871,In_1695,In_3034);
and U7872 (N_7872,In_4395,In_1773);
nand U7873 (N_7873,In_4687,In_3929);
or U7874 (N_7874,In_222,In_1868);
xnor U7875 (N_7875,In_2217,In_3204);
or U7876 (N_7876,In_683,In_4851);
nand U7877 (N_7877,In_3023,In_2530);
xnor U7878 (N_7878,In_3513,In_61);
or U7879 (N_7879,In_4348,In_1807);
and U7880 (N_7880,In_3435,In_1869);
xnor U7881 (N_7881,In_462,In_3696);
nor U7882 (N_7882,In_2403,In_2216);
xor U7883 (N_7883,In_2563,In_1388);
nor U7884 (N_7884,In_130,In_2412);
xnor U7885 (N_7885,In_2671,In_3145);
or U7886 (N_7886,In_4990,In_568);
xnor U7887 (N_7887,In_1623,In_3655);
and U7888 (N_7888,In_2039,In_2288);
xor U7889 (N_7889,In_1687,In_1094);
nand U7890 (N_7890,In_12,In_3308);
nand U7891 (N_7891,In_1853,In_1536);
or U7892 (N_7892,In_1523,In_2373);
or U7893 (N_7893,In_2247,In_1089);
nand U7894 (N_7894,In_4736,In_2857);
or U7895 (N_7895,In_3975,In_4398);
and U7896 (N_7896,In_4515,In_439);
nand U7897 (N_7897,In_813,In_151);
nor U7898 (N_7898,In_2317,In_4756);
and U7899 (N_7899,In_1670,In_1405);
nor U7900 (N_7900,In_702,In_1629);
xor U7901 (N_7901,In_3206,In_1112);
or U7902 (N_7902,In_2897,In_756);
nand U7903 (N_7903,In_2592,In_407);
nand U7904 (N_7904,In_3482,In_3959);
nand U7905 (N_7905,In_2215,In_1861);
and U7906 (N_7906,In_2494,In_41);
xor U7907 (N_7907,In_1757,In_4774);
nand U7908 (N_7908,In_2430,In_1395);
and U7909 (N_7909,In_2240,In_1926);
xnor U7910 (N_7910,In_3716,In_4897);
nor U7911 (N_7911,In_497,In_3733);
xor U7912 (N_7912,In_3305,In_4007);
and U7913 (N_7913,In_353,In_1181);
nand U7914 (N_7914,In_3544,In_3761);
xor U7915 (N_7915,In_3465,In_4466);
xor U7916 (N_7916,In_4666,In_4260);
nand U7917 (N_7917,In_81,In_1348);
xnor U7918 (N_7918,In_3223,In_594);
and U7919 (N_7919,In_478,In_4605);
and U7920 (N_7920,In_3524,In_4941);
nor U7921 (N_7921,In_4567,In_829);
or U7922 (N_7922,In_2056,In_2422);
nor U7923 (N_7923,In_1744,In_1986);
or U7924 (N_7924,In_494,In_4653);
nor U7925 (N_7925,In_4092,In_1584);
and U7926 (N_7926,In_2327,In_4074);
nand U7927 (N_7927,In_237,In_4525);
nand U7928 (N_7928,In_4888,In_2109);
or U7929 (N_7929,In_1824,In_4682);
nand U7930 (N_7930,In_1065,In_3786);
nor U7931 (N_7931,In_586,In_115);
nor U7932 (N_7932,In_1602,In_2551);
nand U7933 (N_7933,In_3009,In_3443);
nand U7934 (N_7934,In_2255,In_863);
xor U7935 (N_7935,In_3205,In_4101);
xor U7936 (N_7936,In_1652,In_4243);
or U7937 (N_7937,In_401,In_4550);
nand U7938 (N_7938,In_1434,In_2793);
nor U7939 (N_7939,In_2432,In_4274);
nand U7940 (N_7940,In_984,In_1248);
nand U7941 (N_7941,In_4207,In_2530);
nand U7942 (N_7942,In_4665,In_245);
or U7943 (N_7943,In_4716,In_1640);
nor U7944 (N_7944,In_64,In_50);
nor U7945 (N_7945,In_2321,In_1838);
xor U7946 (N_7946,In_1114,In_4646);
nor U7947 (N_7947,In_3294,In_4913);
or U7948 (N_7948,In_991,In_935);
nand U7949 (N_7949,In_1640,In_911);
nor U7950 (N_7950,In_3573,In_3603);
or U7951 (N_7951,In_2914,In_4738);
nand U7952 (N_7952,In_1890,In_1404);
xor U7953 (N_7953,In_975,In_2248);
and U7954 (N_7954,In_975,In_2462);
or U7955 (N_7955,In_2960,In_4872);
nor U7956 (N_7956,In_3985,In_3889);
xnor U7957 (N_7957,In_1353,In_1521);
nand U7958 (N_7958,In_1094,In_755);
xor U7959 (N_7959,In_1769,In_2542);
xnor U7960 (N_7960,In_897,In_3883);
nand U7961 (N_7961,In_2734,In_4866);
nor U7962 (N_7962,In_1572,In_4547);
nand U7963 (N_7963,In_161,In_1016);
xnor U7964 (N_7964,In_4726,In_4162);
xnor U7965 (N_7965,In_2622,In_4368);
nand U7966 (N_7966,In_4238,In_2944);
nor U7967 (N_7967,In_1787,In_3077);
or U7968 (N_7968,In_1889,In_79);
and U7969 (N_7969,In_3438,In_1142);
and U7970 (N_7970,In_2533,In_232);
xor U7971 (N_7971,In_330,In_1792);
and U7972 (N_7972,In_2873,In_3975);
or U7973 (N_7973,In_2424,In_1177);
and U7974 (N_7974,In_827,In_2009);
or U7975 (N_7975,In_4886,In_763);
nor U7976 (N_7976,In_1765,In_4469);
or U7977 (N_7977,In_443,In_2947);
and U7978 (N_7978,In_3946,In_4035);
and U7979 (N_7979,In_116,In_4060);
nor U7980 (N_7980,In_257,In_2944);
nor U7981 (N_7981,In_2413,In_3947);
or U7982 (N_7982,In_2516,In_2430);
or U7983 (N_7983,In_1975,In_959);
xor U7984 (N_7984,In_879,In_3777);
nand U7985 (N_7985,In_1169,In_2061);
nor U7986 (N_7986,In_2923,In_2873);
nor U7987 (N_7987,In_2848,In_748);
and U7988 (N_7988,In_2599,In_2710);
or U7989 (N_7989,In_3516,In_680);
and U7990 (N_7990,In_2923,In_4214);
nor U7991 (N_7991,In_3069,In_2287);
and U7992 (N_7992,In_3107,In_4989);
nor U7993 (N_7993,In_4899,In_4240);
nor U7994 (N_7994,In_571,In_3864);
nand U7995 (N_7995,In_1259,In_712);
nor U7996 (N_7996,In_2996,In_3903);
xor U7997 (N_7997,In_4028,In_1120);
nor U7998 (N_7998,In_853,In_4842);
and U7999 (N_7999,In_3856,In_2562);
and U8000 (N_8000,In_1816,In_2113);
nand U8001 (N_8001,In_1500,In_545);
nor U8002 (N_8002,In_1005,In_1810);
nor U8003 (N_8003,In_3858,In_3848);
xor U8004 (N_8004,In_471,In_4337);
nand U8005 (N_8005,In_3259,In_1644);
xor U8006 (N_8006,In_3549,In_2039);
nand U8007 (N_8007,In_3271,In_935);
and U8008 (N_8008,In_1403,In_4543);
and U8009 (N_8009,In_726,In_1936);
nand U8010 (N_8010,In_3168,In_3627);
nand U8011 (N_8011,In_1756,In_3219);
nand U8012 (N_8012,In_3229,In_2780);
and U8013 (N_8013,In_4331,In_1091);
or U8014 (N_8014,In_972,In_771);
xnor U8015 (N_8015,In_4684,In_1710);
nor U8016 (N_8016,In_1539,In_3456);
nor U8017 (N_8017,In_3366,In_1705);
and U8018 (N_8018,In_3427,In_4806);
xnor U8019 (N_8019,In_1490,In_185);
and U8020 (N_8020,In_4493,In_154);
or U8021 (N_8021,In_93,In_777);
xor U8022 (N_8022,In_4857,In_2665);
xnor U8023 (N_8023,In_4306,In_4840);
nor U8024 (N_8024,In_152,In_1737);
xor U8025 (N_8025,In_2192,In_2140);
nand U8026 (N_8026,In_574,In_1540);
nand U8027 (N_8027,In_74,In_4443);
and U8028 (N_8028,In_3134,In_826);
nor U8029 (N_8029,In_2353,In_4202);
nor U8030 (N_8030,In_3151,In_2749);
nor U8031 (N_8031,In_4716,In_1313);
nor U8032 (N_8032,In_4917,In_2547);
or U8033 (N_8033,In_3399,In_4698);
and U8034 (N_8034,In_4206,In_2688);
or U8035 (N_8035,In_4817,In_1644);
nand U8036 (N_8036,In_2385,In_3323);
and U8037 (N_8037,In_3077,In_1298);
or U8038 (N_8038,In_2975,In_3922);
or U8039 (N_8039,In_3124,In_2742);
xnor U8040 (N_8040,In_858,In_2291);
nor U8041 (N_8041,In_1020,In_103);
and U8042 (N_8042,In_2287,In_3005);
nand U8043 (N_8043,In_3579,In_4009);
nor U8044 (N_8044,In_861,In_2436);
nor U8045 (N_8045,In_1604,In_3555);
xor U8046 (N_8046,In_3152,In_4097);
nor U8047 (N_8047,In_2355,In_2420);
nand U8048 (N_8048,In_160,In_828);
and U8049 (N_8049,In_48,In_769);
nand U8050 (N_8050,In_1462,In_4184);
or U8051 (N_8051,In_4977,In_2256);
xor U8052 (N_8052,In_4324,In_367);
and U8053 (N_8053,In_1185,In_3247);
and U8054 (N_8054,In_1820,In_1223);
or U8055 (N_8055,In_437,In_125);
or U8056 (N_8056,In_3269,In_1658);
or U8057 (N_8057,In_62,In_2099);
or U8058 (N_8058,In_2553,In_4247);
nand U8059 (N_8059,In_497,In_1310);
xor U8060 (N_8060,In_2049,In_601);
nor U8061 (N_8061,In_3318,In_4058);
and U8062 (N_8062,In_658,In_2444);
xnor U8063 (N_8063,In_146,In_3538);
xor U8064 (N_8064,In_2656,In_3856);
or U8065 (N_8065,In_4230,In_632);
or U8066 (N_8066,In_1257,In_2380);
and U8067 (N_8067,In_2144,In_4881);
xnor U8068 (N_8068,In_1770,In_1327);
nor U8069 (N_8069,In_755,In_4354);
nor U8070 (N_8070,In_600,In_2433);
nor U8071 (N_8071,In_4505,In_1673);
nor U8072 (N_8072,In_192,In_4769);
or U8073 (N_8073,In_1336,In_2606);
or U8074 (N_8074,In_4468,In_1546);
nor U8075 (N_8075,In_2469,In_966);
nand U8076 (N_8076,In_2767,In_2256);
and U8077 (N_8077,In_1177,In_4212);
nor U8078 (N_8078,In_4068,In_753);
nand U8079 (N_8079,In_2203,In_4946);
and U8080 (N_8080,In_4198,In_2190);
or U8081 (N_8081,In_669,In_2599);
nand U8082 (N_8082,In_3806,In_1051);
nor U8083 (N_8083,In_4110,In_872);
or U8084 (N_8084,In_1394,In_1330);
nor U8085 (N_8085,In_1498,In_255);
and U8086 (N_8086,In_3343,In_1068);
nor U8087 (N_8087,In_3577,In_486);
nor U8088 (N_8088,In_3028,In_460);
xnor U8089 (N_8089,In_3555,In_2353);
or U8090 (N_8090,In_3066,In_1570);
and U8091 (N_8091,In_974,In_215);
nor U8092 (N_8092,In_1032,In_29);
xnor U8093 (N_8093,In_3631,In_4187);
xor U8094 (N_8094,In_2657,In_4013);
and U8095 (N_8095,In_4635,In_4333);
and U8096 (N_8096,In_1259,In_3087);
nand U8097 (N_8097,In_164,In_4370);
nand U8098 (N_8098,In_1110,In_3421);
and U8099 (N_8099,In_3296,In_1506);
nand U8100 (N_8100,In_101,In_321);
nand U8101 (N_8101,In_2171,In_2918);
xor U8102 (N_8102,In_1711,In_542);
nand U8103 (N_8103,In_2360,In_2767);
or U8104 (N_8104,In_4306,In_1586);
nand U8105 (N_8105,In_915,In_2039);
and U8106 (N_8106,In_2017,In_1253);
and U8107 (N_8107,In_1431,In_3340);
or U8108 (N_8108,In_3348,In_2013);
or U8109 (N_8109,In_3732,In_2403);
nand U8110 (N_8110,In_2655,In_3639);
xor U8111 (N_8111,In_33,In_1740);
and U8112 (N_8112,In_3374,In_1077);
nor U8113 (N_8113,In_726,In_2539);
or U8114 (N_8114,In_4750,In_4379);
and U8115 (N_8115,In_798,In_2505);
and U8116 (N_8116,In_3603,In_173);
and U8117 (N_8117,In_4949,In_1387);
or U8118 (N_8118,In_4625,In_1666);
or U8119 (N_8119,In_229,In_118);
nor U8120 (N_8120,In_4392,In_1630);
nand U8121 (N_8121,In_1880,In_2244);
xor U8122 (N_8122,In_4048,In_4394);
nor U8123 (N_8123,In_114,In_4169);
nand U8124 (N_8124,In_1140,In_1783);
nor U8125 (N_8125,In_3480,In_4548);
nand U8126 (N_8126,In_2099,In_3177);
nor U8127 (N_8127,In_4268,In_311);
xor U8128 (N_8128,In_1362,In_2667);
xnor U8129 (N_8129,In_2309,In_3171);
and U8130 (N_8130,In_3826,In_2380);
xnor U8131 (N_8131,In_2907,In_2119);
nand U8132 (N_8132,In_771,In_2738);
xnor U8133 (N_8133,In_2409,In_3226);
and U8134 (N_8134,In_1317,In_2592);
nand U8135 (N_8135,In_591,In_4415);
nand U8136 (N_8136,In_153,In_3218);
and U8137 (N_8137,In_1215,In_3786);
or U8138 (N_8138,In_3333,In_230);
nor U8139 (N_8139,In_4130,In_499);
xor U8140 (N_8140,In_3550,In_3599);
xor U8141 (N_8141,In_2202,In_4796);
nand U8142 (N_8142,In_1316,In_1796);
and U8143 (N_8143,In_1084,In_4404);
xor U8144 (N_8144,In_1052,In_4323);
xnor U8145 (N_8145,In_4816,In_2671);
nand U8146 (N_8146,In_1120,In_4366);
and U8147 (N_8147,In_2664,In_4022);
nor U8148 (N_8148,In_3572,In_2896);
and U8149 (N_8149,In_509,In_750);
nor U8150 (N_8150,In_1700,In_4914);
or U8151 (N_8151,In_193,In_2654);
xor U8152 (N_8152,In_3873,In_2052);
or U8153 (N_8153,In_137,In_3972);
xor U8154 (N_8154,In_4116,In_341);
nor U8155 (N_8155,In_2410,In_1711);
or U8156 (N_8156,In_394,In_2308);
nand U8157 (N_8157,In_659,In_1611);
nor U8158 (N_8158,In_1718,In_2558);
nor U8159 (N_8159,In_2653,In_3795);
xnor U8160 (N_8160,In_1629,In_2335);
and U8161 (N_8161,In_2218,In_2381);
and U8162 (N_8162,In_441,In_748);
and U8163 (N_8163,In_1734,In_4526);
xnor U8164 (N_8164,In_1234,In_294);
nor U8165 (N_8165,In_3328,In_843);
nand U8166 (N_8166,In_1476,In_696);
and U8167 (N_8167,In_1539,In_986);
or U8168 (N_8168,In_694,In_2227);
or U8169 (N_8169,In_3080,In_283);
or U8170 (N_8170,In_148,In_402);
nand U8171 (N_8171,In_1154,In_2075);
xnor U8172 (N_8172,In_687,In_4031);
and U8173 (N_8173,In_2640,In_1468);
and U8174 (N_8174,In_2098,In_963);
nand U8175 (N_8175,In_2834,In_2692);
nand U8176 (N_8176,In_1061,In_3677);
nor U8177 (N_8177,In_1928,In_4462);
nor U8178 (N_8178,In_293,In_4481);
nand U8179 (N_8179,In_2394,In_55);
or U8180 (N_8180,In_173,In_4002);
or U8181 (N_8181,In_1064,In_1895);
and U8182 (N_8182,In_877,In_2964);
and U8183 (N_8183,In_2096,In_2331);
xor U8184 (N_8184,In_1871,In_1599);
and U8185 (N_8185,In_4374,In_2476);
nand U8186 (N_8186,In_2292,In_3882);
nor U8187 (N_8187,In_272,In_1621);
or U8188 (N_8188,In_4510,In_4013);
nor U8189 (N_8189,In_4402,In_4393);
nand U8190 (N_8190,In_4007,In_275);
and U8191 (N_8191,In_2258,In_3322);
xnor U8192 (N_8192,In_4268,In_2812);
or U8193 (N_8193,In_1217,In_912);
and U8194 (N_8194,In_4398,In_420);
or U8195 (N_8195,In_3202,In_1899);
and U8196 (N_8196,In_3434,In_2398);
or U8197 (N_8197,In_1421,In_4248);
nand U8198 (N_8198,In_2386,In_2763);
xnor U8199 (N_8199,In_1020,In_1938);
or U8200 (N_8200,In_3612,In_322);
nor U8201 (N_8201,In_1439,In_4601);
nand U8202 (N_8202,In_2099,In_3029);
nand U8203 (N_8203,In_3891,In_3726);
nor U8204 (N_8204,In_613,In_3103);
nor U8205 (N_8205,In_180,In_4807);
nor U8206 (N_8206,In_10,In_15);
xor U8207 (N_8207,In_2648,In_3799);
xnor U8208 (N_8208,In_1394,In_3965);
xnor U8209 (N_8209,In_460,In_3117);
nand U8210 (N_8210,In_3888,In_2914);
xnor U8211 (N_8211,In_1563,In_512);
nand U8212 (N_8212,In_4093,In_3673);
and U8213 (N_8213,In_3052,In_1366);
xor U8214 (N_8214,In_976,In_3577);
and U8215 (N_8215,In_862,In_2927);
nor U8216 (N_8216,In_4496,In_2390);
nor U8217 (N_8217,In_2612,In_1028);
and U8218 (N_8218,In_1576,In_854);
and U8219 (N_8219,In_2854,In_112);
nor U8220 (N_8220,In_4641,In_1999);
and U8221 (N_8221,In_1222,In_3073);
and U8222 (N_8222,In_1880,In_494);
xor U8223 (N_8223,In_4069,In_1178);
or U8224 (N_8224,In_3614,In_3469);
and U8225 (N_8225,In_3363,In_2755);
nor U8226 (N_8226,In_3511,In_2620);
xnor U8227 (N_8227,In_3198,In_3292);
and U8228 (N_8228,In_2434,In_1257);
or U8229 (N_8229,In_2789,In_2401);
and U8230 (N_8230,In_3860,In_3017);
and U8231 (N_8231,In_3692,In_3909);
xnor U8232 (N_8232,In_2227,In_4699);
or U8233 (N_8233,In_535,In_618);
nand U8234 (N_8234,In_61,In_664);
xnor U8235 (N_8235,In_4395,In_1469);
and U8236 (N_8236,In_1221,In_4101);
xnor U8237 (N_8237,In_883,In_29);
nand U8238 (N_8238,In_4056,In_310);
or U8239 (N_8239,In_844,In_2893);
and U8240 (N_8240,In_3048,In_2626);
nor U8241 (N_8241,In_2461,In_2941);
or U8242 (N_8242,In_235,In_1966);
and U8243 (N_8243,In_757,In_3946);
xnor U8244 (N_8244,In_347,In_4075);
nand U8245 (N_8245,In_2554,In_513);
xor U8246 (N_8246,In_1952,In_1490);
nor U8247 (N_8247,In_2444,In_3530);
nand U8248 (N_8248,In_3537,In_2488);
and U8249 (N_8249,In_2074,In_573);
and U8250 (N_8250,In_1067,In_3517);
nor U8251 (N_8251,In_3215,In_4306);
nor U8252 (N_8252,In_1580,In_179);
or U8253 (N_8253,In_1122,In_1138);
xnor U8254 (N_8254,In_1718,In_2118);
xor U8255 (N_8255,In_2460,In_1187);
xor U8256 (N_8256,In_4372,In_387);
and U8257 (N_8257,In_491,In_4639);
xor U8258 (N_8258,In_897,In_4163);
nor U8259 (N_8259,In_4916,In_909);
nor U8260 (N_8260,In_973,In_419);
nand U8261 (N_8261,In_2776,In_4028);
and U8262 (N_8262,In_2336,In_4136);
nor U8263 (N_8263,In_2591,In_456);
or U8264 (N_8264,In_133,In_4259);
xnor U8265 (N_8265,In_262,In_4444);
or U8266 (N_8266,In_3935,In_2675);
and U8267 (N_8267,In_2337,In_4196);
xor U8268 (N_8268,In_2077,In_3876);
nand U8269 (N_8269,In_3762,In_693);
nor U8270 (N_8270,In_4386,In_4592);
nand U8271 (N_8271,In_135,In_3410);
and U8272 (N_8272,In_3227,In_1877);
xnor U8273 (N_8273,In_456,In_4082);
or U8274 (N_8274,In_4250,In_1376);
or U8275 (N_8275,In_3666,In_4878);
xor U8276 (N_8276,In_3789,In_1930);
nor U8277 (N_8277,In_2,In_1683);
and U8278 (N_8278,In_4109,In_4173);
or U8279 (N_8279,In_1148,In_384);
or U8280 (N_8280,In_2804,In_269);
xor U8281 (N_8281,In_4712,In_4358);
xor U8282 (N_8282,In_2381,In_771);
xor U8283 (N_8283,In_4816,In_3512);
xor U8284 (N_8284,In_1312,In_2529);
and U8285 (N_8285,In_4291,In_2719);
and U8286 (N_8286,In_2470,In_1808);
or U8287 (N_8287,In_97,In_657);
and U8288 (N_8288,In_755,In_4676);
nand U8289 (N_8289,In_4793,In_146);
and U8290 (N_8290,In_1644,In_2766);
nand U8291 (N_8291,In_921,In_670);
or U8292 (N_8292,In_3112,In_1174);
xnor U8293 (N_8293,In_3219,In_2038);
nor U8294 (N_8294,In_608,In_2264);
or U8295 (N_8295,In_4338,In_378);
nand U8296 (N_8296,In_2320,In_4913);
and U8297 (N_8297,In_2554,In_3482);
nand U8298 (N_8298,In_4836,In_622);
xnor U8299 (N_8299,In_4862,In_753);
nor U8300 (N_8300,In_3102,In_1419);
nor U8301 (N_8301,In_3175,In_3268);
nand U8302 (N_8302,In_4356,In_2881);
and U8303 (N_8303,In_3368,In_607);
or U8304 (N_8304,In_3383,In_3863);
or U8305 (N_8305,In_1534,In_3408);
xnor U8306 (N_8306,In_400,In_3404);
or U8307 (N_8307,In_1776,In_1010);
nand U8308 (N_8308,In_4406,In_3686);
nor U8309 (N_8309,In_4973,In_3723);
nand U8310 (N_8310,In_1690,In_4149);
or U8311 (N_8311,In_4119,In_4029);
or U8312 (N_8312,In_3733,In_4127);
and U8313 (N_8313,In_2783,In_544);
or U8314 (N_8314,In_2775,In_3484);
or U8315 (N_8315,In_701,In_3946);
nor U8316 (N_8316,In_1265,In_1008);
nand U8317 (N_8317,In_4795,In_4679);
xnor U8318 (N_8318,In_4180,In_1090);
nor U8319 (N_8319,In_3305,In_3542);
nand U8320 (N_8320,In_1294,In_2430);
nand U8321 (N_8321,In_4589,In_3544);
nand U8322 (N_8322,In_1372,In_4083);
xnor U8323 (N_8323,In_1688,In_3007);
nand U8324 (N_8324,In_4573,In_1093);
or U8325 (N_8325,In_2625,In_3102);
or U8326 (N_8326,In_3089,In_4443);
nor U8327 (N_8327,In_4474,In_3996);
nand U8328 (N_8328,In_4508,In_4340);
xnor U8329 (N_8329,In_481,In_4492);
and U8330 (N_8330,In_1070,In_492);
xor U8331 (N_8331,In_1941,In_268);
and U8332 (N_8332,In_2041,In_3840);
xor U8333 (N_8333,In_322,In_909);
nand U8334 (N_8334,In_904,In_4465);
nor U8335 (N_8335,In_1555,In_4737);
nor U8336 (N_8336,In_4489,In_199);
nand U8337 (N_8337,In_1452,In_4455);
and U8338 (N_8338,In_3778,In_4717);
nor U8339 (N_8339,In_4235,In_4907);
and U8340 (N_8340,In_4103,In_676);
and U8341 (N_8341,In_4587,In_3080);
or U8342 (N_8342,In_4477,In_2013);
xor U8343 (N_8343,In_440,In_2381);
and U8344 (N_8344,In_1509,In_982);
and U8345 (N_8345,In_1728,In_2010);
xnor U8346 (N_8346,In_288,In_4086);
nor U8347 (N_8347,In_3100,In_3025);
xor U8348 (N_8348,In_200,In_859);
nor U8349 (N_8349,In_1034,In_3035);
and U8350 (N_8350,In_2580,In_4460);
xnor U8351 (N_8351,In_2559,In_4661);
nand U8352 (N_8352,In_3600,In_4418);
or U8353 (N_8353,In_284,In_2706);
or U8354 (N_8354,In_3306,In_3055);
and U8355 (N_8355,In_2827,In_1368);
xor U8356 (N_8356,In_1140,In_4887);
nor U8357 (N_8357,In_3827,In_206);
nand U8358 (N_8358,In_3001,In_4300);
or U8359 (N_8359,In_1513,In_2432);
nor U8360 (N_8360,In_4616,In_3362);
nor U8361 (N_8361,In_3619,In_1138);
nor U8362 (N_8362,In_4117,In_2432);
or U8363 (N_8363,In_3282,In_2307);
nor U8364 (N_8364,In_2620,In_1977);
nor U8365 (N_8365,In_822,In_1439);
and U8366 (N_8366,In_2705,In_3951);
and U8367 (N_8367,In_1039,In_987);
nor U8368 (N_8368,In_2053,In_3315);
and U8369 (N_8369,In_3706,In_1575);
or U8370 (N_8370,In_4570,In_2862);
and U8371 (N_8371,In_4186,In_2991);
xor U8372 (N_8372,In_1990,In_1390);
and U8373 (N_8373,In_4072,In_3016);
xnor U8374 (N_8374,In_3634,In_2764);
xnor U8375 (N_8375,In_2861,In_4536);
nand U8376 (N_8376,In_2651,In_2980);
or U8377 (N_8377,In_2198,In_3905);
nor U8378 (N_8378,In_4287,In_3349);
nand U8379 (N_8379,In_901,In_876);
nor U8380 (N_8380,In_3836,In_3133);
and U8381 (N_8381,In_1674,In_2806);
or U8382 (N_8382,In_337,In_278);
nand U8383 (N_8383,In_2135,In_4696);
nor U8384 (N_8384,In_1669,In_4548);
nand U8385 (N_8385,In_2625,In_3662);
or U8386 (N_8386,In_380,In_1227);
or U8387 (N_8387,In_1441,In_2578);
nor U8388 (N_8388,In_1578,In_4774);
or U8389 (N_8389,In_4953,In_4335);
xor U8390 (N_8390,In_1402,In_4321);
and U8391 (N_8391,In_2388,In_2876);
nor U8392 (N_8392,In_3031,In_4457);
nand U8393 (N_8393,In_656,In_3469);
nand U8394 (N_8394,In_3315,In_2972);
or U8395 (N_8395,In_180,In_4778);
and U8396 (N_8396,In_4470,In_958);
xnor U8397 (N_8397,In_2962,In_1183);
or U8398 (N_8398,In_1604,In_4195);
or U8399 (N_8399,In_1227,In_1139);
xnor U8400 (N_8400,In_4112,In_4938);
or U8401 (N_8401,In_3699,In_3560);
nor U8402 (N_8402,In_38,In_2125);
nor U8403 (N_8403,In_1472,In_2785);
nor U8404 (N_8404,In_4668,In_196);
nand U8405 (N_8405,In_334,In_4390);
nor U8406 (N_8406,In_70,In_133);
and U8407 (N_8407,In_4726,In_511);
and U8408 (N_8408,In_1478,In_3496);
or U8409 (N_8409,In_1282,In_2503);
nand U8410 (N_8410,In_3956,In_4956);
nor U8411 (N_8411,In_2682,In_2496);
nand U8412 (N_8412,In_1835,In_4738);
or U8413 (N_8413,In_1632,In_1020);
or U8414 (N_8414,In_3773,In_2354);
nor U8415 (N_8415,In_4566,In_742);
nor U8416 (N_8416,In_1638,In_3270);
or U8417 (N_8417,In_1630,In_2740);
and U8418 (N_8418,In_942,In_3757);
and U8419 (N_8419,In_4948,In_324);
nor U8420 (N_8420,In_1763,In_2879);
or U8421 (N_8421,In_2877,In_160);
xnor U8422 (N_8422,In_1530,In_4866);
or U8423 (N_8423,In_423,In_3516);
and U8424 (N_8424,In_4744,In_594);
xor U8425 (N_8425,In_1467,In_4764);
and U8426 (N_8426,In_1020,In_3767);
and U8427 (N_8427,In_2398,In_2343);
or U8428 (N_8428,In_1296,In_1831);
nor U8429 (N_8429,In_487,In_145);
nand U8430 (N_8430,In_184,In_1520);
nor U8431 (N_8431,In_3574,In_290);
xor U8432 (N_8432,In_2698,In_4068);
xor U8433 (N_8433,In_958,In_960);
xnor U8434 (N_8434,In_1416,In_1937);
xnor U8435 (N_8435,In_2509,In_2814);
and U8436 (N_8436,In_3448,In_4867);
or U8437 (N_8437,In_51,In_1505);
nor U8438 (N_8438,In_3880,In_815);
nor U8439 (N_8439,In_868,In_2933);
nand U8440 (N_8440,In_1446,In_233);
nor U8441 (N_8441,In_4328,In_4641);
nand U8442 (N_8442,In_2320,In_2824);
nor U8443 (N_8443,In_3945,In_2436);
nand U8444 (N_8444,In_376,In_3318);
nand U8445 (N_8445,In_2710,In_1121);
and U8446 (N_8446,In_3267,In_1485);
nand U8447 (N_8447,In_3625,In_684);
and U8448 (N_8448,In_4653,In_3145);
or U8449 (N_8449,In_162,In_1501);
and U8450 (N_8450,In_4426,In_2161);
nand U8451 (N_8451,In_1895,In_4249);
or U8452 (N_8452,In_2690,In_3616);
xor U8453 (N_8453,In_4933,In_1412);
xor U8454 (N_8454,In_4431,In_4698);
xnor U8455 (N_8455,In_3241,In_2949);
nand U8456 (N_8456,In_2391,In_617);
xnor U8457 (N_8457,In_2257,In_2790);
nand U8458 (N_8458,In_3595,In_2451);
nand U8459 (N_8459,In_2008,In_4247);
xor U8460 (N_8460,In_1573,In_4793);
and U8461 (N_8461,In_1453,In_4895);
or U8462 (N_8462,In_922,In_3796);
nand U8463 (N_8463,In_2483,In_668);
xor U8464 (N_8464,In_4732,In_3775);
and U8465 (N_8465,In_4144,In_3772);
nand U8466 (N_8466,In_4830,In_1032);
nor U8467 (N_8467,In_4586,In_2191);
nand U8468 (N_8468,In_3957,In_691);
xnor U8469 (N_8469,In_521,In_623);
and U8470 (N_8470,In_3046,In_3699);
or U8471 (N_8471,In_954,In_1839);
xnor U8472 (N_8472,In_1897,In_3672);
xor U8473 (N_8473,In_4751,In_307);
nand U8474 (N_8474,In_779,In_2304);
and U8475 (N_8475,In_4580,In_2207);
nor U8476 (N_8476,In_3281,In_574);
xnor U8477 (N_8477,In_1726,In_1984);
or U8478 (N_8478,In_3178,In_4137);
and U8479 (N_8479,In_346,In_1072);
xor U8480 (N_8480,In_1605,In_3923);
nor U8481 (N_8481,In_3474,In_388);
and U8482 (N_8482,In_2361,In_1202);
or U8483 (N_8483,In_3708,In_2397);
xor U8484 (N_8484,In_4263,In_60);
nand U8485 (N_8485,In_3723,In_4391);
nand U8486 (N_8486,In_4877,In_17);
nor U8487 (N_8487,In_2364,In_4105);
xnor U8488 (N_8488,In_3787,In_1047);
xor U8489 (N_8489,In_2605,In_2525);
nand U8490 (N_8490,In_468,In_1813);
nor U8491 (N_8491,In_1163,In_3404);
xnor U8492 (N_8492,In_4235,In_3922);
xor U8493 (N_8493,In_1365,In_4823);
nor U8494 (N_8494,In_3028,In_1756);
nand U8495 (N_8495,In_1533,In_58);
nand U8496 (N_8496,In_2173,In_2947);
and U8497 (N_8497,In_2709,In_2745);
nand U8498 (N_8498,In_4465,In_2217);
xnor U8499 (N_8499,In_1226,In_4657);
nand U8500 (N_8500,In_1112,In_859);
nand U8501 (N_8501,In_2784,In_3341);
nor U8502 (N_8502,In_4833,In_938);
nor U8503 (N_8503,In_3759,In_1897);
and U8504 (N_8504,In_2826,In_4424);
nand U8505 (N_8505,In_552,In_3711);
xor U8506 (N_8506,In_2238,In_4617);
and U8507 (N_8507,In_2117,In_4431);
and U8508 (N_8508,In_3136,In_378);
nor U8509 (N_8509,In_1257,In_4041);
xnor U8510 (N_8510,In_4137,In_655);
xnor U8511 (N_8511,In_3591,In_1228);
or U8512 (N_8512,In_3685,In_3099);
nor U8513 (N_8513,In_1999,In_4438);
and U8514 (N_8514,In_3365,In_926);
xor U8515 (N_8515,In_4422,In_1988);
or U8516 (N_8516,In_4820,In_3568);
and U8517 (N_8517,In_4748,In_3165);
nor U8518 (N_8518,In_76,In_2578);
and U8519 (N_8519,In_3624,In_4765);
and U8520 (N_8520,In_3021,In_4766);
or U8521 (N_8521,In_1756,In_2495);
nand U8522 (N_8522,In_576,In_787);
nor U8523 (N_8523,In_2735,In_1573);
nor U8524 (N_8524,In_2460,In_309);
or U8525 (N_8525,In_2624,In_3588);
and U8526 (N_8526,In_1665,In_2978);
xnor U8527 (N_8527,In_858,In_1446);
and U8528 (N_8528,In_4842,In_3712);
nor U8529 (N_8529,In_4333,In_3327);
and U8530 (N_8530,In_2888,In_3136);
or U8531 (N_8531,In_1064,In_2484);
nor U8532 (N_8532,In_1717,In_3113);
xnor U8533 (N_8533,In_690,In_4913);
and U8534 (N_8534,In_368,In_4625);
nand U8535 (N_8535,In_4511,In_4124);
nor U8536 (N_8536,In_84,In_413);
nand U8537 (N_8537,In_4476,In_820);
and U8538 (N_8538,In_373,In_3000);
and U8539 (N_8539,In_4508,In_545);
xor U8540 (N_8540,In_2087,In_773);
or U8541 (N_8541,In_2392,In_1473);
or U8542 (N_8542,In_3507,In_1998);
and U8543 (N_8543,In_985,In_831);
and U8544 (N_8544,In_923,In_1174);
nor U8545 (N_8545,In_1964,In_82);
nor U8546 (N_8546,In_1569,In_1481);
and U8547 (N_8547,In_423,In_3722);
xnor U8548 (N_8548,In_26,In_452);
or U8549 (N_8549,In_3064,In_1398);
nor U8550 (N_8550,In_4436,In_2586);
nand U8551 (N_8551,In_3702,In_2394);
nand U8552 (N_8552,In_4856,In_1376);
nand U8553 (N_8553,In_3492,In_2704);
nor U8554 (N_8554,In_3391,In_1023);
and U8555 (N_8555,In_1846,In_4929);
or U8556 (N_8556,In_4895,In_2521);
or U8557 (N_8557,In_901,In_2064);
and U8558 (N_8558,In_709,In_2867);
or U8559 (N_8559,In_1774,In_2584);
or U8560 (N_8560,In_2490,In_1708);
nor U8561 (N_8561,In_3482,In_798);
xnor U8562 (N_8562,In_474,In_4673);
nor U8563 (N_8563,In_4782,In_779);
xor U8564 (N_8564,In_1807,In_4654);
nand U8565 (N_8565,In_3234,In_2199);
or U8566 (N_8566,In_431,In_4511);
and U8567 (N_8567,In_4387,In_334);
nand U8568 (N_8568,In_2353,In_1705);
nand U8569 (N_8569,In_139,In_792);
or U8570 (N_8570,In_2528,In_3855);
xnor U8571 (N_8571,In_4745,In_1090);
nand U8572 (N_8572,In_1010,In_263);
or U8573 (N_8573,In_4848,In_4729);
xor U8574 (N_8574,In_173,In_2773);
nor U8575 (N_8575,In_4617,In_4089);
or U8576 (N_8576,In_1218,In_2700);
xnor U8577 (N_8577,In_720,In_4569);
xor U8578 (N_8578,In_4141,In_4156);
and U8579 (N_8579,In_3073,In_3203);
nand U8580 (N_8580,In_1261,In_1701);
or U8581 (N_8581,In_1023,In_221);
xnor U8582 (N_8582,In_640,In_782);
and U8583 (N_8583,In_2669,In_3502);
nand U8584 (N_8584,In_1636,In_1294);
and U8585 (N_8585,In_805,In_1289);
and U8586 (N_8586,In_3873,In_205);
xnor U8587 (N_8587,In_1378,In_3310);
and U8588 (N_8588,In_2783,In_3853);
nor U8589 (N_8589,In_2299,In_1851);
xnor U8590 (N_8590,In_621,In_2236);
nand U8591 (N_8591,In_1989,In_1208);
nand U8592 (N_8592,In_2151,In_3125);
xor U8593 (N_8593,In_4532,In_799);
or U8594 (N_8594,In_2338,In_2977);
and U8595 (N_8595,In_4354,In_3175);
nand U8596 (N_8596,In_3884,In_52);
xor U8597 (N_8597,In_1461,In_3410);
xor U8598 (N_8598,In_3650,In_3282);
and U8599 (N_8599,In_912,In_2614);
or U8600 (N_8600,In_1787,In_3168);
nand U8601 (N_8601,In_2752,In_1072);
xnor U8602 (N_8602,In_2652,In_1393);
or U8603 (N_8603,In_4253,In_3353);
xor U8604 (N_8604,In_4959,In_3128);
and U8605 (N_8605,In_1476,In_4212);
nor U8606 (N_8606,In_1202,In_3233);
nand U8607 (N_8607,In_2602,In_1685);
xnor U8608 (N_8608,In_4455,In_4101);
xor U8609 (N_8609,In_711,In_3767);
xnor U8610 (N_8610,In_3121,In_1199);
nor U8611 (N_8611,In_2592,In_2515);
or U8612 (N_8612,In_4041,In_3575);
nor U8613 (N_8613,In_4619,In_334);
nand U8614 (N_8614,In_78,In_221);
or U8615 (N_8615,In_1498,In_2332);
nor U8616 (N_8616,In_1575,In_4515);
or U8617 (N_8617,In_2308,In_2496);
or U8618 (N_8618,In_705,In_4956);
xnor U8619 (N_8619,In_318,In_1347);
and U8620 (N_8620,In_1717,In_1968);
nor U8621 (N_8621,In_3698,In_2974);
and U8622 (N_8622,In_3019,In_3737);
xor U8623 (N_8623,In_120,In_4325);
or U8624 (N_8624,In_4049,In_564);
or U8625 (N_8625,In_564,In_3224);
nor U8626 (N_8626,In_92,In_1926);
nand U8627 (N_8627,In_4227,In_1745);
or U8628 (N_8628,In_1330,In_510);
nand U8629 (N_8629,In_2775,In_2559);
and U8630 (N_8630,In_1481,In_3729);
nor U8631 (N_8631,In_4439,In_594);
or U8632 (N_8632,In_1264,In_1814);
and U8633 (N_8633,In_300,In_563);
nor U8634 (N_8634,In_4892,In_768);
xor U8635 (N_8635,In_3386,In_3185);
and U8636 (N_8636,In_3827,In_173);
nand U8637 (N_8637,In_4681,In_3164);
or U8638 (N_8638,In_2909,In_901);
and U8639 (N_8639,In_2307,In_4253);
nand U8640 (N_8640,In_1503,In_3703);
nand U8641 (N_8641,In_532,In_649);
or U8642 (N_8642,In_2807,In_3605);
nand U8643 (N_8643,In_915,In_2100);
or U8644 (N_8644,In_4558,In_1698);
nand U8645 (N_8645,In_3446,In_836);
or U8646 (N_8646,In_3225,In_266);
and U8647 (N_8647,In_2039,In_1541);
nor U8648 (N_8648,In_3329,In_3825);
and U8649 (N_8649,In_4774,In_59);
nor U8650 (N_8650,In_2509,In_2387);
and U8651 (N_8651,In_1244,In_2152);
or U8652 (N_8652,In_4068,In_3605);
nor U8653 (N_8653,In_2884,In_4750);
or U8654 (N_8654,In_1135,In_3489);
nand U8655 (N_8655,In_278,In_2304);
and U8656 (N_8656,In_4283,In_1586);
nor U8657 (N_8657,In_3131,In_1696);
xor U8658 (N_8658,In_1348,In_4900);
nor U8659 (N_8659,In_3832,In_3758);
and U8660 (N_8660,In_4467,In_305);
nor U8661 (N_8661,In_1762,In_1093);
or U8662 (N_8662,In_3606,In_3047);
nor U8663 (N_8663,In_1695,In_43);
nand U8664 (N_8664,In_2405,In_4347);
and U8665 (N_8665,In_2954,In_612);
nor U8666 (N_8666,In_3057,In_225);
or U8667 (N_8667,In_1119,In_4504);
and U8668 (N_8668,In_1507,In_298);
xor U8669 (N_8669,In_3864,In_1451);
and U8670 (N_8670,In_817,In_3026);
xnor U8671 (N_8671,In_2376,In_1239);
xor U8672 (N_8672,In_3238,In_1548);
nand U8673 (N_8673,In_1907,In_1964);
and U8674 (N_8674,In_284,In_1191);
xnor U8675 (N_8675,In_623,In_901);
nor U8676 (N_8676,In_3260,In_2385);
or U8677 (N_8677,In_1585,In_3938);
nor U8678 (N_8678,In_4287,In_1761);
and U8679 (N_8679,In_4756,In_3218);
xnor U8680 (N_8680,In_1633,In_2679);
xnor U8681 (N_8681,In_3431,In_2317);
xnor U8682 (N_8682,In_1630,In_3831);
or U8683 (N_8683,In_602,In_2532);
xnor U8684 (N_8684,In_4293,In_1964);
and U8685 (N_8685,In_2669,In_60);
nor U8686 (N_8686,In_3902,In_4388);
and U8687 (N_8687,In_3055,In_1576);
or U8688 (N_8688,In_2615,In_1255);
nor U8689 (N_8689,In_2195,In_494);
nor U8690 (N_8690,In_1077,In_1610);
or U8691 (N_8691,In_1656,In_2585);
nand U8692 (N_8692,In_3566,In_3872);
xnor U8693 (N_8693,In_4963,In_3950);
and U8694 (N_8694,In_4892,In_3430);
or U8695 (N_8695,In_4314,In_2869);
or U8696 (N_8696,In_1766,In_575);
or U8697 (N_8697,In_623,In_3569);
and U8698 (N_8698,In_4117,In_4586);
nor U8699 (N_8699,In_2987,In_205);
nand U8700 (N_8700,In_4576,In_2682);
nor U8701 (N_8701,In_4104,In_259);
xnor U8702 (N_8702,In_4552,In_3502);
and U8703 (N_8703,In_2669,In_2419);
nor U8704 (N_8704,In_1356,In_940);
xnor U8705 (N_8705,In_139,In_290);
nor U8706 (N_8706,In_2684,In_2002);
nand U8707 (N_8707,In_3276,In_714);
and U8708 (N_8708,In_3253,In_4066);
nand U8709 (N_8709,In_938,In_2763);
or U8710 (N_8710,In_2343,In_1677);
and U8711 (N_8711,In_1231,In_4975);
nor U8712 (N_8712,In_473,In_3716);
nand U8713 (N_8713,In_4742,In_2471);
xor U8714 (N_8714,In_4268,In_215);
xor U8715 (N_8715,In_4097,In_3801);
nand U8716 (N_8716,In_3453,In_273);
or U8717 (N_8717,In_2071,In_737);
nor U8718 (N_8718,In_1309,In_4629);
nor U8719 (N_8719,In_1978,In_4058);
and U8720 (N_8720,In_2185,In_862);
and U8721 (N_8721,In_3506,In_3762);
or U8722 (N_8722,In_4245,In_1588);
and U8723 (N_8723,In_2899,In_2835);
and U8724 (N_8724,In_1597,In_3420);
nor U8725 (N_8725,In_288,In_4672);
or U8726 (N_8726,In_405,In_20);
and U8727 (N_8727,In_2199,In_3477);
xnor U8728 (N_8728,In_1920,In_3705);
nor U8729 (N_8729,In_2142,In_6);
nor U8730 (N_8730,In_4457,In_2331);
and U8731 (N_8731,In_1729,In_1933);
nor U8732 (N_8732,In_1453,In_2300);
and U8733 (N_8733,In_2618,In_1792);
xor U8734 (N_8734,In_970,In_1269);
or U8735 (N_8735,In_476,In_1154);
xnor U8736 (N_8736,In_1091,In_3834);
nor U8737 (N_8737,In_1829,In_3367);
and U8738 (N_8738,In_4314,In_1732);
nor U8739 (N_8739,In_4411,In_985);
or U8740 (N_8740,In_4485,In_722);
or U8741 (N_8741,In_3779,In_526);
and U8742 (N_8742,In_1857,In_81);
and U8743 (N_8743,In_4127,In_1244);
xor U8744 (N_8744,In_1897,In_801);
nor U8745 (N_8745,In_1844,In_2923);
or U8746 (N_8746,In_2300,In_1112);
and U8747 (N_8747,In_1774,In_419);
xnor U8748 (N_8748,In_381,In_3172);
and U8749 (N_8749,In_2868,In_4152);
nand U8750 (N_8750,In_517,In_4144);
nor U8751 (N_8751,In_2871,In_3573);
and U8752 (N_8752,In_1287,In_554);
xor U8753 (N_8753,In_4072,In_638);
nand U8754 (N_8754,In_2982,In_2109);
xor U8755 (N_8755,In_1504,In_4750);
nor U8756 (N_8756,In_4506,In_1047);
or U8757 (N_8757,In_4325,In_4337);
xnor U8758 (N_8758,In_3383,In_4264);
or U8759 (N_8759,In_998,In_2578);
nor U8760 (N_8760,In_2342,In_3972);
and U8761 (N_8761,In_1807,In_4598);
nor U8762 (N_8762,In_2617,In_1133);
xor U8763 (N_8763,In_1422,In_4068);
nor U8764 (N_8764,In_4584,In_2611);
or U8765 (N_8765,In_1995,In_1166);
and U8766 (N_8766,In_4464,In_4173);
nand U8767 (N_8767,In_3691,In_1322);
or U8768 (N_8768,In_984,In_312);
and U8769 (N_8769,In_2173,In_1708);
or U8770 (N_8770,In_1072,In_2225);
xor U8771 (N_8771,In_4418,In_335);
nand U8772 (N_8772,In_1384,In_2006);
nand U8773 (N_8773,In_3852,In_1055);
or U8774 (N_8774,In_3602,In_2435);
or U8775 (N_8775,In_4979,In_4458);
nor U8776 (N_8776,In_1865,In_3282);
xnor U8777 (N_8777,In_3832,In_4717);
nand U8778 (N_8778,In_2703,In_1601);
or U8779 (N_8779,In_4280,In_610);
nand U8780 (N_8780,In_3986,In_2881);
or U8781 (N_8781,In_1483,In_1413);
or U8782 (N_8782,In_352,In_679);
and U8783 (N_8783,In_3994,In_4613);
nor U8784 (N_8784,In_4250,In_4307);
nor U8785 (N_8785,In_3373,In_750);
nor U8786 (N_8786,In_3146,In_2194);
nor U8787 (N_8787,In_4085,In_2574);
or U8788 (N_8788,In_2240,In_2298);
and U8789 (N_8789,In_2995,In_1528);
and U8790 (N_8790,In_467,In_4148);
xnor U8791 (N_8791,In_149,In_1088);
and U8792 (N_8792,In_3899,In_4506);
xor U8793 (N_8793,In_2859,In_4263);
and U8794 (N_8794,In_2553,In_2272);
xor U8795 (N_8795,In_4597,In_2655);
and U8796 (N_8796,In_1317,In_3289);
nor U8797 (N_8797,In_4287,In_516);
or U8798 (N_8798,In_853,In_3533);
xor U8799 (N_8799,In_2287,In_1289);
nor U8800 (N_8800,In_3578,In_4954);
nand U8801 (N_8801,In_2899,In_2174);
xnor U8802 (N_8802,In_1195,In_2819);
xor U8803 (N_8803,In_1710,In_1311);
and U8804 (N_8804,In_2073,In_3148);
or U8805 (N_8805,In_4398,In_4900);
nor U8806 (N_8806,In_4732,In_3075);
xor U8807 (N_8807,In_1519,In_1651);
or U8808 (N_8808,In_3294,In_2671);
xor U8809 (N_8809,In_958,In_1712);
or U8810 (N_8810,In_4093,In_2348);
or U8811 (N_8811,In_2495,In_267);
or U8812 (N_8812,In_942,In_4209);
nor U8813 (N_8813,In_1289,In_341);
or U8814 (N_8814,In_3281,In_4284);
or U8815 (N_8815,In_2913,In_4695);
nor U8816 (N_8816,In_2951,In_1564);
or U8817 (N_8817,In_1398,In_2680);
xor U8818 (N_8818,In_4038,In_2478);
nand U8819 (N_8819,In_4663,In_3232);
nand U8820 (N_8820,In_4313,In_45);
xor U8821 (N_8821,In_3653,In_18);
or U8822 (N_8822,In_2549,In_4034);
nor U8823 (N_8823,In_2154,In_3875);
and U8824 (N_8824,In_4004,In_1739);
nor U8825 (N_8825,In_2497,In_3709);
nand U8826 (N_8826,In_1575,In_1870);
nor U8827 (N_8827,In_4497,In_1976);
nand U8828 (N_8828,In_4397,In_3675);
and U8829 (N_8829,In_1376,In_3308);
nand U8830 (N_8830,In_414,In_3497);
nand U8831 (N_8831,In_838,In_4586);
or U8832 (N_8832,In_3915,In_4063);
xor U8833 (N_8833,In_1917,In_3933);
or U8834 (N_8834,In_4003,In_2835);
and U8835 (N_8835,In_2579,In_3873);
nor U8836 (N_8836,In_2747,In_1870);
xor U8837 (N_8837,In_2836,In_4879);
xor U8838 (N_8838,In_2221,In_27);
nor U8839 (N_8839,In_3150,In_431);
or U8840 (N_8840,In_3546,In_2805);
and U8841 (N_8841,In_865,In_4532);
nand U8842 (N_8842,In_3743,In_2724);
and U8843 (N_8843,In_4908,In_4410);
or U8844 (N_8844,In_3203,In_4731);
xnor U8845 (N_8845,In_2682,In_456);
nor U8846 (N_8846,In_1625,In_2756);
nor U8847 (N_8847,In_2577,In_1008);
xor U8848 (N_8848,In_4128,In_3088);
nor U8849 (N_8849,In_563,In_1394);
nand U8850 (N_8850,In_4789,In_376);
xnor U8851 (N_8851,In_4297,In_4170);
nand U8852 (N_8852,In_3165,In_4275);
nor U8853 (N_8853,In_3396,In_4226);
nor U8854 (N_8854,In_1397,In_1288);
nor U8855 (N_8855,In_1048,In_2355);
nor U8856 (N_8856,In_4024,In_2642);
and U8857 (N_8857,In_1115,In_2440);
nand U8858 (N_8858,In_1596,In_3428);
or U8859 (N_8859,In_2461,In_3290);
nand U8860 (N_8860,In_2852,In_2024);
or U8861 (N_8861,In_3338,In_1411);
or U8862 (N_8862,In_3627,In_1932);
xnor U8863 (N_8863,In_3448,In_1989);
or U8864 (N_8864,In_2540,In_4276);
nor U8865 (N_8865,In_2125,In_4889);
or U8866 (N_8866,In_2987,In_2999);
nand U8867 (N_8867,In_5,In_1741);
nor U8868 (N_8868,In_436,In_2421);
xnor U8869 (N_8869,In_2438,In_4036);
and U8870 (N_8870,In_957,In_3200);
xnor U8871 (N_8871,In_738,In_524);
and U8872 (N_8872,In_2894,In_3648);
nor U8873 (N_8873,In_1255,In_1594);
xor U8874 (N_8874,In_2362,In_4247);
or U8875 (N_8875,In_2283,In_4362);
xnor U8876 (N_8876,In_931,In_2082);
nor U8877 (N_8877,In_3523,In_1866);
nor U8878 (N_8878,In_2774,In_1662);
or U8879 (N_8879,In_3359,In_1286);
xnor U8880 (N_8880,In_1837,In_935);
or U8881 (N_8881,In_1466,In_1980);
and U8882 (N_8882,In_160,In_1670);
nand U8883 (N_8883,In_4194,In_753);
and U8884 (N_8884,In_496,In_105);
nor U8885 (N_8885,In_2953,In_2524);
nand U8886 (N_8886,In_33,In_1662);
and U8887 (N_8887,In_2731,In_2847);
xor U8888 (N_8888,In_3901,In_186);
or U8889 (N_8889,In_4767,In_1231);
nand U8890 (N_8890,In_4070,In_4907);
nand U8891 (N_8891,In_754,In_1184);
or U8892 (N_8892,In_96,In_31);
nand U8893 (N_8893,In_3507,In_3849);
nor U8894 (N_8894,In_3076,In_2286);
nor U8895 (N_8895,In_3223,In_4741);
nand U8896 (N_8896,In_4352,In_2992);
or U8897 (N_8897,In_1730,In_2617);
nor U8898 (N_8898,In_4398,In_4185);
nand U8899 (N_8899,In_1715,In_4350);
nand U8900 (N_8900,In_496,In_2614);
nand U8901 (N_8901,In_2292,In_525);
xor U8902 (N_8902,In_689,In_2599);
nand U8903 (N_8903,In_3804,In_3298);
nand U8904 (N_8904,In_4566,In_4273);
or U8905 (N_8905,In_2072,In_4106);
xnor U8906 (N_8906,In_1785,In_487);
nor U8907 (N_8907,In_2420,In_4657);
nand U8908 (N_8908,In_4132,In_1021);
nor U8909 (N_8909,In_1955,In_1791);
or U8910 (N_8910,In_2342,In_4448);
or U8911 (N_8911,In_2102,In_2340);
nor U8912 (N_8912,In_3559,In_909);
or U8913 (N_8913,In_4560,In_2444);
or U8914 (N_8914,In_2245,In_2518);
nand U8915 (N_8915,In_94,In_2153);
nor U8916 (N_8916,In_1927,In_4519);
xnor U8917 (N_8917,In_4010,In_4468);
nor U8918 (N_8918,In_2275,In_4976);
nand U8919 (N_8919,In_3607,In_1245);
and U8920 (N_8920,In_1597,In_1478);
nor U8921 (N_8921,In_673,In_3020);
or U8922 (N_8922,In_2634,In_1044);
nor U8923 (N_8923,In_1254,In_2834);
and U8924 (N_8924,In_3177,In_3437);
and U8925 (N_8925,In_1430,In_1698);
nand U8926 (N_8926,In_4837,In_2428);
nor U8927 (N_8927,In_3238,In_3126);
nand U8928 (N_8928,In_694,In_1388);
and U8929 (N_8929,In_2129,In_3335);
nor U8930 (N_8930,In_4752,In_3063);
and U8931 (N_8931,In_1750,In_3435);
nand U8932 (N_8932,In_2275,In_1953);
or U8933 (N_8933,In_1094,In_3055);
and U8934 (N_8934,In_4698,In_2609);
and U8935 (N_8935,In_922,In_4039);
or U8936 (N_8936,In_2703,In_2383);
or U8937 (N_8937,In_1319,In_793);
nand U8938 (N_8938,In_2003,In_87);
and U8939 (N_8939,In_1474,In_1613);
or U8940 (N_8940,In_4718,In_483);
or U8941 (N_8941,In_4282,In_66);
or U8942 (N_8942,In_3934,In_3336);
nand U8943 (N_8943,In_4327,In_1865);
nand U8944 (N_8944,In_2488,In_3317);
xnor U8945 (N_8945,In_1367,In_4469);
xnor U8946 (N_8946,In_2594,In_140);
xnor U8947 (N_8947,In_2620,In_1001);
xor U8948 (N_8948,In_1934,In_151);
and U8949 (N_8949,In_2012,In_761);
nand U8950 (N_8950,In_3477,In_945);
xnor U8951 (N_8951,In_705,In_2552);
nand U8952 (N_8952,In_3481,In_2884);
nand U8953 (N_8953,In_3412,In_3474);
nand U8954 (N_8954,In_853,In_2878);
xnor U8955 (N_8955,In_3150,In_3295);
xnor U8956 (N_8956,In_2776,In_3311);
or U8957 (N_8957,In_2772,In_2696);
nor U8958 (N_8958,In_721,In_557);
nor U8959 (N_8959,In_1878,In_2100);
nor U8960 (N_8960,In_4125,In_319);
and U8961 (N_8961,In_2535,In_1309);
and U8962 (N_8962,In_3266,In_4546);
and U8963 (N_8963,In_3764,In_2044);
nand U8964 (N_8964,In_363,In_1348);
or U8965 (N_8965,In_578,In_4419);
and U8966 (N_8966,In_1621,In_546);
or U8967 (N_8967,In_4690,In_5);
and U8968 (N_8968,In_4161,In_3920);
and U8969 (N_8969,In_1222,In_2866);
or U8970 (N_8970,In_2321,In_3089);
and U8971 (N_8971,In_3097,In_3455);
xor U8972 (N_8972,In_1039,In_4699);
and U8973 (N_8973,In_1359,In_4937);
and U8974 (N_8974,In_1190,In_3953);
or U8975 (N_8975,In_3471,In_807);
nand U8976 (N_8976,In_929,In_2255);
and U8977 (N_8977,In_2476,In_1000);
or U8978 (N_8978,In_544,In_3310);
nor U8979 (N_8979,In_695,In_3949);
and U8980 (N_8980,In_4557,In_1943);
and U8981 (N_8981,In_448,In_3247);
nor U8982 (N_8982,In_384,In_3507);
xnor U8983 (N_8983,In_978,In_3446);
nand U8984 (N_8984,In_1297,In_2747);
and U8985 (N_8985,In_353,In_4468);
and U8986 (N_8986,In_1979,In_910);
and U8987 (N_8987,In_2201,In_643);
nand U8988 (N_8988,In_1329,In_1091);
and U8989 (N_8989,In_3298,In_2106);
nand U8990 (N_8990,In_3091,In_216);
and U8991 (N_8991,In_135,In_3489);
xor U8992 (N_8992,In_1238,In_1381);
xor U8993 (N_8993,In_770,In_1604);
nor U8994 (N_8994,In_136,In_3114);
nor U8995 (N_8995,In_4131,In_1869);
xnor U8996 (N_8996,In_3226,In_4228);
and U8997 (N_8997,In_1131,In_3152);
nand U8998 (N_8998,In_1637,In_1359);
xor U8999 (N_8999,In_2746,In_1750);
nand U9000 (N_9000,In_3724,In_2717);
xnor U9001 (N_9001,In_3736,In_4124);
nand U9002 (N_9002,In_3616,In_1521);
or U9003 (N_9003,In_4063,In_1799);
or U9004 (N_9004,In_910,In_4555);
and U9005 (N_9005,In_4466,In_4177);
nand U9006 (N_9006,In_1711,In_2882);
or U9007 (N_9007,In_1746,In_1010);
xnor U9008 (N_9008,In_3713,In_872);
nor U9009 (N_9009,In_2631,In_1461);
nand U9010 (N_9010,In_3406,In_4855);
nor U9011 (N_9011,In_1317,In_7);
nor U9012 (N_9012,In_4889,In_3718);
or U9013 (N_9013,In_2047,In_122);
xor U9014 (N_9014,In_3508,In_2449);
nand U9015 (N_9015,In_684,In_817);
and U9016 (N_9016,In_769,In_1345);
or U9017 (N_9017,In_3362,In_2495);
xnor U9018 (N_9018,In_1370,In_2700);
and U9019 (N_9019,In_3715,In_1147);
and U9020 (N_9020,In_100,In_3866);
nor U9021 (N_9021,In_657,In_4749);
and U9022 (N_9022,In_4498,In_4619);
nand U9023 (N_9023,In_1190,In_988);
or U9024 (N_9024,In_4946,In_2992);
nor U9025 (N_9025,In_3307,In_3559);
and U9026 (N_9026,In_3853,In_2193);
nand U9027 (N_9027,In_3052,In_3295);
xnor U9028 (N_9028,In_4146,In_149);
nand U9029 (N_9029,In_1956,In_536);
or U9030 (N_9030,In_64,In_978);
or U9031 (N_9031,In_3267,In_2038);
nand U9032 (N_9032,In_2975,In_3523);
or U9033 (N_9033,In_424,In_263);
xor U9034 (N_9034,In_403,In_1190);
nor U9035 (N_9035,In_1533,In_2663);
nand U9036 (N_9036,In_635,In_150);
or U9037 (N_9037,In_1265,In_4970);
or U9038 (N_9038,In_1680,In_3088);
and U9039 (N_9039,In_3598,In_1732);
nand U9040 (N_9040,In_1583,In_4538);
and U9041 (N_9041,In_3577,In_4446);
xor U9042 (N_9042,In_4933,In_1647);
nor U9043 (N_9043,In_836,In_1695);
or U9044 (N_9044,In_2081,In_4616);
or U9045 (N_9045,In_3449,In_1593);
and U9046 (N_9046,In_2093,In_1775);
nor U9047 (N_9047,In_3536,In_1706);
and U9048 (N_9048,In_121,In_3210);
nand U9049 (N_9049,In_956,In_3023);
or U9050 (N_9050,In_2473,In_1933);
xnor U9051 (N_9051,In_2508,In_4956);
xor U9052 (N_9052,In_174,In_1049);
and U9053 (N_9053,In_361,In_1351);
nor U9054 (N_9054,In_2006,In_4268);
nand U9055 (N_9055,In_731,In_4555);
and U9056 (N_9056,In_3004,In_4680);
and U9057 (N_9057,In_4801,In_4836);
or U9058 (N_9058,In_1433,In_1527);
nor U9059 (N_9059,In_245,In_3711);
nor U9060 (N_9060,In_1963,In_4493);
nor U9061 (N_9061,In_2558,In_1294);
nand U9062 (N_9062,In_3971,In_4852);
nand U9063 (N_9063,In_3109,In_626);
and U9064 (N_9064,In_3417,In_3732);
nand U9065 (N_9065,In_1793,In_3215);
or U9066 (N_9066,In_3642,In_669);
nand U9067 (N_9067,In_1384,In_1829);
or U9068 (N_9068,In_1988,In_294);
and U9069 (N_9069,In_1030,In_3155);
nor U9070 (N_9070,In_1317,In_1637);
and U9071 (N_9071,In_2030,In_131);
xnor U9072 (N_9072,In_2478,In_1608);
nor U9073 (N_9073,In_2318,In_3691);
or U9074 (N_9074,In_1817,In_232);
and U9075 (N_9075,In_1112,In_2887);
or U9076 (N_9076,In_150,In_4509);
and U9077 (N_9077,In_2855,In_4715);
nor U9078 (N_9078,In_1771,In_299);
nor U9079 (N_9079,In_4902,In_469);
or U9080 (N_9080,In_3263,In_515);
nor U9081 (N_9081,In_3321,In_1114);
nor U9082 (N_9082,In_1107,In_2141);
nor U9083 (N_9083,In_3099,In_3871);
xnor U9084 (N_9084,In_1182,In_1948);
and U9085 (N_9085,In_2070,In_1523);
nand U9086 (N_9086,In_2307,In_454);
or U9087 (N_9087,In_1377,In_4911);
nor U9088 (N_9088,In_108,In_3587);
xnor U9089 (N_9089,In_3224,In_3083);
xor U9090 (N_9090,In_1640,In_4828);
nand U9091 (N_9091,In_4474,In_3957);
and U9092 (N_9092,In_3520,In_2652);
nand U9093 (N_9093,In_4957,In_2799);
or U9094 (N_9094,In_3810,In_4860);
and U9095 (N_9095,In_1416,In_3051);
nor U9096 (N_9096,In_1155,In_1284);
nor U9097 (N_9097,In_2347,In_2608);
nor U9098 (N_9098,In_1186,In_3323);
xor U9099 (N_9099,In_3825,In_3416);
and U9100 (N_9100,In_37,In_2400);
nand U9101 (N_9101,In_3431,In_3943);
nor U9102 (N_9102,In_1800,In_2436);
or U9103 (N_9103,In_145,In_3016);
nor U9104 (N_9104,In_779,In_3761);
xor U9105 (N_9105,In_1079,In_3052);
and U9106 (N_9106,In_1811,In_3784);
xor U9107 (N_9107,In_3530,In_24);
nand U9108 (N_9108,In_1092,In_4520);
and U9109 (N_9109,In_3595,In_3855);
or U9110 (N_9110,In_478,In_2081);
nor U9111 (N_9111,In_660,In_154);
nor U9112 (N_9112,In_607,In_787);
nor U9113 (N_9113,In_937,In_3133);
nor U9114 (N_9114,In_1490,In_1357);
nor U9115 (N_9115,In_1004,In_1530);
xor U9116 (N_9116,In_1277,In_1264);
or U9117 (N_9117,In_1382,In_3155);
or U9118 (N_9118,In_4022,In_3228);
nor U9119 (N_9119,In_688,In_1527);
or U9120 (N_9120,In_60,In_3004);
nor U9121 (N_9121,In_3138,In_4087);
nor U9122 (N_9122,In_1792,In_1415);
and U9123 (N_9123,In_1353,In_473);
nand U9124 (N_9124,In_3680,In_4647);
nand U9125 (N_9125,In_32,In_951);
or U9126 (N_9126,In_4004,In_873);
and U9127 (N_9127,In_2978,In_2388);
nor U9128 (N_9128,In_2845,In_1740);
nand U9129 (N_9129,In_519,In_2586);
or U9130 (N_9130,In_734,In_3328);
nand U9131 (N_9131,In_3269,In_807);
or U9132 (N_9132,In_3950,In_353);
nor U9133 (N_9133,In_4482,In_1488);
xnor U9134 (N_9134,In_3399,In_2082);
nor U9135 (N_9135,In_4133,In_3376);
or U9136 (N_9136,In_402,In_2662);
xnor U9137 (N_9137,In_1477,In_4563);
xnor U9138 (N_9138,In_3172,In_1828);
and U9139 (N_9139,In_236,In_1418);
xor U9140 (N_9140,In_1307,In_1734);
nor U9141 (N_9141,In_3028,In_2417);
and U9142 (N_9142,In_3126,In_2981);
nand U9143 (N_9143,In_468,In_4595);
nand U9144 (N_9144,In_3138,In_1511);
xor U9145 (N_9145,In_3831,In_196);
or U9146 (N_9146,In_4145,In_1868);
and U9147 (N_9147,In_897,In_4259);
and U9148 (N_9148,In_851,In_50);
nor U9149 (N_9149,In_4646,In_254);
xnor U9150 (N_9150,In_923,In_2270);
nand U9151 (N_9151,In_1684,In_4422);
or U9152 (N_9152,In_4668,In_2616);
and U9153 (N_9153,In_4247,In_4688);
nor U9154 (N_9154,In_65,In_2979);
and U9155 (N_9155,In_24,In_1529);
and U9156 (N_9156,In_2467,In_4957);
nor U9157 (N_9157,In_2702,In_769);
nor U9158 (N_9158,In_4428,In_4598);
and U9159 (N_9159,In_2027,In_3285);
nor U9160 (N_9160,In_414,In_3158);
and U9161 (N_9161,In_4883,In_3537);
nand U9162 (N_9162,In_898,In_3590);
or U9163 (N_9163,In_3741,In_3867);
or U9164 (N_9164,In_4145,In_4376);
or U9165 (N_9165,In_4032,In_4069);
or U9166 (N_9166,In_903,In_1848);
nor U9167 (N_9167,In_0,In_2561);
nor U9168 (N_9168,In_121,In_536);
nor U9169 (N_9169,In_3668,In_3604);
or U9170 (N_9170,In_3811,In_4407);
nand U9171 (N_9171,In_1259,In_2380);
nand U9172 (N_9172,In_2112,In_2104);
and U9173 (N_9173,In_3554,In_227);
xor U9174 (N_9174,In_748,In_3008);
or U9175 (N_9175,In_4155,In_361);
nor U9176 (N_9176,In_309,In_1133);
nor U9177 (N_9177,In_4764,In_3210);
and U9178 (N_9178,In_3991,In_4975);
and U9179 (N_9179,In_2860,In_1574);
nor U9180 (N_9180,In_4603,In_3236);
or U9181 (N_9181,In_3691,In_4702);
xor U9182 (N_9182,In_2271,In_3229);
and U9183 (N_9183,In_2423,In_1063);
nand U9184 (N_9184,In_1025,In_4798);
and U9185 (N_9185,In_500,In_1702);
and U9186 (N_9186,In_2073,In_866);
nor U9187 (N_9187,In_3017,In_2910);
and U9188 (N_9188,In_3840,In_3986);
nor U9189 (N_9189,In_3284,In_2225);
nor U9190 (N_9190,In_2954,In_419);
nand U9191 (N_9191,In_1762,In_3360);
xnor U9192 (N_9192,In_1276,In_661);
and U9193 (N_9193,In_4340,In_4688);
and U9194 (N_9194,In_4200,In_2420);
and U9195 (N_9195,In_4718,In_59);
and U9196 (N_9196,In_2359,In_776);
nor U9197 (N_9197,In_3148,In_3690);
xnor U9198 (N_9198,In_881,In_3243);
and U9199 (N_9199,In_2462,In_4850);
and U9200 (N_9200,In_471,In_784);
or U9201 (N_9201,In_2351,In_4586);
and U9202 (N_9202,In_2082,In_2649);
or U9203 (N_9203,In_4757,In_2802);
nand U9204 (N_9204,In_395,In_2000);
and U9205 (N_9205,In_1278,In_2246);
nand U9206 (N_9206,In_4037,In_3845);
nor U9207 (N_9207,In_3081,In_4174);
nand U9208 (N_9208,In_3929,In_286);
or U9209 (N_9209,In_1614,In_1892);
or U9210 (N_9210,In_117,In_4007);
nor U9211 (N_9211,In_431,In_2002);
xor U9212 (N_9212,In_4471,In_3158);
xor U9213 (N_9213,In_4926,In_4846);
nand U9214 (N_9214,In_43,In_1879);
xnor U9215 (N_9215,In_4889,In_898);
xor U9216 (N_9216,In_500,In_22);
nor U9217 (N_9217,In_217,In_3789);
nor U9218 (N_9218,In_732,In_2611);
or U9219 (N_9219,In_965,In_2600);
or U9220 (N_9220,In_771,In_1536);
nand U9221 (N_9221,In_1918,In_2484);
nand U9222 (N_9222,In_3251,In_1303);
nor U9223 (N_9223,In_768,In_289);
or U9224 (N_9224,In_2161,In_3903);
nor U9225 (N_9225,In_1756,In_4288);
and U9226 (N_9226,In_3976,In_3838);
and U9227 (N_9227,In_4370,In_3472);
and U9228 (N_9228,In_2228,In_671);
and U9229 (N_9229,In_2294,In_2181);
nor U9230 (N_9230,In_4089,In_1276);
nand U9231 (N_9231,In_2814,In_4245);
nand U9232 (N_9232,In_3604,In_4633);
nor U9233 (N_9233,In_1915,In_763);
or U9234 (N_9234,In_2849,In_1366);
xor U9235 (N_9235,In_2622,In_3375);
or U9236 (N_9236,In_1758,In_998);
nor U9237 (N_9237,In_1796,In_1629);
xnor U9238 (N_9238,In_3357,In_1503);
and U9239 (N_9239,In_1370,In_4602);
and U9240 (N_9240,In_3959,In_110);
xnor U9241 (N_9241,In_1596,In_76);
nand U9242 (N_9242,In_4746,In_1084);
or U9243 (N_9243,In_404,In_285);
xor U9244 (N_9244,In_234,In_3901);
or U9245 (N_9245,In_4908,In_986);
and U9246 (N_9246,In_2629,In_471);
and U9247 (N_9247,In_3348,In_2488);
xor U9248 (N_9248,In_4262,In_4766);
and U9249 (N_9249,In_2024,In_4771);
nand U9250 (N_9250,In_4684,In_4522);
or U9251 (N_9251,In_1362,In_4198);
nand U9252 (N_9252,In_4304,In_4801);
nand U9253 (N_9253,In_4340,In_1202);
nor U9254 (N_9254,In_2789,In_3810);
and U9255 (N_9255,In_3885,In_1350);
and U9256 (N_9256,In_1714,In_888);
nor U9257 (N_9257,In_1916,In_571);
nand U9258 (N_9258,In_971,In_2039);
nand U9259 (N_9259,In_1539,In_2014);
or U9260 (N_9260,In_2272,In_1773);
nand U9261 (N_9261,In_36,In_4637);
nor U9262 (N_9262,In_2767,In_2184);
and U9263 (N_9263,In_2623,In_168);
nor U9264 (N_9264,In_843,In_2543);
or U9265 (N_9265,In_191,In_2512);
and U9266 (N_9266,In_4437,In_2076);
and U9267 (N_9267,In_2761,In_2513);
xnor U9268 (N_9268,In_1376,In_355);
nor U9269 (N_9269,In_641,In_1873);
nor U9270 (N_9270,In_1973,In_2567);
nand U9271 (N_9271,In_3539,In_4533);
and U9272 (N_9272,In_6,In_3671);
xor U9273 (N_9273,In_56,In_2389);
or U9274 (N_9274,In_4061,In_1443);
nor U9275 (N_9275,In_3525,In_502);
nor U9276 (N_9276,In_4290,In_3045);
or U9277 (N_9277,In_4648,In_54);
xor U9278 (N_9278,In_196,In_4682);
nor U9279 (N_9279,In_1106,In_370);
and U9280 (N_9280,In_4513,In_2102);
and U9281 (N_9281,In_998,In_1941);
or U9282 (N_9282,In_4492,In_1032);
nor U9283 (N_9283,In_1250,In_3933);
xnor U9284 (N_9284,In_2651,In_3177);
or U9285 (N_9285,In_2672,In_1672);
nor U9286 (N_9286,In_1262,In_3419);
xor U9287 (N_9287,In_4710,In_4367);
or U9288 (N_9288,In_4284,In_4062);
and U9289 (N_9289,In_210,In_4815);
nand U9290 (N_9290,In_4404,In_2096);
nand U9291 (N_9291,In_2959,In_4210);
and U9292 (N_9292,In_2831,In_4391);
nor U9293 (N_9293,In_1924,In_3924);
and U9294 (N_9294,In_3570,In_4864);
and U9295 (N_9295,In_1293,In_2501);
nor U9296 (N_9296,In_1027,In_2618);
and U9297 (N_9297,In_1592,In_74);
nor U9298 (N_9298,In_4507,In_4896);
xnor U9299 (N_9299,In_3898,In_4053);
and U9300 (N_9300,In_1979,In_1048);
or U9301 (N_9301,In_4334,In_2214);
and U9302 (N_9302,In_1731,In_4486);
nand U9303 (N_9303,In_2549,In_3488);
nor U9304 (N_9304,In_2215,In_2718);
nand U9305 (N_9305,In_3747,In_4720);
nor U9306 (N_9306,In_4245,In_2266);
or U9307 (N_9307,In_4518,In_3269);
or U9308 (N_9308,In_352,In_4855);
and U9309 (N_9309,In_2052,In_1465);
or U9310 (N_9310,In_4366,In_1029);
nand U9311 (N_9311,In_4951,In_3245);
or U9312 (N_9312,In_141,In_4526);
and U9313 (N_9313,In_4850,In_3456);
nand U9314 (N_9314,In_4718,In_2180);
xor U9315 (N_9315,In_4822,In_828);
xnor U9316 (N_9316,In_2122,In_450);
or U9317 (N_9317,In_821,In_505);
or U9318 (N_9318,In_4063,In_1698);
xnor U9319 (N_9319,In_3745,In_1548);
xnor U9320 (N_9320,In_1210,In_4844);
and U9321 (N_9321,In_1315,In_4490);
xnor U9322 (N_9322,In_3337,In_1306);
nand U9323 (N_9323,In_1176,In_186);
nor U9324 (N_9324,In_2865,In_3489);
or U9325 (N_9325,In_4955,In_1645);
and U9326 (N_9326,In_4489,In_1932);
or U9327 (N_9327,In_995,In_3443);
nor U9328 (N_9328,In_520,In_758);
nor U9329 (N_9329,In_931,In_868);
xnor U9330 (N_9330,In_3157,In_2332);
xor U9331 (N_9331,In_3745,In_3161);
nand U9332 (N_9332,In_4796,In_3189);
or U9333 (N_9333,In_3448,In_3626);
or U9334 (N_9334,In_2644,In_4707);
and U9335 (N_9335,In_1853,In_527);
or U9336 (N_9336,In_4703,In_3375);
nor U9337 (N_9337,In_3556,In_2690);
xor U9338 (N_9338,In_912,In_1136);
nand U9339 (N_9339,In_175,In_2007);
nand U9340 (N_9340,In_762,In_759);
nand U9341 (N_9341,In_2268,In_855);
nor U9342 (N_9342,In_4609,In_3300);
or U9343 (N_9343,In_4114,In_1661);
or U9344 (N_9344,In_175,In_1497);
nor U9345 (N_9345,In_439,In_512);
nand U9346 (N_9346,In_61,In_3700);
or U9347 (N_9347,In_3268,In_53);
nand U9348 (N_9348,In_1118,In_3259);
nor U9349 (N_9349,In_4995,In_4708);
xnor U9350 (N_9350,In_3339,In_491);
nand U9351 (N_9351,In_4798,In_4111);
nor U9352 (N_9352,In_708,In_1804);
and U9353 (N_9353,In_295,In_1046);
nand U9354 (N_9354,In_1331,In_2726);
and U9355 (N_9355,In_1515,In_3911);
nand U9356 (N_9356,In_4449,In_3414);
xor U9357 (N_9357,In_3130,In_2528);
and U9358 (N_9358,In_1331,In_4744);
or U9359 (N_9359,In_1391,In_1736);
and U9360 (N_9360,In_4669,In_2252);
or U9361 (N_9361,In_1746,In_2043);
nor U9362 (N_9362,In_927,In_1682);
xnor U9363 (N_9363,In_3234,In_812);
xor U9364 (N_9364,In_695,In_1096);
and U9365 (N_9365,In_678,In_482);
or U9366 (N_9366,In_3307,In_1882);
or U9367 (N_9367,In_3354,In_2680);
and U9368 (N_9368,In_3758,In_250);
nand U9369 (N_9369,In_595,In_664);
or U9370 (N_9370,In_3709,In_2750);
or U9371 (N_9371,In_2753,In_2566);
or U9372 (N_9372,In_4746,In_788);
or U9373 (N_9373,In_3027,In_288);
xor U9374 (N_9374,In_1008,In_2769);
or U9375 (N_9375,In_3240,In_4602);
nor U9376 (N_9376,In_4595,In_1202);
nand U9377 (N_9377,In_2700,In_1769);
xnor U9378 (N_9378,In_4684,In_2711);
or U9379 (N_9379,In_3811,In_2101);
xnor U9380 (N_9380,In_627,In_717);
xor U9381 (N_9381,In_3755,In_463);
and U9382 (N_9382,In_2474,In_1653);
or U9383 (N_9383,In_3733,In_2877);
nand U9384 (N_9384,In_3721,In_1028);
nand U9385 (N_9385,In_3391,In_483);
nor U9386 (N_9386,In_2236,In_3419);
nand U9387 (N_9387,In_2908,In_4930);
nand U9388 (N_9388,In_4943,In_1831);
or U9389 (N_9389,In_1728,In_341);
nor U9390 (N_9390,In_4403,In_196);
xnor U9391 (N_9391,In_2326,In_812);
nor U9392 (N_9392,In_651,In_3334);
nor U9393 (N_9393,In_2370,In_4727);
or U9394 (N_9394,In_929,In_1459);
or U9395 (N_9395,In_2974,In_2041);
and U9396 (N_9396,In_2501,In_1414);
nand U9397 (N_9397,In_1581,In_2362);
nor U9398 (N_9398,In_1337,In_255);
and U9399 (N_9399,In_670,In_3673);
and U9400 (N_9400,In_1795,In_4074);
xnor U9401 (N_9401,In_4441,In_3915);
or U9402 (N_9402,In_1733,In_558);
xor U9403 (N_9403,In_4374,In_1910);
nand U9404 (N_9404,In_1119,In_3614);
and U9405 (N_9405,In_1772,In_1012);
xor U9406 (N_9406,In_3191,In_3316);
nor U9407 (N_9407,In_1397,In_3091);
or U9408 (N_9408,In_950,In_3908);
xor U9409 (N_9409,In_2023,In_1606);
and U9410 (N_9410,In_1551,In_3826);
xnor U9411 (N_9411,In_3979,In_4945);
nor U9412 (N_9412,In_4831,In_4722);
and U9413 (N_9413,In_2281,In_2688);
or U9414 (N_9414,In_4808,In_837);
nand U9415 (N_9415,In_3215,In_551);
nand U9416 (N_9416,In_2344,In_2952);
and U9417 (N_9417,In_2828,In_529);
nand U9418 (N_9418,In_4033,In_478);
nand U9419 (N_9419,In_3089,In_1470);
nand U9420 (N_9420,In_1618,In_3683);
xor U9421 (N_9421,In_120,In_841);
and U9422 (N_9422,In_2444,In_1568);
nor U9423 (N_9423,In_3746,In_2765);
nor U9424 (N_9424,In_795,In_3785);
nand U9425 (N_9425,In_3188,In_1238);
and U9426 (N_9426,In_2281,In_150);
and U9427 (N_9427,In_1221,In_3773);
or U9428 (N_9428,In_4910,In_1425);
xor U9429 (N_9429,In_3751,In_2614);
nand U9430 (N_9430,In_3001,In_2814);
nand U9431 (N_9431,In_925,In_1085);
nand U9432 (N_9432,In_2446,In_427);
and U9433 (N_9433,In_3276,In_1217);
nand U9434 (N_9434,In_1061,In_2774);
or U9435 (N_9435,In_521,In_20);
and U9436 (N_9436,In_2109,In_95);
or U9437 (N_9437,In_300,In_3970);
or U9438 (N_9438,In_138,In_105);
and U9439 (N_9439,In_2648,In_622);
xnor U9440 (N_9440,In_704,In_3638);
nand U9441 (N_9441,In_1042,In_1592);
nand U9442 (N_9442,In_691,In_2703);
and U9443 (N_9443,In_3630,In_981);
or U9444 (N_9444,In_10,In_1700);
nor U9445 (N_9445,In_2618,In_2808);
or U9446 (N_9446,In_4933,In_1388);
nor U9447 (N_9447,In_1480,In_2406);
xnor U9448 (N_9448,In_2268,In_2591);
xnor U9449 (N_9449,In_2614,In_3634);
nand U9450 (N_9450,In_4126,In_3251);
nand U9451 (N_9451,In_3469,In_597);
xnor U9452 (N_9452,In_2700,In_1402);
and U9453 (N_9453,In_2225,In_215);
and U9454 (N_9454,In_2438,In_4623);
and U9455 (N_9455,In_3781,In_2335);
and U9456 (N_9456,In_2197,In_102);
or U9457 (N_9457,In_1298,In_4943);
and U9458 (N_9458,In_2936,In_1982);
nor U9459 (N_9459,In_4360,In_3900);
nor U9460 (N_9460,In_1850,In_1260);
or U9461 (N_9461,In_1855,In_4333);
xor U9462 (N_9462,In_2691,In_365);
xor U9463 (N_9463,In_2482,In_4517);
nor U9464 (N_9464,In_2493,In_200);
nor U9465 (N_9465,In_2844,In_2463);
nor U9466 (N_9466,In_2715,In_1241);
xnor U9467 (N_9467,In_2643,In_765);
or U9468 (N_9468,In_4228,In_2646);
nor U9469 (N_9469,In_2915,In_4333);
nand U9470 (N_9470,In_1220,In_1674);
xor U9471 (N_9471,In_3931,In_2414);
or U9472 (N_9472,In_989,In_4255);
nor U9473 (N_9473,In_3085,In_1085);
xnor U9474 (N_9474,In_1021,In_37);
nor U9475 (N_9475,In_2153,In_4663);
or U9476 (N_9476,In_23,In_4578);
and U9477 (N_9477,In_1069,In_4858);
nor U9478 (N_9478,In_3345,In_4096);
and U9479 (N_9479,In_4266,In_4008);
nand U9480 (N_9480,In_3194,In_4371);
nand U9481 (N_9481,In_1628,In_1425);
nor U9482 (N_9482,In_1160,In_818);
and U9483 (N_9483,In_1409,In_1028);
xor U9484 (N_9484,In_1357,In_2240);
nand U9485 (N_9485,In_2685,In_2016);
xnor U9486 (N_9486,In_2734,In_1263);
nand U9487 (N_9487,In_16,In_4608);
and U9488 (N_9488,In_2708,In_119);
xnor U9489 (N_9489,In_1655,In_615);
and U9490 (N_9490,In_1943,In_1228);
and U9491 (N_9491,In_4199,In_4539);
nor U9492 (N_9492,In_2870,In_2905);
and U9493 (N_9493,In_2124,In_4040);
and U9494 (N_9494,In_3338,In_3143);
nand U9495 (N_9495,In_812,In_2564);
xor U9496 (N_9496,In_966,In_3871);
and U9497 (N_9497,In_397,In_4729);
or U9498 (N_9498,In_1615,In_1020);
or U9499 (N_9499,In_290,In_999);
nand U9500 (N_9500,In_1199,In_3896);
xor U9501 (N_9501,In_2779,In_601);
and U9502 (N_9502,In_2900,In_525);
xor U9503 (N_9503,In_3605,In_4518);
nand U9504 (N_9504,In_1688,In_283);
xor U9505 (N_9505,In_4786,In_2134);
or U9506 (N_9506,In_3168,In_2890);
and U9507 (N_9507,In_4845,In_2452);
nand U9508 (N_9508,In_4983,In_2749);
nor U9509 (N_9509,In_4393,In_1803);
xnor U9510 (N_9510,In_4751,In_2331);
and U9511 (N_9511,In_4036,In_4351);
xnor U9512 (N_9512,In_2137,In_1281);
and U9513 (N_9513,In_4068,In_778);
and U9514 (N_9514,In_4521,In_2085);
nand U9515 (N_9515,In_2554,In_465);
nand U9516 (N_9516,In_2559,In_4395);
nor U9517 (N_9517,In_2510,In_2925);
and U9518 (N_9518,In_591,In_697);
nor U9519 (N_9519,In_2996,In_4821);
xnor U9520 (N_9520,In_1457,In_749);
xnor U9521 (N_9521,In_2625,In_1007);
nor U9522 (N_9522,In_1512,In_1470);
and U9523 (N_9523,In_251,In_3390);
xor U9524 (N_9524,In_4619,In_329);
or U9525 (N_9525,In_3468,In_2337);
nor U9526 (N_9526,In_3900,In_2246);
or U9527 (N_9527,In_2010,In_4919);
or U9528 (N_9528,In_881,In_160);
or U9529 (N_9529,In_3819,In_2596);
nor U9530 (N_9530,In_4403,In_787);
nor U9531 (N_9531,In_3941,In_924);
nor U9532 (N_9532,In_3300,In_4399);
and U9533 (N_9533,In_4075,In_1500);
or U9534 (N_9534,In_3767,In_3941);
nor U9535 (N_9535,In_4827,In_0);
xor U9536 (N_9536,In_2872,In_1952);
nor U9537 (N_9537,In_3787,In_1680);
or U9538 (N_9538,In_2579,In_1040);
xor U9539 (N_9539,In_320,In_1796);
nor U9540 (N_9540,In_3186,In_4078);
nor U9541 (N_9541,In_1035,In_1264);
or U9542 (N_9542,In_2155,In_3741);
nor U9543 (N_9543,In_4013,In_3427);
nand U9544 (N_9544,In_2327,In_209);
or U9545 (N_9545,In_2405,In_1581);
xor U9546 (N_9546,In_2239,In_1017);
xnor U9547 (N_9547,In_3771,In_421);
nor U9548 (N_9548,In_4057,In_1249);
xor U9549 (N_9549,In_4265,In_3715);
nand U9550 (N_9550,In_2387,In_4182);
and U9551 (N_9551,In_819,In_2444);
nand U9552 (N_9552,In_3427,In_2628);
and U9553 (N_9553,In_1712,In_3592);
nand U9554 (N_9554,In_1742,In_1028);
xor U9555 (N_9555,In_3747,In_1316);
nor U9556 (N_9556,In_968,In_1733);
or U9557 (N_9557,In_3866,In_637);
or U9558 (N_9558,In_1304,In_2048);
nor U9559 (N_9559,In_3149,In_464);
nor U9560 (N_9560,In_1520,In_1304);
or U9561 (N_9561,In_4644,In_4208);
nand U9562 (N_9562,In_1677,In_2683);
nand U9563 (N_9563,In_4931,In_1890);
or U9564 (N_9564,In_1089,In_1600);
and U9565 (N_9565,In_4215,In_4288);
and U9566 (N_9566,In_2367,In_3168);
nand U9567 (N_9567,In_1302,In_3285);
and U9568 (N_9568,In_4218,In_2236);
nand U9569 (N_9569,In_2547,In_4203);
xor U9570 (N_9570,In_4644,In_2990);
and U9571 (N_9571,In_859,In_4852);
and U9572 (N_9572,In_4624,In_4061);
nand U9573 (N_9573,In_3752,In_511);
nor U9574 (N_9574,In_166,In_657);
nand U9575 (N_9575,In_66,In_4441);
xor U9576 (N_9576,In_4930,In_2525);
xnor U9577 (N_9577,In_2829,In_2910);
nor U9578 (N_9578,In_2440,In_580);
or U9579 (N_9579,In_4839,In_3563);
xor U9580 (N_9580,In_4582,In_4749);
and U9581 (N_9581,In_3488,In_238);
nor U9582 (N_9582,In_2544,In_4903);
nand U9583 (N_9583,In_4893,In_1638);
nand U9584 (N_9584,In_3213,In_891);
xor U9585 (N_9585,In_2027,In_4330);
and U9586 (N_9586,In_4024,In_1541);
nor U9587 (N_9587,In_3532,In_4679);
and U9588 (N_9588,In_4819,In_3475);
nor U9589 (N_9589,In_1257,In_1865);
xor U9590 (N_9590,In_4463,In_982);
and U9591 (N_9591,In_488,In_2106);
nand U9592 (N_9592,In_2494,In_4344);
or U9593 (N_9593,In_4959,In_1026);
nand U9594 (N_9594,In_1218,In_2161);
and U9595 (N_9595,In_3719,In_4538);
nor U9596 (N_9596,In_3085,In_2935);
and U9597 (N_9597,In_4950,In_2178);
nor U9598 (N_9598,In_1321,In_865);
and U9599 (N_9599,In_1054,In_3553);
nand U9600 (N_9600,In_2141,In_499);
and U9601 (N_9601,In_3623,In_121);
or U9602 (N_9602,In_415,In_4249);
or U9603 (N_9603,In_2376,In_245);
nor U9604 (N_9604,In_3211,In_4348);
nand U9605 (N_9605,In_818,In_2859);
xor U9606 (N_9606,In_2701,In_306);
or U9607 (N_9607,In_3055,In_4177);
and U9608 (N_9608,In_3879,In_4862);
nor U9609 (N_9609,In_4121,In_182);
and U9610 (N_9610,In_3595,In_3012);
or U9611 (N_9611,In_2120,In_4019);
or U9612 (N_9612,In_209,In_870);
nand U9613 (N_9613,In_3606,In_2591);
nand U9614 (N_9614,In_4906,In_626);
xor U9615 (N_9615,In_773,In_512);
or U9616 (N_9616,In_1494,In_2996);
nor U9617 (N_9617,In_4662,In_3379);
nor U9618 (N_9618,In_2181,In_3351);
or U9619 (N_9619,In_2512,In_1805);
xor U9620 (N_9620,In_893,In_1147);
or U9621 (N_9621,In_148,In_2696);
or U9622 (N_9622,In_3550,In_3308);
nor U9623 (N_9623,In_1428,In_411);
nand U9624 (N_9624,In_2798,In_381);
nand U9625 (N_9625,In_42,In_4655);
nand U9626 (N_9626,In_33,In_635);
nor U9627 (N_9627,In_4934,In_1977);
nor U9628 (N_9628,In_1242,In_835);
nor U9629 (N_9629,In_3719,In_2093);
or U9630 (N_9630,In_952,In_4302);
xnor U9631 (N_9631,In_4937,In_2707);
and U9632 (N_9632,In_2010,In_2483);
xnor U9633 (N_9633,In_1000,In_3234);
nor U9634 (N_9634,In_306,In_584);
and U9635 (N_9635,In_1274,In_118);
xor U9636 (N_9636,In_2060,In_934);
xnor U9637 (N_9637,In_408,In_3147);
nor U9638 (N_9638,In_892,In_456);
and U9639 (N_9639,In_1641,In_3212);
nor U9640 (N_9640,In_2244,In_4668);
xor U9641 (N_9641,In_2663,In_4902);
and U9642 (N_9642,In_4167,In_4883);
or U9643 (N_9643,In_3155,In_1912);
nand U9644 (N_9644,In_714,In_2792);
or U9645 (N_9645,In_2277,In_2040);
nand U9646 (N_9646,In_21,In_391);
or U9647 (N_9647,In_2514,In_2042);
xor U9648 (N_9648,In_843,In_2563);
nor U9649 (N_9649,In_4621,In_3935);
or U9650 (N_9650,In_3334,In_3572);
nor U9651 (N_9651,In_4306,In_222);
xor U9652 (N_9652,In_419,In_3611);
and U9653 (N_9653,In_2902,In_2948);
xnor U9654 (N_9654,In_1999,In_540);
and U9655 (N_9655,In_493,In_4465);
or U9656 (N_9656,In_2007,In_1522);
xnor U9657 (N_9657,In_381,In_73);
or U9658 (N_9658,In_4797,In_35);
nor U9659 (N_9659,In_2650,In_4205);
and U9660 (N_9660,In_1539,In_999);
or U9661 (N_9661,In_2593,In_4174);
and U9662 (N_9662,In_1146,In_2540);
nand U9663 (N_9663,In_3547,In_780);
nor U9664 (N_9664,In_4298,In_4923);
and U9665 (N_9665,In_2847,In_2177);
and U9666 (N_9666,In_1411,In_1427);
nand U9667 (N_9667,In_4569,In_2068);
nor U9668 (N_9668,In_169,In_396);
nand U9669 (N_9669,In_3126,In_566);
xnor U9670 (N_9670,In_1102,In_1472);
xnor U9671 (N_9671,In_588,In_4393);
xnor U9672 (N_9672,In_1866,In_254);
or U9673 (N_9673,In_4341,In_1937);
xor U9674 (N_9674,In_2300,In_1188);
or U9675 (N_9675,In_439,In_2877);
and U9676 (N_9676,In_2222,In_230);
nand U9677 (N_9677,In_2224,In_1863);
and U9678 (N_9678,In_1980,In_4737);
or U9679 (N_9679,In_1175,In_4325);
nor U9680 (N_9680,In_4898,In_505);
or U9681 (N_9681,In_916,In_2542);
nand U9682 (N_9682,In_1450,In_0);
nor U9683 (N_9683,In_355,In_4564);
xnor U9684 (N_9684,In_3912,In_3168);
or U9685 (N_9685,In_2460,In_1260);
nor U9686 (N_9686,In_4019,In_3156);
and U9687 (N_9687,In_4554,In_1910);
nor U9688 (N_9688,In_1758,In_3676);
xnor U9689 (N_9689,In_447,In_1583);
xnor U9690 (N_9690,In_4858,In_4031);
xnor U9691 (N_9691,In_2383,In_4372);
or U9692 (N_9692,In_2346,In_2733);
xor U9693 (N_9693,In_2289,In_2389);
nand U9694 (N_9694,In_1992,In_1176);
nand U9695 (N_9695,In_4850,In_498);
nand U9696 (N_9696,In_1655,In_4911);
or U9697 (N_9697,In_2701,In_2429);
nand U9698 (N_9698,In_42,In_4616);
nor U9699 (N_9699,In_2016,In_2423);
nand U9700 (N_9700,In_1729,In_259);
or U9701 (N_9701,In_2622,In_4019);
nand U9702 (N_9702,In_4374,In_2098);
nand U9703 (N_9703,In_4622,In_4868);
and U9704 (N_9704,In_1165,In_3983);
xor U9705 (N_9705,In_613,In_3920);
xor U9706 (N_9706,In_4631,In_205);
nor U9707 (N_9707,In_2576,In_4696);
or U9708 (N_9708,In_3327,In_3302);
xor U9709 (N_9709,In_1894,In_2625);
nor U9710 (N_9710,In_4254,In_212);
xor U9711 (N_9711,In_2440,In_538);
or U9712 (N_9712,In_426,In_369);
or U9713 (N_9713,In_988,In_3321);
and U9714 (N_9714,In_2107,In_1090);
xnor U9715 (N_9715,In_4559,In_1121);
nand U9716 (N_9716,In_1033,In_2907);
nor U9717 (N_9717,In_1411,In_908);
nand U9718 (N_9718,In_4049,In_4201);
nand U9719 (N_9719,In_4766,In_4046);
and U9720 (N_9720,In_2032,In_675);
or U9721 (N_9721,In_3200,In_1411);
xnor U9722 (N_9722,In_811,In_2060);
and U9723 (N_9723,In_4639,In_2335);
or U9724 (N_9724,In_4461,In_1741);
nor U9725 (N_9725,In_727,In_629);
nand U9726 (N_9726,In_1127,In_2905);
nor U9727 (N_9727,In_8,In_4277);
nand U9728 (N_9728,In_3907,In_4435);
nor U9729 (N_9729,In_4688,In_3110);
or U9730 (N_9730,In_4553,In_3383);
and U9731 (N_9731,In_1457,In_2385);
xnor U9732 (N_9732,In_1143,In_4875);
xnor U9733 (N_9733,In_2377,In_3439);
or U9734 (N_9734,In_4804,In_4940);
nor U9735 (N_9735,In_2493,In_3211);
xnor U9736 (N_9736,In_2173,In_1750);
and U9737 (N_9737,In_1035,In_2898);
and U9738 (N_9738,In_4577,In_1870);
or U9739 (N_9739,In_1227,In_13);
xnor U9740 (N_9740,In_730,In_4304);
nand U9741 (N_9741,In_2637,In_2095);
xnor U9742 (N_9742,In_387,In_846);
and U9743 (N_9743,In_3068,In_2196);
xor U9744 (N_9744,In_978,In_3325);
or U9745 (N_9745,In_2139,In_3149);
xnor U9746 (N_9746,In_3829,In_3049);
or U9747 (N_9747,In_2653,In_1173);
nand U9748 (N_9748,In_1863,In_3044);
nand U9749 (N_9749,In_1682,In_1910);
nand U9750 (N_9750,In_2271,In_1015);
nor U9751 (N_9751,In_2413,In_223);
nor U9752 (N_9752,In_1211,In_3667);
or U9753 (N_9753,In_3984,In_1562);
or U9754 (N_9754,In_3161,In_547);
and U9755 (N_9755,In_3309,In_1748);
or U9756 (N_9756,In_4826,In_4193);
and U9757 (N_9757,In_3784,In_645);
or U9758 (N_9758,In_2,In_2509);
nor U9759 (N_9759,In_1147,In_4305);
nor U9760 (N_9760,In_3806,In_1557);
nor U9761 (N_9761,In_4977,In_1018);
nor U9762 (N_9762,In_1159,In_2909);
nor U9763 (N_9763,In_4765,In_2827);
and U9764 (N_9764,In_3349,In_728);
and U9765 (N_9765,In_4777,In_4652);
nor U9766 (N_9766,In_573,In_3268);
nor U9767 (N_9767,In_4318,In_1639);
or U9768 (N_9768,In_3179,In_4043);
nor U9769 (N_9769,In_1596,In_2415);
nor U9770 (N_9770,In_774,In_2830);
or U9771 (N_9771,In_4810,In_2090);
or U9772 (N_9772,In_1855,In_2995);
nor U9773 (N_9773,In_2662,In_1125);
nor U9774 (N_9774,In_4967,In_148);
xnor U9775 (N_9775,In_2956,In_2906);
xor U9776 (N_9776,In_3258,In_3612);
and U9777 (N_9777,In_2382,In_3400);
nor U9778 (N_9778,In_4271,In_3049);
nor U9779 (N_9779,In_2168,In_3217);
and U9780 (N_9780,In_1262,In_511);
and U9781 (N_9781,In_338,In_3307);
xor U9782 (N_9782,In_3170,In_260);
xnor U9783 (N_9783,In_4872,In_1124);
and U9784 (N_9784,In_444,In_1217);
nand U9785 (N_9785,In_260,In_1782);
or U9786 (N_9786,In_1494,In_245);
xor U9787 (N_9787,In_1931,In_2898);
nand U9788 (N_9788,In_906,In_2701);
nand U9789 (N_9789,In_475,In_4701);
xnor U9790 (N_9790,In_2786,In_4497);
nand U9791 (N_9791,In_4398,In_2661);
or U9792 (N_9792,In_1869,In_2596);
nand U9793 (N_9793,In_3591,In_342);
nor U9794 (N_9794,In_779,In_1860);
xor U9795 (N_9795,In_48,In_2659);
xor U9796 (N_9796,In_3674,In_966);
or U9797 (N_9797,In_3623,In_3240);
and U9798 (N_9798,In_1766,In_2915);
nor U9799 (N_9799,In_966,In_3857);
nor U9800 (N_9800,In_3367,In_4100);
nand U9801 (N_9801,In_1129,In_12);
nor U9802 (N_9802,In_4658,In_3523);
xnor U9803 (N_9803,In_4190,In_1331);
or U9804 (N_9804,In_356,In_2699);
or U9805 (N_9805,In_1152,In_2541);
xor U9806 (N_9806,In_4474,In_633);
nor U9807 (N_9807,In_1483,In_2383);
nor U9808 (N_9808,In_3312,In_1132);
or U9809 (N_9809,In_1951,In_1113);
xnor U9810 (N_9810,In_1686,In_1049);
nand U9811 (N_9811,In_4437,In_4411);
nand U9812 (N_9812,In_1641,In_1531);
nor U9813 (N_9813,In_2133,In_3273);
nand U9814 (N_9814,In_2565,In_3997);
and U9815 (N_9815,In_1131,In_289);
nor U9816 (N_9816,In_2930,In_2294);
or U9817 (N_9817,In_2789,In_2518);
nand U9818 (N_9818,In_2593,In_2995);
nor U9819 (N_9819,In_718,In_4170);
nor U9820 (N_9820,In_3635,In_4091);
nor U9821 (N_9821,In_340,In_105);
nor U9822 (N_9822,In_4610,In_3043);
nor U9823 (N_9823,In_728,In_3247);
and U9824 (N_9824,In_4702,In_1722);
xor U9825 (N_9825,In_1756,In_3507);
nor U9826 (N_9826,In_867,In_4825);
and U9827 (N_9827,In_1022,In_2378);
xnor U9828 (N_9828,In_1178,In_583);
nand U9829 (N_9829,In_4593,In_3525);
xor U9830 (N_9830,In_1070,In_980);
and U9831 (N_9831,In_4798,In_3589);
and U9832 (N_9832,In_4752,In_1057);
nand U9833 (N_9833,In_4420,In_3500);
nor U9834 (N_9834,In_2995,In_3088);
nor U9835 (N_9835,In_2782,In_1571);
or U9836 (N_9836,In_1530,In_2605);
and U9837 (N_9837,In_2111,In_1761);
nor U9838 (N_9838,In_4986,In_3997);
xnor U9839 (N_9839,In_1023,In_3155);
nor U9840 (N_9840,In_3457,In_921);
or U9841 (N_9841,In_4408,In_2479);
nor U9842 (N_9842,In_2902,In_3786);
nor U9843 (N_9843,In_4417,In_2455);
xnor U9844 (N_9844,In_360,In_1775);
xor U9845 (N_9845,In_3099,In_4538);
and U9846 (N_9846,In_245,In_3623);
xor U9847 (N_9847,In_3129,In_1490);
xnor U9848 (N_9848,In_920,In_3374);
or U9849 (N_9849,In_3813,In_9);
nor U9850 (N_9850,In_2600,In_453);
and U9851 (N_9851,In_4150,In_2661);
and U9852 (N_9852,In_3751,In_3366);
or U9853 (N_9853,In_2026,In_4371);
nor U9854 (N_9854,In_3819,In_3753);
nor U9855 (N_9855,In_1577,In_4606);
nor U9856 (N_9856,In_1948,In_3946);
xor U9857 (N_9857,In_2310,In_4932);
and U9858 (N_9858,In_2407,In_4071);
nand U9859 (N_9859,In_434,In_77);
or U9860 (N_9860,In_2678,In_4511);
xnor U9861 (N_9861,In_3215,In_212);
or U9862 (N_9862,In_3728,In_1063);
and U9863 (N_9863,In_3470,In_2450);
nor U9864 (N_9864,In_110,In_1130);
nor U9865 (N_9865,In_3114,In_4798);
or U9866 (N_9866,In_1714,In_4780);
xnor U9867 (N_9867,In_4944,In_3382);
nand U9868 (N_9868,In_2719,In_2090);
or U9869 (N_9869,In_2975,In_4643);
and U9870 (N_9870,In_1415,In_3058);
and U9871 (N_9871,In_3923,In_647);
nor U9872 (N_9872,In_4744,In_4990);
nand U9873 (N_9873,In_4299,In_1494);
nor U9874 (N_9874,In_2771,In_4048);
nand U9875 (N_9875,In_2640,In_4554);
or U9876 (N_9876,In_1334,In_4221);
nand U9877 (N_9877,In_896,In_191);
nand U9878 (N_9878,In_891,In_4045);
and U9879 (N_9879,In_4562,In_4557);
nor U9880 (N_9880,In_996,In_3793);
or U9881 (N_9881,In_3294,In_2923);
nand U9882 (N_9882,In_4370,In_193);
and U9883 (N_9883,In_635,In_3649);
xnor U9884 (N_9884,In_3975,In_3669);
xnor U9885 (N_9885,In_1296,In_4238);
xor U9886 (N_9886,In_37,In_2570);
or U9887 (N_9887,In_4212,In_1447);
xnor U9888 (N_9888,In_1879,In_3308);
nor U9889 (N_9889,In_90,In_1135);
and U9890 (N_9890,In_2674,In_2758);
nand U9891 (N_9891,In_3532,In_2169);
nor U9892 (N_9892,In_2974,In_405);
nor U9893 (N_9893,In_2427,In_1441);
xor U9894 (N_9894,In_2283,In_548);
and U9895 (N_9895,In_587,In_2565);
xnor U9896 (N_9896,In_2113,In_4807);
and U9897 (N_9897,In_2372,In_636);
nor U9898 (N_9898,In_4218,In_3338);
xor U9899 (N_9899,In_2168,In_790);
or U9900 (N_9900,In_2632,In_779);
nand U9901 (N_9901,In_4234,In_4097);
xnor U9902 (N_9902,In_2874,In_3962);
xor U9903 (N_9903,In_2566,In_2554);
nor U9904 (N_9904,In_538,In_1981);
nand U9905 (N_9905,In_2438,In_3328);
or U9906 (N_9906,In_2464,In_1025);
or U9907 (N_9907,In_3568,In_189);
xnor U9908 (N_9908,In_1289,In_16);
and U9909 (N_9909,In_3785,In_4311);
and U9910 (N_9910,In_1517,In_723);
and U9911 (N_9911,In_4943,In_792);
nor U9912 (N_9912,In_4671,In_4246);
and U9913 (N_9913,In_729,In_3526);
or U9914 (N_9914,In_4189,In_4918);
nor U9915 (N_9915,In_3390,In_3300);
nor U9916 (N_9916,In_2702,In_445);
nand U9917 (N_9917,In_2796,In_2833);
nand U9918 (N_9918,In_1451,In_2900);
and U9919 (N_9919,In_3839,In_3698);
xnor U9920 (N_9920,In_1472,In_4184);
xor U9921 (N_9921,In_2512,In_2080);
nor U9922 (N_9922,In_83,In_1579);
or U9923 (N_9923,In_3992,In_3513);
xnor U9924 (N_9924,In_2779,In_1136);
xnor U9925 (N_9925,In_2086,In_1620);
and U9926 (N_9926,In_3628,In_3333);
or U9927 (N_9927,In_1486,In_196);
nand U9928 (N_9928,In_314,In_1083);
nor U9929 (N_9929,In_2162,In_3427);
nor U9930 (N_9930,In_4742,In_4029);
or U9931 (N_9931,In_58,In_2002);
nor U9932 (N_9932,In_197,In_2296);
nand U9933 (N_9933,In_254,In_4777);
and U9934 (N_9934,In_2200,In_2376);
xor U9935 (N_9935,In_1709,In_652);
nor U9936 (N_9936,In_3182,In_392);
nor U9937 (N_9937,In_1986,In_4419);
or U9938 (N_9938,In_778,In_4269);
or U9939 (N_9939,In_2699,In_4867);
or U9940 (N_9940,In_1992,In_4016);
or U9941 (N_9941,In_2625,In_1227);
and U9942 (N_9942,In_2321,In_2408);
and U9943 (N_9943,In_1087,In_4174);
xor U9944 (N_9944,In_1152,In_1961);
xor U9945 (N_9945,In_1157,In_4608);
nand U9946 (N_9946,In_1420,In_4323);
or U9947 (N_9947,In_3891,In_2748);
xor U9948 (N_9948,In_3261,In_3856);
or U9949 (N_9949,In_4473,In_1796);
or U9950 (N_9950,In_3839,In_67);
xor U9951 (N_9951,In_4498,In_1248);
nor U9952 (N_9952,In_856,In_4782);
nor U9953 (N_9953,In_2261,In_2263);
xor U9954 (N_9954,In_650,In_50);
xor U9955 (N_9955,In_4872,In_2259);
nand U9956 (N_9956,In_1058,In_4632);
or U9957 (N_9957,In_2285,In_4479);
xnor U9958 (N_9958,In_2162,In_4864);
nand U9959 (N_9959,In_961,In_3511);
xnor U9960 (N_9960,In_4553,In_4557);
nor U9961 (N_9961,In_2615,In_1827);
xnor U9962 (N_9962,In_2902,In_1485);
and U9963 (N_9963,In_2939,In_1512);
nand U9964 (N_9964,In_4576,In_1316);
nand U9965 (N_9965,In_1055,In_4705);
and U9966 (N_9966,In_2647,In_1818);
or U9967 (N_9967,In_622,In_1634);
nor U9968 (N_9968,In_1670,In_4823);
xnor U9969 (N_9969,In_506,In_2201);
nand U9970 (N_9970,In_1110,In_1276);
and U9971 (N_9971,In_866,In_2663);
xor U9972 (N_9972,In_4546,In_4353);
and U9973 (N_9973,In_143,In_1505);
and U9974 (N_9974,In_562,In_19);
or U9975 (N_9975,In_3780,In_179);
nand U9976 (N_9976,In_2363,In_37);
or U9977 (N_9977,In_2573,In_2634);
xnor U9978 (N_9978,In_3234,In_20);
nor U9979 (N_9979,In_632,In_1477);
xor U9980 (N_9980,In_4464,In_3937);
nand U9981 (N_9981,In_1706,In_3066);
and U9982 (N_9982,In_2797,In_3730);
and U9983 (N_9983,In_3118,In_1491);
nand U9984 (N_9984,In_2393,In_3899);
xor U9985 (N_9985,In_3241,In_657);
nand U9986 (N_9986,In_2954,In_2180);
xor U9987 (N_9987,In_4553,In_3962);
and U9988 (N_9988,In_2144,In_941);
and U9989 (N_9989,In_3336,In_350);
nand U9990 (N_9990,In_3453,In_4160);
nand U9991 (N_9991,In_1633,In_182);
xnor U9992 (N_9992,In_4160,In_3550);
and U9993 (N_9993,In_3686,In_1011);
nand U9994 (N_9994,In_4776,In_2291);
xor U9995 (N_9995,In_4735,In_424);
and U9996 (N_9996,In_1945,In_2827);
and U9997 (N_9997,In_496,In_2026);
and U9998 (N_9998,In_1574,In_73);
nand U9999 (N_9999,In_1382,In_1689);
xor U10000 (N_10000,N_965,N_4944);
nor U10001 (N_10001,N_7669,N_9119);
nor U10002 (N_10002,N_8342,N_3009);
xor U10003 (N_10003,N_5449,N_9003);
nor U10004 (N_10004,N_2990,N_5584);
and U10005 (N_10005,N_4673,N_5973);
xor U10006 (N_10006,N_4030,N_1473);
xor U10007 (N_10007,N_3208,N_130);
and U10008 (N_10008,N_1850,N_9837);
and U10009 (N_10009,N_3258,N_2404);
or U10010 (N_10010,N_3046,N_5617);
xor U10011 (N_10011,N_5125,N_2931);
nand U10012 (N_10012,N_9930,N_2830);
and U10013 (N_10013,N_9297,N_5732);
xnor U10014 (N_10014,N_2254,N_5667);
nor U10015 (N_10015,N_9693,N_2494);
and U10016 (N_10016,N_3468,N_9536);
nand U10017 (N_10017,N_2809,N_9032);
or U10018 (N_10018,N_8541,N_1938);
nand U10019 (N_10019,N_9324,N_8801);
nand U10020 (N_10020,N_209,N_1841);
or U10021 (N_10021,N_3603,N_2764);
or U10022 (N_10022,N_4273,N_4354);
and U10023 (N_10023,N_895,N_743);
xnor U10024 (N_10024,N_3722,N_7750);
or U10025 (N_10025,N_2166,N_5517);
and U10026 (N_10026,N_2125,N_3538);
or U10027 (N_10027,N_1802,N_2019);
xor U10028 (N_10028,N_2612,N_4027);
and U10029 (N_10029,N_4933,N_4369);
and U10030 (N_10030,N_4500,N_7674);
nand U10031 (N_10031,N_6273,N_6210);
and U10032 (N_10032,N_3660,N_5726);
nand U10033 (N_10033,N_7956,N_9364);
xor U10034 (N_10034,N_4654,N_8688);
nand U10035 (N_10035,N_9627,N_5211);
xnor U10036 (N_10036,N_2514,N_105);
nor U10037 (N_10037,N_9157,N_828);
xor U10038 (N_10038,N_3,N_9701);
and U10039 (N_10039,N_4447,N_0);
nand U10040 (N_10040,N_3813,N_3051);
xor U10041 (N_10041,N_5794,N_4598);
xor U10042 (N_10042,N_3123,N_3186);
nand U10043 (N_10043,N_9772,N_1102);
xor U10044 (N_10044,N_8737,N_4525);
nand U10045 (N_10045,N_2292,N_9635);
xor U10046 (N_10046,N_6139,N_2621);
xnor U10047 (N_10047,N_5679,N_6836);
xnor U10048 (N_10048,N_2093,N_5915);
and U10049 (N_10049,N_2556,N_5312);
nand U10050 (N_10050,N_9156,N_7790);
xor U10051 (N_10051,N_2143,N_6870);
and U10052 (N_10052,N_8225,N_8162);
nor U10053 (N_10053,N_45,N_1664);
nor U10054 (N_10054,N_4633,N_3557);
or U10055 (N_10055,N_6051,N_9608);
nand U10056 (N_10056,N_8927,N_9940);
and U10057 (N_10057,N_6153,N_4863);
and U10058 (N_10058,N_7158,N_7753);
nand U10059 (N_10059,N_2918,N_5146);
or U10060 (N_10060,N_9880,N_9028);
or U10061 (N_10061,N_9495,N_326);
and U10062 (N_10062,N_5480,N_5697);
nor U10063 (N_10063,N_3435,N_8115);
nor U10064 (N_10064,N_6391,N_2785);
nand U10065 (N_10065,N_5583,N_8234);
and U10066 (N_10066,N_8623,N_5468);
nor U10067 (N_10067,N_1344,N_5519);
or U10068 (N_10068,N_5776,N_7567);
nand U10069 (N_10069,N_6242,N_685);
xnor U10070 (N_10070,N_1370,N_2688);
or U10071 (N_10071,N_4743,N_1847);
and U10072 (N_10072,N_1032,N_102);
and U10073 (N_10073,N_9278,N_795);
and U10074 (N_10074,N_4553,N_3755);
and U10075 (N_10075,N_7619,N_6916);
nand U10076 (N_10076,N_8107,N_1732);
and U10077 (N_10077,N_1333,N_5103);
and U10078 (N_10078,N_2564,N_3891);
xnor U10079 (N_10079,N_3529,N_3792);
or U10080 (N_10080,N_1718,N_5147);
nand U10081 (N_10081,N_386,N_3068);
nand U10082 (N_10082,N_7818,N_8475);
nor U10083 (N_10083,N_4821,N_5864);
xor U10084 (N_10084,N_6887,N_3183);
nor U10085 (N_10085,N_9260,N_2988);
and U10086 (N_10086,N_1899,N_1498);
nor U10087 (N_10087,N_8564,N_9974);
xor U10088 (N_10088,N_6117,N_7070);
xnor U10089 (N_10089,N_9418,N_3929);
or U10090 (N_10090,N_4586,N_3428);
and U10091 (N_10091,N_7172,N_885);
nand U10092 (N_10092,N_8991,N_9180);
nand U10093 (N_10093,N_7885,N_1894);
or U10094 (N_10094,N_6027,N_6364);
xnor U10095 (N_10095,N_5887,N_182);
nor U10096 (N_10096,N_9673,N_2579);
nor U10097 (N_10097,N_3243,N_4389);
nand U10098 (N_10098,N_8016,N_7940);
xnor U10099 (N_10099,N_2325,N_5040);
and U10100 (N_10100,N_1050,N_3418);
xnor U10101 (N_10101,N_4861,N_5423);
or U10102 (N_10102,N_5443,N_8183);
xnor U10103 (N_10103,N_6322,N_512);
and U10104 (N_10104,N_2239,N_2220);
nor U10105 (N_10105,N_3425,N_1786);
nand U10106 (N_10106,N_2884,N_8233);
or U10107 (N_10107,N_3732,N_4958);
nor U10108 (N_10108,N_3461,N_4067);
nand U10109 (N_10109,N_3297,N_2369);
xor U10110 (N_10110,N_9247,N_6118);
and U10111 (N_10111,N_4339,N_8748);
nor U10112 (N_10112,N_8866,N_4057);
and U10113 (N_10113,N_2316,N_750);
or U10114 (N_10114,N_7634,N_9077);
xor U10115 (N_10115,N_1129,N_9525);
or U10116 (N_10116,N_9195,N_247);
nor U10117 (N_10117,N_6132,N_4547);
nand U10118 (N_10118,N_6263,N_5552);
nor U10119 (N_10119,N_1235,N_5886);
nor U10120 (N_10120,N_237,N_6740);
nand U10121 (N_10121,N_4597,N_356);
and U10122 (N_10122,N_5326,N_5350);
and U10123 (N_10123,N_6513,N_4953);
and U10124 (N_10124,N_5965,N_1573);
nor U10125 (N_10125,N_8766,N_9116);
xor U10126 (N_10126,N_7913,N_7056);
nand U10127 (N_10127,N_9140,N_9506);
xor U10128 (N_10128,N_1376,N_5009);
xnor U10129 (N_10129,N_7726,N_2018);
and U10130 (N_10130,N_9092,N_1010);
or U10131 (N_10131,N_990,N_6280);
or U10132 (N_10132,N_6743,N_918);
nand U10133 (N_10133,N_7266,N_5404);
xnor U10134 (N_10134,N_2004,N_2845);
or U10135 (N_10135,N_8284,N_7520);
and U10136 (N_10136,N_9395,N_2469);
nor U10137 (N_10137,N_9282,N_9496);
or U10138 (N_10138,N_274,N_5899);
and U10139 (N_10139,N_3867,N_5734);
xnor U10140 (N_10140,N_5045,N_3071);
and U10141 (N_10141,N_865,N_7420);
nand U10142 (N_10142,N_7960,N_1608);
or U10143 (N_10143,N_2246,N_5665);
and U10144 (N_10144,N_7624,N_4559);
nand U10145 (N_10145,N_2952,N_6402);
or U10146 (N_10146,N_4835,N_5635);
or U10147 (N_10147,N_2173,N_3658);
nand U10148 (N_10148,N_3798,N_9569);
nor U10149 (N_10149,N_6438,N_168);
xor U10150 (N_10150,N_8851,N_3482);
or U10151 (N_10151,N_9522,N_7336);
and U10152 (N_10152,N_2695,N_5558);
and U10153 (N_10153,N_7810,N_5591);
xor U10154 (N_10154,N_2328,N_7493);
nand U10155 (N_10155,N_7995,N_2862);
nor U10156 (N_10156,N_9838,N_3040);
xnor U10157 (N_10157,N_7078,N_5600);
nor U10158 (N_10158,N_4956,N_5546);
and U10159 (N_10159,N_3432,N_4371);
nor U10160 (N_10160,N_4342,N_7282);
nor U10161 (N_10161,N_2135,N_434);
or U10162 (N_10162,N_2049,N_7800);
nor U10163 (N_10163,N_6356,N_8759);
nand U10164 (N_10164,N_9558,N_6468);
xnor U10165 (N_10165,N_6232,N_6741);
and U10166 (N_10166,N_2443,N_8007);
or U10167 (N_10167,N_4803,N_2545);
and U10168 (N_10168,N_1578,N_1457);
or U10169 (N_10169,N_5202,N_6604);
nor U10170 (N_10170,N_502,N_7920);
xor U10171 (N_10171,N_8753,N_6727);
nand U10172 (N_10172,N_3153,N_6613);
nor U10173 (N_10173,N_3066,N_9578);
and U10174 (N_10174,N_8572,N_481);
xor U10175 (N_10175,N_6247,N_1643);
nor U10176 (N_10176,N_1428,N_1227);
and U10177 (N_10177,N_549,N_2281);
xor U10178 (N_10178,N_8716,N_4032);
or U10179 (N_10179,N_3905,N_3528);
nor U10180 (N_10180,N_7093,N_692);
xnor U10181 (N_10181,N_5702,N_3246);
nor U10182 (N_10182,N_5150,N_559);
xor U10183 (N_10183,N_9261,N_5076);
and U10184 (N_10184,N_9053,N_5460);
xor U10185 (N_10185,N_1931,N_2327);
xor U10186 (N_10186,N_8656,N_3713);
nand U10187 (N_10187,N_8486,N_3894);
nor U10188 (N_10188,N_4667,N_5230);
nand U10189 (N_10189,N_6233,N_5335);
xnor U10190 (N_10190,N_9223,N_9586);
nand U10191 (N_10191,N_1682,N_4687);
and U10192 (N_10192,N_7397,N_4570);
nor U10193 (N_10193,N_7723,N_6845);
nor U10194 (N_10194,N_6589,N_8336);
nand U10195 (N_10195,N_5920,N_8430);
or U10196 (N_10196,N_4504,N_4441);
nand U10197 (N_10197,N_9492,N_8278);
xor U10198 (N_10198,N_2763,N_2979);
nor U10199 (N_10199,N_6544,N_5269);
nor U10200 (N_10200,N_5588,N_8586);
and U10201 (N_10201,N_6086,N_775);
and U10202 (N_10202,N_6180,N_335);
and U10203 (N_10203,N_7646,N_8076);
xnor U10204 (N_10204,N_5755,N_9800);
or U10205 (N_10205,N_6176,N_6196);
nand U10206 (N_10206,N_4400,N_7602);
nand U10207 (N_10207,N_6899,N_2784);
xor U10208 (N_10208,N_9726,N_3812);
nand U10209 (N_10209,N_8678,N_3512);
nand U10210 (N_10210,N_3061,N_1556);
nand U10211 (N_10211,N_3586,N_7895);
and U10212 (N_10212,N_4359,N_9802);
xnor U10213 (N_10213,N_2757,N_5652);
and U10214 (N_10214,N_7805,N_2727);
nor U10215 (N_10215,N_3730,N_4193);
and U10216 (N_10216,N_6760,N_4170);
nand U10217 (N_10217,N_6819,N_781);
xnor U10218 (N_10218,N_7456,N_8964);
nor U10219 (N_10219,N_7419,N_7804);
nor U10220 (N_10220,N_63,N_6189);
or U10221 (N_10221,N_7111,N_4859);
nand U10222 (N_10222,N_7533,N_7159);
xor U10223 (N_10223,N_2856,N_1331);
nand U10224 (N_10224,N_9758,N_6373);
nor U10225 (N_10225,N_6512,N_8528);
xnor U10226 (N_10226,N_1525,N_9070);
nor U10227 (N_10227,N_5483,N_5270);
or U10228 (N_10228,N_1648,N_5216);
xnor U10229 (N_10229,N_8188,N_9245);
and U10230 (N_10230,N_3176,N_2548);
or U10231 (N_10231,N_6877,N_7907);
xor U10232 (N_10232,N_3513,N_5113);
xnor U10233 (N_10233,N_4086,N_1112);
nor U10234 (N_10234,N_7112,N_9476);
and U10235 (N_10235,N_2759,N_9410);
nor U10236 (N_10236,N_8041,N_1011);
nor U10237 (N_10237,N_9806,N_1913);
xnor U10238 (N_10238,N_2439,N_7984);
or U10239 (N_10239,N_2674,N_3163);
nand U10240 (N_10240,N_4418,N_2907);
or U10241 (N_10241,N_4113,N_2317);
or U10242 (N_10242,N_2732,N_6013);
or U10243 (N_10243,N_7259,N_6747);
nand U10244 (N_10244,N_271,N_5421);
and U10245 (N_10245,N_8556,N_2);
and U10246 (N_10246,N_3687,N_3588);
nand U10247 (N_10247,N_2026,N_979);
and U10248 (N_10248,N_1510,N_8140);
or U10249 (N_10249,N_9985,N_6515);
nand U10250 (N_10250,N_2924,N_6578);
nor U10251 (N_10251,N_3429,N_9799);
xor U10252 (N_10252,N_8840,N_37);
or U10253 (N_10253,N_1845,N_2583);
and U10254 (N_10254,N_2402,N_1955);
xor U10255 (N_10255,N_4980,N_6622);
and U10256 (N_10256,N_9280,N_1554);
xor U10257 (N_10257,N_4129,N_253);
nand U10258 (N_10258,N_6884,N_8271);
xor U10259 (N_10259,N_4957,N_976);
xnor U10260 (N_10260,N_3215,N_6416);
xor U10261 (N_10261,N_6565,N_1228);
nor U10262 (N_10262,N_2415,N_8298);
nand U10263 (N_10263,N_7441,N_3074);
and U10264 (N_10264,N_1557,N_1212);
and U10265 (N_10265,N_1184,N_8847);
or U10266 (N_10266,N_4582,N_6859);
xnor U10267 (N_10267,N_573,N_281);
and U10268 (N_10268,N_2940,N_3772);
or U10269 (N_10269,N_6658,N_8053);
nand U10270 (N_10270,N_8459,N_9513);
xor U10271 (N_10271,N_1884,N_6254);
nor U10272 (N_10272,N_7297,N_2777);
or U10273 (N_10273,N_8913,N_1771);
or U10274 (N_10274,N_5240,N_1051);
and U10275 (N_10275,N_1974,N_438);
xor U10276 (N_10276,N_8922,N_7388);
nand U10277 (N_10277,N_4647,N_2915);
or U10278 (N_10278,N_1917,N_7180);
nand U10279 (N_10279,N_3676,N_9271);
and U10280 (N_10280,N_4130,N_5545);
or U10281 (N_10281,N_824,N_9937);
xnor U10282 (N_10282,N_6155,N_5267);
nor U10283 (N_10283,N_5936,N_923);
nand U10284 (N_10284,N_9750,N_9068);
nand U10285 (N_10285,N_3958,N_6946);
or U10286 (N_10286,N_7584,N_6394);
and U10287 (N_10287,N_8460,N_288);
nand U10288 (N_10288,N_2191,N_8354);
nor U10289 (N_10289,N_2136,N_9186);
and U10290 (N_10290,N_1138,N_7786);
xor U10291 (N_10291,N_9172,N_2701);
nand U10292 (N_10292,N_9317,N_2094);
nand U10293 (N_10293,N_9845,N_2315);
xor U10294 (N_10294,N_4305,N_1704);
nand U10295 (N_10295,N_9965,N_7224);
nor U10296 (N_10296,N_1538,N_5842);
and U10297 (N_10297,N_1672,N_7132);
nand U10298 (N_10298,N_7734,N_5220);
nand U10299 (N_10299,N_1305,N_6299);
and U10300 (N_10300,N_5386,N_6491);
nand U10301 (N_10301,N_1876,N_1513);
nor U10302 (N_10302,N_7554,N_7824);
nand U10303 (N_10303,N_7700,N_6315);
nand U10304 (N_10304,N_1976,N_9878);
nand U10305 (N_10305,N_8424,N_9007);
or U10306 (N_10306,N_5769,N_7604);
xor U10307 (N_10307,N_9855,N_5832);
or U10308 (N_10308,N_2746,N_1202);
or U10309 (N_10309,N_9136,N_6713);
xor U10310 (N_10310,N_2427,N_5670);
nor U10311 (N_10311,N_9605,N_2846);
xor U10312 (N_10312,N_7679,N_1230);
nand U10313 (N_10313,N_1218,N_4247);
xnor U10314 (N_10314,N_8426,N_1666);
nor U10315 (N_10315,N_1155,N_4295);
and U10316 (N_10316,N_7145,N_1208);
xor U10317 (N_10317,N_3525,N_1392);
and U10318 (N_10318,N_6592,N_4607);
or U10319 (N_10319,N_3151,N_2065);
and U10320 (N_10320,N_798,N_6112);
nand U10321 (N_10321,N_4698,N_9060);
xor U10322 (N_10322,N_954,N_4850);
xor U10323 (N_10323,N_1787,N_4238);
and U10324 (N_10324,N_4608,N_9600);
xor U10325 (N_10325,N_4896,N_1741);
xor U10326 (N_10326,N_5063,N_7702);
nand U10327 (N_10327,N_2188,N_7938);
nand U10328 (N_10328,N_1980,N_3787);
or U10329 (N_10329,N_2577,N_5687);
nor U10330 (N_10330,N_2567,N_8496);
xor U10331 (N_10331,N_5087,N_7458);
nand U10332 (N_10332,N_7399,N_7477);
nor U10333 (N_10333,N_8253,N_4603);
xnor U10334 (N_10334,N_8112,N_355);
and U10335 (N_10335,N_8713,N_9900);
and U10336 (N_10336,N_1161,N_3785);
or U10337 (N_10337,N_4520,N_8531);
and U10338 (N_10338,N_2914,N_7539);
or U10339 (N_10339,N_7121,N_4860);
nand U10340 (N_10340,N_1217,N_6370);
xor U10341 (N_10341,N_5084,N_8307);
or U10342 (N_10342,N_9211,N_6114);
nand U10343 (N_10343,N_8351,N_2649);
nand U10344 (N_10344,N_5708,N_417);
xnor U10345 (N_10345,N_8139,N_6992);
and U10346 (N_10346,N_8826,N_7941);
xor U10347 (N_10347,N_344,N_2098);
and U10348 (N_10348,N_321,N_4196);
or U10349 (N_10349,N_2983,N_7064);
nand U10350 (N_10350,N_1361,N_4413);
and U10351 (N_10351,N_6393,N_2035);
nor U10352 (N_10352,N_6959,N_3518);
nor U10353 (N_10353,N_4661,N_56);
or U10354 (N_10354,N_7451,N_6177);
or U10355 (N_10355,N_5838,N_1579);
xnor U10356 (N_10356,N_1086,N_7024);
and U10357 (N_10357,N_4627,N_8048);
nor U10358 (N_10358,N_6973,N_2876);
nand U10359 (N_10359,N_1162,N_3763);
and U10360 (N_10360,N_1970,N_9946);
or U10361 (N_10361,N_3127,N_9689);
or U10362 (N_10362,N_6892,N_4399);
xor U10363 (N_10363,N_1559,N_8329);
or U10364 (N_10364,N_9313,N_1378);
nand U10365 (N_10365,N_8313,N_8050);
or U10366 (N_10366,N_6548,N_6509);
nand U10367 (N_10367,N_9113,N_3521);
and U10368 (N_10368,N_4108,N_6615);
nor U10369 (N_10369,N_3533,N_6849);
nand U10370 (N_10370,N_7350,N_4380);
nor U10371 (N_10371,N_9990,N_34);
and U10372 (N_10372,N_8422,N_2380);
or U10373 (N_10373,N_4682,N_2792);
nand U10374 (N_10374,N_4242,N_4970);
or U10375 (N_10375,N_8983,N_7994);
xnor U10376 (N_10376,N_7245,N_8391);
nor U10377 (N_10377,N_9371,N_2390);
and U10378 (N_10378,N_8002,N_4781);
nand U10379 (N_10379,N_5138,N_4960);
nand U10380 (N_10380,N_8262,N_7768);
nand U10381 (N_10381,N_9676,N_1567);
nand U10382 (N_10382,N_2625,N_2156);
and U10383 (N_10383,N_8989,N_8707);
and U10384 (N_10384,N_2917,N_6381);
nand U10385 (N_10385,N_9559,N_3760);
nand U10386 (N_10386,N_814,N_2363);
and U10387 (N_10387,N_4574,N_2269);
or U10388 (N_10388,N_9819,N_9715);
nand U10389 (N_10389,N_2698,N_3956);
xor U10390 (N_10390,N_5564,N_8571);
and U10391 (N_10391,N_562,N_6150);
nand U10392 (N_10392,N_875,N_7961);
nor U10393 (N_10393,N_9368,N_4874);
or U10394 (N_10394,N_832,N_5436);
xnor U10395 (N_10395,N_8465,N_7534);
and U10396 (N_10396,N_996,N_3870);
nand U10397 (N_10397,N_1571,N_7383);
nand U10398 (N_10398,N_2096,N_3170);
xnor U10399 (N_10399,N_5364,N_6810);
nand U10400 (N_10400,N_5896,N_6938);
xnor U10401 (N_10401,N_3472,N_9415);
xor U10402 (N_10402,N_7535,N_7705);
nor U10403 (N_10403,N_4341,N_2736);
nand U10404 (N_10404,N_2909,N_1546);
nor U10405 (N_10405,N_6262,N_9585);
nand U10406 (N_10406,N_2538,N_5655);
xnor U10407 (N_10407,N_6412,N_8615);
nand U10408 (N_10408,N_1150,N_1183);
or U10409 (N_10409,N_2639,N_8028);
nand U10410 (N_10410,N_4141,N_9685);
or U10411 (N_10411,N_4105,N_9144);
nor U10412 (N_10412,N_6572,N_1432);
and U10413 (N_10413,N_8728,N_192);
nand U10414 (N_10414,N_6925,N_1670);
xor U10415 (N_10415,N_9408,N_7710);
nand U10416 (N_10416,N_9777,N_8256);
nor U10417 (N_10417,N_1404,N_807);
nand U10418 (N_10418,N_9756,N_8032);
and U10419 (N_10419,N_460,N_5762);
nor U10420 (N_10420,N_4004,N_6953);
nor U10421 (N_10421,N_4050,N_2257);
xor U10422 (N_10422,N_9805,N_7086);
or U10423 (N_10423,N_7853,N_3360);
and U10424 (N_10424,N_4577,N_7688);
nor U10425 (N_10425,N_5924,N_205);
xor U10426 (N_10426,N_9887,N_607);
and U10427 (N_10427,N_3375,N_6439);
nor U10428 (N_10428,N_7828,N_4535);
and U10429 (N_10429,N_9447,N_2611);
nor U10430 (N_10430,N_370,N_2962);
xnor U10431 (N_10431,N_5653,N_6066);
nand U10432 (N_10432,N_7730,N_9964);
xor U10433 (N_10433,N_3953,N_6487);
or U10434 (N_10434,N_2082,N_4266);
xor U10435 (N_10435,N_2000,N_2011);
or U10436 (N_10436,N_7432,N_4324);
nor U10437 (N_10437,N_8210,N_9491);
and U10438 (N_10438,N_5725,N_7678);
xnor U10439 (N_10439,N_5373,N_5365);
and U10440 (N_10440,N_9344,N_1780);
nor U10441 (N_10441,N_4111,N_3043);
xnor U10442 (N_10442,N_1790,N_2197);
or U10443 (N_10443,N_2357,N_7716);
or U10444 (N_10444,N_9794,N_2287);
nor U10445 (N_10445,N_854,N_7014);
and U10446 (N_10446,N_3606,N_1744);
nand U10447 (N_10447,N_3541,N_8437);
nand U10448 (N_10448,N_4873,N_8903);
and U10449 (N_10449,N_2165,N_1939);
or U10450 (N_10450,N_6554,N_7067);
and U10451 (N_10451,N_3324,N_4074);
and U10452 (N_10452,N_6268,N_6672);
and U10453 (N_10453,N_9987,N_3598);
nand U10454 (N_10454,N_8887,N_6014);
or U10455 (N_10455,N_4134,N_3317);
xnor U10456 (N_10456,N_6486,N_5486);
xnor U10457 (N_10457,N_7848,N_4033);
and U10458 (N_10458,N_3589,N_147);
nand U10459 (N_10459,N_4954,N_4529);
nor U10460 (N_10460,N_4264,N_9541);
nand U10461 (N_10461,N_2470,N_5967);
or U10462 (N_10462,N_8830,N_1114);
and U10463 (N_10463,N_2050,N_1069);
or U10464 (N_10464,N_9620,N_3268);
xor U10465 (N_10465,N_808,N_4796);
nor U10466 (N_10466,N_3115,N_575);
nor U10467 (N_10467,N_7407,N_799);
xnor U10468 (N_10468,N_1413,N_794);
xnor U10469 (N_10469,N_1948,N_5484);
and U10470 (N_10470,N_2479,N_4376);
xor U10471 (N_10471,N_6540,N_4940);
nand U10472 (N_10472,N_9956,N_2070);
xnor U10473 (N_10473,N_4830,N_1943);
nor U10474 (N_10474,N_8000,N_296);
and U10475 (N_10475,N_1462,N_8120);
nand U10476 (N_10476,N_713,N_1921);
and U10477 (N_10477,N_5970,N_3766);
xor U10478 (N_10478,N_3454,N_677);
or U10479 (N_10479,N_1085,N_7830);
nand U10480 (N_10480,N_8229,N_6036);
or U10481 (N_10481,N_999,N_455);
nor U10482 (N_10482,N_9957,N_3641);
and U10483 (N_10483,N_8818,N_9128);
nand U10484 (N_10484,N_8463,N_6105);
or U10485 (N_10485,N_5662,N_8125);
nor U10486 (N_10486,N_1030,N_3212);
nor U10487 (N_10487,N_6494,N_1665);
or U10488 (N_10488,N_7803,N_495);
xnor U10489 (N_10489,N_2116,N_3818);
and U10490 (N_10490,N_5097,N_190);
and U10491 (N_10491,N_970,N_7273);
nand U10492 (N_10492,N_1128,N_8106);
and U10493 (N_10493,N_7105,N_577);
and U10494 (N_10494,N_1926,N_7708);
and U10495 (N_10495,N_4065,N_9812);
xnor U10496 (N_10496,N_2291,N_4572);
or U10497 (N_10497,N_7378,N_4838);
xnor U10498 (N_10498,N_8580,N_4763);
xor U10499 (N_10499,N_7389,N_3270);
nor U10500 (N_10500,N_7082,N_7091);
nor U10501 (N_10501,N_3885,N_6496);
or U10502 (N_10502,N_4326,N_8619);
or U10503 (N_10503,N_9445,N_3523);
or U10504 (N_10504,N_2273,N_6530);
and U10505 (N_10505,N_7033,N_8532);
nand U10506 (N_10506,N_4314,N_3933);
or U10507 (N_10507,N_1687,N_4826);
nand U10508 (N_10508,N_3964,N_1066);
and U10509 (N_10509,N_8850,N_9303);
or U10510 (N_10510,N_4340,N_5799);
or U10511 (N_10511,N_5172,N_516);
or U10512 (N_10512,N_1187,N_6519);
nand U10513 (N_10513,N_4753,N_2781);
xor U10514 (N_10514,N_4128,N_1616);
and U10515 (N_10515,N_9481,N_5606);
nand U10516 (N_10516,N_7989,N_7760);
xor U10517 (N_10517,N_6081,N_5010);
or U10518 (N_10518,N_1828,N_3459);
nand U10519 (N_10519,N_1297,N_7156);
nor U10520 (N_10520,N_9835,N_3250);
nand U10521 (N_10521,N_2835,N_4383);
xor U10522 (N_10522,N_9020,N_2615);
nand U10523 (N_10523,N_8523,N_8828);
and U10524 (N_10524,N_4472,N_9785);
xnor U10525 (N_10525,N_2320,N_3136);
nand U10526 (N_10526,N_47,N_7170);
nand U10527 (N_10527,N_1748,N_6893);
or U10528 (N_10528,N_2483,N_149);
xor U10529 (N_10529,N_5114,N_8655);
nand U10530 (N_10530,N_7856,N_7392);
and U10531 (N_10531,N_1637,N_8607);
or U10532 (N_10532,N_6827,N_4207);
xor U10533 (N_10533,N_6321,N_6806);
or U10534 (N_10534,N_7507,N_5403);
nor U10535 (N_10535,N_3678,N_5493);
xor U10536 (N_10536,N_8730,N_680);
nor U10537 (N_10537,N_1663,N_2401);
xnor U10538 (N_10538,N_5599,N_4419);
or U10539 (N_10539,N_494,N_8658);
nand U10540 (N_10540,N_4289,N_1826);
xor U10541 (N_10541,N_2466,N_5544);
nand U10542 (N_10542,N_3814,N_7168);
and U10543 (N_10543,N_4076,N_3394);
nand U10544 (N_10544,N_2594,N_5786);
nand U10545 (N_10545,N_5567,N_5446);
nor U10546 (N_10546,N_4833,N_4724);
nor U10547 (N_10547,N_1871,N_7010);
or U10548 (N_10548,N_8738,N_544);
or U10549 (N_10549,N_9192,N_9182);
nand U10550 (N_10550,N_4566,N_9528);
and U10551 (N_10551,N_8795,N_5943);
or U10552 (N_10552,N_1189,N_6525);
nand U10553 (N_10553,N_4772,N_1733);
xor U10554 (N_10554,N_7552,N_754);
nor U10555 (N_10555,N_1799,N_5837);
nand U10556 (N_10556,N_9421,N_7636);
or U10557 (N_10557,N_5579,N_7408);
xor U10558 (N_10558,N_8588,N_4423);
and U10559 (N_10559,N_6733,N_8926);
or U10560 (N_10560,N_9230,N_5348);
or U10561 (N_10561,N_8827,N_6922);
xnor U10562 (N_10562,N_1860,N_8949);
or U10563 (N_10563,N_9959,N_9197);
nor U10564 (N_10564,N_3592,N_1177);
nand U10565 (N_10565,N_1389,N_9279);
and U10566 (N_10566,N_4776,N_4506);
nand U10567 (N_10567,N_2808,N_9889);
nor U10568 (N_10568,N_9325,N_8353);
nand U10569 (N_10569,N_5956,N_8806);
or U10570 (N_10570,N_7195,N_4735);
xor U10571 (N_10571,N_3244,N_4415);
xnor U10572 (N_10572,N_6325,N_6976);
or U10573 (N_10573,N_4568,N_6260);
and U10574 (N_10574,N_3542,N_5511);
nand U10575 (N_10575,N_3677,N_6564);
and U10576 (N_10576,N_3622,N_3398);
nor U10577 (N_10577,N_6497,N_3011);
or U10578 (N_10578,N_784,N_1959);
xnor U10579 (N_10579,N_3034,N_4053);
and U10580 (N_10580,N_8561,N_9078);
xor U10581 (N_10581,N_7594,N_8614);
and U10582 (N_10582,N_5987,N_4750);
and U10583 (N_10583,N_1625,N_4919);
nand U10584 (N_10584,N_8374,N_4160);
nand U10585 (N_10585,N_9059,N_3483);
nand U10586 (N_10586,N_3377,N_9343);
or U10587 (N_10587,N_382,N_8551);
nand U10588 (N_10588,N_8290,N_3897);
nand U10589 (N_10589,N_8813,N_2480);
or U10590 (N_10590,N_2100,N_5372);
xor U10591 (N_10591,N_9100,N_3628);
nor U10592 (N_10592,N_5696,N_153);
nand U10593 (N_10593,N_2182,N_7204);
and U10594 (N_10594,N_6522,N_5342);
xnor U10595 (N_10595,N_2522,N_8570);
nand U10596 (N_10596,N_3880,N_847);
nand U10597 (N_10597,N_723,N_9630);
nand U10598 (N_10598,N_9073,N_8954);
xnor U10599 (N_10599,N_4888,N_5808);
nand U10600 (N_10600,N_2361,N_2738);
nor U10601 (N_10601,N_7592,N_6348);
xnor U10602 (N_10602,N_4268,N_2484);
nand U10603 (N_10603,N_373,N_2650);
or U10604 (N_10604,N_1835,N_1558);
xnor U10605 (N_10605,N_4813,N_9748);
xnor U10606 (N_10606,N_9108,N_1175);
nand U10607 (N_10607,N_3556,N_9288);
nor U10608 (N_10608,N_8471,N_7235);
and U10609 (N_10609,N_2652,N_2885);
xnor U10610 (N_10610,N_7081,N_1543);
xor U10611 (N_10611,N_3931,N_6516);
xnor U10612 (N_10612,N_3828,N_827);
or U10613 (N_10613,N_6237,N_8065);
xnor U10614 (N_10614,N_3386,N_1041);
or U10615 (N_10615,N_1534,N_2827);
nor U10616 (N_10616,N_6184,N_7426);
nand U10617 (N_10617,N_5843,N_4931);
xnor U10618 (N_10618,N_4617,N_6347);
xor U10619 (N_10619,N_830,N_5425);
nor U10620 (N_10620,N_5341,N_9416);
or U10621 (N_10621,N_5962,N_9869);
and U10622 (N_10622,N_2954,N_2656);
xor U10623 (N_10623,N_6895,N_9668);
nor U10624 (N_10624,N_697,N_2271);
nor U10625 (N_10625,N_8335,N_4106);
nor U10626 (N_10626,N_9531,N_7667);
nor U10627 (N_10627,N_3659,N_8963);
xor U10628 (N_10628,N_9854,N_6694);
xnor U10629 (N_10629,N_6505,N_9738);
nand U10630 (N_10630,N_3704,N_506);
nor U10631 (N_10631,N_8392,N_583);
nand U10632 (N_10632,N_839,N_7062);
nand U10633 (N_10633,N_6696,N_7034);
nand U10634 (N_10634,N_7006,N_2298);
nor U10635 (N_10635,N_2149,N_1009);
nand U10636 (N_10636,N_5385,N_5909);
nor U10637 (N_10637,N_5983,N_2778);
and U10638 (N_10638,N_3451,N_5495);
nor U10639 (N_10639,N_1702,N_7766);
nor U10640 (N_10640,N_9083,N_3469);
nand U10641 (N_10641,N_2831,N_7751);
nor U10642 (N_10642,N_8825,N_3050);
nand U10643 (N_10643,N_1427,N_4771);
nand U10644 (N_10644,N_2171,N_4640);
and U10645 (N_10645,N_721,N_6135);
and U10646 (N_10646,N_1332,N_1196);
nor U10647 (N_10647,N_7197,N_7543);
and U10648 (N_10648,N_1730,N_5015);
nor U10649 (N_10649,N_6056,N_8583);
and U10650 (N_10650,N_7516,N_5833);
or U10651 (N_10651,N_5266,N_9857);
nand U10652 (N_10652,N_7437,N_4800);
or U10653 (N_10653,N_1257,N_8155);
xnor U10654 (N_10654,N_463,N_5035);
nand U10655 (N_10655,N_2030,N_7825);
and U10656 (N_10656,N_9731,N_9565);
and U10657 (N_10657,N_4241,N_8714);
and U10658 (N_10658,N_5088,N_491);
xor U10659 (N_10659,N_574,N_6912);
or U10660 (N_10660,N_679,N_2762);
or U10661 (N_10661,N_179,N_5997);
xnor U10662 (N_10662,N_5419,N_3473);
and U10663 (N_10663,N_5654,N_2855);
nor U10664 (N_10664,N_229,N_8481);
nand U10665 (N_10665,N_8652,N_7550);
nand U10666 (N_10666,N_3630,N_9832);
or U10667 (N_10667,N_1599,N_9143);
xor U10668 (N_10668,N_2965,N_1800);
or U10669 (N_10669,N_6476,N_6332);
xor U10670 (N_10670,N_7831,N_5733);
and U10671 (N_10671,N_480,N_3369);
or U10672 (N_10672,N_1283,N_4210);
or U10673 (N_10673,N_3373,N_2566);
or U10674 (N_10674,N_2532,N_184);
xor U10675 (N_10675,N_2558,N_1689);
and U10676 (N_10676,N_7052,N_9190);
xor U10677 (N_10677,N_1831,N_5831);
nand U10678 (N_10678,N_7977,N_1363);
nor U10679 (N_10679,N_159,N_2871);
xor U10680 (N_10680,N_2218,N_6455);
nand U10681 (N_10681,N_4274,N_6574);
nand U10682 (N_10682,N_3832,N_6454);
nand U10683 (N_10683,N_5750,N_8425);
nand U10684 (N_10684,N_3522,N_3493);
xor U10685 (N_10685,N_8988,N_1515);
or U10686 (N_10686,N_7868,N_5390);
or U10687 (N_10687,N_3564,N_5908);
nor U10688 (N_10688,N_4503,N_6188);
xnor U10689 (N_10689,N_9283,N_7548);
and U10690 (N_10690,N_6094,N_3495);
and U10691 (N_10691,N_5328,N_7732);
nor U10692 (N_10692,N_9769,N_9159);
nor U10693 (N_10693,N_4459,N_1635);
nand U10694 (N_10694,N_1581,N_422);
or U10695 (N_10695,N_9398,N_457);
nand U10696 (N_10696,N_3477,N_7812);
xnor U10697 (N_10697,N_9989,N_5064);
or U10698 (N_10698,N_2372,N_6278);
nand U10699 (N_10699,N_383,N_634);
or U10700 (N_10700,N_732,N_3936);
nor U10701 (N_10701,N_1487,N_9874);
or U10702 (N_10702,N_6214,N_5078);
nor U10703 (N_10703,N_4188,N_3731);
and U10704 (N_10704,N_3924,N_1673);
nand U10705 (N_10705,N_9744,N_9400);
nand U10706 (N_10706,N_4442,N_8750);
nor U10707 (N_10707,N_371,N_4453);
or U10708 (N_10708,N_6205,N_5783);
nand U10709 (N_10709,N_1447,N_643);
xor U10710 (N_10710,N_187,N_6712);
and U10711 (N_10711,N_9762,N_3925);
or U10712 (N_10712,N_6460,N_8945);
nand U10713 (N_10713,N_446,N_7761);
nor U10714 (N_10714,N_9858,N_8756);
nor U10715 (N_10715,N_5362,N_4497);
and U10716 (N_10716,N_8096,N_9203);
nand U10717 (N_10717,N_7454,N_4350);
or U10718 (N_10718,N_8040,N_2680);
xor U10719 (N_10719,N_6201,N_1881);
xnor U10720 (N_10720,N_3757,N_2552);
and U10721 (N_10721,N_4963,N_7916);
and U10722 (N_10722,N_9222,N_8202);
or U10723 (N_10723,N_2720,N_4473);
and U10724 (N_10724,N_8539,N_4403);
or U10725 (N_10725,N_1776,N_2419);
and U10726 (N_10726,N_9573,N_1919);
and U10727 (N_10727,N_4110,N_8578);
nand U10728 (N_10728,N_2840,N_318);
and U10729 (N_10729,N_535,N_726);
nand U10730 (N_10730,N_6250,N_9945);
xnor U10731 (N_10731,N_7084,N_1726);
xor U10732 (N_10732,N_9026,N_4523);
nand U10733 (N_10733,N_2139,N_3871);
nand U10734 (N_10734,N_6372,N_4091);
or U10735 (N_10735,N_483,N_8251);
xor U10736 (N_10736,N_9653,N_5590);
nand U10737 (N_10737,N_3333,N_5637);
or U10738 (N_10738,N_3788,N_4900);
xnor U10739 (N_10739,N_4966,N_3062);
xnor U10740 (N_10740,N_2010,N_740);
and U10741 (N_10741,N_7249,N_3855);
nor U10742 (N_10742,N_8624,N_255);
nand U10743 (N_10743,N_9521,N_9935);
xnor U10744 (N_10744,N_5331,N_7965);
nor U10745 (N_10745,N_4959,N_4131);
and U10746 (N_10746,N_2167,N_2436);
or U10747 (N_10747,N_8950,N_8346);
or U10748 (N_10748,N_9464,N_9069);
or U10749 (N_10749,N_2892,N_6298);
or U10750 (N_10750,N_1912,N_599);
nand U10751 (N_10751,N_1686,N_7090);
or U10752 (N_10752,N_1176,N_503);
nor U10753 (N_10753,N_5770,N_2841);
nor U10754 (N_10754,N_8734,N_2972);
nand U10755 (N_10755,N_2925,N_7274);
xor U10756 (N_10756,N_8783,N_2832);
and U10757 (N_10757,N_1053,N_6545);
or U10758 (N_10758,N_9908,N_9241);
xnor U10759 (N_10759,N_8181,N_4790);
xnor U10760 (N_10760,N_8414,N_3655);
nor U10761 (N_10761,N_3194,N_6071);
and U10762 (N_10762,N_3707,N_5415);
xor U10763 (N_10763,N_7357,N_5881);
nand U10764 (N_10764,N_2332,N_9135);
and U10765 (N_10765,N_9112,N_5198);
and U10766 (N_10766,N_7153,N_8340);
or U10767 (N_10767,N_5041,N_6706);
xnor U10768 (N_10768,N_1125,N_4986);
nand U10769 (N_10769,N_6805,N_4573);
nand U10770 (N_10770,N_1505,N_6316);
or U10771 (N_10771,N_2170,N_2694);
xnor U10772 (N_10772,N_7402,N_5408);
nand U10773 (N_10773,N_5632,N_7374);
and U10774 (N_10774,N_7954,N_8260);
or U10775 (N_10775,N_9240,N_9962);
nand U10776 (N_10776,N_6283,N_1719);
xor U10777 (N_10777,N_8081,N_1829);
nor U10778 (N_10778,N_3029,N_7703);
and U10779 (N_10779,N_2729,N_4759);
nor U10780 (N_10780,N_5081,N_3735);
or U10781 (N_10781,N_8123,N_7649);
nor U10782 (N_10782,N_52,N_4528);
nor U10783 (N_10783,N_8855,N_1292);
and U10784 (N_10784,N_7656,N_3727);
or U10785 (N_10785,N_4244,N_7890);
and U10786 (N_10786,N_6789,N_9176);
nor U10787 (N_10787,N_2462,N_5490);
nand U10788 (N_10788,N_2794,N_8821);
xnor U10789 (N_10789,N_8147,N_6808);
nor U10790 (N_10790,N_2243,N_7817);
and U10791 (N_10791,N_2659,N_2666);
and U10792 (N_10792,N_3593,N_8344);
xnor U10793 (N_10793,N_7030,N_917);
or U10794 (N_10794,N_4235,N_1713);
nand U10795 (N_10795,N_3605,N_8520);
and U10796 (N_10796,N_3101,N_9008);
nand U10797 (N_10797,N_4409,N_2459);
xnor U10798 (N_10798,N_16,N_2718);
nand U10799 (N_10799,N_5631,N_4217);
and U10800 (N_10800,N_3171,N_582);
nor U10801 (N_10801,N_6855,N_9788);
nor U10802 (N_10802,N_8628,N_2630);
or U10803 (N_10803,N_6573,N_9027);
nor U10804 (N_10804,N_103,N_719);
nor U10805 (N_10805,N_5101,N_868);
or U10806 (N_10806,N_572,N_659);
and U10807 (N_10807,N_4023,N_9285);
xor U10808 (N_10808,N_9710,N_7261);
nand U10809 (N_10809,N_2241,N_7813);
xor U10810 (N_10810,N_5434,N_7017);
nor U10811 (N_10811,N_9348,N_8549);
xor U10812 (N_10812,N_4254,N_4225);
or U10813 (N_10813,N_7875,N_5656);
nand U10814 (N_10814,N_1451,N_6942);
xor U10815 (N_10815,N_9014,N_9358);
and U10816 (N_10816,N_1533,N_197);
or U10817 (N_10817,N_2935,N_8055);
nor U10818 (N_10818,N_6041,N_2916);
and U10819 (N_10819,N_8357,N_3213);
nor U10820 (N_10820,N_3272,N_7363);
xor U10821 (N_10821,N_3698,N_6088);
nand U10822 (N_10822,N_6478,N_4375);
nand U10823 (N_10823,N_8912,N_8719);
xor U10824 (N_10824,N_4257,N_7097);
or U10825 (N_10825,N_7859,N_2516);
nand U10826 (N_10826,N_5002,N_1307);
xnor U10827 (N_10827,N_6142,N_9019);
or U10828 (N_10828,N_2398,N_5461);
and U10829 (N_10829,N_7329,N_9305);
or U10830 (N_10830,N_4321,N_8567);
and U10831 (N_10831,N_7323,N_1570);
and U10832 (N_10832,N_4621,N_2041);
and U10833 (N_10833,N_8533,N_5893);
nand U10834 (N_10834,N_7527,N_5339);
nand U10835 (N_10835,N_8102,N_8565);
or U10836 (N_10836,N_4905,N_8100);
nand U10837 (N_10837,N_3941,N_9138);
nor U10838 (N_10838,N_880,N_2849);
nand U10839 (N_10839,N_1752,N_3387);
and U10840 (N_10840,N_3649,N_1440);
nor U10841 (N_10841,N_4618,N_4811);
and U10842 (N_10842,N_997,N_1679);
xor U10843 (N_10843,N_8068,N_9490);
nor U10844 (N_10844,N_9686,N_800);
and U10845 (N_10845,N_8566,N_7488);
xnor U10846 (N_10846,N_8979,N_5208);
or U10847 (N_10847,N_9470,N_2224);
or U10848 (N_10848,N_8858,N_1029);
xor U10849 (N_10849,N_4493,N_4149);
or U10850 (N_10850,N_5374,N_5629);
or U10851 (N_10851,N_3041,N_6432);
nor U10852 (N_10852,N_7326,N_2531);
and U10853 (N_10853,N_1727,N_8920);
nand U10854 (N_10854,N_5132,N_5334);
xor U10855 (N_10855,N_6826,N_7008);
nand U10856 (N_10856,N_7237,N_2111);
nor U10857 (N_10857,N_1645,N_3012);
xnor U10858 (N_10858,N_9252,N_44);
nand U10859 (N_10859,N_2400,N_7635);
nor U10860 (N_10860,N_7560,N_6790);
xnor U10861 (N_10861,N_4628,N_4322);
nand U10862 (N_10862,N_8720,N_7131);
nand U10863 (N_10863,N_5507,N_4637);
nor U10864 (N_10864,N_1947,N_6499);
or U10865 (N_10865,N_3550,N_6586);
nor U10866 (N_10866,N_725,N_3471);
nand U10867 (N_10867,N_5311,N_305);
or U10868 (N_10868,N_1439,N_5819);
nand U10869 (N_10869,N_410,N_8314);
xor U10870 (N_10870,N_5804,N_4190);
or U10871 (N_10871,N_2491,N_1074);
and U10872 (N_10872,N_8675,N_8668);
or U10873 (N_10873,N_2346,N_8792);
nor U10874 (N_10874,N_6837,N_7919);
and U10875 (N_10875,N_155,N_501);
nand U10876 (N_10876,N_6524,N_9404);
xnor U10877 (N_10877,N_7928,N_2057);
and U10878 (N_10878,N_3411,N_7136);
nor U10879 (N_10879,N_3150,N_7355);
or U10880 (N_10880,N_9713,N_8812);
nand U10881 (N_10881,N_8516,N_1690);
nand U10882 (N_10882,N_5004,N_9894);
or U10883 (N_10883,N_166,N_4545);
nor U10884 (N_10884,N_219,N_7613);
xnor U10885 (N_10885,N_5959,N_6266);
or U10886 (N_10886,N_8574,N_7193);
nand U10887 (N_10887,N_4422,N_7682);
or U10888 (N_10888,N_418,N_3201);
nand U10889 (N_10889,N_1181,N_1068);
or U10890 (N_10890,N_6011,N_7191);
nand U10891 (N_10891,N_8308,N_8427);
xnor U10892 (N_10892,N_9782,N_982);
xor U10893 (N_10893,N_1796,N_6553);
nand U10894 (N_10894,N_9910,N_6956);
xnor U10895 (N_10895,N_8444,N_4993);
xor U10896 (N_10896,N_3085,N_2121);
or U10897 (N_10897,N_7680,N_3129);
nand U10898 (N_10898,N_4041,N_5128);
nand U10899 (N_10899,N_3879,N_1937);
and U10900 (N_10900,N_380,N_9526);
and U10901 (N_10901,N_9591,N_9351);
and U10902 (N_10902,N_8494,N_225);
and U10903 (N_10903,N_7429,N_8593);
and U10904 (N_10904,N_8497,N_8705);
nor U10905 (N_10905,N_1367,N_7157);
and U10906 (N_10906,N_9009,N_6368);
and U10907 (N_10907,N_5566,N_7489);
nand U10908 (N_10908,N_4536,N_5134);
nor U10909 (N_10909,N_4822,N_9354);
or U10910 (N_10910,N_3614,N_3368);
nor U10911 (N_10911,N_4868,N_5955);
nor U10912 (N_10912,N_9347,N_7841);
xnor U10913 (N_10913,N_2752,N_2455);
and U10914 (N_10914,N_3752,N_275);
nand U10915 (N_10915,N_4842,N_6062);
or U10916 (N_10916,N_43,N_4175);
xor U10917 (N_10917,N_585,N_1103);
nand U10918 (N_10918,N_7918,N_6123);
nor U10919 (N_10919,N_1522,N_8020);
nor U10920 (N_10920,N_2048,N_2403);
or U10921 (N_10921,N_5999,N_8754);
nor U10922 (N_10922,N_9789,N_675);
and U10923 (N_10923,N_6384,N_1814);
xnor U10924 (N_10924,N_6042,N_720);
or U10925 (N_10925,N_5701,N_2877);
and U10926 (N_10926,N_4112,N_7466);
nand U10927 (N_10927,N_7740,N_5512);
nand U10928 (N_10928,N_5301,N_9754);
nand U10929 (N_10929,N_2276,N_962);
and U10930 (N_10930,N_3974,N_935);
nor U10931 (N_10931,N_5573,N_8373);
and U10932 (N_10932,N_3067,N_1808);
nor U10933 (N_10933,N_3674,N_9039);
nand U10934 (N_10934,N_9133,N_2987);
xor U10935 (N_10935,N_9057,N_8591);
and U10936 (N_10936,N_6754,N_4416);
and U10937 (N_10937,N_1677,N_354);
or U10938 (N_10938,N_164,N_6730);
and U10939 (N_10939,N_3852,N_6032);
nand U10940 (N_10940,N_8191,N_2882);
nand U10941 (N_10941,N_3904,N_4590);
and U10942 (N_10942,N_7588,N_1284);
or U10943 (N_10943,N_4307,N_257);
and U10944 (N_10944,N_3193,N_4102);
xnor U10945 (N_10945,N_1236,N_7851);
xnor U10946 (N_10946,N_727,N_6128);
nand U10947 (N_10947,N_7647,N_1371);
nand U10948 (N_10948,N_7262,N_8248);
and U10949 (N_10949,N_320,N_8215);
and U10950 (N_10950,N_2217,N_4119);
and U10951 (N_10951,N_9931,N_1210);
and U10952 (N_10952,N_9926,N_4683);
or U10953 (N_10953,N_4704,N_8981);
nand U10954 (N_10954,N_5659,N_936);
nand U10955 (N_10955,N_9330,N_6624);
and U10956 (N_10956,N_7947,N_6835);
nand U10957 (N_10957,N_3346,N_8395);
nand U10958 (N_10958,N_4306,N_5535);
or U10959 (N_10959,N_15,N_6470);
or U10960 (N_10960,N_8925,N_8408);
nor U10961 (N_10961,N_1160,N_6851);
or U10962 (N_10962,N_555,N_3568);
or U10963 (N_10963,N_4135,N_6526);
and U10964 (N_10964,N_498,N_3448);
or U10965 (N_10965,N_1062,N_9508);
nor U10966 (N_10966,N_5826,N_8304);
and U10967 (N_10967,N_7589,N_7881);
nor U10968 (N_10968,N_3632,N_8735);
nor U10969 (N_10969,N_7869,N_7125);
xor U10970 (N_10970,N_1715,N_2842);
or U10971 (N_10971,N_8349,N_9243);
or U10972 (N_10972,N_3508,N_8128);
nand U10973 (N_10973,N_5363,N_3102);
and U10974 (N_10974,N_9546,N_5359);
nand U10975 (N_10975,N_5154,N_3651);
xnor U10976 (N_10976,N_2710,N_8143);
xnor U10977 (N_10977,N_3221,N_385);
or U10978 (N_10978,N_1927,N_6817);
and U10979 (N_10979,N_5024,N_4236);
and U10980 (N_10980,N_7648,N_891);
nand U10981 (N_10981,N_120,N_70);
nor U10982 (N_10982,N_7333,N_7015);
and U10983 (N_10983,N_3017,N_1337);
or U10984 (N_10984,N_5068,N_597);
and U10985 (N_10985,N_9817,N_4599);
or U10986 (N_10986,N_4517,N_6226);
nand U10987 (N_10987,N_4967,N_4641);
nor U10988 (N_10988,N_4589,N_6428);
nand U10989 (N_10989,N_3159,N_6243);
and U10990 (N_10990,N_4466,N_9023);
nor U10991 (N_10991,N_3551,N_8370);
or U10992 (N_10992,N_6929,N_9338);
nor U10993 (N_10993,N_1488,N_4179);
and U10994 (N_10994,N_1777,N_4489);
nor U10995 (N_10995,N_1059,N_6595);
or U10996 (N_10996,N_3737,N_2431);
xor U10997 (N_10997,N_792,N_9455);
nand U10998 (N_10998,N_5693,N_3294);
nor U10999 (N_10999,N_8809,N_7480);
nor U11000 (N_11000,N_1313,N_6213);
xnor U11001 (N_11001,N_8325,N_8943);
nor U11002 (N_11002,N_5303,N_782);
or U11003 (N_11003,N_4756,N_5038);
and U11004 (N_11004,N_5322,N_4146);
nor U11005 (N_11005,N_6421,N_304);
nor U11006 (N_11006,N_4358,N_1685);
and U11007 (N_11007,N_228,N_2155);
nand U11008 (N_11008,N_2330,N_691);
nor U11009 (N_11009,N_4555,N_5368);
and U11010 (N_11010,N_9570,N_2908);
nand U11011 (N_11011,N_2534,N_409);
nand U11012 (N_11012,N_2713,N_7600);
nor U11013 (N_11013,N_661,N_5209);
or U11014 (N_11014,N_1518,N_8375);
nand U11015 (N_11015,N_4005,N_144);
and U11016 (N_11016,N_8791,N_4832);
nand U11017 (N_11017,N_7631,N_3777);
nand U11018 (N_11018,N_1266,N_9907);
xor U11019 (N_11019,N_7839,N_2213);
nor U11020 (N_11020,N_3363,N_7542);
xnor U11021 (N_11021,N_1512,N_8907);
or U11022 (N_11022,N_4283,N_7089);
nand U11023 (N_11023,N_6181,N_5747);
nor U11024 (N_11024,N_9422,N_8973);
nor U11025 (N_11025,N_8511,N_6010);
xor U11026 (N_11026,N_478,N_3829);
or U11027 (N_11027,N_3906,N_7538);
nor U11028 (N_11028,N_4281,N_1594);
or U11029 (N_11029,N_4785,N_7218);
or U11030 (N_11030,N_9276,N_9884);
nand U11031 (N_11031,N_4711,N_6241);
and U11032 (N_11032,N_8842,N_4914);
or U11033 (N_11033,N_2970,N_9659);
or U11034 (N_11034,N_1204,N_9030);
nand U11035 (N_11035,N_2405,N_9281);
nor U11036 (N_11036,N_8458,N_4087);
or U11037 (N_11037,N_8222,N_3166);
nand U11038 (N_11038,N_5375,N_4174);
and U11039 (N_11039,N_1214,N_4483);
and U11040 (N_11040,N_7865,N_7779);
or U11041 (N_11041,N_6616,N_9181);
or U11042 (N_11042,N_9064,N_1667);
or U11043 (N_11043,N_4450,N_9378);
and U11044 (N_11044,N_1001,N_7499);
nand U11045 (N_11045,N_5137,N_9691);
and U11046 (N_11046,N_3740,N_7553);
or U11047 (N_11047,N_7692,N_7050);
and U11048 (N_11048,N_5382,N_9577);
or U11049 (N_11049,N_2836,N_522);
nand U11050 (N_11050,N_5706,N_5614);
nand U11051 (N_11051,N_9753,N_9406);
xnor U11052 (N_11052,N_9899,N_222);
nand U11053 (N_11053,N_4777,N_74);
nand U11054 (N_11054,N_3754,N_4006);
nand U11055 (N_11055,N_3038,N_8412);
nand U11056 (N_11056,N_7248,N_6791);
nand U11057 (N_11057,N_4652,N_5782);
nand U11058 (N_11058,N_8054,N_2495);
nor U11059 (N_11059,N_4378,N_2163);
nor U11060 (N_11060,N_9543,N_5763);
nand U11061 (N_11061,N_9911,N_4029);
nor U11062 (N_11062,N_2515,N_5822);
nor U11063 (N_11063,N_3057,N_5399);
or U11064 (N_11064,N_3835,N_5638);
nand U11065 (N_11065,N_1843,N_4600);
nand U11066 (N_11066,N_3370,N_1003);
nand U11067 (N_11067,N_2889,N_8594);
nor U11068 (N_11068,N_6221,N_280);
nand U11069 (N_11069,N_4010,N_2951);
nand U11070 (N_11070,N_1480,N_4052);
and U11071 (N_11071,N_5857,N_8608);
xnor U11072 (N_11072,N_8205,N_4604);
and U11073 (N_11073,N_7606,N_7906);
and U11074 (N_11074,N_5548,N_3916);
nand U11075 (N_11075,N_2354,N_9951);
xor U11076 (N_11076,N_6636,N_8680);
nor U11077 (N_11077,N_8418,N_8138);
nand U11078 (N_11078,N_2210,N_9803);
nor U11079 (N_11079,N_9994,N_7985);
or U11080 (N_11080,N_3947,N_505);
or U11081 (N_11081,N_889,N_2767);
nor U11082 (N_11082,N_7038,N_6767);
xor U11083 (N_11083,N_6753,N_8649);
xor U11084 (N_11084,N_4668,N_8544);
xor U11085 (N_11085,N_7278,N_7164);
nand U11086 (N_11086,N_6566,N_4123);
xnor U11087 (N_11087,N_8742,N_8901);
and U11088 (N_11088,N_2671,N_6495);
nor U11089 (N_11089,N_739,N_3969);
or U11090 (N_11090,N_9993,N_7243);
nand U11091 (N_11091,N_3684,N_6414);
or U11092 (N_11092,N_8967,N_9153);
and U11093 (N_11093,N_5151,N_7403);
and U11094 (N_11094,N_7233,N_9353);
nand U11095 (N_11095,N_5553,N_3033);
nor U11096 (N_11096,N_4412,N_2629);
xnor U11097 (N_11097,N_2471,N_1952);
nor U11098 (N_11098,N_2722,N_9212);
nor U11099 (N_11099,N_2910,N_6429);
nor U11100 (N_11100,N_5773,N_5882);
xor U11101 (N_11101,N_7239,N_1900);
xnor U11102 (N_11102,N_4990,N_5046);
or U11103 (N_11103,N_9825,N_8402);
nand U11104 (N_11104,N_4019,N_3098);
nand U11105 (N_11105,N_5159,N_3355);
and U11106 (N_11106,N_9548,N_7540);
xor U11107 (N_11107,N_314,N_7182);
nor U11108 (N_11108,N_5644,N_2179);
or U11109 (N_11109,N_8667,N_9611);
nor U11110 (N_11110,N_8416,N_5713);
and U11111 (N_11111,N_7167,N_8056);
or U11112 (N_11112,N_1956,N_2117);
nor U11113 (N_11113,N_4444,N_3139);
nand U11114 (N_11114,N_1100,N_4348);
xnor U11115 (N_11115,N_681,N_1182);
nor U11116 (N_11116,N_568,N_3500);
nor U11117 (N_11117,N_353,N_8916);
nor U11118 (N_11118,N_4884,N_9185);
or U11119 (N_11119,N_853,N_4948);
nand U11120 (N_11120,N_9006,N_389);
nor U11121 (N_11121,N_3488,N_3122);
xnor U11122 (N_11122,N_4594,N_4544);
and U11123 (N_11123,N_114,N_8306);
xnor U11124 (N_11124,N_3977,N_1133);
xnor U11125 (N_11125,N_1870,N_6304);
nand U11126 (N_11126,N_6695,N_8082);
nand U11127 (N_11127,N_6762,N_6689);
nor U11128 (N_11128,N_6988,N_8512);
or U11129 (N_11129,N_4407,N_7524);
nand U11130 (N_11130,N_3124,N_514);
nand U11131 (N_11131,N_7837,N_5630);
xor U11132 (N_11132,N_8142,N_6255);
and U11133 (N_11133,N_5165,N_7801);
or U11134 (N_11134,N_2387,N_2237);
xor U11135 (N_11135,N_83,N_9214);
or U11136 (N_11136,N_7771,N_287);
and U11137 (N_11137,N_6207,N_1209);
or U11138 (N_11138,N_7706,N_9842);
and U11139 (N_11139,N_8695,N_888);
or U11140 (N_11140,N_398,N_8);
xnor U11141 (N_11141,N_538,N_5957);
nor U11142 (N_11142,N_4318,N_7367);
nor U11143 (N_11143,N_4736,N_9170);
and U11144 (N_11144,N_5998,N_3381);
and U11145 (N_11145,N_3310,N_2396);
or U11146 (N_11146,N_1166,N_9372);
or U11147 (N_11147,N_9882,N_7677);
nand U11148 (N_11148,N_4921,N_6045);
and U11149 (N_11149,N_8787,N_6396);
xor U11150 (N_11150,N_3751,N_6459);
nand U11151 (N_11151,N_2523,N_3053);
xor U11152 (N_11152,N_1430,N_7463);
nand U11153 (N_11153,N_8407,N_4899);
nor U11154 (N_11154,N_8360,N_8621);
or U11155 (N_11155,N_9809,N_8281);
nor U11156 (N_11156,N_2664,N_5611);
and U11157 (N_11157,N_1838,N_5000);
or U11158 (N_11158,N_1393,N_5669);
xor U11159 (N_11159,N_5704,N_7866);
xor U11160 (N_11160,N_6457,N_6294);
and U11161 (N_11161,N_2383,N_1058);
xor U11162 (N_11162,N_20,N_1720);
nor U11163 (N_11163,N_6124,N_4719);
and U11164 (N_11164,N_5905,N_7657);
nand U11165 (N_11165,N_3530,N_9084);
or U11166 (N_11166,N_4917,N_3255);
nand U11167 (N_11167,N_4031,N_5868);
nor U11168 (N_11168,N_9647,N_5692);
nor U11169 (N_11169,N_2825,N_518);
nand U11170 (N_11170,N_125,N_6725);
and U11171 (N_11171,N_1661,N_9304);
nor U11172 (N_11172,N_5800,N_5369);
nand U11173 (N_11173,N_9315,N_2389);
and U11174 (N_11174,N_986,N_985);
or U11175 (N_11175,N_1334,N_3608);
xnor U11176 (N_11176,N_9327,N_2209);
nor U11177 (N_11177,N_2131,N_9234);
xnor U11178 (N_11178,N_8240,N_8918);
nor U11179 (N_11179,N_6225,N_1966);
nand U11180 (N_11180,N_1891,N_7059);
nand U11181 (N_11181,N_365,N_1823);
nor U11182 (N_11182,N_7973,N_8966);
and U11183 (N_11183,N_4202,N_9249);
or U11184 (N_11184,N_2088,N_8915);
or U11185 (N_11185,N_4245,N_357);
and U11186 (N_11186,N_4892,N_6434);
nand U11187 (N_11187,N_4801,N_2038);
or U11188 (N_11188,N_8078,N_3293);
or U11189 (N_11189,N_1179,N_3271);
nor U11190 (N_11190,N_8208,N_7743);
or U11191 (N_11191,N_987,N_9086);
xor U11192 (N_11192,N_7037,N_1267);
xnor U11193 (N_11193,N_7088,N_5917);
xnor U11194 (N_11194,N_4118,N_9790);
or U11195 (N_11195,N_8321,N_1206);
or U11196 (N_11196,N_6994,N_8886);
nor U11197 (N_11197,N_1901,N_8160);
and U11198 (N_11198,N_252,N_2773);
nand U11199 (N_11199,N_53,N_5691);
xnor U11200 (N_11200,N_3112,N_9709);
nor U11201 (N_11201,N_1338,N_7060);
xor U11202 (N_11202,N_5248,N_3008);
nand U11203 (N_11203,N_3903,N_3908);
nor U11204 (N_11204,N_7294,N_7411);
nor U11205 (N_11205,N_7242,N_9485);
xnor U11206 (N_11206,N_2550,N_6514);
nand U11207 (N_11207,N_4153,N_1511);
and U11208 (N_11208,N_7900,N_5093);
or U11209 (N_11209,N_4328,N_2293);
and U11210 (N_11210,N_7791,N_4055);
and U11211 (N_11211,N_6059,N_9594);
nand U11212 (N_11212,N_6750,N_4381);
nand U11213 (N_11213,N_6080,N_3323);
or U11214 (N_11214,N_9121,N_932);
nand U11215 (N_11215,N_8622,N_3248);
xnor U11216 (N_11216,N_6650,N_3047);
and U11217 (N_11217,N_5807,N_6679);
and U11218 (N_11218,N_2958,N_5145);
xnor U11219 (N_11219,N_7492,N_3104);
nand U11220 (N_11220,N_9250,N_4325);
nor U11221 (N_11221,N_7041,N_897);
nor U11222 (N_11222,N_2730,N_6166);
nand U11223 (N_11223,N_8326,N_894);
nor U11224 (N_11224,N_7759,N_2530);
or U11225 (N_11225,N_4096,N_5459);
or U11226 (N_11226,N_6211,N_5189);
nor U11227 (N_11227,N_9903,N_2946);
and U11228 (N_11228,N_6219,N_8706);
or U11229 (N_11229,N_9751,N_23);
and U11230 (N_11230,N_1509,N_3970);
or U11231 (N_11231,N_7241,N_9984);
and U11232 (N_11232,N_945,N_7967);
xnor U11233 (N_11233,N_1094,N_9658);
or U11234 (N_11234,N_7997,N_8568);
nor U11235 (N_11235,N_8369,N_3397);
nand U11236 (N_11236,N_2989,N_1928);
xor U11237 (N_11237,N_7756,N_7189);
or U11238 (N_11238,N_4551,N_2561);
or U11239 (N_11239,N_2853,N_3019);
xor U11240 (N_11240,N_1431,N_1562);
or U11241 (N_11241,N_1365,N_9579);
xnor U11242 (N_11242,N_8439,N_109);
nor U11243 (N_11243,N_2982,N_1504);
nor U11244 (N_11244,N_1191,N_6055);
and U11245 (N_11245,N_6122,N_9200);
nand U11246 (N_11246,N_3003,N_5673);
and U11247 (N_11247,N_8557,N_2883);
or U11248 (N_11248,N_1957,N_7763);
nand U11249 (N_11249,N_1072,N_934);
or U11250 (N_11250,N_7054,N_700);
xnor U11251 (N_11251,N_3918,N_9666);
nor U11252 (N_11252,N_5450,N_9);
nand U11253 (N_11253,N_3216,N_8992);
xor U11254 (N_11254,N_3503,N_2406);
nor U11255 (N_11255,N_5357,N_9155);
and U11256 (N_11256,N_7192,N_892);
nand U11257 (N_11257,N_1701,N_6390);
nor U11258 (N_11258,N_6134,N_7663);
nand U11259 (N_11259,N_7384,N_8319);
nand U11260 (N_11260,N_5218,N_4038);
and U11261 (N_11261,N_5859,N_7287);
nand U11262 (N_11262,N_9960,N_9612);
nand U11263 (N_11263,N_9694,N_4421);
xnor U11264 (N_11264,N_2410,N_6197);
xor U11265 (N_11265,N_5581,N_3331);
or U11266 (N_11266,N_6218,N_1362);
xnor U11267 (N_11267,N_1060,N_2932);
nor U11268 (N_11268,N_92,N_4816);
nor U11269 (N_11269,N_1384,N_3001);
nor U11270 (N_11270,N_9774,N_5839);
and U11271 (N_11271,N_8004,N_8891);
or U11272 (N_11272,N_9860,N_2699);
or U11273 (N_11273,N_6698,N_7177);
and U11274 (N_11274,N_1423,N_9567);
nand U11275 (N_11275,N_3644,N_4061);
and U11276 (N_11276,N_1192,N_3232);
or U11277 (N_11277,N_787,N_7179);
xor U11278 (N_11278,N_6834,N_8330);
nor U11279 (N_11279,N_472,N_8276);
and U11280 (N_11280,N_6555,N_9117);
or U11281 (N_11281,N_8919,N_884);
nor U11282 (N_11282,N_3685,N_367);
nor U11283 (N_11283,N_5841,N_1725);
nand U11284 (N_11284,N_9624,N_4961);
nor U11285 (N_11285,N_7665,N_5646);
or U11286 (N_11286,N_2352,N_5968);
and U11287 (N_11287,N_3402,N_4158);
nor U11288 (N_11288,N_4913,N_6231);
nand U11289 (N_11289,N_2638,N_6446);
nor U11290 (N_11290,N_1909,N_6815);
xor U11291 (N_11291,N_7807,N_1295);
or U11292 (N_11292,N_3341,N_3900);
or U11293 (N_11293,N_9311,N_6186);
or U11294 (N_11294,N_3308,N_4387);
nor U11295 (N_11295,N_8152,N_3414);
xor U11296 (N_11296,N_9688,N_5034);
nand U11297 (N_11297,N_520,N_3909);
nor U11298 (N_11298,N_4169,N_3580);
nand U11299 (N_11299,N_7621,N_9438);
nor U11300 (N_11300,N_7808,N_311);
nand U11301 (N_11301,N_3889,N_9385);
nor U11302 (N_11302,N_3679,N_1478);
xor U11303 (N_11303,N_5510,N_1775);
nand U11304 (N_11304,N_1842,N_9258);
and U11305 (N_11305,N_429,N_647);
or U11306 (N_11306,N_6020,N_7832);
or U11307 (N_11307,N_4218,N_4349);
nor U11308 (N_11308,N_403,N_1696);
xnor U11309 (N_11309,N_5346,N_2711);
nand U11310 (N_11310,N_7998,N_6217);
xnor U11311 (N_11311,N_8790,N_5722);
and U11312 (N_11312,N_3197,N_5932);
and U11313 (N_11313,N_2105,N_1358);
nand U11314 (N_11314,N_9698,N_635);
or U11315 (N_11315,N_3815,N_425);
xnor U11316 (N_11316,N_1466,N_7185);
and U11317 (N_11317,N_9711,N_7826);
and U11318 (N_11318,N_4669,N_2064);
and U11319 (N_11319,N_8204,N_4592);
nand U11320 (N_11320,N_6091,N_5764);
and U11321 (N_11321,N_9232,N_974);
nor U11322 (N_11322,N_8207,N_4706);
or U11323 (N_11323,N_2955,N_9524);
xnor U11324 (N_11324,N_2937,N_9301);
nor U11325 (N_11325,N_524,N_4688);
nor U11326 (N_11326,N_6095,N_8498);
nand U11327 (N_11327,N_4605,N_693);
or U11328 (N_11328,N_117,N_7733);
nor U11329 (N_11329,N_7285,N_6939);
nor U11330 (N_11330,N_4224,N_5946);
or U11331 (N_11331,N_1141,N_4404);
or U11332 (N_11332,N_995,N_7352);
nand U11333 (N_11333,N_1809,N_5031);
nand U11334 (N_11334,N_9293,N_3082);
nand U11335 (N_11335,N_3992,N_9166);
or U11336 (N_11336,N_8136,N_6539);
nor U11337 (N_11337,N_2068,N_1075);
nor U11338 (N_11338,N_8362,N_7946);
or U11339 (N_11339,N_9650,N_2748);
or U11340 (N_11340,N_6935,N_7210);
nor U11341 (N_11341,N_265,N_8179);
and U11342 (N_11342,N_4746,N_3340);
xor U11343 (N_11343,N_1453,N_9360);
and U11344 (N_11344,N_9728,N_7163);
or U11345 (N_11345,N_5020,N_4797);
and U11346 (N_11346,N_2417,N_3393);
xnor U11347 (N_11347,N_1024,N_7069);
and U11348 (N_11348,N_3259,N_5605);
xor U11349 (N_11349,N_327,N_8151);
and U11350 (N_11350,N_6617,N_2524);
xor U11351 (N_11351,N_9362,N_2288);
xnor U11352 (N_11352,N_8582,N_2430);
nand U11353 (N_11353,N_3526,N_7320);
and U11354 (N_11354,N_9405,N_6461);
nand U11355 (N_11355,N_657,N_201);
or U11356 (N_11356,N_3400,N_8315);
xor U11357 (N_11357,N_9602,N_857);
or U11358 (N_11358,N_3781,N_1813);
and U11359 (N_11359,N_9834,N_6261);
nor U11360 (N_11360,N_6162,N_388);
and U11361 (N_11361,N_4679,N_1839);
and U11362 (N_11362,N_9075,N_6582);
nor U11363 (N_11363,N_1501,N_2704);
nand U11364 (N_11364,N_2774,N_5494);
or U11365 (N_11365,N_3739,N_1317);
xor U11366 (N_11366,N_1458,N_1655);
or U11367 (N_11367,N_6444,N_6735);
nor U11368 (N_11368,N_8937,N_7330);
and U11369 (N_11369,N_4955,N_1580);
and U11370 (N_11370,N_4431,N_3654);
or U11371 (N_11371,N_424,N_5565);
xnor U11372 (N_11372,N_306,N_4659);
nor U11373 (N_11373,N_8247,N_1932);
and U11374 (N_11374,N_5397,N_3726);
nor U11375 (N_11375,N_3099,N_1705);
and U11376 (N_11376,N_9018,N_2264);
nand U11377 (N_11377,N_3230,N_5282);
and U11378 (N_11378,N_509,N_7698);
and U11379 (N_11379,N_6608,N_2307);
nor U11380 (N_11380,N_6536,N_4936);
nand U11381 (N_11381,N_8490,N_4045);
or U11382 (N_11382,N_6158,N_1360);
xor U11383 (N_11383,N_941,N_1049);
xor U11384 (N_11384,N_3883,N_9130);
and U11385 (N_11385,N_9356,N_9730);
and U11386 (N_11386,N_2177,N_9082);
xnor U11387 (N_11387,N_143,N_8124);
or U11388 (N_11388,N_4448,N_1090);
nand U11389 (N_11389,N_8522,N_2912);
or U11390 (N_11390,N_8940,N_2743);
nor U11391 (N_11391,N_2536,N_2700);
and U11392 (N_11392,N_376,N_9171);
nand U11393 (N_11393,N_3571,N_8752);
and U11394 (N_11394,N_9610,N_3796);
and U11395 (N_11395,N_802,N_5200);
nand U11396 (N_11396,N_2821,N_2434);
xnor U11397 (N_11397,N_2707,N_2920);
or U11398 (N_11398,N_3097,N_6949);
nand U11399 (N_11399,N_3382,N_2715);
or U11400 (N_11400,N_2313,N_5663);
or U11401 (N_11401,N_8361,N_2858);
nor U11402 (N_11402,N_4116,N_1021);
xor U11403 (N_11403,N_3021,N_3720);
and U11404 (N_11404,N_8687,N_4221);
nor U11405 (N_11405,N_4794,N_4946);
xnor U11406 (N_11406,N_8644,N_5641);
nand U11407 (N_11407,N_2014,N_2034);
or U11408 (N_11408,N_8598,N_5934);
and U11409 (N_11409,N_5089,N_6556);
and U11410 (N_11410,N_9626,N_6490);
or U11411 (N_11411,N_8852,N_849);
or U11412 (N_11412,N_8740,N_4461);
nor U11413 (N_11413,N_1446,N_8327);
xnor U11414 (N_11414,N_7103,N_5409);
or U11415 (N_11415,N_6688,N_3254);
xor U11416 (N_11416,N_258,N_3940);
nor U11417 (N_11417,N_2930,N_3497);
nand U11418 (N_11418,N_5442,N_5840);
nor U11419 (N_11419,N_4278,N_5156);
and U11420 (N_11420,N_7331,N_183);
and U11421 (N_11421,N_9164,N_4214);
xnor U11422 (N_11422,N_185,N_2506);
xor U11423 (N_11423,N_733,N_5304);
or U11424 (N_11424,N_9561,N_554);
nand U11425 (N_11425,N_6803,N_7519);
nand U11426 (N_11426,N_6598,N_5714);
nor U11427 (N_11427,N_8001,N_5928);
or U11428 (N_11428,N_7531,N_7905);
xor U11429 (N_11429,N_9179,N_5527);
or U11430 (N_11430,N_1703,N_8781);
xnor U11431 (N_11431,N_5231,N_6326);
or U11432 (N_11432,N_9332,N_6619);
nor U11433 (N_11433,N_9740,N_1045);
and U11434 (N_11434,N_1885,N_537);
nand U11435 (N_11435,N_948,N_666);
nor U11436 (N_11436,N_4677,N_8285);
and U11437 (N_11437,N_4429,N_777);
and U11438 (N_11438,N_8670,N_920);
and U11439 (N_11439,N_8761,N_9124);
nor U11440 (N_11440,N_7139,N_440);
nor U11441 (N_11441,N_2024,N_9320);
or U11442 (N_11442,N_4657,N_427);
xor U11443 (N_11443,N_533,N_111);
xor U11444 (N_11444,N_6399,N_4847);
or U11445 (N_11445,N_7748,N_6127);
xor U11446 (N_11446,N_4464,N_6228);
and U11447 (N_11447,N_9302,N_858);
nand U11448 (N_11448,N_9665,N_8338);
and U11449 (N_11449,N_5295,N_4492);
nand U11450 (N_11450,N_6193,N_6064);
nor U11451 (N_11451,N_2365,N_3023);
nand U11452 (N_11452,N_1421,N_8026);
xor U11453 (N_11453,N_3546,N_4613);
and U11454 (N_11454,N_5439,N_9450);
nor U11455 (N_11455,N_8091,N_5249);
nor U11456 (N_11456,N_272,N_7366);
and U11457 (N_11457,N_5244,N_1004);
nor U11458 (N_11458,N_5592,N_5122);
nand U11459 (N_11459,N_6645,N_9734);
and U11460 (N_11460,N_4718,N_1391);
or U11461 (N_11461,N_9227,N_5562);
xnor U11462 (N_11462,N_488,N_569);
nand U11463 (N_11463,N_6731,N_4109);
nor U11464 (N_11464,N_6352,N_4191);
xor U11465 (N_11465,N_3486,N_469);
and U11466 (N_11466,N_596,N_774);
nor U11467 (N_11467,N_5077,N_3214);
nand U11468 (N_11468,N_7142,N_8110);
xnor U11469 (N_11469,N_349,N_87);
and U11470 (N_11470,N_7854,N_8944);
nand U11471 (N_11471,N_8299,N_5612);
or U11472 (N_11472,N_2033,N_9377);
nor U11473 (N_11473,N_1659,N_7341);
and U11474 (N_11474,N_2428,N_513);
or U11475 (N_11475,N_8625,N_6649);
or U11476 (N_11476,N_5919,N_7379);
xnor U11477 (N_11477,N_7725,N_3957);
or U11478 (N_11478,N_4094,N_9716);
and U11479 (N_11479,N_6614,N_5117);
or U11480 (N_11480,N_9723,N_4648);
and U11481 (N_11481,N_1958,N_7925);
or U11482 (N_11482,N_4478,N_7577);
nor U11483 (N_11483,N_8930,N_9796);
or U11484 (N_11484,N_2905,N_2095);
nor U11485 (N_11485,N_2244,N_7345);
xor U11486 (N_11486,N_1646,N_8216);
xnor U11487 (N_11487,N_566,N_1918);
and U11488 (N_11488,N_497,N_9722);
nor U11489 (N_11489,N_4144,N_1519);
nand U11490 (N_11490,N_5221,N_6500);
xor U11491 (N_11491,N_8789,N_2571);
xor U11492 (N_11492,N_2619,N_7721);
nand U11493 (N_11493,N_2370,N_4754);
and U11494 (N_11494,N_8951,N_7778);
and U11495 (N_11495,N_8693,N_9970);
and U11496 (N_11496,N_5774,N_2902);
nand U11497 (N_11497,N_5086,N_2374);
nor U11498 (N_11498,N_1830,N_7277);
nor U11499 (N_11499,N_560,N_6119);
nand U11500 (N_11500,N_5981,N_4951);
nand U11501 (N_11501,N_1444,N_6168);
xor U11502 (N_11502,N_2740,N_7629);
or U11503 (N_11503,N_7794,N_2200);
nor U11504 (N_11504,N_1052,N_2673);
and U11505 (N_11505,N_2745,N_1852);
or U11506 (N_11506,N_3484,N_1180);
nor U11507 (N_11507,N_4485,N_6602);
or U11508 (N_11508,N_470,N_6191);
xnor U11509 (N_11509,N_947,N_3769);
nand U11510 (N_11510,N_4220,N_2075);
xnor U11511 (N_11511,N_1380,N_4837);
nand U11512 (N_11512,N_64,N_4192);
and U11513 (N_11513,N_9479,N_1651);
and U11514 (N_11514,N_333,N_2031);
nor U11515 (N_11515,N_6466,N_5593);
and U11516 (N_11516,N_4971,N_9912);
xnor U11517 (N_11517,N_9141,N_7739);
or U11518 (N_11518,N_5787,N_1818);
or U11519 (N_11519,N_2245,N_770);
nor U11520 (N_11520,N_236,N_8287);
or U11521 (N_11521,N_3450,N_2596);
nor U11522 (N_11522,N_8822,N_4695);
nor U11523 (N_11523,N_2463,N_5108);
or U11524 (N_11524,N_6474,N_4437);
or U11525 (N_11525,N_8873,N_4250);
and U11526 (N_11526,N_9414,N_5129);
nand U11527 (N_11527,N_2284,N_1998);
nor U11528 (N_11528,N_2416,N_3773);
nand U11529 (N_11529,N_7858,N_2126);
or U11530 (N_11530,N_2575,N_8318);
or U11531 (N_11531,N_170,N_822);
xor U11532 (N_11532,N_9103,N_890);
nand U11533 (N_11533,N_7325,N_3921);
or U11534 (N_11534,N_8213,N_3237);
nor U11535 (N_11535,N_9741,N_592);
or U11536 (N_11536,N_5676,N_9717);
nand U11537 (N_11537,N_1186,N_3721);
or U11538 (N_11538,N_1309,N_8073);
and U11539 (N_11539,N_6351,N_5785);
nand U11540 (N_11540,N_7670,N_6707);
and U11541 (N_11541,N_6507,N_9430);
nor U11542 (N_11542,N_4252,N_6245);
and U11543 (N_11543,N_9733,N_1397);
or U11544 (N_11544,N_508,N_4487);
and U11545 (N_11545,N_6561,N_7525);
xor U11546 (N_11546,N_9792,N_4836);
nor U11547 (N_11547,N_1684,N_7827);
or U11548 (N_11548,N_8711,N_4013);
nor U11549 (N_11549,N_5891,N_7849);
xor U11550 (N_11550,N_358,N_390);
and U11551 (N_11551,N_3138,N_7495);
or U11552 (N_11552,N_1588,N_5709);
nor U11553 (N_11553,N_4745,N_9446);
nor U11554 (N_11554,N_5401,N_4230);
nand U11555 (N_11555,N_1419,N_4465);
nand U11556 (N_11556,N_8194,N_1174);
nor U11557 (N_11557,N_3109,N_7641);
or U11558 (N_11558,N_3320,N_9542);
xnor U11559 (N_11559,N_5082,N_8834);
nand U11560 (N_11560,N_268,N_1198);
or U11561 (N_11561,N_6079,N_7244);
xnor U11562 (N_11562,N_1548,N_7720);
nor U11563 (N_11563,N_9396,N_4014);
nand U11564 (N_11564,N_9576,N_2042);
and U11565 (N_11565,N_8379,N_6634);
nor U11566 (N_11566,N_337,N_2517);
xnor U11567 (N_11567,N_9033,N_8359);
nor U11568 (N_11568,N_3063,N_8857);
nor U11569 (N_11569,N_1145,N_9308);
nor U11570 (N_11570,N_730,N_3875);
xnor U11571 (N_11571,N_1999,N_3013);
or U11572 (N_11572,N_3266,N_3280);
nand U11573 (N_11573,N_3192,N_1139);
and U11574 (N_11574,N_5158,N_4237);
or U11575 (N_11575,N_8854,N_1415);
xnor U11576 (N_11576,N_9129,N_39);
xnor U11577 (N_11577,N_3952,N_8785);
and U11578 (N_11578,N_9000,N_2250);
or U11579 (N_11579,N_3742,N_2814);
or U11580 (N_11580,N_6229,N_6109);
or U11581 (N_11581,N_9024,N_5);
and U11582 (N_11582,N_638,N_5803);
nand U11583 (N_11583,N_1330,N_4388);
nor U11584 (N_11584,N_2867,N_5835);
xor U11585 (N_11585,N_5058,N_3620);
xnor U11586 (N_11586,N_5497,N_5885);
nor U11587 (N_11587,N_9115,N_173);
nand U11588 (N_11588,N_226,N_3534);
nand U11589 (N_11589,N_7788,N_4638);
or U11590 (N_11590,N_4426,N_8673);
or U11591 (N_11591,N_8199,N_5070);
nor U11592 (N_11592,N_7668,N_1568);
and U11593 (N_11593,N_5320,N_1592);
and U11594 (N_11594,N_9883,N_4774);
xor U11595 (N_11595,N_8230,N_3733);
nor U11596 (N_11596,N_1017,N_2559);
nand U11597 (N_11597,N_7855,N_4107);
and U11598 (N_11598,N_6794,N_2617);
and U11599 (N_11599,N_8969,N_7376);
nor U11600 (N_11600,N_6787,N_2627);
nand U11601 (N_11601,N_5074,N_6271);
xor U11602 (N_11602,N_347,N_9132);
xnor U11603 (N_11603,N_4915,N_5274);
nand U11604 (N_11604,N_5431,N_8731);
xnor U11605 (N_11605,N_6092,N_2555);
nand U11606 (N_11606,N_4979,N_6149);
or U11607 (N_11607,N_7780,N_7373);
xnor U11608 (N_11608,N_3175,N_9757);
xnor U11609 (N_11609,N_2826,N_243);
nor U11610 (N_11610,N_6643,N_9642);
and U11611 (N_11611,N_2636,N_328);
nand U11612 (N_11612,N_6848,N_6272);
xnor U11613 (N_11613,N_3993,N_2233);
xnor U11614 (N_11614,N_3016,N_8562);
xnor U11615 (N_11615,N_9643,N_3998);
nand U11616 (N_11616,N_1449,N_387);
nand U11617 (N_11617,N_10,N_8510);
nor U11618 (N_11618,N_3265,N_4650);
nand U11619 (N_11619,N_4709,N_1872);
and U11620 (N_11620,N_9454,N_9216);
xor U11621 (N_11621,N_3996,N_1250);
nor U11622 (N_11622,N_8810,N_8021);
or U11623 (N_11623,N_1915,N_2897);
nor U11624 (N_11624,N_5336,N_7847);
nor U11625 (N_11625,N_7993,N_1603);
or U11626 (N_11626,N_7572,N_1106);
nor U11627 (N_11627,N_3405,N_5855);
nor U11628 (N_11628,N_2438,N_4997);
nand U11629 (N_11629,N_9262,N_2141);
nand U11630 (N_11630,N_4120,N_6063);
nand U11631 (N_11631,N_6058,N_2529);
xnor U11632 (N_11632,N_7979,N_7581);
xnor U11633 (N_11633,N_8538,N_4502);
xor U11634 (N_11634,N_9933,N_3984);
nand U11635 (N_11635,N_8817,N_3604);
or U11636 (N_11636,N_213,N_396);
nand U11637 (N_11637,N_2286,N_848);
or U11638 (N_11638,N_4645,N_1355);
xnor U11639 (N_11639,N_3196,N_2580);
xor U11640 (N_11640,N_8962,N_3779);
nor U11641 (N_11641,N_5289,N_7959);
or U11642 (N_11642,N_9603,N_8672);
xor U11643 (N_11643,N_8177,N_7450);
and U11644 (N_11644,N_1263,N_1739);
nand U11645 (N_11645,N_7644,N_8440);
nand U11646 (N_11646,N_8867,N_6873);
nor U11647 (N_11647,N_2123,N_9590);
nor U11648 (N_11648,N_5874,N_2547);
and U11649 (N_11649,N_110,N_5634);
or U11650 (N_11650,N_6008,N_8603);
nand U11651 (N_11651,N_7234,N_4542);
or U11652 (N_11652,N_8434,N_7190);
nand U11653 (N_11653,N_2037,N_1647);
xnor U11654 (N_11654,N_1886,N_3544);
nor U11655 (N_11655,N_6425,N_139);
nand U11656 (N_11656,N_8819,N_6838);
or U11657 (N_11657,N_2838,N_1699);
and U11658 (N_11658,N_7882,N_2949);
or U11659 (N_11659,N_2159,N_3963);
xor U11660 (N_11660,N_2801,N_2451);
xor U11661 (N_11661,N_4251,N_1553);
nand U11662 (N_11662,N_7042,N_7416);
nand U11663 (N_11663,N_6847,N_2735);
and U11664 (N_11664,N_1810,N_4088);
or U11665 (N_11665,N_26,N_7501);
or U11666 (N_11666,N_3845,N_5079);
and U11667 (N_11667,N_7666,N_3839);
xor U11668 (N_11668,N_4234,N_711);
xor U11669 (N_11669,N_1507,N_6323);
nand U11670 (N_11670,N_4543,N_598);
nor U11671 (N_11671,N_2865,N_5805);
and U11672 (N_11672,N_2810,N_9641);
xnor U11673 (N_11673,N_6590,N_4578);
nand U11674 (N_11674,N_3907,N_8956);
nor U11675 (N_11675,N_6596,N_3463);
xnor U11676 (N_11676,N_7044,N_7148);
or U11677 (N_11677,N_9971,N_2822);
and U11678 (N_11678,N_2388,N_7930);
nand U11679 (N_11679,N_8005,N_4952);
nor U11680 (N_11680,N_2901,N_9864);
and U11681 (N_11681,N_4945,N_5466);
or U11682 (N_11682,N_3167,N_6409);
nand U11683 (N_11683,N_336,N_7280);
nand U11684 (N_11684,N_9467,N_3514);
nand U11685 (N_11685,N_558,N_1390);
nor U11686 (N_11686,N_5746,N_5453);
nand U11687 (N_11687,N_8618,N_1220);
xor U11688 (N_11688,N_5757,N_623);
and U11689 (N_11689,N_2226,N_1088);
or U11690 (N_11690,N_4397,N_4334);
or U11691 (N_11691,N_581,N_1037);
or U11692 (N_11692,N_1328,N_6797);
nor U11693 (N_11693,N_6508,N_8396);
and U11694 (N_11694,N_8069,N_106);
and U11695 (N_11695,N_9954,N_4663);
or U11696 (N_11696,N_7343,N_59);
and U11697 (N_11697,N_116,N_1491);
xnor U11698 (N_11698,N_4203,N_2452);
xnor U11699 (N_11699,N_2863,N_6605);
xnor U11700 (N_11700,N_3668,N_3389);
and U11701 (N_11701,N_7922,N_1239);
nand U11702 (N_11702,N_7506,N_9902);
nand U11703 (N_11703,N_5410,N_1244);
and U11704 (N_11704,N_3791,N_673);
or U11705 (N_11705,N_7970,N_2943);
nand U11706 (N_11706,N_2733,N_5880);
or U11707 (N_11707,N_3938,N_9672);
xor U11708 (N_11708,N_1530,N_1770);
nor U11709 (N_11709,N_6,N_8385);
nand U11710 (N_11710,N_4249,N_9088);
and U11711 (N_11711,N_1113,N_7075);
or U11712 (N_11712,N_9384,N_5621);
nor U11713 (N_11713,N_1016,N_3552);
xnor U11714 (N_11714,N_3264,N_6116);
nor U11715 (N_11715,N_6374,N_5884);
nor U11716 (N_11716,N_5513,N_1751);
nand U11717 (N_11717,N_211,N_2904);
and U11718 (N_11718,N_7289,N_6581);
nand U11719 (N_11719,N_7503,N_7697);
nor U11720 (N_11720,N_3623,N_2277);
and U11721 (N_11721,N_3045,N_5610);
xor U11722 (N_11722,N_4748,N_9146);
nand U11723 (N_11723,N_2214,N_5140);
and U11724 (N_11724,N_5811,N_6532);
or U11725 (N_11725,N_4386,N_8933);
and U11726 (N_11726,N_7194,N_2795);
xnor U11727 (N_11727,N_1735,N_3131);
and U11728 (N_11728,N_1671,N_9975);
nand U11729 (N_11729,N_6420,N_6048);
xnor U11730 (N_11730,N_8581,N_2407);
nor U11731 (N_11731,N_9867,N_3822);
or U11732 (N_11732,N_1229,N_1738);
or U11733 (N_11733,N_2928,N_7625);
and U11734 (N_11734,N_1279,N_5878);
xnor U11735 (N_11735,N_7181,N_5476);
xnor U11736 (N_11736,N_5379,N_3672);
nor U11737 (N_11737,N_7490,N_4684);
and U11738 (N_11738,N_6963,N_134);
and U11739 (N_11739,N_3173,N_5853);
nor U11740 (N_11740,N_8097,N_2527);
nand U11741 (N_11741,N_7963,N_1792);
xnor U11742 (N_11742,N_9268,N_2686);
or U11743 (N_11743,N_3565,N_9784);
nand U11744 (N_11744,N_1781,N_6981);
or U11745 (N_11745,N_5207,N_5888);
nor U11746 (N_11746,N_6591,N_5432);
nand U11747 (N_11747,N_9409,N_6479);
nand U11748 (N_11748,N_9604,N_6380);
nand U11749 (N_11749,N_6896,N_8513);
and U11750 (N_11750,N_7076,N_8075);
or U11751 (N_11751,N_4165,N_1989);
nand U11752 (N_11752,N_1855,N_341);
and U11753 (N_11753,N_1398,N_2453);
or U11754 (N_11754,N_6290,N_1285);
nor U11755 (N_11755,N_3474,N_7040);
or U11756 (N_11756,N_1628,N_3285);
and U11757 (N_11757,N_9294,N_7563);
nor U11758 (N_11758,N_230,N_1617);
xnor U11759 (N_11759,N_6167,N_1222);
or U11760 (N_11760,N_4490,N_984);
or U11761 (N_11761,N_7348,N_5761);
nand U11762 (N_11762,N_5745,N_402);
xnor U11763 (N_11763,N_5435,N_3211);
nor U11764 (N_11764,N_89,N_2043);
or U11765 (N_11765,N_4530,N_2675);
and U11766 (N_11766,N_5626,N_3036);
and U11767 (N_11767,N_4587,N_9099);
or U11768 (N_11768,N_1805,N_8604);
nand U11769 (N_11769,N_3700,N_8993);
nand U11770 (N_11770,N_9909,N_437);
nor U11771 (N_11771,N_1140,N_195);
xnor U11772 (N_11772,N_8022,N_5139);
nand U11773 (N_11773,N_7152,N_1135);
or U11774 (N_11774,N_4456,N_9051);
xnor U11775 (N_11775,N_368,N_352);
nor U11776 (N_11776,N_4,N_1565);
nand U11777 (N_11777,N_4814,N_2608);
or U11778 (N_11778,N_7585,N_7364);
nand U11779 (N_11779,N_791,N_5603);
xor U11780 (N_11780,N_204,N_8447);
xnor U11781 (N_11781,N_2080,N_5699);
and U11782 (N_11782,N_5568,N_351);
xor U11783 (N_11783,N_5971,N_8554);
and U11784 (N_11784,N_924,N_926);
nand U11785 (N_11785,N_1618,N_1908);
xnor U11786 (N_11786,N_6110,N_1143);
xor U11787 (N_11787,N_1323,N_9523);
and U11788 (N_11788,N_2726,N_7822);
nand U11789 (N_11789,N_8724,N_1290);
or U11790 (N_11790,N_5661,N_1883);
xnor U11791 (N_11791,N_4194,N_9497);
nand U11792 (N_11792,N_1499,N_9781);
or U11793 (N_11793,N_9839,N_71);
nor U11794 (N_11794,N_6965,N_869);
xor U11795 (N_11795,N_5264,N_2029);
or U11796 (N_11796,N_6388,N_734);
nor U11797 (N_11797,N_1120,N_2377);
or U11798 (N_11798,N_7198,N_1815);
nand U11799 (N_11799,N_1949,N_3579);
nand U11800 (N_11800,N_8122,N_2421);
nor U11801 (N_11801,N_4924,N_9690);
and U11802 (N_11802,N_2886,N_6888);
or U11803 (N_11803,N_3547,N_2319);
or U11804 (N_11804,N_1804,N_563);
nor U11805 (N_11805,N_927,N_1503);
and U11806 (N_11806,N_8853,N_7487);
nand U11807 (N_11807,N_4042,N_9474);
nand U11808 (N_11808,N_4246,N_4424);
nand U11809 (N_11809,N_6520,N_7316);
and U11810 (N_11810,N_3804,N_4576);
and U11811 (N_11811,N_1134,N_6880);
xor U11812 (N_11812,N_4596,N_7061);
nor U11813 (N_11813,N_1574,N_3645);
or U11814 (N_11814,N_5232,N_8487);
and U11815 (N_11815,N_9267,N_8874);
xnor U11816 (N_11816,N_2584,N_9199);
or U11817 (N_11817,N_6314,N_9890);
xor U11818 (N_11818,N_9616,N_7742);
and U11819 (N_11819,N_709,N_214);
and U11820 (N_11820,N_9844,N_767);
or U11821 (N_11821,N_2820,N_4769);
xnor U11822 (N_11822,N_5759,N_908);
nand U11823 (N_11823,N_4290,N_91);
xor U11824 (N_11824,N_3703,N_3390);
or U11825 (N_11825,N_181,N_8493);
nand U11826 (N_11826,N_9761,N_7962);
and U11827 (N_11827,N_315,N_1163);
xor U11828 (N_11828,N_7811,N_536);
xnor U11829 (N_11829,N_5858,N_7247);
or U11830 (N_11830,N_6317,N_4362);
xnor U11831 (N_11831,N_7444,N_7945);
xor U11832 (N_11832,N_9394,N_1464);
nor U11833 (N_11833,N_4705,N_3702);
nor U11834 (N_11834,N_510,N_8999);
and U11835 (N_11835,N_8585,N_3652);
or U11836 (N_11836,N_2507,N_4025);
nor U11837 (N_11837,N_6511,N_1527);
nand U11838 (N_11838,N_2342,N_2124);
xnor U11839 (N_11839,N_6077,N_8671);
or U11840 (N_11840,N_4505,N_6663);
nor U11841 (N_11841,N_493,N_381);
or U11842 (N_11842,N_5974,N_3851);
nor U11843 (N_11843,N_244,N_4630);
nand U11844 (N_11844,N_8495,N_7661);
nand U11845 (N_11845,N_671,N_1552);
and U11846 (N_11846,N_2001,N_6293);
and U11847 (N_11847,N_7217,N_2429);
xor U11848 (N_11848,N_5441,N_9502);
and U11849 (N_11849,N_3640,N_4929);
nand U11850 (N_11850,N_2148,N_1394);
xor U11851 (N_11851,N_1296,N_5877);
or U11852 (N_11852,N_342,N_3706);
and U11853 (N_11853,N_588,N_7936);
nand U11854 (N_11854,N_2358,N_6386);
nor U11855 (N_11855,N_9700,N_18);
nand U11856 (N_11856,N_5482,N_4632);
nand U11857 (N_11857,N_1124,N_7494);
xor U11858 (N_11858,N_3291,N_1914);
nor U11859 (N_11859,N_3738,N_180);
or U11860 (N_11860,N_5222,N_7914);
and U11861 (N_11861,N_4882,N_4372);
nand U11862 (N_11862,N_2097,N_2324);
xnor U11863 (N_11863,N_8883,N_9814);
and U11864 (N_11864,N_6170,N_2854);
nor U11865 (N_11865,N_7645,N_4482);
xnor U11866 (N_11866,N_6029,N_3872);
nand U11867 (N_11867,N_7485,N_9273);
nand U11868 (N_11868,N_3049,N_1882);
or U11869 (N_11869,N_531,N_2090);
nor U11870 (N_11870,N_5019,N_8995);
nor U11871 (N_11871,N_3572,N_4969);
and U11872 (N_11872,N_6830,N_206);
nor U11873 (N_11873,N_2393,N_9161);
or U11874 (N_11874,N_2134,N_7655);
and U11875 (N_11875,N_2425,N_9958);
xor U11876 (N_11876,N_8231,N_1078);
nand U11877 (N_11877,N_9163,N_4538);
nor U11878 (N_11878,N_9189,N_9111);
nor U11879 (N_11879,N_5651,N_6856);
nor U11880 (N_11880,N_8163,N_5961);
and U11881 (N_11881,N_1729,N_2379);
nand U11882 (N_11882,N_2644,N_9150);
or U11883 (N_11883,N_8441,N_6699);
xor U11884 (N_11884,N_1132,N_9383);
or U11885 (N_11885,N_4972,N_6647);
xor U11886 (N_11886,N_6991,N_612);
xnor U11887 (N_11887,N_6626,N_146);
or U11888 (N_11888,N_7652,N_4898);
nand U11889 (N_11889,N_5682,N_1920);
nor U11890 (N_11890,N_4451,N_1675);
xnor U11891 (N_11891,N_5549,N_8924);
xnor U11892 (N_11892,N_163,N_7227);
xnor U11893 (N_11893,N_8150,N_2202);
nor U11894 (N_11894,N_1639,N_4197);
nor U11895 (N_11895,N_6668,N_4890);
and U11896 (N_11896,N_3990,N_9034);
nand U11897 (N_11897,N_7469,N_8067);
nor U11898 (N_11898,N_3217,N_2663);
nor U11899 (N_11899,N_3309,N_9583);
nand U11900 (N_11900,N_3563,N_6244);
or U11901 (N_11901,N_8378,N_4233);
nor U11902 (N_11902,N_5018,N_5818);
or U11903 (N_11903,N_7623,N_7556);
and U11904 (N_11904,N_3296,N_1231);
nor U11905 (N_11905,N_8090,N_9881);
nor U11906 (N_11906,N_3692,N_2039);
nand U11907 (N_11907,N_9547,N_5417);
xnor U11908 (N_11908,N_7651,N_2697);
xnor U11909 (N_11909,N_1772,N_5817);
nand U11910 (N_11910,N_4373,N_8646);
nor U11911 (N_11911,N_2839,N_9037);
or U11912 (N_11912,N_2493,N_73);
nor U11913 (N_11913,N_3671,N_2252);
or U11914 (N_11914,N_2903,N_5760);
nor U11915 (N_11915,N_9934,N_2345);
nor U11916 (N_11916,N_6685,N_4911);
xor U11917 (N_11917,N_9683,N_5206);
nor U11918 (N_11918,N_8712,N_8587);
nor U11919 (N_11919,N_7203,N_5982);
and U11920 (N_11920,N_708,N_4715);
or U11921 (N_11921,N_477,N_3717);
nand U11922 (N_11922,N_4070,N_8224);
or U11923 (N_11923,N_4809,N_2040);
and U11924 (N_11924,N_5376,N_7409);
nand U11925 (N_11925,N_6660,N_489);
or U11926 (N_11926,N_6005,N_9471);
nand U11927 (N_11927,N_8198,N_84);
and U11928 (N_11928,N_2006,N_3126);
xnor U11929 (N_11929,N_3967,N_1697);
nor U11930 (N_11930,N_6681,N_1154);
nor U11931 (N_11931,N_6355,N_4176);
and U11932 (N_11932,N_1260,N_7799);
or U11933 (N_11933,N_4296,N_5391);
nand U11934 (N_11934,N_2059,N_3295);
or U11935 (N_11935,N_7891,N_1098);
xnor U11936 (N_11936,N_8838,N_7390);
nor U11937 (N_11937,N_9518,N_4539);
or U11938 (N_11938,N_5050,N_1890);
or U11939 (N_11939,N_9918,N_8758);
or U11940 (N_11940,N_6905,N_9233);
nor U11941 (N_11941,N_1123,N_7127);
and U11942 (N_11942,N_5945,N_3945);
xnor U11943 (N_11943,N_6471,N_6746);
nor U11944 (N_11944,N_2242,N_3841);
or U11945 (N_11945,N_3354,N_1211);
nor U11946 (N_11946,N_9049,N_7505);
or U11947 (N_11947,N_5498,N_6038);
nand U11948 (N_11948,N_5173,N_5212);
or U11949 (N_11949,N_4184,N_1782);
nor U11950 (N_11950,N_6163,N_4484);
nor U11951 (N_11951,N_2304,N_5806);
xor U11952 (N_11952,N_9555,N_1354);
or U11953 (N_11953,N_2344,N_840);
nor U11954 (N_11954,N_3135,N_5715);
nor U11955 (N_11955,N_749,N_4527);
nor U11956 (N_11956,N_3147,N_9499);
and U11957 (N_11957,N_8739,N_656);
nor U11958 (N_11958,N_6361,N_6534);
xor U11959 (N_11959,N_3307,N_4831);
and U11960 (N_11960,N_8871,N_9743);
xor U11961 (N_11961,N_1896,N_66);
and U11962 (N_11962,N_1905,N_5201);
xnor U11963 (N_11963,N_4060,N_7597);
xnor U11964 (N_11964,N_5929,N_9997);
and U11965 (N_11965,N_9553,N_836);
or U11966 (N_11966,N_7754,N_4187);
nor U11967 (N_11967,N_2528,N_4021);
xor U11968 (N_11968,N_3888,N_6882);
or U11969 (N_11969,N_8435,N_1142);
xor U11970 (N_11970,N_1249,N_9904);
or U11971 (N_11971,N_3774,N_4664);
and U11972 (N_11972,N_8889,N_1452);
nor U11973 (N_11973,N_9169,N_7216);
nand U11974 (N_11974,N_4028,N_7717);
and U11975 (N_11975,N_7976,N_1902);
or U11976 (N_11976,N_7952,N_7878);
nor U11977 (N_11977,N_2610,N_4730);
nor U11978 (N_11978,N_6875,N_8238);
and U11979 (N_11979,N_4164,N_75);
and U11980 (N_11980,N_1159,N_3095);
or U11981 (N_11981,N_9807,N_4140);
or U11982 (N_11982,N_1351,N_2414);
and U11983 (N_11983,N_4015,N_2570);
xnor U11984 (N_11984,N_1095,N_4425);
or U11985 (N_11985,N_8704,N_9359);
nand U11986 (N_11986,N_4690,N_6641);
and U11987 (N_11987,N_9042,N_8228);
nor U11988 (N_11988,N_8499,N_9919);
or U11989 (N_11989,N_1846,N_5897);
nor U11990 (N_11990,N_6900,N_1216);
or U11991 (N_11991,N_9631,N_9979);
nand U11992 (N_11992,N_6501,N_9927);
and U11993 (N_11993,N_9373,N_7386);
xnor U11994 (N_11994,N_9797,N_4150);
xor U11995 (N_11995,N_5083,N_3553);
nand U11996 (N_11996,N_9652,N_1589);
nor U11997 (N_11997,N_2635,N_4902);
nand U11998 (N_11998,N_3108,N_7518);
xnor U11999 (N_11999,N_7377,N_5075);
nor U12000 (N_12000,N_1372,N_5448);
nand U12001 (N_12001,N_8077,N_4909);
xor U12002 (N_12002,N_1593,N_5813);
nand U12003 (N_12003,N_394,N_6862);
or U12004 (N_12004,N_5547,N_4720);
nor U12005 (N_12005,N_4795,N_1327);
nor U12006 (N_12006,N_7833,N_7149);
and U12007 (N_12007,N_6035,N_4180);
nand U12008 (N_12008,N_7729,N_8547);
xor U12009 (N_12009,N_2301,N_1550);
and U12010 (N_12010,N_9318,N_4616);
and U12011 (N_12011,N_9312,N_3821);
nor U12012 (N_12012,N_4392,N_1822);
and U12013 (N_12013,N_2776,N_4624);
xor U12014 (N_12014,N_7433,N_6061);
xnor U12015 (N_12015,N_738,N_442);
nor U12016 (N_12016,N_5027,N_4151);
xor U12017 (N_12017,N_9735,N_1028);
nand U12018 (N_12018,N_4907,N_5178);
and U12019 (N_12019,N_4932,N_254);
xor U12020 (N_12020,N_6968,N_3960);
nand U12021 (N_12021,N_1026,N_9021);
xor U12022 (N_12022,N_4678,N_3253);
xor U12023 (N_12023,N_3744,N_289);
nand U12024 (N_12024,N_1674,N_1402);
or U12025 (N_12025,N_790,N_5871);
nor U12026 (N_12026,N_9625,N_5984);
or U12027 (N_12027,N_4938,N_5854);
or U12028 (N_12028,N_6506,N_8786);
or U12029 (N_12029,N_5022,N_8303);
or U12030 (N_12030,N_6378,N_7291);
and U12031 (N_12031,N_7640,N_375);
nor U12032 (N_12032,N_1888,N_5332);
or U12033 (N_12033,N_856,N_4327);
nand U12034 (N_12034,N_6868,N_3746);
nand U12035 (N_12035,N_9955,N_466);
or U12036 (N_12036,N_2634,N_7209);
xor U12037 (N_12037,N_3868,N_3965);
xor U12038 (N_12038,N_7819,N_5688);
nor U12039 (N_12039,N_4258,N_2939);
or U12040 (N_12040,N_543,N_479);
nand U12041 (N_12041,N_9820,N_7251);
nor U12042 (N_12042,N_9623,N_4143);
or U12043 (N_12043,N_717,N_773);
and U12044 (N_12044,N_7290,N_8666);
xnor U12045 (N_12045,N_5772,N_6295);
nand U12046 (N_12046,N_8049,N_9104);
nor U12047 (N_12047,N_4081,N_2378);
and U12048 (N_12048,N_419,N_7314);
or U12049 (N_12049,N_6060,N_876);
nand U12050 (N_12050,N_1972,N_2806);
nor U12051 (N_12051,N_3005,N_4288);
nand U12052 (N_12052,N_2628,N_1109);
xor U12053 (N_12053,N_7897,N_8906);
and U12054 (N_12054,N_7434,N_3590);
nor U12055 (N_12055,N_6726,N_8066);
nand U12056 (N_12056,N_5526,N_2573);
or U12057 (N_12057,N_8650,N_2804);
or U12058 (N_12058,N_2212,N_2816);
xor U12059 (N_12059,N_8629,N_2492);
nand U12060 (N_12060,N_6267,N_4934);
or U12061 (N_12061,N_5824,N_421);
nor U12062 (N_12062,N_8896,N_4697);
nand U12063 (N_12063,N_6972,N_3417);
or U12064 (N_12064,N_8997,N_9660);
or U12065 (N_12065,N_6424,N_9365);
nand U12066 (N_12066,N_8525,N_6285);
and U12067 (N_12067,N_9087,N_7109);
or U12068 (N_12068,N_8796,N_9187);
and U12069 (N_12069,N_9609,N_5235);
xnor U12070 (N_12070,N_9633,N_4137);
nand U12071 (N_12071,N_8012,N_7650);
and U12072 (N_12072,N_3342,N_9379);
xor U12073 (N_12073,N_5501,N_5809);
nand U12074 (N_12074,N_8504,N_2553);
nor U12075 (N_12075,N_8743,N_5427);
xnor U12076 (N_12076,N_525,N_5790);
xnor U12077 (N_12077,N_5161,N_3838);
nor U12078 (N_12078,N_4916,N_194);
nor U12079 (N_12079,N_3805,N_9079);
and U12080 (N_12080,N_5263,N_4930);
or U12081 (N_12081,N_5337,N_6736);
xnor U12082 (N_12082,N_1992,N_3701);
or U12083 (N_12083,N_8167,N_312);
and U12084 (N_12084,N_8839,N_1551);
xnor U12085 (N_12085,N_4865,N_1940);
and U12086 (N_12086,N_9096,N_2891);
xnor U12087 (N_12087,N_7874,N_6376);
xnor U12088 (N_12088,N_2158,N_4356);
nor U12089 (N_12089,N_6977,N_2017);
nor U12090 (N_12090,N_1895,N_6697);
or U12091 (N_12091,N_6140,N_1756);
or U12092 (N_12092,N_4280,N_9089);
or U12093 (N_12093,N_458,N_5428);
nor U12094 (N_12094,N_1898,N_8701);
and U12095 (N_12095,N_7063,N_4927);
nor U12096 (N_12096,N_9102,N_7653);
or U12097 (N_12097,N_9255,N_3635);
and U12098 (N_12098,N_7472,N_9615);
nor U12099 (N_12099,N_2418,N_5153);
or U12100 (N_12100,N_994,N_4546);
nor U12101 (N_12101,N_2268,N_5197);
or U12102 (N_12102,N_8252,N_2923);
xnor U12103 (N_12103,N_4526,N_2963);
and U12104 (N_12104,N_3177,N_3133);
or U12105 (N_12105,N_966,N_3689);
and U12106 (N_12106,N_4947,N_1335);
nor U12107 (N_12107,N_2231,N_2947);
xnor U12108 (N_12108,N_9942,N_2828);
xnor U12109 (N_12109,N_6481,N_4139);
xor U12110 (N_12110,N_4764,N_6964);
nor U12111 (N_12111,N_1467,N_3231);
xnor U12112 (N_12112,N_9827,N_7510);
or U12113 (N_12113,N_826,N_7566);
or U12114 (N_12114,N_5740,N_6443);
or U12115 (N_12115,N_4733,N_9580);
xnor U12116 (N_12116,N_1476,N_8577);
and U12117 (N_12117,N_922,N_2618);
and U12118 (N_12118,N_1484,N_9556);
and U12119 (N_12119,N_7955,N_4644);
or U12120 (N_12120,N_6362,N_3901);
xor U12121 (N_12121,N_1172,N_9928);
or U12122 (N_12122,N_5184,N_7228);
nand U12123 (N_12123,N_8694,N_5109);
xnor U12124 (N_12124,N_9617,N_174);
or U12125 (N_12125,N_7143,N_6918);
or U12126 (N_12126,N_5996,N_2183);
nand U12127 (N_12127,N_2107,N_8343);
xor U12128 (N_12128,N_8236,N_9714);
nand U12129 (N_12129,N_9527,N_5601);
nor U12130 (N_12130,N_9331,N_2187);
nor U12131 (N_12131,N_9498,N_8865);
and U12132 (N_12132,N_652,N_4020);
nor U12133 (N_12133,N_2385,N_6333);
nand U12134 (N_12134,N_2844,N_8149);
nor U12135 (N_12135,N_5279,N_901);
nand U12136 (N_12136,N_5518,N_7903);
and U12137 (N_12137,N_8985,N_5923);
and U12138 (N_12138,N_7271,N_3262);
xor U12139 (N_12139,N_2626,N_7741);
nor U12140 (N_12140,N_1747,N_2953);
nand U12141 (N_12141,N_5360,N_5530);
nand U12142 (N_12142,N_1520,N_4565);
nor U12143 (N_12143,N_4222,N_415);
nor U12144 (N_12144,N_5597,N_7943);
or U12145 (N_12145,N_169,N_171);
nor U12146 (N_12146,N_4093,N_1766);
or U12147 (N_12147,N_907,N_5642);
nand U12148 (N_12148,N_2067,N_7934);
and U12149 (N_12149,N_2591,N_1099);
and U12150 (N_12150,N_4805,N_8773);
xor U12151 (N_12151,N_7406,N_4226);
nand U12152 (N_12152,N_8275,N_7902);
nand U12153 (N_12153,N_4744,N_629);
nor U12154 (N_12154,N_1540,N_9549);
nand U12155 (N_12155,N_50,N_2071);
and U12156 (N_12156,N_5836,N_5875);
nand U12157 (N_12157,N_817,N_6215);
xnor U12158 (N_12158,N_6693,N_9142);
nor U12159 (N_12159,N_7448,N_626);
or U12160 (N_12160,N_2637,N_9775);
nand U12161 (N_12161,N_7820,N_3595);
nor U12162 (N_12162,N_2142,N_2874);
xnor U12163 (N_12163,N_5728,N_1350);
xor U12164 (N_12164,N_1368,N_8088);
nor U12165 (N_12165,N_3226,N_9456);
nor U12166 (N_12166,N_809,N_2927);
nor U12167 (N_12167,N_7083,N_3110);
nand U12168 (N_12168,N_3337,N_1349);
and U12169 (N_12169,N_1054,N_2473);
nand U12170 (N_12170,N_6795,N_6173);
nand U12171 (N_12171,N_4406,N_4716);
nor U12172 (N_12172,N_7713,N_4366);
xnor U12173 (N_12173,N_7256,N_7654);
or U12174 (N_12174,N_292,N_119);
nand U12175 (N_12175,N_9929,N_8010);
nor U12176 (N_12176,N_7299,N_9017);
or U12177 (N_12177,N_6445,N_9072);
nand U12178 (N_12178,N_4263,N_1769);
or U12179 (N_12179,N_3954,N_4090);
xnor U12180 (N_12180,N_9776,N_8280);
and U12181 (N_12181,N_5071,N_698);
xor U12182 (N_12182,N_813,N_8502);
and U12183 (N_12183,N_5044,N_2894);
and U12184 (N_12184,N_7022,N_69);
nand U12185 (N_12185,N_7770,N_4818);
nand U12186 (N_12186,N_3775,N_8760);
xor U12187 (N_12187,N_762,N_9266);
nor U12188 (N_12188,N_2600,N_7161);
and U12189 (N_12189,N_6700,N_55);
and U12190 (N_12190,N_407,N_4864);
nand U12191 (N_12191,N_9636,N_5327);
and U12192 (N_12192,N_450,N_6330);
or U12193 (N_12193,N_8881,N_5522);
nor U12194 (N_12194,N_2742,N_7283);
nor U12195 (N_12195,N_5371,N_3535);
and U12196 (N_12196,N_3169,N_6823);
xor U12197 (N_12197,N_9340,N_3060);
nand U12198 (N_12198,N_7187,N_3634);
or U12199 (N_12199,N_2409,N_3878);
nor U12200 (N_12200,N_8689,N_9097);
xnor U12201 (N_12201,N_745,N_641);
nor U12202 (N_12202,N_5685,N_9818);
nor U12203 (N_12203,N_5445,N_2448);
xor U12204 (N_12204,N_3088,N_6664);
nor U12205 (N_12205,N_7526,N_7188);
nand U12206 (N_12206,N_8820,N_9465);
and U12207 (N_12207,N_4646,N_763);
nand U12208 (N_12208,N_703,N_2020);
or U12209 (N_12209,N_1968,N_2693);
nand U12210 (N_12210,N_447,N_3602);
and U12211 (N_12211,N_8044,N_8415);
or U12212 (N_12212,N_4308,N_8878);
and U12213 (N_12213,N_1930,N_8540);
nand U12214 (N_12214,N_1082,N_8904);
xor U12215 (N_12215,N_4741,N_7541);
and U12216 (N_12216,N_33,N_2168);
nand U12217 (N_12217,N_6222,N_7744);
and U12218 (N_12218,N_3128,N_7917);
or U12219 (N_12219,N_1693,N_3682);
and U12220 (N_12220,N_4783,N_9054);
xor U12221 (N_12221,N_6493,N_223);
nand U12222 (N_12222,N_620,N_8774);
or U12223 (N_12223,N_7401,N_4209);
nor U12224 (N_12224,N_3968,N_7675);
nor U12225 (N_12225,N_3191,N_5313);
nand U12226 (N_12226,N_4309,N_1600);
or U12227 (N_12227,N_7268,N_5294);
nand U12228 (N_12228,N_4707,N_8130);
and U12229 (N_12229,N_9999,N_3283);
nor U12230 (N_12230,N_188,N_4100);
and U12231 (N_12231,N_5879,N_900);
nor U12232 (N_12232,N_4877,N_6967);
or U12233 (N_12233,N_8709,N_5214);
or U12234 (N_12234,N_825,N_7005);
nand U12235 (N_12235,N_6936,N_6190);
nor U12236 (N_12236,N_5707,N_8484);
nand U12237 (N_12237,N_7559,N_3479);
or U12238 (N_12238,N_3856,N_1096);
nor U12239 (N_12239,N_5664,N_760);
nor U12240 (N_12240,N_9967,N_6341);
and U12241 (N_12241,N_3269,N_9953);
or U12242 (N_12242,N_8514,N_3507);
and U12243 (N_12243,N_665,N_298);
or U12244 (N_12244,N_2869,N_1710);
and U12245 (N_12245,N_8527,N_5681);
xor U12246 (N_12246,N_3155,N_7369);
or U12247 (N_12247,N_7108,N_521);
and U12248 (N_12248,N_221,N_2053);
xnor U12249 (N_12249,N_6334,N_3912);
and U12250 (N_12250,N_2321,N_8808);
nor U12251 (N_12251,N_283,N_6259);
or U12252 (N_12252,N_3710,N_804);
or U12253 (N_12253,N_8779,N_499);
xnor U12254 (N_12254,N_6782,N_3284);
or U12255 (N_12255,N_7611,N_5758);
xnor U12256 (N_12256,N_9346,N_9791);
and U12257 (N_12257,N_8736,N_8165);
nor U12258 (N_12258,N_1698,N_2749);
xnor U12259 (N_12259,N_7738,N_4499);
and U12260 (N_12260,N_788,N_8832);
or U12261 (N_12261,N_6472,N_5781);
or U12262 (N_12262,N_1692,N_4046);
or U12263 (N_12263,N_649,N_6467);
nand U12264 (N_12264,N_4666,N_6103);
and U12265 (N_12265,N_3617,N_8364);
xnor U12266 (N_12266,N_2153,N_5846);
or U12267 (N_12267,N_3601,N_4115);
nor U12268 (N_12268,N_1144,N_1073);
nand U12269 (N_12269,N_3140,N_1286);
nor U12270 (N_12270,N_2747,N_7877);
or U12271 (N_12271,N_1044,N_1626);
and U12272 (N_12272,N_3646,N_1015);
nor U12273 (N_12273,N_51,N_7694);
and U12274 (N_12274,N_5351,N_216);
or U12275 (N_12275,N_2047,N_838);
nor U12276 (N_12276,N_7173,N_8909);
nand U12277 (N_12277,N_7418,N_1043);
nor U12278 (N_12278,N_9875,N_8175);
nor U12279 (N_12279,N_3330,N_1127);
or U12280 (N_12280,N_3527,N_593);
nand U12281 (N_12281,N_871,N_670);
or U12282 (N_12282,N_1988,N_3688);
and U12283 (N_12283,N_9298,N_6737);
nand U12284 (N_12284,N_8553,N_3199);
xor U12285 (N_12285,N_1056,N_7021);
and U12286 (N_12286,N_2322,N_5922);
and U12287 (N_12287,N_4436,N_8174);
nor U12288 (N_12288,N_1289,N_2991);
and U12289 (N_12289,N_1941,N_5118);
nor U12290 (N_12290,N_3146,N_1591);
nand U12291 (N_12291,N_978,N_5246);
nand U12292 (N_12292,N_8472,N_3404);
nand U12293 (N_12293,N_3315,N_928);
xor U12294 (N_12294,N_5472,N_8849);
nand U12295 (N_12295,N_8158,N_5433);
nand U12296 (N_12296,N_9963,N_2682);
and U12297 (N_12297,N_7638,N_6597);
and U12298 (N_12298,N_4602,N_1609);
xnor U12299 (N_12299,N_3831,N_3759);
nor U12300 (N_12300,N_3982,N_2609);
nand U12301 (N_12301,N_527,N_3385);
xnor U12302 (N_12302,N_5473,N_490);
nor U12303 (N_12303,N_8267,N_6811);
xor U12304 (N_12304,N_8273,N_1221);
nor U12305 (N_12305,N_861,N_6251);
xnor U12306 (N_12306,N_2085,N_5992);
xnor U12307 (N_12307,N_3761,N_9587);
nand U12308 (N_12308,N_5215,N_1610);
and U12309 (N_12309,N_8099,N_8453);
or U12310 (N_12310,N_8960,N_2449);
xnor U12311 (N_12311,N_1607,N_4725);
and U12312 (N_12312,N_3915,N_7711);
xor U12313 (N_12313,N_9101,N_5650);
or U12314 (N_12314,N_5300,N_8626);
and U12315 (N_12315,N_3848,N_2981);
and U12316 (N_12316,N_391,N_7747);
xnor U12317 (N_12317,N_7371,N_8103);
nand U12318 (N_12318,N_6990,N_1606);
or U12319 (N_12319,N_7045,N_3809);
or U12320 (N_12320,N_8126,N_5550);
xor U12321 (N_12321,N_3729,N_2843);
nand U12322 (N_12322,N_2375,N_3711);
xnor U12323 (N_12323,N_5171,N_8692);
xnor U12324 (N_12324,N_3134,N_5195);
xnor U12325 (N_12325,N_646,N_6850);
and U12326 (N_12326,N_2741,N_76);
nand U12327 (N_12327,N_1981,N_9982);
xor U12328 (N_12328,N_2721,N_2996);
and U12329 (N_12329,N_3305,N_7026);
nor U12330 (N_12330,N_7354,N_8685);
xor U12331 (N_12331,N_3125,N_2647);
and U12332 (N_12332,N_8265,N_8534);
or U12333 (N_12333,N_5465,N_9393);
and U12334 (N_12334,N_9739,N_1794);
xnor U12335 (N_12335,N_8211,N_6296);
and U12336 (N_12336,N_9742,N_5377);
or U12337 (N_12337,N_8144,N_9198);
nor U12338 (N_12338,N_1547,N_6350);
nor U12339 (N_12339,N_5640,N_2995);
nor U12340 (N_12340,N_7110,N_7630);
and U12341 (N_12341,N_7966,N_1406);
xnor U12342 (N_12342,N_5798,N_3697);
nor U12343 (N_12343,N_4995,N_5949);
nor U12344 (N_12344,N_5536,N_2475);
and U12345 (N_12345,N_1798,N_9326);
or U12346 (N_12346,N_1479,N_6108);
nand U12347 (N_12347,N_2518,N_6354);
nor U12348 (N_12348,N_1754,N_564);
or U12349 (N_12349,N_4564,N_362);
xnor U12350 (N_12350,N_6527,N_7911);
or U12351 (N_12351,N_7850,N_6415);
xnor U12352 (N_12352,N_7671,N_1014);
or U12353 (N_12353,N_1820,N_1524);
nor U12354 (N_12354,N_9568,N_5609);
and U12355 (N_12355,N_904,N_860);
or U12356 (N_12356,N_7071,N_4626);
nor U12357 (N_12357,N_9783,N_233);
nand U12358 (N_12358,N_8643,N_7335);
or U12359 (N_12359,N_8223,N_4457);
nand U12360 (N_12360,N_5361,N_4943);
or U12361 (N_12361,N_4377,N_6107);
and U12362 (N_12362,N_4286,N_4829);
and U12363 (N_12363,N_5396,N_5952);
and U12364 (N_12364,N_1903,N_5735);
or U12365 (N_12365,N_9968,N_3597);
nand U12366 (N_12366,N_2582,N_2186);
or U12367 (N_12367,N_2440,N_8923);
nor U12368 (N_12368,N_6788,N_2802);
xor U12369 (N_12369,N_9110,N_7515);
nor U12370 (N_12370,N_8118,N_7737);
nor U12371 (N_12371,N_8617,N_4738);
nor U12372 (N_12372,N_4984,N_2631);
and U12373 (N_12373,N_3042,N_7028);
and U12374 (N_12374,N_8971,N_4332);
xnor U12375 (N_12375,N_2974,N_8863);
nor U12376 (N_12376,N_7894,N_1858);
and U12377 (N_12377,N_2339,N_6288);
nor U12378 (N_12378,N_7475,N_4989);
or U12379 (N_12379,N_2309,N_2079);
and U12380 (N_12380,N_7969,N_6303);
and U12381 (N_12381,N_3873,N_433);
nand U12382 (N_12382,N_1979,N_2120);
or U12383 (N_12383,N_3083,N_6025);
or U12384 (N_12384,N_9105,N_4799);
and U12385 (N_12385,N_2604,N_7066);
and U12386 (N_12386,N_8677,N_3569);
and U12387 (N_12387,N_5253,N_3204);
nor U12388 (N_12388,N_8929,N_2464);
or U12389 (N_12389,N_1111,N_6030);
and U12390 (N_12390,N_496,N_4062);
or U12391 (N_12391,N_5317,N_1008);
xnor U12392 (N_12392,N_9574,N_2259);
and U12393 (N_12393,N_7915,N_9998);
nand U12394 (N_12394,N_8584,N_1864);
and U12395 (N_12395,N_5440,N_735);
and U12396 (N_12396,N_7138,N_1761);
or U12397 (N_12397,N_7382,N_7549);
nor U12398 (N_12398,N_556,N_7471);
xnor U12399 (N_12399,N_1526,N_5850);
and U12400 (N_12400,N_1079,N_6911);
and U12401 (N_12401,N_6607,N_2751);
nor U12402 (N_12402,N_1165,N_6143);
nand U12403 (N_12403,N_6171,N_4162);
xnor U12404 (N_12404,N_9434,N_5739);
nand U12405 (N_12405,N_7942,N_2394);
xor U12406 (N_12406,N_8317,N_2852);
xor U12407 (N_12407,N_627,N_3747);
nand U12408 (N_12408,N_4855,N_7949);
and U12409 (N_12409,N_2310,N_6465);
xor U12410 (N_12410,N_6969,N_1137);
nand U12411 (N_12411,N_6431,N_1745);
or U12412 (N_12412,N_8942,N_121);
and U12413 (N_12413,N_5092,N_7410);
nand U12414 (N_12414,N_8456,N_2036);
or U12415 (N_12415,N_7569,N_3972);
xnor U12416 (N_12416,N_9554,N_7718);
or U12417 (N_12417,N_909,N_5537);
nor U12418 (N_12418,N_2076,N_624);
nand U12419 (N_12419,N_5481,N_7002);
and U12420 (N_12420,N_4142,N_3314);
or U12421 (N_12421,N_7909,N_7884);
and U12422 (N_12422,N_7169,N_3858);
nand U12423 (N_12423,N_6238,N_4034);
and U12424 (N_12424,N_4694,N_7950);
nand U12425 (N_12425,N_6379,N_4213);
or U12426 (N_12426,N_1862,N_731);
nand U12427 (N_12427,N_2334,N_191);
xnor U12428 (N_12428,N_2133,N_1791);
nand U12429 (N_12429,N_5224,N_1409);
xnor U12430 (N_12430,N_806,N_7436);
and U12431 (N_12431,N_8653,N_7596);
nor U12432 (N_12432,N_4301,N_9165);
nand U12433 (N_12433,N_9452,N_7460);
xor U12434 (N_12434,N_8093,N_1622);
xnor U12435 (N_12435,N_137,N_7474);
nor U12436 (N_12436,N_4994,N_5777);
or U12437 (N_12437,N_2823,N_4770);
nand U12438 (N_12438,N_6277,N_7860);
or U12439 (N_12439,N_8530,N_4721);
nor U12440 (N_12440,N_6950,N_3780);
xor U12441 (N_12441,N_6248,N_1101);
xor U12442 (N_12442,N_6897,N_3585);
xnor U12443 (N_12443,N_7551,N_4852);
xor U12444 (N_12444,N_7119,N_7863);
and U12445 (N_12445,N_3087,N_8166);
nand U12446 (N_12446,N_4567,N_1065);
or U12447 (N_12447,N_5057,N_2015);
nand U12448 (N_12448,N_9341,N_8113);
nand U12449 (N_12449,N_1801,N_7362);
nor U12450 (N_12450,N_6065,N_8452);
and U12451 (N_12451,N_9219,N_1694);
or U12452 (N_12452,N_4368,N_6096);
xor U12453 (N_12453,N_1728,N_1612);
nor U12454 (N_12454,N_5862,N_1352);
nor U12455 (N_12455,N_2592,N_1386);
nor U12456 (N_12456,N_4132,N_1105);
and U12457 (N_12457,N_3442,N_1170);
nor U12458 (N_12458,N_2248,N_8266);
nor U12459 (N_12459,N_8394,N_4876);
nor U12460 (N_12460,N_4269,N_6074);
nor U12461 (N_12461,N_4610,N_6921);
and U12462 (N_12462,N_8755,N_7513);
and U12463 (N_12463,N_2395,N_9851);
nor U12464 (N_12464,N_2130,N_453);
or U12465 (N_12465,N_6842,N_1638);
or U12466 (N_12466,N_4606,N_6632);
nor U12467 (N_12467,N_9876,N_5115);
or U12468 (N_12468,N_468,N_5577);
xnor U12469 (N_12469,N_8401,N_135);
or U12470 (N_12470,N_3666,N_855);
or U12471 (N_12471,N_7798,N_9601);
or U12472 (N_12472,N_2335,N_8996);
xnor U12473 (N_12473,N_8116,N_6057);
nor U12474 (N_12474,N_7774,N_4906);
and U12475 (N_12475,N_9973,N_9737);
or U12476 (N_12476,N_5402,N_1650);
nor U12477 (N_12477,N_2323,N_2247);
and U12478 (N_12478,N_8059,N_8961);
and U12479 (N_12479,N_4810,N_392);
nand U12480 (N_12480,N_1806,N_5767);
nand U12481 (N_12481,N_547,N_9226);
or U12482 (N_12482,N_8300,N_5633);
nand U12483 (N_12483,N_8640,N_8836);
nand U12484 (N_12484,N_7359,N_1711);
and U12485 (N_12485,N_5475,N_6769);
nand U12486 (N_12486,N_4411,N_7288);
xnor U12487 (N_12487,N_6952,N_4063);
nand U12488 (N_12488,N_8148,N_4514);
and U12489 (N_12489,N_2115,N_571);
or U12490 (N_12490,N_5847,N_7453);
nor U12491 (N_12491,N_212,N_9932);
and U12492 (N_12492,N_7836,N_5827);
nand U12493 (N_12493,N_2537,N_7455);
and U12494 (N_12494,N_5898,N_3642);
xor U12495 (N_12495,N_3516,N_2504);
and U12496 (N_12496,N_4762,N_9841);
nand U12497 (N_12497,N_9681,N_3052);
nor U12498 (N_12498,N_3847,N_6329);
xnor U12499 (N_12499,N_2110,N_2933);
nand U12500 (N_12500,N_4595,N_4563);
xnor U12501 (N_12501,N_2956,N_6423);
and U12502 (N_12502,N_4000,N_8908);
nor U12503 (N_12503,N_9826,N_3287);
or U12504 (N_12504,N_662,N_431);
nor U12505 (N_12505,N_9355,N_1164);
nor U12506 (N_12506,N_2562,N_6858);
and U12507 (N_12507,N_3555,N_1379);
or U12508 (N_12508,N_46,N_4239);
nand U12509 (N_12509,N_699,N_3178);
and U12510 (N_12510,N_8182,N_8589);
xor U12511 (N_12511,N_6194,N_3863);
or U12512 (N_12512,N_7186,N_8094);
or U12513 (N_12513,N_1977,N_7971);
and U12514 (N_12514,N_2613,N_9906);
and U12515 (N_12515,N_286,N_3105);
or U12516 (N_12516,N_3100,N_4185);
xor U12517 (N_12517,N_5257,N_4068);
nand U12518 (N_12518,N_1061,N_4449);
or U12519 (N_12519,N_6611,N_8074);
or U12520 (N_12520,N_4374,N_2692);
nand U12521 (N_12521,N_9977,N_2367);
nand U12522 (N_12522,N_6620,N_841);
nand U12523 (N_12523,N_9137,N_4985);
xnor U12524 (N_12524,N_9175,N_4788);
xnor U12525 (N_12525,N_844,N_4729);
xor U12526 (N_12526,N_5672,N_3184);
or U12527 (N_12527,N_9679,N_1318);
nand U12528 (N_12528,N_8064,N_7214);
nand U12529 (N_12529,N_5048,N_756);
nor U12530 (N_12530,N_2297,N_2648);
xor U12531 (N_12531,N_4703,N_1356);
xor U12532 (N_12532,N_5555,N_5444);
and U12533 (N_12533,N_7483,N_5870);
nor U12534 (N_12534,N_471,N_9417);
xor U12535 (N_12535,N_8292,N_7222);
xor U12536 (N_12536,N_1316,N_251);
or U12537 (N_12537,N_2180,N_5106);
or U12538 (N_12538,N_7981,N_3106);
and U12539 (N_12539,N_8535,N_6480);
nand U12540 (N_12540,N_4867,N_6987);
xnor U12541 (N_12541,N_3647,N_3980);
and U12542 (N_12542,N_6999,N_6146);
nand U12543 (N_12543,N_729,N_8297);
xnor U12544 (N_12544,N_614,N_5623);
nor U12545 (N_12545,N_2500,N_7719);
xnor U12546 (N_12546,N_8765,N_5684);
or U12547 (N_12547,N_3561,N_9381);
and U12548 (N_12548,N_4920,N_2605);
and U12549 (N_12549,N_7536,N_9949);
nor U12550 (N_12550,N_8768,N_2539);
and U12551 (N_12551,N_4962,N_2519);
nor U12552 (N_12552,N_2857,N_1149);
or U12553 (N_12553,N_4200,N_7358);
nand U12554 (N_12554,N_11,N_5073);
and U12555 (N_12555,N_6926,N_6503);
or U12556 (N_12556,N_6716,N_5602);
nand U12557 (N_12557,N_8034,N_113);
nand U12558 (N_12558,N_6798,N_8691);
xor U12559 (N_12559,N_4926,N_5055);
nand U12560 (N_12560,N_9420,N_1844);
xor U12561 (N_12561,N_2347,N_1193);
nand U12562 (N_12562,N_9718,N_3480);
or U12563 (N_12563,N_6682,N_343);
nor U12564 (N_12564,N_833,N_4265);
nor U12565 (N_12565,N_8101,N_6090);
nand U12566 (N_12566,N_1324,N_8974);
and U12567 (N_12567,N_631,N_6371);
nor U12568 (N_12568,N_9184,N_2262);
and U12569 (N_12569,N_5213,N_2960);
or U12570 (N_12570,N_3499,N_4364);
xnor U12571 (N_12571,N_6049,N_4685);
nor U12572 (N_12572,N_9435,N_5784);
nor U12573 (N_12573,N_2563,N_2478);
or U12574 (N_12574,N_1269,N_7467);
nor U12575 (N_12575,N_5395,N_6630);
xor U12576 (N_12576,N_2665,N_7004);
or U12577 (N_12577,N_3388,N_6665);
xnor U12578 (N_12578,N_4333,N_7281);
or U12579 (N_12579,N_6018,N_2444);
or U12580 (N_12580,N_6183,N_7605);
nor U12581 (N_12581,N_484,N_2696);
or U12582 (N_12582,N_9329,N_5329);
xor U12583 (N_12583,N_2420,N_883);
nand U12584 (N_12584,N_9503,N_4345);
or U12585 (N_12585,N_1951,N_983);
nor U12586 (N_12586,N_663,N_5914);
and U12587 (N_12587,N_5030,N_3343);
and U12588 (N_12588,N_1280,N_915);
nor U12589 (N_12589,N_3443,N_4815);
nand U12590 (N_12590,N_956,N_9595);
xor U12591 (N_12591,N_3103,N_6282);
nand U12592 (N_12592,N_17,N_7144);
xor U12593 (N_12593,N_8470,N_8596);
xnor U12594 (N_12594,N_5268,N_178);
nor U12595 (N_12595,N_1944,N_4352);
nand U12596 (N_12596,N_1385,N_2199);
nor U12597 (N_12597,N_6076,N_303);
and U12598 (N_12598,N_6458,N_1493);
or U12599 (N_12599,N_9678,N_5276);
nor U12600 (N_12600,N_5012,N_1986);
nand U12601 (N_12601,N_1046,N_8710);
or U12602 (N_12602,N_1420,N_5525);
xnor U12603 (N_12603,N_9509,N_4581);
nor U12604 (N_12604,N_4740,N_8980);
xnor U12605 (N_12605,N_28,N_5309);
or U12606 (N_12606,N_2337,N_3002);
or U12607 (N_12607,N_6657,N_4509);
and U12608 (N_12608,N_1080,N_2798);
nor U12609 (N_12609,N_9309,N_5574);
or U12610 (N_12610,N_6807,N_8762);
xor U12611 (N_12611,N_3055,N_3073);
or U12612 (N_12612,N_2866,N_9256);
nor U12613 (N_12613,N_7178,N_701);
or U12614 (N_12614,N_9295,N_8879);
or U12615 (N_12615,N_6131,N_3846);
xor U12616 (N_12616,N_1990,N_2295);
nor U12617 (N_12617,N_4255,N_3926);
and U12618 (N_12618,N_1502,N_4779);
or U12619 (N_12619,N_3509,N_761);
nand U12620 (N_12620,N_4849,N_3616);
and U12621 (N_12621,N_3224,N_2685);
and U12622 (N_12622,N_6302,N_989);
and U12623 (N_12623,N_5492,N_9389);
xor U12624 (N_12624,N_653,N_6732);
nand U12625 (N_12625,N_9533,N_2235);
nand U12626 (N_12626,N_3865,N_9544);
and U12627 (N_12627,N_302,N_2229);
xor U12628 (N_12628,N_3611,N_8423);
or U12629 (N_12629,N_746,N_8717);
and U12630 (N_12630,N_8119,N_5578);
xnor U12631 (N_12631,N_4117,N_7699);
nand U12632 (N_12632,N_5185,N_7609);
nor U12633 (N_12633,N_8011,N_2851);
xnor U12634 (N_12634,N_9618,N_8811);
nor U12635 (N_12635,N_1396,N_8729);
xnor U12636 (N_12636,N_7982,N_5524);
or U12637 (N_12637,N_5315,N_6993);
nand U12638 (N_12638,N_3185,N_9510);
nand U12639 (N_12639,N_8769,N_5958);
xnor U12640 (N_12640,N_5496,N_1566);
or U12641 (N_12641,N_452,N_5186);
nand U12642 (N_12642,N_3657,N_4541);
or U12643 (N_12643,N_7196,N_7226);
nor U12644 (N_12644,N_5062,N_8648);
xnor U12645 (N_12645,N_2282,N_8442);
and U12646 (N_12646,N_57,N_6343);
xnor U12647 (N_12647,N_6307,N_8841);
xnor U12648 (N_12648,N_529,N_1042);
and U12649 (N_12649,N_6179,N_3882);
nor U12650 (N_12650,N_5384,N_5104);
xnor U12651 (N_12651,N_361,N_2681);
nor U12652 (N_12652,N_6360,N_1306);
xnor U12653 (N_12653,N_9399,N_6046);
and U12654 (N_12654,N_748,N_2780);
nand U12655 (N_12655,N_3624,N_561);
xnor U12656 (N_12656,N_4336,N_8800);
nor U12657 (N_12657,N_818,N_9387);
or U12658 (N_12658,N_3834,N_6718);
nor U12659 (N_12659,N_5330,N_991);
nor U12660 (N_12660,N_4145,N_8870);
xor U12661 (N_12661,N_5624,N_2084);
nor U12662 (N_12662,N_6073,N_8451);
and U12663 (N_12663,N_3249,N_5608);
and U12664 (N_12664,N_4026,N_9871);
or U12665 (N_12665,N_2543,N_1013);
xor U12666 (N_12666,N_7601,N_6411);
nor U12667 (N_12667,N_5489,N_4885);
nor U12668 (N_12668,N_1712,N_1215);
nor U12669 (N_12669,N_7334,N_8890);
xnor U12670 (N_12670,N_9938,N_6560);
xor U12671 (N_12671,N_6703,N_3313);
or U12672 (N_12672,N_9749,N_9322);
or U12673 (N_12673,N_6861,N_1583);
nor U12674 (N_12674,N_702,N_5812);
nor U12675 (N_12675,N_8902,N_2207);
nand U12676 (N_12676,N_3995,N_5272);
or U12677 (N_12677,N_5554,N_2091);
xnor U12678 (N_12678,N_3869,N_5677);
or U12679 (N_12679,N_2174,N_9530);
xor U12680 (N_12680,N_852,N_1416);
and U12681 (N_12681,N_4857,N_8178);
or U12682 (N_12682,N_5751,N_8606);
nor U12683 (N_12683,N_8036,N_2118);
and U12684 (N_12684,N_7208,N_2348);
and U12685 (N_12685,N_248,N_3419);
nand U12686 (N_12686,N_2616,N_1984);
nor U12687 (N_12687,N_8310,N_5705);
and U12688 (N_12688,N_2679,N_203);
nor U12689 (N_12689,N_9363,N_1226);
xnor U12690 (N_12690,N_8722,N_9272);
or U12691 (N_12691,N_3724,N_1407);
xnor U12692 (N_12692,N_4439,N_1348);
and U12693 (N_12693,N_3978,N_3081);
and U12694 (N_12694,N_6462,N_9515);
xnor U12695 (N_12695,N_6944,N_32);
nor U12696 (N_12696,N_7304,N_1040);
nor U12697 (N_12697,N_5032,N_9065);
nor U12698 (N_12698,N_3636,N_5080);
nor U12699 (N_12699,N_8072,N_2633);
nor U12700 (N_12700,N_753,N_8141);
nand U12701 (N_12701,N_6441,N_8793);
nand U12702 (N_12702,N_3504,N_21);
nand U12703 (N_12703,N_4853,N_715);
and U12704 (N_12704,N_6464,N_126);
xnor U12705 (N_12705,N_263,N_772);
or U12706 (N_12706,N_3840,N_5142);
nand U12707 (N_12707,N_1341,N_3338);
nor U12708 (N_12708,N_2837,N_3078);
xor U12709 (N_12709,N_2151,N_443);
nor U12710 (N_12710,N_8038,N_2992);
or U12711 (N_12711,N_7491,N_2104);
and U12712 (N_12712,N_3024,N_7576);
xor U12713 (N_12713,N_9677,N_5136);
nand U12714 (N_12714,N_5243,N_2260);
and U12715 (N_12715,N_360,N_5828);
or U12716 (N_12716,N_5177,N_5736);
nand U12717 (N_12717,N_4495,N_2289);
xnor U12718 (N_12718,N_6720,N_2227);
nor U12719 (N_12719,N_3741,N_1683);
xor U12720 (N_12720,N_7728,N_9545);
nand U12721 (N_12721,N_2942,N_1783);
and U12722 (N_12722,N_8399,N_6691);
nor U12723 (N_12723,N_8935,N_7660);
nand U12724 (N_12724,N_2714,N_7001);
nand U12725 (N_12725,N_8466,N_7486);
or U12726 (N_12726,N_8477,N_8829);
nand U12727 (N_12727,N_8153,N_6623);
nor U12728 (N_12728,N_2285,N_6567);
and U12729 (N_12729,N_1092,N_9131);
nand U12730 (N_12730,N_4396,N_428);
or U12731 (N_12731,N_4114,N_8639);
or U12732 (N_12732,N_3207,N_6328);
xnor U12733 (N_12733,N_8609,N_2887);
or U12734 (N_12734,N_9829,N_4035);
nand U12735 (N_12735,N_2270,N_6773);
nand U12736 (N_12736,N_9436,N_8339);
or U12737 (N_12737,N_8676,N_4672);
nor U12738 (N_12738,N_1542,N_7009);
nor U12739 (N_12739,N_3917,N_5141);
or U12740 (N_12740,N_4508,N_5292);
nor U12741 (N_12741,N_859,N_3764);
or U12742 (N_12742,N_2705,N_5719);
and U12743 (N_12743,N_873,N_9046);
or U12744 (N_12744,N_6757,N_6908);
and U12745 (N_12745,N_1340,N_4229);
nand U12746 (N_12746,N_8035,N_6160);
nor U12747 (N_12747,N_3548,N_6982);
or U12748 (N_12748,N_372,N_2873);
xnor U12749 (N_12749,N_68,N_9466);
or U12750 (N_12750,N_6577,N_9411);
or U12751 (N_12751,N_2603,N_8814);
or U12752 (N_12752,N_4760,N_2102);
xor U12753 (N_12753,N_3143,N_6521);
or U12754 (N_12754,N_7896,N_1273);
nand U12755 (N_12755,N_2760,N_5569);
and U12756 (N_12756,N_6752,N_7932);
or U12757 (N_12757,N_8986,N_7327);
and U12758 (N_12758,N_3367,N_9236);
nand U12759 (N_12759,N_6043,N_2520);
nor U12760 (N_12760,N_5488,N_7003);
nor U12761 (N_12761,N_6297,N_19);
or U12762 (N_12762,N_694,N_3357);
xnor U12763 (N_12763,N_1925,N_8200);
or U12764 (N_12764,N_8062,N_8455);
nor U12765 (N_12765,N_4470,N_6484);
nand U12766 (N_12766,N_2290,N_5273);
nand U12767 (N_12767,N_4481,N_1833);
and U12768 (N_12768,N_9259,N_6717);
and U12769 (N_12769,N_9244,N_5014);
and U12770 (N_12770,N_1472,N_6137);
and U12771 (N_12771,N_7931,N_5941);
and U12772 (N_12772,N_3475,N_7150);
nand U12773 (N_12773,N_2101,N_6869);
xor U12774 (N_12774,N_5598,N_4828);
nand U12775 (N_12775,N_9944,N_9978);
and U12776 (N_12776,N_8835,N_9489);
or U12777 (N_12777,N_7055,N_3910);
nor U12778 (N_12778,N_9158,N_4585);
nand U12779 (N_12779,N_3881,N_906);
xnor U12780 (N_12780,N_3576,N_3203);
nor U12781 (N_12781,N_6552,N_9801);
xor U12782 (N_12782,N_3756,N_2112);
xor U12783 (N_12783,N_4201,N_2872);
xor U12784 (N_12784,N_4988,N_2236);
xor U12785 (N_12785,N_4615,N_3257);
nand U12786 (N_12786,N_3054,N_3753);
and U12787 (N_12787,N_7267,N_9846);
or U12788 (N_12788,N_5305,N_9342);
and U12789 (N_12789,N_1878,N_4642);
and U12790 (N_12790,N_6583,N_8355);
nand U12791 (N_12791,N_716,N_5778);
nand U12792 (N_12792,N_9300,N_1345);
and U12793 (N_12793,N_1954,N_1424);
nand U12794 (N_12794,N_2766,N_8404);
and U12795 (N_12795,N_940,N_9238);
nand U12796 (N_12796,N_7765,N_7025);
nor U12797 (N_12797,N_3080,N_5580);
and U12798 (N_12798,N_7215,N_9916);
and U12799 (N_12799,N_1325,N_9058);
nand U12800 (N_12800,N_94,N_7254);
xnor U12801 (N_12801,N_2240,N_7749);
nor U12802 (N_12802,N_6724,N_7023);
xnor U12803 (N_12803,N_8856,N_364);
or U12804 (N_12804,N_5017,N_5217);
nor U12805 (N_12805,N_5175,N_971);
xor U12806 (N_12806,N_3319,N_6864);
and U12807 (N_12807,N_8815,N_3380);
nand U12808 (N_12808,N_4942,N_2961);
and U12809 (N_12809,N_9458,N_3445);
nor U12810 (N_12810,N_5183,N_6159);
xnor U12811 (N_12811,N_6395,N_399);
nand U12812 (N_12812,N_7892,N_658);
or U12813 (N_12813,N_4243,N_9885);
xor U12814 (N_12814,N_9253,N_9336);
xor U12815 (N_12815,N_8921,N_589);
nor U12816 (N_12816,N_5724,N_2457);
nand U12817 (N_12817,N_9167,N_2653);
xnor U12818 (N_12818,N_8955,N_1721);
nor U12819 (N_12819,N_5400,N_4696);
nor U12820 (N_12820,N_7007,N_2993);
nand U12821 (N_12821,N_921,N_5090);
xnor U12822 (N_12822,N_151,N_1339);
and U12823 (N_12823,N_9218,N_3288);
xnor U12824 (N_12824,N_4878,N_4292);
xor U12825 (N_12825,N_6319,N_6227);
and U12826 (N_12826,N_3890,N_1326);
xor U12827 (N_12827,N_3496,N_9823);
or U12828 (N_12828,N_3895,N_5861);
nor U12829 (N_12829,N_539,N_9473);
nand U12830 (N_12830,N_4619,N_8259);
or U12831 (N_12831,N_81,N_3247);
xor U12832 (N_12832,N_6164,N_2461);
xnor U12833 (N_12833,N_4232,N_7986);
nor U12834 (N_12834,N_4533,N_1353);
nand U12835 (N_12835,N_8145,N_4293);
xor U12836 (N_12836,N_2426,N_1460);
nand U12837 (N_12837,N_7555,N_5455);
nor U12838 (N_12838,N_2737,N_6814);
xnor U12839 (N_12839,N_9897,N_9350);
nand U12840 (N_12840,N_8953,N_2642);
or U12841 (N_12841,N_4569,N_8684);
or U12842 (N_12842,N_9424,N_3065);
xnor U12843 (N_12843,N_5979,N_8526);
and U12844 (N_12844,N_7165,N_6828);
xor U12845 (N_12845,N_7128,N_5438);
or U12846 (N_12846,N_1875,N_3379);
nand U12847 (N_12847,N_7658,N_5344);
nor U12848 (N_12848,N_6089,N_7643);
nor U12849 (N_12849,N_1097,N_668);
nand U12850 (N_12850,N_2568,N_4784);
or U12851 (N_12851,N_5491,N_6886);
or U12852 (N_12852,N_3515,N_1742);
or U12853 (N_12853,N_4351,N_5613);
xor U12854 (N_12854,N_5700,N_8117);
and U12855 (N_12855,N_5742,N_5192);
nand U12856 (N_12856,N_2485,N_6338);
nand U12857 (N_12857,N_1023,N_7122);
nand U12858 (N_12858,N_3783,N_3896);
nor U12859 (N_12859,N_1481,N_1261);
nand U12860 (N_12860,N_3187,N_6728);
nand U12861 (N_12861,N_8928,N_5883);
nand U12862 (N_12862,N_2503,N_938);
nand U12863 (N_12863,N_2587,N_7684);
xor U12864 (N_12864,N_6776,N_695);
nand U12865 (N_12865,N_4370,N_2811);
or U12866 (N_12866,N_4092,N_9487);
nor U12867 (N_12867,N_1797,N_874);
or U12868 (N_12868,N_5520,N_3395);
and U12869 (N_12869,N_958,N_6203);
nor U12870 (N_12870,N_8613,N_8030);
or U12871 (N_12871,N_2770,N_6165);
nand U12872 (N_12872,N_3070,N_6234);
or U12873 (N_12873,N_449,N_8579);
or U12874 (N_12874,N_5575,N_411);
and U12875 (N_12875,N_5867,N_4820);
xor U12876 (N_12876,N_6489,N_959);
or U12877 (N_12877,N_8293,N_2813);
xor U12878 (N_12878,N_2509,N_2670);
and U12879 (N_12879,N_8239,N_4992);
and U12880 (N_12880,N_6646,N_6023);
nand U12881 (N_12881,N_4438,N_9370);
xnor U12882 (N_12882,N_6453,N_504);
or U12883 (N_12883,N_7068,N_2450);
or U12884 (N_12884,N_1108,N_9560);
nor U12885 (N_12885,N_8645,N_6485);
and U12886 (N_12886,N_220,N_9265);
nor U12887 (N_12887,N_8084,N_4691);
or U12888 (N_12888,N_4227,N_5255);
xnor U12889 (N_12889,N_7610,N_690);
or U12890 (N_12890,N_1991,N_1000);
xor U12891 (N_12891,N_5414,N_2314);
or U12892 (N_12892,N_6546,N_6161);
nand U12893 (N_12893,N_7587,N_4189);
or U12894 (N_12894,N_462,N_1399);
and U12895 (N_12895,N_6839,N_2651);
or U12896 (N_12896,N_6878,N_6710);
nand U12897 (N_12897,N_3037,N_9621);
nor U12898 (N_12898,N_1560,N_1978);
xor U12899 (N_12899,N_4300,N_1717);
nor U12900 (N_12900,N_2893,N_5845);
or U12901 (N_12901,N_2196,N_2447);
or U12902 (N_12902,N_5619,N_7622);
nand U12903 (N_12903,N_8382,N_8982);
nand U12904 (N_12904,N_5437,N_4531);
and U12905 (N_12905,N_2959,N_7672);
xnor U12906 (N_12906,N_912,N_9335);
nand U12907 (N_12907,N_3693,N_5239);
nor U12908 (N_12908,N_8537,N_1869);
or U12909 (N_12909,N_8192,N_5066);
nor U12910 (N_12910,N_8105,N_6239);
xor U12911 (N_12911,N_9494,N_6678);
nand U12912 (N_12912,N_3278,N_3441);
nand U12913 (N_12913,N_3599,N_6971);
and U12914 (N_12914,N_3229,N_9237);
nor U12915 (N_12915,N_688,N_8702);
nor U12916 (N_12916,N_949,N_5411);
and U12917 (N_12917,N_8642,N_3491);
xor U12918 (N_12918,N_7029,N_8323);
xnor U12919 (N_12919,N_6274,N_5989);
xor U12920 (N_12920,N_7365,N_9778);
or U12921 (N_12921,N_2632,N_9804);
xor U12922 (N_12922,N_1575,N_975);
nor U12923 (N_12923,N_5110,N_141);
or U12924 (N_12924,N_1521,N_8934);
xor U12925 (N_12925,N_8681,N_5643);
and U12926 (N_12926,N_2256,N_1746);
and U12927 (N_12927,N_1907,N_1070);
nor U12928 (N_12928,N_6430,N_1964);
and U12929 (N_12929,N_5422,N_9793);
nor U12930 (N_12930,N_7279,N_9645);
xnor U12931 (N_12931,N_7051,N_9674);
nor U12932 (N_12932,N_4205,N_5765);
xor U12933 (N_12933,N_3455,N_7593);
and U12934 (N_12934,N_2296,N_9257);
nand U12935 (N_12935,N_1993,N_645);
xor U12936 (N_12936,N_1395,N_3460);
nand U12937 (N_12937,N_1965,N_7255);
xor U12938 (N_12938,N_3157,N_475);
and U12939 (N_12939,N_7616,N_9296);
nor U12940 (N_12940,N_8263,N_8428);
and U12941 (N_12941,N_2465,N_4827);
and U12942 (N_12942,N_93,N_8161);
nor U12943 (N_12943,N_487,N_3161);
nor U12944 (N_12944,N_8784,N_1678);
or U12945 (N_12945,N_5005,N_4231);
and U12946 (N_12946,N_3558,N_27);
xnor U12947 (N_12947,N_285,N_3939);
nor U12948 (N_12948,N_4808,N_2178);
and U12949 (N_12949,N_8134,N_9664);
nor U12950 (N_12950,N_9950,N_8190);
nor U12951 (N_12951,N_2146,N_2147);
xnor U12952 (N_12952,N_5907,N_3911);
nand U12953 (N_12953,N_7213,N_3545);
or U12954 (N_12954,N_8559,N_8227);
and U12955 (N_12955,N_7709,N_4580);
or U12956 (N_12956,N_9654,N_7072);
or U12957 (N_12957,N_9557,N_7929);
nand U12958 (N_12958,N_1987,N_9798);
or U12959 (N_12959,N_1047,N_9564);
nand U12960 (N_12960,N_7762,N_5995);
and U12961 (N_12961,N_829,N_5039);
xor U12962 (N_12962,N_960,N_2490);
nand U12963 (N_12963,N_3302,N_6389);
xnor U12964 (N_12964,N_9229,N_6026);
nor U12965 (N_12965,N_5256,N_8479);
nand U12966 (N_12966,N_7449,N_9662);
and U12967 (N_12967,N_6537,N_2482);
nand U12968 (N_12968,N_1936,N_3465);
nand U12969 (N_12969,N_8133,N_2164);
and U12970 (N_12970,N_872,N_7843);
xnor U12971 (N_12971,N_1605,N_1922);
or U12972 (N_12972,N_6206,N_3519);
or U12973 (N_12973,N_2512,N_6312);
or U12974 (N_12974,N_9306,N_8419);
or U12975 (N_12975,N_3436,N_369);
nor U12976 (N_12976,N_2526,N_3160);
nor U12977 (N_12977,N_7470,N_2127);
xor U12978 (N_12978,N_7,N_9323);
and U12979 (N_12979,N_4302,N_4786);
nand U12980 (N_12980,N_6666,N_2864);
or U12981 (N_12981,N_3765,N_6340);
and U12982 (N_12982,N_8366,N_5860);
nand U12983 (N_12983,N_9584,N_3600);
and U12984 (N_12984,N_1657,N_3383);
xnor U12985 (N_12985,N_232,N_2756);
xnor U12986 (N_12986,N_6785,N_3225);
and U12987 (N_12987,N_4486,N_5049);
nand U12988 (N_12988,N_4311,N_1169);
or U12989 (N_12989,N_7972,N_6874);
nand U12990 (N_12990,N_3189,N_6099);
or U12991 (N_12991,N_9246,N_3152);
and U12992 (N_12992,N_2712,N_6223);
or U12993 (N_12993,N_3637,N_7704);
and U12994 (N_12994,N_8039,N_145);
and U12995 (N_12995,N_1083,N_4084);
or U12996 (N_12996,N_4713,N_439);
or U12997 (N_12997,N_7693,N_845);
xor U12998 (N_12998,N_6914,N_615);
or U12999 (N_12999,N_5741,N_2660);
xor U13000 (N_13000,N_4198,N_1602);
and U13001 (N_13001,N_5356,N_5910);
nand U13002 (N_13002,N_9208,N_6000);
or U13003 (N_13003,N_6998,N_9532);
nor U13004 (N_13004,N_5487,N_465);
or U13005 (N_13005,N_6275,N_3554);
nor U13006 (N_13006,N_4601,N_747);
nor U13007 (N_13007,N_5310,N_9684);
or U13008 (N_13008,N_1022,N_9613);
nor U13009 (N_13009,N_6209,N_2502);
nor U13010 (N_13010,N_6890,N_4126);
nor U13011 (N_13011,N_1412,N_7722);
xor U13012 (N_13012,N_7319,N_793);
nor U13013 (N_13013,N_4270,N_6075);
xnor U13014 (N_13014,N_3922,N_8521);
xnor U13015 (N_13015,N_8590,N_3899);
or U13016 (N_13016,N_2027,N_3719);
and U13017 (N_13017,N_445,N_7317);
or U13018 (N_13018,N_2657,N_3321);
and U13019 (N_13019,N_9055,N_5903);
and U13020 (N_13020,N_7992,N_6053);
nor U13021 (N_13021,N_2723,N_6764);
and U13022 (N_13022,N_8877,N_3044);
nand U13023 (N_13023,N_5814,N_881);
xnor U13024 (N_13024,N_8665,N_9764);
or U13025 (N_13025,N_3874,N_9924);
or U13026 (N_13026,N_9888,N_4912);
xor U13027 (N_13027,N_887,N_3378);
and U13028 (N_13028,N_3318,N_8911);
or U13029 (N_13029,N_4303,N_7590);
or U13030 (N_13030,N_6659,N_4007);
xor U13031 (N_13031,N_7532,N_3206);
xor U13032 (N_13032,N_5683,N_6256);
or U13033 (N_13033,N_7921,N_8445);
nand U13034 (N_13034,N_669,N_8987);
and U13035 (N_13035,N_8947,N_5668);
xnor U13036 (N_13036,N_8837,N_2672);
nor U13037 (N_13037,N_7232,N_5797);
nand U13038 (N_13038,N_4048,N_5429);
or U13039 (N_13039,N_5834,N_167);
and U13040 (N_13040,N_9106,N_238);
nand U13041 (N_13041,N_551,N_6017);
xnor U13042 (N_13042,N_9269,N_2376);
xnor U13043 (N_13043,N_7201,N_7528);
nor U13044 (N_13044,N_9667,N_737);
nand U13045 (N_13045,N_8519,N_8970);
and U13046 (N_13046,N_131,N_5718);
nor U13047 (N_13047,N_2412,N_4320);
nor U13048 (N_13048,N_7546,N_605);
nor U13049 (N_13049,N_3728,N_5155);
xnor U13050 (N_13050,N_7035,N_8746);
nand U13051 (N_13051,N_3300,N_4880);
nor U13052 (N_13052,N_7767,N_2074);
xor U13053 (N_13053,N_7685,N_8770);
nor U13054 (N_13054,N_8305,N_4127);
xnor U13055 (N_13055,N_2589,N_8869);
xor U13056 (N_13056,N_2724,N_49);
and U13057 (N_13057,N_8898,N_4556);
and U13058 (N_13058,N_7987,N_5616);
xor U13059 (N_13059,N_6473,N_5830);
nor U13060 (N_13060,N_6037,N_4710);
nand U13061 (N_13061,N_6843,N_8914);
xnor U13062 (N_13062,N_150,N_8218);
nand U13063 (N_13063,N_3336,N_4680);
or U13064 (N_13064,N_4824,N_1171);
nand U13065 (N_13065,N_4304,N_5061);
xor U13066 (N_13066,N_8432,N_5098);
xor U13067 (N_13067,N_1264,N_796);
or U13068 (N_13068,N_8421,N_7452);
xnor U13069 (N_13069,N_5622,N_1620);
and U13070 (N_13070,N_1288,N_6783);
nand U13071 (N_13071,N_5054,N_6780);
or U13072 (N_13072,N_4012,N_6287);
or U13073 (N_13073,N_1837,N_7712);
or U13074 (N_13074,N_8027,N_9632);
or U13075 (N_13075,N_3612,N_4016);
or U13076 (N_13076,N_4166,N_4889);
or U13077 (N_13077,N_4148,N_8757);
and U13078 (N_13078,N_2069,N_4082);
or U13079 (N_13079,N_4501,N_8388);
and U13080 (N_13080,N_8506,N_7752);
or U13081 (N_13081,N_2169,N_9588);
nand U13082 (N_13082,N_9062,N_1680);
nor U13083 (N_13083,N_2985,N_1089);
nor U13084 (N_13084,N_1630,N_6889);
nand U13085 (N_13085,N_752,N_1734);
and U13086 (N_13086,N_5181,N_6148);
xnor U13087 (N_13087,N_7975,N_4287);
nand U13088 (N_13088,N_6078,N_4903);
nand U13089 (N_13089,N_1178,N_6824);
xor U13090 (N_13090,N_9002,N_5977);
and U13091 (N_13091,N_4402,N_420);
and U13092 (N_13092,N_3857,N_5163);
nand U13093 (N_13093,N_515,N_4125);
and U13094 (N_13094,N_3365,N_4588);
and U13095 (N_13095,N_8242,N_5416);
nand U13096 (N_13096,N_40,N_423);
xor U13097 (N_13097,N_3348,N_279);
nor U13098 (N_13098,N_7999,N_9572);
nand U13099 (N_13099,N_7626,N_5210);
and U13100 (N_13100,N_4941,N_4124);
nor U13101 (N_13101,N_2458,N_6901);
nor U13102 (N_13102,N_9451,N_8745);
and U13103 (N_13103,N_9824,N_3803);
or U13104 (N_13104,N_412,N_2753);
xnor U13105 (N_13105,N_1463,N_5457);
or U13106 (N_13106,N_913,N_4262);
nand U13107 (N_13107,N_8686,N_6576);
or U13108 (N_13108,N_5927,N_235);
nor U13109 (N_13109,N_408,N_696);
or U13110 (N_13110,N_9025,N_4474);
or U13111 (N_13111,N_7558,N_7707);
or U13112 (N_13112,N_8631,N_6702);
or U13113 (N_13113,N_5576,N_7013);
or U13114 (N_13114,N_3950,N_6477);
xnor U13115 (N_13115,N_3937,N_142);
xor U13116 (N_13116,N_2007,N_4562);
nor U13117 (N_13117,N_2796,N_426);
nor U13118 (N_13118,N_2986,N_9193);
and U13119 (N_13119,N_3817,N_1450);
xor U13120 (N_13120,N_6185,N_2219);
and U13121 (N_13121,N_6050,N_3943);
and U13122 (N_13122,N_8939,N_902);
nor U13123 (N_13123,N_4513,N_4337);
nor U13124 (N_13124,N_1537,N_2161);
nand U13125 (N_13125,N_7829,N_260);
and U13126 (N_13126,N_9044,N_3431);
nand U13127 (N_13127,N_955,N_5900);
xor U13128 (N_13128,N_9215,N_3810);
nand U13129 (N_13129,N_7714,N_6252);
nand U13130 (N_13130,N_9729,N_684);
xnor U13131 (N_13131,N_5144,N_1759);
xor U13132 (N_13132,N_4182,N_8612);
or U13133 (N_13133,N_5284,N_9905);
nor U13134 (N_13134,N_8611,N_1985);
nand U13135 (N_13135,N_3625,N_1475);
and U13136 (N_13136,N_5639,N_7360);
and U13137 (N_13137,N_9457,N_3849);
and U13138 (N_13138,N_9879,N_4856);
xor U13139 (N_13139,N_8156,N_1788);
nand U13140 (N_13140,N_9127,N_1714);
or U13141 (N_13141,N_7545,N_9649);
nand U13142 (N_13142,N_8910,N_4973);
nor U13143 (N_13143,N_8176,N_9941);
nand U13144 (N_13144,N_7395,N_5723);
xnor U13145 (N_13145,N_9118,N_3223);
or U13146 (N_13146,N_1688,N_8726);
nor U13147 (N_13147,N_7307,N_4674);
or U13148 (N_13148,N_4037,N_3403);
nor U13149 (N_13149,N_9936,N_552);
xnor U13150 (N_13150,N_1197,N_4737);
or U13151 (N_13151,N_2895,N_8033);
nor U13152 (N_13152,N_1119,N_755);
and U13153 (N_13153,N_2597,N_1418);
xor U13154 (N_13154,N_5241,N_2676);
nand U13155 (N_13155,N_1374,N_7603);
and U13156 (N_13156,N_6654,N_3673);
or U13157 (N_13157,N_8006,N_9488);
xnor U13158 (N_13158,N_4382,N_3141);
xor U13159 (N_13159,N_8371,N_2541);
and U13160 (N_13160,N_6866,N_7988);
nor U13161 (N_13161,N_9501,N_1874);
xnor U13162 (N_13162,N_1034,N_8483);
and U13163 (N_13163,N_9551,N_6832);
nand U13164 (N_13164,N_5505,N_5539);
xnor U13165 (N_13165,N_6951,N_7757);
or U13166 (N_13166,N_4211,N_308);
nand U13167 (N_13167,N_4886,N_8071);
nand U13168 (N_13168,N_8804,N_916);
and U13169 (N_13169,N_6766,N_8575);
xor U13170 (N_13170,N_7512,N_8052);
xor U13171 (N_13171,N_4329,N_6320);
nand U13172 (N_13172,N_8700,N_1400);
nor U13173 (N_13173,N_9511,N_1033);
nor U13174 (N_13174,N_2371,N_2919);
nand U13175 (N_13175,N_231,N_345);
xor U13176 (N_13176,N_8449,N_8406);
xnor U13177 (N_13177,N_517,N_2581);
or U13178 (N_13178,N_5585,N_6603);
nand U13179 (N_13179,N_7381,N_650);
or U13180 (N_13180,N_2510,N_6111);
nand U13181 (N_13181,N_2646,N_8771);
nand U13182 (N_13182,N_3691,N_4825);
nand U13183 (N_13183,N_7047,N_8333);
xnor U13184 (N_13184,N_5916,N_7927);
nor U13185 (N_13185,N_157,N_507);
and U13186 (N_13186,N_2058,N_1455);
or U13187 (N_13187,N_5872,N_2089);
xor U13188 (N_13188,N_3316,N_9050);
and U13189 (N_13189,N_9639,N_3631);
nand U13190 (N_13190,N_128,N_8154);
nor U13191 (N_13191,N_7155,N_1544);
xnor U13192 (N_13192,N_805,N_2870);
or U13193 (N_13193,N_1470,N_2819);
and U13194 (N_13194,N_5065,N_609);
or U13195 (N_13195,N_5686,N_2238);
nor U13196 (N_13196,N_2868,N_2817);
and U13197 (N_13197,N_2119,N_8051);
nor U13198 (N_13198,N_7745,N_7211);
nor U13199 (N_13199,N_7154,N_877);
nand U13200 (N_13200,N_4636,N_567);
nor U13201 (N_13201,N_9571,N_9015);
xor U13202 (N_13202,N_6309,N_2667);
or U13203 (N_13203,N_2793,N_62);
and U13204 (N_13204,N_8900,N_7746);
and U13205 (N_13205,N_6585,N_3116);
and U13206 (N_13206,N_1631,N_3750);
and U13207 (N_13207,N_9695,N_2411);
xnor U13208 (N_13208,N_1763,N_294);
xor U13209 (N_13209,N_5727,N_6759);
or U13210 (N_13210,N_7202,N_3430);
nor U13211 (N_13211,N_3227,N_7225);
and U13212 (N_13212,N_8803,N_7899);
nand U13213 (N_13213,N_9519,N_3156);
nand U13214 (N_13214,N_1633,N_8597);
nor U13215 (N_13215,N_3256,N_5169);
nand U13216 (N_13216,N_393,N_4018);
xor U13217 (N_13217,N_3240,N_3384);
or U13218 (N_13218,N_5458,N_931);
and U13219 (N_13219,N_4653,N_202);
nor U13220 (N_13220,N_5254,N_594);
and U13221 (N_13221,N_5127,N_8823);
or U13222 (N_13222,N_4752,N_2373);
nand U13223 (N_13223,N_7615,N_2099);
nor U13224 (N_13224,N_2899,N_3235);
or U13225 (N_13225,N_2968,N_3347);
xor U13226 (N_13226,N_4634,N_8859);
or U13227 (N_13227,N_4346,N_7731);
or U13228 (N_13228,N_1388,N_1707);
or U13229 (N_13229,N_7473,N_8563);
xnor U13230 (N_13230,N_2205,N_8931);
xor U13231 (N_13231,N_4479,N_9640);
nor U13232 (N_13232,N_1865,N_878);
xor U13233 (N_13233,N_7562,N_1946);
or U13234 (N_13234,N_2160,N_9427);
xor U13235 (N_13235,N_9983,N_6661);
nor U13236 (N_13236,N_9593,N_6960);
nand U13237 (N_13237,N_3158,N_765);
nor U13238 (N_13238,N_9917,N_378);
and U13239 (N_13239,N_7910,N_1057);
nor U13240 (N_13240,N_6300,N_963);
nor U13241 (N_13241,N_7842,N_78);
xor U13242 (N_13242,N_3988,N_2661);
and U13243 (N_13243,N_7031,N_8548);
nand U13244 (N_13244,N_2274,N_7662);
and U13245 (N_13245,N_7815,N_3281);
or U13246 (N_13246,N_4172,N_3955);
xnor U13247 (N_13247,N_4643,N_6670);
nor U13248 (N_13248,N_7394,N_6662);
xnor U13249 (N_13249,N_9988,N_473);
and U13250 (N_13250,N_2054,N_129);
nor U13251 (N_13251,N_4778,N_384);
and U13252 (N_13252,N_6904,N_1251);
nor U13253 (N_13253,N_7715,N_6705);
nand U13254 (N_13254,N_5193,N_3492);
and U13255 (N_13255,N_2717,N_5325);
xor U13256 (N_13256,N_3251,N_7027);
or U13257 (N_13257,N_8592,N_8214);
and U13258 (N_13258,N_6711,N_2456);
and U13259 (N_13259,N_3113,N_7923);
and U13260 (N_13260,N_5281,N_1194);
and U13261 (N_13261,N_9697,N_5586);
nor U13262 (N_13262,N_2557,N_8505);
nand U13263 (N_13263,N_12,N_7391);
and U13264 (N_13264,N_6385,N_9865);
and U13265 (N_13265,N_9598,N_4405);
or U13266 (N_13266,N_6765,N_6249);
nand U13267 (N_13267,N_241,N_6291);
xor U13268 (N_13268,N_9493,N_6975);
nand U13269 (N_13269,N_4297,N_7246);
xor U13270 (N_13270,N_1564,N_1224);
xor U13271 (N_13271,N_8892,N_9638);
xnor U13272 (N_13272,N_8083,N_6915);
nor U13273 (N_13273,N_1007,N_4840);
or U13274 (N_13274,N_1621,N_2012);
xnor U13275 (N_13275,N_7221,N_651);
nor U13276 (N_13276,N_7792,N_3987);
xor U13277 (N_13277,N_4420,N_6930);
xor U13278 (N_13278,N_9847,N_8708);
xor U13279 (N_13279,N_2775,N_7175);
xnor U13280 (N_13280,N_1310,N_1793);
nand U13281 (N_13281,N_8250,N_2189);
or U13282 (N_13282,N_3949,N_2128);
nand U13283 (N_13283,N_5006,N_3356);
or U13284 (N_13284,N_6569,N_9048);
and U13285 (N_13285,N_1859,N_1482);
nand U13286 (N_13286,N_2645,N_7096);
and U13287 (N_13287,N_4894,N_4440);
xor U13288 (N_13288,N_4103,N_4022);
xor U13289 (N_13289,N_48,N_4395);
or U13290 (N_13290,N_6363,N_2569);
xor U13291 (N_13291,N_2221,N_6529);
nand U13292 (N_13292,N_6562,N_5352);
nor U13293 (N_13293,N_8959,N_9206);
and U13294 (N_13294,N_980,N_6208);
and U13295 (N_13295,N_6902,N_4579);
or U13296 (N_13296,N_2152,N_7579);
xor U13297 (N_13297,N_3361,N_4977);
xnor U13298 (N_13298,N_7785,N_5056);
and U13299 (N_13299,N_542,N_9732);
nor U13300 (N_13300,N_993,N_9923);
and U13301 (N_13301,N_6721,N_1572);
nor U13302 (N_13302,N_5190,N_1812);
nand U13303 (N_13303,N_591,N_3362);
nand U13304 (N_13304,N_5100,N_4879);
nand U13305 (N_13305,N_3844,N_5469);
and U13306 (N_13306,N_8255,N_4391);
nor U13307 (N_13307,N_5559,N_3705);
nand U13308 (N_13308,N_3406,N_8312);
nand U13309 (N_13309,N_1027,N_3675);
and U13310 (N_13310,N_6543,N_5615);
and U13311 (N_13311,N_2800,N_6891);
xnor U13312 (N_13312,N_6549,N_5072);
nand U13313 (N_13313,N_3866,N_6860);
and U13314 (N_13314,N_8098,N_6927);
nor U13315 (N_13315,N_7351,N_981);
nand U13316 (N_13316,N_4998,N_7043);
nor U13317 (N_13317,N_4469,N_5123);
nand U13318 (N_13318,N_290,N_8047);
xor U13319 (N_13319,N_6928,N_1036);
nor U13320 (N_13320,N_6125,N_6138);
or U13321 (N_13321,N_9859,N_8009);
nand U13322 (N_13322,N_6618,N_2175);
or U13323 (N_13323,N_4622,N_7481);
and U13324 (N_13324,N_3490,N_2362);
and U13325 (N_13325,N_7845,N_7769);
or U13326 (N_13326,N_9310,N_7514);
or U13327 (N_13327,N_8226,N_6121);
or U13328 (N_13328,N_5738,N_2194);
or U13329 (N_13329,N_929,N_5978);
xor U13330 (N_13330,N_886,N_3372);
nand U13331 (N_13331,N_8634,N_1081);
nor U13332 (N_13332,N_3930,N_837);
or U13333 (N_13333,N_9390,N_1760);
and U13334 (N_13334,N_5508,N_9178);
or U13335 (N_13335,N_9486,N_5203);
xor U13336 (N_13336,N_3335,N_7846);
xor U13337 (N_13337,N_9992,N_5043);
nand U13338 (N_13338,N_5618,N_9922);
xnor U13339 (N_13339,N_5514,N_3374);
or U13340 (N_13340,N_8732,N_8884);
nand U13341 (N_13341,N_7872,N_1942);
nand U13342 (N_13342,N_5485,N_8864);
xnor U13343 (N_13343,N_8015,N_1867);
or U13344 (N_13344,N_9337,N_7777);
and U13345 (N_13345,N_678,N_6353);
xnor U13346 (N_13346,N_7461,N_3358);
xor U13347 (N_13347,N_6867,N_7312);
nand U13348 (N_13348,N_9162,N_98);
xor U13349 (N_13349,N_1369,N_8417);
or U13350 (N_13350,N_3619,N_8086);
nand U13351 (N_13351,N_1063,N_9036);
or U13352 (N_13352,N_1469,N_2606);
and U13353 (N_13353,N_7789,N_4279);
nor U13354 (N_13354,N_4675,N_1486);
nand U13355 (N_13355,N_835,N_7387);
nor U13356 (N_13356,N_3794,N_5848);
and U13357 (N_13357,N_7835,N_9581);
nor U13358 (N_13358,N_8023,N_3058);
and U13359 (N_13359,N_714,N_6039);
and U13360 (N_13360,N_8187,N_9307);
xor U13361 (N_13361,N_3376,N_2654);
or U13362 (N_13362,N_2351,N_3806);
and U13363 (N_13363,N_7775,N_2442);
and U13364 (N_13364,N_1087,N_363);
nor U13365 (N_13365,N_9898,N_2474);
or U13366 (N_13366,N_4458,N_5756);
xnor U13367 (N_13367,N_4104,N_6345);
xnor U13368 (N_13368,N_4313,N_4216);
and U13369 (N_13369,N_6558,N_5130);
nand U13370 (N_13370,N_1084,N_1660);
xnor U13371 (N_13371,N_5366,N_8546);
or U13372 (N_13372,N_3650,N_5085);
and U13373 (N_13373,N_5479,N_9810);
and U13374 (N_13374,N_3421,N_1778);
xnor U13375 (N_13375,N_4079,N_7886);
xor U13376 (N_13376,N_968,N_239);
and U13377 (N_13377,N_7948,N_6652);
nor U13378 (N_13378,N_2272,N_5318);
or U13379 (N_13379,N_1234,N_3449);
nor U13380 (N_13380,N_3776,N_6821);
and U13381 (N_13381,N_4631,N_1213);
nor U13382 (N_13382,N_6069,N_6881);
or U13383 (N_13383,N_2586,N_6504);
nand U13384 (N_13384,N_186,N_7864);
and U13385 (N_13385,N_339,N_234);
or U13386 (N_13386,N_4699,N_2911);
nor U13387 (N_13387,N_9986,N_4950);
and U13388 (N_13388,N_7337,N_5528);
nand U13389 (N_13389,N_5148,N_7773);
or U13390 (N_13390,N_8998,N_4259);
nand U13391 (N_13391,N_3239,N_6216);
nor U13392 (N_13392,N_5347,N_8288);
or U13393 (N_13393,N_1840,N_9516);
and U13394 (N_13394,N_2834,N_6436);
nor U13395 (N_13395,N_1765,N_6009);
nand U13396 (N_13396,N_6397,N_2215);
nand U13397 (N_13397,N_1287,N_2230);
and U13398 (N_13398,N_9242,N_3762);
xor U13399 (N_13399,N_8529,N_2114);
xnor U13400 (N_13400,N_5572,N_104);
xnor U13401 (N_13401,N_9596,N_2137);
nor U13402 (N_13402,N_8782,N_8429);
and U13403 (N_13403,N_9575,N_1203);
and U13404 (N_13404,N_4427,N_6269);
and U13405 (N_13405,N_9745,N_124);
nor U13406 (N_13406,N_4620,N_3366);
xnor U13407 (N_13407,N_2934,N_6637);
and U13408 (N_13408,N_9292,N_7772);
nand U13409 (N_13409,N_9375,N_5752);
nand U13410 (N_13410,N_7764,N_1136);
xnor U13411 (N_13411,N_379,N_5571);
and U13412 (N_13412,N_4524,N_3301);
nor U13413 (N_13413,N_5570,N_316);
or U13414 (N_13414,N_803,N_9961);
and U13415 (N_13415,N_6612,N_6651);
nand U13416 (N_13416,N_441,N_5251);
xnor U13417 (N_13417,N_1445,N_6253);
xor U13418 (N_13418,N_541,N_256);
nand U13419 (N_13419,N_3453,N_7867);
or U13420 (N_13420,N_8431,N_4897);
nand U13421 (N_13421,N_5904,N_6085);
and U13422 (N_13422,N_6492,N_5388);
and U13423 (N_13423,N_611,N_7372);
xor U13424 (N_13424,N_88,N_3712);
nand U13425 (N_13425,N_96,N_8433);
or U13426 (N_13426,N_9191,N_112);
nor U13427 (N_13427,N_2585,N_4806);
and U13428 (N_13428,N_4072,N_4475);
or U13429 (N_13429,N_9067,N_950);
nor U13430 (N_13430,N_9813,N_8268);
xnor U13431 (N_13431,N_8352,N_8476);
and U13432 (N_13432,N_6178,N_6917);
or U13433 (N_13433,N_7561,N_3114);
nor U13434 (N_13434,N_3117,N_5966);
or U13435 (N_13435,N_4152,N_9566);
or U13436 (N_13436,N_4056,N_619);
xnor U13437 (N_13437,N_744,N_3416);
nor U13438 (N_13438,N_5418,N_3638);
or U13439 (N_13439,N_1200,N_5226);
and U13440 (N_13440,N_9861,N_8219);
nor U13441 (N_13441,N_8185,N_4276);
or U13442 (N_13442,N_6559,N_8193);
nand U13443 (N_13443,N_5948,N_9040);
or U13444 (N_13444,N_175,N_3326);
nand U13445 (N_13445,N_7840,N_6382);
or U13446 (N_13446,N_8390,N_648);
nand U13447 (N_13447,N_5037,N_8241);
or U13448 (N_13448,N_3771,N_4085);
or U13449 (N_13449,N_2432,N_2062);
nand U13450 (N_13450,N_1268,N_724);
or U13451 (N_13451,N_3594,N_5333);
or U13452 (N_13452,N_2103,N_133);
xor U13453 (N_13453,N_7309,N_3470);
or U13454 (N_13454,N_6447,N_3680);
nand U13455 (N_13455,N_138,N_8400);
nor U13456 (N_13456,N_4433,N_4593);
nor U13457 (N_13457,N_9980,N_2381);
nor U13458 (N_13458,N_1861,N_7100);
nor U13459 (N_13459,N_3517,N_5287);
nor U13460 (N_13460,N_7462,N_9475);
or U13461 (N_13461,N_6883,N_6344);
or U13462 (N_13462,N_5534,N_1640);
or U13463 (N_13463,N_4611,N_957);
or U13464 (N_13464,N_7862,N_7413);
nand U13465 (N_13465,N_3219,N_9107);
xor U13466 (N_13466,N_6635,N_1414);
xor U13467 (N_13467,N_8669,N_1240);
nand U13468 (N_13468,N_8184,N_4463);
nand U13469 (N_13469,N_3531,N_4839);
nand U13470 (N_13470,N_6677,N_942);
xnor U13471 (N_13471,N_5789,N_2678);
nand U13472 (N_13472,N_1975,N_2193);
nand U13473 (N_13473,N_1924,N_9423);
nand U13474 (N_13474,N_2211,N_1983);
xor U13475 (N_13475,N_325,N_1205);
xnor U13476 (N_13476,N_7690,N_2976);
xor U13477 (N_13477,N_6535,N_6906);
or U13478 (N_13478,N_3820,N_2978);
nand U13479 (N_13479,N_5252,N_7137);
nand U13480 (N_13480,N_4862,N_6934);
or U13481 (N_13481,N_9773,N_2595);
or U13482 (N_13482,N_2326,N_8636);
nor U13483 (N_13483,N_7296,N_7642);
nor U13484 (N_13484,N_3220,N_6169);
and U13485 (N_13485,N_4782,N_97);
and U13486 (N_13486,N_1311,N_7129);
nor U13487 (N_13487,N_8749,N_7094);
or U13488 (N_13488,N_1055,N_5451);
and U13489 (N_13489,N_3447,N_4978);
and U13490 (N_13490,N_4939,N_2623);
nand U13491 (N_13491,N_9437,N_7530);
nand U13492 (N_13492,N_3145,N_2973);
xnor U13493 (N_13493,N_4271,N_6768);
or U13494 (N_13494,N_6909,N_2791);
nor U13495 (N_13495,N_459,N_6667);
nand U13496 (N_13496,N_9755,N_7586);
or U13497 (N_13497,N_3610,N_2318);
and U13498 (N_13498,N_6349,N_2998);
nand U13499 (N_13499,N_1762,N_2223);
and U13500 (N_13500,N_6628,N_9780);
or U13501 (N_13501,N_4689,N_3004);
xor U13502 (N_13502,N_8632,N_776);
or U13503 (N_13503,N_5938,N_4807);
nand U13504 (N_13504,N_3975,N_208);
and U13505 (N_13505,N_7102,N_6375);
nor U13506 (N_13506,N_3824,N_8485);
and U13507 (N_13507,N_8776,N_330);
nand U13508 (N_13508,N_9047,N_4999);
nand U13509 (N_13509,N_3537,N_1401);
nand U13510 (N_13510,N_8063,N_7147);
nor U13511 (N_13511,N_7276,N_2308);
nor U13512 (N_13512,N_405,N_2601);
or U13513 (N_13513,N_4982,N_4454);
nand U13514 (N_13514,N_5194,N_7311);
nand U13515 (N_13515,N_579,N_6016);
nand U13516 (N_13516,N_6621,N_4468);
nor U13517 (N_13517,N_7342,N_3681);
or U13518 (N_13518,N_4550,N_1454);
nand U13519 (N_13519,N_3629,N_5105);
nand U13520 (N_13520,N_2340,N_618);
nand U13521 (N_13521,N_6894,N_8682);
nor U13522 (N_13522,N_8478,N_925);
xor U13523 (N_13523,N_815,N_6550);
xor U13524 (N_13524,N_3854,N_946);
xor U13525 (N_13525,N_1091,N_2702);
and U13526 (N_13526,N_7065,N_1298);
or U13527 (N_13527,N_1819,N_8657);
nor U13528 (N_13528,N_3130,N_3574);
nor U13529 (N_13529,N_1825,N_1910);
nand U13530 (N_13530,N_1342,N_2203);
and U13531 (N_13531,N_8616,N_621);
nor U13532 (N_13532,N_332,N_4355);
or U13533 (N_13533,N_7424,N_5196);
or U13534 (N_13534,N_2769,N_1492);
nor U13535 (N_13535,N_395,N_2969);
nor U13536 (N_13536,N_7113,N_2279);
and U13537 (N_13537,N_1377,N_9093);
xor U13538 (N_13538,N_4775,N_5890);
and U13539 (N_13539,N_7101,N_2703);
nor U13540 (N_13540,N_5247,N_9896);
xnor U13541 (N_13541,N_4625,N_5531);
xnor U13542 (N_13542,N_8358,N_1767);
and U13543 (N_13543,N_4011,N_6305);
nor U13544 (N_13544,N_2061,N_29);
nor U13545 (N_13545,N_8235,N_7873);
and U13546 (N_13546,N_6174,N_8332);
nor U13547 (N_13547,N_4518,N_6068);
or U13548 (N_13548,N_7957,N_4758);
xor U13549 (N_13549,N_9286,N_4078);
nand U13550 (N_13550,N_5596,N_1619);
and U13551 (N_13551,N_8788,N_152);
nand U13552 (N_13552,N_3304,N_5383);
xor U13553 (N_13553,N_6133,N_5394);
or U13554 (N_13554,N_676,N_1658);
nand U13555 (N_13555,N_2771,N_3696);
xnor U13556 (N_13556,N_2878,N_1740);
and U13557 (N_13557,N_951,N_8383);
nor U13558 (N_13558,N_8917,N_6236);
nor U13559 (N_13559,N_148,N_9217);
nor U13560 (N_13560,N_6265,N_4540);
nor U13561 (N_13561,N_8209,N_5324);
nand U13562 (N_13562,N_2706,N_4080);
xnor U13563 (N_13563,N_8508,N_9622);
xor U13564 (N_13564,N_6433,N_1265);
nand U13565 (N_13565,N_5711,N_8443);
or U13566 (N_13566,N_7944,N_13);
nand U13567 (N_13567,N_6279,N_7755);
nor U13568 (N_13568,N_5720,N_6313);
nand U13569 (N_13569,N_580,N_7324);
or U13570 (N_13570,N_1456,N_5744);
nor U13571 (N_13571,N_2046,N_617);
or U13572 (N_13572,N_72,N_8172);
nand U13573 (N_13573,N_8257,N_1012);
xnor U13574 (N_13574,N_7464,N_8620);
or U13575 (N_13575,N_3234,N_1383);
xor U13576 (N_13576,N_8777,N_3985);
xnor U13577 (N_13577,N_1405,N_4338);
and U13578 (N_13578,N_3627,N_7286);
xnor U13579 (N_13579,N_7322,N_1911);
xor U13580 (N_13580,N_6336,N_2423);
and U13581 (N_13581,N_644,N_6885);
xor U13582 (N_13582,N_2880,N_1148);
and U13583 (N_13583,N_3587,N_8393);
and U13584 (N_13584,N_1611,N_9469);
nand U13585 (N_13585,N_1897,N_6448);
nor U13586 (N_13586,N_8696,N_36);
xnor U13587 (N_13587,N_5199,N_9529);
and U13588 (N_13588,N_6784,N_704);
xor U13589 (N_13589,N_6690,N_9277);
xor U13590 (N_13590,N_2329,N_3914);
or U13591 (N_13591,N_4460,N_6517);
or U13592 (N_13592,N_7781,N_8545);
nand U13593 (N_13593,N_9702,N_6192);
nor U13594 (N_13594,N_2815,N_6692);
and U13595 (N_13595,N_3786,N_6997);
xnor U13596 (N_13596,N_4766,N_4875);
nand U13597 (N_13597,N_6408,N_8337);
and U13598 (N_13598,N_154,N_801);
nand U13599 (N_13599,N_3069,N_534);
or U13600 (N_13600,N_1277,N_2013);
xor U13601 (N_13601,N_3833,N_5180);
nor U13602 (N_13602,N_1706,N_4761);
nor U13603 (N_13603,N_1642,N_4347);
nor U13604 (N_13604,N_1613,N_6779);
or U13605 (N_13605,N_3409,N_4693);
nor U13606 (N_13606,N_4147,N_340);
or U13607 (N_13607,N_9004,N_751);
xor U13608 (N_13608,N_780,N_1889);
nor U13609 (N_13609,N_9333,N_4284);
and U13610 (N_13610,N_3424,N_6502);
or U13611 (N_13611,N_2303,N_6840);
and U13612 (N_13612,N_9482,N_3228);
nand U13613 (N_13613,N_3971,N_8845);
or U13614 (N_13614,N_9699,N_1731);
nand U13615 (N_13615,N_9892,N_374);
xnor U13616 (N_13616,N_8555,N_8311);
and U13617 (N_13617,N_2805,N_3862);
nor U13618 (N_13618,N_7074,N_3743);
or U13619 (N_13619,N_3559,N_2496);
nor U13620 (N_13620,N_8723,N_3422);
and U13621 (N_13621,N_9386,N_366);
and U13622 (N_13622,N_1254,N_1403);
and U13623 (N_13623,N_595,N_8610);
or U13624 (N_13624,N_4895,N_6377);
or U13625 (N_13625,N_1873,N_2232);
or U13626 (N_13626,N_1039,N_630);
and U13627 (N_13627,N_2847,N_4379);
nor U13628 (N_13628,N_7417,N_3334);
xnor U13629 (N_13629,N_8721,N_565);
xor U13630 (N_13630,N_3501,N_4714);
nand U13631 (N_13631,N_8127,N_7898);
nor U13632 (N_13632,N_9507,N_9012);
xor U13633 (N_13633,N_7400,N_3218);
and U13634 (N_13634,N_5869,N_8994);
or U13635 (N_13635,N_3633,N_5467);
or U13636 (N_13636,N_3951,N_8637);
and U13637 (N_13637,N_3444,N_6200);
and U13638 (N_13638,N_245,N_8464);
nand U13639 (N_13639,N_9913,N_3210);
or U13640 (N_13640,N_5380,N_3819);
nand U13641 (N_13641,N_8627,N_4168);
nor U13642 (N_13642,N_6403,N_5166);
nor U13643 (N_13643,N_3876,N_6809);
or U13644 (N_13644,N_6028,N_3549);
xor U13645 (N_13645,N_867,N_6876);
or U13646 (N_13646,N_5595,N_7889);
and U13647 (N_13647,N_9746,N_7614);
and U13648 (N_13648,N_603,N_2353);
nand U13649 (N_13649,N_5543,N_602);
or U13650 (N_13650,N_5994,N_3510);
or U13651 (N_13651,N_5926,N_7257);
nor U13652 (N_13652,N_8043,N_3758);
or U13653 (N_13653,N_4260,N_8936);
and U13654 (N_13654,N_9123,N_2216);
xor U13655 (N_13655,N_7339,N_546);
and U13656 (N_13656,N_988,N_482);
or U13657 (N_13657,N_6437,N_9514);
nand U13658 (N_13658,N_77,N_9719);
and U13659 (N_13659,N_1038,N_4949);
or U13660 (N_13660,N_4665,N_9862);
xnor U13661 (N_13661,N_1067,N_2022);
xnor U13662 (N_13662,N_5516,N_3797);
nor U13663 (N_13663,N_8972,N_5532);
nor U13664 (N_13664,N_9582,N_1320);
nor U13665 (N_13665,N_2181,N_9221);
xor U13666 (N_13666,N_2614,N_3524);
and U13667 (N_13667,N_6346,N_2052);
nand U13668 (N_13668,N_9357,N_2498);
and U13669 (N_13669,N_742,N_9453);
and U13670 (N_13670,N_25,N_3077);
xnor U13671 (N_13671,N_8173,N_2172);
nand U13672 (N_13672,N_4571,N_952);
nor U13673 (N_13673,N_2554,N_3748);
nor U13674 (N_13674,N_3282,N_4253);
or U13675 (N_13675,N_6230,N_969);
nand U13676 (N_13676,N_3830,N_1233);
nor U13677 (N_13677,N_6822,N_1429);
or U13678 (N_13678,N_5260,N_2945);
and U13679 (N_13679,N_3877,N_8282);
nor U13680 (N_13680,N_4047,N_1669);
nor U13681 (N_13681,N_8469,N_3328);
or U13682 (N_13682,N_3261,N_8386);
xor U13683 (N_13683,N_2391,N_7439);
nor U13684 (N_13684,N_9925,N_6417);
and U13685 (N_13685,N_7123,N_7482);
and U13686 (N_13686,N_3768,N_1774);
nor U13687 (N_13687,N_1232,N_5703);
and U13688 (N_13688,N_6404,N_60);
nand U13689 (N_13689,N_2599,N_5067);
nand U13690 (N_13690,N_3784,N_2768);
xnor U13691 (N_13691,N_9085,N_5288);
and U13692 (N_13692,N_937,N_7236);
or U13693 (N_13693,N_2140,N_9552);
nand U13694 (N_13694,N_4732,N_4002);
nand U13695 (N_13695,N_9316,N_2386);
nor U13696 (N_13696,N_4261,N_7077);
xnor U13697 (N_13697,N_414,N_5387);
and U13698 (N_13698,N_1064,N_8747);
xor U13699 (N_13699,N_5680,N_6937);
xnor U13700 (N_13700,N_5964,N_8775);
and U13701 (N_13701,N_3596,N_5716);
or U13702 (N_13702,N_1199,N_4928);
xor U13703 (N_13703,N_3976,N_7250);
and U13704 (N_13704,N_6995,N_5355);
xnor U13705 (N_13705,N_9401,N_7574);
nand U13706 (N_13706,N_5876,N_1586);
and U13707 (N_13707,N_6714,N_1516);
or U13708 (N_13708,N_7683,N_548);
nor U13709 (N_13709,N_616,N_7347);
nand U13710 (N_13710,N_8045,N_3944);
and U13711 (N_13711,N_317,N_639);
or U13712 (N_13712,N_8291,N_7120);
and U13713 (N_13713,N_2228,N_4793);
and U13714 (N_13714,N_1795,N_404);
nand U13715 (N_13715,N_1709,N_4881);
or U13716 (N_13716,N_9948,N_1757);
nand U13717 (N_13717,N_9505,N_7687);
or U13718 (N_13718,N_3276,N_606);
nor U13719 (N_13719,N_590,N_176);
or U13720 (N_13720,N_8114,N_9821);
nand U13721 (N_13721,N_3252,N_8254);
nand U13722 (N_13722,N_4629,N_2944);
and U13723 (N_13723,N_9328,N_9063);
and U13724 (N_13724,N_5059,N_2204);
or U13725 (N_13725,N_526,N_9538);
nor U13726 (N_13726,N_2655,N_476);
nor U13727 (N_13727,N_8085,N_7529);
xnor U13728 (N_13728,N_540,N_7735);
xor U13729 (N_13729,N_4511,N_584);
xor U13730 (N_13730,N_8868,N_67);
xor U13731 (N_13731,N_9248,N_7443);
nor U13732 (N_13732,N_6044,N_467);
xor U13733 (N_13733,N_1681,N_9736);
xor U13734 (N_13734,N_5149,N_259);
xnor U13735 (N_13735,N_4660,N_5710);
xor U13736 (N_13736,N_3695,N_4455);
xor U13737 (N_13737,N_6786,N_7570);
nand U13738 (N_13738,N_8368,N_8654);
and U13739 (N_13739,N_3699,N_8662);
xnor U13740 (N_13740,N_5556,N_1517);
nor U13741 (N_13741,N_8413,N_5011);
nor U13742 (N_13742,N_6580,N_9443);
nor U13743 (N_13743,N_189,N_1821);
and U13744 (N_13744,N_9207,N_6771);
or U13745 (N_13745,N_2833,N_2129);
xor U13746 (N_13746,N_196,N_5791);
and U13747 (N_13747,N_5721,N_7793);
and U13748 (N_13748,N_24,N_1923);
nand U13749 (N_13749,N_4845,N_172);
xnor U13750 (N_13750,N_5323,N_9038);
and U13751 (N_13751,N_1117,N_6687);
nand U13752 (N_13752,N_3799,N_1152);
and U13753 (N_13753,N_4727,N_2782);
nor U13754 (N_13754,N_6452,N_5844);
and U13755 (N_13755,N_4317,N_2848);
xor U13756 (N_13756,N_3670,N_4780);
or U13757 (N_13757,N_9275,N_2950);
nor U13758 (N_13758,N_5029,N_456);
and U13759 (N_13759,N_5990,N_9562);
and U13760 (N_13760,N_4792,N_9013);
or U13761 (N_13761,N_3618,N_3089);
xnor U13762 (N_13762,N_8387,N_5277);
nand U13763 (N_13763,N_4315,N_7627);
nor U13764 (N_13764,N_8095,N_6187);
or U13765 (N_13765,N_5258,N_2521);
or U13766 (N_13766,N_4671,N_2056);
xnor U13767 (N_13767,N_8270,N_8573);
nand U13768 (N_13768,N_6147,N_3322);
or U13769 (N_13769,N_6570,N_9448);
xor U13770 (N_13770,N_2936,N_5008);
xnor U13771 (N_13771,N_6954,N_7174);
nor U13772 (N_13772,N_930,N_4394);
or U13773 (N_13773,N_655,N_9629);
xor U13774 (N_13774,N_5112,N_4467);
and U13775 (N_13775,N_5627,N_4043);
nor U13776 (N_13776,N_8024,N_5675);
nor U13777 (N_13777,N_246,N_6751);
and U13778 (N_13778,N_4515,N_9707);
nand U13779 (N_13779,N_7939,N_276);
xor U13780 (N_13780,N_6734,N_9352);
xnor U13781 (N_13781,N_1877,N_284);
or U13782 (N_13782,N_9402,N_3165);
and U13783 (N_13783,N_5091,N_1301);
and U13784 (N_13784,N_8946,N_9550);
xor U13785 (N_13785,N_8880,N_9361);
or U13786 (N_13786,N_500,N_7838);
nand U13787 (N_13787,N_961,N_2055);
and U13788 (N_13788,N_3059,N_4883);
nand U13789 (N_13789,N_5671,N_2364);
nand U13790 (N_13790,N_1624,N_4869);
nor U13791 (N_13791,N_4904,N_9943);
xnor U13792 (N_13792,N_4819,N_7116);
or U13793 (N_13793,N_9696,N_9080);
nand U13794 (N_13794,N_914,N_6015);
or U13795 (N_13795,N_7857,N_1662);
xnor U13796 (N_13796,N_9391,N_9972);
nor U13797 (N_13797,N_9209,N_1749);
xor U13798 (N_13798,N_1879,N_7425);
nand U13799 (N_13799,N_613,N_797);
or U13800 (N_13800,N_9392,N_3149);
and U13801 (N_13801,N_4651,N_6113);
nor U13802 (N_13802,N_3086,N_2731);
nand U13803 (N_13803,N_8888,N_5695);
and U13804 (N_13804,N_8108,N_5286);
xor U13805 (N_13805,N_5960,N_7787);
nor U13806 (N_13806,N_8372,N_1857);
or U13807 (N_13807,N_242,N_9205);
and U13808 (N_13808,N_122,N_1314);
or U13809 (N_13809,N_8965,N_1676);
nand U13810 (N_13810,N_7599,N_198);
or U13811 (N_13811,N_7020,N_728);
nand U13812 (N_13812,N_2750,N_7431);
and U13813 (N_13813,N_1807,N_5095);
or U13814 (N_13814,N_4256,N_7888);
or U13815 (N_13815,N_7039,N_2002);
and U13816 (N_13816,N_4009,N_2109);
xor U13817 (N_13817,N_9634,N_6857);
nand U13818 (N_13818,N_6571,N_9795);
xnor U13819 (N_13819,N_1426,N_2144);
or U13820 (N_13820,N_266,N_8977);
nor U13821 (N_13821,N_5748,N_5551);
xor U13822 (N_13822,N_1736,N_4681);
nor U13823 (N_13823,N_757,N_2338);
and U13824 (N_13824,N_939,N_851);
or U13825 (N_13825,N_1271,N_5280);
and U13826 (N_13826,N_2501,N_4040);
nor U13827 (N_13827,N_300,N_8659);
and U13828 (N_13828,N_2786,N_7344);
and U13829 (N_13829,N_6405,N_6818);
nor U13830 (N_13830,N_6719,N_6024);
nor U13831 (N_13831,N_454,N_7887);
nor U13832 (N_13832,N_9289,N_5674);
nand U13833 (N_13833,N_2331,N_870);
nor U13834 (N_13834,N_608,N_2382);
xor U13835 (N_13835,N_162,N_5016);
nand U13836 (N_13836,N_5233,N_7000);
nand U13837 (N_13837,N_5976,N_7380);
nand U13838 (N_13838,N_6120,N_6157);
and U13839 (N_13839,N_5345,N_3811);
and U13840 (N_13840,N_7598,N_2572);
nand U13841 (N_13841,N_7968,N_7695);
nor U13842 (N_13842,N_1523,N_6182);
xnor U13843 (N_13843,N_8159,N_2201);
and U13844 (N_13844,N_1104,N_9850);
xor U13845 (N_13845,N_8978,N_277);
or U13846 (N_13846,N_2072,N_8272);
nand U13847 (N_13847,N_8249,N_6286);
and U13848 (N_13848,N_6518,N_7019);
nor U13849 (N_13849,N_6359,N_7422);
nor U13850 (N_13850,N_6542,N_6310);
nor U13851 (N_13851,N_3437,N_8019);
xor U13852 (N_13852,N_8448,N_9412);
nor U13853 (N_13853,N_6019,N_3485);
or U13854 (N_13854,N_8322,N_2113);
nor U13855 (N_13855,N_7935,N_8031);
xnor U13856 (N_13856,N_1753,N_4357);
or U13857 (N_13857,N_7595,N_3478);
or U13858 (N_13858,N_570,N_5541);
xor U13859 (N_13859,N_99,N_5454);
or U13860 (N_13860,N_1994,N_3026);
nand U13861 (N_13861,N_3014,N_9425);
and U13862 (N_13862,N_1585,N_9264);
or U13863 (N_13863,N_578,N_9440);
nand U13864 (N_13864,N_6339,N_309);
xor U13865 (N_13865,N_5187,N_1653);
and U13866 (N_13866,N_8377,N_1188);
and U13867 (N_13867,N_7580,N_1255);
nor U13868 (N_13868,N_9704,N_7212);
or U13869 (N_13869,N_4319,N_3770);
and U13870 (N_13870,N_240,N_9231);
or U13871 (N_13871,N_4491,N_6775);
xor U13872 (N_13872,N_4575,N_224);
xnor U13873 (N_13873,N_8833,N_3312);
or U13874 (N_13874,N_9263,N_1737);
and U13875 (N_13875,N_8295,N_9687);
nand U13876 (N_13876,N_6763,N_5933);
and U13877 (N_13877,N_9366,N_8087);
and U13878 (N_13878,N_7428,N_7983);
or U13879 (N_13879,N_416,N_4017);
xor U13880 (N_13880,N_9995,N_3245);
nand U13881 (N_13881,N_977,N_2341);
or U13882 (N_13882,N_1312,N_282);
nor U13883 (N_13883,N_3714,N_7229);
nor U13884 (N_13884,N_4291,N_1945);
nand U13885 (N_13885,N_1425,N_6281);
and U13886 (N_13886,N_1436,N_1387);
or U13887 (N_13887,N_9367,N_2922);
nor U13888 (N_13888,N_2360,N_6584);
xnor U13889 (N_13889,N_3539,N_511);
or U13890 (N_13890,N_6154,N_6644);
nor U13891 (N_13891,N_3190,N_5007);
nand U13892 (N_13892,N_5636,N_2789);
or U13893 (N_13893,N_998,N_3000);
xnor U13894 (N_13894,N_2190,N_4700);
or U13895 (N_13895,N_7591,N_8221);
xnor U13896 (N_13896,N_5754,N_8802);
xnor U13897 (N_13897,N_5381,N_1410);
xor U13898 (N_13898,N_6801,N_6872);
nand U13899 (N_13899,N_3391,N_1541);
nand U13900 (N_13900,N_7691,N_6983);
xnor U13901 (N_13901,N_5471,N_9656);
nand U13902 (N_13902,N_3532,N_7107);
nand U13903 (N_13903,N_8129,N_7521);
xnor U13904 (N_13904,N_8799,N_9779);
nand U13905 (N_13905,N_310,N_3948);
or U13906 (N_13906,N_898,N_7557);
nand U13907 (N_13907,N_3290,N_1118);
nor U13908 (N_13908,N_7353,N_6781);
or U13909 (N_13909,N_4922,N_3350);
and U13910 (N_13910,N_3476,N_5795);
or U13911 (N_13911,N_8489,N_3120);
nand U13912 (N_13912,N_165,N_5133);
and U13913 (N_13913,N_9407,N_718);
xnor U13914 (N_13914,N_3327,N_3667);
nand U13915 (N_13915,N_1005,N_2525);
nor U13916 (N_13916,N_2206,N_4122);
or U13917 (N_13917,N_7583,N_687);
nor U13918 (N_13918,N_430,N_9848);
and U13919 (N_13919,N_1779,N_2941);
and U13920 (N_13920,N_5689,N_4723);
xor U13921 (N_13921,N_3339,N_8718);
and U13922 (N_13922,N_9828,N_758);
nor U13923 (N_13923,N_4154,N_9041);
xor U13924 (N_13924,N_5698,N_5285);
xor U13925 (N_13925,N_9770,N_8605);
or U13926 (N_13926,N_2590,N_3962);
nand U13927 (N_13927,N_8131,N_7608);
nand U13928 (N_13928,N_1508,N_2349);
xnor U13929 (N_13929,N_3072,N_9914);
xnor U13930 (N_13930,N_5407,N_9463);
nand U13931 (N_13931,N_7404,N_1115);
nand U13932 (N_13932,N_6052,N_2999);
nor U13933 (N_13933,N_1768,N_9284);
and U13934 (N_13934,N_5026,N_3401);
and U13935 (N_13935,N_5563,N_2162);
nand U13936 (N_13936,N_4476,N_3413);
nor U13937 (N_13937,N_4435,N_911);
nor U13938 (N_13938,N_7953,N_7879);
nand U13939 (N_13939,N_1528,N_3006);
and U13940 (N_13940,N_1863,N_2818);
nand U13941 (N_13941,N_7681,N_3581);
or U13942 (N_13942,N_4717,N_1468);
nor U13943 (N_13943,N_2790,N_2266);
and U13944 (N_13944,N_7564,N_4887);
xnor U13945 (N_13945,N_1967,N_1649);
xnor U13946 (N_13946,N_3277,N_9010);
and U13947 (N_13947,N_2505,N_1849);
and U13948 (N_13948,N_722,N_5851);
xnor U13949 (N_13949,N_7166,N_2755);
nand U13950 (N_13950,N_5509,N_7415);
and U13951 (N_13951,N_5290,N_3279);
nor U13952 (N_13952,N_7303,N_1563);
or U13953 (N_13953,N_4323,N_7498);
nand U13954 (N_13954,N_9606,N_1448);
or U13955 (N_13955,N_6198,N_5694);
nand U13956 (N_13956,N_6557,N_3181);
nand U13957 (N_13957,N_5560,N_5225);
nand U13958 (N_13958,N_786,N_2454);
and U13959 (N_13959,N_7032,N_2234);
xor U13960 (N_13960,N_5649,N_864);
or U13961 (N_13961,N_1364,N_3311);
and U13962 (N_13962,N_3864,N_7338);
and U13963 (N_13963,N_9188,N_3607);
and U13964 (N_13964,N_6087,N_8212);
nand U13965 (N_13965,N_4384,N_3639);
and U13966 (N_13966,N_1322,N_7230);
or U13967 (N_13967,N_7346,N_4344);
nor U13968 (N_13968,N_5988,N_5792);
or U13969 (N_13969,N_4051,N_1315);
nor U13970 (N_13970,N_3609,N_3274);
xor U13971 (N_13971,N_7114,N_6101);
and U13972 (N_13972,N_7996,N_3162);
and U13973 (N_13973,N_1438,N_7782);
nor U13974 (N_13974,N_35,N_5013);
nand U13975 (N_13975,N_8507,N_7219);
or U13976 (N_13976,N_8411,N_7200);
or U13977 (N_13977,N_5424,N_2896);
nor U13978 (N_13978,N_2551,N_7575);
or U13979 (N_13979,N_5993,N_7176);
and U13980 (N_13980,N_1853,N_7612);
nand U13981 (N_13981,N_7502,N_6804);
and U13982 (N_13982,N_7951,N_5951);
xnor U13983 (N_13983,N_5283,N_406);
nor U13984 (N_13984,N_1596,N_6204);
and U13985 (N_13985,N_7053,N_3961);
and U13986 (N_13986,N_9891,N_5262);
xnor U13987 (N_13987,N_557,N_4768);
nor U13988 (N_13988,N_3222,N_3286);
nor U13989 (N_13989,N_6031,N_5176);
or U13990 (N_13990,N_789,N_7079);
xor U13991 (N_13991,N_5242,N_8403);
and U13992 (N_13992,N_4335,N_7912);
and U13993 (N_13993,N_2929,N_4987);
nand U13994 (N_13994,N_9592,N_3020);
or U13995 (N_13995,N_1278,N_7292);
and U13996 (N_13996,N_278,N_8468);
and U13997 (N_13997,N_5236,N_6406);
xnor U13998 (N_13998,N_5297,N_1020);
nand U13999 (N_13999,N_5338,N_3686);
nand U14000 (N_14000,N_9076,N_1623);
xnor U14001 (N_14001,N_2716,N_3010);
nand U14002 (N_14002,N_9478,N_6770);
nand U14003 (N_14003,N_903,N_4532);
or U14004 (N_14004,N_6955,N_1291);
or U14005 (N_14005,N_7776,N_5340);
nand U14006 (N_14006,N_8893,N_8518);
xor U14007 (N_14007,N_6084,N_8018);
nand U14008 (N_14008,N_7199,N_3241);
nor U14009 (N_14009,N_953,N_7547);
and U14010 (N_14010,N_4996,N_2198);
nand U14011 (N_14011,N_1459,N_4866);
nor U14012 (N_14012,N_1506,N_9090);
nor U14013 (N_14013,N_5126,N_1293);
or U14014 (N_14014,N_7130,N_2593);
or U14015 (N_14015,N_8079,N_9419);
nor U14016 (N_14016,N_9428,N_8246);
nand U14017 (N_14017,N_7300,N_3466);
xnor U14018 (N_14018,N_7484,N_4390);
and U14019 (N_14019,N_5238,N_5678);
or U14020 (N_14020,N_8968,N_9766);
or U14021 (N_14021,N_9996,N_7133);
nand U14022 (N_14022,N_7861,N_2016);
or U14023 (N_14023,N_1960,N_8244);
or U14024 (N_14024,N_2185,N_587);
nor U14025 (N_14025,N_5152,N_2662);
and U14026 (N_14026,N_7504,N_7509);
xnor U14027 (N_14027,N_7264,N_7412);
or U14028 (N_14028,N_8816,N_7618);
nor U14029 (N_14029,N_9836,N_2255);
and U14030 (N_14030,N_2807,N_6331);
and U14031 (N_14031,N_6669,N_4095);
or U14032 (N_14032,N_6606,N_4521);
nand U14033 (N_14033,N_4267,N_5557);
nand U14034 (N_14034,N_3205,N_4097);
xor U14035 (N_14035,N_9480,N_3502);
xor U14036 (N_14036,N_2333,N_1303);
nand U14037 (N_14037,N_6913,N_1281);
and U14038 (N_14038,N_7398,N_8491);
nor U14039 (N_14039,N_4817,N_1961);
nand U14040 (N_14040,N_9433,N_6684);
or U14041 (N_14041,N_3456,N_4066);
nand U14042 (N_14042,N_1615,N_7405);
xnor U14043 (N_14043,N_1549,N_8488);
and U14044 (N_14044,N_1002,N_6007);
nand U14045 (N_14045,N_2948,N_4854);
xor U14046 (N_14046,N_5802,N_9235);
and U14047 (N_14047,N_1006,N_5801);
nand U14048 (N_14048,N_3452,N_6932);
and U14049 (N_14049,N_1121,N_9477);
or U14050 (N_14050,N_2533,N_1465);
or U14051 (N_14051,N_3789,N_4477);
and U14052 (N_14052,N_9224,N_7701);
xnor U14053 (N_14053,N_785,N_4401);
or U14054 (N_14054,N_8436,N_4554);
nor U14055 (N_14055,N_1359,N_8013);
or U14056 (N_14056,N_5234,N_140);
and U14057 (N_14057,N_2643,N_8334);
or U14058 (N_14058,N_2900,N_3027);
nand U14059 (N_14059,N_3079,N_6270);
xnor U14060 (N_14060,N_5028,N_8576);
nor U14061 (N_14061,N_3665,N_4462);
nand U14062 (N_14062,N_1834,N_6258);
and U14063 (N_14063,N_4552,N_5229);
or U14064 (N_14064,N_8848,N_972);
and U14065 (N_14065,N_3031,N_3188);
or U14066 (N_14066,N_3615,N_1259);
xnor U14067 (N_14067,N_1035,N_2005);
nand U14068 (N_14068,N_9439,N_810);
xnor U14069 (N_14069,N_5894,N_2008);
xor U14070 (N_14070,N_2253,N_331);
or U14071 (N_14071,N_5538,N_3669);
nor U14072 (N_14072,N_5503,N_1716);
xor U14073 (N_14073,N_5873,N_2263);
nor U14074 (N_14074,N_8524,N_8331);
or U14075 (N_14075,N_9001,N_8885);
or U14076 (N_14076,N_5293,N_3093);
or U14077 (N_14077,N_9966,N_4186);
nand U14078 (N_14078,N_6923,N_9483);
and U14079 (N_14079,N_3983,N_115);
or U14080 (N_14080,N_9056,N_9868);
nand U14081 (N_14081,N_4734,N_4558);
and U14082 (N_14082,N_4557,N_4183);
or U14083 (N_14083,N_7140,N_5052);
and U14084 (N_14084,N_5825,N_8017);
and U14085 (N_14085,N_8294,N_604);
and U14086 (N_14086,N_2275,N_6070);
and U14087 (N_14087,N_9213,N_9151);
or U14088 (N_14088,N_1241,N_5111);
xnor U14089 (N_14089,N_1962,N_4591);
xor U14090 (N_14090,N_5969,N_9460);
nand U14091 (N_14091,N_5972,N_6202);
xor U14092 (N_14092,N_5124,N_5447);
or U14093 (N_14093,N_6600,N_3292);
nand U14094 (N_14094,N_1848,N_6510);
or U14095 (N_14095,N_4609,N_1577);
nand U14096 (N_14096,N_8862,N_3096);
or U14097 (N_14097,N_4173,N_5771);
or U14098 (N_14098,N_1107,N_3825);
nand U14099 (N_14099,N_492,N_8245);
and U14100 (N_14100,N_3795,N_2957);
nand U14101 (N_14101,N_9225,N_3853);
nand U14102 (N_14102,N_4692,N_2078);
nand U14103 (N_14103,N_9091,N_6610);
and U14104 (N_14104,N_9160,N_3836);
or U14105 (N_14105,N_7497,N_967);
xor U14106 (N_14106,N_6324,N_1691);
or U14107 (N_14107,N_7758,N_3440);
and U14108 (N_14108,N_4702,N_7080);
nor U14109 (N_14109,N_7511,N_8975);
xnor U14110 (N_14110,N_7802,N_1411);
nand U14111 (N_14111,N_2540,N_8492);
nor U14112 (N_14112,N_9787,N_2803);
or U14113 (N_14113,N_7423,N_5298);
nand U14114 (N_14114,N_4965,N_9853);
nand U14115 (N_14115,N_2799,N_6653);
or U14116 (N_14116,N_4935,N_1122);
nand U14117 (N_14117,N_7171,N_4075);
xnor U14118 (N_14118,N_1329,N_3329);
and U14119 (N_14119,N_2278,N_6482);
xnor U14120 (N_14120,N_3048,N_8180);
and U14121 (N_14121,N_9535,N_8397);
xor U14122 (N_14122,N_3745,N_6796);
nor U14123 (N_14123,N_9921,N_9644);
nand U14124 (N_14124,N_9339,N_6979);
nand U14125 (N_14125,N_2063,N_6547);
nand U14126 (N_14126,N_4662,N_2690);
nand U14127 (N_14127,N_6440,N_5657);
and U14128 (N_14128,N_5815,N_9873);
and U14129 (N_14129,N_9504,N_943);
or U14130 (N_14130,N_9815,N_667);
nor U14131 (N_14131,N_7087,N_1933);
xnor U14132 (N_14132,N_5462,N_9145);
xor U14133 (N_14133,N_6933,N_3091);
nand U14134 (N_14134,N_6387,N_1590);
nor U14135 (N_14135,N_2225,N_2598);
nand U14136 (N_14136,N_7447,N_8384);
nand U14137 (N_14137,N_3457,N_4432);
or U14138 (N_14138,N_6422,N_6054);
nand U14139 (N_14139,N_3179,N_7349);
xor U14140 (N_14140,N_1489,N_9706);
nand U14141 (N_14141,N_273,N_2576);
nand U14142 (N_14142,N_2222,N_4834);
nand U14143 (N_14143,N_4471,N_4925);
nor U14144 (N_14144,N_9520,N_6738);
nor U14145 (N_14145,N_1252,N_2073);
and U14146 (N_14146,N_5003,N_8201);
xnor U14147 (N_14147,N_741,N_6342);
xnor U14148 (N_14148,N_8104,N_8350);
nor U14149 (N_14149,N_8405,N_1668);
nand U14150 (N_14150,N_5470,N_3030);
nand U14151 (N_14151,N_9628,N_3626);
nor U14152 (N_14152,N_5168,N_5271);
xor U14153 (N_14153,N_3793,N_7795);
xnor U14154 (N_14154,N_766,N_9168);
and U14155 (N_14155,N_7057,N_2280);
nor U14156 (N_14156,N_8341,N_7396);
nand U14157 (N_14157,N_2195,N_736);
or U14158 (N_14158,N_1276,N_1495);
xnor U14159 (N_14159,N_2898,N_8195);
xnor U14160 (N_14160,N_9290,N_3007);
nor U14161 (N_14161,N_3420,N_323);
or U14162 (N_14162,N_1854,N_7141);
and U14163 (N_14163,N_1382,N_6392);
nor U14164 (N_14164,N_8157,N_3015);
nand U14165 (N_14165,N_5645,N_6852);
and U14166 (N_14166,N_9461,N_3663);
nor U14167 (N_14167,N_8286,N_6407);
xor U14168 (N_14168,N_6680,N_1536);
and U14169 (N_14169,N_8952,N_7893);
xnor U14170 (N_14170,N_7958,N_7937);
nand U14171 (N_14171,N_3932,N_4204);
or U14172 (N_14172,N_6538,N_2355);
and U14173 (N_14173,N_6264,N_9177);
and U14174 (N_14174,N_8111,N_3575);
nor U14175 (N_14175,N_3892,N_1934);
xor U14176 (N_14176,N_4851,N_600);
and U14177 (N_14177,N_7258,N_6575);
or U14178 (N_14178,N_8899,N_9831);
nor U14179 (N_14179,N_9413,N_7736);
nand U14180 (N_14180,N_2032,N_8764);
xor U14181 (N_14181,N_3121,N_3536);
or U14182 (N_14182,N_5939,N_9939);
nor U14183 (N_14183,N_2641,N_1300);
or U14184 (N_14184,N_8638,N_9534);
xor U14185 (N_14185,N_4901,N_1851);
or U14186 (N_14186,N_6456,N_7816);
nand U14187 (N_14187,N_1373,N_5023);
xnor U14188 (N_14188,N_4548,N_8438);
and U14189 (N_14189,N_5963,N_2708);
and U14190 (N_14190,N_4584,N_9095);
and U14191 (N_14191,N_7991,N_550);
and U14192 (N_14192,N_2150,N_7361);
and U14193 (N_14193,N_5950,N_5413);
nor U14194 (N_14194,N_8261,N_6367);
xor U14195 (N_14195,N_9646,N_2028);
xor U14196 (N_14196,N_397,N_9472);
nand U14197 (N_14197,N_1893,N_9449);
xnor U14198 (N_14198,N_8699,N_42);
and U14199 (N_14199,N_8316,N_4923);
nor U14200 (N_14200,N_1434,N_6924);
xnor U14201 (N_14201,N_82,N_1803);
and U14202 (N_14202,N_5587,N_1743);
nor U14203 (N_14203,N_6152,N_4331);
nor U14204 (N_14204,N_9786,N_3407);
nor U14205 (N_14205,N_4039,N_7978);
nand U14206 (N_14206,N_9661,N_6919);
or U14207 (N_14207,N_5296,N_1302);
and U14208 (N_14208,N_6418,N_9122);
nand U14209 (N_14209,N_377,N_9720);
xor U14210 (N_14210,N_6910,N_346);
nor U14211 (N_14211,N_4199,N_6022);
xnor U14212 (N_14212,N_9109,N_1636);
or U14213 (N_14213,N_6761,N_9512);
and U14214 (N_14214,N_7797,N_9607);
nor U14215 (N_14215,N_7438,N_8569);
nand U14216 (N_14216,N_7924,N_3267);
nand U14217 (N_14217,N_9334,N_9204);
xor U14218 (N_14218,N_1272,N_4398);
xor U14219 (N_14219,N_6958,N_5452);
nand U14220 (N_14220,N_7537,N_6419);
nand U14221 (N_14221,N_8976,N_2535);
nor U14222 (N_14222,N_5542,N_3494);
nor U14223 (N_14223,N_4071,N_1973);
and U14224 (N_14224,N_7880,N_3643);
or U14225 (N_14225,N_1652,N_1569);
and U14226 (N_14226,N_5307,N_8674);
nand U14227 (N_14227,N_6841,N_22);
xnor U14228 (N_14228,N_9125,N_6115);
xnor U14229 (N_14229,N_4791,N_3022);
and U14230 (N_14230,N_9459,N_6337);
or U14231 (N_14231,N_1077,N_177);
or U14232 (N_14232,N_1076,N_6609);
nand U14233 (N_14233,N_816,N_4272);
and U14234 (N_14234,N_8170,N_3927);
or U14235 (N_14235,N_8948,N_4428);
and U14236 (N_14236,N_9863,N_6943);
and U14237 (N_14237,N_4964,N_6625);
nand U14238 (N_14238,N_1,N_7664);
nand U14239 (N_14239,N_5170,N_5042);
nor U14240 (N_14240,N_8984,N_4846);
and U14241 (N_14241,N_6941,N_5314);
nor U14242 (N_14242,N_3648,N_8003);
nor U14243 (N_14243,N_3345,N_7092);
or U14244 (N_14244,N_1595,N_1248);
or U14245 (N_14245,N_1832,N_811);
nor U14246 (N_14246,N_2994,N_3994);
or U14247 (N_14247,N_6945,N_9071);
xor U14248 (N_14248,N_210,N_2861);
nor U14249 (N_14249,N_6587,N_4434);
xnor U14250 (N_14250,N_5829,N_8875);
xnor U14251 (N_14251,N_9866,N_8296);
or U14252 (N_14252,N_6744,N_7356);
and U14253 (N_14253,N_1785,N_1969);
and U14254 (N_14254,N_2758,N_6655);
or U14255 (N_14255,N_5182,N_5901);
and U14256 (N_14256,N_4275,N_4726);
nand U14257 (N_14257,N_8938,N_3935);
nor U14258 (N_14258,N_90,N_2305);
and U14259 (N_14259,N_3107,N_1817);
xor U14260 (N_14260,N_227,N_8420);
nor U14261 (N_14261,N_5935,N_1816);
xnor U14262 (N_14262,N_9239,N_7238);
or U14263 (N_14263,N_9895,N_5504);
nor U14264 (N_14264,N_3298,N_6541);
nor U14265 (N_14265,N_7018,N_1614);
or U14266 (N_14266,N_1207,N_6318);
nand U14267 (N_14267,N_7183,N_1173);
and U14268 (N_14268,N_7295,N_4789);
and U14269 (N_14269,N_2106,N_3913);
and U14270 (N_14270,N_6749,N_2850);
nand U14271 (N_14271,N_5912,N_269);
and U14272 (N_14272,N_6594,N_4365);
nand U14273 (N_14273,N_5174,N_9148);
nor U14274 (N_14274,N_2359,N_654);
xor U14275 (N_14275,N_6246,N_9431);
nand U14276 (N_14276,N_9655,N_8109);
nand U14277 (N_14277,N_3808,N_6853);
or U14278 (N_14278,N_3273,N_7240);
or U14279 (N_14279,N_5690,N_8861);
and U14280 (N_14280,N_3506,N_5278);
nand U14281 (N_14281,N_4639,N_7253);
or U14282 (N_14282,N_5343,N_519);
and U14283 (N_14283,N_5406,N_1485);
or U14284 (N_14284,N_299,N_8367);
nand U14285 (N_14285,N_3715,N_3182);
and U14286 (N_14286,N_8733,N_3860);
and U14287 (N_14287,N_4728,N_4316);
xnor U14288 (N_14288,N_7457,N_2489);
xor U14289 (N_14289,N_435,N_7117);
nor U14290 (N_14290,N_6104,N_6980);
or U14291 (N_14291,N_9251,N_5540);
nand U14292 (N_14292,N_2888,N_1433);
and U14293 (N_14293,N_9614,N_261);
or U14294 (N_14294,N_2725,N_3118);
nor U14295 (N_14295,N_1644,N_6102);
nor U14296 (N_14296,N_4159,N_866);
and U14297 (N_14297,N_6640,N_2350);
nor U14298 (N_14298,N_7440,N_3399);
or U14299 (N_14299,N_7085,N_9114);
or U14300 (N_14300,N_7231,N_1375);
nor U14301 (N_14301,N_3661,N_1381);
nand U14302 (N_14302,N_3694,N_9856);
and U14303 (N_14303,N_8279,N_2549);
nor U14304 (N_14304,N_5389,N_8767);
nor U14305 (N_14305,N_9403,N_79);
nor U14306 (N_14306,N_6126,N_8990);
nor U14307 (N_14307,N_3303,N_4195);
nand U14308 (N_14308,N_834,N_319);
and U14309 (N_14309,N_2624,N_3520);
xnor U14310 (N_14310,N_9220,N_8715);
and U14311 (N_14311,N_2783,N_5753);
nor U14312 (N_14312,N_9500,N_14);
and U14313 (N_14313,N_9173,N_9843);
or U14314 (N_14314,N_1126,N_9771);
and U14315 (N_14315,N_3734,N_5167);
xnor U14316 (N_14316,N_8503,N_2023);
and U14317 (N_14317,N_4755,N_9849);
and U14318 (N_14318,N_8283,N_8844);
nand U14319 (N_14319,N_1963,N_8831);
or U14320 (N_14320,N_6365,N_9016);
xnor U14321 (N_14321,N_7689,N_5793);
nor U14322 (N_14322,N_4823,N_2829);
and U14323 (N_14323,N_4708,N_5354);
nand U14324 (N_14324,N_2343,N_9877);
nand U14325 (N_14325,N_5500,N_896);
xor U14326 (N_14326,N_8543,N_2477);
and U14327 (N_14327,N_8328,N_5456);
nand U14328 (N_14328,N_5533,N_6748);
nand U14329 (N_14329,N_1190,N_9822);
xnor U14330 (N_14330,N_674,N_5561);
and U14331 (N_14331,N_7206,N_6475);
or U14332 (N_14332,N_2087,N_9035);
and U14333 (N_14333,N_5529,N_2445);
nand U14334 (N_14334,N_1219,N_8882);
nand U14335 (N_14335,N_7298,N_2544);
xor U14336 (N_14336,N_2176,N_3653);
nor U14337 (N_14337,N_863,N_5135);
xor U14338 (N_14338,N_3959,N_2497);
nand U14339 (N_14339,N_2009,N_6130);
and U14340 (N_14340,N_3823,N_8070);
xor U14341 (N_14341,N_161,N_4083);
and U14342 (N_14342,N_5521,N_7901);
nand U14343 (N_14343,N_5025,N_8348);
or U14344 (N_14344,N_9005,N_6829);
nor U14345 (N_14345,N_5302,N_7990);
or U14346 (N_14346,N_9397,N_8824);
nand U14347 (N_14347,N_5892,N_4208);
nand U14348 (N_14348,N_5120,N_6633);
or U14349 (N_14349,N_2788,N_5944);
xor U14350 (N_14350,N_6410,N_8664);
and U14351 (N_14351,N_7980,N_9947);
nand U14352 (N_14352,N_4445,N_769);
nand U14353 (N_14353,N_9270,N_1237);
nand U14354 (N_14354,N_7974,N_3200);
xor U14355 (N_14355,N_9043,N_1357);
or U14356 (N_14356,N_3412,N_2658);
or U14357 (N_14357,N_8092,N_1724);
nand U14358 (N_14358,N_7523,N_3439);
and U14359 (N_14359,N_2668,N_2511);
nand U14360 (N_14360,N_3893,N_823);
nor U14361 (N_14361,N_3132,N_3716);
or U14362 (N_14362,N_5349,N_5902);
nor U14363 (N_14363,N_8132,N_2574);
or U14364 (N_14364,N_8542,N_7393);
nor U14365 (N_14365,N_2397,N_1950);
nand U14366 (N_14366,N_8958,N_6871);
xor U14367 (N_14367,N_1500,N_7184);
nand U14368 (N_14368,N_9274,N_4656);
xor U14369 (N_14369,N_7632,N_5749);
nor U14370 (N_14370,N_2122,N_3708);
nor U14371 (N_14371,N_4049,N_4001);
xor U14372 (N_14372,N_6793,N_8197);
nor U14373 (N_14373,N_1442,N_8277);
xnor U14374 (N_14374,N_8690,N_5506);
xnor U14375 (N_14375,N_4843,N_1441);
or U14376 (N_14376,N_359,N_444);
and U14377 (N_14377,N_7016,N_8550);
and U14378 (N_14378,N_8121,N_2437);
and U14379 (N_14379,N_5358,N_1474);
nor U14380 (N_14380,N_4981,N_3560);
or U14381 (N_14381,N_1153,N_1836);
or U14382 (N_14382,N_6648,N_6739);
nand U14383 (N_14383,N_7573,N_899);
xor U14384 (N_14384,N_9669,N_7012);
nand U14385 (N_14385,N_3364,N_6715);
nor U14386 (N_14386,N_65,N_249);
and U14387 (N_14387,N_215,N_5849);
or U14388 (N_14388,N_5367,N_5660);
nor U14389 (N_14389,N_820,N_1561);
nand U14390 (N_14390,N_8778,N_532);
xnor U14391 (N_14391,N_2499,N_8876);
nor U14392 (N_14392,N_8060,N_3999);
xnor U14393 (N_14393,N_3242,N_127);
nand U14394 (N_14394,N_9201,N_7821);
xor U14395 (N_14395,N_2081,N_5796);
xor U14396 (N_14396,N_9345,N_5729);
or U14397 (N_14397,N_9202,N_3613);
or U14398 (N_14398,N_5743,N_1996);
xnor U14399 (N_14399,N_8080,N_3111);
nor U14400 (N_14400,N_1238,N_2302);
or U14401 (N_14401,N_3736,N_3148);
nor U14402 (N_14402,N_7205,N_5863);
and U14403 (N_14403,N_7305,N_1887);
or U14404 (N_14404,N_2967,N_2913);
and U14405 (N_14405,N_5099,N_3426);
nand U14406 (N_14406,N_307,N_4098);
or U14407 (N_14407,N_474,N_2824);
or U14408 (N_14408,N_9517,N_270);
xor U14409 (N_14409,N_5157,N_3802);
nor U14410 (N_14410,N_640,N_6756);
nand U14411 (N_14411,N_2306,N_8037);
nand U14412 (N_14412,N_632,N_1916);
xnor U14413 (N_14413,N_2691,N_160);
xnor U14414 (N_14414,N_2486,N_8843);
nand U14415 (N_14415,N_6854,N_8356);
or U14416 (N_14416,N_8189,N_6722);
or U14417 (N_14417,N_6426,N_6001);
or U14418 (N_14418,N_8763,N_2025);
nand U14419 (N_14419,N_2154,N_2921);
nor U14420 (N_14420,N_8309,N_3056);
xnor U14421 (N_14421,N_6802,N_1880);
nor U14422 (N_14422,N_4044,N_8560);
nand U14423 (N_14423,N_7834,N_207);
nor U14424 (N_14424,N_2300,N_8186);
xnor U14425 (N_14425,N_5779,N_4767);
xor U14426 (N_14426,N_5775,N_7783);
or U14427 (N_14427,N_4138,N_9045);
and U14428 (N_14428,N_8365,N_1437);
and U14429 (N_14429,N_6686,N_9537);
nand U14430 (N_14430,N_4430,N_156);
and U14431 (N_14431,N_8794,N_9029);
or U14432 (N_14432,N_1243,N_7446);
nor U14433 (N_14433,N_4446,N_5895);
nand U14434 (N_14434,N_1443,N_295);
or U14435 (N_14435,N_7308,N_6144);
and U14436 (N_14436,N_1582,N_8302);
or U14437 (N_14437,N_6629,N_2192);
and U14438 (N_14438,N_7385,N_7908);
and U14439 (N_14439,N_54,N_5515);
nor U14440 (N_14440,N_9432,N_2433);
or U14441 (N_14441,N_1982,N_4537);
nor U14442 (N_14442,N_633,N_3075);
nand U14443 (N_14443,N_9210,N_5353);
xnor U14444 (N_14444,N_3934,N_3966);
and U14445 (N_14445,N_297,N_7368);
nand U14446 (N_14446,N_2684,N_5291);
nor U14447 (N_14447,N_7036,N_9680);
nand U14448 (N_14448,N_3886,N_4614);
or U14449 (N_14449,N_7115,N_9599);
xnor U14450 (N_14450,N_6083,N_123);
xnor U14451 (N_14451,N_2977,N_6306);
and U14452 (N_14452,N_4367,N_1167);
or U14453 (N_14453,N_1700,N_1242);
xnor U14454 (N_14454,N_5931,N_5420);
nand U14455 (N_14455,N_1158,N_6528);
or U14456 (N_14456,N_3236,N_5119);
nor U14457 (N_14457,N_1247,N_107);
xor U14458 (N_14458,N_5975,N_1262);
nor U14459 (N_14459,N_6235,N_8595);
or U14460 (N_14460,N_3142,N_4891);
nand U14461 (N_14461,N_4858,N_2812);
and U14462 (N_14462,N_3174,N_1422);
xor U14463 (N_14463,N_7260,N_6006);
nand U14464 (N_14464,N_3359,N_642);
xor U14465 (N_14465,N_6674,N_7435);
xnor U14466 (N_14466,N_6989,N_6224);
or U14467 (N_14467,N_2779,N_850);
xnor U14468 (N_14468,N_8515,N_5620);
or U14469 (N_14469,N_3467,N_9126);
xnor U14470 (N_14470,N_9721,N_7964);
nor U14471 (N_14471,N_3800,N_4073);
xnor U14472 (N_14472,N_4408,N_4893);
nor U14473 (N_14473,N_683,N_7871);
nand U14474 (N_14474,N_3511,N_3092);
and U14475 (N_14475,N_267,N_8651);
xnor U14476 (N_14476,N_1555,N_4452);
xor U14477 (N_14477,N_7876,N_4312);
nand U14478 (N_14478,N_2728,N_5102);
nand U14479 (N_14479,N_8164,N_4101);
xor U14480 (N_14480,N_2508,N_4177);
nor U14481 (N_14481,N_4560,N_193);
nor U14482 (N_14482,N_8454,N_6800);
nand U14483 (N_14483,N_7375,N_8501);
and U14484 (N_14484,N_1245,N_905);
nand U14485 (N_14485,N_8480,N_8467);
nor U14486 (N_14486,N_3567,N_8679);
or U14487 (N_14487,N_545,N_5316);
xnor U14488 (N_14488,N_1018,N_2488);
nand U14489 (N_14489,N_2772,N_7315);
nor U14490 (N_14490,N_6136,N_8683);
nor U14491 (N_14491,N_9663,N_1256);
or U14492 (N_14492,N_4747,N_8289);
xor U14493 (N_14493,N_7099,N_3566);
or U14494 (N_14494,N_6948,N_5925);
nand U14495 (N_14495,N_2060,N_1201);
or U14496 (N_14496,N_778,N_1258);
xor U14497 (N_14497,N_9539,N_5261);
nand U14498 (N_14498,N_8042,N_2336);
or U14499 (N_14499,N_4731,N_1811);
and U14500 (N_14500,N_1168,N_8058);
xor U14501 (N_14501,N_8320,N_8741);
xnor U14502 (N_14502,N_4871,N_1116);
nor U14503 (N_14503,N_8536,N_5947);
nor U14504 (N_14504,N_7607,N_2966);
nor U14505 (N_14505,N_250,N_1497);
nor U14506 (N_14506,N_1824,N_6308);
nand U14507 (N_14507,N_5810,N_9765);
or U14508 (N_14508,N_3427,N_9830);
or U14509 (N_14509,N_6966,N_313);
and U14510 (N_14510,N_1587,N_1195);
and U14511 (N_14511,N_6903,N_5265);
nor U14512 (N_14512,N_5121,N_6593);
xnor U14513 (N_14513,N_6498,N_4976);
nand U14514 (N_14514,N_7318,N_3119);
nor U14515 (N_14515,N_2472,N_1773);
or U14516 (N_14516,N_5259,N_6040);
or U14517 (N_14517,N_8057,N_7421);
or U14518 (N_14518,N_8798,N_6673);
xor U14519 (N_14519,N_8630,N_1627);
nor U14520 (N_14520,N_6723,N_6082);
and U14521 (N_14521,N_2906,N_4701);
and U14522 (N_14522,N_3997,N_8517);
or U14523 (N_14523,N_8461,N_8797);
xor U14524 (N_14524,N_4722,N_9670);
nor U14525 (N_14525,N_9692,N_7479);
nor U14526 (N_14526,N_3090,N_9708);
nor U14527 (N_14527,N_8237,N_7926);
or U14528 (N_14528,N_3861,N_4215);
and U14529 (N_14529,N_4798,N_217);
nand U14530 (N_14530,N_1246,N_1304);
or U14531 (N_14531,N_7809,N_3505);
nand U14532 (N_14532,N_7571,N_8169);
nor U14533 (N_14533,N_5308,N_8509);
or U14534 (N_14534,N_3837,N_95);
nor U14535 (N_14535,N_1598,N_1366);
nand U14536 (N_14536,N_5821,N_2368);
or U14537 (N_14537,N_2265,N_1634);
or U14538 (N_14538,N_3656,N_6846);
xor U14539 (N_14539,N_6398,N_2487);
and U14540 (N_14540,N_5223,N_9759);
and U14541 (N_14541,N_4181,N_9081);
nand U14542 (N_14542,N_7306,N_2413);
nand U14543 (N_14543,N_4155,N_2424);
and U14544 (N_14544,N_4219,N_7500);
and U14545 (N_14545,N_2051,N_8410);
or U14546 (N_14546,N_7118,N_5227);
nor U14547 (N_14547,N_5712,N_9747);
and U14548 (N_14548,N_3025,N_9319);
and U14549 (N_14549,N_8633,N_6961);
nor U14550 (N_14550,N_7686,N_8601);
nand U14551 (N_14551,N_2734,N_6631);
or U14552 (N_14552,N_8860,N_6072);
nor U14553 (N_14553,N_6002,N_879);
or U14554 (N_14554,N_9682,N_2964);
nor U14555 (N_14555,N_1723,N_9852);
xor U14556 (N_14556,N_80,N_9619);
nand U14557 (N_14557,N_7293,N_301);
nand U14558 (N_14558,N_9382,N_6755);
xnor U14559 (N_14559,N_1048,N_6820);
nand U14560 (N_14560,N_6212,N_38);
xor U14561 (N_14561,N_4655,N_4385);
and U14562 (N_14562,N_264,N_628);
or U14563 (N_14563,N_4294,N_2890);
nor U14564 (N_14564,N_218,N_660);
nand U14565 (N_14565,N_5392,N_9442);
nor U14566 (N_14566,N_9703,N_8780);
nand U14567 (N_14567,N_5464,N_8380);
nand U14568 (N_14568,N_7476,N_2157);
nand U14569 (N_14569,N_199,N_3392);
xnor U14570 (N_14570,N_1632,N_6671);
and U14571 (N_14571,N_6106,N_3344);
nand U14572 (N_14572,N_9540,N_6488);
nand U14573 (N_14573,N_4812,N_9444);
xnor U14574 (N_14574,N_413,N_7151);
nand U14575 (N_14575,N_3942,N_4064);
and U14576 (N_14576,N_9376,N_2132);
xor U14577 (N_14577,N_7844,N_1274);
nand U14578 (N_14578,N_58,N_4121);
or U14579 (N_14579,N_9886,N_86);
nand U14580 (N_14580,N_3371,N_5589);
xnor U14581 (N_14581,N_3396,N_4133);
or U14582 (N_14582,N_8061,N_910);
nor U14583 (N_14583,N_2021,N_5107);
nor U14584 (N_14584,N_5647,N_6483);
nor U14585 (N_14585,N_4510,N_3582);
and U14586 (N_14586,N_1347,N_1071);
and U14587 (N_14587,N_2744,N_6986);
nand U14588 (N_14588,N_5604,N_610);
or U14589 (N_14589,N_5499,N_846);
xor U14590 (N_14590,N_9380,N_1223);
and U14591 (N_14591,N_4872,N_3180);
or U14592 (N_14592,N_6931,N_682);
and U14593 (N_14593,N_1576,N_6701);
xnor U14594 (N_14594,N_5918,N_9597);
nor U14595 (N_14595,N_3540,N_3725);
and U14596 (N_14596,N_1299,N_5502);
and U14597 (N_14597,N_5852,N_5788);
nand U14598 (N_14598,N_8232,N_6813);
or U14599 (N_14599,N_3423,N_9426);
nand U14600 (N_14600,N_553,N_2283);
xor U14601 (N_14601,N_3351,N_8895);
nor U14602 (N_14602,N_9808,N_2546);
nor U14603 (N_14603,N_7639,N_2875);
xor U14604 (N_14604,N_992,N_9374);
xnor U14605 (N_14605,N_3164,N_4561);
xnor U14606 (N_14606,N_8046,N_3723);
or U14607 (N_14607,N_7628,N_324);
and U14608 (N_14608,N_7269,N_8663);
nor U14609 (N_14609,N_5986,N_4975);
and U14610 (N_14610,N_3233,N_5299);
nand U14611 (N_14611,N_2602,N_9872);
nand U14612 (N_14612,N_4549,N_6145);
or U14613 (N_14613,N_6311,N_6098);
nand U14614 (N_14614,N_2739,N_4361);
xor U14615 (N_14615,N_1294,N_7522);
nor U14616 (N_14616,N_1629,N_764);
nor U14617 (N_14617,N_8089,N_8744);
and U14618 (N_14618,N_5913,N_5321);
xor U14619 (N_14619,N_8473,N_2860);
and U14620 (N_14620,N_1935,N_8872);
nand U14621 (N_14621,N_3578,N_5942);
xnor U14622 (N_14622,N_7620,N_6413);
or U14623 (N_14623,N_3238,N_2513);
xnor U14624 (N_14624,N_8301,N_2312);
nand U14625 (N_14625,N_3850,N_3433);
or U14626 (N_14626,N_8217,N_7272);
and U14627 (N_14627,N_2938,N_6172);
or U14628 (N_14628,N_7073,N_5370);
and U14629 (N_14629,N_2294,N_4363);
nor U14630 (N_14630,N_1604,N_5865);
xor U14631 (N_14631,N_2249,N_4156);
xor U14632 (N_14632,N_3826,N_1532);
or U14633 (N_14633,N_7544,N_8220);
or U14634 (N_14634,N_7011,N_4003);
nor U14635 (N_14635,N_7275,N_1708);
xor U14636 (N_14636,N_6683,N_2476);
xnor U14637 (N_14637,N_9484,N_4024);
nor U14638 (N_14638,N_8389,N_6563);
nor U14639 (N_14639,N_9768,N_8725);
nor U14640 (N_14640,N_5717,N_1758);
or U14641 (N_14641,N_6799,N_9094);
xnor U14642 (N_14642,N_486,N_7098);
xnor U14643 (N_14643,N_9254,N_3991);
or U14644 (N_14644,N_6463,N_1490);
xnor U14645 (N_14645,N_4223,N_1997);
and U14646 (N_14646,N_6284,N_8029);
and U14647 (N_14647,N_6778,N_5953);
and U14648 (N_14648,N_5730,N_2077);
nor U14649 (N_14649,N_8345,N_5275);
xnor U14650 (N_14650,N_7883,N_1147);
or U14651 (N_14651,N_6974,N_200);
nor U14652 (N_14652,N_2481,N_8599);
xor U14653 (N_14653,N_8635,N_4417);
or U14654 (N_14654,N_6825,N_5625);
nor U14655 (N_14655,N_4036,N_842);
nor U14656 (N_14656,N_8703,N_1856);
or U14657 (N_14657,N_7340,N_9675);
nand U14658 (N_14658,N_4228,N_3438);
nand U14659 (N_14659,N_4054,N_1892);
or U14660 (N_14660,N_6996,N_1866);
xnor U14661 (N_14661,N_3782,N_6220);
xnor U14662 (N_14662,N_528,N_7727);
xnor U14663 (N_14663,N_7370,N_8196);
xnor U14664 (N_14664,N_1784,N_2251);
nor U14665 (N_14665,N_586,N_4443);
or U14666 (N_14666,N_9767,N_6327);
nand U14667 (N_14667,N_8660,N_1019);
and U14668 (N_14668,N_7135,N_6335);
nand U14669 (N_14669,N_9152,N_4534);
nand U14670 (N_14670,N_4841,N_6523);
xnor U14671 (N_14671,N_601,N_9074);
nor U14672 (N_14672,N_6844,N_1408);
nand U14673 (N_14673,N_8641,N_4498);
nor U14674 (N_14674,N_3979,N_6898);
and U14675 (N_14675,N_3709,N_6704);
and U14676 (N_14676,N_8697,N_4870);
and U14677 (N_14677,N_2620,N_9196);
or U14678 (N_14678,N_637,N_7852);
or U14679 (N_14679,N_2578,N_108);
nand U14680 (N_14680,N_5889,N_7696);
or U14681 (N_14681,N_9031,N_9299);
xor U14682 (N_14682,N_3306,N_2108);
or U14683 (N_14683,N_3573,N_9388);
nand U14684 (N_14684,N_7582,N_6984);
and U14685 (N_14685,N_8014,N_3920);
or U14686 (N_14686,N_1417,N_6383);
xor U14687 (N_14687,N_771,N_8727);
nand U14688 (N_14688,N_3884,N_3790);
xnor U14689 (N_14689,N_3084,N_5474);
nor U14690 (N_14690,N_8146,N_4240);
and U14691 (N_14691,N_5053,N_2879);
and U14692 (N_14692,N_6195,N_6100);
nor U14693 (N_14693,N_1654,N_1695);
or U14694 (N_14694,N_8381,N_964);
nand U14695 (N_14695,N_6865,N_9657);
or U14696 (N_14696,N_8805,N_7870);
nor U14697 (N_14697,N_9760,N_783);
xor U14698 (N_14698,N_6758,N_6257);
nand U14699 (N_14699,N_3289,N_4751);
xnor U14700 (N_14700,N_7104,N_6792);
or U14701 (N_14701,N_136,N_821);
or U14702 (N_14702,N_7414,N_7637);
or U14703 (N_14703,N_664,N_9915);
and U14704 (N_14704,N_1597,N_1764);
xor U14705 (N_14705,N_9287,N_8905);
nor U14706 (N_14706,N_625,N_9314);
nor U14707 (N_14707,N_8932,N_5648);
or U14708 (N_14708,N_400,N_686);
nor U14709 (N_14709,N_9174,N_7220);
nand U14710 (N_14710,N_4299,N_7252);
nor U14711 (N_14711,N_6289,N_4360);
nor U14712 (N_14712,N_8171,N_4077);
xor U14713 (N_14713,N_9637,N_7496);
xnor U14714 (N_14714,N_2622,N_7058);
nand U14715 (N_14715,N_3168,N_4212);
or U14716 (N_14716,N_5991,N_6012);
nor U14717 (N_14717,N_7445,N_6451);
nand U14718 (N_14718,N_401,N_5426);
xor U14719 (N_14719,N_2261,N_4330);
nand U14720 (N_14720,N_8807,N_6427);
and U14721 (N_14721,N_4488,N_4908);
nand U14722 (N_14722,N_448,N_1346);
nand U14723 (N_14723,N_2542,N_2859);
and U14724 (N_14724,N_2980,N_5937);
or U14725 (N_14725,N_334,N_2392);
nor U14726 (N_14726,N_4749,N_3487);
nand U14727 (N_14727,N_5816,N_672);
xor U14728 (N_14728,N_9816,N_1929);
or U14729 (N_14729,N_6675,N_7442);
nand U14730 (N_14730,N_3144,N_7270);
or U14731 (N_14731,N_2797,N_6175);
nor U14732 (N_14732,N_8347,N_1496);
xnor U14733 (N_14733,N_6156,N_3986);
or U14734 (N_14734,N_6531,N_6920);
nand U14735 (N_14735,N_2044,N_7095);
and U14736 (N_14736,N_7904,N_9870);
nor U14737 (N_14737,N_3718,N_1146);
or U14738 (N_14738,N_1319,N_7124);
xor U14739 (N_14739,N_7134,N_8446);
nor U14740 (N_14740,N_3275,N_6093);
xor U14741 (N_14741,N_451,N_8846);
xor U14742 (N_14742,N_3498,N_9840);
xnor U14743 (N_14743,N_6450,N_7676);
xnor U14744 (N_14744,N_3591,N_636);
nand U14745 (N_14745,N_1275,N_8274);
xnor U14746 (N_14746,N_6469,N_5820);
and U14747 (N_14747,N_8897,N_2435);
or U14748 (N_14748,N_4494,N_9705);
nand U14749 (N_14749,N_5160,N_6638);
xor U14750 (N_14750,N_8243,N_2683);
and U14751 (N_14751,N_5188,N_9011);
nand U14752 (N_14752,N_2984,N_1755);
nand U14753 (N_14753,N_3923,N_9061);
or U14754 (N_14754,N_6742,N_9022);
xor U14755 (N_14755,N_9893,N_461);
xnor U14756 (N_14756,N_4635,N_3816);
nand U14757 (N_14757,N_4773,N_1750);
nand U14758 (N_14758,N_5131,N_3902);
and U14759 (N_14759,N_8137,N_1601);
and U14760 (N_14760,N_4248,N_7160);
nand U14761 (N_14761,N_3209,N_5047);
and U14762 (N_14762,N_1253,N_4058);
nor U14763 (N_14763,N_2208,N_4787);
xnor U14764 (N_14764,N_3973,N_3981);
nand U14765 (N_14765,N_2138,N_1343);
nand U14766 (N_14766,N_9291,N_2971);
xor U14767 (N_14767,N_5164,N_9671);
nor U14768 (N_14768,N_3332,N_5191);
nand U14769 (N_14769,N_4612,N_4353);
nand U14770 (N_14770,N_5985,N_1995);
nor U14771 (N_14771,N_9969,N_5980);
nand U14772 (N_14772,N_6774,N_812);
or U14773 (N_14773,N_329,N_5405);
and U14774 (N_14774,N_2092,N_4658);
nor U14775 (N_14775,N_7459,N_2399);
nand U14776 (N_14776,N_6579,N_530);
xor U14777 (N_14777,N_3464,N_9727);
nand U14778 (N_14778,N_6435,N_4089);
xor U14779 (N_14779,N_919,N_9724);
and U14780 (N_14780,N_2267,N_1282);
nor U14781 (N_14781,N_3778,N_3489);
nand U14782 (N_14782,N_4991,N_9228);
nor U14783 (N_14783,N_3989,N_5001);
or U14784 (N_14784,N_4496,N_8206);
xnor U14785 (N_14785,N_5954,N_3137);
xnor U14786 (N_14786,N_5430,N_9811);
and U14787 (N_14787,N_1539,N_2045);
nand U14788 (N_14788,N_3481,N_4686);
nor U14789 (N_14789,N_5204,N_3202);
nor U14790 (N_14790,N_5393,N_3039);
nand U14791 (N_14791,N_8168,N_3664);
xnor U14792 (N_14792,N_1531,N_6709);
and U14793 (N_14793,N_1336,N_7430);
or U14794 (N_14794,N_9651,N_6962);
xnor U14795 (N_14795,N_2754,N_705);
nor U14796 (N_14796,N_9369,N_1270);
xor U14797 (N_14797,N_9952,N_3843);
xor U14798 (N_14798,N_3028,N_6401);
xor U14799 (N_14799,N_2640,N_7263);
and U14800 (N_14800,N_6003,N_768);
and U14801 (N_14801,N_3801,N_6831);
nor U14802 (N_14802,N_576,N_2588);
and U14803 (N_14803,N_9120,N_5766);
and U14804 (N_14804,N_5666,N_6533);
and U14805 (N_14805,N_7046,N_4178);
nor U14806 (N_14806,N_6141,N_4623);
xnor U14807 (N_14807,N_1789,N_8363);
xor U14808 (N_14808,N_8324,N_7328);
nand U14809 (N_14809,N_1151,N_6772);
nand U14810 (N_14810,N_9149,N_7796);
or U14811 (N_14811,N_4848,N_118);
and U14812 (N_14812,N_882,N_5237);
xor U14813 (N_14813,N_8600,N_2607);
nand U14814 (N_14814,N_4844,N_6449);
xnor U14815 (N_14815,N_5594,N_6588);
and U14816 (N_14816,N_4136,N_7427);
and U14817 (N_14817,N_1953,N_8482);
xor U14818 (N_14818,N_8135,N_1656);
and U14819 (N_14819,N_5658,N_7568);
and U14820 (N_14820,N_3299,N_8552);
nand U14821 (N_14821,N_4171,N_2975);
xor U14822 (N_14822,N_4163,N_779);
xnor U14823 (N_14823,N_759,N_1130);
xor U14824 (N_14824,N_3898,N_5219);
and U14825 (N_14825,N_9462,N_338);
nor U14826 (N_14826,N_6656,N_1025);
xor U14827 (N_14827,N_322,N_4670);
nor U14828 (N_14828,N_5478,N_4298);
and U14829 (N_14829,N_6004,N_6812);
nand U14830 (N_14830,N_9429,N_2460);
nor U14831 (N_14831,N_1641,N_9154);
nor U14832 (N_14832,N_2003,N_4937);
and U14833 (N_14833,N_6627,N_30);
nand U14834 (N_14834,N_2384,N_41);
xor U14835 (N_14835,N_2086,N_4167);
nand U14836 (N_14836,N_7724,N_4206);
xor U14837 (N_14837,N_7508,N_5731);
or U14838 (N_14838,N_1868,N_31);
nor U14839 (N_14839,N_4918,N_8474);
and U14840 (N_14840,N_1156,N_4414);
nand U14841 (N_14841,N_5582,N_2258);
nand U14842 (N_14842,N_2441,N_7146);
xor U14843 (N_14843,N_7313,N_1321);
or U14844 (N_14844,N_9098,N_432);
or U14845 (N_14845,N_6021,N_4983);
xnor U14846 (N_14846,N_7106,N_3408);
nor U14847 (N_14847,N_1971,N_7565);
nand U14848 (N_14848,N_4310,N_4507);
and U14849 (N_14849,N_1225,N_5306);
nand U14850 (N_14850,N_3035,N_8661);
nor U14851 (N_14851,N_8409,N_7814);
nand U14852 (N_14852,N_6129,N_7465);
xnor U14853 (N_14853,N_973,N_464);
and U14854 (N_14854,N_5228,N_1722);
nand U14855 (N_14855,N_6970,N_5866);
nand U14856 (N_14856,N_2446,N_1904);
nand U14857 (N_14857,N_4757,N_1535);
and U14858 (N_14858,N_4393,N_8008);
or U14859 (N_14859,N_101,N_1435);
nor U14860 (N_14860,N_7049,N_8258);
or U14861 (N_14861,N_3172,N_4161);
nor U14862 (N_14862,N_6957,N_3690);
nand U14863 (N_14863,N_6940,N_3154);
nand U14864 (N_14864,N_2422,N_3410);
nand U14865 (N_14865,N_132,N_4277);
and U14866 (N_14866,N_5911,N_2669);
or U14867 (N_14867,N_933,N_262);
or U14868 (N_14868,N_9321,N_7332);
and U14869 (N_14869,N_9991,N_9648);
xor U14870 (N_14870,N_3683,N_7617);
nor U14871 (N_14871,N_2560,N_1157);
nor U14872 (N_14872,N_5051,N_6639);
nand U14873 (N_14873,N_9725,N_2997);
or U14874 (N_14874,N_6879,N_1461);
xnor U14875 (N_14875,N_8457,N_7162);
xor U14876 (N_14876,N_5143,N_4099);
and U14877 (N_14877,N_1827,N_5060);
nand U14878 (N_14878,N_9052,N_436);
or U14879 (N_14879,N_4512,N_7478);
or U14880 (N_14880,N_3807,N_8957);
xnor U14881 (N_14881,N_9147,N_6978);
nor U14882 (N_14882,N_2719,N_6745);
nor U14883 (N_14883,N_622,N_2184);
or U14884 (N_14884,N_1494,N_6568);
or U14885 (N_14885,N_5096,N_1131);
and U14886 (N_14886,N_4968,N_4583);
nor U14887 (N_14887,N_2083,N_8558);
and U14888 (N_14888,N_6777,N_6601);
and U14889 (N_14889,N_8376,N_7633);
and U14890 (N_14890,N_7301,N_5921);
and U14891 (N_14891,N_4974,N_7673);
or U14892 (N_14892,N_6369,N_3584);
nor U14893 (N_14893,N_2565,N_3352);
nor U14894 (N_14894,N_5737,N_3621);
xor U14895 (N_14895,N_6985,N_6067);
or U14896 (N_14896,N_6097,N_5768);
nor U14897 (N_14897,N_8450,N_5477);
nand U14898 (N_14898,N_8025,N_3434);
nor U14899 (N_14899,N_100,N_4410);
nor U14900 (N_14900,N_5607,N_4910);
xnor U14901 (N_14901,N_9139,N_9833);
or U14902 (N_14902,N_8894,N_3353);
xor U14903 (N_14903,N_4519,N_4480);
nand U14904 (N_14904,N_3662,N_3562);
and U14905 (N_14905,N_3887,N_6033);
nand U14906 (N_14906,N_5162,N_7823);
and U14907 (N_14907,N_5205,N_6301);
xor U14908 (N_14908,N_843,N_710);
and U14909 (N_14909,N_5906,N_5940);
nor U14910 (N_14910,N_5245,N_3032);
or U14911 (N_14911,N_7284,N_6729);
nand U14912 (N_14912,N_2787,N_158);
nor U14913 (N_14913,N_5033,N_3543);
xnor U14914 (N_14914,N_9194,N_6833);
nand U14915 (N_14915,N_6947,N_9920);
or U14916 (N_14916,N_3928,N_5179);
nand U14917 (N_14917,N_706,N_6642);
or U14918 (N_14918,N_1514,N_3446);
nor U14919 (N_14919,N_6907,N_7321);
xor U14920 (N_14920,N_9563,N_689);
nor U14921 (N_14921,N_7265,N_1110);
nor U14922 (N_14922,N_2356,N_3018);
or U14923 (N_14923,N_5378,N_6357);
or U14924 (N_14924,N_6400,N_5116);
and U14925 (N_14925,N_9134,N_4649);
nor U14926 (N_14926,N_293,N_3325);
nand U14927 (N_14927,N_6442,N_9589);
nor U14928 (N_14928,N_831,N_7517);
nand U14929 (N_14929,N_3570,N_3767);
and U14930 (N_14930,N_2467,N_3577);
nor U14931 (N_14931,N_6599,N_5523);
nor U14932 (N_14932,N_3842,N_1545);
nand U14933 (N_14933,N_6676,N_348);
xor U14934 (N_14934,N_291,N_2468);
and U14935 (N_14935,N_2311,N_6276);
or U14936 (N_14936,N_3415,N_5398);
xnor U14937 (N_14937,N_2145,N_3094);
xor U14938 (N_14938,N_5412,N_9712);
nor U14939 (N_14939,N_3859,N_85);
nor U14940 (N_14940,N_4802,N_6199);
and U14941 (N_14941,N_4059,N_3946);
and U14942 (N_14942,N_5856,N_3076);
nor U14943 (N_14943,N_350,N_4522);
or U14944 (N_14944,N_61,N_1471);
nor U14945 (N_14945,N_6151,N_6358);
nand U14946 (N_14946,N_3349,N_4516);
and U14947 (N_14947,N_8751,N_7468);
nand U14948 (N_14948,N_2761,N_4804);
xnor U14949 (N_14949,N_9976,N_4285);
and U14950 (N_14950,N_3919,N_8772);
xnor U14951 (N_14951,N_7126,N_1185);
nand U14952 (N_14952,N_4712,N_7806);
or U14953 (N_14953,N_8462,N_7223);
or U14954 (N_14954,N_485,N_862);
nor U14955 (N_14955,N_6816,N_523);
or U14956 (N_14956,N_1906,N_8698);
xor U14957 (N_14957,N_3260,N_6240);
nand U14958 (N_14958,N_7659,N_3195);
nor U14959 (N_14959,N_2677,N_9066);
xnor U14960 (N_14960,N_5930,N_8602);
or U14961 (N_14961,N_9763,N_712);
nand U14962 (N_14962,N_707,N_5250);
or U14963 (N_14963,N_1093,N_6551);
nand U14964 (N_14964,N_2299,N_1483);
or U14965 (N_14965,N_3583,N_4765);
nor U14966 (N_14966,N_819,N_9183);
or U14967 (N_14967,N_5823,N_2689);
or U14968 (N_14968,N_9981,N_4739);
nor U14969 (N_14969,N_6863,N_2709);
or U14970 (N_14970,N_7578,N_1584);
nor U14971 (N_14971,N_2881,N_8269);
nand U14972 (N_14972,N_1529,N_2066);
or U14973 (N_14973,N_8398,N_4157);
nand U14974 (N_14974,N_944,N_3462);
or U14975 (N_14975,N_3458,N_3263);
or U14976 (N_14976,N_8941,N_9468);
nand U14977 (N_14977,N_5780,N_4282);
xnor U14978 (N_14978,N_1031,N_8647);
nand U14979 (N_14979,N_5069,N_4742);
nor U14980 (N_14980,N_7207,N_8264);
nand U14981 (N_14981,N_1308,N_893);
xor U14982 (N_14982,N_5021,N_2408);
and U14983 (N_14983,N_4676,N_4069);
nor U14984 (N_14984,N_1477,N_6366);
or U14985 (N_14985,N_7784,N_6047);
and U14986 (N_14986,N_5319,N_3749);
and U14987 (N_14987,N_2926,N_3198);
nand U14988 (N_14988,N_9901,N_9349);
nand U14989 (N_14989,N_4343,N_5036);
nor U14990 (N_14990,N_2765,N_7048);
and U14991 (N_14991,N_6034,N_5463);
nand U14992 (N_14992,N_8203,N_7302);
nor U14993 (N_14993,N_9752,N_7933);
xor U14994 (N_14994,N_2687,N_3827);
xor U14995 (N_14995,N_3064,N_6708);
xor U14996 (N_14996,N_2366,N_7310);
nand U14997 (N_14997,N_9441,N_4008);
and U14998 (N_14998,N_6292,N_5628);
and U14999 (N_14999,N_5094,N_8500);
nand U15000 (N_15000,N_690,N_6441);
nor U15001 (N_15001,N_6744,N_4983);
or U15002 (N_15002,N_1534,N_6095);
or U15003 (N_15003,N_4634,N_4586);
nor U15004 (N_15004,N_5983,N_9295);
nor U15005 (N_15005,N_322,N_3283);
xor U15006 (N_15006,N_9518,N_7806);
nor U15007 (N_15007,N_126,N_1081);
or U15008 (N_15008,N_9232,N_2033);
nor U15009 (N_15009,N_6537,N_6190);
or U15010 (N_15010,N_7705,N_8960);
nor U15011 (N_15011,N_3815,N_6589);
xor U15012 (N_15012,N_2130,N_2926);
or U15013 (N_15013,N_612,N_8685);
nand U15014 (N_15014,N_9217,N_5084);
nand U15015 (N_15015,N_8621,N_1106);
nor U15016 (N_15016,N_8993,N_9855);
or U15017 (N_15017,N_9383,N_9660);
xor U15018 (N_15018,N_5267,N_2308);
or U15019 (N_15019,N_481,N_1454);
xor U15020 (N_15020,N_9874,N_5969);
nand U15021 (N_15021,N_892,N_7538);
nor U15022 (N_15022,N_4992,N_4965);
and U15023 (N_15023,N_8185,N_3729);
or U15024 (N_15024,N_4282,N_83);
nand U15025 (N_15025,N_9721,N_9547);
xor U15026 (N_15026,N_6492,N_9224);
nand U15027 (N_15027,N_8633,N_2476);
or U15028 (N_15028,N_4951,N_5155);
nor U15029 (N_15029,N_3840,N_2270);
and U15030 (N_15030,N_7467,N_8556);
and U15031 (N_15031,N_9935,N_2239);
xnor U15032 (N_15032,N_301,N_2654);
nand U15033 (N_15033,N_8905,N_6384);
or U15034 (N_15034,N_7923,N_7199);
nor U15035 (N_15035,N_6251,N_7905);
or U15036 (N_15036,N_2646,N_840);
nand U15037 (N_15037,N_6739,N_5701);
nor U15038 (N_15038,N_2406,N_5965);
nor U15039 (N_15039,N_5642,N_3119);
nor U15040 (N_15040,N_8156,N_3109);
nand U15041 (N_15041,N_3499,N_830);
nand U15042 (N_15042,N_3727,N_6106);
nor U15043 (N_15043,N_2869,N_1935);
nor U15044 (N_15044,N_1015,N_736);
or U15045 (N_15045,N_3269,N_2318);
nand U15046 (N_15046,N_9474,N_2589);
and U15047 (N_15047,N_3883,N_4033);
xnor U15048 (N_15048,N_7394,N_6021);
and U15049 (N_15049,N_314,N_8489);
nand U15050 (N_15050,N_1145,N_2680);
nor U15051 (N_15051,N_3798,N_2852);
xor U15052 (N_15052,N_5937,N_8448);
or U15053 (N_15053,N_7936,N_1985);
and U15054 (N_15054,N_2947,N_5935);
or U15055 (N_15055,N_8205,N_8453);
or U15056 (N_15056,N_5236,N_3865);
nand U15057 (N_15057,N_836,N_5609);
xnor U15058 (N_15058,N_4091,N_8319);
or U15059 (N_15059,N_3524,N_807);
nor U15060 (N_15060,N_4839,N_2842);
or U15061 (N_15061,N_506,N_9039);
or U15062 (N_15062,N_5473,N_8095);
nor U15063 (N_15063,N_6952,N_1814);
nor U15064 (N_15064,N_5280,N_6781);
nand U15065 (N_15065,N_9471,N_7915);
nor U15066 (N_15066,N_861,N_6102);
nand U15067 (N_15067,N_8606,N_8762);
nand U15068 (N_15068,N_5911,N_8609);
and U15069 (N_15069,N_6485,N_7158);
xor U15070 (N_15070,N_8218,N_6105);
nand U15071 (N_15071,N_8630,N_3339);
xnor U15072 (N_15072,N_9062,N_7666);
nand U15073 (N_15073,N_5692,N_3939);
nand U15074 (N_15074,N_7456,N_3765);
nor U15075 (N_15075,N_9026,N_7630);
xor U15076 (N_15076,N_6559,N_698);
nor U15077 (N_15077,N_1519,N_8258);
nand U15078 (N_15078,N_5549,N_8280);
and U15079 (N_15079,N_3588,N_6096);
nand U15080 (N_15080,N_2604,N_1915);
xor U15081 (N_15081,N_2264,N_2427);
nand U15082 (N_15082,N_1657,N_4234);
nand U15083 (N_15083,N_2488,N_3979);
xor U15084 (N_15084,N_4478,N_7646);
nor U15085 (N_15085,N_9372,N_9255);
or U15086 (N_15086,N_3282,N_9247);
or U15087 (N_15087,N_7062,N_6260);
nand U15088 (N_15088,N_6141,N_8379);
nand U15089 (N_15089,N_4503,N_7776);
or U15090 (N_15090,N_5942,N_3119);
and U15091 (N_15091,N_9328,N_5524);
xor U15092 (N_15092,N_1553,N_2054);
xnor U15093 (N_15093,N_1849,N_6480);
and U15094 (N_15094,N_1150,N_9748);
nor U15095 (N_15095,N_535,N_9023);
xnor U15096 (N_15096,N_9537,N_9497);
nor U15097 (N_15097,N_7064,N_4590);
nor U15098 (N_15098,N_1016,N_6450);
xnor U15099 (N_15099,N_9770,N_1054);
or U15100 (N_15100,N_6570,N_6476);
or U15101 (N_15101,N_1314,N_3301);
nand U15102 (N_15102,N_5154,N_7049);
nand U15103 (N_15103,N_454,N_9581);
nand U15104 (N_15104,N_1291,N_9388);
xnor U15105 (N_15105,N_441,N_5347);
and U15106 (N_15106,N_4948,N_6576);
and U15107 (N_15107,N_5643,N_3949);
nand U15108 (N_15108,N_1188,N_7326);
nor U15109 (N_15109,N_5006,N_5716);
xor U15110 (N_15110,N_5792,N_526);
nand U15111 (N_15111,N_9898,N_5256);
and U15112 (N_15112,N_3905,N_176);
nor U15113 (N_15113,N_8295,N_9191);
nor U15114 (N_15114,N_749,N_4192);
nor U15115 (N_15115,N_464,N_9356);
or U15116 (N_15116,N_6520,N_4158);
and U15117 (N_15117,N_3669,N_4948);
nand U15118 (N_15118,N_7563,N_7581);
nand U15119 (N_15119,N_2430,N_4804);
nand U15120 (N_15120,N_2490,N_559);
and U15121 (N_15121,N_7934,N_146);
or U15122 (N_15122,N_3475,N_5612);
nor U15123 (N_15123,N_7233,N_660);
and U15124 (N_15124,N_6331,N_3102);
nand U15125 (N_15125,N_3101,N_394);
xor U15126 (N_15126,N_4356,N_393);
or U15127 (N_15127,N_4720,N_8735);
or U15128 (N_15128,N_2226,N_7333);
or U15129 (N_15129,N_3742,N_5927);
xor U15130 (N_15130,N_9898,N_2307);
nor U15131 (N_15131,N_4748,N_1822);
xnor U15132 (N_15132,N_7489,N_5512);
nor U15133 (N_15133,N_3451,N_9244);
or U15134 (N_15134,N_3455,N_901);
xnor U15135 (N_15135,N_9806,N_8582);
and U15136 (N_15136,N_4367,N_6067);
nand U15137 (N_15137,N_1826,N_5516);
nor U15138 (N_15138,N_9274,N_1838);
or U15139 (N_15139,N_2991,N_3866);
nor U15140 (N_15140,N_7480,N_6078);
nand U15141 (N_15141,N_7169,N_4475);
and U15142 (N_15142,N_8036,N_2445);
nor U15143 (N_15143,N_2677,N_5584);
xor U15144 (N_15144,N_2453,N_981);
or U15145 (N_15145,N_8989,N_692);
or U15146 (N_15146,N_2585,N_2032);
and U15147 (N_15147,N_7995,N_4049);
and U15148 (N_15148,N_2989,N_8002);
nand U15149 (N_15149,N_6721,N_9097);
and U15150 (N_15150,N_5616,N_4953);
nor U15151 (N_15151,N_2569,N_8329);
nand U15152 (N_15152,N_9414,N_5936);
or U15153 (N_15153,N_3887,N_767);
nand U15154 (N_15154,N_7477,N_6089);
xor U15155 (N_15155,N_1945,N_588);
xor U15156 (N_15156,N_5831,N_6869);
nor U15157 (N_15157,N_8337,N_4477);
nand U15158 (N_15158,N_8670,N_8204);
nand U15159 (N_15159,N_3467,N_9672);
or U15160 (N_15160,N_2521,N_8230);
nor U15161 (N_15161,N_2362,N_2201);
and U15162 (N_15162,N_8321,N_3897);
nor U15163 (N_15163,N_629,N_4322);
or U15164 (N_15164,N_4138,N_2165);
and U15165 (N_15165,N_6566,N_7560);
and U15166 (N_15166,N_8928,N_4957);
nand U15167 (N_15167,N_2563,N_8298);
or U15168 (N_15168,N_1825,N_4963);
and U15169 (N_15169,N_7885,N_7416);
nor U15170 (N_15170,N_9729,N_711);
nor U15171 (N_15171,N_2169,N_6561);
or U15172 (N_15172,N_4455,N_6552);
xor U15173 (N_15173,N_6776,N_6113);
or U15174 (N_15174,N_1022,N_228);
nand U15175 (N_15175,N_9208,N_7140);
xnor U15176 (N_15176,N_1121,N_4418);
or U15177 (N_15177,N_8360,N_2250);
or U15178 (N_15178,N_7628,N_933);
xnor U15179 (N_15179,N_9151,N_6739);
xor U15180 (N_15180,N_247,N_3026);
or U15181 (N_15181,N_8236,N_4615);
nand U15182 (N_15182,N_5032,N_4623);
xor U15183 (N_15183,N_3337,N_807);
nand U15184 (N_15184,N_2101,N_8531);
nand U15185 (N_15185,N_457,N_4137);
xor U15186 (N_15186,N_2032,N_9268);
nor U15187 (N_15187,N_502,N_9209);
or U15188 (N_15188,N_4762,N_5998);
xnor U15189 (N_15189,N_2375,N_3204);
xor U15190 (N_15190,N_6674,N_4095);
xor U15191 (N_15191,N_9816,N_8050);
or U15192 (N_15192,N_7169,N_7088);
nor U15193 (N_15193,N_6549,N_3078);
and U15194 (N_15194,N_8054,N_4820);
or U15195 (N_15195,N_1072,N_1030);
and U15196 (N_15196,N_588,N_8875);
nand U15197 (N_15197,N_1921,N_6556);
and U15198 (N_15198,N_1297,N_2007);
and U15199 (N_15199,N_5043,N_4516);
xnor U15200 (N_15200,N_1285,N_6121);
and U15201 (N_15201,N_8921,N_5440);
nand U15202 (N_15202,N_1953,N_4181);
nand U15203 (N_15203,N_6494,N_1716);
nor U15204 (N_15204,N_7117,N_493);
or U15205 (N_15205,N_4963,N_3157);
nor U15206 (N_15206,N_8761,N_1546);
or U15207 (N_15207,N_2416,N_7621);
xnor U15208 (N_15208,N_265,N_7361);
nand U15209 (N_15209,N_3910,N_6875);
nand U15210 (N_15210,N_6415,N_5774);
xnor U15211 (N_15211,N_403,N_4742);
nor U15212 (N_15212,N_3225,N_1104);
xnor U15213 (N_15213,N_7327,N_4080);
or U15214 (N_15214,N_7946,N_4792);
or U15215 (N_15215,N_6980,N_5124);
or U15216 (N_15216,N_7051,N_9059);
xor U15217 (N_15217,N_5044,N_8210);
xor U15218 (N_15218,N_3299,N_7398);
and U15219 (N_15219,N_7653,N_9956);
xor U15220 (N_15220,N_9013,N_1301);
nor U15221 (N_15221,N_1104,N_2871);
xnor U15222 (N_15222,N_2852,N_153);
and U15223 (N_15223,N_454,N_3995);
or U15224 (N_15224,N_3538,N_129);
or U15225 (N_15225,N_8126,N_6045);
xor U15226 (N_15226,N_2391,N_7333);
xor U15227 (N_15227,N_8311,N_406);
nor U15228 (N_15228,N_5131,N_3999);
and U15229 (N_15229,N_8676,N_2267);
and U15230 (N_15230,N_2881,N_9518);
nand U15231 (N_15231,N_600,N_9574);
nor U15232 (N_15232,N_7287,N_7432);
nand U15233 (N_15233,N_5035,N_5801);
or U15234 (N_15234,N_3414,N_1308);
or U15235 (N_15235,N_667,N_8807);
nand U15236 (N_15236,N_4266,N_8506);
or U15237 (N_15237,N_3166,N_9814);
nor U15238 (N_15238,N_1627,N_2248);
nand U15239 (N_15239,N_9933,N_8653);
nand U15240 (N_15240,N_1290,N_1041);
nand U15241 (N_15241,N_6345,N_6348);
nor U15242 (N_15242,N_6554,N_8994);
or U15243 (N_15243,N_6818,N_5650);
nor U15244 (N_15244,N_5983,N_7240);
xnor U15245 (N_15245,N_8724,N_6012);
xnor U15246 (N_15246,N_4834,N_1641);
or U15247 (N_15247,N_3502,N_1135);
nand U15248 (N_15248,N_537,N_8543);
xor U15249 (N_15249,N_5296,N_6647);
and U15250 (N_15250,N_6791,N_4416);
nand U15251 (N_15251,N_5713,N_4892);
nor U15252 (N_15252,N_5498,N_6953);
and U15253 (N_15253,N_9638,N_5669);
or U15254 (N_15254,N_5167,N_500);
xnor U15255 (N_15255,N_9483,N_1001);
and U15256 (N_15256,N_4314,N_164);
nor U15257 (N_15257,N_6444,N_1700);
nor U15258 (N_15258,N_2676,N_9014);
nand U15259 (N_15259,N_4548,N_5201);
nand U15260 (N_15260,N_6259,N_2347);
nor U15261 (N_15261,N_9978,N_8809);
xor U15262 (N_15262,N_9023,N_1935);
xnor U15263 (N_15263,N_8692,N_2912);
nor U15264 (N_15264,N_4623,N_2040);
or U15265 (N_15265,N_4225,N_510);
and U15266 (N_15266,N_4435,N_2158);
nor U15267 (N_15267,N_4180,N_5347);
nand U15268 (N_15268,N_4445,N_1190);
nor U15269 (N_15269,N_4429,N_312);
nand U15270 (N_15270,N_611,N_5525);
xnor U15271 (N_15271,N_2600,N_4282);
or U15272 (N_15272,N_9922,N_6923);
xnor U15273 (N_15273,N_4230,N_3576);
nor U15274 (N_15274,N_4231,N_5805);
and U15275 (N_15275,N_813,N_8877);
and U15276 (N_15276,N_2679,N_6745);
xor U15277 (N_15277,N_8568,N_548);
nor U15278 (N_15278,N_4500,N_8068);
or U15279 (N_15279,N_5326,N_2595);
xnor U15280 (N_15280,N_335,N_9064);
nor U15281 (N_15281,N_52,N_2325);
xor U15282 (N_15282,N_7664,N_8651);
nor U15283 (N_15283,N_1852,N_9101);
nand U15284 (N_15284,N_1674,N_7470);
nor U15285 (N_15285,N_4334,N_3943);
and U15286 (N_15286,N_4109,N_3833);
nand U15287 (N_15287,N_4322,N_9672);
nand U15288 (N_15288,N_1032,N_1695);
and U15289 (N_15289,N_6046,N_9453);
nor U15290 (N_15290,N_6289,N_4343);
nand U15291 (N_15291,N_9363,N_7863);
or U15292 (N_15292,N_1746,N_5775);
nor U15293 (N_15293,N_9802,N_3751);
and U15294 (N_15294,N_5543,N_6933);
nand U15295 (N_15295,N_1326,N_1968);
nor U15296 (N_15296,N_8823,N_6613);
or U15297 (N_15297,N_5428,N_2021);
nor U15298 (N_15298,N_3548,N_6361);
or U15299 (N_15299,N_5283,N_7001);
xor U15300 (N_15300,N_7235,N_5213);
nor U15301 (N_15301,N_4445,N_8699);
and U15302 (N_15302,N_2554,N_8513);
and U15303 (N_15303,N_5223,N_5538);
nor U15304 (N_15304,N_9978,N_5473);
or U15305 (N_15305,N_8804,N_974);
nor U15306 (N_15306,N_2158,N_3857);
and U15307 (N_15307,N_750,N_5527);
nand U15308 (N_15308,N_3066,N_2527);
nand U15309 (N_15309,N_8857,N_1182);
or U15310 (N_15310,N_4730,N_2450);
nor U15311 (N_15311,N_5523,N_5192);
or U15312 (N_15312,N_5385,N_1843);
or U15313 (N_15313,N_19,N_3038);
nand U15314 (N_15314,N_3340,N_1779);
and U15315 (N_15315,N_6863,N_447);
and U15316 (N_15316,N_7008,N_2414);
xor U15317 (N_15317,N_9273,N_1383);
nor U15318 (N_15318,N_843,N_2400);
nor U15319 (N_15319,N_6985,N_1994);
nor U15320 (N_15320,N_7740,N_3855);
or U15321 (N_15321,N_4820,N_7735);
xnor U15322 (N_15322,N_2818,N_8031);
nor U15323 (N_15323,N_5785,N_5988);
or U15324 (N_15324,N_8850,N_8646);
or U15325 (N_15325,N_6892,N_1615);
or U15326 (N_15326,N_9612,N_1635);
and U15327 (N_15327,N_7139,N_3523);
xnor U15328 (N_15328,N_9657,N_6775);
nand U15329 (N_15329,N_8087,N_5429);
nor U15330 (N_15330,N_2136,N_8335);
nand U15331 (N_15331,N_7587,N_5569);
or U15332 (N_15332,N_8708,N_7361);
or U15333 (N_15333,N_5833,N_3010);
nor U15334 (N_15334,N_1215,N_8566);
or U15335 (N_15335,N_5605,N_4223);
and U15336 (N_15336,N_8593,N_1524);
xor U15337 (N_15337,N_4272,N_7927);
nor U15338 (N_15338,N_1028,N_5590);
and U15339 (N_15339,N_2041,N_596);
xor U15340 (N_15340,N_9455,N_7477);
nand U15341 (N_15341,N_4911,N_2993);
nand U15342 (N_15342,N_3946,N_2027);
nand U15343 (N_15343,N_5608,N_6197);
or U15344 (N_15344,N_2860,N_6214);
or U15345 (N_15345,N_3503,N_9805);
or U15346 (N_15346,N_532,N_2339);
nor U15347 (N_15347,N_2328,N_6891);
nor U15348 (N_15348,N_6504,N_7498);
and U15349 (N_15349,N_8156,N_7858);
nor U15350 (N_15350,N_5983,N_7663);
nand U15351 (N_15351,N_5990,N_9233);
nand U15352 (N_15352,N_7122,N_6719);
and U15353 (N_15353,N_8987,N_9374);
and U15354 (N_15354,N_22,N_4841);
or U15355 (N_15355,N_8286,N_8016);
nor U15356 (N_15356,N_8724,N_562);
nor U15357 (N_15357,N_9112,N_5497);
and U15358 (N_15358,N_8534,N_5519);
and U15359 (N_15359,N_8583,N_7058);
nand U15360 (N_15360,N_6976,N_5120);
and U15361 (N_15361,N_846,N_9742);
or U15362 (N_15362,N_1145,N_9272);
and U15363 (N_15363,N_5259,N_3051);
nand U15364 (N_15364,N_7191,N_2460);
nor U15365 (N_15365,N_7718,N_5518);
and U15366 (N_15366,N_6289,N_6864);
and U15367 (N_15367,N_6873,N_6595);
or U15368 (N_15368,N_4544,N_3708);
nor U15369 (N_15369,N_3576,N_1667);
nor U15370 (N_15370,N_7566,N_8363);
nand U15371 (N_15371,N_9117,N_9292);
xnor U15372 (N_15372,N_7070,N_2888);
nor U15373 (N_15373,N_1752,N_155);
or U15374 (N_15374,N_2071,N_9753);
or U15375 (N_15375,N_3163,N_3845);
or U15376 (N_15376,N_4166,N_8676);
or U15377 (N_15377,N_3852,N_3107);
nand U15378 (N_15378,N_9145,N_8343);
or U15379 (N_15379,N_9954,N_8474);
or U15380 (N_15380,N_6684,N_1101);
nand U15381 (N_15381,N_3214,N_48);
nor U15382 (N_15382,N_8124,N_6880);
or U15383 (N_15383,N_647,N_6934);
nand U15384 (N_15384,N_8981,N_9312);
or U15385 (N_15385,N_236,N_6974);
or U15386 (N_15386,N_5669,N_1973);
xnor U15387 (N_15387,N_5744,N_6408);
xor U15388 (N_15388,N_1040,N_7430);
nand U15389 (N_15389,N_6789,N_3280);
and U15390 (N_15390,N_6008,N_3608);
nor U15391 (N_15391,N_8998,N_7699);
or U15392 (N_15392,N_980,N_7624);
xor U15393 (N_15393,N_8646,N_248);
xor U15394 (N_15394,N_2022,N_1555);
xnor U15395 (N_15395,N_6745,N_6791);
nor U15396 (N_15396,N_3625,N_1600);
and U15397 (N_15397,N_6549,N_879);
nand U15398 (N_15398,N_8342,N_9621);
xnor U15399 (N_15399,N_2564,N_9089);
nand U15400 (N_15400,N_1028,N_3336);
xor U15401 (N_15401,N_3081,N_3);
nor U15402 (N_15402,N_6473,N_6244);
or U15403 (N_15403,N_6275,N_756);
and U15404 (N_15404,N_9679,N_872);
or U15405 (N_15405,N_5520,N_1417);
xor U15406 (N_15406,N_3326,N_5902);
nor U15407 (N_15407,N_8841,N_5054);
nor U15408 (N_15408,N_8177,N_7424);
nor U15409 (N_15409,N_6473,N_278);
nor U15410 (N_15410,N_88,N_72);
nor U15411 (N_15411,N_4976,N_3895);
nor U15412 (N_15412,N_5951,N_6186);
xor U15413 (N_15413,N_3373,N_7579);
nand U15414 (N_15414,N_3169,N_2541);
and U15415 (N_15415,N_3928,N_2344);
nor U15416 (N_15416,N_6123,N_5007);
or U15417 (N_15417,N_9766,N_7789);
nand U15418 (N_15418,N_4365,N_4261);
and U15419 (N_15419,N_8989,N_3606);
nor U15420 (N_15420,N_5261,N_4578);
xnor U15421 (N_15421,N_8200,N_6560);
or U15422 (N_15422,N_2031,N_6626);
and U15423 (N_15423,N_8275,N_7252);
or U15424 (N_15424,N_5880,N_2170);
nor U15425 (N_15425,N_315,N_8462);
or U15426 (N_15426,N_7142,N_815);
nor U15427 (N_15427,N_3015,N_5468);
nand U15428 (N_15428,N_1269,N_1319);
and U15429 (N_15429,N_4796,N_94);
and U15430 (N_15430,N_1534,N_2971);
nand U15431 (N_15431,N_2379,N_9911);
nor U15432 (N_15432,N_3635,N_2641);
xnor U15433 (N_15433,N_5863,N_7971);
xor U15434 (N_15434,N_2068,N_1863);
xor U15435 (N_15435,N_3837,N_4724);
or U15436 (N_15436,N_8109,N_6573);
nand U15437 (N_15437,N_3030,N_510);
nor U15438 (N_15438,N_1524,N_3064);
nand U15439 (N_15439,N_685,N_5609);
nor U15440 (N_15440,N_2733,N_1511);
xnor U15441 (N_15441,N_8498,N_2804);
and U15442 (N_15442,N_7326,N_3404);
or U15443 (N_15443,N_3186,N_5544);
or U15444 (N_15444,N_1328,N_8591);
and U15445 (N_15445,N_2955,N_301);
nand U15446 (N_15446,N_1722,N_3321);
xor U15447 (N_15447,N_830,N_4303);
xnor U15448 (N_15448,N_136,N_1798);
xnor U15449 (N_15449,N_1983,N_4573);
xnor U15450 (N_15450,N_9279,N_6555);
or U15451 (N_15451,N_5584,N_1870);
nor U15452 (N_15452,N_4033,N_8511);
or U15453 (N_15453,N_5955,N_3950);
nor U15454 (N_15454,N_747,N_3685);
or U15455 (N_15455,N_3956,N_4307);
or U15456 (N_15456,N_9375,N_5082);
nand U15457 (N_15457,N_512,N_6873);
nor U15458 (N_15458,N_1696,N_1230);
and U15459 (N_15459,N_5990,N_5556);
and U15460 (N_15460,N_8122,N_6686);
and U15461 (N_15461,N_7064,N_7114);
or U15462 (N_15462,N_9666,N_3808);
or U15463 (N_15463,N_681,N_2540);
nor U15464 (N_15464,N_6888,N_8163);
xor U15465 (N_15465,N_1563,N_206);
nor U15466 (N_15466,N_8763,N_1786);
nand U15467 (N_15467,N_2130,N_6389);
nand U15468 (N_15468,N_5133,N_8378);
xor U15469 (N_15469,N_5727,N_8461);
nor U15470 (N_15470,N_4780,N_4456);
nand U15471 (N_15471,N_6331,N_370);
nor U15472 (N_15472,N_9809,N_5121);
and U15473 (N_15473,N_9569,N_4423);
nor U15474 (N_15474,N_1581,N_1135);
or U15475 (N_15475,N_2492,N_6051);
xor U15476 (N_15476,N_8167,N_5322);
or U15477 (N_15477,N_4381,N_9903);
and U15478 (N_15478,N_5327,N_7060);
xnor U15479 (N_15479,N_8392,N_4672);
and U15480 (N_15480,N_8845,N_448);
nor U15481 (N_15481,N_938,N_8208);
and U15482 (N_15482,N_5394,N_5845);
nor U15483 (N_15483,N_1751,N_7995);
xor U15484 (N_15484,N_1899,N_6585);
or U15485 (N_15485,N_8220,N_4944);
nand U15486 (N_15486,N_3053,N_1126);
and U15487 (N_15487,N_298,N_5934);
xnor U15488 (N_15488,N_3733,N_4604);
and U15489 (N_15489,N_5687,N_286);
or U15490 (N_15490,N_7220,N_6067);
xnor U15491 (N_15491,N_8941,N_2217);
and U15492 (N_15492,N_1655,N_7559);
xor U15493 (N_15493,N_71,N_7299);
or U15494 (N_15494,N_7626,N_1529);
xor U15495 (N_15495,N_3281,N_7286);
nor U15496 (N_15496,N_2963,N_9268);
nand U15497 (N_15497,N_1685,N_4402);
nand U15498 (N_15498,N_1838,N_4640);
nor U15499 (N_15499,N_3551,N_967);
nor U15500 (N_15500,N_8932,N_9627);
and U15501 (N_15501,N_9403,N_1693);
nor U15502 (N_15502,N_9123,N_4800);
or U15503 (N_15503,N_9041,N_902);
nand U15504 (N_15504,N_2423,N_2574);
and U15505 (N_15505,N_3120,N_3755);
nand U15506 (N_15506,N_6310,N_1939);
nand U15507 (N_15507,N_2329,N_6605);
xnor U15508 (N_15508,N_485,N_9233);
nor U15509 (N_15509,N_5784,N_3132);
nor U15510 (N_15510,N_3792,N_2696);
nand U15511 (N_15511,N_3443,N_700);
nor U15512 (N_15512,N_5868,N_6883);
nand U15513 (N_15513,N_5708,N_1173);
nor U15514 (N_15514,N_1740,N_2077);
and U15515 (N_15515,N_8461,N_1679);
xnor U15516 (N_15516,N_1730,N_606);
xnor U15517 (N_15517,N_6168,N_8560);
xor U15518 (N_15518,N_9979,N_8768);
and U15519 (N_15519,N_124,N_93);
xnor U15520 (N_15520,N_6435,N_6580);
and U15521 (N_15521,N_4685,N_3534);
xor U15522 (N_15522,N_4586,N_5672);
nor U15523 (N_15523,N_7488,N_6204);
and U15524 (N_15524,N_881,N_6309);
or U15525 (N_15525,N_5919,N_6333);
nor U15526 (N_15526,N_2239,N_4179);
xor U15527 (N_15527,N_5703,N_932);
or U15528 (N_15528,N_7700,N_7747);
xnor U15529 (N_15529,N_9259,N_7602);
nand U15530 (N_15530,N_3514,N_459);
nand U15531 (N_15531,N_7965,N_2613);
nand U15532 (N_15532,N_4287,N_4229);
xor U15533 (N_15533,N_8651,N_6744);
nand U15534 (N_15534,N_8537,N_8203);
nor U15535 (N_15535,N_0,N_1095);
nor U15536 (N_15536,N_9141,N_3264);
or U15537 (N_15537,N_2983,N_2567);
nand U15538 (N_15538,N_2987,N_5579);
nand U15539 (N_15539,N_3382,N_6985);
nor U15540 (N_15540,N_3464,N_6054);
xor U15541 (N_15541,N_2555,N_2898);
or U15542 (N_15542,N_8371,N_6995);
nor U15543 (N_15543,N_1401,N_1060);
xor U15544 (N_15544,N_839,N_824);
nor U15545 (N_15545,N_7420,N_1199);
nand U15546 (N_15546,N_4443,N_8134);
nand U15547 (N_15547,N_6601,N_162);
nand U15548 (N_15548,N_7530,N_2795);
nand U15549 (N_15549,N_4540,N_8406);
xor U15550 (N_15550,N_7734,N_5022);
xor U15551 (N_15551,N_2426,N_4121);
xor U15552 (N_15552,N_5177,N_3216);
nor U15553 (N_15553,N_7122,N_9502);
nor U15554 (N_15554,N_3162,N_1036);
nand U15555 (N_15555,N_7205,N_3158);
or U15556 (N_15556,N_7935,N_4042);
or U15557 (N_15557,N_6741,N_648);
and U15558 (N_15558,N_5251,N_2388);
nor U15559 (N_15559,N_5682,N_4494);
nand U15560 (N_15560,N_7521,N_7908);
nand U15561 (N_15561,N_9247,N_3577);
or U15562 (N_15562,N_719,N_975);
or U15563 (N_15563,N_2464,N_7248);
nand U15564 (N_15564,N_8513,N_1724);
and U15565 (N_15565,N_5033,N_4979);
xor U15566 (N_15566,N_9514,N_6227);
nand U15567 (N_15567,N_786,N_7927);
and U15568 (N_15568,N_8505,N_2137);
and U15569 (N_15569,N_5212,N_216);
nand U15570 (N_15570,N_4099,N_3084);
nor U15571 (N_15571,N_7332,N_4885);
nor U15572 (N_15572,N_2261,N_2974);
or U15573 (N_15573,N_62,N_9320);
nand U15574 (N_15574,N_6830,N_1720);
nand U15575 (N_15575,N_7366,N_8441);
and U15576 (N_15576,N_5137,N_2298);
nand U15577 (N_15577,N_991,N_3070);
nand U15578 (N_15578,N_427,N_3139);
and U15579 (N_15579,N_6736,N_87);
or U15580 (N_15580,N_6530,N_2688);
nand U15581 (N_15581,N_5863,N_6931);
or U15582 (N_15582,N_9781,N_5490);
nor U15583 (N_15583,N_5131,N_4924);
or U15584 (N_15584,N_462,N_1771);
and U15585 (N_15585,N_191,N_3927);
nor U15586 (N_15586,N_5503,N_9486);
nand U15587 (N_15587,N_3479,N_2284);
nor U15588 (N_15588,N_9780,N_4916);
and U15589 (N_15589,N_2551,N_1247);
and U15590 (N_15590,N_5178,N_7225);
xnor U15591 (N_15591,N_9603,N_4036);
and U15592 (N_15592,N_4691,N_9795);
nand U15593 (N_15593,N_3824,N_804);
xnor U15594 (N_15594,N_8114,N_4174);
nand U15595 (N_15595,N_3472,N_5571);
or U15596 (N_15596,N_8290,N_3201);
xnor U15597 (N_15597,N_2956,N_18);
nor U15598 (N_15598,N_1080,N_3199);
nand U15599 (N_15599,N_7674,N_5947);
nor U15600 (N_15600,N_4791,N_9261);
or U15601 (N_15601,N_9538,N_9971);
or U15602 (N_15602,N_4804,N_5102);
and U15603 (N_15603,N_2256,N_7486);
and U15604 (N_15604,N_8523,N_1750);
or U15605 (N_15605,N_3276,N_5131);
and U15606 (N_15606,N_8668,N_6833);
nand U15607 (N_15607,N_5508,N_6436);
nand U15608 (N_15608,N_7104,N_2403);
nor U15609 (N_15609,N_8470,N_9458);
nor U15610 (N_15610,N_278,N_8806);
or U15611 (N_15611,N_684,N_7378);
or U15612 (N_15612,N_6800,N_6950);
nor U15613 (N_15613,N_9966,N_5975);
nand U15614 (N_15614,N_5662,N_7708);
or U15615 (N_15615,N_5620,N_1543);
or U15616 (N_15616,N_1366,N_5932);
xnor U15617 (N_15617,N_7088,N_9375);
and U15618 (N_15618,N_8425,N_2490);
xor U15619 (N_15619,N_1314,N_4198);
nand U15620 (N_15620,N_2564,N_7046);
or U15621 (N_15621,N_7209,N_588);
and U15622 (N_15622,N_6271,N_1003);
xor U15623 (N_15623,N_1773,N_662);
nand U15624 (N_15624,N_7929,N_1457);
nor U15625 (N_15625,N_5320,N_4078);
xnor U15626 (N_15626,N_2250,N_8609);
nor U15627 (N_15627,N_4961,N_7889);
or U15628 (N_15628,N_6857,N_7828);
nor U15629 (N_15629,N_268,N_7524);
or U15630 (N_15630,N_6615,N_2520);
nand U15631 (N_15631,N_7116,N_6146);
nor U15632 (N_15632,N_5331,N_5008);
nor U15633 (N_15633,N_6171,N_8525);
xnor U15634 (N_15634,N_9700,N_7567);
nand U15635 (N_15635,N_7085,N_5842);
nor U15636 (N_15636,N_5858,N_4209);
nand U15637 (N_15637,N_1701,N_8518);
and U15638 (N_15638,N_7194,N_9922);
xnor U15639 (N_15639,N_1368,N_5703);
nand U15640 (N_15640,N_8639,N_8923);
or U15641 (N_15641,N_871,N_3953);
nand U15642 (N_15642,N_8718,N_6601);
nor U15643 (N_15643,N_7547,N_783);
or U15644 (N_15644,N_4334,N_628);
and U15645 (N_15645,N_2790,N_7237);
and U15646 (N_15646,N_740,N_6184);
xor U15647 (N_15647,N_6839,N_3648);
xnor U15648 (N_15648,N_4712,N_1784);
nand U15649 (N_15649,N_1588,N_5667);
nand U15650 (N_15650,N_6517,N_837);
or U15651 (N_15651,N_652,N_4021);
nand U15652 (N_15652,N_3314,N_6249);
xnor U15653 (N_15653,N_2114,N_8118);
or U15654 (N_15654,N_2465,N_9669);
xor U15655 (N_15655,N_2396,N_2398);
nor U15656 (N_15656,N_5121,N_7876);
and U15657 (N_15657,N_5394,N_1492);
xor U15658 (N_15658,N_728,N_3100);
xor U15659 (N_15659,N_7486,N_5556);
and U15660 (N_15660,N_8675,N_775);
nor U15661 (N_15661,N_7056,N_6785);
xnor U15662 (N_15662,N_8125,N_610);
xnor U15663 (N_15663,N_7275,N_7847);
xnor U15664 (N_15664,N_3022,N_411);
xor U15665 (N_15665,N_2066,N_9915);
nor U15666 (N_15666,N_9374,N_8231);
nor U15667 (N_15667,N_7505,N_6530);
or U15668 (N_15668,N_376,N_5717);
nand U15669 (N_15669,N_5638,N_7285);
or U15670 (N_15670,N_5324,N_9004);
and U15671 (N_15671,N_1354,N_5728);
nor U15672 (N_15672,N_6464,N_4161);
xnor U15673 (N_15673,N_2601,N_981);
or U15674 (N_15674,N_6458,N_6910);
xor U15675 (N_15675,N_196,N_3988);
xor U15676 (N_15676,N_2166,N_5437);
nor U15677 (N_15677,N_6872,N_3186);
nor U15678 (N_15678,N_9469,N_2546);
or U15679 (N_15679,N_7641,N_7681);
or U15680 (N_15680,N_5958,N_660);
and U15681 (N_15681,N_5031,N_6762);
and U15682 (N_15682,N_5682,N_32);
xor U15683 (N_15683,N_1735,N_1463);
nand U15684 (N_15684,N_9120,N_2673);
xor U15685 (N_15685,N_6108,N_625);
nand U15686 (N_15686,N_1614,N_6015);
xor U15687 (N_15687,N_140,N_6666);
xor U15688 (N_15688,N_5422,N_7189);
nor U15689 (N_15689,N_9807,N_3115);
nand U15690 (N_15690,N_9296,N_6022);
and U15691 (N_15691,N_4818,N_8530);
and U15692 (N_15692,N_5846,N_5613);
or U15693 (N_15693,N_7763,N_1494);
xnor U15694 (N_15694,N_4721,N_7522);
nand U15695 (N_15695,N_9727,N_9173);
xnor U15696 (N_15696,N_4065,N_1562);
nand U15697 (N_15697,N_6893,N_1701);
and U15698 (N_15698,N_6173,N_4621);
nor U15699 (N_15699,N_9693,N_8948);
nor U15700 (N_15700,N_73,N_5363);
and U15701 (N_15701,N_6854,N_9628);
xnor U15702 (N_15702,N_5404,N_493);
and U15703 (N_15703,N_2735,N_9578);
or U15704 (N_15704,N_2356,N_9656);
xor U15705 (N_15705,N_3735,N_100);
or U15706 (N_15706,N_5956,N_8134);
and U15707 (N_15707,N_4900,N_5201);
and U15708 (N_15708,N_4214,N_3980);
nor U15709 (N_15709,N_5043,N_9234);
and U15710 (N_15710,N_5182,N_8817);
nor U15711 (N_15711,N_8209,N_5377);
nand U15712 (N_15712,N_5723,N_7394);
nand U15713 (N_15713,N_3298,N_1421);
nor U15714 (N_15714,N_5341,N_4242);
xor U15715 (N_15715,N_1903,N_5921);
nand U15716 (N_15716,N_2526,N_2528);
xnor U15717 (N_15717,N_3760,N_4250);
or U15718 (N_15718,N_8759,N_2078);
nand U15719 (N_15719,N_4603,N_652);
xor U15720 (N_15720,N_9443,N_8035);
nor U15721 (N_15721,N_679,N_120);
nand U15722 (N_15722,N_6231,N_287);
or U15723 (N_15723,N_4397,N_7057);
or U15724 (N_15724,N_5843,N_3504);
xnor U15725 (N_15725,N_1282,N_517);
or U15726 (N_15726,N_8105,N_8572);
nand U15727 (N_15727,N_7392,N_6173);
and U15728 (N_15728,N_4490,N_8483);
nand U15729 (N_15729,N_8184,N_9081);
and U15730 (N_15730,N_7883,N_3598);
and U15731 (N_15731,N_5074,N_2600);
xor U15732 (N_15732,N_1141,N_960);
xnor U15733 (N_15733,N_8430,N_8156);
and U15734 (N_15734,N_9239,N_8383);
xor U15735 (N_15735,N_8318,N_1130);
and U15736 (N_15736,N_7415,N_6267);
nand U15737 (N_15737,N_5882,N_5128);
nor U15738 (N_15738,N_5567,N_9784);
and U15739 (N_15739,N_3566,N_7378);
nor U15740 (N_15740,N_9424,N_935);
or U15741 (N_15741,N_3020,N_8114);
and U15742 (N_15742,N_4244,N_1978);
and U15743 (N_15743,N_3541,N_8456);
xnor U15744 (N_15744,N_6559,N_9802);
or U15745 (N_15745,N_8626,N_1099);
nor U15746 (N_15746,N_1049,N_7792);
and U15747 (N_15747,N_6226,N_9551);
xnor U15748 (N_15748,N_7593,N_7889);
nand U15749 (N_15749,N_421,N_2890);
nand U15750 (N_15750,N_2496,N_1430);
nand U15751 (N_15751,N_5449,N_3405);
nand U15752 (N_15752,N_3631,N_7236);
nor U15753 (N_15753,N_5139,N_2377);
nand U15754 (N_15754,N_5006,N_3768);
nor U15755 (N_15755,N_8811,N_83);
nand U15756 (N_15756,N_6268,N_8836);
or U15757 (N_15757,N_4948,N_5130);
or U15758 (N_15758,N_2011,N_1233);
xnor U15759 (N_15759,N_6451,N_7782);
nor U15760 (N_15760,N_1410,N_8178);
nor U15761 (N_15761,N_5640,N_875);
and U15762 (N_15762,N_1088,N_5667);
and U15763 (N_15763,N_4526,N_1834);
or U15764 (N_15764,N_7574,N_9545);
nand U15765 (N_15765,N_8567,N_7067);
nand U15766 (N_15766,N_4921,N_9246);
nand U15767 (N_15767,N_2462,N_3277);
nor U15768 (N_15768,N_1122,N_703);
nor U15769 (N_15769,N_3218,N_6755);
nor U15770 (N_15770,N_1577,N_7559);
and U15771 (N_15771,N_9698,N_6077);
and U15772 (N_15772,N_1373,N_1958);
xor U15773 (N_15773,N_9964,N_306);
or U15774 (N_15774,N_8131,N_5651);
nor U15775 (N_15775,N_7531,N_678);
nand U15776 (N_15776,N_5430,N_5287);
or U15777 (N_15777,N_4878,N_1598);
or U15778 (N_15778,N_8825,N_4772);
nor U15779 (N_15779,N_9733,N_971);
xnor U15780 (N_15780,N_1852,N_1499);
xnor U15781 (N_15781,N_8371,N_9823);
xor U15782 (N_15782,N_1506,N_7908);
or U15783 (N_15783,N_9190,N_1391);
xnor U15784 (N_15784,N_9449,N_9495);
or U15785 (N_15785,N_1642,N_6088);
nor U15786 (N_15786,N_813,N_2041);
xnor U15787 (N_15787,N_1310,N_4249);
nand U15788 (N_15788,N_9788,N_3220);
and U15789 (N_15789,N_4896,N_8081);
and U15790 (N_15790,N_2857,N_9809);
xor U15791 (N_15791,N_8902,N_2753);
xor U15792 (N_15792,N_7341,N_4135);
or U15793 (N_15793,N_8725,N_5121);
nor U15794 (N_15794,N_5207,N_2557);
and U15795 (N_15795,N_6239,N_1630);
or U15796 (N_15796,N_5216,N_2665);
or U15797 (N_15797,N_3224,N_4582);
xnor U15798 (N_15798,N_930,N_6343);
nor U15799 (N_15799,N_4649,N_5354);
or U15800 (N_15800,N_5182,N_4161);
xnor U15801 (N_15801,N_3024,N_8596);
and U15802 (N_15802,N_8998,N_6569);
and U15803 (N_15803,N_4684,N_1660);
nand U15804 (N_15804,N_160,N_1314);
xor U15805 (N_15805,N_3601,N_4305);
nand U15806 (N_15806,N_8111,N_2962);
nand U15807 (N_15807,N_8197,N_8025);
and U15808 (N_15808,N_6150,N_9585);
and U15809 (N_15809,N_1118,N_8148);
or U15810 (N_15810,N_2894,N_252);
or U15811 (N_15811,N_211,N_9169);
nor U15812 (N_15812,N_7072,N_1574);
nand U15813 (N_15813,N_3913,N_7988);
and U15814 (N_15814,N_1059,N_1980);
nor U15815 (N_15815,N_4656,N_8352);
or U15816 (N_15816,N_9379,N_2618);
nor U15817 (N_15817,N_6406,N_9495);
or U15818 (N_15818,N_5370,N_6299);
xnor U15819 (N_15819,N_6014,N_220);
xnor U15820 (N_15820,N_675,N_26);
nor U15821 (N_15821,N_5170,N_5363);
nand U15822 (N_15822,N_9445,N_2558);
and U15823 (N_15823,N_5175,N_6575);
nor U15824 (N_15824,N_3564,N_792);
xnor U15825 (N_15825,N_1128,N_2344);
and U15826 (N_15826,N_7298,N_527);
nand U15827 (N_15827,N_2029,N_5514);
nor U15828 (N_15828,N_9091,N_9136);
nand U15829 (N_15829,N_9166,N_5652);
nand U15830 (N_15830,N_9739,N_3775);
or U15831 (N_15831,N_1554,N_4960);
xor U15832 (N_15832,N_6260,N_960);
and U15833 (N_15833,N_8561,N_7553);
xnor U15834 (N_15834,N_2545,N_9155);
nor U15835 (N_15835,N_5587,N_3453);
or U15836 (N_15836,N_7220,N_1434);
xnor U15837 (N_15837,N_4741,N_2129);
and U15838 (N_15838,N_4327,N_455);
xnor U15839 (N_15839,N_6770,N_1628);
and U15840 (N_15840,N_9143,N_5497);
nand U15841 (N_15841,N_117,N_7397);
nor U15842 (N_15842,N_9316,N_4201);
nor U15843 (N_15843,N_3622,N_4669);
nand U15844 (N_15844,N_4397,N_4149);
nor U15845 (N_15845,N_5570,N_438);
xnor U15846 (N_15846,N_7976,N_5731);
or U15847 (N_15847,N_6342,N_7210);
nand U15848 (N_15848,N_3258,N_7153);
and U15849 (N_15849,N_6678,N_6664);
or U15850 (N_15850,N_7848,N_1037);
or U15851 (N_15851,N_2467,N_2551);
and U15852 (N_15852,N_6475,N_3722);
nand U15853 (N_15853,N_5406,N_7366);
xor U15854 (N_15854,N_8904,N_7187);
xor U15855 (N_15855,N_9788,N_4092);
and U15856 (N_15856,N_8336,N_3641);
nand U15857 (N_15857,N_2446,N_4790);
or U15858 (N_15858,N_8647,N_5814);
nand U15859 (N_15859,N_517,N_8770);
and U15860 (N_15860,N_6797,N_4585);
and U15861 (N_15861,N_9059,N_4740);
or U15862 (N_15862,N_8385,N_1314);
nor U15863 (N_15863,N_2492,N_1113);
and U15864 (N_15864,N_8022,N_6750);
and U15865 (N_15865,N_5835,N_8366);
and U15866 (N_15866,N_5874,N_1189);
and U15867 (N_15867,N_5073,N_1534);
and U15868 (N_15868,N_5492,N_9025);
nand U15869 (N_15869,N_6777,N_8531);
and U15870 (N_15870,N_1978,N_3582);
nor U15871 (N_15871,N_7617,N_2670);
xnor U15872 (N_15872,N_570,N_6173);
or U15873 (N_15873,N_736,N_6163);
and U15874 (N_15874,N_5090,N_2619);
xor U15875 (N_15875,N_4976,N_9140);
and U15876 (N_15876,N_1275,N_4929);
nand U15877 (N_15877,N_883,N_7743);
nor U15878 (N_15878,N_4785,N_6566);
xnor U15879 (N_15879,N_7703,N_7037);
nor U15880 (N_15880,N_8653,N_4165);
nand U15881 (N_15881,N_3577,N_3653);
nand U15882 (N_15882,N_6305,N_3753);
xnor U15883 (N_15883,N_1637,N_8946);
nor U15884 (N_15884,N_7992,N_4228);
nor U15885 (N_15885,N_52,N_9288);
nand U15886 (N_15886,N_6705,N_4451);
and U15887 (N_15887,N_750,N_8918);
nor U15888 (N_15888,N_7663,N_1785);
or U15889 (N_15889,N_5247,N_4084);
xnor U15890 (N_15890,N_2941,N_7037);
nand U15891 (N_15891,N_8463,N_8182);
or U15892 (N_15892,N_9366,N_1807);
and U15893 (N_15893,N_1807,N_1830);
nand U15894 (N_15894,N_3547,N_1318);
nand U15895 (N_15895,N_7050,N_5599);
xnor U15896 (N_15896,N_4973,N_6050);
and U15897 (N_15897,N_7181,N_4034);
nor U15898 (N_15898,N_4345,N_1208);
xnor U15899 (N_15899,N_7509,N_904);
nor U15900 (N_15900,N_2901,N_6630);
and U15901 (N_15901,N_2596,N_321);
xnor U15902 (N_15902,N_8872,N_9604);
or U15903 (N_15903,N_9930,N_2938);
xor U15904 (N_15904,N_2299,N_3913);
nor U15905 (N_15905,N_9996,N_9129);
nand U15906 (N_15906,N_9381,N_3001);
and U15907 (N_15907,N_2597,N_2840);
nor U15908 (N_15908,N_2088,N_6630);
and U15909 (N_15909,N_6244,N_2666);
nor U15910 (N_15910,N_9662,N_7574);
nor U15911 (N_15911,N_4187,N_2705);
and U15912 (N_15912,N_223,N_4854);
nor U15913 (N_15913,N_8703,N_9611);
xnor U15914 (N_15914,N_7222,N_5981);
and U15915 (N_15915,N_3623,N_7897);
xor U15916 (N_15916,N_1417,N_4330);
and U15917 (N_15917,N_9641,N_2970);
xor U15918 (N_15918,N_4465,N_3385);
or U15919 (N_15919,N_5329,N_9241);
or U15920 (N_15920,N_2737,N_5219);
nor U15921 (N_15921,N_6980,N_5743);
nand U15922 (N_15922,N_3323,N_1108);
and U15923 (N_15923,N_4344,N_4022);
or U15924 (N_15924,N_7195,N_6926);
and U15925 (N_15925,N_5263,N_6237);
and U15926 (N_15926,N_3994,N_259);
nand U15927 (N_15927,N_6664,N_9728);
or U15928 (N_15928,N_3333,N_5783);
nand U15929 (N_15929,N_4716,N_9743);
or U15930 (N_15930,N_9307,N_5455);
or U15931 (N_15931,N_9759,N_3844);
and U15932 (N_15932,N_5382,N_1201);
nor U15933 (N_15933,N_9705,N_7394);
nor U15934 (N_15934,N_5031,N_4708);
nor U15935 (N_15935,N_3834,N_7129);
and U15936 (N_15936,N_6923,N_5542);
xor U15937 (N_15937,N_7994,N_5888);
nand U15938 (N_15938,N_5422,N_6935);
nor U15939 (N_15939,N_3763,N_1448);
nand U15940 (N_15940,N_3890,N_3000);
or U15941 (N_15941,N_4662,N_484);
xor U15942 (N_15942,N_6365,N_3578);
or U15943 (N_15943,N_2222,N_2243);
xnor U15944 (N_15944,N_530,N_7927);
xnor U15945 (N_15945,N_148,N_5085);
nor U15946 (N_15946,N_9866,N_6824);
or U15947 (N_15947,N_2042,N_8681);
nor U15948 (N_15948,N_2854,N_3809);
and U15949 (N_15949,N_4393,N_8052);
nor U15950 (N_15950,N_7331,N_5915);
nand U15951 (N_15951,N_1024,N_2777);
nand U15952 (N_15952,N_5080,N_7740);
or U15953 (N_15953,N_1258,N_8635);
xor U15954 (N_15954,N_1893,N_795);
or U15955 (N_15955,N_6759,N_7942);
xnor U15956 (N_15956,N_3671,N_4989);
nand U15957 (N_15957,N_247,N_8693);
and U15958 (N_15958,N_6805,N_9956);
nor U15959 (N_15959,N_3789,N_7508);
nand U15960 (N_15960,N_6829,N_3155);
and U15961 (N_15961,N_8946,N_461);
and U15962 (N_15962,N_1042,N_5564);
nand U15963 (N_15963,N_5957,N_2084);
xor U15964 (N_15964,N_652,N_3750);
and U15965 (N_15965,N_8978,N_3671);
nor U15966 (N_15966,N_5761,N_8794);
nor U15967 (N_15967,N_2684,N_1860);
nor U15968 (N_15968,N_705,N_9188);
nand U15969 (N_15969,N_9201,N_8622);
and U15970 (N_15970,N_1596,N_2743);
and U15971 (N_15971,N_5776,N_8064);
and U15972 (N_15972,N_5715,N_8829);
nor U15973 (N_15973,N_9516,N_1482);
xor U15974 (N_15974,N_4753,N_2572);
or U15975 (N_15975,N_8801,N_5011);
or U15976 (N_15976,N_964,N_4074);
nor U15977 (N_15977,N_9522,N_8971);
and U15978 (N_15978,N_9781,N_7328);
nand U15979 (N_15979,N_6031,N_1);
xnor U15980 (N_15980,N_9517,N_1629);
xnor U15981 (N_15981,N_4584,N_1470);
nand U15982 (N_15982,N_7936,N_5798);
xor U15983 (N_15983,N_8371,N_8782);
and U15984 (N_15984,N_3310,N_304);
and U15985 (N_15985,N_3265,N_5209);
xor U15986 (N_15986,N_7741,N_3013);
xnor U15987 (N_15987,N_8470,N_7298);
xnor U15988 (N_15988,N_9313,N_9144);
and U15989 (N_15989,N_5792,N_8133);
and U15990 (N_15990,N_976,N_3225);
xnor U15991 (N_15991,N_9548,N_7005);
nor U15992 (N_15992,N_2619,N_7778);
xor U15993 (N_15993,N_868,N_6061);
xor U15994 (N_15994,N_4520,N_5615);
xor U15995 (N_15995,N_8830,N_2523);
nand U15996 (N_15996,N_7698,N_3778);
xnor U15997 (N_15997,N_1465,N_2610);
and U15998 (N_15998,N_4883,N_6745);
and U15999 (N_15999,N_2560,N_8431);
and U16000 (N_16000,N_4270,N_6354);
or U16001 (N_16001,N_1230,N_3385);
nand U16002 (N_16002,N_5241,N_5728);
and U16003 (N_16003,N_3821,N_1467);
nand U16004 (N_16004,N_49,N_6483);
xor U16005 (N_16005,N_8051,N_6801);
nor U16006 (N_16006,N_3153,N_2918);
or U16007 (N_16007,N_1246,N_4692);
or U16008 (N_16008,N_4552,N_8371);
xnor U16009 (N_16009,N_4816,N_4830);
nor U16010 (N_16010,N_3770,N_1916);
xor U16011 (N_16011,N_1862,N_8440);
or U16012 (N_16012,N_2277,N_428);
nor U16013 (N_16013,N_9117,N_5508);
nand U16014 (N_16014,N_2159,N_8806);
xnor U16015 (N_16015,N_3987,N_1856);
nor U16016 (N_16016,N_5085,N_919);
nor U16017 (N_16017,N_9339,N_6314);
xnor U16018 (N_16018,N_5769,N_6088);
or U16019 (N_16019,N_9691,N_5591);
xnor U16020 (N_16020,N_6453,N_5930);
xor U16021 (N_16021,N_2349,N_2369);
nand U16022 (N_16022,N_6902,N_3732);
nor U16023 (N_16023,N_5162,N_5141);
nand U16024 (N_16024,N_7340,N_2784);
nand U16025 (N_16025,N_8468,N_6144);
or U16026 (N_16026,N_64,N_2183);
xnor U16027 (N_16027,N_5779,N_5581);
or U16028 (N_16028,N_9543,N_8669);
or U16029 (N_16029,N_1156,N_4383);
nor U16030 (N_16030,N_3663,N_8897);
or U16031 (N_16031,N_1277,N_3661);
nand U16032 (N_16032,N_4375,N_7901);
xor U16033 (N_16033,N_3433,N_3381);
nor U16034 (N_16034,N_9094,N_1815);
and U16035 (N_16035,N_6823,N_8952);
or U16036 (N_16036,N_844,N_5725);
xnor U16037 (N_16037,N_7630,N_1289);
nand U16038 (N_16038,N_7162,N_9003);
or U16039 (N_16039,N_415,N_9685);
nor U16040 (N_16040,N_6721,N_6761);
nor U16041 (N_16041,N_1279,N_7074);
or U16042 (N_16042,N_2023,N_3166);
nor U16043 (N_16043,N_4507,N_1259);
and U16044 (N_16044,N_5406,N_2245);
nand U16045 (N_16045,N_3464,N_4226);
xnor U16046 (N_16046,N_1835,N_8689);
nand U16047 (N_16047,N_5736,N_3308);
nand U16048 (N_16048,N_8001,N_8277);
and U16049 (N_16049,N_5005,N_7002);
or U16050 (N_16050,N_9125,N_3501);
and U16051 (N_16051,N_1806,N_5314);
nand U16052 (N_16052,N_6150,N_7640);
xnor U16053 (N_16053,N_5532,N_4270);
nor U16054 (N_16054,N_1250,N_2363);
and U16055 (N_16055,N_3672,N_1411);
xnor U16056 (N_16056,N_3639,N_4137);
or U16057 (N_16057,N_4474,N_9773);
or U16058 (N_16058,N_2007,N_6596);
or U16059 (N_16059,N_7962,N_2163);
or U16060 (N_16060,N_3083,N_3901);
nor U16061 (N_16061,N_6427,N_7504);
xor U16062 (N_16062,N_7074,N_6404);
xor U16063 (N_16063,N_6797,N_6733);
or U16064 (N_16064,N_8147,N_1737);
nand U16065 (N_16065,N_4482,N_6915);
xnor U16066 (N_16066,N_6291,N_457);
xnor U16067 (N_16067,N_1623,N_512);
xnor U16068 (N_16068,N_3336,N_4401);
and U16069 (N_16069,N_3320,N_9500);
or U16070 (N_16070,N_4173,N_6285);
and U16071 (N_16071,N_6862,N_4889);
nand U16072 (N_16072,N_6443,N_5226);
nand U16073 (N_16073,N_1012,N_8155);
or U16074 (N_16074,N_2279,N_1956);
xor U16075 (N_16075,N_2390,N_9908);
nand U16076 (N_16076,N_7587,N_8948);
xnor U16077 (N_16077,N_7426,N_2234);
or U16078 (N_16078,N_5954,N_1736);
nand U16079 (N_16079,N_4248,N_6853);
nor U16080 (N_16080,N_9280,N_5764);
and U16081 (N_16081,N_1565,N_8708);
xor U16082 (N_16082,N_3109,N_5563);
nand U16083 (N_16083,N_5884,N_1404);
or U16084 (N_16084,N_1334,N_4212);
xnor U16085 (N_16085,N_1214,N_7335);
nor U16086 (N_16086,N_8195,N_1827);
and U16087 (N_16087,N_9597,N_4678);
or U16088 (N_16088,N_86,N_2143);
xnor U16089 (N_16089,N_2192,N_8773);
or U16090 (N_16090,N_8478,N_5198);
nor U16091 (N_16091,N_6800,N_9836);
and U16092 (N_16092,N_2782,N_2689);
and U16093 (N_16093,N_8857,N_2856);
xnor U16094 (N_16094,N_4033,N_8213);
or U16095 (N_16095,N_3338,N_6958);
nand U16096 (N_16096,N_7356,N_211);
and U16097 (N_16097,N_1542,N_9327);
or U16098 (N_16098,N_6783,N_3946);
and U16099 (N_16099,N_393,N_6551);
and U16100 (N_16100,N_4465,N_3241);
nand U16101 (N_16101,N_6910,N_4521);
nand U16102 (N_16102,N_4219,N_3624);
nor U16103 (N_16103,N_5470,N_22);
nor U16104 (N_16104,N_9663,N_6104);
nor U16105 (N_16105,N_3368,N_5919);
nor U16106 (N_16106,N_735,N_8894);
or U16107 (N_16107,N_1266,N_3187);
and U16108 (N_16108,N_553,N_8060);
xor U16109 (N_16109,N_3089,N_2557);
and U16110 (N_16110,N_6948,N_2271);
nor U16111 (N_16111,N_8038,N_6501);
nor U16112 (N_16112,N_2277,N_3750);
or U16113 (N_16113,N_9731,N_8953);
nor U16114 (N_16114,N_4676,N_4819);
and U16115 (N_16115,N_2475,N_3889);
nor U16116 (N_16116,N_3764,N_1167);
nor U16117 (N_16117,N_4985,N_913);
xor U16118 (N_16118,N_9441,N_806);
nor U16119 (N_16119,N_1891,N_3269);
xor U16120 (N_16120,N_7039,N_2805);
and U16121 (N_16121,N_277,N_1470);
and U16122 (N_16122,N_2750,N_2517);
xnor U16123 (N_16123,N_9420,N_5194);
xnor U16124 (N_16124,N_7683,N_2584);
nor U16125 (N_16125,N_7274,N_285);
or U16126 (N_16126,N_5262,N_408);
or U16127 (N_16127,N_5548,N_3974);
and U16128 (N_16128,N_9937,N_7671);
and U16129 (N_16129,N_3074,N_1234);
nand U16130 (N_16130,N_3763,N_1919);
nor U16131 (N_16131,N_3185,N_5759);
and U16132 (N_16132,N_8848,N_7840);
nand U16133 (N_16133,N_3269,N_4309);
and U16134 (N_16134,N_6003,N_8620);
nand U16135 (N_16135,N_3674,N_896);
nor U16136 (N_16136,N_5064,N_8002);
and U16137 (N_16137,N_9683,N_6619);
and U16138 (N_16138,N_1431,N_9311);
nand U16139 (N_16139,N_8545,N_653);
xnor U16140 (N_16140,N_5912,N_4739);
nor U16141 (N_16141,N_606,N_9790);
nor U16142 (N_16142,N_3841,N_153);
xor U16143 (N_16143,N_4669,N_388);
nor U16144 (N_16144,N_3030,N_2345);
or U16145 (N_16145,N_8291,N_2372);
xnor U16146 (N_16146,N_51,N_388);
or U16147 (N_16147,N_2180,N_9765);
nand U16148 (N_16148,N_3527,N_4655);
or U16149 (N_16149,N_4721,N_9354);
xnor U16150 (N_16150,N_4612,N_5275);
xnor U16151 (N_16151,N_9116,N_3926);
and U16152 (N_16152,N_6665,N_23);
nor U16153 (N_16153,N_2051,N_8811);
nand U16154 (N_16154,N_8448,N_1899);
nand U16155 (N_16155,N_9731,N_8492);
xor U16156 (N_16156,N_7217,N_6372);
and U16157 (N_16157,N_3227,N_6926);
xor U16158 (N_16158,N_7013,N_1232);
xor U16159 (N_16159,N_4898,N_1833);
xor U16160 (N_16160,N_2641,N_7629);
nor U16161 (N_16161,N_3306,N_595);
or U16162 (N_16162,N_4555,N_9361);
or U16163 (N_16163,N_6931,N_2751);
xnor U16164 (N_16164,N_1020,N_8049);
xor U16165 (N_16165,N_9375,N_6582);
or U16166 (N_16166,N_2163,N_5656);
and U16167 (N_16167,N_1764,N_6576);
or U16168 (N_16168,N_7591,N_1096);
nand U16169 (N_16169,N_2828,N_3638);
or U16170 (N_16170,N_2699,N_5758);
xor U16171 (N_16171,N_3313,N_5267);
xor U16172 (N_16172,N_6957,N_7810);
nor U16173 (N_16173,N_3856,N_8375);
nand U16174 (N_16174,N_937,N_2718);
or U16175 (N_16175,N_4855,N_962);
or U16176 (N_16176,N_2238,N_9751);
and U16177 (N_16177,N_5640,N_5368);
or U16178 (N_16178,N_9639,N_1475);
nand U16179 (N_16179,N_3401,N_4961);
nor U16180 (N_16180,N_5034,N_3943);
xnor U16181 (N_16181,N_599,N_6453);
nor U16182 (N_16182,N_187,N_1335);
xor U16183 (N_16183,N_6704,N_3951);
xnor U16184 (N_16184,N_6505,N_6060);
or U16185 (N_16185,N_8835,N_4431);
or U16186 (N_16186,N_9577,N_1954);
nand U16187 (N_16187,N_6652,N_6641);
nor U16188 (N_16188,N_9920,N_2092);
or U16189 (N_16189,N_2344,N_9895);
or U16190 (N_16190,N_5021,N_5909);
nand U16191 (N_16191,N_9298,N_1413);
or U16192 (N_16192,N_3797,N_5790);
nand U16193 (N_16193,N_5900,N_5711);
xor U16194 (N_16194,N_9143,N_8948);
xnor U16195 (N_16195,N_6016,N_83);
and U16196 (N_16196,N_4130,N_2971);
nand U16197 (N_16197,N_6900,N_8323);
nand U16198 (N_16198,N_9592,N_2583);
nand U16199 (N_16199,N_2639,N_78);
xnor U16200 (N_16200,N_4065,N_7509);
nand U16201 (N_16201,N_5834,N_745);
nor U16202 (N_16202,N_6624,N_7780);
nor U16203 (N_16203,N_8487,N_7124);
xnor U16204 (N_16204,N_2536,N_6369);
nor U16205 (N_16205,N_6108,N_7892);
nand U16206 (N_16206,N_3359,N_1989);
or U16207 (N_16207,N_9253,N_7290);
xor U16208 (N_16208,N_9285,N_9615);
or U16209 (N_16209,N_8122,N_5242);
or U16210 (N_16210,N_1624,N_2261);
nand U16211 (N_16211,N_3933,N_194);
nor U16212 (N_16212,N_6095,N_7608);
nor U16213 (N_16213,N_2807,N_1795);
nand U16214 (N_16214,N_1457,N_6743);
or U16215 (N_16215,N_6330,N_8471);
nand U16216 (N_16216,N_5153,N_7758);
or U16217 (N_16217,N_2031,N_6842);
or U16218 (N_16218,N_3561,N_3353);
or U16219 (N_16219,N_7741,N_7134);
and U16220 (N_16220,N_995,N_2802);
nand U16221 (N_16221,N_4802,N_8898);
or U16222 (N_16222,N_7942,N_224);
or U16223 (N_16223,N_800,N_3001);
and U16224 (N_16224,N_9895,N_9102);
nand U16225 (N_16225,N_2516,N_8938);
and U16226 (N_16226,N_2648,N_6547);
xor U16227 (N_16227,N_8777,N_2370);
xor U16228 (N_16228,N_2387,N_9025);
nand U16229 (N_16229,N_6108,N_2924);
nand U16230 (N_16230,N_5682,N_3539);
and U16231 (N_16231,N_5754,N_9451);
and U16232 (N_16232,N_9425,N_854);
nor U16233 (N_16233,N_2547,N_5348);
and U16234 (N_16234,N_1278,N_7163);
nor U16235 (N_16235,N_3018,N_6469);
nand U16236 (N_16236,N_4812,N_2701);
nor U16237 (N_16237,N_6636,N_1387);
nor U16238 (N_16238,N_5173,N_1985);
nand U16239 (N_16239,N_4528,N_8211);
nor U16240 (N_16240,N_3913,N_3976);
nand U16241 (N_16241,N_5688,N_4206);
nor U16242 (N_16242,N_738,N_852);
nand U16243 (N_16243,N_2733,N_3427);
xnor U16244 (N_16244,N_8129,N_6302);
xnor U16245 (N_16245,N_8150,N_9066);
and U16246 (N_16246,N_9958,N_8994);
or U16247 (N_16247,N_7236,N_4194);
xor U16248 (N_16248,N_8073,N_6757);
or U16249 (N_16249,N_3730,N_5617);
nand U16250 (N_16250,N_5263,N_3294);
or U16251 (N_16251,N_1282,N_4926);
nor U16252 (N_16252,N_1344,N_3199);
nand U16253 (N_16253,N_4928,N_6591);
xnor U16254 (N_16254,N_1944,N_2062);
nor U16255 (N_16255,N_108,N_2886);
and U16256 (N_16256,N_5101,N_4168);
nand U16257 (N_16257,N_8620,N_529);
nor U16258 (N_16258,N_3554,N_1124);
nor U16259 (N_16259,N_2717,N_10);
and U16260 (N_16260,N_1037,N_4669);
xnor U16261 (N_16261,N_6179,N_8242);
nor U16262 (N_16262,N_4430,N_4232);
or U16263 (N_16263,N_2086,N_285);
and U16264 (N_16264,N_9372,N_9223);
nor U16265 (N_16265,N_8771,N_336);
xor U16266 (N_16266,N_9506,N_9602);
and U16267 (N_16267,N_957,N_6990);
or U16268 (N_16268,N_4563,N_5570);
and U16269 (N_16269,N_5681,N_5172);
nand U16270 (N_16270,N_8278,N_8258);
or U16271 (N_16271,N_4350,N_4403);
xnor U16272 (N_16272,N_2786,N_6796);
or U16273 (N_16273,N_5165,N_8972);
xnor U16274 (N_16274,N_2996,N_216);
nand U16275 (N_16275,N_576,N_7783);
nor U16276 (N_16276,N_2303,N_7834);
xor U16277 (N_16277,N_8969,N_5800);
or U16278 (N_16278,N_8943,N_1475);
or U16279 (N_16279,N_4431,N_5605);
nor U16280 (N_16280,N_1012,N_8814);
nor U16281 (N_16281,N_5570,N_1320);
nor U16282 (N_16282,N_7230,N_3910);
or U16283 (N_16283,N_1356,N_3732);
nor U16284 (N_16284,N_7181,N_4381);
and U16285 (N_16285,N_7111,N_2717);
xnor U16286 (N_16286,N_2209,N_6053);
nand U16287 (N_16287,N_8656,N_6851);
xnor U16288 (N_16288,N_7288,N_3724);
xor U16289 (N_16289,N_3729,N_273);
or U16290 (N_16290,N_6826,N_6591);
nor U16291 (N_16291,N_854,N_5566);
or U16292 (N_16292,N_7271,N_9842);
or U16293 (N_16293,N_8713,N_9422);
and U16294 (N_16294,N_3754,N_861);
and U16295 (N_16295,N_1860,N_6544);
or U16296 (N_16296,N_3528,N_9476);
xnor U16297 (N_16297,N_4237,N_1648);
nor U16298 (N_16298,N_338,N_8110);
nand U16299 (N_16299,N_7337,N_1246);
nand U16300 (N_16300,N_8334,N_1918);
nand U16301 (N_16301,N_1744,N_8380);
or U16302 (N_16302,N_2770,N_4377);
or U16303 (N_16303,N_387,N_1609);
xor U16304 (N_16304,N_9164,N_4641);
xnor U16305 (N_16305,N_9819,N_4464);
and U16306 (N_16306,N_2883,N_1447);
xor U16307 (N_16307,N_863,N_7042);
and U16308 (N_16308,N_2065,N_7593);
nor U16309 (N_16309,N_5718,N_7038);
nor U16310 (N_16310,N_5991,N_4842);
xnor U16311 (N_16311,N_3062,N_950);
nor U16312 (N_16312,N_8232,N_3635);
or U16313 (N_16313,N_7864,N_2589);
nand U16314 (N_16314,N_3207,N_7135);
or U16315 (N_16315,N_654,N_2196);
and U16316 (N_16316,N_6973,N_6259);
xor U16317 (N_16317,N_9722,N_3800);
nand U16318 (N_16318,N_5872,N_6168);
nand U16319 (N_16319,N_8809,N_87);
or U16320 (N_16320,N_7057,N_8916);
or U16321 (N_16321,N_8810,N_1753);
or U16322 (N_16322,N_1872,N_8040);
and U16323 (N_16323,N_8832,N_983);
nor U16324 (N_16324,N_7548,N_5059);
and U16325 (N_16325,N_5615,N_7036);
or U16326 (N_16326,N_6206,N_9783);
nor U16327 (N_16327,N_9219,N_8769);
nor U16328 (N_16328,N_7385,N_913);
xnor U16329 (N_16329,N_5931,N_4653);
or U16330 (N_16330,N_4463,N_2901);
and U16331 (N_16331,N_495,N_1664);
nor U16332 (N_16332,N_7472,N_638);
nand U16333 (N_16333,N_484,N_6826);
or U16334 (N_16334,N_7260,N_6313);
xor U16335 (N_16335,N_1140,N_1826);
nand U16336 (N_16336,N_2795,N_6546);
nor U16337 (N_16337,N_768,N_880);
and U16338 (N_16338,N_4714,N_6255);
nand U16339 (N_16339,N_6573,N_1001);
xor U16340 (N_16340,N_392,N_5720);
and U16341 (N_16341,N_4233,N_3050);
nor U16342 (N_16342,N_3438,N_954);
nand U16343 (N_16343,N_3123,N_240);
and U16344 (N_16344,N_6368,N_6212);
nor U16345 (N_16345,N_6351,N_9446);
and U16346 (N_16346,N_2326,N_6978);
or U16347 (N_16347,N_5418,N_3797);
and U16348 (N_16348,N_1750,N_4328);
nor U16349 (N_16349,N_3518,N_4225);
xnor U16350 (N_16350,N_1153,N_5566);
and U16351 (N_16351,N_9152,N_183);
nand U16352 (N_16352,N_9498,N_5576);
nor U16353 (N_16353,N_3488,N_9441);
and U16354 (N_16354,N_3360,N_3275);
or U16355 (N_16355,N_164,N_7464);
or U16356 (N_16356,N_5049,N_6675);
and U16357 (N_16357,N_8006,N_8038);
nor U16358 (N_16358,N_4579,N_1165);
or U16359 (N_16359,N_180,N_760);
and U16360 (N_16360,N_467,N_217);
xor U16361 (N_16361,N_7733,N_3371);
and U16362 (N_16362,N_8874,N_7449);
or U16363 (N_16363,N_2419,N_7847);
nand U16364 (N_16364,N_9531,N_1496);
and U16365 (N_16365,N_5388,N_4337);
xor U16366 (N_16366,N_4985,N_140);
xor U16367 (N_16367,N_8643,N_2628);
nor U16368 (N_16368,N_7112,N_7122);
nand U16369 (N_16369,N_443,N_9836);
and U16370 (N_16370,N_1022,N_74);
or U16371 (N_16371,N_1574,N_7794);
or U16372 (N_16372,N_8714,N_22);
or U16373 (N_16373,N_4629,N_8685);
or U16374 (N_16374,N_3768,N_926);
xnor U16375 (N_16375,N_5740,N_9390);
nor U16376 (N_16376,N_2074,N_4240);
or U16377 (N_16377,N_2173,N_9180);
xnor U16378 (N_16378,N_7597,N_5692);
or U16379 (N_16379,N_2613,N_9003);
nor U16380 (N_16380,N_7839,N_9471);
nand U16381 (N_16381,N_7700,N_656);
and U16382 (N_16382,N_2509,N_952);
xnor U16383 (N_16383,N_2099,N_670);
xor U16384 (N_16384,N_6544,N_5400);
or U16385 (N_16385,N_9850,N_6112);
and U16386 (N_16386,N_3128,N_6122);
or U16387 (N_16387,N_7498,N_8969);
and U16388 (N_16388,N_4002,N_6243);
and U16389 (N_16389,N_2276,N_665);
or U16390 (N_16390,N_6023,N_5501);
and U16391 (N_16391,N_1185,N_7815);
xnor U16392 (N_16392,N_8739,N_6454);
nor U16393 (N_16393,N_7642,N_1506);
nor U16394 (N_16394,N_6010,N_7026);
and U16395 (N_16395,N_813,N_3227);
and U16396 (N_16396,N_6328,N_2587);
nand U16397 (N_16397,N_4189,N_4753);
or U16398 (N_16398,N_3457,N_5892);
xnor U16399 (N_16399,N_1537,N_3283);
and U16400 (N_16400,N_5120,N_469);
or U16401 (N_16401,N_4425,N_5719);
nand U16402 (N_16402,N_7534,N_2548);
or U16403 (N_16403,N_1476,N_3248);
and U16404 (N_16404,N_6337,N_9557);
or U16405 (N_16405,N_6497,N_6077);
or U16406 (N_16406,N_6880,N_1229);
nor U16407 (N_16407,N_6499,N_3669);
and U16408 (N_16408,N_4099,N_6872);
nor U16409 (N_16409,N_2751,N_1574);
and U16410 (N_16410,N_9004,N_2130);
xor U16411 (N_16411,N_658,N_34);
nor U16412 (N_16412,N_4321,N_6759);
nor U16413 (N_16413,N_9455,N_2377);
or U16414 (N_16414,N_3313,N_9874);
and U16415 (N_16415,N_7484,N_1384);
nor U16416 (N_16416,N_9455,N_691);
or U16417 (N_16417,N_6659,N_7254);
nand U16418 (N_16418,N_6881,N_128);
and U16419 (N_16419,N_998,N_5939);
and U16420 (N_16420,N_4264,N_7434);
and U16421 (N_16421,N_7914,N_2112);
or U16422 (N_16422,N_5952,N_541);
xnor U16423 (N_16423,N_614,N_910);
or U16424 (N_16424,N_6808,N_1353);
nand U16425 (N_16425,N_7346,N_4134);
nand U16426 (N_16426,N_4460,N_3958);
nor U16427 (N_16427,N_6115,N_6308);
nand U16428 (N_16428,N_8476,N_2093);
nand U16429 (N_16429,N_3451,N_2403);
xnor U16430 (N_16430,N_9632,N_561);
or U16431 (N_16431,N_2793,N_7952);
or U16432 (N_16432,N_3595,N_4085);
or U16433 (N_16433,N_9596,N_8598);
and U16434 (N_16434,N_7506,N_7966);
and U16435 (N_16435,N_9597,N_8791);
nand U16436 (N_16436,N_9305,N_5900);
nor U16437 (N_16437,N_2871,N_363);
or U16438 (N_16438,N_626,N_7675);
and U16439 (N_16439,N_6652,N_4684);
nand U16440 (N_16440,N_5399,N_3595);
or U16441 (N_16441,N_2274,N_5104);
or U16442 (N_16442,N_2300,N_1932);
or U16443 (N_16443,N_4910,N_6630);
or U16444 (N_16444,N_602,N_382);
and U16445 (N_16445,N_7886,N_3977);
and U16446 (N_16446,N_5101,N_7527);
nor U16447 (N_16447,N_3382,N_9405);
or U16448 (N_16448,N_2709,N_9946);
and U16449 (N_16449,N_7671,N_8369);
nand U16450 (N_16450,N_3445,N_9822);
nand U16451 (N_16451,N_1959,N_3888);
xnor U16452 (N_16452,N_8707,N_1882);
or U16453 (N_16453,N_689,N_3976);
nor U16454 (N_16454,N_2068,N_4871);
nand U16455 (N_16455,N_2444,N_1462);
nand U16456 (N_16456,N_8217,N_9812);
or U16457 (N_16457,N_5100,N_2230);
and U16458 (N_16458,N_8017,N_1702);
nand U16459 (N_16459,N_9614,N_2119);
or U16460 (N_16460,N_8101,N_8377);
or U16461 (N_16461,N_7741,N_5973);
and U16462 (N_16462,N_4269,N_2064);
and U16463 (N_16463,N_3729,N_8725);
nand U16464 (N_16464,N_4245,N_3887);
nor U16465 (N_16465,N_5644,N_5244);
and U16466 (N_16466,N_6849,N_2533);
xor U16467 (N_16467,N_9050,N_9608);
nor U16468 (N_16468,N_6044,N_4132);
or U16469 (N_16469,N_9924,N_2187);
and U16470 (N_16470,N_3875,N_2442);
xor U16471 (N_16471,N_1416,N_5868);
nand U16472 (N_16472,N_6880,N_5356);
nor U16473 (N_16473,N_5808,N_2787);
or U16474 (N_16474,N_9019,N_4852);
xnor U16475 (N_16475,N_9881,N_1804);
and U16476 (N_16476,N_8834,N_3127);
and U16477 (N_16477,N_8455,N_2465);
and U16478 (N_16478,N_3905,N_3188);
or U16479 (N_16479,N_1539,N_6883);
nand U16480 (N_16480,N_6743,N_4141);
nor U16481 (N_16481,N_679,N_5944);
and U16482 (N_16482,N_6985,N_9440);
xnor U16483 (N_16483,N_3606,N_463);
and U16484 (N_16484,N_9562,N_3512);
and U16485 (N_16485,N_3104,N_9556);
nand U16486 (N_16486,N_582,N_1369);
and U16487 (N_16487,N_664,N_9546);
nand U16488 (N_16488,N_4494,N_415);
or U16489 (N_16489,N_3218,N_7914);
and U16490 (N_16490,N_265,N_2168);
xor U16491 (N_16491,N_3857,N_4391);
or U16492 (N_16492,N_8820,N_3286);
and U16493 (N_16493,N_5424,N_4745);
and U16494 (N_16494,N_2013,N_6552);
xor U16495 (N_16495,N_3502,N_4724);
nor U16496 (N_16496,N_9896,N_3118);
or U16497 (N_16497,N_616,N_7664);
nand U16498 (N_16498,N_3016,N_8059);
or U16499 (N_16499,N_5100,N_9939);
or U16500 (N_16500,N_1933,N_4370);
nand U16501 (N_16501,N_2394,N_9423);
and U16502 (N_16502,N_2672,N_5279);
or U16503 (N_16503,N_5062,N_735);
nand U16504 (N_16504,N_4605,N_4871);
nor U16505 (N_16505,N_1455,N_7591);
nor U16506 (N_16506,N_762,N_6559);
or U16507 (N_16507,N_7039,N_3293);
nor U16508 (N_16508,N_2067,N_3174);
or U16509 (N_16509,N_7747,N_8904);
nand U16510 (N_16510,N_2251,N_7804);
and U16511 (N_16511,N_853,N_9052);
xnor U16512 (N_16512,N_3457,N_6134);
nand U16513 (N_16513,N_9323,N_4812);
xnor U16514 (N_16514,N_7285,N_2085);
nor U16515 (N_16515,N_2616,N_34);
or U16516 (N_16516,N_99,N_7195);
nor U16517 (N_16517,N_5399,N_5521);
nor U16518 (N_16518,N_6671,N_6519);
xnor U16519 (N_16519,N_8502,N_2727);
nor U16520 (N_16520,N_7768,N_1815);
nor U16521 (N_16521,N_6342,N_7446);
nand U16522 (N_16522,N_7614,N_4706);
nand U16523 (N_16523,N_141,N_171);
or U16524 (N_16524,N_7008,N_1360);
and U16525 (N_16525,N_9883,N_7077);
and U16526 (N_16526,N_690,N_4240);
nand U16527 (N_16527,N_1752,N_1985);
and U16528 (N_16528,N_7193,N_1952);
or U16529 (N_16529,N_9759,N_5729);
nand U16530 (N_16530,N_6292,N_1553);
nor U16531 (N_16531,N_2446,N_976);
or U16532 (N_16532,N_855,N_9308);
nor U16533 (N_16533,N_564,N_3107);
nand U16534 (N_16534,N_3188,N_65);
xor U16535 (N_16535,N_28,N_3119);
and U16536 (N_16536,N_6897,N_6310);
xnor U16537 (N_16537,N_242,N_5553);
or U16538 (N_16538,N_7983,N_2255);
nor U16539 (N_16539,N_848,N_6693);
nand U16540 (N_16540,N_7163,N_571);
nand U16541 (N_16541,N_3581,N_951);
nand U16542 (N_16542,N_4737,N_5284);
and U16543 (N_16543,N_7224,N_8445);
nor U16544 (N_16544,N_5060,N_2008);
nor U16545 (N_16545,N_5625,N_4504);
and U16546 (N_16546,N_3764,N_9374);
xor U16547 (N_16547,N_788,N_6322);
xnor U16548 (N_16548,N_9933,N_8085);
nor U16549 (N_16549,N_5031,N_221);
xor U16550 (N_16550,N_881,N_437);
nand U16551 (N_16551,N_7586,N_5456);
and U16552 (N_16552,N_4428,N_4224);
nor U16553 (N_16553,N_1356,N_9852);
xor U16554 (N_16554,N_9031,N_4305);
or U16555 (N_16555,N_7651,N_4723);
nor U16556 (N_16556,N_3795,N_7774);
and U16557 (N_16557,N_8451,N_8786);
and U16558 (N_16558,N_7003,N_6604);
nand U16559 (N_16559,N_6260,N_8802);
or U16560 (N_16560,N_6281,N_5420);
and U16561 (N_16561,N_1843,N_9538);
nand U16562 (N_16562,N_3517,N_1230);
xnor U16563 (N_16563,N_2514,N_4160);
or U16564 (N_16564,N_5734,N_6666);
and U16565 (N_16565,N_3072,N_2352);
nor U16566 (N_16566,N_8847,N_5609);
nor U16567 (N_16567,N_5438,N_3919);
and U16568 (N_16568,N_8962,N_8310);
nand U16569 (N_16569,N_3997,N_7265);
xnor U16570 (N_16570,N_7563,N_3416);
nor U16571 (N_16571,N_6054,N_6966);
or U16572 (N_16572,N_9422,N_2943);
xnor U16573 (N_16573,N_1392,N_1310);
and U16574 (N_16574,N_6619,N_1832);
nor U16575 (N_16575,N_1818,N_210);
nand U16576 (N_16576,N_7914,N_9417);
and U16577 (N_16577,N_6121,N_9684);
and U16578 (N_16578,N_3157,N_3755);
and U16579 (N_16579,N_7078,N_8477);
xor U16580 (N_16580,N_9814,N_6139);
xnor U16581 (N_16581,N_5897,N_3819);
xor U16582 (N_16582,N_4087,N_9217);
and U16583 (N_16583,N_1363,N_8398);
and U16584 (N_16584,N_5329,N_4426);
nand U16585 (N_16585,N_2840,N_4329);
nor U16586 (N_16586,N_59,N_7654);
and U16587 (N_16587,N_4577,N_6831);
and U16588 (N_16588,N_9949,N_5726);
xor U16589 (N_16589,N_497,N_7917);
or U16590 (N_16590,N_851,N_6588);
and U16591 (N_16591,N_5574,N_5653);
nand U16592 (N_16592,N_2090,N_41);
xnor U16593 (N_16593,N_5771,N_6849);
nand U16594 (N_16594,N_1420,N_7217);
nand U16595 (N_16595,N_1321,N_8833);
nor U16596 (N_16596,N_1832,N_5271);
and U16597 (N_16597,N_9344,N_1675);
and U16598 (N_16598,N_2842,N_4537);
nand U16599 (N_16599,N_9825,N_7678);
xnor U16600 (N_16600,N_1916,N_7051);
or U16601 (N_16601,N_4669,N_7786);
or U16602 (N_16602,N_3611,N_5826);
xor U16603 (N_16603,N_6544,N_9672);
xor U16604 (N_16604,N_7194,N_2909);
or U16605 (N_16605,N_2718,N_4283);
xor U16606 (N_16606,N_3761,N_2300);
and U16607 (N_16607,N_4111,N_6721);
nand U16608 (N_16608,N_6731,N_3999);
or U16609 (N_16609,N_6872,N_4415);
or U16610 (N_16610,N_5020,N_5250);
nand U16611 (N_16611,N_5800,N_1220);
nand U16612 (N_16612,N_6139,N_7760);
nor U16613 (N_16613,N_6161,N_9806);
nor U16614 (N_16614,N_6702,N_2461);
xor U16615 (N_16615,N_5439,N_6011);
xor U16616 (N_16616,N_8216,N_738);
nor U16617 (N_16617,N_6738,N_4669);
nor U16618 (N_16618,N_6487,N_142);
and U16619 (N_16619,N_9551,N_1157);
or U16620 (N_16620,N_1733,N_7802);
and U16621 (N_16621,N_5079,N_7531);
or U16622 (N_16622,N_2761,N_4490);
nor U16623 (N_16623,N_5018,N_6178);
or U16624 (N_16624,N_6303,N_9078);
nand U16625 (N_16625,N_2623,N_9022);
nor U16626 (N_16626,N_6228,N_5542);
xor U16627 (N_16627,N_7472,N_4798);
and U16628 (N_16628,N_1748,N_9754);
or U16629 (N_16629,N_3560,N_1835);
xnor U16630 (N_16630,N_103,N_1055);
xor U16631 (N_16631,N_7918,N_1954);
xnor U16632 (N_16632,N_3117,N_6580);
nor U16633 (N_16633,N_9304,N_5163);
xnor U16634 (N_16634,N_1959,N_4908);
or U16635 (N_16635,N_2408,N_1605);
xor U16636 (N_16636,N_8971,N_508);
xor U16637 (N_16637,N_9062,N_2707);
and U16638 (N_16638,N_4916,N_4719);
xnor U16639 (N_16639,N_479,N_4693);
xor U16640 (N_16640,N_3196,N_1840);
nand U16641 (N_16641,N_2278,N_9906);
and U16642 (N_16642,N_4622,N_54);
nor U16643 (N_16643,N_8759,N_999);
nand U16644 (N_16644,N_4237,N_4433);
nand U16645 (N_16645,N_6972,N_9777);
nand U16646 (N_16646,N_2201,N_9974);
nor U16647 (N_16647,N_3384,N_1846);
and U16648 (N_16648,N_7055,N_2994);
or U16649 (N_16649,N_4715,N_1876);
nor U16650 (N_16650,N_445,N_876);
and U16651 (N_16651,N_6740,N_3363);
xnor U16652 (N_16652,N_6523,N_9320);
nand U16653 (N_16653,N_3084,N_2381);
nor U16654 (N_16654,N_9346,N_4110);
and U16655 (N_16655,N_3659,N_1339);
xnor U16656 (N_16656,N_8070,N_436);
nor U16657 (N_16657,N_441,N_7467);
xor U16658 (N_16658,N_4598,N_8514);
and U16659 (N_16659,N_3347,N_2419);
xnor U16660 (N_16660,N_1192,N_2886);
nand U16661 (N_16661,N_1950,N_5766);
and U16662 (N_16662,N_1126,N_7301);
nor U16663 (N_16663,N_3689,N_3282);
nor U16664 (N_16664,N_6285,N_6293);
nand U16665 (N_16665,N_9506,N_8124);
or U16666 (N_16666,N_7369,N_6763);
xnor U16667 (N_16667,N_1007,N_9122);
and U16668 (N_16668,N_7882,N_8040);
xor U16669 (N_16669,N_4608,N_648);
xnor U16670 (N_16670,N_7953,N_5403);
and U16671 (N_16671,N_3637,N_9764);
nor U16672 (N_16672,N_1195,N_3170);
and U16673 (N_16673,N_9032,N_1395);
or U16674 (N_16674,N_5703,N_2678);
and U16675 (N_16675,N_610,N_2322);
or U16676 (N_16676,N_3883,N_4688);
or U16677 (N_16677,N_7430,N_4404);
and U16678 (N_16678,N_6232,N_8337);
nor U16679 (N_16679,N_6978,N_3972);
nand U16680 (N_16680,N_7107,N_1093);
and U16681 (N_16681,N_409,N_7050);
and U16682 (N_16682,N_845,N_6599);
or U16683 (N_16683,N_4049,N_3737);
and U16684 (N_16684,N_7296,N_8391);
nand U16685 (N_16685,N_1389,N_8892);
and U16686 (N_16686,N_1938,N_4192);
nand U16687 (N_16687,N_867,N_3186);
xnor U16688 (N_16688,N_5423,N_5793);
xnor U16689 (N_16689,N_2739,N_4866);
nor U16690 (N_16690,N_8569,N_1097);
nor U16691 (N_16691,N_5440,N_9175);
xnor U16692 (N_16692,N_7887,N_5690);
nand U16693 (N_16693,N_9037,N_7305);
nor U16694 (N_16694,N_2055,N_3720);
xnor U16695 (N_16695,N_4571,N_7603);
nor U16696 (N_16696,N_2613,N_7334);
xor U16697 (N_16697,N_5700,N_4409);
xor U16698 (N_16698,N_4867,N_1530);
and U16699 (N_16699,N_9068,N_4248);
nor U16700 (N_16700,N_8486,N_9492);
xor U16701 (N_16701,N_8289,N_5060);
and U16702 (N_16702,N_6952,N_7085);
and U16703 (N_16703,N_9931,N_6639);
nor U16704 (N_16704,N_249,N_4066);
or U16705 (N_16705,N_4504,N_3366);
or U16706 (N_16706,N_6274,N_8695);
nor U16707 (N_16707,N_516,N_3871);
nand U16708 (N_16708,N_906,N_5671);
and U16709 (N_16709,N_9413,N_8230);
nor U16710 (N_16710,N_4685,N_6694);
and U16711 (N_16711,N_5223,N_2089);
nand U16712 (N_16712,N_2928,N_7017);
xnor U16713 (N_16713,N_4226,N_3430);
nand U16714 (N_16714,N_5029,N_2271);
or U16715 (N_16715,N_2644,N_3818);
xnor U16716 (N_16716,N_7097,N_4126);
xnor U16717 (N_16717,N_1303,N_4119);
xor U16718 (N_16718,N_8371,N_9817);
xor U16719 (N_16719,N_4264,N_6013);
nor U16720 (N_16720,N_2483,N_7451);
nand U16721 (N_16721,N_9068,N_673);
and U16722 (N_16722,N_8158,N_7418);
nand U16723 (N_16723,N_4465,N_7656);
nand U16724 (N_16724,N_1715,N_6886);
and U16725 (N_16725,N_6818,N_5996);
nand U16726 (N_16726,N_915,N_2949);
xnor U16727 (N_16727,N_7525,N_8364);
and U16728 (N_16728,N_7394,N_2466);
or U16729 (N_16729,N_2037,N_744);
nand U16730 (N_16730,N_1923,N_4764);
or U16731 (N_16731,N_7506,N_2952);
or U16732 (N_16732,N_407,N_4493);
and U16733 (N_16733,N_3794,N_3815);
xor U16734 (N_16734,N_3352,N_1900);
nor U16735 (N_16735,N_3844,N_2815);
nor U16736 (N_16736,N_3818,N_9304);
nor U16737 (N_16737,N_1731,N_6995);
nand U16738 (N_16738,N_2851,N_6195);
and U16739 (N_16739,N_8016,N_8700);
xor U16740 (N_16740,N_6723,N_7378);
or U16741 (N_16741,N_9633,N_6314);
xor U16742 (N_16742,N_5212,N_92);
and U16743 (N_16743,N_6678,N_6491);
or U16744 (N_16744,N_4314,N_6089);
xor U16745 (N_16745,N_119,N_6046);
or U16746 (N_16746,N_55,N_696);
xnor U16747 (N_16747,N_6537,N_7833);
nand U16748 (N_16748,N_5456,N_572);
xor U16749 (N_16749,N_6199,N_9511);
nand U16750 (N_16750,N_7004,N_5341);
nor U16751 (N_16751,N_296,N_4906);
and U16752 (N_16752,N_2933,N_4597);
xor U16753 (N_16753,N_4248,N_7944);
xnor U16754 (N_16754,N_2131,N_9077);
and U16755 (N_16755,N_4383,N_4858);
xnor U16756 (N_16756,N_4271,N_8764);
or U16757 (N_16757,N_8560,N_3006);
nand U16758 (N_16758,N_3605,N_9491);
xor U16759 (N_16759,N_7634,N_5373);
and U16760 (N_16760,N_5387,N_890);
or U16761 (N_16761,N_3830,N_9667);
xor U16762 (N_16762,N_3586,N_939);
or U16763 (N_16763,N_9341,N_3521);
and U16764 (N_16764,N_7186,N_4078);
xor U16765 (N_16765,N_2549,N_6665);
nor U16766 (N_16766,N_6642,N_3197);
nand U16767 (N_16767,N_5382,N_8580);
xnor U16768 (N_16768,N_5087,N_6993);
or U16769 (N_16769,N_2295,N_9410);
nor U16770 (N_16770,N_3709,N_2602);
or U16771 (N_16771,N_9374,N_1281);
nor U16772 (N_16772,N_9333,N_9480);
xnor U16773 (N_16773,N_118,N_1702);
xnor U16774 (N_16774,N_6427,N_7055);
or U16775 (N_16775,N_3740,N_9923);
and U16776 (N_16776,N_9994,N_6687);
and U16777 (N_16777,N_974,N_2797);
and U16778 (N_16778,N_7142,N_7567);
and U16779 (N_16779,N_5667,N_5313);
nand U16780 (N_16780,N_2716,N_4783);
and U16781 (N_16781,N_3001,N_1499);
nand U16782 (N_16782,N_1821,N_9793);
nor U16783 (N_16783,N_5071,N_8855);
nand U16784 (N_16784,N_7579,N_5956);
and U16785 (N_16785,N_4763,N_7181);
and U16786 (N_16786,N_313,N_2739);
nand U16787 (N_16787,N_719,N_2291);
or U16788 (N_16788,N_2984,N_3881);
xor U16789 (N_16789,N_7389,N_1808);
nand U16790 (N_16790,N_9589,N_1582);
nor U16791 (N_16791,N_8513,N_9716);
nand U16792 (N_16792,N_8681,N_8830);
or U16793 (N_16793,N_6572,N_1033);
nor U16794 (N_16794,N_9496,N_9571);
or U16795 (N_16795,N_7486,N_7946);
xnor U16796 (N_16796,N_5866,N_4586);
or U16797 (N_16797,N_7871,N_7810);
or U16798 (N_16798,N_2783,N_4145);
xnor U16799 (N_16799,N_7523,N_9641);
or U16800 (N_16800,N_437,N_1123);
nand U16801 (N_16801,N_4214,N_2220);
nor U16802 (N_16802,N_2561,N_1427);
xnor U16803 (N_16803,N_6512,N_8960);
and U16804 (N_16804,N_6072,N_9140);
nor U16805 (N_16805,N_9053,N_2825);
and U16806 (N_16806,N_7575,N_1511);
xnor U16807 (N_16807,N_418,N_7985);
xor U16808 (N_16808,N_9396,N_5521);
nand U16809 (N_16809,N_1510,N_2588);
nor U16810 (N_16810,N_2732,N_1843);
nand U16811 (N_16811,N_3426,N_6676);
xnor U16812 (N_16812,N_2062,N_8704);
xor U16813 (N_16813,N_3232,N_6317);
nor U16814 (N_16814,N_3006,N_4814);
and U16815 (N_16815,N_8335,N_1305);
and U16816 (N_16816,N_8773,N_851);
or U16817 (N_16817,N_1455,N_8858);
nor U16818 (N_16818,N_4602,N_7388);
and U16819 (N_16819,N_4600,N_8093);
nor U16820 (N_16820,N_7648,N_6049);
or U16821 (N_16821,N_733,N_3409);
or U16822 (N_16822,N_4640,N_4121);
nand U16823 (N_16823,N_6117,N_6322);
xor U16824 (N_16824,N_9997,N_9675);
or U16825 (N_16825,N_6325,N_4132);
nand U16826 (N_16826,N_2345,N_3002);
nand U16827 (N_16827,N_4229,N_6048);
and U16828 (N_16828,N_1135,N_2694);
or U16829 (N_16829,N_4002,N_946);
nor U16830 (N_16830,N_2706,N_6172);
nor U16831 (N_16831,N_9202,N_8375);
or U16832 (N_16832,N_9336,N_1359);
nor U16833 (N_16833,N_661,N_9508);
nand U16834 (N_16834,N_9935,N_7663);
nand U16835 (N_16835,N_1573,N_6591);
and U16836 (N_16836,N_6964,N_652);
or U16837 (N_16837,N_8776,N_3613);
xor U16838 (N_16838,N_931,N_274);
nand U16839 (N_16839,N_3728,N_7594);
nand U16840 (N_16840,N_1484,N_8033);
nand U16841 (N_16841,N_5183,N_852);
or U16842 (N_16842,N_664,N_3096);
or U16843 (N_16843,N_3180,N_3876);
nor U16844 (N_16844,N_5371,N_9344);
xor U16845 (N_16845,N_2036,N_1035);
or U16846 (N_16846,N_7255,N_6490);
nand U16847 (N_16847,N_1728,N_2962);
and U16848 (N_16848,N_2547,N_4969);
xnor U16849 (N_16849,N_6256,N_447);
nand U16850 (N_16850,N_8958,N_7002);
or U16851 (N_16851,N_7750,N_7892);
and U16852 (N_16852,N_2869,N_5216);
nor U16853 (N_16853,N_1485,N_5242);
xnor U16854 (N_16854,N_6532,N_5869);
xnor U16855 (N_16855,N_5393,N_1392);
and U16856 (N_16856,N_9706,N_6388);
nand U16857 (N_16857,N_542,N_8086);
nor U16858 (N_16858,N_5786,N_365);
nor U16859 (N_16859,N_9953,N_8115);
nand U16860 (N_16860,N_189,N_7044);
or U16861 (N_16861,N_887,N_2979);
or U16862 (N_16862,N_7665,N_8567);
xnor U16863 (N_16863,N_554,N_7642);
nor U16864 (N_16864,N_3246,N_5501);
or U16865 (N_16865,N_4661,N_110);
nor U16866 (N_16866,N_4565,N_2896);
nor U16867 (N_16867,N_2213,N_45);
or U16868 (N_16868,N_7321,N_4612);
xnor U16869 (N_16869,N_8301,N_2199);
and U16870 (N_16870,N_5384,N_6476);
xor U16871 (N_16871,N_7242,N_1969);
and U16872 (N_16872,N_7015,N_7911);
nand U16873 (N_16873,N_5993,N_4604);
and U16874 (N_16874,N_4444,N_3013);
and U16875 (N_16875,N_723,N_4990);
xor U16876 (N_16876,N_8123,N_3735);
nand U16877 (N_16877,N_8380,N_5322);
and U16878 (N_16878,N_809,N_4609);
nor U16879 (N_16879,N_2751,N_8145);
and U16880 (N_16880,N_8561,N_7066);
or U16881 (N_16881,N_6422,N_3586);
or U16882 (N_16882,N_6728,N_4481);
nand U16883 (N_16883,N_8527,N_5121);
or U16884 (N_16884,N_3293,N_5349);
nor U16885 (N_16885,N_4349,N_7266);
and U16886 (N_16886,N_995,N_1302);
nor U16887 (N_16887,N_6854,N_6213);
nand U16888 (N_16888,N_42,N_2619);
xnor U16889 (N_16889,N_5871,N_4663);
nand U16890 (N_16890,N_9249,N_7);
xor U16891 (N_16891,N_3005,N_4167);
and U16892 (N_16892,N_4698,N_3147);
xnor U16893 (N_16893,N_9153,N_5302);
xnor U16894 (N_16894,N_8473,N_3545);
or U16895 (N_16895,N_3657,N_3741);
or U16896 (N_16896,N_4748,N_8448);
xnor U16897 (N_16897,N_7573,N_3932);
nand U16898 (N_16898,N_6054,N_1469);
nand U16899 (N_16899,N_5554,N_402);
nor U16900 (N_16900,N_3607,N_5394);
or U16901 (N_16901,N_2025,N_9485);
nand U16902 (N_16902,N_2459,N_3420);
or U16903 (N_16903,N_4254,N_5226);
nand U16904 (N_16904,N_6041,N_1180);
xor U16905 (N_16905,N_2547,N_2616);
and U16906 (N_16906,N_8497,N_2255);
xnor U16907 (N_16907,N_4806,N_7608);
nor U16908 (N_16908,N_113,N_6591);
xor U16909 (N_16909,N_5956,N_3059);
nor U16910 (N_16910,N_627,N_1276);
nand U16911 (N_16911,N_7253,N_5434);
nand U16912 (N_16912,N_3996,N_5801);
and U16913 (N_16913,N_4928,N_6664);
or U16914 (N_16914,N_9263,N_2174);
or U16915 (N_16915,N_6862,N_5117);
xor U16916 (N_16916,N_5700,N_5451);
and U16917 (N_16917,N_9060,N_6045);
xor U16918 (N_16918,N_6495,N_2621);
xor U16919 (N_16919,N_3467,N_6375);
and U16920 (N_16920,N_5260,N_4122);
xnor U16921 (N_16921,N_5117,N_5152);
nor U16922 (N_16922,N_8395,N_8384);
or U16923 (N_16923,N_5309,N_7161);
and U16924 (N_16924,N_6203,N_7959);
xor U16925 (N_16925,N_9084,N_6748);
or U16926 (N_16926,N_4658,N_8125);
nand U16927 (N_16927,N_2954,N_316);
nor U16928 (N_16928,N_6448,N_4723);
nor U16929 (N_16929,N_4521,N_3858);
or U16930 (N_16930,N_2824,N_4052);
nor U16931 (N_16931,N_8852,N_9925);
nor U16932 (N_16932,N_9863,N_7924);
and U16933 (N_16933,N_8602,N_4086);
or U16934 (N_16934,N_5668,N_394);
and U16935 (N_16935,N_4528,N_5376);
xor U16936 (N_16936,N_9227,N_9285);
xor U16937 (N_16937,N_5545,N_3977);
xnor U16938 (N_16938,N_8345,N_8483);
or U16939 (N_16939,N_1618,N_7899);
and U16940 (N_16940,N_4830,N_7256);
nor U16941 (N_16941,N_8702,N_3161);
or U16942 (N_16942,N_2117,N_9233);
or U16943 (N_16943,N_2572,N_2574);
nor U16944 (N_16944,N_1097,N_9996);
or U16945 (N_16945,N_3113,N_9226);
nand U16946 (N_16946,N_3798,N_7621);
or U16947 (N_16947,N_5422,N_227);
xor U16948 (N_16948,N_6729,N_6728);
xor U16949 (N_16949,N_840,N_3417);
xnor U16950 (N_16950,N_5256,N_501);
xnor U16951 (N_16951,N_8901,N_2513);
nand U16952 (N_16952,N_7669,N_8147);
xor U16953 (N_16953,N_5591,N_2592);
or U16954 (N_16954,N_6676,N_6609);
or U16955 (N_16955,N_9531,N_9047);
xnor U16956 (N_16956,N_4339,N_1298);
xnor U16957 (N_16957,N_5615,N_1716);
or U16958 (N_16958,N_2757,N_2412);
nor U16959 (N_16959,N_4053,N_8225);
and U16960 (N_16960,N_8781,N_7300);
nand U16961 (N_16961,N_5024,N_2122);
nand U16962 (N_16962,N_767,N_6288);
nor U16963 (N_16963,N_753,N_9053);
and U16964 (N_16964,N_9913,N_3035);
nor U16965 (N_16965,N_6635,N_5842);
or U16966 (N_16966,N_2321,N_5229);
nor U16967 (N_16967,N_4419,N_9355);
nand U16968 (N_16968,N_4654,N_4414);
xor U16969 (N_16969,N_5243,N_6404);
nor U16970 (N_16970,N_5249,N_9612);
nand U16971 (N_16971,N_6319,N_7874);
or U16972 (N_16972,N_8612,N_1202);
nand U16973 (N_16973,N_7117,N_9023);
or U16974 (N_16974,N_4871,N_4890);
or U16975 (N_16975,N_2703,N_3118);
xnor U16976 (N_16976,N_567,N_2572);
and U16977 (N_16977,N_1116,N_7254);
nor U16978 (N_16978,N_5243,N_9781);
or U16979 (N_16979,N_215,N_7452);
xor U16980 (N_16980,N_558,N_2695);
or U16981 (N_16981,N_7314,N_1308);
or U16982 (N_16982,N_7237,N_1319);
nand U16983 (N_16983,N_9517,N_1721);
nand U16984 (N_16984,N_5005,N_5580);
nand U16985 (N_16985,N_7605,N_7099);
or U16986 (N_16986,N_8215,N_1888);
nor U16987 (N_16987,N_6964,N_7213);
or U16988 (N_16988,N_5000,N_6861);
xnor U16989 (N_16989,N_912,N_8926);
xnor U16990 (N_16990,N_7654,N_6928);
xnor U16991 (N_16991,N_4393,N_437);
or U16992 (N_16992,N_7534,N_6989);
or U16993 (N_16993,N_7714,N_5362);
or U16994 (N_16994,N_3566,N_3503);
nor U16995 (N_16995,N_7185,N_9297);
and U16996 (N_16996,N_2349,N_590);
nand U16997 (N_16997,N_9900,N_8939);
or U16998 (N_16998,N_6347,N_8995);
nand U16999 (N_16999,N_7790,N_9960);
and U17000 (N_17000,N_7320,N_4788);
or U17001 (N_17001,N_1188,N_7857);
nor U17002 (N_17002,N_6317,N_3161);
nor U17003 (N_17003,N_1887,N_6154);
xor U17004 (N_17004,N_4382,N_2740);
and U17005 (N_17005,N_4412,N_7730);
xor U17006 (N_17006,N_8501,N_2133);
nand U17007 (N_17007,N_8461,N_8161);
or U17008 (N_17008,N_8651,N_6702);
nor U17009 (N_17009,N_1156,N_1505);
and U17010 (N_17010,N_2730,N_1517);
nor U17011 (N_17011,N_1473,N_6136);
or U17012 (N_17012,N_7686,N_8567);
nand U17013 (N_17013,N_9314,N_652);
nand U17014 (N_17014,N_6268,N_742);
nor U17015 (N_17015,N_6928,N_6122);
nand U17016 (N_17016,N_1010,N_7135);
and U17017 (N_17017,N_1232,N_5806);
nor U17018 (N_17018,N_9526,N_760);
and U17019 (N_17019,N_4324,N_8983);
xnor U17020 (N_17020,N_5646,N_7539);
xor U17021 (N_17021,N_8740,N_8781);
xnor U17022 (N_17022,N_6129,N_2387);
or U17023 (N_17023,N_2203,N_3062);
and U17024 (N_17024,N_7049,N_5011);
xnor U17025 (N_17025,N_311,N_5908);
and U17026 (N_17026,N_7605,N_686);
and U17027 (N_17027,N_7373,N_8718);
nor U17028 (N_17028,N_7993,N_2918);
and U17029 (N_17029,N_9303,N_909);
nor U17030 (N_17030,N_3380,N_3447);
or U17031 (N_17031,N_5322,N_6468);
nor U17032 (N_17032,N_3690,N_7135);
xnor U17033 (N_17033,N_9535,N_7516);
nand U17034 (N_17034,N_7229,N_6554);
xnor U17035 (N_17035,N_9334,N_2365);
and U17036 (N_17036,N_1555,N_6642);
or U17037 (N_17037,N_3422,N_7512);
nand U17038 (N_17038,N_8270,N_885);
xor U17039 (N_17039,N_6714,N_7184);
and U17040 (N_17040,N_7218,N_605);
or U17041 (N_17041,N_2583,N_2191);
and U17042 (N_17042,N_4364,N_7295);
nor U17043 (N_17043,N_9856,N_6629);
nand U17044 (N_17044,N_3085,N_9991);
and U17045 (N_17045,N_2615,N_6720);
xnor U17046 (N_17046,N_790,N_4943);
xor U17047 (N_17047,N_3190,N_3932);
nor U17048 (N_17048,N_7325,N_6464);
nand U17049 (N_17049,N_1821,N_9832);
nand U17050 (N_17050,N_6264,N_9194);
nand U17051 (N_17051,N_1148,N_1098);
nor U17052 (N_17052,N_3291,N_3014);
nor U17053 (N_17053,N_691,N_227);
and U17054 (N_17054,N_7838,N_7623);
or U17055 (N_17055,N_1098,N_3375);
and U17056 (N_17056,N_6439,N_582);
or U17057 (N_17057,N_6471,N_1382);
or U17058 (N_17058,N_4622,N_9240);
nand U17059 (N_17059,N_6494,N_2461);
or U17060 (N_17060,N_6227,N_7890);
xor U17061 (N_17061,N_4043,N_2908);
and U17062 (N_17062,N_5206,N_5713);
and U17063 (N_17063,N_2894,N_7613);
xor U17064 (N_17064,N_7481,N_5658);
nor U17065 (N_17065,N_6617,N_4246);
or U17066 (N_17066,N_9532,N_3386);
and U17067 (N_17067,N_7265,N_4114);
nand U17068 (N_17068,N_5692,N_9673);
nor U17069 (N_17069,N_6088,N_9065);
xnor U17070 (N_17070,N_5671,N_4917);
or U17071 (N_17071,N_3626,N_1035);
or U17072 (N_17072,N_5640,N_2707);
and U17073 (N_17073,N_1018,N_3455);
nor U17074 (N_17074,N_8260,N_5630);
or U17075 (N_17075,N_9284,N_9602);
xor U17076 (N_17076,N_1406,N_8674);
xnor U17077 (N_17077,N_475,N_4610);
and U17078 (N_17078,N_1767,N_9580);
nand U17079 (N_17079,N_2252,N_7198);
nor U17080 (N_17080,N_9196,N_9297);
nand U17081 (N_17081,N_4410,N_9871);
and U17082 (N_17082,N_8626,N_2070);
xor U17083 (N_17083,N_2100,N_5566);
and U17084 (N_17084,N_4532,N_2313);
and U17085 (N_17085,N_6990,N_810);
nand U17086 (N_17086,N_7139,N_3521);
nand U17087 (N_17087,N_2224,N_9953);
nor U17088 (N_17088,N_2830,N_2034);
xnor U17089 (N_17089,N_4010,N_8220);
xor U17090 (N_17090,N_4160,N_1880);
nor U17091 (N_17091,N_995,N_3353);
nor U17092 (N_17092,N_2789,N_8951);
xnor U17093 (N_17093,N_7829,N_7172);
nand U17094 (N_17094,N_7916,N_4358);
nor U17095 (N_17095,N_3562,N_2093);
nor U17096 (N_17096,N_2794,N_9858);
nand U17097 (N_17097,N_5343,N_2768);
nand U17098 (N_17098,N_6431,N_7011);
nand U17099 (N_17099,N_9212,N_1511);
nand U17100 (N_17100,N_1762,N_9722);
nand U17101 (N_17101,N_4261,N_852);
and U17102 (N_17102,N_1713,N_2838);
and U17103 (N_17103,N_3502,N_3348);
nand U17104 (N_17104,N_59,N_177);
xor U17105 (N_17105,N_7657,N_2551);
nand U17106 (N_17106,N_1729,N_3581);
nand U17107 (N_17107,N_6257,N_8560);
xnor U17108 (N_17108,N_7130,N_2707);
nor U17109 (N_17109,N_5725,N_537);
or U17110 (N_17110,N_8998,N_5383);
nand U17111 (N_17111,N_3810,N_3564);
xor U17112 (N_17112,N_2608,N_8480);
or U17113 (N_17113,N_4103,N_2118);
nand U17114 (N_17114,N_2601,N_8957);
or U17115 (N_17115,N_6339,N_7232);
xnor U17116 (N_17116,N_3471,N_7569);
xnor U17117 (N_17117,N_1676,N_1241);
xor U17118 (N_17118,N_3295,N_5725);
xor U17119 (N_17119,N_1474,N_594);
xor U17120 (N_17120,N_8251,N_6809);
nor U17121 (N_17121,N_8299,N_5743);
or U17122 (N_17122,N_9859,N_3602);
nand U17123 (N_17123,N_7369,N_5068);
xor U17124 (N_17124,N_3309,N_3215);
and U17125 (N_17125,N_6026,N_102);
or U17126 (N_17126,N_4466,N_1940);
nor U17127 (N_17127,N_5173,N_8689);
or U17128 (N_17128,N_5152,N_9835);
and U17129 (N_17129,N_7513,N_6352);
and U17130 (N_17130,N_7049,N_4437);
and U17131 (N_17131,N_3108,N_3074);
xor U17132 (N_17132,N_5168,N_888);
nor U17133 (N_17133,N_9003,N_3115);
nor U17134 (N_17134,N_4416,N_3194);
nand U17135 (N_17135,N_9000,N_4158);
and U17136 (N_17136,N_1967,N_6740);
xor U17137 (N_17137,N_8709,N_2978);
nand U17138 (N_17138,N_1854,N_3562);
xor U17139 (N_17139,N_7986,N_6216);
nand U17140 (N_17140,N_3412,N_9866);
xnor U17141 (N_17141,N_3975,N_318);
xor U17142 (N_17142,N_4076,N_919);
nor U17143 (N_17143,N_6544,N_9685);
xnor U17144 (N_17144,N_1916,N_2320);
nand U17145 (N_17145,N_3007,N_4200);
nand U17146 (N_17146,N_3214,N_6678);
nor U17147 (N_17147,N_4123,N_1788);
xor U17148 (N_17148,N_7519,N_3210);
or U17149 (N_17149,N_5286,N_6245);
and U17150 (N_17150,N_9731,N_3541);
nand U17151 (N_17151,N_47,N_8975);
xor U17152 (N_17152,N_4065,N_126);
nor U17153 (N_17153,N_590,N_9306);
xor U17154 (N_17154,N_1543,N_3771);
nor U17155 (N_17155,N_6989,N_8923);
nor U17156 (N_17156,N_2598,N_4332);
or U17157 (N_17157,N_7696,N_2496);
nand U17158 (N_17158,N_5467,N_7008);
or U17159 (N_17159,N_3412,N_5557);
xnor U17160 (N_17160,N_5796,N_2988);
or U17161 (N_17161,N_3415,N_6407);
or U17162 (N_17162,N_9207,N_9734);
xor U17163 (N_17163,N_685,N_5383);
and U17164 (N_17164,N_197,N_103);
xnor U17165 (N_17165,N_5464,N_52);
or U17166 (N_17166,N_5652,N_5313);
and U17167 (N_17167,N_1543,N_129);
nand U17168 (N_17168,N_8222,N_559);
nor U17169 (N_17169,N_6663,N_401);
nor U17170 (N_17170,N_5144,N_5212);
or U17171 (N_17171,N_6820,N_2364);
or U17172 (N_17172,N_171,N_161);
nor U17173 (N_17173,N_8406,N_2684);
xnor U17174 (N_17174,N_6483,N_6358);
nand U17175 (N_17175,N_5254,N_4339);
nor U17176 (N_17176,N_466,N_8879);
xor U17177 (N_17177,N_905,N_9090);
and U17178 (N_17178,N_7132,N_1784);
xnor U17179 (N_17179,N_5326,N_4801);
nand U17180 (N_17180,N_5633,N_9409);
and U17181 (N_17181,N_4393,N_4253);
or U17182 (N_17182,N_4013,N_205);
nor U17183 (N_17183,N_8137,N_9338);
nor U17184 (N_17184,N_1631,N_235);
nor U17185 (N_17185,N_773,N_644);
or U17186 (N_17186,N_1183,N_2628);
xor U17187 (N_17187,N_4836,N_4520);
xor U17188 (N_17188,N_8388,N_3905);
xnor U17189 (N_17189,N_2131,N_9597);
nor U17190 (N_17190,N_9336,N_7713);
nor U17191 (N_17191,N_2273,N_206);
and U17192 (N_17192,N_4775,N_2622);
nor U17193 (N_17193,N_9849,N_6413);
or U17194 (N_17194,N_6615,N_3592);
nand U17195 (N_17195,N_1255,N_9330);
nor U17196 (N_17196,N_8154,N_7773);
xor U17197 (N_17197,N_9498,N_3327);
xnor U17198 (N_17198,N_499,N_8719);
nand U17199 (N_17199,N_485,N_2721);
nor U17200 (N_17200,N_411,N_1915);
xnor U17201 (N_17201,N_2629,N_2586);
and U17202 (N_17202,N_9111,N_1479);
xnor U17203 (N_17203,N_5071,N_1205);
and U17204 (N_17204,N_8022,N_4878);
nor U17205 (N_17205,N_7286,N_6994);
xnor U17206 (N_17206,N_6345,N_4014);
xor U17207 (N_17207,N_9364,N_419);
xnor U17208 (N_17208,N_9353,N_255);
xor U17209 (N_17209,N_3064,N_881);
nor U17210 (N_17210,N_389,N_430);
nand U17211 (N_17211,N_5089,N_7774);
xor U17212 (N_17212,N_9703,N_7156);
nand U17213 (N_17213,N_4310,N_3357);
nand U17214 (N_17214,N_8193,N_5459);
or U17215 (N_17215,N_6302,N_4536);
nand U17216 (N_17216,N_834,N_2758);
and U17217 (N_17217,N_5033,N_2724);
and U17218 (N_17218,N_9269,N_2211);
nand U17219 (N_17219,N_251,N_1454);
xnor U17220 (N_17220,N_8653,N_9035);
or U17221 (N_17221,N_1474,N_2091);
nor U17222 (N_17222,N_9306,N_2653);
nor U17223 (N_17223,N_6941,N_5173);
or U17224 (N_17224,N_6633,N_4713);
xnor U17225 (N_17225,N_4952,N_2394);
or U17226 (N_17226,N_6341,N_1520);
xor U17227 (N_17227,N_52,N_3357);
xor U17228 (N_17228,N_6509,N_784);
and U17229 (N_17229,N_9800,N_3423);
or U17230 (N_17230,N_6538,N_8991);
nor U17231 (N_17231,N_6234,N_2748);
or U17232 (N_17232,N_7003,N_6736);
or U17233 (N_17233,N_3016,N_6483);
xnor U17234 (N_17234,N_186,N_9057);
nor U17235 (N_17235,N_2979,N_6491);
nor U17236 (N_17236,N_2329,N_8908);
nor U17237 (N_17237,N_7521,N_7632);
nand U17238 (N_17238,N_9834,N_939);
nand U17239 (N_17239,N_1436,N_6378);
or U17240 (N_17240,N_5716,N_13);
or U17241 (N_17241,N_9831,N_9528);
nand U17242 (N_17242,N_5298,N_4385);
xor U17243 (N_17243,N_4560,N_564);
nor U17244 (N_17244,N_7611,N_9076);
xor U17245 (N_17245,N_4422,N_916);
nor U17246 (N_17246,N_9218,N_5752);
nor U17247 (N_17247,N_1647,N_11);
xor U17248 (N_17248,N_1636,N_354);
nor U17249 (N_17249,N_5311,N_7413);
nor U17250 (N_17250,N_1571,N_8845);
and U17251 (N_17251,N_1679,N_3328);
xor U17252 (N_17252,N_5003,N_7056);
nand U17253 (N_17253,N_4777,N_8049);
and U17254 (N_17254,N_1828,N_802);
and U17255 (N_17255,N_5424,N_4701);
xnor U17256 (N_17256,N_7261,N_1328);
nand U17257 (N_17257,N_1988,N_1524);
nor U17258 (N_17258,N_5678,N_5039);
nand U17259 (N_17259,N_1970,N_8053);
and U17260 (N_17260,N_3590,N_7607);
or U17261 (N_17261,N_5538,N_7444);
nor U17262 (N_17262,N_6322,N_689);
nand U17263 (N_17263,N_9971,N_4003);
nor U17264 (N_17264,N_9642,N_5424);
nand U17265 (N_17265,N_4561,N_8972);
xnor U17266 (N_17266,N_875,N_4176);
or U17267 (N_17267,N_9101,N_5222);
nor U17268 (N_17268,N_4661,N_5759);
or U17269 (N_17269,N_1616,N_8156);
nor U17270 (N_17270,N_8586,N_4461);
nor U17271 (N_17271,N_8308,N_7675);
nand U17272 (N_17272,N_9501,N_8593);
and U17273 (N_17273,N_2342,N_6997);
nor U17274 (N_17274,N_4748,N_2469);
xor U17275 (N_17275,N_4716,N_2217);
xor U17276 (N_17276,N_1819,N_1789);
xnor U17277 (N_17277,N_1053,N_5731);
and U17278 (N_17278,N_3897,N_8839);
xor U17279 (N_17279,N_5117,N_4994);
nand U17280 (N_17280,N_4745,N_3651);
nor U17281 (N_17281,N_2537,N_4269);
nand U17282 (N_17282,N_8493,N_7857);
or U17283 (N_17283,N_3745,N_1612);
nand U17284 (N_17284,N_106,N_8506);
xor U17285 (N_17285,N_2597,N_3014);
xnor U17286 (N_17286,N_4539,N_1852);
nor U17287 (N_17287,N_2585,N_2877);
or U17288 (N_17288,N_3794,N_4089);
and U17289 (N_17289,N_532,N_6171);
xor U17290 (N_17290,N_2372,N_83);
nor U17291 (N_17291,N_29,N_3226);
xnor U17292 (N_17292,N_5225,N_5701);
nor U17293 (N_17293,N_7319,N_9604);
nand U17294 (N_17294,N_6645,N_4449);
and U17295 (N_17295,N_9969,N_4063);
xnor U17296 (N_17296,N_5182,N_612);
and U17297 (N_17297,N_2734,N_6478);
or U17298 (N_17298,N_2709,N_6147);
or U17299 (N_17299,N_9067,N_8111);
or U17300 (N_17300,N_8954,N_7921);
or U17301 (N_17301,N_1989,N_6968);
nor U17302 (N_17302,N_7521,N_6427);
nor U17303 (N_17303,N_8990,N_6331);
nor U17304 (N_17304,N_211,N_2390);
xnor U17305 (N_17305,N_5143,N_9868);
xnor U17306 (N_17306,N_133,N_9784);
and U17307 (N_17307,N_3486,N_8570);
and U17308 (N_17308,N_4434,N_8521);
xnor U17309 (N_17309,N_7936,N_4122);
or U17310 (N_17310,N_5113,N_722);
and U17311 (N_17311,N_3372,N_7841);
nand U17312 (N_17312,N_6981,N_3105);
xor U17313 (N_17313,N_1043,N_6673);
nor U17314 (N_17314,N_8291,N_7116);
nor U17315 (N_17315,N_6517,N_4043);
or U17316 (N_17316,N_7702,N_540);
and U17317 (N_17317,N_5898,N_5216);
and U17318 (N_17318,N_6781,N_9574);
nand U17319 (N_17319,N_1476,N_7076);
nand U17320 (N_17320,N_7402,N_7453);
and U17321 (N_17321,N_6799,N_7372);
nand U17322 (N_17322,N_5338,N_7517);
and U17323 (N_17323,N_5258,N_2730);
or U17324 (N_17324,N_5328,N_8978);
nand U17325 (N_17325,N_8384,N_1554);
or U17326 (N_17326,N_351,N_953);
xnor U17327 (N_17327,N_8777,N_9093);
or U17328 (N_17328,N_5383,N_2606);
nor U17329 (N_17329,N_1565,N_5279);
xor U17330 (N_17330,N_493,N_1333);
and U17331 (N_17331,N_1603,N_280);
xnor U17332 (N_17332,N_2102,N_6897);
nand U17333 (N_17333,N_4773,N_7743);
xor U17334 (N_17334,N_1553,N_4635);
and U17335 (N_17335,N_6441,N_455);
nor U17336 (N_17336,N_7637,N_7566);
nand U17337 (N_17337,N_5608,N_60);
nor U17338 (N_17338,N_1607,N_9148);
nor U17339 (N_17339,N_4890,N_6583);
or U17340 (N_17340,N_1334,N_778);
or U17341 (N_17341,N_267,N_1175);
nor U17342 (N_17342,N_9558,N_9050);
and U17343 (N_17343,N_4909,N_904);
and U17344 (N_17344,N_3010,N_296);
and U17345 (N_17345,N_7466,N_5382);
or U17346 (N_17346,N_8595,N_5234);
nand U17347 (N_17347,N_6455,N_3594);
or U17348 (N_17348,N_6701,N_5189);
or U17349 (N_17349,N_4667,N_3976);
or U17350 (N_17350,N_8591,N_4800);
nor U17351 (N_17351,N_9351,N_5491);
nand U17352 (N_17352,N_5648,N_6064);
xor U17353 (N_17353,N_5770,N_6515);
nand U17354 (N_17354,N_899,N_8946);
and U17355 (N_17355,N_9073,N_546);
nand U17356 (N_17356,N_7971,N_4048);
nand U17357 (N_17357,N_6274,N_9417);
nand U17358 (N_17358,N_6777,N_7801);
xnor U17359 (N_17359,N_93,N_2596);
nor U17360 (N_17360,N_6893,N_7860);
and U17361 (N_17361,N_371,N_6280);
nor U17362 (N_17362,N_8736,N_9057);
and U17363 (N_17363,N_9393,N_7878);
xor U17364 (N_17364,N_5698,N_2696);
and U17365 (N_17365,N_6487,N_3741);
and U17366 (N_17366,N_8374,N_6371);
xnor U17367 (N_17367,N_2154,N_2329);
xor U17368 (N_17368,N_4683,N_3752);
nor U17369 (N_17369,N_6861,N_4363);
or U17370 (N_17370,N_5376,N_4777);
nand U17371 (N_17371,N_1395,N_9521);
nand U17372 (N_17372,N_7076,N_7440);
nand U17373 (N_17373,N_9611,N_3127);
nor U17374 (N_17374,N_6369,N_3202);
and U17375 (N_17375,N_5359,N_8799);
and U17376 (N_17376,N_5210,N_379);
and U17377 (N_17377,N_8813,N_1234);
nand U17378 (N_17378,N_3220,N_61);
and U17379 (N_17379,N_1776,N_8495);
and U17380 (N_17380,N_1772,N_8523);
or U17381 (N_17381,N_268,N_2358);
xor U17382 (N_17382,N_2091,N_8391);
and U17383 (N_17383,N_7677,N_2245);
xor U17384 (N_17384,N_228,N_8368);
nand U17385 (N_17385,N_4064,N_5417);
nor U17386 (N_17386,N_4412,N_2946);
xnor U17387 (N_17387,N_986,N_1728);
and U17388 (N_17388,N_462,N_4549);
nor U17389 (N_17389,N_3459,N_8115);
and U17390 (N_17390,N_8268,N_1327);
and U17391 (N_17391,N_7643,N_3835);
xnor U17392 (N_17392,N_721,N_1902);
nor U17393 (N_17393,N_2936,N_8405);
or U17394 (N_17394,N_751,N_4045);
xnor U17395 (N_17395,N_4499,N_1921);
xnor U17396 (N_17396,N_2831,N_2460);
nor U17397 (N_17397,N_7382,N_5575);
and U17398 (N_17398,N_7861,N_1986);
and U17399 (N_17399,N_2347,N_3516);
nand U17400 (N_17400,N_442,N_4817);
or U17401 (N_17401,N_1833,N_7020);
and U17402 (N_17402,N_8600,N_1448);
or U17403 (N_17403,N_5080,N_1599);
or U17404 (N_17404,N_5193,N_6807);
nand U17405 (N_17405,N_4502,N_9833);
xnor U17406 (N_17406,N_6023,N_3651);
or U17407 (N_17407,N_8934,N_5179);
and U17408 (N_17408,N_3138,N_7958);
xnor U17409 (N_17409,N_3633,N_4903);
nor U17410 (N_17410,N_5855,N_8019);
xnor U17411 (N_17411,N_7421,N_3979);
nand U17412 (N_17412,N_7258,N_7378);
nor U17413 (N_17413,N_9971,N_796);
nor U17414 (N_17414,N_3281,N_2836);
xnor U17415 (N_17415,N_1339,N_1057);
and U17416 (N_17416,N_4328,N_8234);
or U17417 (N_17417,N_8692,N_4636);
nand U17418 (N_17418,N_700,N_4233);
nand U17419 (N_17419,N_4736,N_268);
nand U17420 (N_17420,N_9697,N_7321);
nand U17421 (N_17421,N_4607,N_2807);
nand U17422 (N_17422,N_7324,N_4803);
nor U17423 (N_17423,N_9922,N_4124);
and U17424 (N_17424,N_2149,N_5177);
and U17425 (N_17425,N_5222,N_7876);
xnor U17426 (N_17426,N_6117,N_1841);
or U17427 (N_17427,N_5160,N_5346);
nand U17428 (N_17428,N_6831,N_2735);
or U17429 (N_17429,N_6436,N_5525);
or U17430 (N_17430,N_104,N_8420);
and U17431 (N_17431,N_5231,N_6590);
xnor U17432 (N_17432,N_2245,N_2653);
nand U17433 (N_17433,N_9758,N_5226);
xnor U17434 (N_17434,N_7661,N_2893);
and U17435 (N_17435,N_2139,N_5101);
nand U17436 (N_17436,N_9703,N_1116);
and U17437 (N_17437,N_3408,N_6858);
xor U17438 (N_17438,N_8626,N_7469);
nand U17439 (N_17439,N_7875,N_5576);
and U17440 (N_17440,N_9167,N_7034);
xnor U17441 (N_17441,N_427,N_9834);
xor U17442 (N_17442,N_9522,N_2414);
nand U17443 (N_17443,N_7859,N_372);
nor U17444 (N_17444,N_3356,N_2184);
nand U17445 (N_17445,N_6090,N_1723);
xnor U17446 (N_17446,N_314,N_105);
or U17447 (N_17447,N_9148,N_8605);
nor U17448 (N_17448,N_9767,N_1900);
nor U17449 (N_17449,N_383,N_8280);
xnor U17450 (N_17450,N_322,N_4039);
or U17451 (N_17451,N_7977,N_6030);
xor U17452 (N_17452,N_5184,N_7619);
nor U17453 (N_17453,N_4064,N_2902);
nor U17454 (N_17454,N_2101,N_4266);
and U17455 (N_17455,N_527,N_802);
and U17456 (N_17456,N_1004,N_7587);
nand U17457 (N_17457,N_159,N_8184);
or U17458 (N_17458,N_1083,N_8635);
or U17459 (N_17459,N_4222,N_4698);
nand U17460 (N_17460,N_7246,N_9985);
nand U17461 (N_17461,N_1803,N_6099);
xnor U17462 (N_17462,N_8516,N_5629);
nor U17463 (N_17463,N_1675,N_6183);
xor U17464 (N_17464,N_4352,N_6439);
xnor U17465 (N_17465,N_272,N_2101);
or U17466 (N_17466,N_620,N_3169);
or U17467 (N_17467,N_140,N_2855);
xor U17468 (N_17468,N_4875,N_6361);
nand U17469 (N_17469,N_212,N_7176);
nor U17470 (N_17470,N_244,N_1410);
and U17471 (N_17471,N_2481,N_3132);
nor U17472 (N_17472,N_2829,N_4492);
nand U17473 (N_17473,N_8165,N_8607);
and U17474 (N_17474,N_2448,N_2806);
and U17475 (N_17475,N_6180,N_8309);
nor U17476 (N_17476,N_9723,N_3038);
and U17477 (N_17477,N_102,N_9103);
or U17478 (N_17478,N_5103,N_8461);
and U17479 (N_17479,N_6492,N_7696);
or U17480 (N_17480,N_4086,N_3359);
xor U17481 (N_17481,N_7483,N_7492);
xnor U17482 (N_17482,N_3011,N_6210);
or U17483 (N_17483,N_7601,N_2281);
nor U17484 (N_17484,N_8407,N_6888);
and U17485 (N_17485,N_5542,N_1098);
and U17486 (N_17486,N_2151,N_4026);
and U17487 (N_17487,N_8757,N_8879);
nor U17488 (N_17488,N_7027,N_8223);
xnor U17489 (N_17489,N_7156,N_9543);
and U17490 (N_17490,N_5159,N_5594);
or U17491 (N_17491,N_3352,N_3953);
and U17492 (N_17492,N_3495,N_3133);
nand U17493 (N_17493,N_5101,N_6788);
xnor U17494 (N_17494,N_3655,N_9499);
nand U17495 (N_17495,N_685,N_6011);
xnor U17496 (N_17496,N_3549,N_6921);
xnor U17497 (N_17497,N_541,N_3745);
nor U17498 (N_17498,N_3276,N_1538);
xnor U17499 (N_17499,N_4285,N_2113);
xnor U17500 (N_17500,N_3704,N_1796);
nand U17501 (N_17501,N_3709,N_6691);
nor U17502 (N_17502,N_2285,N_8604);
nor U17503 (N_17503,N_6094,N_6826);
and U17504 (N_17504,N_6118,N_4626);
and U17505 (N_17505,N_5254,N_984);
or U17506 (N_17506,N_2596,N_3872);
xor U17507 (N_17507,N_7527,N_1365);
nand U17508 (N_17508,N_1815,N_8637);
nand U17509 (N_17509,N_7311,N_6711);
or U17510 (N_17510,N_2764,N_7180);
and U17511 (N_17511,N_8630,N_534);
or U17512 (N_17512,N_4106,N_4968);
xor U17513 (N_17513,N_7325,N_2847);
nand U17514 (N_17514,N_322,N_8396);
and U17515 (N_17515,N_4068,N_5785);
xor U17516 (N_17516,N_1876,N_1163);
xor U17517 (N_17517,N_8439,N_801);
nor U17518 (N_17518,N_6820,N_3328);
nor U17519 (N_17519,N_3810,N_7979);
xnor U17520 (N_17520,N_9329,N_2197);
nor U17521 (N_17521,N_6245,N_4982);
nor U17522 (N_17522,N_5570,N_1342);
or U17523 (N_17523,N_1414,N_6159);
and U17524 (N_17524,N_461,N_3091);
or U17525 (N_17525,N_7808,N_3864);
or U17526 (N_17526,N_2228,N_463);
nand U17527 (N_17527,N_543,N_5134);
and U17528 (N_17528,N_626,N_4692);
or U17529 (N_17529,N_5414,N_5687);
and U17530 (N_17530,N_382,N_8788);
nand U17531 (N_17531,N_9425,N_7860);
nor U17532 (N_17532,N_3646,N_1214);
nor U17533 (N_17533,N_8538,N_2669);
xnor U17534 (N_17534,N_6676,N_5561);
or U17535 (N_17535,N_9362,N_3131);
nand U17536 (N_17536,N_2122,N_322);
or U17537 (N_17537,N_5573,N_6971);
nand U17538 (N_17538,N_6638,N_163);
nor U17539 (N_17539,N_9689,N_6220);
or U17540 (N_17540,N_627,N_4359);
and U17541 (N_17541,N_5107,N_4892);
and U17542 (N_17542,N_2117,N_3583);
xor U17543 (N_17543,N_6538,N_2892);
xnor U17544 (N_17544,N_4226,N_5294);
or U17545 (N_17545,N_5967,N_4755);
or U17546 (N_17546,N_3412,N_9381);
and U17547 (N_17547,N_5672,N_8305);
nand U17548 (N_17548,N_6735,N_2554);
nor U17549 (N_17549,N_8944,N_2205);
or U17550 (N_17550,N_4014,N_9626);
nand U17551 (N_17551,N_2548,N_3010);
nand U17552 (N_17552,N_1529,N_2433);
and U17553 (N_17553,N_2554,N_3971);
nand U17554 (N_17554,N_9114,N_3890);
or U17555 (N_17555,N_8128,N_9979);
xnor U17556 (N_17556,N_1867,N_9056);
xnor U17557 (N_17557,N_1181,N_1932);
and U17558 (N_17558,N_6116,N_9695);
nand U17559 (N_17559,N_1638,N_3379);
nand U17560 (N_17560,N_7291,N_2544);
nand U17561 (N_17561,N_8558,N_6004);
and U17562 (N_17562,N_8352,N_6624);
or U17563 (N_17563,N_9190,N_5784);
or U17564 (N_17564,N_1026,N_218);
xnor U17565 (N_17565,N_3842,N_4663);
nand U17566 (N_17566,N_8834,N_4264);
nor U17567 (N_17567,N_8283,N_8979);
nor U17568 (N_17568,N_3285,N_3156);
xor U17569 (N_17569,N_2495,N_9910);
nor U17570 (N_17570,N_3382,N_810);
nand U17571 (N_17571,N_2348,N_3926);
nor U17572 (N_17572,N_5491,N_1875);
nand U17573 (N_17573,N_8025,N_971);
and U17574 (N_17574,N_9285,N_3576);
or U17575 (N_17575,N_4920,N_4998);
or U17576 (N_17576,N_3054,N_7322);
xnor U17577 (N_17577,N_6234,N_3057);
xor U17578 (N_17578,N_4256,N_2150);
and U17579 (N_17579,N_5537,N_3418);
or U17580 (N_17580,N_6083,N_9233);
nor U17581 (N_17581,N_354,N_4583);
nor U17582 (N_17582,N_2962,N_7797);
xor U17583 (N_17583,N_8510,N_9654);
nor U17584 (N_17584,N_3915,N_3268);
nor U17585 (N_17585,N_7619,N_1445);
nand U17586 (N_17586,N_1133,N_7848);
xor U17587 (N_17587,N_6866,N_7910);
nor U17588 (N_17588,N_4663,N_5825);
or U17589 (N_17589,N_9108,N_4959);
and U17590 (N_17590,N_2579,N_8124);
nor U17591 (N_17591,N_4101,N_2252);
nand U17592 (N_17592,N_2583,N_3556);
and U17593 (N_17593,N_5232,N_4986);
xor U17594 (N_17594,N_2523,N_7190);
nand U17595 (N_17595,N_954,N_9392);
nand U17596 (N_17596,N_6324,N_9539);
nand U17597 (N_17597,N_6351,N_7220);
xnor U17598 (N_17598,N_1520,N_5086);
nand U17599 (N_17599,N_744,N_216);
and U17600 (N_17600,N_21,N_4650);
xnor U17601 (N_17601,N_5144,N_4450);
nor U17602 (N_17602,N_3175,N_9254);
and U17603 (N_17603,N_4417,N_912);
or U17604 (N_17604,N_7278,N_2380);
nand U17605 (N_17605,N_7395,N_6577);
nor U17606 (N_17606,N_2840,N_9695);
or U17607 (N_17607,N_1004,N_6078);
nor U17608 (N_17608,N_541,N_7885);
or U17609 (N_17609,N_6643,N_6768);
nand U17610 (N_17610,N_7672,N_4264);
or U17611 (N_17611,N_5053,N_317);
and U17612 (N_17612,N_8729,N_4341);
nand U17613 (N_17613,N_7740,N_9677);
and U17614 (N_17614,N_8821,N_3603);
xor U17615 (N_17615,N_7220,N_1355);
nand U17616 (N_17616,N_3160,N_9092);
or U17617 (N_17617,N_4067,N_2512);
nand U17618 (N_17618,N_6450,N_6799);
xor U17619 (N_17619,N_5879,N_5186);
and U17620 (N_17620,N_2183,N_1463);
or U17621 (N_17621,N_3469,N_8631);
xnor U17622 (N_17622,N_8088,N_5237);
or U17623 (N_17623,N_9333,N_3289);
nand U17624 (N_17624,N_9399,N_8360);
and U17625 (N_17625,N_3293,N_4404);
nor U17626 (N_17626,N_203,N_456);
nand U17627 (N_17627,N_8499,N_3481);
or U17628 (N_17628,N_337,N_2587);
nand U17629 (N_17629,N_5662,N_6802);
nor U17630 (N_17630,N_3774,N_8559);
and U17631 (N_17631,N_4829,N_2781);
nand U17632 (N_17632,N_270,N_2447);
nand U17633 (N_17633,N_3450,N_7323);
xor U17634 (N_17634,N_1817,N_9278);
and U17635 (N_17635,N_3840,N_6795);
and U17636 (N_17636,N_2312,N_4761);
and U17637 (N_17637,N_8160,N_1814);
or U17638 (N_17638,N_1113,N_4819);
nand U17639 (N_17639,N_9155,N_9599);
xor U17640 (N_17640,N_8616,N_9020);
nand U17641 (N_17641,N_4643,N_6761);
nand U17642 (N_17642,N_2083,N_3);
nor U17643 (N_17643,N_5190,N_2130);
xnor U17644 (N_17644,N_7214,N_4903);
and U17645 (N_17645,N_8779,N_8068);
and U17646 (N_17646,N_4689,N_3132);
nand U17647 (N_17647,N_2306,N_5533);
nand U17648 (N_17648,N_1044,N_6709);
nor U17649 (N_17649,N_7865,N_2890);
nor U17650 (N_17650,N_9766,N_9285);
nor U17651 (N_17651,N_4232,N_2141);
nand U17652 (N_17652,N_5257,N_2237);
or U17653 (N_17653,N_751,N_2253);
or U17654 (N_17654,N_8511,N_7117);
or U17655 (N_17655,N_6229,N_203);
and U17656 (N_17656,N_1008,N_1557);
nor U17657 (N_17657,N_6006,N_3208);
xor U17658 (N_17658,N_5040,N_5422);
and U17659 (N_17659,N_250,N_3351);
xnor U17660 (N_17660,N_8752,N_1014);
nor U17661 (N_17661,N_7488,N_7413);
xnor U17662 (N_17662,N_6084,N_3863);
or U17663 (N_17663,N_6858,N_6083);
or U17664 (N_17664,N_6325,N_1991);
nor U17665 (N_17665,N_2150,N_5148);
xnor U17666 (N_17666,N_147,N_3726);
xor U17667 (N_17667,N_8612,N_9359);
nand U17668 (N_17668,N_4130,N_4058);
or U17669 (N_17669,N_5666,N_9663);
nand U17670 (N_17670,N_9224,N_9775);
and U17671 (N_17671,N_1177,N_4480);
or U17672 (N_17672,N_4930,N_9321);
nor U17673 (N_17673,N_3037,N_6100);
and U17674 (N_17674,N_489,N_3068);
and U17675 (N_17675,N_8494,N_1061);
nand U17676 (N_17676,N_4532,N_4860);
xnor U17677 (N_17677,N_4893,N_9476);
xor U17678 (N_17678,N_1344,N_5541);
nand U17679 (N_17679,N_4097,N_9421);
nand U17680 (N_17680,N_6581,N_6482);
xor U17681 (N_17681,N_3149,N_1652);
and U17682 (N_17682,N_1352,N_4237);
nor U17683 (N_17683,N_4889,N_1644);
and U17684 (N_17684,N_3210,N_7813);
nor U17685 (N_17685,N_5075,N_596);
or U17686 (N_17686,N_3306,N_9925);
or U17687 (N_17687,N_2412,N_1835);
nor U17688 (N_17688,N_6876,N_5683);
nand U17689 (N_17689,N_1151,N_932);
or U17690 (N_17690,N_3795,N_2413);
nand U17691 (N_17691,N_7478,N_756);
nor U17692 (N_17692,N_9532,N_3258);
nand U17693 (N_17693,N_46,N_8158);
xor U17694 (N_17694,N_7967,N_59);
xor U17695 (N_17695,N_6181,N_7168);
xnor U17696 (N_17696,N_6216,N_325);
or U17697 (N_17697,N_791,N_5527);
nand U17698 (N_17698,N_9415,N_9450);
and U17699 (N_17699,N_9382,N_6665);
or U17700 (N_17700,N_4314,N_2807);
nor U17701 (N_17701,N_3409,N_7041);
or U17702 (N_17702,N_276,N_7462);
nand U17703 (N_17703,N_7576,N_2275);
and U17704 (N_17704,N_6662,N_4580);
xor U17705 (N_17705,N_5056,N_8282);
xor U17706 (N_17706,N_9335,N_1067);
or U17707 (N_17707,N_1615,N_6734);
xor U17708 (N_17708,N_4421,N_7968);
nand U17709 (N_17709,N_2510,N_4381);
nand U17710 (N_17710,N_9295,N_2225);
nor U17711 (N_17711,N_2209,N_8108);
nand U17712 (N_17712,N_7968,N_3893);
or U17713 (N_17713,N_9031,N_8432);
and U17714 (N_17714,N_7147,N_1203);
and U17715 (N_17715,N_8286,N_221);
and U17716 (N_17716,N_1864,N_2225);
nand U17717 (N_17717,N_8393,N_7331);
or U17718 (N_17718,N_4320,N_964);
nand U17719 (N_17719,N_5814,N_807);
or U17720 (N_17720,N_5049,N_9438);
nand U17721 (N_17721,N_1105,N_200);
and U17722 (N_17722,N_2599,N_3561);
xor U17723 (N_17723,N_9034,N_1768);
and U17724 (N_17724,N_2163,N_6059);
and U17725 (N_17725,N_9673,N_2090);
nor U17726 (N_17726,N_9697,N_8493);
and U17727 (N_17727,N_7013,N_1919);
and U17728 (N_17728,N_9579,N_1213);
nand U17729 (N_17729,N_6989,N_2341);
nand U17730 (N_17730,N_1585,N_4240);
or U17731 (N_17731,N_4609,N_1463);
nor U17732 (N_17732,N_5033,N_3516);
nor U17733 (N_17733,N_6053,N_1178);
or U17734 (N_17734,N_850,N_6754);
or U17735 (N_17735,N_2503,N_2817);
or U17736 (N_17736,N_6196,N_7210);
nand U17737 (N_17737,N_4985,N_4519);
or U17738 (N_17738,N_6913,N_2617);
xor U17739 (N_17739,N_8686,N_3469);
or U17740 (N_17740,N_4203,N_410);
xor U17741 (N_17741,N_881,N_2717);
xor U17742 (N_17742,N_8266,N_9753);
nand U17743 (N_17743,N_3379,N_3545);
nor U17744 (N_17744,N_4802,N_1954);
xor U17745 (N_17745,N_1203,N_4664);
and U17746 (N_17746,N_301,N_1182);
nand U17747 (N_17747,N_7560,N_4129);
nor U17748 (N_17748,N_9825,N_9912);
nor U17749 (N_17749,N_392,N_3293);
nor U17750 (N_17750,N_9242,N_7835);
and U17751 (N_17751,N_690,N_3413);
nor U17752 (N_17752,N_3198,N_5164);
xor U17753 (N_17753,N_5655,N_5921);
or U17754 (N_17754,N_1867,N_1656);
xor U17755 (N_17755,N_1005,N_6101);
nand U17756 (N_17756,N_9401,N_3865);
and U17757 (N_17757,N_5987,N_6461);
and U17758 (N_17758,N_5272,N_1386);
xor U17759 (N_17759,N_9898,N_1244);
or U17760 (N_17760,N_5551,N_5368);
nor U17761 (N_17761,N_3811,N_4019);
and U17762 (N_17762,N_4029,N_255);
or U17763 (N_17763,N_8041,N_6540);
and U17764 (N_17764,N_8203,N_1059);
nor U17765 (N_17765,N_1806,N_8002);
or U17766 (N_17766,N_2544,N_6578);
and U17767 (N_17767,N_181,N_2890);
and U17768 (N_17768,N_2675,N_8496);
xor U17769 (N_17769,N_7572,N_404);
xor U17770 (N_17770,N_1710,N_7367);
nor U17771 (N_17771,N_8502,N_3038);
and U17772 (N_17772,N_2572,N_6242);
nand U17773 (N_17773,N_136,N_5084);
xor U17774 (N_17774,N_1673,N_8876);
nor U17775 (N_17775,N_2674,N_78);
and U17776 (N_17776,N_9097,N_290);
xnor U17777 (N_17777,N_2959,N_5976);
nand U17778 (N_17778,N_8556,N_3407);
or U17779 (N_17779,N_4405,N_5086);
xor U17780 (N_17780,N_5250,N_9144);
xor U17781 (N_17781,N_5652,N_3733);
and U17782 (N_17782,N_4628,N_1401);
nor U17783 (N_17783,N_4184,N_3903);
nor U17784 (N_17784,N_4620,N_7137);
nor U17785 (N_17785,N_2885,N_9780);
and U17786 (N_17786,N_2934,N_6462);
and U17787 (N_17787,N_8827,N_3150);
and U17788 (N_17788,N_8599,N_7224);
nor U17789 (N_17789,N_5063,N_6723);
xor U17790 (N_17790,N_3776,N_4416);
xor U17791 (N_17791,N_4751,N_2892);
nand U17792 (N_17792,N_2495,N_5574);
or U17793 (N_17793,N_3160,N_6940);
or U17794 (N_17794,N_2930,N_6510);
xnor U17795 (N_17795,N_2441,N_3005);
or U17796 (N_17796,N_4933,N_3032);
nor U17797 (N_17797,N_2397,N_2754);
nor U17798 (N_17798,N_4780,N_6616);
and U17799 (N_17799,N_3881,N_5938);
xor U17800 (N_17800,N_8223,N_8134);
and U17801 (N_17801,N_5633,N_3510);
or U17802 (N_17802,N_7418,N_2841);
nand U17803 (N_17803,N_9731,N_9410);
nor U17804 (N_17804,N_101,N_1084);
nor U17805 (N_17805,N_909,N_488);
nand U17806 (N_17806,N_6738,N_5587);
xnor U17807 (N_17807,N_1125,N_9381);
nor U17808 (N_17808,N_5784,N_7352);
or U17809 (N_17809,N_19,N_4913);
xor U17810 (N_17810,N_8191,N_4742);
or U17811 (N_17811,N_362,N_8074);
or U17812 (N_17812,N_9035,N_1105);
nand U17813 (N_17813,N_4395,N_2133);
nor U17814 (N_17814,N_4490,N_6249);
and U17815 (N_17815,N_2456,N_5291);
or U17816 (N_17816,N_9919,N_652);
and U17817 (N_17817,N_6305,N_9530);
nand U17818 (N_17818,N_5808,N_1980);
and U17819 (N_17819,N_8283,N_9185);
or U17820 (N_17820,N_1743,N_9162);
xnor U17821 (N_17821,N_4527,N_2538);
and U17822 (N_17822,N_3826,N_5569);
xor U17823 (N_17823,N_9163,N_6879);
nand U17824 (N_17824,N_2306,N_4292);
or U17825 (N_17825,N_2633,N_4953);
nor U17826 (N_17826,N_1034,N_1510);
nor U17827 (N_17827,N_6369,N_2691);
nor U17828 (N_17828,N_2378,N_7710);
xnor U17829 (N_17829,N_6164,N_5968);
or U17830 (N_17830,N_6896,N_6371);
xnor U17831 (N_17831,N_3534,N_5558);
nand U17832 (N_17832,N_1048,N_8372);
nand U17833 (N_17833,N_7011,N_3897);
xnor U17834 (N_17834,N_1365,N_5331);
or U17835 (N_17835,N_3180,N_5471);
nand U17836 (N_17836,N_1425,N_9153);
or U17837 (N_17837,N_2778,N_8998);
and U17838 (N_17838,N_634,N_9877);
nor U17839 (N_17839,N_3490,N_8244);
or U17840 (N_17840,N_1742,N_9679);
or U17841 (N_17841,N_4867,N_7585);
nor U17842 (N_17842,N_3216,N_8168);
nor U17843 (N_17843,N_84,N_2942);
and U17844 (N_17844,N_5509,N_2615);
xor U17845 (N_17845,N_8870,N_3587);
nand U17846 (N_17846,N_7363,N_2172);
nand U17847 (N_17847,N_4848,N_9835);
or U17848 (N_17848,N_9766,N_5203);
nor U17849 (N_17849,N_6877,N_8287);
nor U17850 (N_17850,N_7070,N_815);
or U17851 (N_17851,N_1152,N_5817);
and U17852 (N_17852,N_9162,N_7932);
xor U17853 (N_17853,N_2891,N_9452);
nor U17854 (N_17854,N_8876,N_871);
or U17855 (N_17855,N_2097,N_8966);
or U17856 (N_17856,N_4899,N_9567);
and U17857 (N_17857,N_309,N_9813);
and U17858 (N_17858,N_9146,N_1921);
nand U17859 (N_17859,N_1916,N_2371);
nand U17860 (N_17860,N_3716,N_8924);
and U17861 (N_17861,N_9801,N_9644);
xor U17862 (N_17862,N_7951,N_6956);
nand U17863 (N_17863,N_4349,N_5283);
xor U17864 (N_17864,N_3540,N_2711);
xnor U17865 (N_17865,N_5184,N_5617);
xnor U17866 (N_17866,N_817,N_753);
and U17867 (N_17867,N_2139,N_4964);
xor U17868 (N_17868,N_5763,N_8296);
and U17869 (N_17869,N_4009,N_5836);
xor U17870 (N_17870,N_5694,N_5805);
nand U17871 (N_17871,N_8999,N_6601);
nor U17872 (N_17872,N_6691,N_5402);
nor U17873 (N_17873,N_6619,N_6131);
nor U17874 (N_17874,N_2890,N_739);
and U17875 (N_17875,N_7869,N_221);
nor U17876 (N_17876,N_5955,N_9922);
and U17877 (N_17877,N_3784,N_4787);
nor U17878 (N_17878,N_2100,N_3744);
and U17879 (N_17879,N_7610,N_2579);
and U17880 (N_17880,N_262,N_76);
xor U17881 (N_17881,N_614,N_455);
nor U17882 (N_17882,N_2060,N_5025);
xor U17883 (N_17883,N_3613,N_469);
or U17884 (N_17884,N_4767,N_676);
nor U17885 (N_17885,N_3068,N_9664);
and U17886 (N_17886,N_2984,N_3235);
nand U17887 (N_17887,N_577,N_4572);
xnor U17888 (N_17888,N_8424,N_9446);
and U17889 (N_17889,N_522,N_3730);
nand U17890 (N_17890,N_1045,N_2956);
xor U17891 (N_17891,N_3599,N_1671);
and U17892 (N_17892,N_3863,N_6940);
and U17893 (N_17893,N_1799,N_8029);
nand U17894 (N_17894,N_5324,N_9825);
nor U17895 (N_17895,N_5367,N_1204);
and U17896 (N_17896,N_1300,N_3776);
nand U17897 (N_17897,N_5793,N_3500);
nor U17898 (N_17898,N_5607,N_8031);
nor U17899 (N_17899,N_9406,N_1764);
xnor U17900 (N_17900,N_3808,N_8961);
xor U17901 (N_17901,N_4292,N_1139);
nand U17902 (N_17902,N_5574,N_1462);
nand U17903 (N_17903,N_455,N_9271);
nor U17904 (N_17904,N_1274,N_1877);
or U17905 (N_17905,N_231,N_3454);
and U17906 (N_17906,N_3203,N_7370);
xor U17907 (N_17907,N_2563,N_5019);
nor U17908 (N_17908,N_5739,N_1232);
or U17909 (N_17909,N_2544,N_2760);
nor U17910 (N_17910,N_4524,N_584);
xor U17911 (N_17911,N_1122,N_2943);
xnor U17912 (N_17912,N_1160,N_1891);
nand U17913 (N_17913,N_5515,N_2555);
nand U17914 (N_17914,N_8875,N_2948);
nand U17915 (N_17915,N_941,N_3084);
nand U17916 (N_17916,N_2242,N_971);
xnor U17917 (N_17917,N_1105,N_3132);
nor U17918 (N_17918,N_3794,N_1515);
nand U17919 (N_17919,N_4202,N_3487);
xnor U17920 (N_17920,N_9713,N_2578);
nand U17921 (N_17921,N_4515,N_5100);
nor U17922 (N_17922,N_3047,N_7653);
nor U17923 (N_17923,N_5470,N_4888);
nand U17924 (N_17924,N_9892,N_5317);
and U17925 (N_17925,N_7507,N_3130);
or U17926 (N_17926,N_7567,N_2458);
or U17927 (N_17927,N_4679,N_795);
nand U17928 (N_17928,N_5746,N_6785);
nor U17929 (N_17929,N_7207,N_8855);
xnor U17930 (N_17930,N_1220,N_9823);
nand U17931 (N_17931,N_7482,N_6071);
nand U17932 (N_17932,N_2183,N_2131);
nor U17933 (N_17933,N_7983,N_2686);
nand U17934 (N_17934,N_5209,N_1772);
or U17935 (N_17935,N_4564,N_1073);
nand U17936 (N_17936,N_5034,N_3844);
xor U17937 (N_17937,N_4674,N_2810);
nand U17938 (N_17938,N_5493,N_5289);
nor U17939 (N_17939,N_5080,N_8770);
nor U17940 (N_17940,N_4591,N_729);
and U17941 (N_17941,N_2578,N_4843);
and U17942 (N_17942,N_6333,N_4264);
and U17943 (N_17943,N_9249,N_9212);
or U17944 (N_17944,N_7269,N_187);
or U17945 (N_17945,N_2831,N_7162);
or U17946 (N_17946,N_6391,N_3198);
nand U17947 (N_17947,N_1797,N_2341);
nor U17948 (N_17948,N_4190,N_1979);
or U17949 (N_17949,N_4142,N_7900);
and U17950 (N_17950,N_8662,N_5804);
or U17951 (N_17951,N_1073,N_8110);
nand U17952 (N_17952,N_7800,N_7724);
nor U17953 (N_17953,N_1179,N_755);
xor U17954 (N_17954,N_9619,N_8305);
or U17955 (N_17955,N_4571,N_8606);
nor U17956 (N_17956,N_9020,N_2644);
nand U17957 (N_17957,N_6406,N_9895);
or U17958 (N_17958,N_3368,N_2869);
xnor U17959 (N_17959,N_6062,N_1418);
nand U17960 (N_17960,N_6343,N_455);
nand U17961 (N_17961,N_352,N_773);
nor U17962 (N_17962,N_2769,N_1622);
xnor U17963 (N_17963,N_731,N_7559);
nor U17964 (N_17964,N_1115,N_8183);
or U17965 (N_17965,N_9631,N_9018);
and U17966 (N_17966,N_1149,N_4666);
xnor U17967 (N_17967,N_7752,N_5778);
and U17968 (N_17968,N_9855,N_5302);
or U17969 (N_17969,N_3480,N_4072);
nand U17970 (N_17970,N_9149,N_1441);
nand U17971 (N_17971,N_5951,N_5622);
nand U17972 (N_17972,N_4662,N_4641);
xor U17973 (N_17973,N_3457,N_6613);
xnor U17974 (N_17974,N_3515,N_5463);
or U17975 (N_17975,N_1610,N_7198);
and U17976 (N_17976,N_1363,N_3106);
nor U17977 (N_17977,N_4436,N_7601);
and U17978 (N_17978,N_3185,N_6917);
or U17979 (N_17979,N_3996,N_1798);
nor U17980 (N_17980,N_5750,N_8489);
nand U17981 (N_17981,N_8706,N_6448);
nand U17982 (N_17982,N_4133,N_2333);
nor U17983 (N_17983,N_202,N_741);
nor U17984 (N_17984,N_1453,N_3896);
and U17985 (N_17985,N_167,N_9210);
xor U17986 (N_17986,N_1754,N_2338);
nor U17987 (N_17987,N_6348,N_3232);
nand U17988 (N_17988,N_1094,N_7360);
or U17989 (N_17989,N_4064,N_7213);
nor U17990 (N_17990,N_4569,N_3436);
or U17991 (N_17991,N_1518,N_5726);
nand U17992 (N_17992,N_1808,N_1316);
nor U17993 (N_17993,N_8492,N_7343);
or U17994 (N_17994,N_2641,N_4393);
or U17995 (N_17995,N_7445,N_7436);
nand U17996 (N_17996,N_2617,N_7968);
xor U17997 (N_17997,N_3667,N_5615);
nand U17998 (N_17998,N_6251,N_2672);
or U17999 (N_17999,N_5436,N_9043);
nor U18000 (N_18000,N_500,N_9859);
nand U18001 (N_18001,N_5466,N_6739);
and U18002 (N_18002,N_9489,N_6912);
nand U18003 (N_18003,N_4453,N_9236);
nor U18004 (N_18004,N_5322,N_5263);
and U18005 (N_18005,N_3506,N_4866);
or U18006 (N_18006,N_3538,N_6982);
and U18007 (N_18007,N_4480,N_5571);
or U18008 (N_18008,N_4155,N_3792);
nand U18009 (N_18009,N_928,N_2063);
xor U18010 (N_18010,N_6311,N_4111);
and U18011 (N_18011,N_8647,N_961);
and U18012 (N_18012,N_4699,N_4235);
nand U18013 (N_18013,N_5147,N_3803);
and U18014 (N_18014,N_1521,N_1222);
nor U18015 (N_18015,N_9464,N_5493);
and U18016 (N_18016,N_8984,N_7266);
xnor U18017 (N_18017,N_796,N_2059);
xor U18018 (N_18018,N_9815,N_4592);
nand U18019 (N_18019,N_647,N_6289);
or U18020 (N_18020,N_3557,N_8792);
or U18021 (N_18021,N_687,N_50);
or U18022 (N_18022,N_5532,N_5415);
nand U18023 (N_18023,N_7751,N_381);
xor U18024 (N_18024,N_539,N_4418);
xnor U18025 (N_18025,N_6354,N_2010);
nand U18026 (N_18026,N_4184,N_6736);
xor U18027 (N_18027,N_3109,N_1147);
nand U18028 (N_18028,N_7887,N_123);
and U18029 (N_18029,N_3157,N_5021);
nand U18030 (N_18030,N_2936,N_8182);
nor U18031 (N_18031,N_1916,N_1063);
and U18032 (N_18032,N_1918,N_5143);
xnor U18033 (N_18033,N_5498,N_420);
xor U18034 (N_18034,N_141,N_7199);
nand U18035 (N_18035,N_9238,N_4231);
nor U18036 (N_18036,N_8010,N_1964);
or U18037 (N_18037,N_7401,N_9719);
and U18038 (N_18038,N_7087,N_8543);
xor U18039 (N_18039,N_2010,N_2294);
nand U18040 (N_18040,N_5707,N_9032);
and U18041 (N_18041,N_3287,N_1911);
xor U18042 (N_18042,N_4632,N_5118);
and U18043 (N_18043,N_903,N_7348);
nand U18044 (N_18044,N_7919,N_5017);
nor U18045 (N_18045,N_4134,N_1073);
or U18046 (N_18046,N_6264,N_8186);
nor U18047 (N_18047,N_7183,N_6268);
xor U18048 (N_18048,N_5826,N_3617);
nor U18049 (N_18049,N_2010,N_7944);
nor U18050 (N_18050,N_708,N_7780);
xnor U18051 (N_18051,N_4825,N_5147);
nand U18052 (N_18052,N_6979,N_2761);
nand U18053 (N_18053,N_7287,N_4634);
and U18054 (N_18054,N_232,N_6450);
xor U18055 (N_18055,N_9969,N_3478);
nor U18056 (N_18056,N_9861,N_877);
nand U18057 (N_18057,N_2562,N_521);
xor U18058 (N_18058,N_1722,N_3690);
or U18059 (N_18059,N_7517,N_9893);
xor U18060 (N_18060,N_8192,N_3938);
nand U18061 (N_18061,N_9975,N_2835);
nand U18062 (N_18062,N_7821,N_6616);
nand U18063 (N_18063,N_4762,N_5082);
nor U18064 (N_18064,N_6264,N_8026);
xnor U18065 (N_18065,N_4348,N_3582);
xor U18066 (N_18066,N_4697,N_4950);
nor U18067 (N_18067,N_5982,N_9131);
and U18068 (N_18068,N_5829,N_7470);
and U18069 (N_18069,N_7207,N_3292);
nor U18070 (N_18070,N_3476,N_7481);
or U18071 (N_18071,N_6998,N_6572);
xor U18072 (N_18072,N_7255,N_4047);
xor U18073 (N_18073,N_9700,N_4445);
or U18074 (N_18074,N_6129,N_4098);
or U18075 (N_18075,N_5648,N_5437);
nand U18076 (N_18076,N_7935,N_6509);
and U18077 (N_18077,N_666,N_7186);
or U18078 (N_18078,N_7391,N_9358);
xor U18079 (N_18079,N_5342,N_5238);
nor U18080 (N_18080,N_7177,N_4716);
or U18081 (N_18081,N_9697,N_1379);
nand U18082 (N_18082,N_932,N_5070);
nand U18083 (N_18083,N_3367,N_6057);
and U18084 (N_18084,N_9711,N_5624);
or U18085 (N_18085,N_9974,N_1140);
or U18086 (N_18086,N_7909,N_2772);
nor U18087 (N_18087,N_3137,N_939);
nand U18088 (N_18088,N_3704,N_4600);
xor U18089 (N_18089,N_3358,N_8451);
nand U18090 (N_18090,N_1162,N_4183);
xnor U18091 (N_18091,N_8673,N_4085);
nand U18092 (N_18092,N_7526,N_8146);
nor U18093 (N_18093,N_5100,N_46);
or U18094 (N_18094,N_1641,N_3006);
and U18095 (N_18095,N_8041,N_273);
nor U18096 (N_18096,N_2976,N_4382);
nor U18097 (N_18097,N_6126,N_5333);
nand U18098 (N_18098,N_7088,N_8024);
nor U18099 (N_18099,N_775,N_4423);
or U18100 (N_18100,N_7146,N_6701);
nor U18101 (N_18101,N_274,N_6515);
nand U18102 (N_18102,N_9836,N_5021);
or U18103 (N_18103,N_13,N_8489);
xnor U18104 (N_18104,N_5616,N_4380);
nand U18105 (N_18105,N_5344,N_3410);
and U18106 (N_18106,N_4644,N_1756);
or U18107 (N_18107,N_9314,N_1313);
and U18108 (N_18108,N_5332,N_9181);
nand U18109 (N_18109,N_9945,N_5329);
xnor U18110 (N_18110,N_7445,N_8534);
xor U18111 (N_18111,N_111,N_5398);
nor U18112 (N_18112,N_9502,N_6420);
and U18113 (N_18113,N_723,N_4689);
nand U18114 (N_18114,N_9802,N_1216);
and U18115 (N_18115,N_1078,N_8704);
or U18116 (N_18116,N_997,N_6432);
and U18117 (N_18117,N_6205,N_9517);
nand U18118 (N_18118,N_1288,N_2285);
nand U18119 (N_18119,N_9308,N_3931);
nand U18120 (N_18120,N_3737,N_3452);
nand U18121 (N_18121,N_4111,N_6714);
and U18122 (N_18122,N_7134,N_263);
nor U18123 (N_18123,N_5190,N_3705);
nor U18124 (N_18124,N_892,N_6539);
nand U18125 (N_18125,N_7586,N_1404);
xor U18126 (N_18126,N_6498,N_5101);
xnor U18127 (N_18127,N_7133,N_3622);
xor U18128 (N_18128,N_9414,N_8727);
nor U18129 (N_18129,N_9104,N_4812);
nor U18130 (N_18130,N_9940,N_3529);
nand U18131 (N_18131,N_326,N_9405);
nand U18132 (N_18132,N_4999,N_8054);
or U18133 (N_18133,N_6677,N_3186);
xor U18134 (N_18134,N_4698,N_2885);
and U18135 (N_18135,N_9393,N_5577);
or U18136 (N_18136,N_5496,N_6243);
or U18137 (N_18137,N_4989,N_6927);
xnor U18138 (N_18138,N_6062,N_2968);
or U18139 (N_18139,N_9524,N_4166);
and U18140 (N_18140,N_7991,N_7401);
and U18141 (N_18141,N_9513,N_1150);
or U18142 (N_18142,N_6562,N_2738);
xnor U18143 (N_18143,N_5669,N_1711);
xor U18144 (N_18144,N_6399,N_8404);
nor U18145 (N_18145,N_3216,N_585);
or U18146 (N_18146,N_9720,N_7572);
xnor U18147 (N_18147,N_1365,N_8682);
xnor U18148 (N_18148,N_4874,N_9197);
nand U18149 (N_18149,N_1103,N_2799);
and U18150 (N_18150,N_1705,N_2731);
xnor U18151 (N_18151,N_9776,N_4217);
nor U18152 (N_18152,N_4142,N_860);
or U18153 (N_18153,N_6269,N_7128);
and U18154 (N_18154,N_9432,N_8986);
and U18155 (N_18155,N_2530,N_2048);
xnor U18156 (N_18156,N_4280,N_7777);
nor U18157 (N_18157,N_9454,N_9313);
and U18158 (N_18158,N_5898,N_8962);
nor U18159 (N_18159,N_5921,N_2660);
nor U18160 (N_18160,N_8010,N_8881);
or U18161 (N_18161,N_7412,N_8264);
or U18162 (N_18162,N_6863,N_5014);
xnor U18163 (N_18163,N_7678,N_9451);
or U18164 (N_18164,N_6082,N_4340);
nand U18165 (N_18165,N_2171,N_2233);
and U18166 (N_18166,N_9044,N_9898);
and U18167 (N_18167,N_8096,N_8134);
xor U18168 (N_18168,N_870,N_5929);
nand U18169 (N_18169,N_6189,N_4461);
or U18170 (N_18170,N_4561,N_8781);
or U18171 (N_18171,N_9985,N_9035);
or U18172 (N_18172,N_6851,N_6569);
nor U18173 (N_18173,N_9067,N_8435);
xor U18174 (N_18174,N_3180,N_7969);
xor U18175 (N_18175,N_2678,N_1545);
or U18176 (N_18176,N_1443,N_6216);
and U18177 (N_18177,N_9371,N_5668);
and U18178 (N_18178,N_4999,N_2441);
xor U18179 (N_18179,N_3979,N_5098);
nand U18180 (N_18180,N_7396,N_6711);
or U18181 (N_18181,N_9166,N_7945);
nor U18182 (N_18182,N_7619,N_3723);
and U18183 (N_18183,N_523,N_6526);
and U18184 (N_18184,N_7418,N_2079);
nor U18185 (N_18185,N_4234,N_1619);
and U18186 (N_18186,N_5067,N_676);
and U18187 (N_18187,N_7247,N_5921);
nand U18188 (N_18188,N_9134,N_8089);
xnor U18189 (N_18189,N_1686,N_5742);
xor U18190 (N_18190,N_9615,N_3784);
nand U18191 (N_18191,N_4121,N_1485);
nor U18192 (N_18192,N_2164,N_3953);
and U18193 (N_18193,N_3745,N_3779);
nor U18194 (N_18194,N_2335,N_9652);
nor U18195 (N_18195,N_9443,N_4402);
and U18196 (N_18196,N_1963,N_5661);
nor U18197 (N_18197,N_4432,N_1141);
nor U18198 (N_18198,N_1544,N_7018);
or U18199 (N_18199,N_6162,N_7115);
xor U18200 (N_18200,N_5815,N_9388);
and U18201 (N_18201,N_7477,N_8505);
xnor U18202 (N_18202,N_5889,N_5912);
nand U18203 (N_18203,N_3482,N_3006);
or U18204 (N_18204,N_9928,N_4081);
and U18205 (N_18205,N_1180,N_4213);
nor U18206 (N_18206,N_4756,N_9643);
and U18207 (N_18207,N_6436,N_2715);
or U18208 (N_18208,N_7497,N_8709);
nand U18209 (N_18209,N_4478,N_712);
or U18210 (N_18210,N_3762,N_7949);
or U18211 (N_18211,N_2316,N_1515);
xor U18212 (N_18212,N_588,N_2225);
nor U18213 (N_18213,N_4987,N_1041);
nor U18214 (N_18214,N_4352,N_6809);
and U18215 (N_18215,N_5519,N_5014);
nand U18216 (N_18216,N_9042,N_887);
xnor U18217 (N_18217,N_1296,N_4152);
nand U18218 (N_18218,N_557,N_413);
nor U18219 (N_18219,N_4137,N_9964);
nand U18220 (N_18220,N_763,N_4314);
and U18221 (N_18221,N_5902,N_6703);
nor U18222 (N_18222,N_9253,N_9503);
xor U18223 (N_18223,N_9447,N_8892);
and U18224 (N_18224,N_5577,N_5475);
nand U18225 (N_18225,N_9065,N_7295);
and U18226 (N_18226,N_6936,N_3301);
nand U18227 (N_18227,N_4944,N_3451);
nor U18228 (N_18228,N_5760,N_2656);
nor U18229 (N_18229,N_4459,N_3300);
nor U18230 (N_18230,N_920,N_3540);
nor U18231 (N_18231,N_220,N_8185);
nor U18232 (N_18232,N_7703,N_3891);
nand U18233 (N_18233,N_8941,N_4097);
nor U18234 (N_18234,N_4953,N_878);
nor U18235 (N_18235,N_2505,N_1454);
xor U18236 (N_18236,N_16,N_6133);
nor U18237 (N_18237,N_7392,N_3574);
nand U18238 (N_18238,N_2528,N_3021);
nor U18239 (N_18239,N_7208,N_3171);
xnor U18240 (N_18240,N_3484,N_8961);
nand U18241 (N_18241,N_8540,N_3550);
and U18242 (N_18242,N_3403,N_2136);
nand U18243 (N_18243,N_675,N_2035);
nor U18244 (N_18244,N_4028,N_1101);
or U18245 (N_18245,N_8123,N_5546);
nand U18246 (N_18246,N_92,N_547);
nor U18247 (N_18247,N_3163,N_5478);
xnor U18248 (N_18248,N_1788,N_1737);
and U18249 (N_18249,N_2399,N_6933);
xnor U18250 (N_18250,N_3085,N_671);
nand U18251 (N_18251,N_9734,N_329);
and U18252 (N_18252,N_6838,N_3329);
and U18253 (N_18253,N_1403,N_732);
or U18254 (N_18254,N_1994,N_1913);
or U18255 (N_18255,N_8467,N_1442);
and U18256 (N_18256,N_717,N_7632);
nand U18257 (N_18257,N_8427,N_951);
or U18258 (N_18258,N_6081,N_861);
nor U18259 (N_18259,N_6066,N_4490);
and U18260 (N_18260,N_7191,N_6698);
nand U18261 (N_18261,N_3716,N_3964);
xnor U18262 (N_18262,N_9572,N_6374);
xnor U18263 (N_18263,N_5211,N_3028);
or U18264 (N_18264,N_1320,N_3798);
xor U18265 (N_18265,N_807,N_3356);
nor U18266 (N_18266,N_1727,N_6511);
and U18267 (N_18267,N_1211,N_5442);
and U18268 (N_18268,N_3577,N_8658);
xor U18269 (N_18269,N_9100,N_1795);
nor U18270 (N_18270,N_8880,N_4818);
and U18271 (N_18271,N_1251,N_5500);
nor U18272 (N_18272,N_9132,N_4097);
nand U18273 (N_18273,N_4101,N_6032);
and U18274 (N_18274,N_6393,N_7189);
nand U18275 (N_18275,N_8865,N_5680);
nand U18276 (N_18276,N_8972,N_8896);
or U18277 (N_18277,N_3539,N_3301);
xnor U18278 (N_18278,N_3911,N_5539);
nand U18279 (N_18279,N_8571,N_5957);
nand U18280 (N_18280,N_2659,N_7423);
xor U18281 (N_18281,N_4421,N_6312);
nor U18282 (N_18282,N_2741,N_7337);
nand U18283 (N_18283,N_6448,N_8827);
nand U18284 (N_18284,N_7737,N_8522);
nand U18285 (N_18285,N_6730,N_9140);
nand U18286 (N_18286,N_1793,N_868);
xnor U18287 (N_18287,N_9546,N_87);
xnor U18288 (N_18288,N_3496,N_548);
nor U18289 (N_18289,N_5879,N_4594);
nor U18290 (N_18290,N_9271,N_2502);
and U18291 (N_18291,N_4891,N_4974);
nor U18292 (N_18292,N_8659,N_5557);
nand U18293 (N_18293,N_2558,N_7231);
nor U18294 (N_18294,N_672,N_7496);
or U18295 (N_18295,N_3677,N_8851);
and U18296 (N_18296,N_3949,N_8266);
nor U18297 (N_18297,N_7250,N_442);
or U18298 (N_18298,N_2798,N_2248);
xnor U18299 (N_18299,N_6169,N_1040);
xnor U18300 (N_18300,N_6777,N_9973);
nor U18301 (N_18301,N_7719,N_9176);
nand U18302 (N_18302,N_4444,N_8786);
or U18303 (N_18303,N_4787,N_3737);
nand U18304 (N_18304,N_4775,N_2481);
nor U18305 (N_18305,N_4937,N_6038);
nor U18306 (N_18306,N_8479,N_2736);
or U18307 (N_18307,N_464,N_7462);
or U18308 (N_18308,N_53,N_1093);
nand U18309 (N_18309,N_4485,N_2960);
xor U18310 (N_18310,N_4602,N_9636);
xor U18311 (N_18311,N_445,N_3475);
nor U18312 (N_18312,N_6272,N_9811);
and U18313 (N_18313,N_9646,N_2927);
nor U18314 (N_18314,N_3809,N_6594);
nor U18315 (N_18315,N_6676,N_3476);
or U18316 (N_18316,N_5982,N_5150);
nand U18317 (N_18317,N_8600,N_937);
xnor U18318 (N_18318,N_8964,N_6197);
nor U18319 (N_18319,N_2759,N_3049);
nor U18320 (N_18320,N_7248,N_8791);
or U18321 (N_18321,N_5882,N_3586);
xor U18322 (N_18322,N_7477,N_1654);
nor U18323 (N_18323,N_6902,N_2845);
and U18324 (N_18324,N_5516,N_2455);
xor U18325 (N_18325,N_2812,N_8876);
nand U18326 (N_18326,N_4035,N_7612);
or U18327 (N_18327,N_3163,N_7510);
xor U18328 (N_18328,N_6366,N_6032);
and U18329 (N_18329,N_9763,N_4640);
or U18330 (N_18330,N_5625,N_4659);
nor U18331 (N_18331,N_3257,N_2074);
or U18332 (N_18332,N_1733,N_8753);
and U18333 (N_18333,N_5395,N_7475);
xnor U18334 (N_18334,N_5654,N_8772);
or U18335 (N_18335,N_7888,N_6743);
xor U18336 (N_18336,N_1173,N_6059);
xnor U18337 (N_18337,N_5411,N_1974);
or U18338 (N_18338,N_1078,N_2770);
and U18339 (N_18339,N_7578,N_912);
xnor U18340 (N_18340,N_9005,N_9586);
or U18341 (N_18341,N_3089,N_691);
nor U18342 (N_18342,N_5275,N_3435);
nor U18343 (N_18343,N_7501,N_7259);
and U18344 (N_18344,N_4878,N_324);
nor U18345 (N_18345,N_9822,N_180);
nor U18346 (N_18346,N_7862,N_9844);
xnor U18347 (N_18347,N_6195,N_3541);
nor U18348 (N_18348,N_783,N_4903);
nor U18349 (N_18349,N_933,N_6523);
or U18350 (N_18350,N_8308,N_5712);
or U18351 (N_18351,N_1997,N_4365);
or U18352 (N_18352,N_2922,N_638);
xnor U18353 (N_18353,N_6620,N_5726);
xor U18354 (N_18354,N_36,N_4922);
or U18355 (N_18355,N_8838,N_1668);
or U18356 (N_18356,N_2538,N_2132);
xor U18357 (N_18357,N_446,N_5413);
or U18358 (N_18358,N_8529,N_3706);
nand U18359 (N_18359,N_9438,N_8377);
nand U18360 (N_18360,N_1699,N_4267);
xor U18361 (N_18361,N_8659,N_8693);
xor U18362 (N_18362,N_8843,N_1377);
nand U18363 (N_18363,N_5609,N_6158);
nor U18364 (N_18364,N_1228,N_3274);
nor U18365 (N_18365,N_4542,N_150);
xor U18366 (N_18366,N_6462,N_6196);
xnor U18367 (N_18367,N_444,N_4424);
or U18368 (N_18368,N_5671,N_6774);
or U18369 (N_18369,N_6896,N_3498);
nand U18370 (N_18370,N_2589,N_4286);
or U18371 (N_18371,N_6080,N_1876);
nor U18372 (N_18372,N_1325,N_2174);
nand U18373 (N_18373,N_7324,N_7890);
and U18374 (N_18374,N_9549,N_492);
nor U18375 (N_18375,N_5587,N_47);
nor U18376 (N_18376,N_1950,N_8202);
or U18377 (N_18377,N_110,N_3674);
nand U18378 (N_18378,N_9140,N_4187);
nor U18379 (N_18379,N_446,N_1948);
nand U18380 (N_18380,N_3498,N_4440);
nand U18381 (N_18381,N_8131,N_7169);
or U18382 (N_18382,N_9123,N_9156);
nor U18383 (N_18383,N_1676,N_6455);
and U18384 (N_18384,N_6379,N_5931);
or U18385 (N_18385,N_4853,N_5199);
nor U18386 (N_18386,N_9518,N_9845);
xnor U18387 (N_18387,N_8712,N_3583);
nor U18388 (N_18388,N_9925,N_2024);
or U18389 (N_18389,N_2856,N_8094);
nor U18390 (N_18390,N_6587,N_9048);
nand U18391 (N_18391,N_1112,N_6012);
nor U18392 (N_18392,N_7008,N_5316);
nand U18393 (N_18393,N_4104,N_7161);
nor U18394 (N_18394,N_4883,N_2645);
nor U18395 (N_18395,N_8486,N_1525);
nand U18396 (N_18396,N_8549,N_6484);
or U18397 (N_18397,N_2409,N_6128);
xor U18398 (N_18398,N_8353,N_9699);
nand U18399 (N_18399,N_7132,N_2325);
xor U18400 (N_18400,N_2551,N_3224);
nand U18401 (N_18401,N_9858,N_3944);
and U18402 (N_18402,N_6290,N_1780);
and U18403 (N_18403,N_3710,N_5231);
or U18404 (N_18404,N_9711,N_7865);
nor U18405 (N_18405,N_5674,N_549);
nor U18406 (N_18406,N_3276,N_2748);
nor U18407 (N_18407,N_7951,N_4980);
or U18408 (N_18408,N_7846,N_4302);
nor U18409 (N_18409,N_7082,N_2873);
xor U18410 (N_18410,N_6327,N_9252);
and U18411 (N_18411,N_7447,N_2364);
or U18412 (N_18412,N_9021,N_9105);
nand U18413 (N_18413,N_3345,N_5163);
xor U18414 (N_18414,N_6586,N_4503);
nor U18415 (N_18415,N_3988,N_6683);
nor U18416 (N_18416,N_652,N_249);
and U18417 (N_18417,N_8100,N_5840);
nor U18418 (N_18418,N_3849,N_5326);
xor U18419 (N_18419,N_9757,N_4072);
nand U18420 (N_18420,N_9250,N_7182);
or U18421 (N_18421,N_9260,N_55);
and U18422 (N_18422,N_4125,N_222);
and U18423 (N_18423,N_353,N_5418);
and U18424 (N_18424,N_8394,N_6167);
xor U18425 (N_18425,N_6956,N_5491);
xor U18426 (N_18426,N_1582,N_9131);
and U18427 (N_18427,N_9824,N_1345);
nand U18428 (N_18428,N_2524,N_882);
or U18429 (N_18429,N_1696,N_3635);
and U18430 (N_18430,N_3351,N_8510);
xor U18431 (N_18431,N_6353,N_2984);
and U18432 (N_18432,N_4722,N_1356);
nand U18433 (N_18433,N_5227,N_7417);
nor U18434 (N_18434,N_9401,N_1636);
nand U18435 (N_18435,N_4197,N_6429);
and U18436 (N_18436,N_4346,N_8830);
nand U18437 (N_18437,N_2043,N_5897);
nand U18438 (N_18438,N_4338,N_4980);
nand U18439 (N_18439,N_8987,N_5539);
nand U18440 (N_18440,N_2144,N_534);
or U18441 (N_18441,N_4046,N_7932);
xnor U18442 (N_18442,N_1040,N_1019);
and U18443 (N_18443,N_9642,N_6434);
nand U18444 (N_18444,N_6455,N_1307);
and U18445 (N_18445,N_6787,N_4832);
nand U18446 (N_18446,N_3590,N_8298);
nor U18447 (N_18447,N_7154,N_3242);
and U18448 (N_18448,N_1749,N_6489);
nor U18449 (N_18449,N_9561,N_1488);
and U18450 (N_18450,N_3011,N_8351);
xor U18451 (N_18451,N_2940,N_4182);
nor U18452 (N_18452,N_3181,N_394);
nand U18453 (N_18453,N_6646,N_9543);
xor U18454 (N_18454,N_5059,N_1324);
xnor U18455 (N_18455,N_2469,N_8600);
or U18456 (N_18456,N_2437,N_7754);
xor U18457 (N_18457,N_3675,N_2746);
nand U18458 (N_18458,N_2820,N_7670);
nor U18459 (N_18459,N_1017,N_2480);
nor U18460 (N_18460,N_5340,N_7250);
nor U18461 (N_18461,N_7093,N_2630);
xor U18462 (N_18462,N_2590,N_926);
nand U18463 (N_18463,N_2900,N_2159);
and U18464 (N_18464,N_9904,N_3076);
nand U18465 (N_18465,N_2140,N_6824);
xnor U18466 (N_18466,N_4900,N_8576);
nor U18467 (N_18467,N_5103,N_8454);
and U18468 (N_18468,N_7911,N_2625);
and U18469 (N_18469,N_4244,N_7562);
or U18470 (N_18470,N_3065,N_9589);
or U18471 (N_18471,N_2623,N_6250);
and U18472 (N_18472,N_7361,N_6649);
and U18473 (N_18473,N_9094,N_4438);
or U18474 (N_18474,N_117,N_7607);
nand U18475 (N_18475,N_9290,N_2958);
and U18476 (N_18476,N_7762,N_8745);
xnor U18477 (N_18477,N_960,N_1764);
nand U18478 (N_18478,N_3815,N_2236);
nand U18479 (N_18479,N_8822,N_2937);
or U18480 (N_18480,N_9946,N_6321);
nand U18481 (N_18481,N_4671,N_2430);
nor U18482 (N_18482,N_3135,N_9647);
and U18483 (N_18483,N_72,N_6449);
or U18484 (N_18484,N_7651,N_2294);
nor U18485 (N_18485,N_1580,N_6884);
nand U18486 (N_18486,N_7740,N_3358);
and U18487 (N_18487,N_4922,N_2986);
nor U18488 (N_18488,N_9659,N_8471);
and U18489 (N_18489,N_8993,N_1339);
nor U18490 (N_18490,N_6938,N_2973);
xor U18491 (N_18491,N_1980,N_1483);
xnor U18492 (N_18492,N_5028,N_6548);
or U18493 (N_18493,N_9764,N_1195);
or U18494 (N_18494,N_703,N_7820);
nand U18495 (N_18495,N_9087,N_8851);
nand U18496 (N_18496,N_2273,N_2439);
or U18497 (N_18497,N_6972,N_5199);
xor U18498 (N_18498,N_8270,N_7619);
nand U18499 (N_18499,N_6596,N_644);
nand U18500 (N_18500,N_765,N_4094);
xnor U18501 (N_18501,N_2529,N_1172);
nand U18502 (N_18502,N_9301,N_1699);
xnor U18503 (N_18503,N_9041,N_2314);
nand U18504 (N_18504,N_8096,N_5148);
or U18505 (N_18505,N_9493,N_37);
and U18506 (N_18506,N_6917,N_4073);
nand U18507 (N_18507,N_3385,N_4808);
nand U18508 (N_18508,N_3944,N_4650);
nand U18509 (N_18509,N_6407,N_6550);
or U18510 (N_18510,N_9637,N_184);
xor U18511 (N_18511,N_7898,N_4805);
nand U18512 (N_18512,N_6417,N_4940);
or U18513 (N_18513,N_9472,N_1130);
xor U18514 (N_18514,N_6073,N_5606);
and U18515 (N_18515,N_233,N_1002);
nor U18516 (N_18516,N_5986,N_8059);
or U18517 (N_18517,N_5661,N_3905);
or U18518 (N_18518,N_3735,N_1518);
nand U18519 (N_18519,N_1180,N_4177);
xor U18520 (N_18520,N_9482,N_2525);
xnor U18521 (N_18521,N_7334,N_7242);
nor U18522 (N_18522,N_7833,N_2405);
nand U18523 (N_18523,N_5725,N_8270);
xnor U18524 (N_18524,N_9766,N_3785);
nor U18525 (N_18525,N_6866,N_4779);
nand U18526 (N_18526,N_7881,N_8564);
nand U18527 (N_18527,N_9576,N_5189);
xnor U18528 (N_18528,N_7051,N_631);
nor U18529 (N_18529,N_6104,N_6375);
or U18530 (N_18530,N_3508,N_817);
xor U18531 (N_18531,N_479,N_5695);
and U18532 (N_18532,N_1246,N_124);
xnor U18533 (N_18533,N_567,N_1333);
nor U18534 (N_18534,N_7964,N_2521);
nand U18535 (N_18535,N_2732,N_5014);
or U18536 (N_18536,N_6193,N_2851);
xor U18537 (N_18537,N_5247,N_6685);
xnor U18538 (N_18538,N_533,N_4644);
or U18539 (N_18539,N_3036,N_3633);
xor U18540 (N_18540,N_281,N_2494);
nand U18541 (N_18541,N_4005,N_8731);
and U18542 (N_18542,N_8044,N_1583);
xor U18543 (N_18543,N_7830,N_6025);
and U18544 (N_18544,N_2959,N_2743);
nand U18545 (N_18545,N_3178,N_79);
or U18546 (N_18546,N_3653,N_8338);
and U18547 (N_18547,N_7662,N_7749);
nor U18548 (N_18548,N_548,N_7507);
or U18549 (N_18549,N_158,N_116);
or U18550 (N_18550,N_1821,N_8442);
nand U18551 (N_18551,N_2517,N_6732);
nor U18552 (N_18552,N_887,N_7781);
and U18553 (N_18553,N_8730,N_8272);
or U18554 (N_18554,N_1670,N_4389);
xnor U18555 (N_18555,N_1051,N_1850);
and U18556 (N_18556,N_2726,N_7902);
nor U18557 (N_18557,N_1560,N_2037);
nor U18558 (N_18558,N_2857,N_6956);
or U18559 (N_18559,N_7179,N_3557);
and U18560 (N_18560,N_5089,N_6085);
nand U18561 (N_18561,N_327,N_7786);
or U18562 (N_18562,N_6132,N_8042);
nor U18563 (N_18563,N_632,N_6847);
nand U18564 (N_18564,N_390,N_7002);
or U18565 (N_18565,N_2889,N_9838);
or U18566 (N_18566,N_1957,N_5794);
nor U18567 (N_18567,N_802,N_1500);
nor U18568 (N_18568,N_4615,N_2499);
nor U18569 (N_18569,N_2118,N_6685);
xnor U18570 (N_18570,N_9842,N_6653);
and U18571 (N_18571,N_2088,N_4963);
xnor U18572 (N_18572,N_8766,N_3309);
and U18573 (N_18573,N_7536,N_8938);
or U18574 (N_18574,N_4846,N_3231);
nand U18575 (N_18575,N_382,N_4029);
or U18576 (N_18576,N_1285,N_4920);
xor U18577 (N_18577,N_8867,N_3739);
nor U18578 (N_18578,N_9555,N_9527);
and U18579 (N_18579,N_2215,N_3519);
nor U18580 (N_18580,N_1447,N_9633);
xnor U18581 (N_18581,N_3945,N_7666);
xor U18582 (N_18582,N_8371,N_9129);
and U18583 (N_18583,N_9731,N_1651);
xor U18584 (N_18584,N_6416,N_1331);
xnor U18585 (N_18585,N_1140,N_9990);
nand U18586 (N_18586,N_3476,N_3607);
xor U18587 (N_18587,N_9760,N_6316);
or U18588 (N_18588,N_8238,N_143);
xor U18589 (N_18589,N_6496,N_6486);
nor U18590 (N_18590,N_986,N_5739);
nand U18591 (N_18591,N_474,N_4721);
or U18592 (N_18592,N_3526,N_3322);
xor U18593 (N_18593,N_4418,N_6433);
nand U18594 (N_18594,N_8370,N_1086);
and U18595 (N_18595,N_6888,N_3420);
or U18596 (N_18596,N_4127,N_9380);
nand U18597 (N_18597,N_5284,N_7483);
nor U18598 (N_18598,N_8606,N_3677);
xnor U18599 (N_18599,N_5028,N_9921);
and U18600 (N_18600,N_9977,N_7685);
xnor U18601 (N_18601,N_2363,N_3231);
nor U18602 (N_18602,N_1451,N_7114);
and U18603 (N_18603,N_2092,N_8572);
nand U18604 (N_18604,N_3962,N_9728);
nor U18605 (N_18605,N_593,N_3773);
nand U18606 (N_18606,N_2517,N_6476);
nand U18607 (N_18607,N_3231,N_6002);
nor U18608 (N_18608,N_6408,N_1401);
nand U18609 (N_18609,N_7241,N_8060);
or U18610 (N_18610,N_7170,N_9708);
xnor U18611 (N_18611,N_4238,N_5575);
nand U18612 (N_18612,N_8734,N_8152);
xor U18613 (N_18613,N_8414,N_7943);
and U18614 (N_18614,N_295,N_4063);
nor U18615 (N_18615,N_548,N_9451);
and U18616 (N_18616,N_8808,N_7511);
nor U18617 (N_18617,N_7062,N_7906);
and U18618 (N_18618,N_5448,N_4754);
or U18619 (N_18619,N_240,N_1410);
xnor U18620 (N_18620,N_568,N_2192);
xor U18621 (N_18621,N_532,N_5021);
nand U18622 (N_18622,N_9653,N_1257);
or U18623 (N_18623,N_3779,N_187);
nand U18624 (N_18624,N_2774,N_6941);
xnor U18625 (N_18625,N_6258,N_3182);
and U18626 (N_18626,N_3003,N_4983);
and U18627 (N_18627,N_6600,N_5315);
and U18628 (N_18628,N_2993,N_8420);
nand U18629 (N_18629,N_2360,N_541);
nor U18630 (N_18630,N_5778,N_9355);
xnor U18631 (N_18631,N_7147,N_5549);
or U18632 (N_18632,N_2391,N_9119);
xnor U18633 (N_18633,N_4620,N_4523);
xor U18634 (N_18634,N_6094,N_1175);
or U18635 (N_18635,N_7223,N_194);
xnor U18636 (N_18636,N_7314,N_2748);
nand U18637 (N_18637,N_2139,N_4172);
or U18638 (N_18638,N_8050,N_9892);
or U18639 (N_18639,N_7450,N_3714);
and U18640 (N_18640,N_5585,N_7286);
and U18641 (N_18641,N_8887,N_308);
xnor U18642 (N_18642,N_8806,N_1259);
and U18643 (N_18643,N_8918,N_1473);
and U18644 (N_18644,N_7025,N_8028);
or U18645 (N_18645,N_9533,N_6847);
and U18646 (N_18646,N_1343,N_3768);
xor U18647 (N_18647,N_4283,N_3773);
nand U18648 (N_18648,N_2760,N_6856);
and U18649 (N_18649,N_5024,N_9255);
or U18650 (N_18650,N_4401,N_4919);
nand U18651 (N_18651,N_4967,N_3548);
xor U18652 (N_18652,N_4008,N_3514);
xnor U18653 (N_18653,N_6241,N_5998);
or U18654 (N_18654,N_1349,N_1257);
nor U18655 (N_18655,N_3144,N_7100);
xor U18656 (N_18656,N_8308,N_141);
nor U18657 (N_18657,N_2429,N_817);
nor U18658 (N_18658,N_1219,N_6063);
or U18659 (N_18659,N_6185,N_6384);
or U18660 (N_18660,N_3398,N_7809);
and U18661 (N_18661,N_9078,N_5212);
and U18662 (N_18662,N_857,N_8549);
and U18663 (N_18663,N_2539,N_3798);
xor U18664 (N_18664,N_3189,N_138);
nor U18665 (N_18665,N_841,N_4397);
or U18666 (N_18666,N_7814,N_9533);
and U18667 (N_18667,N_7783,N_4367);
nand U18668 (N_18668,N_5365,N_431);
nand U18669 (N_18669,N_4129,N_6815);
nand U18670 (N_18670,N_6420,N_84);
nand U18671 (N_18671,N_1004,N_890);
nand U18672 (N_18672,N_7799,N_187);
or U18673 (N_18673,N_5703,N_3962);
nor U18674 (N_18674,N_8799,N_5953);
and U18675 (N_18675,N_7122,N_2093);
nand U18676 (N_18676,N_5727,N_2864);
and U18677 (N_18677,N_7892,N_3280);
nor U18678 (N_18678,N_4343,N_8995);
xor U18679 (N_18679,N_3860,N_2659);
and U18680 (N_18680,N_670,N_5741);
nand U18681 (N_18681,N_9696,N_4514);
xor U18682 (N_18682,N_9831,N_4126);
and U18683 (N_18683,N_8428,N_578);
nand U18684 (N_18684,N_47,N_2986);
or U18685 (N_18685,N_7527,N_2689);
or U18686 (N_18686,N_5193,N_6012);
nor U18687 (N_18687,N_3644,N_1717);
xor U18688 (N_18688,N_7138,N_4481);
and U18689 (N_18689,N_3336,N_1965);
xnor U18690 (N_18690,N_6862,N_4993);
or U18691 (N_18691,N_8638,N_103);
and U18692 (N_18692,N_6221,N_7327);
xor U18693 (N_18693,N_1288,N_6119);
xor U18694 (N_18694,N_5210,N_9704);
or U18695 (N_18695,N_2341,N_1555);
nand U18696 (N_18696,N_9310,N_5772);
or U18697 (N_18697,N_5134,N_9078);
and U18698 (N_18698,N_2081,N_1696);
xor U18699 (N_18699,N_558,N_3544);
or U18700 (N_18700,N_5649,N_6538);
or U18701 (N_18701,N_5444,N_1026);
and U18702 (N_18702,N_1240,N_5088);
and U18703 (N_18703,N_8794,N_8912);
and U18704 (N_18704,N_8001,N_9896);
or U18705 (N_18705,N_7738,N_1635);
xnor U18706 (N_18706,N_2525,N_2811);
nor U18707 (N_18707,N_8345,N_4625);
and U18708 (N_18708,N_7699,N_7766);
nand U18709 (N_18709,N_5259,N_7315);
or U18710 (N_18710,N_5348,N_261);
nand U18711 (N_18711,N_6995,N_5734);
nand U18712 (N_18712,N_7828,N_1218);
and U18713 (N_18713,N_4864,N_5980);
and U18714 (N_18714,N_5409,N_6227);
xnor U18715 (N_18715,N_9539,N_1454);
nand U18716 (N_18716,N_6717,N_2203);
nor U18717 (N_18717,N_8301,N_9433);
xor U18718 (N_18718,N_2743,N_9706);
or U18719 (N_18719,N_7386,N_7084);
nor U18720 (N_18720,N_6129,N_6053);
or U18721 (N_18721,N_8357,N_4972);
xnor U18722 (N_18722,N_4157,N_8136);
nand U18723 (N_18723,N_1376,N_6698);
or U18724 (N_18724,N_7435,N_7389);
nor U18725 (N_18725,N_7494,N_1191);
or U18726 (N_18726,N_3024,N_6860);
nor U18727 (N_18727,N_3865,N_3517);
nor U18728 (N_18728,N_7260,N_1463);
xor U18729 (N_18729,N_8644,N_569);
or U18730 (N_18730,N_2479,N_8111);
nor U18731 (N_18731,N_5803,N_9623);
or U18732 (N_18732,N_3008,N_4317);
and U18733 (N_18733,N_2349,N_2672);
nor U18734 (N_18734,N_6506,N_7077);
nor U18735 (N_18735,N_2421,N_2761);
or U18736 (N_18736,N_9143,N_5273);
nand U18737 (N_18737,N_7869,N_9553);
xor U18738 (N_18738,N_7289,N_4673);
or U18739 (N_18739,N_688,N_9294);
and U18740 (N_18740,N_8034,N_5048);
xor U18741 (N_18741,N_795,N_5405);
or U18742 (N_18742,N_986,N_5492);
or U18743 (N_18743,N_5215,N_5037);
nor U18744 (N_18744,N_7459,N_1352);
nand U18745 (N_18745,N_8536,N_7217);
or U18746 (N_18746,N_3546,N_2994);
or U18747 (N_18747,N_548,N_487);
nor U18748 (N_18748,N_4937,N_593);
nor U18749 (N_18749,N_6513,N_4729);
xnor U18750 (N_18750,N_9537,N_9155);
xnor U18751 (N_18751,N_9503,N_1579);
xnor U18752 (N_18752,N_2704,N_7315);
nor U18753 (N_18753,N_7356,N_4368);
and U18754 (N_18754,N_6428,N_1852);
or U18755 (N_18755,N_6007,N_4706);
nand U18756 (N_18756,N_225,N_4855);
and U18757 (N_18757,N_6557,N_2015);
nand U18758 (N_18758,N_2035,N_9615);
or U18759 (N_18759,N_4446,N_1813);
xor U18760 (N_18760,N_7037,N_3734);
xnor U18761 (N_18761,N_9227,N_8845);
xor U18762 (N_18762,N_3692,N_621);
or U18763 (N_18763,N_4719,N_1629);
and U18764 (N_18764,N_7670,N_1543);
or U18765 (N_18765,N_7926,N_5643);
and U18766 (N_18766,N_503,N_5015);
nor U18767 (N_18767,N_4844,N_9884);
or U18768 (N_18768,N_8805,N_5599);
xnor U18769 (N_18769,N_8724,N_3520);
or U18770 (N_18770,N_313,N_5748);
xor U18771 (N_18771,N_1214,N_4881);
and U18772 (N_18772,N_8407,N_2496);
or U18773 (N_18773,N_7592,N_137);
nand U18774 (N_18774,N_8292,N_4292);
nor U18775 (N_18775,N_6407,N_3990);
and U18776 (N_18776,N_3515,N_9888);
or U18777 (N_18777,N_9212,N_7577);
or U18778 (N_18778,N_8440,N_1581);
xor U18779 (N_18779,N_6011,N_2628);
xnor U18780 (N_18780,N_2356,N_6643);
nand U18781 (N_18781,N_1365,N_8213);
nand U18782 (N_18782,N_8490,N_8164);
or U18783 (N_18783,N_2887,N_2483);
xnor U18784 (N_18784,N_8550,N_716);
nor U18785 (N_18785,N_8416,N_2003);
xnor U18786 (N_18786,N_8738,N_2127);
nand U18787 (N_18787,N_4146,N_2981);
and U18788 (N_18788,N_8468,N_222);
or U18789 (N_18789,N_4527,N_447);
xor U18790 (N_18790,N_3225,N_6093);
or U18791 (N_18791,N_9727,N_8193);
nor U18792 (N_18792,N_9312,N_1359);
nand U18793 (N_18793,N_5845,N_1687);
nand U18794 (N_18794,N_3676,N_4415);
xnor U18795 (N_18795,N_4875,N_165);
nor U18796 (N_18796,N_260,N_2842);
nor U18797 (N_18797,N_1384,N_2863);
or U18798 (N_18798,N_8369,N_5502);
and U18799 (N_18799,N_7665,N_4546);
nand U18800 (N_18800,N_3305,N_9753);
nor U18801 (N_18801,N_6394,N_757);
and U18802 (N_18802,N_6457,N_2093);
xor U18803 (N_18803,N_15,N_3571);
nand U18804 (N_18804,N_9218,N_8689);
nand U18805 (N_18805,N_9024,N_7156);
xnor U18806 (N_18806,N_4533,N_2365);
nand U18807 (N_18807,N_9701,N_8249);
xor U18808 (N_18808,N_1248,N_2559);
xor U18809 (N_18809,N_686,N_9827);
nor U18810 (N_18810,N_4179,N_4261);
and U18811 (N_18811,N_3127,N_718);
nor U18812 (N_18812,N_3105,N_6739);
nor U18813 (N_18813,N_3563,N_8189);
xor U18814 (N_18814,N_7685,N_1889);
or U18815 (N_18815,N_2397,N_5992);
and U18816 (N_18816,N_4973,N_1352);
and U18817 (N_18817,N_7608,N_9570);
and U18818 (N_18818,N_7495,N_9957);
or U18819 (N_18819,N_8442,N_2122);
and U18820 (N_18820,N_202,N_4923);
and U18821 (N_18821,N_4219,N_3975);
and U18822 (N_18822,N_8840,N_4187);
or U18823 (N_18823,N_8751,N_4528);
xor U18824 (N_18824,N_6757,N_457);
nand U18825 (N_18825,N_1801,N_3289);
or U18826 (N_18826,N_2627,N_9671);
xor U18827 (N_18827,N_3296,N_3301);
nor U18828 (N_18828,N_6438,N_5725);
xnor U18829 (N_18829,N_1422,N_3646);
and U18830 (N_18830,N_4048,N_2240);
nor U18831 (N_18831,N_2024,N_5335);
xor U18832 (N_18832,N_2759,N_4332);
xor U18833 (N_18833,N_6378,N_6980);
nand U18834 (N_18834,N_363,N_8048);
xor U18835 (N_18835,N_1350,N_9241);
nand U18836 (N_18836,N_5141,N_8534);
xnor U18837 (N_18837,N_3158,N_8094);
and U18838 (N_18838,N_2156,N_6563);
and U18839 (N_18839,N_3687,N_1681);
xor U18840 (N_18840,N_5789,N_1237);
or U18841 (N_18841,N_2540,N_2092);
nand U18842 (N_18842,N_1149,N_5538);
and U18843 (N_18843,N_1738,N_1653);
nor U18844 (N_18844,N_8851,N_5752);
or U18845 (N_18845,N_4276,N_6579);
or U18846 (N_18846,N_1797,N_4893);
and U18847 (N_18847,N_1166,N_5620);
and U18848 (N_18848,N_2381,N_826);
nand U18849 (N_18849,N_2588,N_7558);
and U18850 (N_18850,N_8716,N_1132);
xnor U18851 (N_18851,N_9200,N_9019);
nand U18852 (N_18852,N_2646,N_2616);
and U18853 (N_18853,N_3807,N_9664);
and U18854 (N_18854,N_8394,N_4875);
or U18855 (N_18855,N_9126,N_8732);
or U18856 (N_18856,N_1742,N_7754);
and U18857 (N_18857,N_7373,N_9125);
or U18858 (N_18858,N_9277,N_2940);
or U18859 (N_18859,N_698,N_373);
nor U18860 (N_18860,N_6694,N_3373);
xor U18861 (N_18861,N_7174,N_7544);
or U18862 (N_18862,N_2731,N_592);
or U18863 (N_18863,N_9923,N_7770);
nor U18864 (N_18864,N_3855,N_6643);
or U18865 (N_18865,N_7117,N_6988);
xnor U18866 (N_18866,N_5046,N_5690);
xnor U18867 (N_18867,N_1316,N_2518);
or U18868 (N_18868,N_5405,N_6523);
xor U18869 (N_18869,N_5229,N_1713);
nand U18870 (N_18870,N_3465,N_3610);
or U18871 (N_18871,N_2956,N_4047);
nor U18872 (N_18872,N_560,N_4717);
or U18873 (N_18873,N_8758,N_546);
and U18874 (N_18874,N_20,N_1310);
and U18875 (N_18875,N_2585,N_7911);
nor U18876 (N_18876,N_5812,N_2124);
and U18877 (N_18877,N_6823,N_6890);
nand U18878 (N_18878,N_5590,N_3727);
or U18879 (N_18879,N_2299,N_2888);
or U18880 (N_18880,N_2276,N_9658);
xnor U18881 (N_18881,N_9931,N_5558);
or U18882 (N_18882,N_1351,N_5910);
and U18883 (N_18883,N_3784,N_107);
xor U18884 (N_18884,N_5889,N_4721);
and U18885 (N_18885,N_3280,N_3429);
nor U18886 (N_18886,N_2805,N_3566);
nand U18887 (N_18887,N_2378,N_771);
nand U18888 (N_18888,N_1570,N_7102);
or U18889 (N_18889,N_6092,N_9171);
and U18890 (N_18890,N_6353,N_876);
xor U18891 (N_18891,N_6015,N_3992);
nand U18892 (N_18892,N_9626,N_3554);
and U18893 (N_18893,N_8879,N_2764);
xnor U18894 (N_18894,N_7595,N_6073);
nor U18895 (N_18895,N_8487,N_2552);
nor U18896 (N_18896,N_1913,N_7265);
nand U18897 (N_18897,N_9147,N_3112);
or U18898 (N_18898,N_4013,N_3984);
nor U18899 (N_18899,N_5373,N_6344);
nor U18900 (N_18900,N_7827,N_5320);
or U18901 (N_18901,N_7418,N_578);
xor U18902 (N_18902,N_7408,N_3175);
nand U18903 (N_18903,N_5305,N_1468);
nand U18904 (N_18904,N_8955,N_7385);
or U18905 (N_18905,N_8160,N_9835);
nor U18906 (N_18906,N_9773,N_9298);
nand U18907 (N_18907,N_6954,N_223);
or U18908 (N_18908,N_2591,N_677);
or U18909 (N_18909,N_4015,N_6132);
nand U18910 (N_18910,N_1088,N_9081);
xor U18911 (N_18911,N_7091,N_4608);
or U18912 (N_18912,N_8729,N_2129);
or U18913 (N_18913,N_2773,N_900);
or U18914 (N_18914,N_3991,N_970);
or U18915 (N_18915,N_9143,N_3064);
and U18916 (N_18916,N_5492,N_1520);
nor U18917 (N_18917,N_9777,N_4133);
xor U18918 (N_18918,N_5234,N_8465);
nor U18919 (N_18919,N_9889,N_9977);
or U18920 (N_18920,N_4548,N_9500);
or U18921 (N_18921,N_9398,N_8245);
nor U18922 (N_18922,N_7212,N_5961);
xor U18923 (N_18923,N_492,N_6170);
and U18924 (N_18924,N_3193,N_9937);
xor U18925 (N_18925,N_659,N_4952);
nand U18926 (N_18926,N_3810,N_497);
or U18927 (N_18927,N_1656,N_3775);
or U18928 (N_18928,N_6858,N_6516);
xnor U18929 (N_18929,N_3643,N_9625);
xnor U18930 (N_18930,N_1470,N_5550);
and U18931 (N_18931,N_1959,N_23);
xnor U18932 (N_18932,N_964,N_8574);
nand U18933 (N_18933,N_2678,N_4603);
nand U18934 (N_18934,N_5477,N_3965);
xnor U18935 (N_18935,N_7101,N_3258);
or U18936 (N_18936,N_2447,N_9210);
and U18937 (N_18937,N_4542,N_5256);
or U18938 (N_18938,N_5902,N_3845);
xnor U18939 (N_18939,N_9870,N_685);
or U18940 (N_18940,N_9980,N_9825);
nor U18941 (N_18941,N_495,N_7365);
nor U18942 (N_18942,N_796,N_8210);
xnor U18943 (N_18943,N_1992,N_7325);
xnor U18944 (N_18944,N_1105,N_3219);
nand U18945 (N_18945,N_4824,N_6830);
nor U18946 (N_18946,N_3063,N_4883);
nand U18947 (N_18947,N_7678,N_9668);
or U18948 (N_18948,N_595,N_6698);
and U18949 (N_18949,N_23,N_8463);
or U18950 (N_18950,N_5367,N_5288);
nand U18951 (N_18951,N_4710,N_7562);
or U18952 (N_18952,N_8354,N_2539);
and U18953 (N_18953,N_3182,N_4237);
and U18954 (N_18954,N_6945,N_1089);
xnor U18955 (N_18955,N_4386,N_2821);
and U18956 (N_18956,N_8192,N_9652);
or U18957 (N_18957,N_7181,N_231);
xnor U18958 (N_18958,N_6376,N_7930);
nand U18959 (N_18959,N_6574,N_7171);
nand U18960 (N_18960,N_1324,N_7484);
nor U18961 (N_18961,N_7303,N_2335);
or U18962 (N_18962,N_4312,N_3397);
nand U18963 (N_18963,N_1074,N_9281);
or U18964 (N_18964,N_1872,N_2132);
xor U18965 (N_18965,N_950,N_1854);
and U18966 (N_18966,N_8689,N_8669);
or U18967 (N_18967,N_6196,N_7144);
nand U18968 (N_18968,N_1930,N_4222);
xor U18969 (N_18969,N_6867,N_7725);
and U18970 (N_18970,N_9231,N_8904);
nand U18971 (N_18971,N_9393,N_7846);
xnor U18972 (N_18972,N_6943,N_7385);
nand U18973 (N_18973,N_3310,N_4189);
nand U18974 (N_18974,N_7339,N_6098);
and U18975 (N_18975,N_2979,N_1093);
nor U18976 (N_18976,N_8605,N_8193);
or U18977 (N_18977,N_5597,N_7650);
xor U18978 (N_18978,N_6167,N_2927);
nand U18979 (N_18979,N_6695,N_3626);
nand U18980 (N_18980,N_2730,N_4546);
nand U18981 (N_18981,N_764,N_7850);
nor U18982 (N_18982,N_230,N_7718);
nor U18983 (N_18983,N_5531,N_4911);
xor U18984 (N_18984,N_1797,N_2446);
and U18985 (N_18985,N_5403,N_2451);
nor U18986 (N_18986,N_6237,N_1028);
xor U18987 (N_18987,N_4824,N_4989);
and U18988 (N_18988,N_9819,N_9201);
or U18989 (N_18989,N_790,N_833);
or U18990 (N_18990,N_7645,N_8451);
nand U18991 (N_18991,N_8868,N_5005);
nand U18992 (N_18992,N_5734,N_485);
nand U18993 (N_18993,N_8726,N_2516);
and U18994 (N_18994,N_5902,N_5798);
xor U18995 (N_18995,N_2673,N_1913);
and U18996 (N_18996,N_9466,N_2824);
nor U18997 (N_18997,N_5703,N_235);
xor U18998 (N_18998,N_1513,N_178);
nand U18999 (N_18999,N_7585,N_9678);
nor U19000 (N_19000,N_7613,N_4194);
nor U19001 (N_19001,N_6940,N_1616);
and U19002 (N_19002,N_1250,N_6146);
or U19003 (N_19003,N_3182,N_1130);
or U19004 (N_19004,N_9620,N_7938);
and U19005 (N_19005,N_7355,N_8802);
and U19006 (N_19006,N_9210,N_1473);
nand U19007 (N_19007,N_6652,N_7647);
nor U19008 (N_19008,N_1401,N_6938);
and U19009 (N_19009,N_6383,N_1156);
xor U19010 (N_19010,N_3408,N_5568);
or U19011 (N_19011,N_7551,N_8977);
xor U19012 (N_19012,N_5527,N_533);
nor U19013 (N_19013,N_5609,N_9259);
xor U19014 (N_19014,N_680,N_1925);
xnor U19015 (N_19015,N_3631,N_48);
xnor U19016 (N_19016,N_1823,N_8211);
nand U19017 (N_19017,N_7469,N_1816);
and U19018 (N_19018,N_7947,N_3637);
nand U19019 (N_19019,N_9679,N_7036);
and U19020 (N_19020,N_833,N_1383);
nand U19021 (N_19021,N_3139,N_1542);
nor U19022 (N_19022,N_4249,N_6311);
nand U19023 (N_19023,N_8414,N_2331);
or U19024 (N_19024,N_7016,N_3855);
nor U19025 (N_19025,N_785,N_2958);
xnor U19026 (N_19026,N_8399,N_9361);
xnor U19027 (N_19027,N_4618,N_5422);
and U19028 (N_19028,N_9186,N_7648);
or U19029 (N_19029,N_9412,N_3901);
nand U19030 (N_19030,N_5815,N_5788);
xor U19031 (N_19031,N_8780,N_3466);
and U19032 (N_19032,N_8720,N_2989);
or U19033 (N_19033,N_8025,N_5098);
or U19034 (N_19034,N_6662,N_5727);
nor U19035 (N_19035,N_8737,N_3529);
xnor U19036 (N_19036,N_5208,N_3047);
xnor U19037 (N_19037,N_8311,N_8775);
nand U19038 (N_19038,N_3384,N_4863);
nand U19039 (N_19039,N_2492,N_184);
and U19040 (N_19040,N_7070,N_8309);
nor U19041 (N_19041,N_5186,N_2055);
and U19042 (N_19042,N_5502,N_5184);
and U19043 (N_19043,N_7712,N_5215);
and U19044 (N_19044,N_9515,N_52);
nor U19045 (N_19045,N_2727,N_3377);
nand U19046 (N_19046,N_7821,N_5665);
and U19047 (N_19047,N_9254,N_7490);
nor U19048 (N_19048,N_1470,N_5263);
xnor U19049 (N_19049,N_4708,N_8179);
nand U19050 (N_19050,N_2860,N_2846);
nand U19051 (N_19051,N_3207,N_9961);
xnor U19052 (N_19052,N_6110,N_2393);
or U19053 (N_19053,N_8681,N_6452);
xor U19054 (N_19054,N_4893,N_5574);
xor U19055 (N_19055,N_9677,N_3071);
and U19056 (N_19056,N_7643,N_729);
or U19057 (N_19057,N_2308,N_5339);
or U19058 (N_19058,N_6313,N_1286);
and U19059 (N_19059,N_9827,N_8804);
and U19060 (N_19060,N_5306,N_6093);
or U19061 (N_19061,N_9672,N_5650);
nor U19062 (N_19062,N_9471,N_2790);
or U19063 (N_19063,N_7578,N_156);
nand U19064 (N_19064,N_9022,N_1258);
nand U19065 (N_19065,N_1264,N_8314);
nand U19066 (N_19066,N_5858,N_8153);
xor U19067 (N_19067,N_9889,N_3956);
xor U19068 (N_19068,N_2268,N_3904);
and U19069 (N_19069,N_368,N_8762);
and U19070 (N_19070,N_9159,N_4896);
and U19071 (N_19071,N_8620,N_3075);
nor U19072 (N_19072,N_353,N_8381);
nor U19073 (N_19073,N_7850,N_1969);
nor U19074 (N_19074,N_2913,N_4284);
and U19075 (N_19075,N_806,N_9622);
nor U19076 (N_19076,N_7444,N_7874);
nor U19077 (N_19077,N_5739,N_9596);
or U19078 (N_19078,N_1907,N_238);
and U19079 (N_19079,N_2590,N_1375);
nor U19080 (N_19080,N_6984,N_1567);
and U19081 (N_19081,N_551,N_5580);
or U19082 (N_19082,N_1716,N_3619);
and U19083 (N_19083,N_4088,N_1146);
xor U19084 (N_19084,N_9497,N_1744);
or U19085 (N_19085,N_6684,N_4597);
nand U19086 (N_19086,N_3304,N_6968);
or U19087 (N_19087,N_9281,N_3309);
xnor U19088 (N_19088,N_5465,N_5975);
or U19089 (N_19089,N_7816,N_3112);
nand U19090 (N_19090,N_3980,N_3117);
or U19091 (N_19091,N_8964,N_3030);
nand U19092 (N_19092,N_8656,N_7197);
and U19093 (N_19093,N_733,N_9015);
nand U19094 (N_19094,N_8515,N_2299);
nor U19095 (N_19095,N_2374,N_3577);
xnor U19096 (N_19096,N_2766,N_2278);
nand U19097 (N_19097,N_3437,N_8454);
xnor U19098 (N_19098,N_5009,N_1662);
nor U19099 (N_19099,N_3502,N_2955);
or U19100 (N_19100,N_4725,N_1052);
nor U19101 (N_19101,N_9725,N_5772);
or U19102 (N_19102,N_3788,N_8374);
and U19103 (N_19103,N_9627,N_5157);
or U19104 (N_19104,N_5173,N_6613);
and U19105 (N_19105,N_5332,N_3344);
and U19106 (N_19106,N_3094,N_1116);
or U19107 (N_19107,N_7425,N_6100);
or U19108 (N_19108,N_2991,N_6270);
xnor U19109 (N_19109,N_4977,N_8013);
nand U19110 (N_19110,N_5999,N_4866);
nor U19111 (N_19111,N_7523,N_1610);
nand U19112 (N_19112,N_491,N_6920);
or U19113 (N_19113,N_4334,N_8106);
and U19114 (N_19114,N_9562,N_2493);
xnor U19115 (N_19115,N_6982,N_5212);
or U19116 (N_19116,N_1145,N_2473);
and U19117 (N_19117,N_1705,N_7602);
and U19118 (N_19118,N_5047,N_1584);
nand U19119 (N_19119,N_6163,N_3003);
and U19120 (N_19120,N_2531,N_2690);
nor U19121 (N_19121,N_1512,N_9928);
nand U19122 (N_19122,N_2992,N_9202);
nor U19123 (N_19123,N_7608,N_6520);
or U19124 (N_19124,N_2740,N_8763);
nor U19125 (N_19125,N_7827,N_6621);
or U19126 (N_19126,N_4639,N_8039);
nor U19127 (N_19127,N_2477,N_2010);
and U19128 (N_19128,N_1866,N_5487);
xnor U19129 (N_19129,N_9081,N_6213);
nand U19130 (N_19130,N_5665,N_3113);
or U19131 (N_19131,N_3071,N_3834);
nor U19132 (N_19132,N_5287,N_1492);
or U19133 (N_19133,N_1945,N_4990);
nand U19134 (N_19134,N_3163,N_9796);
nor U19135 (N_19135,N_8205,N_5368);
xor U19136 (N_19136,N_7403,N_6527);
or U19137 (N_19137,N_1291,N_6418);
xnor U19138 (N_19138,N_1934,N_6632);
and U19139 (N_19139,N_117,N_2014);
and U19140 (N_19140,N_5537,N_6973);
nor U19141 (N_19141,N_4386,N_3552);
xnor U19142 (N_19142,N_5347,N_913);
or U19143 (N_19143,N_9788,N_2561);
or U19144 (N_19144,N_3705,N_4111);
and U19145 (N_19145,N_8272,N_4276);
xnor U19146 (N_19146,N_2611,N_7587);
and U19147 (N_19147,N_6360,N_4407);
or U19148 (N_19148,N_851,N_3233);
nor U19149 (N_19149,N_6629,N_7053);
and U19150 (N_19150,N_2987,N_4270);
nor U19151 (N_19151,N_5247,N_529);
or U19152 (N_19152,N_3217,N_2152);
xor U19153 (N_19153,N_7474,N_2747);
nor U19154 (N_19154,N_4976,N_3134);
nand U19155 (N_19155,N_7922,N_330);
or U19156 (N_19156,N_9970,N_5308);
nand U19157 (N_19157,N_9549,N_9429);
nor U19158 (N_19158,N_5556,N_3226);
nor U19159 (N_19159,N_5417,N_390);
nand U19160 (N_19160,N_6106,N_633);
nand U19161 (N_19161,N_2837,N_3424);
nor U19162 (N_19162,N_3766,N_9684);
nand U19163 (N_19163,N_3260,N_9391);
nor U19164 (N_19164,N_205,N_1063);
nand U19165 (N_19165,N_5483,N_2810);
and U19166 (N_19166,N_4664,N_3623);
and U19167 (N_19167,N_5382,N_9424);
or U19168 (N_19168,N_5544,N_6529);
nand U19169 (N_19169,N_7700,N_9);
nor U19170 (N_19170,N_2957,N_8926);
and U19171 (N_19171,N_8172,N_9433);
xor U19172 (N_19172,N_1404,N_5179);
nand U19173 (N_19173,N_5971,N_3082);
or U19174 (N_19174,N_8941,N_442);
xnor U19175 (N_19175,N_9005,N_3854);
xor U19176 (N_19176,N_2016,N_6812);
and U19177 (N_19177,N_2825,N_2902);
nand U19178 (N_19178,N_6797,N_8938);
and U19179 (N_19179,N_4786,N_2355);
nor U19180 (N_19180,N_9521,N_8467);
nor U19181 (N_19181,N_4131,N_3661);
xor U19182 (N_19182,N_1473,N_4486);
or U19183 (N_19183,N_7906,N_2663);
nand U19184 (N_19184,N_9205,N_226);
xor U19185 (N_19185,N_8780,N_4743);
nand U19186 (N_19186,N_1728,N_7288);
and U19187 (N_19187,N_8839,N_4469);
or U19188 (N_19188,N_3539,N_3072);
and U19189 (N_19189,N_4754,N_7435);
and U19190 (N_19190,N_294,N_8314);
nand U19191 (N_19191,N_6895,N_2889);
and U19192 (N_19192,N_4045,N_6083);
and U19193 (N_19193,N_6755,N_8286);
nor U19194 (N_19194,N_1883,N_814);
and U19195 (N_19195,N_3095,N_7746);
or U19196 (N_19196,N_8410,N_5637);
and U19197 (N_19197,N_6657,N_732);
and U19198 (N_19198,N_6124,N_7352);
nor U19199 (N_19199,N_5735,N_1558);
or U19200 (N_19200,N_6182,N_4668);
or U19201 (N_19201,N_2922,N_560);
and U19202 (N_19202,N_8849,N_6340);
xnor U19203 (N_19203,N_6992,N_1262);
nor U19204 (N_19204,N_4539,N_3390);
or U19205 (N_19205,N_3046,N_8179);
or U19206 (N_19206,N_412,N_1086);
and U19207 (N_19207,N_3415,N_5528);
xor U19208 (N_19208,N_3497,N_3974);
or U19209 (N_19209,N_7366,N_1881);
or U19210 (N_19210,N_1036,N_3925);
nor U19211 (N_19211,N_9867,N_6170);
nand U19212 (N_19212,N_3056,N_8345);
or U19213 (N_19213,N_4264,N_1818);
or U19214 (N_19214,N_8149,N_6935);
xor U19215 (N_19215,N_3698,N_4945);
or U19216 (N_19216,N_6773,N_1179);
nor U19217 (N_19217,N_5450,N_2880);
nor U19218 (N_19218,N_4568,N_294);
nand U19219 (N_19219,N_9206,N_6388);
or U19220 (N_19220,N_4275,N_1091);
nor U19221 (N_19221,N_4599,N_5024);
or U19222 (N_19222,N_227,N_1722);
or U19223 (N_19223,N_7420,N_1234);
nand U19224 (N_19224,N_9326,N_2529);
and U19225 (N_19225,N_2545,N_8608);
and U19226 (N_19226,N_1013,N_80);
and U19227 (N_19227,N_9402,N_9050);
xnor U19228 (N_19228,N_6031,N_752);
nor U19229 (N_19229,N_918,N_5636);
xor U19230 (N_19230,N_3510,N_6858);
or U19231 (N_19231,N_908,N_3001);
or U19232 (N_19232,N_6883,N_9052);
xor U19233 (N_19233,N_691,N_3375);
xnor U19234 (N_19234,N_9262,N_72);
nor U19235 (N_19235,N_6301,N_1299);
nor U19236 (N_19236,N_6743,N_9188);
nor U19237 (N_19237,N_973,N_1351);
nor U19238 (N_19238,N_1611,N_3685);
or U19239 (N_19239,N_15,N_7960);
xnor U19240 (N_19240,N_143,N_3895);
xor U19241 (N_19241,N_2745,N_5141);
xor U19242 (N_19242,N_8872,N_337);
and U19243 (N_19243,N_2874,N_7977);
and U19244 (N_19244,N_5191,N_8178);
xor U19245 (N_19245,N_9776,N_5175);
and U19246 (N_19246,N_8335,N_2622);
and U19247 (N_19247,N_8244,N_229);
nand U19248 (N_19248,N_5908,N_2640);
and U19249 (N_19249,N_8858,N_4904);
and U19250 (N_19250,N_6220,N_5231);
nand U19251 (N_19251,N_955,N_1705);
nand U19252 (N_19252,N_6900,N_6112);
or U19253 (N_19253,N_112,N_5412);
nand U19254 (N_19254,N_530,N_8205);
xor U19255 (N_19255,N_8259,N_6364);
nand U19256 (N_19256,N_2449,N_460);
and U19257 (N_19257,N_1475,N_9872);
and U19258 (N_19258,N_9591,N_2686);
nand U19259 (N_19259,N_9499,N_7300);
and U19260 (N_19260,N_7173,N_4672);
xor U19261 (N_19261,N_2712,N_9124);
xnor U19262 (N_19262,N_5185,N_3890);
or U19263 (N_19263,N_966,N_8237);
nand U19264 (N_19264,N_4119,N_6583);
nor U19265 (N_19265,N_8167,N_6818);
nor U19266 (N_19266,N_7931,N_8415);
nor U19267 (N_19267,N_1433,N_6474);
nand U19268 (N_19268,N_3760,N_7654);
or U19269 (N_19269,N_9355,N_6979);
nor U19270 (N_19270,N_3160,N_4735);
nand U19271 (N_19271,N_1075,N_8293);
nor U19272 (N_19272,N_1544,N_7153);
and U19273 (N_19273,N_7919,N_1972);
nand U19274 (N_19274,N_322,N_622);
xnor U19275 (N_19275,N_3133,N_959);
or U19276 (N_19276,N_6423,N_8097);
xor U19277 (N_19277,N_6611,N_9231);
xor U19278 (N_19278,N_9276,N_1189);
xnor U19279 (N_19279,N_2240,N_3831);
and U19280 (N_19280,N_9763,N_3074);
nand U19281 (N_19281,N_8253,N_2872);
nor U19282 (N_19282,N_7364,N_5085);
xor U19283 (N_19283,N_750,N_4002);
or U19284 (N_19284,N_7058,N_6036);
xor U19285 (N_19285,N_1679,N_2720);
nand U19286 (N_19286,N_4628,N_3183);
and U19287 (N_19287,N_7786,N_4706);
nand U19288 (N_19288,N_3888,N_3577);
nand U19289 (N_19289,N_3830,N_3909);
nand U19290 (N_19290,N_4642,N_2566);
xnor U19291 (N_19291,N_5783,N_8481);
nand U19292 (N_19292,N_6284,N_538);
nor U19293 (N_19293,N_3909,N_5293);
xnor U19294 (N_19294,N_2413,N_1143);
nand U19295 (N_19295,N_95,N_2484);
xnor U19296 (N_19296,N_1348,N_5755);
or U19297 (N_19297,N_9534,N_6045);
or U19298 (N_19298,N_7051,N_5648);
xor U19299 (N_19299,N_6673,N_8682);
nor U19300 (N_19300,N_1671,N_6228);
nor U19301 (N_19301,N_7259,N_1692);
nand U19302 (N_19302,N_6286,N_9772);
xnor U19303 (N_19303,N_2846,N_6755);
xor U19304 (N_19304,N_4671,N_8490);
nand U19305 (N_19305,N_3878,N_186);
and U19306 (N_19306,N_9192,N_9631);
nor U19307 (N_19307,N_4666,N_6611);
xor U19308 (N_19308,N_7683,N_6407);
nand U19309 (N_19309,N_6116,N_9647);
and U19310 (N_19310,N_7518,N_1994);
and U19311 (N_19311,N_8328,N_2329);
and U19312 (N_19312,N_1483,N_9119);
nor U19313 (N_19313,N_9213,N_4668);
nand U19314 (N_19314,N_6315,N_6692);
nor U19315 (N_19315,N_4247,N_1055);
xor U19316 (N_19316,N_7499,N_312);
and U19317 (N_19317,N_9562,N_7657);
nor U19318 (N_19318,N_6898,N_2846);
nand U19319 (N_19319,N_2238,N_8382);
or U19320 (N_19320,N_6588,N_4018);
or U19321 (N_19321,N_9367,N_7791);
xor U19322 (N_19322,N_2826,N_1504);
nor U19323 (N_19323,N_3473,N_6444);
nand U19324 (N_19324,N_5581,N_2468);
and U19325 (N_19325,N_8013,N_3584);
nand U19326 (N_19326,N_4316,N_2988);
and U19327 (N_19327,N_5886,N_1085);
nand U19328 (N_19328,N_2511,N_5989);
and U19329 (N_19329,N_2980,N_4084);
or U19330 (N_19330,N_8959,N_1520);
nand U19331 (N_19331,N_7654,N_7616);
xnor U19332 (N_19332,N_7496,N_2631);
nand U19333 (N_19333,N_4626,N_5085);
nand U19334 (N_19334,N_6619,N_4264);
or U19335 (N_19335,N_8342,N_2536);
xnor U19336 (N_19336,N_9509,N_2749);
xnor U19337 (N_19337,N_2070,N_4199);
nand U19338 (N_19338,N_679,N_5843);
nor U19339 (N_19339,N_7930,N_8029);
or U19340 (N_19340,N_9977,N_5871);
nand U19341 (N_19341,N_5188,N_771);
nand U19342 (N_19342,N_3848,N_7935);
or U19343 (N_19343,N_3931,N_9817);
or U19344 (N_19344,N_9187,N_4405);
nand U19345 (N_19345,N_6299,N_9094);
xor U19346 (N_19346,N_3326,N_1947);
nor U19347 (N_19347,N_6092,N_542);
nand U19348 (N_19348,N_8376,N_9055);
and U19349 (N_19349,N_2045,N_987);
nor U19350 (N_19350,N_7463,N_4906);
nor U19351 (N_19351,N_7512,N_6834);
and U19352 (N_19352,N_7613,N_7273);
and U19353 (N_19353,N_5772,N_4286);
nor U19354 (N_19354,N_3984,N_1485);
xnor U19355 (N_19355,N_7622,N_2310);
and U19356 (N_19356,N_4607,N_880);
and U19357 (N_19357,N_9362,N_6520);
nor U19358 (N_19358,N_3382,N_9430);
xor U19359 (N_19359,N_4443,N_7331);
nand U19360 (N_19360,N_8198,N_9412);
and U19361 (N_19361,N_9997,N_7249);
and U19362 (N_19362,N_9101,N_5578);
nor U19363 (N_19363,N_3469,N_219);
xnor U19364 (N_19364,N_2562,N_8283);
or U19365 (N_19365,N_5821,N_6921);
xor U19366 (N_19366,N_8862,N_4646);
nor U19367 (N_19367,N_9292,N_6911);
and U19368 (N_19368,N_3172,N_7746);
and U19369 (N_19369,N_2408,N_4234);
nand U19370 (N_19370,N_7160,N_9388);
and U19371 (N_19371,N_7073,N_1658);
nor U19372 (N_19372,N_2072,N_5744);
xor U19373 (N_19373,N_3496,N_3817);
or U19374 (N_19374,N_3382,N_4177);
and U19375 (N_19375,N_9659,N_9318);
xnor U19376 (N_19376,N_841,N_4007);
xor U19377 (N_19377,N_886,N_6048);
or U19378 (N_19378,N_1577,N_3474);
nand U19379 (N_19379,N_4607,N_8906);
nor U19380 (N_19380,N_7234,N_9337);
or U19381 (N_19381,N_8217,N_4206);
nor U19382 (N_19382,N_4091,N_1499);
or U19383 (N_19383,N_9100,N_9700);
or U19384 (N_19384,N_5467,N_3852);
xor U19385 (N_19385,N_9479,N_7390);
nor U19386 (N_19386,N_4308,N_453);
nand U19387 (N_19387,N_6208,N_985);
nand U19388 (N_19388,N_858,N_8202);
nor U19389 (N_19389,N_5340,N_4818);
nand U19390 (N_19390,N_1589,N_5400);
and U19391 (N_19391,N_7365,N_4072);
xor U19392 (N_19392,N_9461,N_9930);
nor U19393 (N_19393,N_6301,N_9554);
nand U19394 (N_19394,N_5797,N_2751);
or U19395 (N_19395,N_5474,N_7219);
nor U19396 (N_19396,N_2914,N_3113);
nor U19397 (N_19397,N_7415,N_2614);
nor U19398 (N_19398,N_4812,N_6638);
or U19399 (N_19399,N_8838,N_3737);
nand U19400 (N_19400,N_7215,N_366);
and U19401 (N_19401,N_1354,N_5967);
xnor U19402 (N_19402,N_5831,N_8406);
xor U19403 (N_19403,N_4514,N_4800);
or U19404 (N_19404,N_6934,N_5808);
or U19405 (N_19405,N_7459,N_4033);
nor U19406 (N_19406,N_2754,N_8744);
and U19407 (N_19407,N_4628,N_3422);
nand U19408 (N_19408,N_4178,N_3624);
nor U19409 (N_19409,N_3790,N_2292);
nand U19410 (N_19410,N_5866,N_8648);
nand U19411 (N_19411,N_6046,N_5939);
nor U19412 (N_19412,N_8071,N_6902);
nand U19413 (N_19413,N_1556,N_1586);
nand U19414 (N_19414,N_134,N_582);
or U19415 (N_19415,N_4167,N_4413);
nor U19416 (N_19416,N_8104,N_3833);
nor U19417 (N_19417,N_1916,N_287);
or U19418 (N_19418,N_560,N_8768);
or U19419 (N_19419,N_9863,N_5520);
nor U19420 (N_19420,N_6305,N_8868);
nand U19421 (N_19421,N_6417,N_1094);
and U19422 (N_19422,N_3497,N_3125);
nor U19423 (N_19423,N_3523,N_3349);
or U19424 (N_19424,N_9636,N_1950);
and U19425 (N_19425,N_6128,N_7918);
nor U19426 (N_19426,N_6542,N_1447);
nor U19427 (N_19427,N_9108,N_821);
nor U19428 (N_19428,N_6817,N_1071);
xor U19429 (N_19429,N_8401,N_1752);
xnor U19430 (N_19430,N_4557,N_5285);
xor U19431 (N_19431,N_6529,N_7989);
nand U19432 (N_19432,N_1573,N_8259);
and U19433 (N_19433,N_5182,N_1236);
and U19434 (N_19434,N_4774,N_9845);
xnor U19435 (N_19435,N_6067,N_8371);
or U19436 (N_19436,N_1718,N_2176);
and U19437 (N_19437,N_1721,N_5976);
or U19438 (N_19438,N_8199,N_5851);
xnor U19439 (N_19439,N_9228,N_2497);
nor U19440 (N_19440,N_615,N_5816);
xnor U19441 (N_19441,N_9140,N_8641);
or U19442 (N_19442,N_3029,N_1783);
nor U19443 (N_19443,N_1785,N_5745);
or U19444 (N_19444,N_8629,N_7327);
and U19445 (N_19445,N_3170,N_2792);
xor U19446 (N_19446,N_904,N_3580);
xor U19447 (N_19447,N_7301,N_8953);
nand U19448 (N_19448,N_2120,N_5462);
or U19449 (N_19449,N_3581,N_2937);
nor U19450 (N_19450,N_2462,N_6068);
nor U19451 (N_19451,N_2825,N_5478);
nand U19452 (N_19452,N_1664,N_3795);
nor U19453 (N_19453,N_8048,N_3958);
or U19454 (N_19454,N_7298,N_1590);
xnor U19455 (N_19455,N_3242,N_603);
or U19456 (N_19456,N_2580,N_1945);
and U19457 (N_19457,N_5410,N_9619);
xnor U19458 (N_19458,N_8194,N_3421);
nand U19459 (N_19459,N_7335,N_4395);
and U19460 (N_19460,N_4240,N_3957);
nand U19461 (N_19461,N_5860,N_544);
nor U19462 (N_19462,N_4182,N_4932);
xor U19463 (N_19463,N_2650,N_7518);
nand U19464 (N_19464,N_7262,N_1781);
or U19465 (N_19465,N_6741,N_377);
xor U19466 (N_19466,N_4729,N_6383);
nand U19467 (N_19467,N_989,N_4109);
nand U19468 (N_19468,N_1391,N_1754);
nand U19469 (N_19469,N_1530,N_547);
nor U19470 (N_19470,N_2736,N_6285);
nand U19471 (N_19471,N_7957,N_2319);
nand U19472 (N_19472,N_9272,N_9415);
nand U19473 (N_19473,N_6861,N_3664);
and U19474 (N_19474,N_8219,N_595);
or U19475 (N_19475,N_6090,N_154);
and U19476 (N_19476,N_5215,N_2933);
and U19477 (N_19477,N_7352,N_3154);
nand U19478 (N_19478,N_5006,N_8199);
nor U19479 (N_19479,N_1559,N_9349);
and U19480 (N_19480,N_8843,N_7834);
nand U19481 (N_19481,N_728,N_1872);
nor U19482 (N_19482,N_5567,N_4107);
xor U19483 (N_19483,N_4634,N_5033);
nor U19484 (N_19484,N_1274,N_1642);
nor U19485 (N_19485,N_2410,N_2548);
or U19486 (N_19486,N_8276,N_4635);
xor U19487 (N_19487,N_9440,N_3252);
nand U19488 (N_19488,N_7341,N_9489);
nand U19489 (N_19489,N_6827,N_921);
xnor U19490 (N_19490,N_2707,N_9421);
nand U19491 (N_19491,N_3837,N_7986);
nand U19492 (N_19492,N_5428,N_99);
or U19493 (N_19493,N_1881,N_6577);
nor U19494 (N_19494,N_7702,N_2894);
xnor U19495 (N_19495,N_3919,N_4811);
nor U19496 (N_19496,N_4411,N_4767);
and U19497 (N_19497,N_1960,N_9850);
or U19498 (N_19498,N_7008,N_1011);
xnor U19499 (N_19499,N_5024,N_6735);
xnor U19500 (N_19500,N_2366,N_5286);
and U19501 (N_19501,N_562,N_7417);
xnor U19502 (N_19502,N_686,N_4509);
nand U19503 (N_19503,N_713,N_1185);
or U19504 (N_19504,N_8986,N_3336);
or U19505 (N_19505,N_1411,N_1015);
and U19506 (N_19506,N_4482,N_6603);
or U19507 (N_19507,N_4249,N_4353);
nor U19508 (N_19508,N_2368,N_6954);
nand U19509 (N_19509,N_7966,N_6711);
nand U19510 (N_19510,N_1518,N_6427);
nand U19511 (N_19511,N_8213,N_6309);
nand U19512 (N_19512,N_3770,N_9571);
nand U19513 (N_19513,N_3081,N_6562);
or U19514 (N_19514,N_2788,N_3638);
xnor U19515 (N_19515,N_2642,N_9180);
nand U19516 (N_19516,N_9446,N_5638);
xor U19517 (N_19517,N_9255,N_649);
or U19518 (N_19518,N_2370,N_1137);
or U19519 (N_19519,N_3750,N_5);
or U19520 (N_19520,N_2828,N_891);
nor U19521 (N_19521,N_3370,N_684);
and U19522 (N_19522,N_3965,N_1837);
nor U19523 (N_19523,N_1156,N_4085);
or U19524 (N_19524,N_5392,N_9580);
xnor U19525 (N_19525,N_206,N_2030);
nand U19526 (N_19526,N_3770,N_4726);
nor U19527 (N_19527,N_2818,N_5698);
nor U19528 (N_19528,N_3285,N_4492);
and U19529 (N_19529,N_9383,N_9292);
nand U19530 (N_19530,N_1969,N_7399);
nand U19531 (N_19531,N_1644,N_4357);
or U19532 (N_19532,N_7461,N_9972);
and U19533 (N_19533,N_787,N_2535);
and U19534 (N_19534,N_6990,N_4045);
xnor U19535 (N_19535,N_7837,N_255);
xnor U19536 (N_19536,N_4430,N_7235);
xor U19537 (N_19537,N_1763,N_4180);
and U19538 (N_19538,N_9650,N_9420);
and U19539 (N_19539,N_5392,N_4408);
and U19540 (N_19540,N_1963,N_4143);
nand U19541 (N_19541,N_7884,N_2399);
nor U19542 (N_19542,N_5832,N_3493);
xnor U19543 (N_19543,N_3657,N_5819);
xor U19544 (N_19544,N_2585,N_5070);
xnor U19545 (N_19545,N_4814,N_4319);
xnor U19546 (N_19546,N_4795,N_4036);
and U19547 (N_19547,N_802,N_6100);
or U19548 (N_19548,N_9091,N_5861);
and U19549 (N_19549,N_2384,N_3020);
or U19550 (N_19550,N_2985,N_8552);
and U19551 (N_19551,N_2439,N_3930);
xor U19552 (N_19552,N_1971,N_4669);
or U19553 (N_19553,N_4769,N_3065);
nand U19554 (N_19554,N_5908,N_790);
nor U19555 (N_19555,N_1775,N_7282);
nand U19556 (N_19556,N_8013,N_8918);
or U19557 (N_19557,N_5867,N_8713);
or U19558 (N_19558,N_3743,N_9877);
nand U19559 (N_19559,N_2069,N_6570);
nor U19560 (N_19560,N_2060,N_8098);
xor U19561 (N_19561,N_8719,N_7297);
and U19562 (N_19562,N_2250,N_7138);
nand U19563 (N_19563,N_9767,N_1964);
nor U19564 (N_19564,N_5264,N_1347);
xnor U19565 (N_19565,N_9469,N_6098);
nor U19566 (N_19566,N_1586,N_5203);
xnor U19567 (N_19567,N_8641,N_5930);
nor U19568 (N_19568,N_3572,N_955);
and U19569 (N_19569,N_3594,N_7207);
nand U19570 (N_19570,N_5820,N_7869);
and U19571 (N_19571,N_9619,N_1806);
or U19572 (N_19572,N_8713,N_3742);
and U19573 (N_19573,N_3747,N_3653);
nor U19574 (N_19574,N_3291,N_4744);
or U19575 (N_19575,N_242,N_7141);
or U19576 (N_19576,N_530,N_2756);
and U19577 (N_19577,N_3843,N_5868);
nand U19578 (N_19578,N_2459,N_9981);
nor U19579 (N_19579,N_2553,N_1592);
and U19580 (N_19580,N_8985,N_1035);
or U19581 (N_19581,N_9702,N_4984);
or U19582 (N_19582,N_4581,N_4892);
xnor U19583 (N_19583,N_5795,N_6488);
nand U19584 (N_19584,N_1723,N_2415);
nand U19585 (N_19585,N_1354,N_1506);
or U19586 (N_19586,N_3213,N_3586);
and U19587 (N_19587,N_3662,N_6921);
nor U19588 (N_19588,N_2498,N_1554);
or U19589 (N_19589,N_3645,N_33);
nor U19590 (N_19590,N_6186,N_9732);
xnor U19591 (N_19591,N_8721,N_8657);
or U19592 (N_19592,N_2754,N_5439);
or U19593 (N_19593,N_2425,N_4355);
nor U19594 (N_19594,N_4128,N_1013);
nor U19595 (N_19595,N_9482,N_6549);
and U19596 (N_19596,N_8221,N_1677);
and U19597 (N_19597,N_7152,N_6965);
xnor U19598 (N_19598,N_1347,N_7997);
nor U19599 (N_19599,N_5443,N_5819);
nand U19600 (N_19600,N_1565,N_5154);
nand U19601 (N_19601,N_6178,N_8530);
or U19602 (N_19602,N_2846,N_3270);
and U19603 (N_19603,N_3401,N_7153);
nand U19604 (N_19604,N_4013,N_8193);
or U19605 (N_19605,N_8258,N_1103);
and U19606 (N_19606,N_6677,N_4188);
and U19607 (N_19607,N_9546,N_9840);
nor U19608 (N_19608,N_8479,N_7215);
nand U19609 (N_19609,N_3289,N_8163);
xor U19610 (N_19610,N_5233,N_6713);
and U19611 (N_19611,N_2136,N_6007);
xor U19612 (N_19612,N_9205,N_4335);
and U19613 (N_19613,N_9144,N_1793);
nand U19614 (N_19614,N_6481,N_4554);
and U19615 (N_19615,N_9488,N_8223);
or U19616 (N_19616,N_1311,N_5764);
and U19617 (N_19617,N_7888,N_2179);
nand U19618 (N_19618,N_1927,N_8185);
or U19619 (N_19619,N_1453,N_1555);
xnor U19620 (N_19620,N_5102,N_8187);
nor U19621 (N_19621,N_1207,N_1922);
nand U19622 (N_19622,N_8935,N_8132);
nand U19623 (N_19623,N_2315,N_8494);
nor U19624 (N_19624,N_3851,N_8362);
nand U19625 (N_19625,N_3217,N_9322);
and U19626 (N_19626,N_2600,N_5865);
nand U19627 (N_19627,N_8397,N_8382);
or U19628 (N_19628,N_7866,N_4790);
nand U19629 (N_19629,N_6390,N_1233);
and U19630 (N_19630,N_8520,N_6228);
and U19631 (N_19631,N_9406,N_6156);
xnor U19632 (N_19632,N_145,N_7782);
or U19633 (N_19633,N_8075,N_6231);
and U19634 (N_19634,N_5675,N_8504);
xnor U19635 (N_19635,N_4480,N_9916);
xor U19636 (N_19636,N_4779,N_1982);
nand U19637 (N_19637,N_8715,N_9501);
or U19638 (N_19638,N_2623,N_1015);
and U19639 (N_19639,N_4914,N_7707);
nor U19640 (N_19640,N_9393,N_2896);
and U19641 (N_19641,N_7500,N_7225);
xor U19642 (N_19642,N_789,N_6061);
nor U19643 (N_19643,N_7271,N_7585);
nor U19644 (N_19644,N_7665,N_4145);
nor U19645 (N_19645,N_1522,N_7225);
nor U19646 (N_19646,N_8723,N_8690);
and U19647 (N_19647,N_3586,N_4348);
or U19648 (N_19648,N_6216,N_6431);
nand U19649 (N_19649,N_775,N_3210);
or U19650 (N_19650,N_1357,N_5174);
xnor U19651 (N_19651,N_8742,N_1252);
and U19652 (N_19652,N_2500,N_2876);
or U19653 (N_19653,N_7482,N_4722);
xnor U19654 (N_19654,N_6244,N_9490);
nor U19655 (N_19655,N_6781,N_5489);
nand U19656 (N_19656,N_3238,N_9937);
xor U19657 (N_19657,N_1112,N_8688);
or U19658 (N_19658,N_5908,N_334);
xnor U19659 (N_19659,N_9695,N_227);
nand U19660 (N_19660,N_7524,N_3377);
nor U19661 (N_19661,N_6047,N_3571);
or U19662 (N_19662,N_1148,N_8731);
nor U19663 (N_19663,N_3323,N_8162);
xnor U19664 (N_19664,N_7532,N_3533);
xor U19665 (N_19665,N_4834,N_6886);
or U19666 (N_19666,N_228,N_8847);
or U19667 (N_19667,N_6167,N_7285);
or U19668 (N_19668,N_9975,N_5028);
nand U19669 (N_19669,N_867,N_9942);
or U19670 (N_19670,N_7214,N_6200);
nand U19671 (N_19671,N_2634,N_6659);
and U19672 (N_19672,N_6312,N_1919);
nor U19673 (N_19673,N_7010,N_117);
and U19674 (N_19674,N_3543,N_2022);
xnor U19675 (N_19675,N_5143,N_3510);
nor U19676 (N_19676,N_2387,N_8754);
and U19677 (N_19677,N_1503,N_1302);
nand U19678 (N_19678,N_897,N_2698);
and U19679 (N_19679,N_1857,N_3283);
nor U19680 (N_19680,N_1552,N_8693);
nor U19681 (N_19681,N_9891,N_8348);
nand U19682 (N_19682,N_6182,N_481);
or U19683 (N_19683,N_6935,N_76);
nor U19684 (N_19684,N_8271,N_101);
nor U19685 (N_19685,N_6625,N_8369);
nor U19686 (N_19686,N_2244,N_9129);
or U19687 (N_19687,N_8931,N_8621);
xor U19688 (N_19688,N_6002,N_5175);
nor U19689 (N_19689,N_8648,N_1512);
nand U19690 (N_19690,N_5745,N_163);
or U19691 (N_19691,N_984,N_9898);
nand U19692 (N_19692,N_9547,N_9710);
nor U19693 (N_19693,N_6470,N_8605);
xor U19694 (N_19694,N_428,N_3819);
nor U19695 (N_19695,N_5611,N_2124);
nor U19696 (N_19696,N_4350,N_4104);
nand U19697 (N_19697,N_9604,N_3015);
nand U19698 (N_19698,N_447,N_4325);
and U19699 (N_19699,N_5446,N_2013);
nor U19700 (N_19700,N_5629,N_9365);
xor U19701 (N_19701,N_7293,N_3792);
nand U19702 (N_19702,N_249,N_2546);
or U19703 (N_19703,N_2680,N_1956);
nor U19704 (N_19704,N_7691,N_3352);
nor U19705 (N_19705,N_8123,N_3926);
xor U19706 (N_19706,N_2485,N_9291);
nand U19707 (N_19707,N_9504,N_4131);
and U19708 (N_19708,N_7120,N_8426);
nand U19709 (N_19709,N_4684,N_729);
nor U19710 (N_19710,N_8001,N_564);
xnor U19711 (N_19711,N_7986,N_8710);
nor U19712 (N_19712,N_134,N_6817);
and U19713 (N_19713,N_3643,N_4328);
xor U19714 (N_19714,N_1912,N_9286);
nand U19715 (N_19715,N_9720,N_4264);
xnor U19716 (N_19716,N_3758,N_9916);
xor U19717 (N_19717,N_3424,N_9888);
or U19718 (N_19718,N_456,N_5799);
or U19719 (N_19719,N_2006,N_6721);
xor U19720 (N_19720,N_3222,N_4060);
nand U19721 (N_19721,N_3666,N_2426);
and U19722 (N_19722,N_5320,N_7427);
nor U19723 (N_19723,N_9976,N_5297);
xor U19724 (N_19724,N_9056,N_4536);
and U19725 (N_19725,N_9919,N_3068);
xnor U19726 (N_19726,N_1934,N_4893);
and U19727 (N_19727,N_1393,N_6255);
and U19728 (N_19728,N_8234,N_657);
nand U19729 (N_19729,N_1757,N_3222);
nor U19730 (N_19730,N_5994,N_8836);
or U19731 (N_19731,N_8699,N_6609);
or U19732 (N_19732,N_657,N_8093);
xor U19733 (N_19733,N_156,N_2475);
and U19734 (N_19734,N_896,N_7878);
or U19735 (N_19735,N_5212,N_6028);
or U19736 (N_19736,N_5746,N_9504);
or U19737 (N_19737,N_3780,N_7929);
or U19738 (N_19738,N_723,N_3710);
nand U19739 (N_19739,N_3256,N_9678);
nand U19740 (N_19740,N_685,N_7795);
or U19741 (N_19741,N_2899,N_7908);
and U19742 (N_19742,N_3197,N_16);
and U19743 (N_19743,N_8253,N_8165);
or U19744 (N_19744,N_9353,N_2641);
and U19745 (N_19745,N_1809,N_4783);
nor U19746 (N_19746,N_8603,N_8509);
nand U19747 (N_19747,N_3629,N_2542);
xor U19748 (N_19748,N_3235,N_9416);
nand U19749 (N_19749,N_1431,N_1829);
and U19750 (N_19750,N_4306,N_4006);
nand U19751 (N_19751,N_9254,N_1489);
or U19752 (N_19752,N_3660,N_3165);
and U19753 (N_19753,N_7396,N_9613);
nor U19754 (N_19754,N_1150,N_7709);
xor U19755 (N_19755,N_3518,N_2541);
xnor U19756 (N_19756,N_4482,N_7137);
nand U19757 (N_19757,N_2217,N_7881);
and U19758 (N_19758,N_1035,N_7420);
nor U19759 (N_19759,N_6420,N_9991);
nor U19760 (N_19760,N_8145,N_8409);
nand U19761 (N_19761,N_1805,N_5930);
nor U19762 (N_19762,N_4309,N_6163);
nor U19763 (N_19763,N_820,N_4228);
nand U19764 (N_19764,N_3104,N_2000);
nand U19765 (N_19765,N_7773,N_1551);
nor U19766 (N_19766,N_8927,N_5022);
xnor U19767 (N_19767,N_4884,N_2003);
and U19768 (N_19768,N_9227,N_8423);
xnor U19769 (N_19769,N_8185,N_4599);
or U19770 (N_19770,N_558,N_2199);
nor U19771 (N_19771,N_7682,N_4149);
nand U19772 (N_19772,N_9399,N_3184);
nand U19773 (N_19773,N_7058,N_7161);
nand U19774 (N_19774,N_3922,N_8284);
nand U19775 (N_19775,N_9050,N_4580);
xnor U19776 (N_19776,N_6265,N_9846);
nor U19777 (N_19777,N_5232,N_2395);
nand U19778 (N_19778,N_7832,N_3047);
and U19779 (N_19779,N_754,N_5326);
nand U19780 (N_19780,N_658,N_7016);
xnor U19781 (N_19781,N_6602,N_5276);
and U19782 (N_19782,N_2110,N_4303);
nand U19783 (N_19783,N_2133,N_6321);
or U19784 (N_19784,N_6836,N_6739);
nor U19785 (N_19785,N_815,N_702);
nor U19786 (N_19786,N_8174,N_1094);
or U19787 (N_19787,N_2431,N_9178);
or U19788 (N_19788,N_7840,N_445);
or U19789 (N_19789,N_6649,N_2286);
nand U19790 (N_19790,N_4404,N_8781);
nor U19791 (N_19791,N_1664,N_6285);
xnor U19792 (N_19792,N_9108,N_5844);
and U19793 (N_19793,N_6405,N_776);
xor U19794 (N_19794,N_9634,N_8221);
xor U19795 (N_19795,N_9855,N_8882);
nand U19796 (N_19796,N_6902,N_8067);
nand U19797 (N_19797,N_1709,N_8281);
nand U19798 (N_19798,N_6442,N_9195);
nand U19799 (N_19799,N_4094,N_5800);
xnor U19800 (N_19800,N_4283,N_7563);
xor U19801 (N_19801,N_1013,N_3850);
and U19802 (N_19802,N_2110,N_710);
and U19803 (N_19803,N_8240,N_9056);
nand U19804 (N_19804,N_7576,N_4583);
nand U19805 (N_19805,N_5132,N_8878);
or U19806 (N_19806,N_9104,N_9121);
and U19807 (N_19807,N_7328,N_764);
xor U19808 (N_19808,N_7921,N_3135);
xor U19809 (N_19809,N_5859,N_1509);
and U19810 (N_19810,N_5618,N_7017);
xnor U19811 (N_19811,N_3856,N_6050);
and U19812 (N_19812,N_2173,N_4561);
nor U19813 (N_19813,N_1342,N_7852);
and U19814 (N_19814,N_8645,N_7100);
or U19815 (N_19815,N_238,N_8132);
or U19816 (N_19816,N_7514,N_2846);
nand U19817 (N_19817,N_2438,N_2373);
and U19818 (N_19818,N_5653,N_6906);
xnor U19819 (N_19819,N_8851,N_8560);
or U19820 (N_19820,N_722,N_7637);
and U19821 (N_19821,N_4570,N_2029);
nand U19822 (N_19822,N_5005,N_885);
and U19823 (N_19823,N_4332,N_5066);
xnor U19824 (N_19824,N_5597,N_5861);
nand U19825 (N_19825,N_8077,N_3922);
xnor U19826 (N_19826,N_4647,N_1995);
nor U19827 (N_19827,N_1767,N_4814);
nor U19828 (N_19828,N_9862,N_8178);
and U19829 (N_19829,N_3088,N_8385);
and U19830 (N_19830,N_2362,N_2658);
xor U19831 (N_19831,N_6429,N_3528);
and U19832 (N_19832,N_8987,N_1188);
nor U19833 (N_19833,N_1724,N_6040);
and U19834 (N_19834,N_8084,N_4848);
xor U19835 (N_19835,N_3506,N_4029);
nand U19836 (N_19836,N_5093,N_7508);
and U19837 (N_19837,N_4430,N_2563);
xor U19838 (N_19838,N_1802,N_191);
nand U19839 (N_19839,N_3072,N_7483);
nand U19840 (N_19840,N_1081,N_5164);
nor U19841 (N_19841,N_3482,N_878);
xor U19842 (N_19842,N_5269,N_1981);
and U19843 (N_19843,N_5546,N_6297);
nor U19844 (N_19844,N_6678,N_9025);
nor U19845 (N_19845,N_9139,N_7763);
nor U19846 (N_19846,N_8746,N_7075);
nand U19847 (N_19847,N_8877,N_6880);
nand U19848 (N_19848,N_3863,N_2497);
xnor U19849 (N_19849,N_3133,N_6901);
nor U19850 (N_19850,N_8962,N_9125);
and U19851 (N_19851,N_6917,N_6362);
nor U19852 (N_19852,N_1114,N_6631);
nor U19853 (N_19853,N_5958,N_335);
nor U19854 (N_19854,N_4719,N_2018);
nand U19855 (N_19855,N_9433,N_9462);
or U19856 (N_19856,N_4096,N_1002);
and U19857 (N_19857,N_6335,N_6385);
xor U19858 (N_19858,N_6587,N_5351);
nor U19859 (N_19859,N_2380,N_6991);
or U19860 (N_19860,N_8198,N_4901);
xor U19861 (N_19861,N_6689,N_8457);
nor U19862 (N_19862,N_1210,N_2457);
or U19863 (N_19863,N_6002,N_1531);
and U19864 (N_19864,N_9916,N_3160);
xnor U19865 (N_19865,N_8690,N_9440);
and U19866 (N_19866,N_7613,N_2694);
xor U19867 (N_19867,N_5438,N_5684);
nand U19868 (N_19868,N_5044,N_5805);
or U19869 (N_19869,N_538,N_8815);
nand U19870 (N_19870,N_9743,N_1988);
and U19871 (N_19871,N_8544,N_4974);
xor U19872 (N_19872,N_1437,N_720);
nand U19873 (N_19873,N_6915,N_1837);
nand U19874 (N_19874,N_4938,N_2257);
xnor U19875 (N_19875,N_3100,N_9271);
and U19876 (N_19876,N_7322,N_5136);
nand U19877 (N_19877,N_658,N_9077);
nand U19878 (N_19878,N_5008,N_7416);
nand U19879 (N_19879,N_9041,N_2067);
nand U19880 (N_19880,N_3057,N_6236);
nor U19881 (N_19881,N_8057,N_8175);
nor U19882 (N_19882,N_6944,N_7704);
xor U19883 (N_19883,N_7302,N_1144);
nand U19884 (N_19884,N_5271,N_2429);
and U19885 (N_19885,N_7469,N_2599);
nand U19886 (N_19886,N_6410,N_4927);
or U19887 (N_19887,N_950,N_2982);
nor U19888 (N_19888,N_7941,N_9774);
xnor U19889 (N_19889,N_5680,N_1777);
or U19890 (N_19890,N_4382,N_5410);
and U19891 (N_19891,N_671,N_9749);
nor U19892 (N_19892,N_8008,N_9358);
and U19893 (N_19893,N_4,N_2643);
nand U19894 (N_19894,N_8856,N_1557);
nor U19895 (N_19895,N_752,N_1396);
nand U19896 (N_19896,N_4404,N_5318);
nor U19897 (N_19897,N_7380,N_8561);
nand U19898 (N_19898,N_8056,N_7184);
and U19899 (N_19899,N_2815,N_416);
nand U19900 (N_19900,N_4797,N_4309);
xor U19901 (N_19901,N_4745,N_4704);
nor U19902 (N_19902,N_1247,N_7204);
nor U19903 (N_19903,N_6099,N_5827);
or U19904 (N_19904,N_520,N_2092);
nor U19905 (N_19905,N_9676,N_5467);
or U19906 (N_19906,N_518,N_5467);
nand U19907 (N_19907,N_8794,N_3170);
nor U19908 (N_19908,N_4434,N_3164);
nor U19909 (N_19909,N_1887,N_5598);
and U19910 (N_19910,N_3245,N_2276);
nor U19911 (N_19911,N_855,N_6996);
and U19912 (N_19912,N_4432,N_4592);
nor U19913 (N_19913,N_5042,N_5828);
nand U19914 (N_19914,N_8266,N_3451);
and U19915 (N_19915,N_3065,N_3139);
and U19916 (N_19916,N_9439,N_2801);
xnor U19917 (N_19917,N_441,N_5083);
and U19918 (N_19918,N_21,N_7675);
nor U19919 (N_19919,N_5063,N_7365);
nand U19920 (N_19920,N_979,N_92);
nand U19921 (N_19921,N_1696,N_2378);
xnor U19922 (N_19922,N_3437,N_1289);
or U19923 (N_19923,N_5679,N_5333);
nor U19924 (N_19924,N_2543,N_3480);
xor U19925 (N_19925,N_1567,N_8890);
xor U19926 (N_19926,N_5514,N_3223);
nand U19927 (N_19927,N_9235,N_638);
or U19928 (N_19928,N_2023,N_3754);
nor U19929 (N_19929,N_5856,N_1795);
and U19930 (N_19930,N_8633,N_8104);
xor U19931 (N_19931,N_9660,N_7141);
and U19932 (N_19932,N_1710,N_4661);
and U19933 (N_19933,N_4109,N_6543);
and U19934 (N_19934,N_5980,N_9200);
xor U19935 (N_19935,N_4031,N_9013);
and U19936 (N_19936,N_2511,N_6593);
or U19937 (N_19937,N_4310,N_6138);
nor U19938 (N_19938,N_3470,N_7040);
or U19939 (N_19939,N_7565,N_2531);
nor U19940 (N_19940,N_9014,N_8471);
nor U19941 (N_19941,N_50,N_4532);
xnor U19942 (N_19942,N_936,N_9030);
xnor U19943 (N_19943,N_1009,N_3676);
xor U19944 (N_19944,N_2921,N_2988);
nand U19945 (N_19945,N_5350,N_5252);
nand U19946 (N_19946,N_6074,N_5457);
xnor U19947 (N_19947,N_4988,N_824);
and U19948 (N_19948,N_896,N_6035);
nand U19949 (N_19949,N_9356,N_9668);
and U19950 (N_19950,N_7950,N_3989);
nand U19951 (N_19951,N_9546,N_9291);
nand U19952 (N_19952,N_4672,N_8913);
and U19953 (N_19953,N_5892,N_899);
xnor U19954 (N_19954,N_7063,N_8325);
and U19955 (N_19955,N_4408,N_4963);
xnor U19956 (N_19956,N_9369,N_6613);
or U19957 (N_19957,N_6779,N_8253);
and U19958 (N_19958,N_6442,N_6358);
and U19959 (N_19959,N_3615,N_7738);
xnor U19960 (N_19960,N_1321,N_850);
and U19961 (N_19961,N_4706,N_9146);
xor U19962 (N_19962,N_7458,N_2723);
nand U19963 (N_19963,N_9519,N_166);
xnor U19964 (N_19964,N_8228,N_1834);
xor U19965 (N_19965,N_4678,N_2936);
nor U19966 (N_19966,N_9745,N_9749);
or U19967 (N_19967,N_6953,N_8511);
nor U19968 (N_19968,N_3196,N_8336);
and U19969 (N_19969,N_2572,N_526);
and U19970 (N_19970,N_7813,N_3475);
nand U19971 (N_19971,N_6512,N_5877);
and U19972 (N_19972,N_8481,N_5299);
and U19973 (N_19973,N_4480,N_5090);
and U19974 (N_19974,N_9329,N_1099);
and U19975 (N_19975,N_9524,N_3990);
xor U19976 (N_19976,N_4500,N_3030);
and U19977 (N_19977,N_9405,N_2367);
nand U19978 (N_19978,N_248,N_1643);
nand U19979 (N_19979,N_9312,N_5696);
nand U19980 (N_19980,N_6661,N_3996);
and U19981 (N_19981,N_7166,N_4652);
nor U19982 (N_19982,N_1150,N_7485);
xor U19983 (N_19983,N_6616,N_2949);
nor U19984 (N_19984,N_5100,N_6483);
or U19985 (N_19985,N_8823,N_7987);
nand U19986 (N_19986,N_6540,N_4536);
xor U19987 (N_19987,N_9641,N_6804);
xor U19988 (N_19988,N_9896,N_8010);
or U19989 (N_19989,N_5528,N_4354);
xnor U19990 (N_19990,N_8629,N_8718);
nor U19991 (N_19991,N_9927,N_8083);
or U19992 (N_19992,N_3408,N_3249);
and U19993 (N_19993,N_4044,N_3535);
xor U19994 (N_19994,N_8167,N_8621);
nor U19995 (N_19995,N_2765,N_6043);
xnor U19996 (N_19996,N_9515,N_3795);
xnor U19997 (N_19997,N_1467,N_64);
or U19998 (N_19998,N_9613,N_8343);
or U19999 (N_19999,N_5521,N_5324);
and U20000 (N_20000,N_18848,N_15375);
xor U20001 (N_20001,N_15521,N_13624);
or U20002 (N_20002,N_10044,N_18607);
and U20003 (N_20003,N_15263,N_13856);
or U20004 (N_20004,N_12290,N_19998);
xor U20005 (N_20005,N_10089,N_16644);
nand U20006 (N_20006,N_19419,N_11130);
nor U20007 (N_20007,N_13467,N_10333);
xnor U20008 (N_20008,N_19296,N_18686);
xor U20009 (N_20009,N_14025,N_10829);
and U20010 (N_20010,N_13562,N_16455);
xnor U20011 (N_20011,N_14421,N_13530);
nor U20012 (N_20012,N_13379,N_19269);
xnor U20013 (N_20013,N_10518,N_13312);
nand U20014 (N_20014,N_18498,N_10175);
nand U20015 (N_20015,N_17788,N_19765);
and U20016 (N_20016,N_14053,N_10011);
xnor U20017 (N_20017,N_14510,N_14165);
and U20018 (N_20018,N_14909,N_19201);
or U20019 (N_20019,N_11108,N_12618);
or U20020 (N_20020,N_18541,N_16888);
xor U20021 (N_20021,N_11372,N_15420);
xor U20022 (N_20022,N_11453,N_18101);
or U20023 (N_20023,N_18378,N_10022);
xnor U20024 (N_20024,N_10894,N_10784);
and U20025 (N_20025,N_12366,N_12992);
nand U20026 (N_20026,N_19508,N_10657);
and U20027 (N_20027,N_19217,N_17275);
and U20028 (N_20028,N_13577,N_16034);
xor U20029 (N_20029,N_10016,N_16614);
or U20030 (N_20030,N_15585,N_19443);
nor U20031 (N_20031,N_14580,N_15247);
xor U20032 (N_20032,N_15900,N_18871);
nand U20033 (N_20033,N_19152,N_14584);
xnor U20034 (N_20034,N_17768,N_14319);
nor U20035 (N_20035,N_18055,N_17205);
or U20036 (N_20036,N_13987,N_11471);
or U20037 (N_20037,N_15135,N_14862);
nor U20038 (N_20038,N_13043,N_16787);
and U20039 (N_20039,N_13405,N_19773);
xnor U20040 (N_20040,N_17847,N_16178);
or U20041 (N_20041,N_14291,N_13186);
nand U20042 (N_20042,N_12873,N_11807);
nand U20043 (N_20043,N_17649,N_17490);
nor U20044 (N_20044,N_13414,N_19386);
xor U20045 (N_20045,N_13035,N_12509);
or U20046 (N_20046,N_11623,N_14920);
or U20047 (N_20047,N_17307,N_19602);
and U20048 (N_20048,N_12317,N_18641);
and U20049 (N_20049,N_12904,N_12253);
xor U20050 (N_20050,N_13171,N_19367);
and U20051 (N_20051,N_15362,N_12938);
nor U20052 (N_20052,N_13950,N_12976);
nor U20053 (N_20053,N_18954,N_10469);
nand U20054 (N_20054,N_17338,N_17744);
nand U20055 (N_20055,N_10420,N_10500);
nor U20056 (N_20056,N_18271,N_10755);
or U20057 (N_20057,N_17472,N_14570);
and U20058 (N_20058,N_11451,N_19830);
nand U20059 (N_20059,N_15041,N_19319);
nand U20060 (N_20060,N_13773,N_10931);
and U20061 (N_20061,N_11088,N_14576);
xnor U20062 (N_20062,N_13589,N_18391);
nand U20063 (N_20063,N_18643,N_16198);
nor U20064 (N_20064,N_14978,N_18792);
nor U20065 (N_20065,N_13462,N_19637);
and U20066 (N_20066,N_14710,N_19513);
and U20067 (N_20067,N_17745,N_18885);
and U20068 (N_20068,N_12959,N_13311);
nand U20069 (N_20069,N_19060,N_10691);
xor U20070 (N_20070,N_10260,N_17132);
and U20071 (N_20071,N_16006,N_11027);
nand U20072 (N_20072,N_17729,N_18809);
nand U20073 (N_20073,N_15191,N_11485);
nand U20074 (N_20074,N_16810,N_13585);
nand U20075 (N_20075,N_11004,N_11581);
or U20076 (N_20076,N_10320,N_15818);
nor U20077 (N_20077,N_16633,N_15566);
or U20078 (N_20078,N_13072,N_18382);
nand U20079 (N_20079,N_18236,N_16463);
xnor U20080 (N_20080,N_19091,N_11072);
nor U20081 (N_20081,N_16871,N_16691);
nor U20082 (N_20082,N_13803,N_13018);
and U20083 (N_20083,N_15483,N_10674);
or U20084 (N_20084,N_10009,N_17262);
xnor U20085 (N_20085,N_12206,N_11102);
nand U20086 (N_20086,N_11111,N_19702);
and U20087 (N_20087,N_19487,N_12002);
nand U20088 (N_20088,N_12439,N_19234);
xnor U20089 (N_20089,N_19591,N_18093);
nand U20090 (N_20090,N_18937,N_16383);
and U20091 (N_20091,N_11860,N_18366);
nor U20092 (N_20092,N_13274,N_15810);
nor U20093 (N_20093,N_18152,N_10813);
or U20094 (N_20094,N_18808,N_13886);
nand U20095 (N_20095,N_10986,N_19354);
xnor U20096 (N_20096,N_10872,N_18026);
nor U20097 (N_20097,N_17356,N_18276);
nand U20098 (N_20098,N_15581,N_18802);
nand U20099 (N_20099,N_19992,N_17207);
or U20100 (N_20100,N_10082,N_18274);
xnor U20101 (N_20101,N_15685,N_13353);
nor U20102 (N_20102,N_17754,N_19155);
and U20103 (N_20103,N_11517,N_15291);
or U20104 (N_20104,N_14480,N_16983);
nand U20105 (N_20105,N_12636,N_16379);
nand U20106 (N_20106,N_13871,N_11913);
xnor U20107 (N_20107,N_12321,N_16547);
and U20108 (N_20108,N_19633,N_19696);
xnor U20109 (N_20109,N_13255,N_14339);
xnor U20110 (N_20110,N_15609,N_19608);
or U20111 (N_20111,N_12149,N_12764);
or U20112 (N_20112,N_16853,N_13867);
or U20113 (N_20113,N_11985,N_13791);
and U20114 (N_20114,N_14342,N_17229);
nand U20115 (N_20115,N_10882,N_13744);
or U20116 (N_20116,N_15535,N_18151);
and U20117 (N_20117,N_17198,N_10847);
xor U20118 (N_20118,N_10771,N_19105);
or U20119 (N_20119,N_13512,N_11405);
nand U20120 (N_20120,N_10144,N_14756);
or U20121 (N_20121,N_15804,N_18009);
xor U20122 (N_20122,N_19982,N_10358);
nand U20123 (N_20123,N_11957,N_12405);
nor U20124 (N_20124,N_15542,N_12041);
nand U20125 (N_20125,N_12586,N_11119);
and U20126 (N_20126,N_17365,N_12255);
and U20127 (N_20127,N_12358,N_15207);
nor U20128 (N_20128,N_11177,N_17871);
or U20129 (N_20129,N_16799,N_16013);
nor U20130 (N_20130,N_10249,N_11916);
xnor U20131 (N_20131,N_19022,N_17054);
nor U20132 (N_20132,N_19940,N_14378);
or U20133 (N_20133,N_14937,N_16084);
xnor U20134 (N_20134,N_13842,N_12660);
nor U20135 (N_20135,N_18963,N_19870);
nand U20136 (N_20136,N_11971,N_10529);
nand U20137 (N_20137,N_11840,N_15443);
xor U20138 (N_20138,N_17656,N_12663);
and U20139 (N_20139,N_11235,N_19810);
and U20140 (N_20140,N_11513,N_18086);
nor U20141 (N_20141,N_19483,N_12236);
and U20142 (N_20142,N_12156,N_15619);
nor U20143 (N_20143,N_17727,N_16385);
and U20144 (N_20144,N_15402,N_19016);
or U20145 (N_20145,N_16228,N_11995);
or U20146 (N_20146,N_15596,N_15989);
nand U20147 (N_20147,N_16591,N_18278);
nor U20148 (N_20148,N_12784,N_19154);
xnor U20149 (N_20149,N_17520,N_14672);
and U20150 (N_20150,N_11690,N_14059);
nand U20151 (N_20151,N_16821,N_19262);
and U20152 (N_20152,N_17920,N_15767);
nand U20153 (N_20153,N_17936,N_14405);
xor U20154 (N_20154,N_12843,N_14693);
or U20155 (N_20155,N_15532,N_12188);
nor U20156 (N_20156,N_18570,N_13696);
nor U20157 (N_20157,N_13887,N_18080);
xor U20158 (N_20158,N_16457,N_13317);
xnor U20159 (N_20159,N_10487,N_14435);
nand U20160 (N_20160,N_14821,N_15725);
or U20161 (N_20161,N_12883,N_12258);
nor U20162 (N_20162,N_14316,N_19576);
and U20163 (N_20163,N_12563,N_10719);
nor U20164 (N_20164,N_17769,N_10941);
xnor U20165 (N_20165,N_18175,N_18129);
nand U20166 (N_20166,N_16253,N_10522);
nand U20167 (N_20167,N_15719,N_18784);
and U20168 (N_20168,N_13592,N_13559);
and U20169 (N_20169,N_10241,N_15370);
nor U20170 (N_20170,N_16890,N_11564);
or U20171 (N_20171,N_10593,N_15478);
xnor U20172 (N_20172,N_16265,N_19132);
or U20173 (N_20173,N_15755,N_10669);
nand U20174 (N_20174,N_19281,N_10770);
or U20175 (N_20175,N_13646,N_14958);
nor U20176 (N_20176,N_11773,N_13799);
and U20177 (N_20177,N_10666,N_10966);
xnor U20178 (N_20178,N_16128,N_15228);
or U20179 (N_20179,N_17455,N_19212);
and U20180 (N_20180,N_13970,N_15788);
and U20181 (N_20181,N_19037,N_12845);
or U20182 (N_20182,N_18311,N_13385);
xnor U20183 (N_20183,N_12034,N_15357);
and U20184 (N_20184,N_15882,N_10468);
nand U20185 (N_20185,N_19561,N_12497);
and U20186 (N_20186,N_19975,N_18838);
nor U20187 (N_20187,N_17879,N_13941);
and U20188 (N_20188,N_16293,N_13563);
nor U20189 (N_20189,N_19473,N_13541);
or U20190 (N_20190,N_19656,N_17381);
nand U20191 (N_20191,N_11988,N_16107);
or U20192 (N_20192,N_12861,N_11364);
nand U20193 (N_20193,N_10906,N_13925);
nand U20194 (N_20194,N_13805,N_13220);
nand U20195 (N_20195,N_17406,N_15242);
or U20196 (N_20196,N_11394,N_12640);
xor U20197 (N_20197,N_14562,N_18429);
and U20198 (N_20198,N_16192,N_14949);
nand U20199 (N_20199,N_15187,N_11450);
and U20200 (N_20200,N_12708,N_12713);
nor U20201 (N_20201,N_14599,N_19002);
nor U20202 (N_20202,N_14020,N_18662);
xor U20203 (N_20203,N_17679,N_19548);
and U20204 (N_20204,N_15143,N_13721);
nand U20205 (N_20205,N_10244,N_19424);
or U20206 (N_20206,N_13812,N_13611);
nand U20207 (N_20207,N_13239,N_16448);
xor U20208 (N_20208,N_11225,N_17096);
nor U20209 (N_20209,N_14335,N_12650);
xnor U20210 (N_20210,N_19965,N_14998);
or U20211 (N_20211,N_11932,N_12948);
and U20212 (N_20212,N_16584,N_10722);
nor U20213 (N_20213,N_15648,N_12858);
nor U20214 (N_20214,N_11839,N_15363);
xor U20215 (N_20215,N_17341,N_12593);
nand U20216 (N_20216,N_15970,N_16069);
and U20217 (N_20217,N_10887,N_15064);
nand U20218 (N_20218,N_16194,N_19138);
nor U20219 (N_20219,N_13675,N_15346);
or U20220 (N_20220,N_10866,N_19542);
or U20221 (N_20221,N_17439,N_11008);
or U20222 (N_20222,N_18901,N_12846);
nor U20223 (N_20223,N_13109,N_14670);
nand U20224 (N_20224,N_11866,N_16165);
nor U20225 (N_20225,N_12373,N_16273);
and U20226 (N_20226,N_12607,N_18824);
and U20227 (N_20227,N_13590,N_14747);
nand U20228 (N_20228,N_16921,N_14945);
nor U20229 (N_20229,N_19912,N_19874);
nor U20230 (N_20230,N_16943,N_12176);
and U20231 (N_20231,N_15917,N_10289);
xor U20232 (N_20232,N_12098,N_12595);
or U20233 (N_20233,N_11144,N_16312);
nor U20234 (N_20234,N_15372,N_15087);
and U20235 (N_20235,N_18102,N_18341);
nor U20236 (N_20236,N_15642,N_15728);
and U20237 (N_20237,N_14608,N_16226);
or U20238 (N_20238,N_18604,N_14509);
xor U20239 (N_20239,N_11469,N_15851);
or U20240 (N_20240,N_14057,N_19507);
nor U20241 (N_20241,N_15688,N_12322);
nor U20242 (N_20242,N_14241,N_11347);
nor U20243 (N_20243,N_11110,N_14321);
nor U20244 (N_20244,N_15634,N_10348);
nor U20245 (N_20245,N_14234,N_16735);
or U20246 (N_20246,N_13518,N_12643);
or U20247 (N_20247,N_14248,N_12289);
and U20248 (N_20248,N_13301,N_12263);
xor U20249 (N_20249,N_10331,N_11656);
nand U20250 (N_20250,N_13900,N_11104);
xor U20251 (N_20251,N_19793,N_15042);
and U20252 (N_20252,N_15673,N_14163);
nand U20253 (N_20253,N_19514,N_17720);
nand U20254 (N_20254,N_18756,N_19260);
nand U20255 (N_20255,N_12407,N_15697);
xnor U20256 (N_20256,N_14432,N_16125);
or U20257 (N_20257,N_17784,N_18976);
and U20258 (N_20258,N_17601,N_15835);
and U20259 (N_20259,N_19191,N_18281);
xor U20260 (N_20260,N_16298,N_18258);
xor U20261 (N_20261,N_15414,N_13163);
and U20262 (N_20262,N_10551,N_12173);
and U20263 (N_20263,N_11121,N_14591);
and U20264 (N_20264,N_18098,N_18229);
nor U20265 (N_20265,N_12981,N_16077);
nand U20266 (N_20266,N_19534,N_19088);
xor U20267 (N_20267,N_12983,N_17952);
nand U20268 (N_20268,N_15326,N_15229);
nand U20269 (N_20269,N_18315,N_19397);
and U20270 (N_20270,N_17104,N_10751);
or U20271 (N_20271,N_18805,N_19334);
or U20272 (N_20272,N_11767,N_11246);
xnor U20273 (N_20273,N_11555,N_15855);
nor U20274 (N_20274,N_14875,N_16284);
or U20275 (N_20275,N_11022,N_17990);
nand U20276 (N_20276,N_18602,N_12572);
nor U20277 (N_20277,N_15962,N_17009);
xnor U20278 (N_20278,N_14589,N_11185);
or U20279 (N_20279,N_11789,N_12574);
xnor U20280 (N_20280,N_18185,N_18493);
xnor U20281 (N_20281,N_18438,N_18922);
and U20282 (N_20282,N_15223,N_19127);
and U20283 (N_20283,N_17058,N_17231);
or U20284 (N_20284,N_11987,N_15633);
and U20285 (N_20285,N_10231,N_14547);
xnor U20286 (N_20286,N_12575,N_10546);
or U20287 (N_20287,N_18711,N_14112);
or U20288 (N_20288,N_10652,N_13252);
nand U20289 (N_20289,N_13352,N_12658);
nor U20290 (N_20290,N_10062,N_16710);
or U20291 (N_20291,N_19404,N_15961);
xor U20292 (N_20292,N_16904,N_11481);
xnor U20293 (N_20293,N_10631,N_16335);
xnor U20294 (N_20294,N_16123,N_14644);
nand U20295 (N_20295,N_11176,N_19661);
nor U20296 (N_20296,N_17705,N_14802);
and U20297 (N_20297,N_10767,N_17459);
and U20298 (N_20298,N_18089,N_17133);
and U20299 (N_20299,N_16225,N_19849);
xor U20300 (N_20300,N_14075,N_15932);
and U20301 (N_20301,N_11715,N_12727);
nand U20302 (N_20302,N_15897,N_12081);
and U20303 (N_20303,N_18169,N_13465);
nor U20304 (N_20304,N_18964,N_15213);
or U20305 (N_20305,N_10801,N_15551);
or U20306 (N_20306,N_13781,N_11215);
nand U20307 (N_20307,N_11747,N_10810);
and U20308 (N_20308,N_19044,N_17176);
xnor U20309 (N_20309,N_19612,N_14305);
or U20310 (N_20310,N_14209,N_17522);
nor U20311 (N_20311,N_14720,N_10133);
nand U20312 (N_20312,N_18702,N_14237);
xor U20313 (N_20313,N_17978,N_10393);
or U20314 (N_20314,N_12682,N_18396);
xnor U20315 (N_20315,N_15976,N_13620);
nor U20316 (N_20316,N_18589,N_16764);
xor U20317 (N_20317,N_12882,N_10643);
or U20318 (N_20318,N_15626,N_10425);
or U20319 (N_20319,N_16079,N_15829);
nand U20320 (N_20320,N_19246,N_18989);
xor U20321 (N_20321,N_10735,N_19890);
nand U20322 (N_20322,N_14734,N_10356);
nand U20323 (N_20323,N_15762,N_11175);
xnor U20324 (N_20324,N_11470,N_12428);
or U20325 (N_20325,N_10627,N_17498);
nor U20326 (N_20326,N_19736,N_12309);
and U20327 (N_20327,N_17991,N_16407);
or U20328 (N_20328,N_10846,N_17721);
or U20329 (N_20329,N_12089,N_14751);
nor U20330 (N_20330,N_16637,N_11781);
or U20331 (N_20331,N_16444,N_18861);
and U20332 (N_20332,N_12064,N_12624);
nor U20333 (N_20333,N_17036,N_11685);
or U20334 (N_20334,N_17576,N_17322);
nor U20335 (N_20335,N_12684,N_19589);
nor U20336 (N_20336,N_10772,N_14356);
and U20337 (N_20337,N_10938,N_11787);
nor U20338 (N_20338,N_16752,N_18322);
nor U20339 (N_20339,N_15875,N_15003);
xnor U20340 (N_20340,N_15654,N_10999);
nand U20341 (N_20341,N_11818,N_19350);
or U20342 (N_20342,N_16849,N_12299);
xor U20343 (N_20343,N_19598,N_18273);
nor U20344 (N_20344,N_13720,N_10806);
or U20345 (N_20345,N_16096,N_14116);
and U20346 (N_20346,N_15779,N_18330);
nand U20347 (N_20347,N_16474,N_18645);
nand U20348 (N_20348,N_19550,N_15845);
nor U20349 (N_20349,N_16778,N_12349);
nand U20350 (N_20350,N_14568,N_16222);
and U20351 (N_20351,N_19658,N_15756);
nand U20352 (N_20352,N_17103,N_19179);
and U20353 (N_20353,N_11019,N_10435);
nor U20354 (N_20354,N_19705,N_15331);
nor U20355 (N_20355,N_18028,N_13157);
nor U20356 (N_20356,N_12185,N_12065);
and U20357 (N_20357,N_11295,N_18985);
xnor U20358 (N_20358,N_10922,N_15466);
nor U20359 (N_20359,N_11896,N_11780);
or U20360 (N_20360,N_17874,N_14289);
nor U20361 (N_20361,N_13212,N_16057);
nor U20362 (N_20362,N_15416,N_10245);
xor U20363 (N_20363,N_16450,N_10178);
and U20364 (N_20364,N_10740,N_18067);
nor U20365 (N_20365,N_15713,N_10193);
xnor U20366 (N_20366,N_14859,N_14564);
nor U20367 (N_20367,N_15614,N_17570);
nand U20368 (N_20368,N_18543,N_14496);
xnor U20369 (N_20369,N_13709,N_14352);
nor U20370 (N_20370,N_15863,N_17429);
nand U20371 (N_20371,N_12294,N_12061);
nand U20372 (N_20372,N_12436,N_14865);
nand U20373 (N_20373,N_18346,N_15392);
xor U20374 (N_20374,N_14008,N_17476);
and U20375 (N_20375,N_15983,N_10439);
nand U20376 (N_20376,N_16598,N_16862);
or U20377 (N_20377,N_15737,N_16617);
nor U20378 (N_20378,N_14755,N_17357);
and U20379 (N_20379,N_16671,N_16418);
nor U20380 (N_20380,N_12559,N_14842);
and U20381 (N_20381,N_17614,N_16356);
nand U20382 (N_20382,N_17010,N_12855);
xor U20383 (N_20383,N_10893,N_14686);
nor U20384 (N_20384,N_10980,N_15373);
xor U20385 (N_20385,N_18694,N_15162);
nand U20386 (N_20386,N_15987,N_18038);
nand U20387 (N_20387,N_15903,N_11499);
nor U20388 (N_20388,N_16558,N_10912);
nor U20389 (N_20389,N_15333,N_10036);
nand U20390 (N_20390,N_14395,N_10296);
nor U20391 (N_20391,N_11509,N_13933);
nor U20392 (N_20392,N_15965,N_17443);
or U20393 (N_20393,N_12755,N_17861);
nand U20394 (N_20394,N_16609,N_17344);
and U20395 (N_20395,N_18692,N_10203);
nor U20396 (N_20396,N_10592,N_10381);
and U20397 (N_20397,N_16022,N_16882);
and U20398 (N_20398,N_19848,N_13490);
and U20399 (N_20399,N_16982,N_16135);
nand U20400 (N_20400,N_18490,N_18059);
xnor U20401 (N_20401,N_18971,N_14249);
nor U20402 (N_20402,N_18136,N_16186);
nor U20403 (N_20403,N_16785,N_10209);
or U20404 (N_20404,N_10268,N_17597);
xnor U20405 (N_20405,N_17667,N_12320);
or U20406 (N_20406,N_15978,N_18567);
nand U20407 (N_20407,N_15474,N_10649);
and U20408 (N_20408,N_16394,N_12054);
and U20409 (N_20409,N_17624,N_12694);
xor U20410 (N_20410,N_10037,N_15047);
or U20411 (N_20411,N_16641,N_13656);
xnor U20412 (N_20412,N_19629,N_11657);
nor U20413 (N_20413,N_14145,N_16314);
nor U20414 (N_20414,N_12218,N_15209);
xnor U20415 (N_20415,N_12612,N_11068);
and U20416 (N_20416,N_13387,N_10694);
nor U20417 (N_20417,N_15645,N_17316);
nand U20418 (N_20418,N_13818,N_19532);
nand U20419 (N_20419,N_15872,N_11299);
or U20420 (N_20420,N_15178,N_16830);
nand U20421 (N_20421,N_10901,N_10447);
nor U20422 (N_20422,N_10001,N_19796);
nand U20423 (N_20423,N_13881,N_17144);
or U20424 (N_20424,N_17514,N_10147);
or U20425 (N_20425,N_18109,N_17175);
nand U20426 (N_20426,N_14083,N_16566);
xnor U20427 (N_20427,N_11480,N_17972);
and U20428 (N_20428,N_18364,N_12757);
or U20429 (N_20429,N_17200,N_10717);
nand U20430 (N_20430,N_11447,N_11148);
or U20431 (N_20431,N_12820,N_15269);
nand U20432 (N_20432,N_12239,N_13122);
xnor U20433 (N_20433,N_16244,N_10781);
or U20434 (N_20434,N_12674,N_19389);
xnor U20435 (N_20435,N_15594,N_10330);
xor U20436 (N_20436,N_17731,N_18446);
xor U20437 (N_20437,N_17318,N_17219);
xor U20438 (N_20438,N_14223,N_15530);
nand U20439 (N_20439,N_18728,N_14299);
xnor U20440 (N_20440,N_14135,N_16951);
nand U20441 (N_20441,N_13898,N_19040);
nor U20442 (N_20442,N_15421,N_14201);
and U20443 (N_20443,N_19906,N_12911);
nand U20444 (N_20444,N_11160,N_12745);
or U20445 (N_20445,N_16323,N_12274);
xnor U20446 (N_20446,N_10206,N_18994);
and U20447 (N_20447,N_19503,N_11126);
xor U20448 (N_20448,N_11039,N_12395);
and U20449 (N_20449,N_17793,N_11674);
xor U20450 (N_20450,N_11038,N_19136);
nor U20451 (N_20451,N_19193,N_14677);
or U20452 (N_20452,N_11187,N_12376);
and U20453 (N_20453,N_17894,N_16941);
nor U20454 (N_20454,N_12148,N_19407);
xnor U20455 (N_20455,N_19676,N_14424);
xnor U20456 (N_20456,N_15819,N_10841);
nor U20457 (N_20457,N_13703,N_10171);
or U20458 (N_20458,N_18673,N_19632);
and U20459 (N_20459,N_17330,N_18367);
and U20460 (N_20460,N_14888,N_16581);
xnor U20461 (N_20461,N_14073,N_19059);
xor U20462 (N_20462,N_13661,N_12984);
nand U20463 (N_20463,N_14619,N_17212);
and U20464 (N_20464,N_10629,N_18622);
xnor U20465 (N_20465,N_14681,N_10967);
and U20466 (N_20466,N_18495,N_12493);
nand U20467 (N_20467,N_16618,N_11232);
and U20468 (N_20468,N_10863,N_12530);
and U20469 (N_20469,N_15177,N_18196);
nand U20470 (N_20470,N_10883,N_17506);
nor U20471 (N_20471,N_12929,N_17655);
nor U20472 (N_20472,N_19968,N_11244);
and U20473 (N_20473,N_12402,N_13928);
nand U20474 (N_20474,N_16203,N_18342);
nand U20475 (N_20475,N_14336,N_14313);
and U20476 (N_20476,N_15815,N_19741);
xnor U20477 (N_20477,N_13341,N_13308);
xnor U20478 (N_20478,N_13189,N_12866);
nor U20479 (N_20479,N_12004,N_15194);
nor U20480 (N_20480,N_18083,N_18938);
or U20481 (N_20481,N_17153,N_10664);
nand U20482 (N_20482,N_17918,N_11615);
and U20483 (N_20483,N_16115,N_19749);
and U20484 (N_20484,N_12827,N_12388);
nor U20485 (N_20485,N_10379,N_18426);
or U20486 (N_20486,N_19709,N_14373);
and U20487 (N_20487,N_19596,N_17622);
and U20488 (N_20488,N_15461,N_12026);
nor U20489 (N_20489,N_10928,N_11449);
nor U20490 (N_20490,N_17710,N_15934);
nor U20491 (N_20491,N_19601,N_15007);
or U20492 (N_20492,N_16279,N_18483);
and U20493 (N_20493,N_19048,N_13923);
xnor U20494 (N_20494,N_18592,N_16595);
nand U20495 (N_20495,N_15351,N_10179);
and U20496 (N_20496,N_17867,N_14680);
nor U20497 (N_20497,N_13521,N_11356);
nand U20498 (N_20498,N_11297,N_11737);
xnor U20499 (N_20499,N_10314,N_14097);
nand U20500 (N_20500,N_14296,N_18338);
or U20501 (N_20501,N_12828,N_16255);
nor U20502 (N_20502,N_19394,N_18251);
nor U20503 (N_20503,N_16091,N_13517);
xor U20504 (N_20504,N_16413,N_16898);
and U20505 (N_20505,N_15743,N_12251);
nand U20506 (N_20506,N_14220,N_18724);
xnor U20507 (N_20507,N_13981,N_12397);
xor U20508 (N_20508,N_12750,N_11428);
nor U20509 (N_20509,N_14572,N_11385);
and U20510 (N_20510,N_15843,N_17294);
or U20511 (N_20511,N_12554,N_12103);
or U20512 (N_20512,N_11935,N_16087);
or U20513 (N_20513,N_12130,N_15118);
or U20514 (N_20514,N_12151,N_12224);
xnor U20515 (N_20515,N_16152,N_15639);
nand U20516 (N_20516,N_19939,N_12193);
nor U20517 (N_20517,N_18324,N_17892);
and U20518 (N_20518,N_16149,N_17210);
nand U20519 (N_20519,N_14955,N_18731);
xnor U20520 (N_20520,N_12000,N_19945);
nor U20521 (N_20521,N_13634,N_19308);
or U20522 (N_20522,N_13929,N_16932);
or U20523 (N_20523,N_19546,N_12112);
xor U20524 (N_20524,N_13116,N_10430);
nor U20525 (N_20525,N_19058,N_16012);
and U20526 (N_20526,N_12653,N_17260);
nor U20527 (N_20527,N_15110,N_19816);
nand U20528 (N_20528,N_14122,N_10466);
xor U20529 (N_20529,N_16775,N_16606);
nand U20530 (N_20530,N_10586,N_11003);
nand U20531 (N_20531,N_17343,N_18799);
and U20532 (N_20532,N_12262,N_11386);
and U20533 (N_20533,N_14425,N_18184);
nand U20534 (N_20534,N_11464,N_10997);
nor U20535 (N_20535,N_15475,N_12834);
nand U20536 (N_20536,N_16332,N_16143);
nor U20537 (N_20537,N_17881,N_12057);
nor U20538 (N_20538,N_17093,N_11168);
and U20539 (N_20539,N_19772,N_12074);
nand U20540 (N_20540,N_14561,N_16183);
nand U20541 (N_20541,N_14966,N_12998);
nand U20542 (N_20542,N_12095,N_16685);
and U20543 (N_20543,N_19805,N_14592);
xnor U20544 (N_20544,N_11240,N_14011);
or U20545 (N_20545,N_19937,N_16583);
xor U20546 (N_20546,N_15400,N_10160);
and U20547 (N_20547,N_10575,N_11219);
xnor U20548 (N_20548,N_11421,N_14387);
or U20549 (N_20549,N_12347,N_14906);
or U20550 (N_20550,N_18800,N_15085);
xor U20551 (N_20551,N_19670,N_13680);
nand U20552 (N_20552,N_10739,N_19496);
nor U20553 (N_20553,N_18593,N_17251);
nor U20554 (N_20554,N_16569,N_15950);
nor U20555 (N_20555,N_19821,N_12494);
or U20556 (N_20556,N_16766,N_16501);
or U20557 (N_20557,N_13145,N_18707);
or U20558 (N_20558,N_17977,N_13511);
and U20559 (N_20559,N_19151,N_17897);
nor U20560 (N_20560,N_18889,N_15928);
xnor U20561 (N_20561,N_10747,N_15267);
nor U20562 (N_20562,N_16758,N_18647);
xnor U20563 (N_20563,N_15741,N_11081);
xor U20564 (N_20564,N_16765,N_19677);
nor U20565 (N_20565,N_12547,N_10744);
nor U20566 (N_20566,N_17862,N_11601);
nor U20567 (N_20567,N_18039,N_15899);
nand U20568 (N_20568,N_15303,N_13524);
nand U20569 (N_20569,N_15144,N_15497);
and U20570 (N_20570,N_11082,N_10342);
or U20571 (N_20571,N_11025,N_16719);
nor U20572 (N_20572,N_10805,N_16597);
xor U20573 (N_20573,N_16272,N_18508);
nor U20574 (N_20574,N_12925,N_14062);
nand U20575 (N_20575,N_14890,N_17470);
nor U20576 (N_20576,N_16792,N_19423);
or U20577 (N_20577,N_16108,N_14153);
nor U20578 (N_20578,N_14362,N_12909);
and U20579 (N_20579,N_17621,N_18168);
and U20580 (N_20580,N_12831,N_16487);
or U20581 (N_20581,N_13951,N_12738);
or U20582 (N_20582,N_11642,N_13632);
or U20583 (N_20583,N_18682,N_14247);
nand U20584 (N_20584,N_11745,N_15629);
or U20585 (N_20585,N_16967,N_14303);
or U20586 (N_20586,N_17491,N_15625);
xor U20587 (N_20587,N_10180,N_13367);
or U20588 (N_20588,N_18590,N_10039);
nor U20589 (N_20589,N_11726,N_13420);
nor U20590 (N_20590,N_13069,N_17303);
or U20591 (N_20591,N_17589,N_10655);
xnor U20592 (N_20592,N_15494,N_15853);
or U20593 (N_20593,N_13595,N_17477);
nand U20594 (N_20594,N_13962,N_14758);
nand U20595 (N_20595,N_18770,N_19330);
nor U20596 (N_20596,N_11399,N_15710);
or U20597 (N_20597,N_13489,N_14052);
nand U20598 (N_20598,N_10251,N_13401);
and U20599 (N_20599,N_11799,N_11525);
or U20600 (N_20600,N_10734,N_19948);
or U20601 (N_20601,N_15190,N_15814);
xnor U20602 (N_20602,N_13944,N_10597);
or U20603 (N_20603,N_18851,N_16481);
or U20604 (N_20604,N_11328,N_16621);
or U20605 (N_20605,N_15681,N_14825);
xnor U20606 (N_20606,N_17348,N_10613);
or U20607 (N_20607,N_16027,N_19449);
and U20608 (N_20608,N_12838,N_18591);
nand U20609 (N_20609,N_11628,N_13123);
or U20610 (N_20610,N_13034,N_10365);
nor U20611 (N_20611,N_17163,N_11558);
nor U20612 (N_20612,N_12486,N_17062);
or U20613 (N_20613,N_12538,N_17707);
or U20614 (N_20614,N_14244,N_11174);
nor U20615 (N_20615,N_19157,N_19686);
nor U20616 (N_20616,N_15054,N_13846);
nor U20617 (N_20617,N_16527,N_13016);
and U20618 (N_20618,N_17868,N_10405);
or U20619 (N_20619,N_17927,N_10132);
and U20620 (N_20620,N_16600,N_11051);
nor U20621 (N_20621,N_15149,N_17762);
nor U20622 (N_20622,N_14857,N_11992);
nor U20623 (N_20623,N_19909,N_10509);
and U20624 (N_20624,N_15080,N_17717);
xor U20625 (N_20625,N_19663,N_17818);
nor U20626 (N_20626,N_17078,N_14149);
xnor U20627 (N_20627,N_11692,N_17304);
or U20628 (N_20628,N_16426,N_12829);
or U20629 (N_20629,N_11610,N_16497);
xnor U20630 (N_20630,N_17254,N_14723);
xnor U20631 (N_20631,N_17538,N_15259);
nand U20632 (N_20632,N_16525,N_15258);
or U20633 (N_20633,N_16389,N_14793);
nor U20634 (N_20634,N_18598,N_19771);
nand U20635 (N_20635,N_11439,N_14064);
and U20636 (N_20636,N_11218,N_11588);
nand U20637 (N_20637,N_15501,N_10831);
and U20638 (N_20638,N_19235,N_12629);
nor U20639 (N_20639,N_10471,N_16592);
or U20640 (N_20640,N_17807,N_19288);
or U20641 (N_20641,N_16408,N_11589);
nor U20642 (N_20642,N_13645,N_12967);
or U20643 (N_20643,N_12029,N_14101);
xor U20644 (N_20644,N_13501,N_15328);
xor U20645 (N_20645,N_11096,N_12551);
xnor U20646 (N_20646,N_14506,N_11868);
and U20647 (N_20647,N_10043,N_10319);
nor U20648 (N_20648,N_16002,N_12021);
xor U20649 (N_20649,N_13491,N_16280);
and U20650 (N_20650,N_17194,N_10720);
nand U20651 (N_20651,N_10851,N_18408);
xnor U20652 (N_20652,N_14961,N_13682);
xor U20653 (N_20653,N_13966,N_12328);
and U20654 (N_20654,N_10107,N_17391);
nor U20655 (N_20655,N_17196,N_18706);
nor U20656 (N_20656,N_19017,N_13267);
or U20657 (N_20657,N_16295,N_19299);
xor U20658 (N_20658,N_12235,N_16173);
and U20659 (N_20659,N_11330,N_14167);
and U20660 (N_20660,N_15453,N_14529);
and U20661 (N_20661,N_15995,N_14784);
nor U20662 (N_20662,N_18340,N_19255);
or U20663 (N_20663,N_16021,N_18286);
and U20664 (N_20664,N_15982,N_14202);
nand U20665 (N_20665,N_14491,N_17384);
nand U20666 (N_20666,N_11487,N_17063);
or U20667 (N_20667,N_14158,N_18449);
or U20668 (N_20668,N_15717,N_14417);
and U20669 (N_20669,N_12963,N_10540);
or U20670 (N_20670,N_19994,N_18934);
or U20671 (N_20671,N_10164,N_11748);
nand U20672 (N_20672,N_11713,N_17708);
or U20673 (N_20673,N_13655,N_14633);
nand U20674 (N_20674,N_12673,N_10714);
nand U20675 (N_20675,N_14544,N_19004);
or U20676 (N_20676,N_11977,N_11543);
or U20677 (N_20677,N_19436,N_16154);
and U20678 (N_20678,N_19064,N_17528);
or U20679 (N_20679,N_11652,N_10269);
nand U20680 (N_20680,N_12584,N_15547);
xnor U20681 (N_20681,N_13411,N_13685);
xnor U20682 (N_20682,N_10394,N_15198);
or U20683 (N_20683,N_15044,N_15428);
and U20684 (N_20684,N_10557,N_16924);
and U20685 (N_20685,N_17172,N_13778);
or U20686 (N_20686,N_10814,N_13207);
nand U20687 (N_20687,N_19630,N_10977);
nand U20688 (N_20688,N_11793,N_15705);
and U20689 (N_20689,N_11413,N_14667);
and U20690 (N_20690,N_13438,N_14962);
xnor U20691 (N_20691,N_15698,N_11529);
and U20692 (N_20692,N_10085,N_17342);
nand U20693 (N_20693,N_18132,N_13979);
and U20694 (N_20694,N_16936,N_16103);
nor U20695 (N_20695,N_18000,N_15791);
nand U20696 (N_20696,N_11740,N_16340);
xor U20697 (N_20697,N_15310,N_11261);
xor U20698 (N_20698,N_16116,N_19042);
nor U20699 (N_20699,N_11978,N_16992);
nor U20700 (N_20700,N_10759,N_14698);
and U20701 (N_20701,N_11946,N_10384);
or U20702 (N_20702,N_13310,N_11928);
nand U20703 (N_20703,N_11202,N_13533);
and U20704 (N_20704,N_19333,N_13125);
nand U20705 (N_20705,N_14990,N_13183);
nor U20706 (N_20706,N_12443,N_16915);
xor U20707 (N_20707,N_10421,N_13075);
and U20708 (N_20708,N_16552,N_15955);
nor U20709 (N_20709,N_12610,N_18411);
nor U20710 (N_20710,N_17431,N_15381);
or U20711 (N_20711,N_19452,N_19902);
or U20712 (N_20712,N_19859,N_14047);
and U20713 (N_20713,N_10571,N_14783);
xnor U20714 (N_20714,N_18270,N_18125);
xnor U20715 (N_20715,N_10873,N_12604);
nand U20716 (N_20716,N_19412,N_17148);
or U20717 (N_20717,N_16304,N_14662);
or U20718 (N_20718,N_11775,N_18049);
xor U20719 (N_20719,N_18845,N_12042);
nand U20720 (N_20720,N_16827,N_18401);
or U20721 (N_20721,N_19899,N_15132);
nand U20722 (N_20722,N_16756,N_17249);
nor U20723 (N_20723,N_11960,N_13152);
or U20724 (N_20724,N_13061,N_18335);
nand U20725 (N_20725,N_10402,N_19922);
nor U20726 (N_20726,N_14294,N_10483);
nand U20727 (N_20727,N_16494,N_15215);
nor U20728 (N_20728,N_18837,N_11965);
nor U20729 (N_20729,N_12955,N_14527);
nand U20730 (N_20730,N_10146,N_17402);
or U20731 (N_20731,N_17625,N_13874);
xnor U20732 (N_20732,N_14484,N_12508);
xnor U20733 (N_20733,N_14504,N_15033);
nor U20734 (N_20734,N_18667,N_11779);
nand U20735 (N_20735,N_11212,N_19030);
xnor U20736 (N_20736,N_11842,N_11432);
xnor U20737 (N_20737,N_16506,N_13108);
nand U20738 (N_20738,N_19227,N_12177);
or U20739 (N_20739,N_14398,N_10899);
or U20740 (N_20740,N_10576,N_15929);
and U20741 (N_20741,N_16895,N_13637);
or U20742 (N_20742,N_17527,N_17517);
xor U20743 (N_20743,N_12852,N_14597);
nand U20744 (N_20744,N_12296,N_13078);
nor U20745 (N_20745,N_12312,N_18506);
xnor U20746 (N_20746,N_16770,N_12522);
nand U20747 (N_20747,N_10670,N_17672);
and U20748 (N_20748,N_17670,N_10207);
xor U20749 (N_20749,N_12722,N_10960);
nand U20750 (N_20750,N_18571,N_12055);
nand U20751 (N_20751,N_16182,N_13935);
nand U20752 (N_20752,N_12539,N_12085);
nand U20753 (N_20753,N_13346,N_14797);
nor U20754 (N_20754,N_18094,N_10828);
and U20755 (N_20755,N_14605,N_15553);
or U20756 (N_20756,N_13383,N_15752);
nand U20757 (N_20757,N_12622,N_17554);
xnor U20758 (N_20758,N_11521,N_13049);
nor U20759 (N_20759,N_15541,N_15582);
nor U20760 (N_20760,N_11491,N_10682);
nor U20761 (N_20761,N_16276,N_10804);
and U20762 (N_20762,N_10005,N_12119);
nand U20763 (N_20763,N_14070,N_19499);
and U20764 (N_20764,N_16940,N_13953);
nor U20765 (N_20765,N_17209,N_14268);
nor U20766 (N_20766,N_19358,N_15831);
or U20767 (N_20767,N_11238,N_15611);
nor U20768 (N_20768,N_12445,N_13246);
and U20769 (N_20769,N_17647,N_14671);
nor U20770 (N_20770,N_17992,N_13096);
nor U20771 (N_20771,N_15376,N_19956);
xnor U20772 (N_20772,N_19435,N_18675);
nand U20773 (N_20773,N_16242,N_11352);
xor U20774 (N_20774,N_12009,N_10741);
nor U20775 (N_20775,N_11819,N_10876);
or U20776 (N_20776,N_13262,N_12115);
nor U20777 (N_20777,N_16465,N_17412);
or U20778 (N_20778,N_14517,N_15173);
or U20779 (N_20779,N_11204,N_15669);
and U20780 (N_20780,N_13686,N_14656);
xor U20781 (N_20781,N_14975,N_10208);
nor U20782 (N_20782,N_18943,N_18939);
nand U20783 (N_20783,N_16336,N_15802);
nor U20784 (N_20784,N_17087,N_13920);
xor U20785 (N_20785,N_17626,N_19520);
nor U20786 (N_20786,N_18422,N_19486);
xnor U20787 (N_20787,N_10263,N_12346);
or U20788 (N_20788,N_13699,N_10007);
or U20789 (N_20789,N_17676,N_18562);
xnor U20790 (N_20790,N_19882,N_15898);
or U20791 (N_20791,N_11359,N_19118);
nor U20792 (N_20792,N_13322,N_12783);
nand U20793 (N_20793,N_19699,N_17099);
and U20794 (N_20794,N_13814,N_12351);
or U20795 (N_20795,N_12979,N_15514);
nand U20796 (N_20796,N_10006,N_16639);
or U20797 (N_20797,N_12069,N_18084);
or U20798 (N_20798,N_10825,N_16275);
nand U20799 (N_20799,N_14456,N_12649);
nand U20800 (N_20800,N_14594,N_17789);
xor U20801 (N_20801,N_17530,N_11976);
nand U20802 (N_20802,N_18032,N_14679);
nand U20803 (N_20803,N_11472,N_16682);
nor U20804 (N_20804,N_15318,N_15518);
nand U20805 (N_20805,N_10083,N_16004);
or U20806 (N_20806,N_11560,N_13730);
xor U20807 (N_20807,N_15967,N_18473);
nand U20808 (N_20808,N_17277,N_18664);
nor U20809 (N_20809,N_17376,N_15840);
or U20810 (N_20810,N_16791,N_19730);
and U20811 (N_20811,N_14182,N_17962);
nand U20812 (N_20812,N_11134,N_12666);
and U20813 (N_20813,N_19344,N_18478);
and U20814 (N_20814,N_18226,N_14007);
nor U20815 (N_20815,N_10515,N_16975);
xor U20816 (N_20816,N_19056,N_15963);
or U20817 (N_20817,N_17809,N_10661);
nor U20818 (N_20818,N_10895,N_17461);
xnor U20819 (N_20819,N_11966,N_17686);
and U20820 (N_20820,N_10463,N_14359);
or U20821 (N_20821,N_11600,N_17296);
nand U20822 (N_20822,N_12187,N_12485);
nor U20823 (N_20823,N_15394,N_18224);
xnor U20824 (N_20824,N_10187,N_16708);
nor U20825 (N_20825,N_18470,N_16257);
nor U20826 (N_20826,N_14844,N_15472);
xnor U20827 (N_20827,N_12626,N_10301);
nand U20828 (N_20828,N_11846,N_13044);
and U20829 (N_20829,N_11285,N_15602);
xnor U20830 (N_20830,N_12217,N_15343);
or U20831 (N_20831,N_11375,N_11647);
and U20832 (N_20832,N_19029,N_11343);
xnor U20833 (N_20833,N_11037,N_10293);
nand U20834 (N_20834,N_15391,N_10041);
xnor U20835 (N_20835,N_11095,N_19967);
nor U20836 (N_20836,N_16662,N_14087);
or U20837 (N_20837,N_14391,N_15164);
or U20838 (N_20838,N_18659,N_10989);
xor U20839 (N_20839,N_10236,N_17805);
xor U20840 (N_20840,N_15866,N_14060);
nor U20841 (N_20841,N_11043,N_18467);
or U20842 (N_20842,N_18898,N_18961);
xor U20843 (N_20843,N_17291,N_12389);
or U20844 (N_20844,N_18677,N_12420);
or U20845 (N_20845,N_19014,N_12355);
xnor U20846 (N_20846,N_12150,N_19631);
xor U20847 (N_20847,N_17692,N_15906);
nand U20848 (N_20848,N_19332,N_13359);
nand U20849 (N_20849,N_14869,N_16857);
or U20850 (N_20850,N_10272,N_14498);
nor U20851 (N_20851,N_12710,N_12114);
nand U20852 (N_20852,N_19976,N_13976);
nor U20853 (N_20853,N_11041,N_15218);
and U20854 (N_20854,N_12654,N_19329);
or U20855 (N_20855,N_13297,N_14815);
xor U20856 (N_20856,N_12378,N_12008);
nand U20857 (N_20857,N_14206,N_15911);
nand U20858 (N_20858,N_19605,N_16210);
nand U20859 (N_20859,N_12797,N_13537);
nand U20860 (N_20860,N_17645,N_11365);
and U20861 (N_20861,N_12451,N_11455);
nor U20862 (N_20862,N_15957,N_16828);
nor U20863 (N_20863,N_15850,N_14982);
nand U20864 (N_20864,N_14200,N_14041);
xnor U20865 (N_20865,N_12363,N_16721);
or U20866 (N_20866,N_11776,N_17206);
nand U20867 (N_20867,N_14852,N_19669);
nand U20868 (N_20868,N_19754,N_12491);
xnor U20869 (N_20869,N_12790,N_18496);
nand U20870 (N_20870,N_11911,N_17363);
nor U20871 (N_20871,N_15732,N_13447);
and U20872 (N_20872,N_14304,N_15325);
xor U20873 (N_20873,N_15116,N_11479);
or U20874 (N_20874,N_11731,N_14753);
or U20875 (N_20875,N_12950,N_16966);
and U20876 (N_20876,N_17736,N_12327);
and U20877 (N_20877,N_14757,N_13345);
nor U20878 (N_20878,N_18430,N_13195);
or U20879 (N_20879,N_12916,N_10410);
or U20880 (N_20880,N_14050,N_16996);
nand U20881 (N_20881,N_11433,N_14994);
xnor U20882 (N_20882,N_16024,N_18235);
xnor U20883 (N_20883,N_10247,N_12280);
or U20884 (N_20884,N_11042,N_16409);
or U20885 (N_20885,N_10662,N_17882);
and U20886 (N_20886,N_13870,N_15871);
and U20887 (N_20887,N_14718,N_11149);
and U20888 (N_20888,N_16724,N_17761);
or U20889 (N_20889,N_14549,N_11638);
nand U20890 (N_20890,N_10639,N_12997);
xnor U20891 (N_20891,N_14831,N_14026);
xor U20892 (N_20892,N_17804,N_18045);
nand U20893 (N_20893,N_15288,N_17113);
nor U20894 (N_20894,N_11231,N_10757);
nand U20895 (N_20895,N_13967,N_19742);
and U20896 (N_20896,N_11339,N_13640);
and U20897 (N_20897,N_18868,N_11704);
nor U20898 (N_20898,N_16833,N_19024);
or U20899 (N_20899,N_11242,N_18951);
xor U20900 (N_20900,N_15603,N_17253);
and U20901 (N_20901,N_16207,N_13292);
and U20902 (N_20902,N_18537,N_11484);
nand U20903 (N_20903,N_13687,N_13666);
nand U20904 (N_20904,N_11832,N_17080);
nand U20905 (N_20905,N_18842,N_15450);
and U20906 (N_20906,N_17135,N_11933);
xnor U20907 (N_20907,N_19497,N_16739);
or U20908 (N_20908,N_18691,N_17558);
or U20909 (N_20909,N_15056,N_14845);
nand U20910 (N_20910,N_18252,N_10881);
nor U20911 (N_20911,N_15516,N_12252);
nand U20912 (N_20912,N_12659,N_15297);
or U20913 (N_20913,N_15051,N_14861);
nand U20914 (N_20914,N_13866,N_14281);
and U20915 (N_20915,N_17411,N_12913);
nand U20916 (N_20916,N_13319,N_17239);
or U20917 (N_20917,N_12985,N_19477);
and U20918 (N_20918,N_14143,N_15445);
xnor U20919 (N_20919,N_11329,N_15330);
nor U20920 (N_20920,N_16893,N_14388);
and U20921 (N_20921,N_10538,N_12045);
nand U20922 (N_20922,N_10403,N_10622);
nand U20923 (N_20923,N_10167,N_18509);
nor U20924 (N_20924,N_19174,N_15768);
and U20925 (N_20925,N_15508,N_17899);
or U20926 (N_20926,N_19878,N_16737);
xor U20927 (N_20927,N_17505,N_10138);
xor U20928 (N_20928,N_18900,N_13974);
xor U20929 (N_20929,N_11936,N_15748);
nor U20930 (N_20930,N_16176,N_12298);
nand U20931 (N_20931,N_16524,N_18310);
or U20932 (N_20932,N_10176,N_18780);
or U20933 (N_20933,N_12429,N_15250);
and U20934 (N_20934,N_13616,N_13707);
and U20935 (N_20935,N_19357,N_11828);
nor U20936 (N_20936,N_18581,N_12070);
and U20937 (N_20937,N_17600,N_11566);
nor U20938 (N_20938,N_16044,N_11054);
or U20939 (N_20939,N_15812,N_13233);
nand U20940 (N_20940,N_14493,N_10172);
nor U20941 (N_20941,N_16232,N_10963);
xnor U20942 (N_20942,N_15236,N_16555);
nor U20943 (N_20943,N_19450,N_17315);
or U20944 (N_20944,N_17002,N_15058);
nand U20945 (N_20945,N_19525,N_17856);
xnor U20946 (N_20946,N_10605,N_10444);
nor U20947 (N_20947,N_12145,N_11319);
or U20948 (N_20948,N_17379,N_18081);
nand U20949 (N_20949,N_16029,N_19495);
and U20950 (N_20950,N_14374,N_15595);
and U20951 (N_20951,N_15809,N_18709);
nand U20952 (N_20952,N_14924,N_12590);
nand U20953 (N_20953,N_18167,N_18982);
or U20954 (N_20954,N_12865,N_15703);
xor U20955 (N_20955,N_10516,N_15309);
nor U20956 (N_20956,N_15837,N_19891);
nor U20957 (N_20957,N_16949,N_11836);
or U20958 (N_20958,N_17136,N_15749);
nand U20959 (N_20959,N_15423,N_17186);
and U20960 (N_20960,N_15766,N_10267);
and U20961 (N_20961,N_13745,N_10973);
nor U20962 (N_20962,N_16899,N_17529);
nand U20963 (N_20963,N_18720,N_14381);
nand U20964 (N_20964,N_17526,N_10303);
xnor U20965 (N_20965,N_13064,N_13914);
nand U20966 (N_20966,N_14684,N_17953);
and U20967 (N_20967,N_18227,N_17387);
nand U20968 (N_20968,N_11855,N_17613);
nand U20969 (N_20969,N_17042,N_19777);
and U20970 (N_20970,N_14548,N_11577);
and U20971 (N_20971,N_18714,N_16005);
nand U20972 (N_20972,N_15935,N_15000);
nor U20973 (N_20973,N_13568,N_15066);
nand U20974 (N_20974,N_10165,N_17378);
nor U20975 (N_20975,N_11435,N_13429);
and U20976 (N_20976,N_17267,N_13667);
nor U20977 (N_20977,N_13132,N_17236);
nand U20978 (N_20978,N_11862,N_16615);
and U20979 (N_20979,N_12679,N_13120);
nor U20980 (N_20980,N_12930,N_11290);
nand U20981 (N_20981,N_12075,N_14492);
or U20982 (N_20982,N_15457,N_17340);
xnor U20983 (N_20983,N_13623,N_18320);
and U20984 (N_20984,N_15656,N_13610);
and U20985 (N_20985,N_15129,N_17130);
nor U20986 (N_20986,N_15998,N_15396);
xnor U20987 (N_20987,N_13845,N_17436);
xnor U20988 (N_20988,N_18044,N_15010);
and U20989 (N_20989,N_17832,N_15185);
and U20990 (N_20990,N_12316,N_12875);
xor U20991 (N_20991,N_17795,N_12284);
and U20992 (N_20992,N_16083,N_18755);
nor U20993 (N_20993,N_19374,N_15512);
nor U20994 (N_20994,N_14279,N_11872);
nand U20995 (N_20995,N_18923,N_12350);
nand U20996 (N_20996,N_19961,N_17581);
nor U20997 (N_20997,N_10283,N_15112);
nand U20998 (N_20998,N_17730,N_10550);
nor U20999 (N_20999,N_13790,N_14147);
or U21000 (N_21000,N_17437,N_11722);
nand U21001 (N_21001,N_12072,N_12214);
xor U21002 (N_21002,N_10572,N_12333);
nand U21003 (N_21003,N_15050,N_13579);
nor U21004 (N_21004,N_13110,N_16391);
nand U21005 (N_21005,N_17758,N_19636);
nor U21006 (N_21006,N_16654,N_16665);
and U21007 (N_21007,N_17725,N_19498);
xnor U21008 (N_21008,N_10491,N_16825);
xor U21009 (N_21009,N_15870,N_10511);
nand U21010 (N_21010,N_16628,N_13062);
nor U21011 (N_21011,N_17863,N_11696);
or U21012 (N_21012,N_15447,N_18279);
or U21013 (N_21013,N_16159,N_18246);
nand U21014 (N_21014,N_18753,N_14649);
nand U21015 (N_21015,N_18915,N_10632);
and U21016 (N_21016,N_15926,N_10505);
nor U21017 (N_21017,N_15610,N_10530);
and U21018 (N_21018,N_10958,N_18103);
or U21019 (N_21019,N_13476,N_18474);
and U21020 (N_21020,N_12524,N_19181);
nand U21021 (N_21021,N_16344,N_10227);
xnor U21022 (N_21022,N_15613,N_18771);
or U21023 (N_21023,N_17232,N_11281);
and U21024 (N_21024,N_19206,N_10679);
or U21025 (N_21025,N_15268,N_11571);
nand U21026 (N_21026,N_16428,N_17418);
xor U21027 (N_21027,N_16805,N_16977);
or U21028 (N_21028,N_10442,N_18066);
nor U21029 (N_21029,N_15909,N_14838);
nor U21030 (N_21030,N_18940,N_10411);
or U21031 (N_21031,N_14874,N_11016);
nor U21032 (N_21032,N_16142,N_19916);
nand U21033 (N_21033,N_11467,N_13362);
xnor U21034 (N_21034,N_18337,N_19843);
and U21035 (N_21035,N_17445,N_12359);
nor U21036 (N_21036,N_13014,N_14377);
nand U21037 (N_21037,N_17540,N_19883);
and U21038 (N_21038,N_12168,N_16368);
and U21039 (N_21039,N_13960,N_11222);
xor U21040 (N_21040,N_17541,N_18482);
or U21041 (N_21041,N_12969,N_11897);
nand U21042 (N_21042,N_13251,N_16788);
nand U21043 (N_21043,N_11031,N_13316);
or U21044 (N_21044,N_10821,N_17924);
nand U21045 (N_21045,N_12140,N_13879);
and U21046 (N_21046,N_16462,N_15278);
or U21047 (N_21047,N_15757,N_18942);
nand U21048 (N_21048,N_17574,N_18856);
nor U21049 (N_21049,N_18577,N_17796);
nand U21050 (N_21050,N_19242,N_13187);
and U21051 (N_21051,N_15244,N_17299);
nor U21052 (N_21052,N_11221,N_16360);
and U21053 (N_21053,N_15842,N_10281);
nor U21054 (N_21054,N_11079,N_14277);
or U21055 (N_21055,N_19521,N_14159);
and U21056 (N_21056,N_12012,N_18993);
nand U21057 (N_21057,N_15940,N_12887);
nor U21058 (N_21058,N_18674,N_12340);
and U21059 (N_21059,N_18410,N_19478);
xnor U21060 (N_21060,N_12589,N_18646);
nand U21061 (N_21061,N_16157,N_11434);
xnor U21062 (N_21062,N_16696,N_18833);
nor U21063 (N_21063,N_13100,N_19083);
and U21064 (N_21064,N_19566,N_14461);
or U21065 (N_21065,N_17542,N_11311);
xor U21066 (N_21066,N_11888,N_11677);
nand U21067 (N_21067,N_17713,N_19564);
and U21068 (N_21068,N_10990,N_14366);
xnor U21069 (N_21069,N_17259,N_19770);
or U21070 (N_21070,N_11165,N_18250);
xnor U21071 (N_21071,N_15720,N_14726);
nand U21072 (N_21072,N_16260,N_16769);
nor U21073 (N_21073,N_11419,N_12446);
xnor U21074 (N_21074,N_14601,N_14164);
or U21075 (N_21075,N_15021,N_15985);
nand U21076 (N_21076,N_14430,N_18126);
nand U21077 (N_21077,N_11135,N_12146);
or U21078 (N_21078,N_12357,N_11336);
xnor U21079 (N_21079,N_16216,N_13021);
or U21080 (N_21080,N_17488,N_12697);
and U21081 (N_21081,N_14467,N_10725);
nor U21082 (N_21082,N_19679,N_17326);
or U21083 (N_21083,N_18249,N_15289);
or U21084 (N_21084,N_10397,N_13643);
nor U21085 (N_21085,N_13444,N_13130);
and U21086 (N_21086,N_19960,N_19163);
or U21087 (N_21087,N_10478,N_19026);
and U21088 (N_21088,N_12161,N_19177);
and U21089 (N_21089,N_18757,N_18925);
nand U21090 (N_21090,N_14385,N_10197);
nand U21091 (N_21091,N_17012,N_16098);
and U21092 (N_21092,N_12326,N_16947);
and U21093 (N_21093,N_15801,N_10304);
and U21094 (N_21094,N_15111,N_16601);
nor U21095 (N_21095,N_18090,N_13277);
nor U21096 (N_21096,N_13097,N_11598);
and U21097 (N_21097,N_13621,N_12212);
nor U21098 (N_21098,N_14873,N_19376);
xor U21099 (N_21099,N_13550,N_13751);
and U21100 (N_21100,N_19619,N_18123);
nand U21101 (N_21101,N_10035,N_13495);
nor U21102 (N_21102,N_18888,N_15075);
nor U21103 (N_21103,N_14160,N_17280);
or U21104 (N_21104,N_14552,N_11369);
xnor U21105 (N_21105,N_18027,N_14217);
and U21106 (N_21106,N_19655,N_19011);
nand U21107 (N_21107,N_15452,N_19370);
or U21108 (N_21108,N_14763,N_16282);
nor U21109 (N_21109,N_13102,N_16880);
xnor U21110 (N_21110,N_17779,N_16933);
nor U21111 (N_21111,N_17742,N_17845);
xnor U21112 (N_21112,N_16575,N_16425);
or U21113 (N_21113,N_18814,N_17585);
nand U21114 (N_21114,N_12132,N_10749);
xor U21115 (N_21115,N_15128,N_16711);
nor U21116 (N_21116,N_17399,N_19124);
or U21117 (N_21117,N_11156,N_13631);
nor U21118 (N_21118,N_11920,N_10556);
and U21119 (N_21119,N_12475,N_19827);
or U21120 (N_21120,N_14565,N_14215);
xnor U21121 (N_21121,N_15742,N_12549);
and U21122 (N_21122,N_17967,N_19023);
and U21123 (N_21123,N_18902,N_10756);
and U21124 (N_21124,N_13082,N_17935);
nand U21125 (N_21125,N_17266,N_16345);
xnor U21126 (N_21126,N_12760,N_14393);
xor U21127 (N_21127,N_16041,N_10327);
nand U21128 (N_21128,N_14174,N_17919);
or U21129 (N_21129,N_15439,N_13649);
nand U21130 (N_21130,N_15781,N_15407);
nor U21131 (N_21131,N_13290,N_15480);
xnor U21132 (N_21132,N_12957,N_11390);
or U21133 (N_21133,N_10028,N_13895);
nor U21134 (N_21134,N_13162,N_15107);
nor U21135 (N_21135,N_17981,N_11029);
xnor U21136 (N_21136,N_17181,N_12199);
and U21137 (N_21137,N_17889,N_13576);
and U21138 (N_21138,N_17502,N_18146);
and U21139 (N_21139,N_19547,N_18352);
nand U21140 (N_21140,N_15763,N_13402);
xor U21141 (N_21141,N_16121,N_14518);
nand U21142 (N_21142,N_18073,N_16897);
or U21143 (N_21143,N_18243,N_14133);
nor U21144 (N_21144,N_14082,N_17605);
or U21145 (N_21145,N_15503,N_10993);
and U21146 (N_21146,N_15916,N_17038);
nand U21147 (N_21147,N_16373,N_14636);
or U21148 (N_21148,N_19923,N_16206);
nand U21149 (N_21149,N_14625,N_19993);
or U21150 (N_21150,N_10423,N_18668);
or U21151 (N_21151,N_16144,N_14571);
xor U21152 (N_21152,N_16401,N_12390);
or U21153 (N_21153,N_16141,N_12775);
xnor U21154 (N_21154,N_19102,N_10563);
and U21155 (N_21155,N_19164,N_18356);
nor U21156 (N_21156,N_14808,N_15413);
xor U21157 (N_21157,N_19538,N_10218);
and U21158 (N_21158,N_15671,N_13470);
xor U21159 (N_21159,N_15800,N_13142);
or U21160 (N_21160,N_13651,N_13369);
xnor U21161 (N_21161,N_13253,N_11801);
and U21162 (N_21162,N_19010,N_14658);
nand U21163 (N_21163,N_15481,N_10611);
nor U21164 (N_21164,N_16854,N_15913);
nand U21165 (N_21165,N_10027,N_16754);
nand U21166 (N_21166,N_18578,N_17146);
xor U21167 (N_21167,N_10726,N_15181);
and U21168 (N_21168,N_10408,N_14964);
or U21169 (N_21169,N_18913,N_17256);
nor U21170 (N_21170,N_13599,N_17081);
and U21171 (N_21171,N_17817,N_13978);
and U21172 (N_21172,N_19639,N_11885);
or U21173 (N_21173,N_11764,N_15468);
xnor U21174 (N_21174,N_19800,N_14338);
or U21175 (N_21175,N_19779,N_17866);
or U21176 (N_21176,N_19952,N_18153);
or U21177 (N_21177,N_17369,N_19996);
nor U21178 (N_21178,N_16952,N_16855);
nand U21179 (N_21179,N_16291,N_16252);
nand U21180 (N_21180,N_18587,N_12512);
and U21181 (N_21181,N_18439,N_11515);
and U21182 (N_21182,N_15822,N_16234);
nand U21183 (N_21183,N_17850,N_13375);
nor U21184 (N_21184,N_16549,N_18843);
and U21185 (N_21185,N_16548,N_16261);
and U21186 (N_21186,N_19430,N_13980);
and U21187 (N_21187,N_11970,N_10848);
nand U21188 (N_21188,N_10388,N_17095);
xor U21189 (N_21189,N_19897,N_15537);
or U21190 (N_21190,N_11233,N_14178);
nand U21191 (N_21191,N_18176,N_16650);
nor U21192 (N_21192,N_19684,N_17352);
xnor U21193 (N_21193,N_16712,N_17035);
xnor U21194 (N_21194,N_11409,N_12123);
xor U21195 (N_21195,N_17167,N_10008);
and U21196 (N_21196,N_14741,N_12511);
nand U21197 (N_21197,N_14190,N_15490);
and U21198 (N_21198,N_17347,N_16743);
nand U21199 (N_21199,N_16922,N_11284);
nor U21200 (N_21200,N_19616,N_15491);
nand U21201 (N_21201,N_15387,N_18762);
and U21202 (N_21202,N_15182,N_10120);
nor U21203 (N_21203,N_11909,N_19036);
xor U21204 (N_21204,N_13691,N_12117);
or U21205 (N_21205,N_14532,N_16371);
and U21206 (N_21206,N_15098,N_12219);
and U21207 (N_21207,N_17855,N_15736);
nor U21208 (N_21208,N_18505,N_15841);
and U21209 (N_21209,N_11641,N_16320);
nor U21210 (N_21210,N_17368,N_17134);
nor U21211 (N_21211,N_16175,N_16726);
xnor U21212 (N_21212,N_18052,N_10902);
and U21213 (N_21213,N_11058,N_17202);
nand U21214 (N_21214,N_13884,N_19041);
nand U21215 (N_21215,N_12027,N_16651);
or U21216 (N_21216,N_13003,N_19978);
or U21217 (N_21217,N_18648,N_10780);
nand U21218 (N_21218,N_19529,N_19858);
or U21219 (N_21219,N_12200,N_17474);
or U21220 (N_21220,N_10010,N_11857);
and U21221 (N_21221,N_18416,N_12753);
and U21222 (N_21222,N_16530,N_16878);
nor U21223 (N_21223,N_17801,N_14702);
or U21224 (N_21224,N_12377,N_12860);
and U21225 (N_21225,N_16605,N_12606);
xor U21226 (N_21226,N_12232,N_14085);
nor U21227 (N_21227,N_18452,N_17559);
nand U21228 (N_21228,N_13917,N_18998);
nor U21229 (N_21229,N_17065,N_10998);
nor U21230 (N_21230,N_13147,N_14034);
and U21231 (N_21231,N_12483,N_14650);
or U21232 (N_21232,N_18139,N_19279);
xnor U21233 (N_21233,N_16942,N_12905);
nor U21234 (N_21234,N_11151,N_11182);
and U21235 (N_21235,N_12609,N_18004);
nand U21236 (N_21236,N_14657,N_19481);
xor U21237 (N_21237,N_15999,N_15828);
or U21238 (N_21238,N_18815,N_16950);
or U21239 (N_21239,N_15293,N_13712);
or U21240 (N_21240,N_10051,N_16544);
nand U21241 (N_21241,N_14740,N_17723);
nand U21242 (N_21242,N_18268,N_13079);
or U21243 (N_21243,N_18823,N_12342);
or U21244 (N_21244,N_11673,N_12084);
nand U21245 (N_21245,N_11827,N_18529);
or U21246 (N_21246,N_11276,N_17419);
or U21247 (N_21247,N_19893,N_15918);
xor U21248 (N_21248,N_14521,N_17851);
nand U21249 (N_21249,N_19826,N_18082);
and U21250 (N_21250,N_16460,N_13493);
and U21251 (N_21251,N_11411,N_16051);
or U21252 (N_21252,N_14728,N_13955);
nor U21253 (N_21253,N_16109,N_13894);
nand U21254 (N_21254,N_18399,N_12504);
xor U21255 (N_21255,N_11639,N_19920);
nand U21256 (N_21256,N_13357,N_13185);
nor U21257 (N_21257,N_11046,N_14822);
nor U21258 (N_21258,N_14971,N_13823);
or U21259 (N_21259,N_11380,N_15575);
nand U21260 (N_21260,N_14236,N_19714);
nand U21261 (N_21261,N_14583,N_19646);
or U21262 (N_21262,N_16759,N_12741);
and U21263 (N_21263,N_13407,N_15988);
xnor U21264 (N_21264,N_12412,N_10076);
and U21265 (N_21265,N_19895,N_17595);
nand U21266 (N_21266,N_13891,N_17524);
and U21267 (N_21267,N_10926,N_17544);
nand U21268 (N_21268,N_18475,N_18558);
or U21269 (N_21269,N_19074,N_13432);
nand U21270 (N_21270,N_15492,N_15777);
and U21271 (N_21271,N_11230,N_18057);
or U21272 (N_21272,N_18201,N_10730);
nand U21273 (N_21273,N_18638,N_11335);
and U21274 (N_21274,N_15543,N_14470);
and U21275 (N_21275,N_16626,N_11552);
nor U21276 (N_21276,N_10395,N_11676);
xor U21277 (N_21277,N_13482,N_16396);
or U21278 (N_21278,N_12580,N_10525);
and U21279 (N_21279,N_12724,N_15462);
nand U21280 (N_21280,N_10981,N_16843);
and U21281 (N_21281,N_15442,N_12186);
or U21282 (N_21282,N_15359,N_19685);
nand U21283 (N_21283,N_14963,N_17567);
nor U21284 (N_21284,N_19121,N_19408);
xnor U21285 (N_21285,N_18513,N_10616);
nand U21286 (N_21286,N_10790,N_18140);
and U21287 (N_21287,N_19785,N_19082);
nand U21288 (N_21288,N_14853,N_19896);
and U21289 (N_21289,N_14546,N_11263);
nand U21290 (N_21290,N_19889,N_13939);
and U21291 (N_21291,N_13392,N_15313);
or U21292 (N_21292,N_19393,N_13099);
or U21293 (N_21293,N_16729,N_19935);
nand U21294 (N_21294,N_19359,N_14935);
or U21295 (N_21295,N_13302,N_19721);
and U21296 (N_21296,N_15371,N_16370);
xor U21297 (N_21297,N_19253,N_14454);
xnor U21298 (N_21298,N_14275,N_14084);
or U21299 (N_21299,N_14500,N_10185);
xor U21300 (N_21300,N_16082,N_17555);
and U21301 (N_21301,N_10069,N_15876);
nand U21302 (N_21302,N_13786,N_17082);
and U21303 (N_21303,N_12477,N_11569);
xor U21304 (N_21304,N_16271,N_18735);
and U21305 (N_21305,N_15601,N_15574);
nand U21306 (N_21306,N_15894,N_17709);
nor U21307 (N_21307,N_17328,N_17998);
and U21308 (N_21308,N_14638,N_17949);
and U21309 (N_21309,N_10075,N_10595);
nand U21310 (N_21310,N_18708,N_17831);
or U21311 (N_21311,N_16449,N_14205);
or U21312 (N_21312,N_11590,N_12155);
xnor U21313 (N_21313,N_17951,N_16374);
nand U21314 (N_21314,N_19200,N_14093);
nor U21315 (N_21315,N_19778,N_19316);
and U21316 (N_21316,N_12468,N_17973);
nand U21317 (N_21317,N_16962,N_18011);
nand U21318 (N_21318,N_14854,N_12427);
or U21319 (N_21319,N_14015,N_12353);
xor U21320 (N_21320,N_16891,N_17208);
and U21321 (N_21321,N_12681,N_15859);
xnor U21322 (N_21322,N_10640,N_16850);
xor U21323 (N_21323,N_19558,N_14105);
nand U21324 (N_21324,N_14598,N_16442);
xnor U21325 (N_21325,N_18970,N_10817);
xnor U21326 (N_21326,N_16235,N_19600);
nand U21327 (N_21327,N_13625,N_14634);
nand U21328 (N_21328,N_15479,N_19556);
nand U21329 (N_21329,N_14358,N_11109);
nand U21330 (N_21330,N_13710,N_18017);
xor U21331 (N_21331,N_16205,N_10033);
and U21332 (N_21332,N_12894,N_12796);
nand U21333 (N_21333,N_16839,N_11346);
nor U21334 (N_21334,N_13733,N_12500);
nor U21335 (N_21335,N_10188,N_18618);
or U21336 (N_21336,N_13057,N_13536);
xor U21337 (N_21337,N_16039,N_17765);
nor U21338 (N_21338,N_12479,N_14764);
and U21339 (N_21339,N_14794,N_11997);
xnor U21340 (N_21340,N_19373,N_12577);
nand U21341 (N_21341,N_18121,N_14866);
nor U21342 (N_21342,N_17827,N_19806);
xnor U21343 (N_21343,N_13351,N_16826);
xor U21344 (N_21344,N_18516,N_17965);
xnor U21345 (N_21345,N_19581,N_14905);
or U21346 (N_21346,N_18981,N_13236);
nand U21347 (N_21347,N_11133,N_17329);
nand U21348 (N_21348,N_16292,N_10840);
or U21349 (N_21349,N_10549,N_18144);
xnor U21350 (N_21350,N_17193,N_12977);
or U21351 (N_21351,N_16635,N_16568);
nand U21352 (N_21352,N_14210,N_14881);
and U21353 (N_21353,N_16980,N_14899);
and U21354 (N_21354,N_14250,N_12699);
xor U21355 (N_21355,N_11015,N_13394);
nand U21356 (N_21356,N_17289,N_19518);
nand U21357 (N_21357,N_18051,N_11719);
nor U21358 (N_21358,N_10137,N_12063);
nand U21359 (N_21359,N_18693,N_13591);
nand U21360 (N_21360,N_12847,N_13785);
nand U21361 (N_21361,N_13281,N_14221);
and U21362 (N_21362,N_17271,N_16640);
nor U21363 (N_21363,N_11140,N_18782);
nand U21364 (N_21364,N_13218,N_16968);
xnor U21365 (N_21365,N_16562,N_16118);
xor U21366 (N_21366,N_11318,N_16905);
nand U21367 (N_21367,N_19203,N_15972);
nor U21368 (N_21368,N_10761,N_10417);
xor U21369 (N_21369,N_16219,N_17659);
nor U21370 (N_21370,N_17853,N_13339);
nand U21371 (N_21371,N_19991,N_12676);
xnor U21372 (N_21372,N_11503,N_11055);
nor U21373 (N_21373,N_18594,N_17891);
nor U21374 (N_21374,N_12723,N_16793);
xnor U21375 (N_21375,N_19410,N_14884);
nand U21376 (N_21376,N_18434,N_16285);
and U21377 (N_21377,N_19267,N_10457);
xor U21378 (N_21378,N_19809,N_19211);
nor U21379 (N_21379,N_15507,N_12715);
and U21380 (N_21380,N_16355,N_12447);
xnor U21381 (N_21381,N_19590,N_17933);
nor U21382 (N_21382,N_10460,N_15498);
or U21383 (N_21383,N_15256,N_16343);
nor U21384 (N_21384,N_15984,N_19536);
xnor U21385 (N_21385,N_17665,N_12432);
and U21386 (N_21386,N_19804,N_15053);
and U21387 (N_21387,N_11023,N_14972);
nor U21388 (N_21388,N_10696,N_19506);
and U21389 (N_21389,N_18882,N_13762);
and U21390 (N_21390,N_19875,N_17606);
nand U21391 (N_21391,N_19306,N_15676);
xor U21392 (N_21392,N_15271,N_16902);
and U21393 (N_21393,N_14870,N_18406);
or U21394 (N_21394,N_17562,N_16801);
nor U21395 (N_21395,N_12053,N_11191);
xnor U21396 (N_21396,N_18534,N_15502);
and U21397 (N_21397,N_11837,N_10157);
or U21398 (N_21398,N_11765,N_18435);
nor U21399 (N_21399,N_15025,N_15959);
nand U21400 (N_21400,N_10449,N_11089);
xnor U21401 (N_21401,N_14199,N_12300);
nor U21402 (N_21402,N_19321,N_19150);
and U21403 (N_21403,N_15925,N_16411);
xor U21404 (N_21404,N_18373,N_17582);
and U21405 (N_21405,N_19725,N_17097);
nor U21406 (N_21406,N_17386,N_18793);
xnor U21407 (N_21407,N_12431,N_10802);
xnor U21408 (N_21408,N_11506,N_14067);
or U21409 (N_21409,N_13876,N_15385);
or U21410 (N_21410,N_18414,N_11973);
nand U21411 (N_21411,N_14603,N_10057);
or U21412 (N_21412,N_11348,N_10531);
nand U21413 (N_21413,N_12079,N_13926);
xnor U21414 (N_21414,N_18586,N_14324);
or U21415 (N_21415,N_12049,N_12642);
or U21416 (N_21416,N_19213,N_19814);
nor U21417 (N_21417,N_13056,N_11157);
nor U21418 (N_21418,N_13009,N_15043);
xnor U21419 (N_21419,N_17806,N_11173);
nand U21420 (N_21420,N_15665,N_16509);
or U21421 (N_21421,N_14876,N_18621);
xnor U21422 (N_21422,N_14000,N_15404);
and U21423 (N_21423,N_13540,N_11854);
and U21424 (N_21424,N_11002,N_11048);
xor U21425 (N_21425,N_19502,N_12744);
nor U21426 (N_21426,N_12648,N_12993);
and U21427 (N_21427,N_16237,N_13174);
or U21428 (N_21428,N_19020,N_18179);
or U21429 (N_21429,N_13795,N_14769);
and U21430 (N_21430,N_14819,N_12656);
nand U21431 (N_21431,N_16723,N_19734);
and U21432 (N_21432,N_12469,N_19634);
xor U21433 (N_21433,N_13010,N_10854);
xnor U21434 (N_21434,N_16001,N_13767);
and U21435 (N_21435,N_16761,N_17963);
or U21436 (N_21436,N_15947,N_13905);
nor U21437 (N_21437,N_18120,N_11211);
xor U21438 (N_21438,N_14089,N_17748);
nor U21439 (N_21439,N_13190,N_19360);
or U21440 (N_21440,N_15980,N_10308);
nor U21441 (N_21441,N_16647,N_16267);
and U21442 (N_21442,N_14179,N_19726);
or U21443 (N_21443,N_18332,N_12664);
xor U21444 (N_21444,N_19693,N_18209);
or U21445 (N_21445,N_14410,N_11258);
or U21446 (N_21446,N_16906,N_14074);
or U21447 (N_21447,N_18486,N_10368);
nand U21448 (N_21448,N_12401,N_11743);
nand U21449 (N_21449,N_16877,N_17055);
nor U21450 (N_21450,N_11834,N_16469);
nor U21451 (N_21451,N_12288,N_13607);
nor U21452 (N_21452,N_13873,N_17044);
and U21453 (N_21453,N_17070,N_13679);
or U21454 (N_21454,N_10888,N_11357);
nand U21455 (N_21455,N_16133,N_19463);
nor U21456 (N_21456,N_15298,N_16068);
nor U21457 (N_21457,N_11441,N_15243);
and U21458 (N_21458,N_14776,N_18582);
xor U21459 (N_21459,N_12685,N_19953);
or U21460 (N_21460,N_11795,N_12157);
nand U21461 (N_21461,N_17447,N_16337);
nor U21462 (N_21462,N_15852,N_12535);
nand U21463 (N_21463,N_10490,N_11736);
or U21464 (N_21464,N_12743,N_10748);
nor U21465 (N_21465,N_10437,N_15062);
nor U21466 (N_21466,N_11084,N_15526);
xor U21467 (N_21467,N_12481,N_17359);
nand U21468 (N_21468,N_10778,N_11466);
or U21469 (N_21469,N_10585,N_15592);
nor U21470 (N_21470,N_15150,N_14315);
and U21471 (N_21471,N_18886,N_18788);
and U21472 (N_21472,N_15795,N_13140);
or U21473 (N_21473,N_13000,N_10612);
or U21474 (N_21474,N_10210,N_16534);
and U21475 (N_21475,N_15621,N_10174);
nor U21476 (N_21476,N_17221,N_15704);
nand U21477 (N_21477,N_18935,N_19647);
and U21478 (N_21478,N_19847,N_11255);
or U21479 (N_21479,N_19788,N_10336);
nand U21480 (N_21480,N_16066,N_14043);
xnor U21481 (N_21481,N_14952,N_14659);
or U21482 (N_21482,N_14274,N_10288);
xnor U21483 (N_21483,N_18826,N_14276);
or U21484 (N_21484,N_14810,N_12689);
nor U21485 (N_21485,N_15199,N_11763);
xnor U21486 (N_21486,N_16259,N_18603);
xnor U21487 (N_21487,N_18927,N_10642);
or U21488 (N_21488,N_11431,N_10429);
xor U21489 (N_21489,N_11770,N_15210);
and U21490 (N_21490,N_11083,N_11858);
nand U21491 (N_21491,N_11492,N_17519);
nand U21492 (N_21492,N_17389,N_13615);
and U21493 (N_21493,N_18599,N_11060);
nand U21494 (N_21494,N_13820,N_18263);
nor U21495 (N_21495,N_19739,N_11984);
xnor U21496 (N_21496,N_12415,N_12995);
nor U21497 (N_21497,N_17174,N_10844);
nand U21498 (N_21498,N_11234,N_15924);
xor U21499 (N_21499,N_16604,N_13896);
xor U21500 (N_21500,N_14772,N_12153);
or U21501 (N_21501,N_16161,N_15589);
xor U21502 (N_21502,N_16803,N_12665);
nand U21503 (N_21503,N_13083,N_17902);
and U21504 (N_21504,N_11619,N_15529);
xor U21505 (N_21505,N_15166,N_18760);
xor U21506 (N_21506,N_16334,N_14226);
xnor U21507 (N_21507,N_13054,N_18544);
nor U21508 (N_21508,N_15653,N_13956);
xnor U21509 (N_21509,N_18442,N_17244);
nor U21510 (N_21510,N_13154,N_10712);
or U21511 (N_21511,N_15290,N_15544);
xor U21512 (N_21512,N_17138,N_18512);
xor U21513 (N_21513,N_16017,N_11752);
nand U21514 (N_21514,N_19034,N_14557);
nand U21515 (N_21515,N_16934,N_18588);
xnor U21516 (N_21516,N_16872,N_15939);
and U21517 (N_21517,N_16419,N_19970);
nand U21518 (N_21518,N_17794,N_19112);
xor U21519 (N_21519,N_17620,N_14346);
nor U21520 (N_21520,N_13889,N_14412);
nand U21521 (N_21521,N_13554,N_15525);
and U21522 (N_21522,N_13510,N_13606);
or U21523 (N_21523,N_18040,N_13774);
and U21524 (N_21524,N_19554,N_19839);
nor U21525 (N_21525,N_10995,N_11033);
and U21526 (N_21526,N_14989,N_14545);
nor U21527 (N_21527,N_10676,N_12192);
or U21528 (N_21528,N_16917,N_16510);
xnor U21529 (N_21529,N_17961,N_18074);
xnor U21530 (N_21530,N_13410,N_13764);
nor U21531 (N_21531,N_11362,N_10648);
or U21532 (N_21532,N_18867,N_13077);
or U21533 (N_21533,N_14440,N_18046);
and U21534 (N_21534,N_10855,N_17125);
xnor U21535 (N_21535,N_12020,N_16018);
and U21536 (N_21536,N_16738,N_12136);
nor U21537 (N_21537,N_18193,N_11947);
xor U21538 (N_21538,N_11190,N_12229);
nor U21539 (N_21539,N_11870,N_17766);
nor U21540 (N_21540,N_19400,N_12051);
xor U21541 (N_21541,N_19143,N_10163);
xor U21542 (N_21542,N_18745,N_15607);
nor U21543 (N_21543,N_12958,N_15807);
nand U21544 (N_21544,N_12732,N_16342);
and U21545 (N_21545,N_15459,N_15324);
nor U21546 (N_21546,N_19620,N_12223);
xor U21547 (N_21547,N_14760,N_17604);
or U21548 (N_21548,N_19484,N_10650);
nand U21549 (N_21549,N_17830,N_13358);
nor U21550 (N_21550,N_18087,N_13200);
or U21551 (N_21551,N_19318,N_15227);
or U21552 (N_21552,N_14024,N_12837);
nor U21553 (N_21553,N_12569,N_11518);
xnor U21554 (N_21554,N_18765,N_14039);
and U21555 (N_21555,N_14252,N_14343);
and U21556 (N_21556,N_14651,N_13832);
and U21557 (N_21557,N_16153,N_18289);
and U21558 (N_21558,N_19808,N_19209);
nor U21559 (N_21559,N_13719,N_19829);
and U21560 (N_21560,N_14501,N_19295);
xnor U21561 (N_21561,N_14832,N_15827);
or U21562 (N_21562,N_17970,N_17681);
xnor U21563 (N_21563,N_13948,N_10607);
or U21564 (N_21564,N_11461,N_19106);
and U21565 (N_21565,N_16518,N_13216);
xnor U21566 (N_21566,N_15522,N_12396);
and U21567 (N_21567,N_18110,N_12799);
or U21568 (N_21568,N_10689,N_13203);
nor U21569 (N_21569,N_19775,N_16631);
nor U21570 (N_21570,N_15092,N_18897);
nand U21571 (N_21571,N_16632,N_13487);
nor U21572 (N_21572,N_17494,N_16500);
and U21573 (N_21573,N_11714,N_19090);
nand U21574 (N_21574,N_15200,N_11118);
nand U21575 (N_21575,N_18642,N_12550);
xor U21576 (N_21576,N_17345,N_17594);
and U21577 (N_21577,N_15838,N_11397);
xnor U21578 (N_21578,N_16458,N_13500);
nor U21579 (N_21579,N_10800,N_17915);
nand U21580 (N_21580,N_12687,N_10340);
nand U21581 (N_21581,N_12879,N_18272);
nor U21582 (N_21582,N_15718,N_19261);
nor U21583 (N_21583,N_19700,N_14100);
or U21584 (N_21584,N_15125,N_19951);
nor U21585 (N_21585,N_17596,N_15096);
xnor U21586 (N_21586,N_12804,N_17092);
nor U21587 (N_21587,N_10795,N_15593);
and U21588 (N_21588,N_17226,N_11090);
or U21589 (N_21589,N_18908,N_18150);
nand U21590 (N_21590,N_10418,N_17746);
or U21591 (N_21591,N_17823,N_16366);
or U21592 (N_21592,N_19731,N_15161);
nor U21593 (N_21593,N_10400,N_16163);
nand U21594 (N_21594,N_11000,N_15964);
nand U21595 (N_21595,N_12052,N_11930);
nand U21596 (N_21596,N_19173,N_15093);
and U21597 (N_21597,N_19776,N_12190);
or U21598 (N_21598,N_17466,N_17534);
nand U21599 (N_21599,N_19844,N_17896);
xnor U21600 (N_21600,N_12987,N_19642);
and U21601 (N_21601,N_19031,N_15122);
nand U21602 (N_21602,N_16088,N_17539);
or U21603 (N_21603,N_12105,N_18822);
or U21604 (N_21604,N_13238,N_16835);
and U21605 (N_21605,N_19811,N_17046);
and U21606 (N_21606,N_10351,N_17140);
and U21607 (N_21607,N_13513,N_19988);
and U21608 (N_21608,N_10683,N_14824);
nor U21609 (N_21609,N_10329,N_10118);
xor U21610 (N_21610,N_14936,N_15448);
nand U21611 (N_21611,N_19651,N_13888);
or U21612 (N_21612,N_16023,N_11611);
xor U21613 (N_21613,N_16806,N_12964);
xor U21614 (N_21614,N_13665,N_17478);
nand U21615 (N_21615,N_13366,N_17117);
or U21616 (N_21616,N_12133,N_11498);
and U21617 (N_21617,N_14155,N_15039);
nand U21618 (N_21618,N_17513,N_12836);
nand U21619 (N_21619,N_17776,N_17003);
xor U21620 (N_21620,N_19641,N_15504);
or U21621 (N_21621,N_14029,N_17496);
nand U21622 (N_21622,N_16658,N_14400);
nand U21623 (N_21623,N_12160,N_17825);
xor U21624 (N_21624,N_13453,N_11603);
nand U21625 (N_21625,N_16753,N_16043);
xnor U21626 (N_21626,N_12221,N_12791);
nand U21627 (N_21627,N_14428,N_10688);
xnor U21628 (N_21628,N_14699,N_13883);
or U21629 (N_21629,N_10399,N_14357);
nor U21630 (N_21630,N_10123,N_12943);
or U21631 (N_21631,N_17377,N_10554);
and U21632 (N_21632,N_12772,N_16846);
or U21633 (N_21633,N_14830,N_10426);
or U21634 (N_21634,N_17738,N_10564);
or U21635 (N_21635,N_15769,N_12798);
nor U21636 (N_21636,N_13173,N_16388);
or U21637 (N_21637,N_16554,N_14351);
nor U21638 (N_21638,N_13975,N_12043);
xor U21639 (N_21639,N_17311,N_15833);
xor U21640 (N_21640,N_10117,N_18584);
nand U21641 (N_21641,N_15138,N_16848);
xor U21642 (N_21642,N_12565,N_12915);
or U21643 (N_21643,N_16814,N_19223);
xnor U21644 (N_21644,N_17486,N_15986);
nand U21645 (N_21645,N_10014,N_11373);
nand U21646 (N_21646,N_11908,N_18492);
or U21647 (N_21647,N_18354,N_11473);
xor U21648 (N_21648,N_11899,N_13718);
nand U21649 (N_21649,N_19182,N_15360);
nor U21650 (N_21650,N_15441,N_11166);
and U21651 (N_21651,N_10577,N_19946);
and U21652 (N_21652,N_13406,N_15878);
nor U21653 (N_21653,N_14744,N_13350);
nand U21654 (N_21654,N_19027,N_16020);
nand U21655 (N_21655,N_13335,N_16900);
nor U21656 (N_21656,N_11879,N_11845);
and U21657 (N_21657,N_10896,N_14648);
xnor U21658 (N_21658,N_10508,N_13217);
and U21659 (N_21659,N_17834,N_14900);
nor U21660 (N_21660,N_19479,N_19248);
xnor U21661 (N_21661,N_10496,N_18056);
xnor U21662 (N_21662,N_18919,N_16119);
nand U21663 (N_21663,N_18157,N_14489);
nand U21664 (N_21664,N_18895,N_11097);
xnor U21665 (N_21665,N_13159,N_17704);
nand U21666 (N_21666,N_13067,N_17233);
xnor U21667 (N_21667,N_12570,N_19543);
or U21668 (N_21668,N_14746,N_19219);
nand U21669 (N_21669,N_14066,N_18312);
nand U21670 (N_21670,N_11006,N_18105);
nor U21671 (N_21671,N_18331,N_13986);
and U21672 (N_21672,N_19093,N_12619);
nand U21673 (N_21673,N_17838,N_13743);
or U21674 (N_21674,N_13614,N_13443);
nand U21675 (N_21675,N_14196,N_19763);
or U21676 (N_21676,N_12406,N_15068);
or U21677 (N_21677,N_14887,N_10628);
nor U21678 (N_21678,N_13028,N_19266);
xnor U21679 (N_21679,N_15706,N_18983);
nand U21680 (N_21680,N_16620,N_19990);
or U21681 (N_21681,N_18656,N_11892);
nand U21682 (N_21682,N_19624,N_17575);
and U21683 (N_21683,N_15011,N_14207);
or U21684 (N_21684,N_14503,N_11462);
and U21685 (N_21685,N_10445,N_16879);
nand U21686 (N_21686,N_16730,N_13880);
and U21687 (N_21687,N_10983,N_12227);
and U21688 (N_21688,N_13005,N_18010);
or U21689 (N_21689,N_12305,N_12421);
or U21690 (N_21690,N_10724,N_19928);
xnor U21691 (N_21691,N_18091,N_16201);
xor U21692 (N_21692,N_17561,N_19977);
xor U21693 (N_21693,N_16126,N_17954);
and U21694 (N_21694,N_16545,N_13996);
and U21695 (N_21695,N_11236,N_17147);
xor U21696 (N_21696,N_19653,N_11321);
nor U21697 (N_21697,N_19208,N_17824);
nor U21698 (N_21698,N_18846,N_19363);
nand U21699 (N_21699,N_16179,N_13997);
nand U21700 (N_21700,N_13356,N_10223);
nand U21701 (N_21701,N_10106,N_16797);
xor U21702 (N_21702,N_18975,N_19427);
and U21703 (N_21703,N_12954,N_10523);
nand U21704 (N_21704,N_14893,N_19085);
nor U21705 (N_21705,N_16412,N_16507);
nor U21706 (N_21706,N_19580,N_11223);
and U21707 (N_21707,N_19345,N_16217);
nor U21708 (N_21708,N_11124,N_17360);
nand U21709 (N_21709,N_13662,N_17214);
nand U21710 (N_21710,N_16172,N_12670);
nor U21711 (N_21711,N_14462,N_13816);
and U21712 (N_21712,N_13551,N_15992);
and U21713 (N_21713,N_17155,N_14314);
and U21714 (N_21714,N_13039,N_17007);
nor U21715 (N_21715,N_13464,N_13143);
xnor U21716 (N_21716,N_11607,N_10924);
nor U21717 (N_21717,N_16576,N_10514);
nor U21718 (N_21718,N_19406,N_12766);
nand U21719 (N_21719,N_16166,N_18385);
xor U21720 (N_21720,N_10699,N_13708);
and U21721 (N_21721,N_18880,N_13045);
xnor U21722 (N_21722,N_15796,N_13566);
nand U21723 (N_21723,N_19170,N_17865);
and U21724 (N_21724,N_14790,N_12946);
nor U21725 (N_21725,N_11486,N_10502);
and U21726 (N_21726,N_13911,N_12099);
or U21727 (N_21727,N_12582,N_17331);
or U21728 (N_21728,N_19068,N_10234);
nor U21729 (N_21729,N_14434,N_10675);
or U21730 (N_21730,N_13857,N_18386);
nor U21731 (N_21731,N_19153,N_12257);
nand U21732 (N_21732,N_15991,N_16169);
nor U21733 (N_21733,N_16988,N_13169);
xor U21734 (N_21734,N_17775,N_16505);
xor U21735 (N_21735,N_13514,N_17584);
nor U21736 (N_21736,N_13104,N_16532);
nor U21737 (N_21737,N_11831,N_18280);
or U21738 (N_21738,N_12014,N_10101);
xnor U21739 (N_21739,N_19327,N_19128);
and U21740 (N_21740,N_18715,N_17264);
and U21741 (N_21741,N_15337,N_16327);
or U21742 (N_21742,N_11757,N_10433);
xnor U21743 (N_21743,N_13181,N_18402);
nand U21744 (N_21744,N_10668,N_15224);
xor U21745 (N_21745,N_10100,N_18463);
nand U21746 (N_21746,N_12970,N_19549);
and U21747 (N_21747,N_10827,N_10764);
nor U21748 (N_21748,N_11172,N_18776);
nand U21749 (N_21749,N_16751,N_14695);
or U21750 (N_21750,N_16230,N_15052);
xor U21751 (N_21751,N_11593,N_15139);
and U21752 (N_21752,N_19738,N_12409);
and U21753 (N_21753,N_18485,N_17168);
nor U21754 (N_21754,N_13498,N_18053);
nand U21755 (N_21755,N_18238,N_12739);
or U21756 (N_21756,N_19533,N_11898);
nand U21757 (N_21757,N_15145,N_19837);
nor U21758 (N_21758,N_13608,N_12170);
xnor U21759 (N_21759,N_19962,N_15615);
nor U21760 (N_21760,N_17145,N_19457);
or U21761 (N_21761,N_10309,N_19325);
xnor U21762 (N_21762,N_19446,N_17028);
or U21763 (N_21763,N_19382,N_19021);
nand U21764 (N_21764,N_12077,N_14707);
and U21765 (N_21765,N_14111,N_15605);
xnor U21766 (N_21766,N_17912,N_15663);
and U21767 (N_21767,N_13724,N_11635);
nor U21768 (N_21768,N_16672,N_15571);
or U21769 (N_21769,N_17630,N_16750);
nor U21770 (N_21770,N_18984,N_13497);
and U21771 (N_21771,N_14162,N_18415);
xor U21772 (N_21772,N_10954,N_12769);
or U21773 (N_21773,N_17467,N_19850);
nor U21774 (N_21774,N_15661,N_19522);
nand U21775 (N_21775,N_13668,N_15554);
or U21776 (N_21776,N_14943,N_12314);
nand U21777 (N_21777,N_18769,N_12782);
and U21778 (N_21778,N_12331,N_16965);
nor U21779 (N_21779,N_15188,N_19052);
nand U21780 (N_21780,N_11556,N_19322);
nor U21781 (N_21781,N_11251,N_19545);
nand U21782 (N_21782,N_16400,N_11241);
or U21783 (N_21783,N_10853,N_17811);
or U21784 (N_21784,N_12090,N_15612);
nor U21785 (N_21785,N_11861,N_18393);
and U21786 (N_21786,N_15651,N_15799);
and U21787 (N_21787,N_16491,N_13670);
nand U21788 (N_21788,N_10539,N_11938);
xnor U21789 (N_21789,N_19617,N_19652);
or U21790 (N_21790,N_10280,N_10644);
and U21791 (N_21791,N_10686,N_10971);
or U21792 (N_21792,N_10198,N_18247);
xnor U21793 (N_21793,N_11994,N_19276);
nand U21794 (N_21794,N_12735,N_18128);
nor U21795 (N_21795,N_17364,N_10310);
nor U21796 (N_21796,N_13170,N_19877);
nor U21797 (N_21797,N_15352,N_13741);
and U21798 (N_21798,N_10042,N_17390);
nor U21799 (N_21799,N_18921,N_17842);
and U21800 (N_21800,N_16305,N_18327);
nand U21801 (N_21801,N_12655,N_13287);
xnor U21802 (N_21802,N_16247,N_17173);
or U21803 (N_21803,N_17185,N_17305);
and U21804 (N_21804,N_16989,N_19753);
nand U21805 (N_21805,N_18627,N_10136);
xor U21806 (N_21806,N_12413,N_17988);
and U21807 (N_21807,N_10141,N_13757);
nor U21808 (N_21808,N_16489,N_19790);
or U21809 (N_21809,N_16432,N_18980);
and U21810 (N_21810,N_16819,N_13930);
and U21811 (N_21811,N_13435,N_13022);
or U21812 (N_21812,N_17072,N_11841);
nand U21813 (N_21813,N_19076,N_17370);
or U21814 (N_21814,N_12442,N_12994);
nand U21815 (N_21815,N_19297,N_17821);
nand U21816 (N_21816,N_11279,N_16266);
nand U21817 (N_21817,N_17550,N_14996);
or U21818 (N_21818,N_16657,N_18299);
or U21819 (N_21819,N_12100,N_15036);
and U21820 (N_21820,N_19228,N_11427);
xnor U21821 (N_21821,N_12129,N_10084);
and U21822 (N_21822,N_10143,N_12371);
xor U21823 (N_21823,N_18803,N_18503);
xnor U21824 (N_21824,N_13700,N_15454);
or U21825 (N_21825,N_17432,N_10908);
nor U21826 (N_21826,N_14404,N_10434);
nand U21827 (N_21827,N_17553,N_13828);
xnor U21828 (N_21828,N_10856,N_16131);
nor U21829 (N_21829,N_18979,N_18950);
nand U21830 (N_21830,N_12794,N_15072);
or U21831 (N_21831,N_10591,N_10312);
nand U21832 (N_21832,N_14355,N_19610);
xor U21833 (N_21833,N_16957,N_17668);
or U21834 (N_21834,N_17583,N_14775);
nand U21835 (N_21835,N_10885,N_19510);
and U21836 (N_21836,N_12480,N_13534);
or U21837 (N_21837,N_16019,N_16241);
nor U21838 (N_21838,N_15754,N_19451);
xor U21839 (N_21839,N_18321,N_17346);
nor U21840 (N_21840,N_14645,N_19835);
nand U21841 (N_21841,N_10609,N_12047);
nor U21842 (N_21842,N_18829,N_14922);
or U21843 (N_21843,N_17980,N_10353);
and U21844 (N_21844,N_19530,N_10476);
or U21845 (N_21845,N_10936,N_19385);
xor U21846 (N_21846,N_16929,N_16250);
and U21847 (N_21847,N_12101,N_14820);
nand U21848 (N_21848,N_12800,N_11751);
nand U21849 (N_21849,N_17361,N_17250);
nand U21850 (N_21850,N_11280,N_17238);
and U21851 (N_21851,N_19268,N_15914);
xnor U21852 (N_21852,N_13087,N_15008);
xnor U21853 (N_21853,N_17182,N_14931);
xor U21854 (N_21854,N_12936,N_12237);
and U21855 (N_21855,N_18383,N_18412);
nand U21856 (N_21856,N_14263,N_13999);
and U21857 (N_21857,N_19123,N_13477);
nor U21858 (N_21858,N_19876,N_19414);
nor U21859 (N_21859,N_17408,N_10139);
nand U21860 (N_21860,N_16669,N_16642);
or U21861 (N_21861,N_10822,N_12945);
nand U21862 (N_21862,N_13912,N_14156);
and U21863 (N_21863,N_10528,N_18924);
nand U21864 (N_21864,N_16398,N_15196);
or U21865 (N_21865,N_16602,N_11643);
nor U21866 (N_21866,N_12718,N_13006);
nor U21867 (N_21867,N_18468,N_12379);
nand U21868 (N_21868,N_19722,N_11883);
nand U21869 (N_21869,N_13117,N_11903);
or U21870 (N_21870,N_18510,N_15073);
or U21871 (N_21871,N_18732,N_10697);
nor U21872 (N_21872,N_17684,N_13153);
or U21873 (N_21873,N_17240,N_11811);
or U21874 (N_21874,N_19303,N_18821);
or U21875 (N_21875,N_15192,N_11592);
nand U21876 (N_21876,N_13134,N_10709);
nor U21877 (N_21877,N_18947,N_11317);
and U21878 (N_21878,N_18917,N_17637);
or U21879 (N_21879,N_13819,N_13107);
nor U21880 (N_21880,N_19783,N_17813);
xor U21881 (N_21881,N_16105,N_10992);
and U21882 (N_21882,N_18559,N_15301);
or U21883 (N_21883,N_11755,N_15264);
xnor U21884 (N_21884,N_11474,N_11661);
or U21885 (N_21885,N_14629,N_14239);
nor U21886 (N_21886,N_16560,N_12652);
nor U21887 (N_21887,N_10777,N_18628);
and U21888 (N_21888,N_18665,N_10166);
nand U21889 (N_21889,N_16567,N_13158);
nand U21890 (N_21890,N_18949,N_14036);
and U21891 (N_21891,N_18318,N_16324);
and U21892 (N_21892,N_10839,N_11824);
xnor U21893 (N_21893,N_17800,N_10222);
xnor U21894 (N_21894,N_17573,N_12872);
nand U21895 (N_21895,N_15627,N_14469);
and U21896 (N_21896,N_10078,N_12506);
or U21897 (N_21897,N_18806,N_10116);
xnor U21898 (N_21898,N_19552,N_11766);
and U21899 (N_21899,N_17975,N_14902);
xor U21900 (N_21900,N_10273,N_19511);
nor U21901 (N_21901,N_13342,N_10716);
xor U21902 (N_21902,N_15867,N_12011);
nor U21903 (N_21903,N_12857,N_16974);
or U21904 (N_21904,N_17615,N_15477);
nand U21905 (N_21905,N_19792,N_10019);
xnor U21906 (N_21906,N_18200,N_18611);
nor U21907 (N_21907,N_11750,N_12714);
and U21908 (N_21908,N_10499,N_18069);
or U21909 (N_21909,N_10258,N_13539);
and U21910 (N_21910,N_12416,N_10242);
or U21911 (N_21911,N_14706,N_16670);
or U21912 (N_21912,N_15750,N_11306);
and U21913 (N_21913,N_12198,N_10464);
xnor U21914 (N_21914,N_11887,N_10128);
and U21915 (N_21915,N_16523,N_19289);
or U21916 (N_21916,N_12677,N_13761);
nor U21917 (N_21917,N_11702,N_15790);
nand U21918 (N_21918,N_17349,N_10594);
nand U21919 (N_21919,N_16353,N_12768);
nand U21920 (N_21920,N_14908,N_13575);
nand U21921 (N_21921,N_13304,N_16573);
nor U21922 (N_21922,N_15214,N_17564);
and U21923 (N_21923,N_10861,N_10625);
or U21924 (N_21924,N_17677,N_13225);
xnor U21925 (N_21925,N_15408,N_18629);
nand U21926 (N_21926,N_13433,N_16539);
nand U21927 (N_21927,N_13618,N_18554);
or U21928 (N_21928,N_13390,N_15304);
and U21929 (N_21929,N_12030,N_13272);
xnor U21930 (N_21930,N_11426,N_19831);
or U21931 (N_21931,N_16847,N_12383);
nand U21932 (N_21932,N_12264,N_16313);
nor U21933 (N_21933,N_17696,N_18944);
xnor U21934 (N_21934,N_13334,N_14987);
nor U21935 (N_21935,N_15220,N_18494);
or U21936 (N_21936,N_12719,N_17141);
xnor U21937 (N_21937,N_13503,N_18690);
nor U21938 (N_21938,N_14676,N_12308);
and U21939 (N_21939,N_16415,N_14433);
xnor U21940 (N_21940,N_12571,N_10104);
xnor U21941 (N_21941,N_14934,N_14420);
or U21942 (N_21942,N_15019,N_16137);
nor U21943 (N_21943,N_11444,N_13095);
and U21944 (N_21944,N_16326,N_11939);
xor U21945 (N_21945,N_14798,N_13314);
nand U21946 (N_21946,N_18260,N_18905);
nand U21947 (N_21947,N_15027,N_18316);
and U21948 (N_21948,N_16471,N_16239);
and U21949 (N_21949,N_19341,N_16521);
xnor U21950 (N_21950,N_13415,N_10170);
nor U21951 (N_21951,N_16931,N_14513);
or U21952 (N_21952,N_14523,N_10286);
nand U21953 (N_21953,N_11826,N_16484);
nand U21954 (N_21954,N_10968,N_18127);
or U21955 (N_21955,N_12686,N_18381);
or U21956 (N_21956,N_11852,N_10454);
nor U21957 (N_21957,N_19537,N_18104);
and U21958 (N_21958,N_19364,N_12345);
nand U21959 (N_21959,N_18215,N_13299);
xor U21960 (N_21960,N_15650,N_19156);
nor U21961 (N_21961,N_18029,N_11816);
nor U21962 (N_21962,N_11425,N_13885);
nor U21963 (N_21963,N_13454,N_19094);
nand U21964 (N_21964,N_15949,N_17986);
nor U21965 (N_21965,N_10453,N_19244);
nor U21966 (N_21966,N_13837,N_17640);
nand U21967 (N_21967,N_12109,N_16262);
and U21968 (N_21968,N_14856,N_14030);
or U21969 (N_21969,N_13701,N_15273);
and U21970 (N_21970,N_18240,N_14431);
xnor U21971 (N_21971,N_10097,N_15436);
nor U21972 (N_21972,N_17641,N_18334);
and U21973 (N_21973,N_18573,N_14901);
or U21974 (N_21974,N_15299,N_18297);
nor U21975 (N_21975,N_17085,N_18653);
xnor U21976 (N_21976,N_18230,N_19462);
nand U21977 (N_21977,N_11520,N_12022);
xnor U21978 (N_21978,N_11332,N_18118);
and U21979 (N_21979,N_13969,N_13247);
nand U21980 (N_21980,N_11617,N_16447);
nor U21981 (N_21981,N_12975,N_10023);
and U21982 (N_21982,N_13918,N_19254);
nand U21983 (N_21983,N_10317,N_11867);
xor U21984 (N_21984,N_11106,N_10387);
and U21985 (N_21985,N_14828,N_16954);
xnor U21986 (N_21986,N_16511,N_17282);
or U21987 (N_21987,N_14399,N_10125);
or U21988 (N_21988,N_12507,N_19900);
nand U21989 (N_21989,N_12297,N_14685);
and U21990 (N_21990,N_17177,N_12463);
xnor U21991 (N_21991,N_10892,N_19517);
nand U21992 (N_21992,N_19335,N_13810);
or U21993 (N_21993,N_16794,N_15335);
nand U21994 (N_21994,N_18525,N_13847);
or U21995 (N_21995,N_17446,N_13441);
xnor U21996 (N_21996,N_17512,N_16981);
and U21997 (N_21997,N_14246,N_15193);
nor U21998 (N_21998,N_16111,N_10190);
xor U21999 (N_21999,N_13333,N_13172);
and U22000 (N_22000,N_14310,N_12166);
and U22001 (N_22001,N_10923,N_18488);
xnor U22002 (N_22002,N_19555,N_11445);
nor U22003 (N_22003,N_11197,N_10507);
nor U22004 (N_22004,N_12776,N_19799);
or U22005 (N_22005,N_16776,N_10927);
nand U22006 (N_22006,N_13192,N_14295);
xor U22007 (N_22007,N_14560,N_15915);
nor U22008 (N_22008,N_14375,N_18047);
and U22009 (N_22009,N_13188,N_10879);
and U22010 (N_22010,N_19304,N_19609);
or U22011 (N_22011,N_17245,N_19399);
or U22012 (N_22012,N_10184,N_12696);
and U22013 (N_22013,N_19047,N_13380);
and U22014 (N_22014,N_12856,N_19426);
or U22015 (N_22015,N_13038,N_16199);
nor U22016 (N_22016,N_17747,N_10948);
or U22017 (N_22017,N_11507,N_16331);
or U22018 (N_22018,N_16286,N_11772);
or U22019 (N_22019,N_15560,N_15587);
nor U22020 (N_22020,N_19908,N_14019);
nand U22021 (N_22021,N_15902,N_13261);
nor U22022 (N_22022,N_14642,N_12691);
and U22023 (N_22023,N_13090,N_14525);
and U22024 (N_22024,N_14001,N_16923);
nor U22025 (N_22025,N_17798,N_15270);
and U22026 (N_22026,N_13973,N_10239);
nor U22027 (N_22027,N_12335,N_16423);
nand U22028 (N_22028,N_19947,N_14439);
and U22029 (N_22029,N_15509,N_19379);
xor U22030 (N_22030,N_12291,N_17069);
or U22031 (N_22031,N_18527,N_17685);
nor U22032 (N_22032,N_11358,N_13150);
xnor U22033 (N_22033,N_16572,N_16227);
nand U22034 (N_22034,N_14904,N_12505);
and U22035 (N_22035,N_15341,N_14370);
and U22036 (N_22036,N_12207,N_15672);
or U22037 (N_22037,N_19468,N_16908);
or U22038 (N_22038,N_18071,N_11523);
or U22039 (N_22039,N_19710,N_13048);
nand U22040 (N_22040,N_15880,N_14715);
and U22041 (N_22041,N_14309,N_17018);
or U22042 (N_22042,N_14176,N_17822);
nand U22043 (N_22043,N_16470,N_18661);
and U22044 (N_22044,N_19392,N_18164);
xnor U22045 (N_22045,N_13050,N_11684);
nand U22046 (N_22046,N_13199,N_16498);
nand U22047 (N_22047,N_17642,N_16744);
xnor U22048 (N_22048,N_18015,N_13103);
or U22049 (N_22049,N_18585,N_16184);
nor U22050 (N_22050,N_19077,N_18881);
nor U22051 (N_22051,N_14703,N_11821);
and U22052 (N_22052,N_10095,N_17629);
and U22053 (N_22053,N_12488,N_10634);
or U22054 (N_22054,N_14969,N_17947);
nor U22055 (N_22055,N_19079,N_14010);
nand U22056 (N_22056,N_16596,N_16653);
and U22057 (N_22057,N_10704,N_14266);
xor U22058 (N_22058,N_19504,N_14809);
nor U22059 (N_22059,N_12544,N_14078);
xor U22060 (N_22060,N_11032,N_16171);
nor U22061 (N_22061,N_10974,N_17760);
or U22062 (N_22062,N_18390,N_14022);
nand U22063 (N_22063,N_19904,N_18191);
and U22064 (N_22064,N_15694,N_16080);
and U22065 (N_22065,N_13897,N_15026);
xnor U22066 (N_22066,N_10479,N_17110);
nor U22067 (N_22067,N_12567,N_11305);
xnor U22068 (N_22068,N_14782,N_19735);
or U22069 (N_22069,N_11040,N_14426);
xor U22070 (N_22070,N_12078,N_12920);
nor U22071 (N_22071,N_10705,N_10796);
xnor U22072 (N_22072,N_12261,N_11597);
xnor U22073 (N_22073,N_11594,N_17170);
or U22074 (N_22074,N_14455,N_11700);
xor U22075 (N_22075,N_10480,N_15770);
and U22076 (N_22076,N_19903,N_18579);
or U22077 (N_22077,N_16727,N_12805);
or U22078 (N_22078,N_17608,N_19236);
nor U22079 (N_22079,N_10074,N_14403);
xor U22080 (N_22080,N_15470,N_13959);
and U22081 (N_22081,N_15347,N_14353);
nand U22082 (N_22082,N_15109,N_13516);
or U22083 (N_22083,N_19782,N_15277);
nor U22084 (N_22084,N_13660,N_13295);
nand U22085 (N_22085,N_13496,N_15563);
xnor U22086 (N_22086,N_15095,N_10842);
nand U22087 (N_22087,N_11345,N_19570);
and U22088 (N_22088,N_11648,N_17495);
and U22089 (N_22089,N_10809,N_12250);
xor U22090 (N_22090,N_17999,N_11944);
or U22091 (N_22091,N_17189,N_13739);
xnor U22092 (N_22092,N_19664,N_16963);
nand U22093 (N_22093,N_12044,N_18727);
or U22094 (N_22094,N_10562,N_10646);
or U22095 (N_22095,N_10555,N_12747);
and U22096 (N_22096,N_15353,N_16920);
nor U22097 (N_22097,N_14109,N_11951);
or U22098 (N_22098,N_13398,N_13092);
nand U22099 (N_22099,N_16365,N_11608);
nand U22100 (N_22100,N_19957,N_16807);
xnor U22101 (N_22101,N_13738,N_17164);
and U22102 (N_22102,N_15930,N_12880);
and U22103 (N_22103,N_11307,N_18783);
nand U22104 (N_22104,N_11915,N_16705);
nand U22105 (N_22105,N_11382,N_13065);
and U22106 (N_22106,N_12454,N_14478);
nand U22107 (N_22107,N_19349,N_16993);
and U22108 (N_22108,N_18672,N_15237);
nor U22109 (N_22109,N_13204,N_14216);
nor U22110 (N_22110,N_11921,N_14238);
or U22111 (N_22111,N_18912,N_12788);
nor U22112 (N_22112,N_13694,N_14534);
xor U22113 (N_22113,N_19781,N_13141);
or U22114 (N_22114,N_10647,N_17420);
nor U22115 (N_22115,N_13060,N_15623);
nand U22116 (N_22116,N_14505,N_15816);
xnor U22117 (N_22117,N_18796,N_12818);
and U22118 (N_22118,N_17903,N_16030);
nor U22119 (N_22119,N_14626,N_16338);
xnor U22120 (N_22120,N_13047,N_11296);
and U22121 (N_22121,N_13399,N_18907);
or U22122 (N_22122,N_16045,N_13118);
xor U22123 (N_22123,N_16346,N_18910);
or U22124 (N_22124,N_12152,N_11949);
or U22125 (N_22125,N_14834,N_11085);
nor U22126 (N_22126,N_10857,N_12158);
nand U22127 (N_22127,N_18758,N_14573);
and U22128 (N_22128,N_10122,N_19065);
and U22129 (N_22129,N_19966,N_19272);
nand U22130 (N_22130,N_14543,N_13843);
xor U22131 (N_22131,N_17880,N_12492);
nor U22132 (N_22132,N_15890,N_13389);
and U22133 (N_22133,N_17763,N_12854);
nand U22134 (N_22134,N_12422,N_12361);
and U22135 (N_22135,N_15690,N_10129);
and U22136 (N_22136,N_13001,N_16533);
and U22137 (N_22137,N_15046,N_10996);
nand U22138 (N_22138,N_12001,N_11398);
nand U22139 (N_22139,N_12248,N_11774);
and U22140 (N_22140,N_11620,N_19425);
and U22141 (N_22141,N_10004,N_13947);
xnor U22142 (N_22142,N_10638,N_14184);
nand U22143 (N_22143,N_15495,N_18376);
nor U22144 (N_22144,N_11387,N_11815);
and U22145 (N_22145,N_15140,N_16329);
and U22146 (N_22146,N_16064,N_17312);
and U22147 (N_22147,N_14864,N_13085);
nor U22148 (N_22148,N_15460,N_19291);
or U22149 (N_22149,N_12226,N_17695);
xnor U22150 (N_22150,N_14023,N_13119);
and U22151 (N_22151,N_13355,N_19218);
nor U22152 (N_22152,N_18712,N_19954);
and U22153 (N_22153,N_10452,N_14272);
xnor U22154 (N_22154,N_14524,N_17886);
or U22155 (N_22155,N_16245,N_10254);
nand U22156 (N_22156,N_15366,N_14141);
xor U22157 (N_22157,N_15379,N_12059);
nor U22158 (N_22158,N_10013,N_11396);
nor U22159 (N_22159,N_18597,N_12039);
nand U22160 (N_22160,N_16062,N_16747);
and U22161 (N_22161,N_16832,N_14891);
xor U22162 (N_22162,N_17733,N_17700);
nor U22163 (N_22163,N_19273,N_12806);
xor U22164 (N_22164,N_12362,N_17127);
and U22165 (N_22165,N_15885,N_13824);
nand U22166 (N_22166,N_15912,N_16440);
and U22167 (N_22167,N_19707,N_13053);
xor U22168 (N_22168,N_16570,N_16845);
and U22169 (N_22169,N_19807,N_10582);
nand U22170 (N_22170,N_15336,N_15104);
xnor U22171 (N_22171,N_11993,N_18857);
xnor U22172 (N_22172,N_17272,N_19894);
nor U22173 (N_22173,N_16070,N_13755);
or U22174 (N_22174,N_17064,N_15559);
nor U22175 (N_22175,N_16516,N_13221);
and U22176 (N_22176,N_19813,N_17643);
nand U22177 (N_22177,N_16325,N_11200);
and U22178 (N_22178,N_15315,N_17557);
nand U22179 (N_22179,N_12171,N_10763);
and U22180 (N_22180,N_19339,N_16372);
xnor U22181 (N_22181,N_10506,N_15329);
nand U22182 (N_22182,N_14742,N_11214);
and U22183 (N_22183,N_11626,N_19459);
and U22184 (N_22184,N_13556,N_12279);
and U22185 (N_22185,N_11941,N_17438);
xnor U22186 (N_22186,N_12940,N_11099);
nand U22187 (N_22187,N_10427,N_15552);
nand U22188 (N_22188,N_17066,N_11113);
nand U22189 (N_22189,N_10391,N_16294);
and U22190 (N_22190,N_11076,N_16577);
or U22191 (N_22191,N_15067,N_10328);
nor U22192 (N_22192,N_12334,N_19053);
or U22193 (N_22193,N_13913,N_14860);
xnor U22194 (N_22194,N_16048,N_14180);
and U22195 (N_22195,N_13659,N_10905);
and U22196 (N_22196,N_19080,N_15789);
nor U22197 (N_22197,N_10930,N_11539);
nand U22198 (N_22198,N_12690,N_14267);
nand U22199 (N_22199,N_17362,N_11101);
or U22200 (N_22200,N_19038,N_11259);
nand U22201 (N_22201,N_17184,N_15451);
or U22202 (N_22202,N_11732,N_19797);
xor U22203 (N_22203,N_17281,N_15579);
nand U22204 (N_22204,N_17908,N_19101);
nand U22205 (N_22205,N_19375,N_19007);
or U22206 (N_22206,N_18899,N_15239);
nand U22207 (N_22207,N_19009,N_14103);
or U22208 (N_22208,N_17452,N_15641);
nand U22209 (N_22209,N_14879,N_11344);
and U22210 (N_22210,N_10250,N_13479);
and U22211 (N_22211,N_18518,N_18916);
nand U22212 (N_22212,N_10407,N_15393);
or U22213 (N_22213,N_13695,N_19035);
and U22214 (N_22214,N_15137,N_15323);
and U22215 (N_22215,N_15974,N_10413);
nand U22216 (N_22216,N_17300,N_16258);
xor U22217 (N_22217,N_11542,N_12444);
or U22218 (N_22218,N_15059,N_18718);
and U22219 (N_22219,N_13765,N_14855);
nand U22220 (N_22220,N_11533,N_10261);
or U22221 (N_22221,N_11760,N_11894);
xnor U22222 (N_22222,N_18163,N_13875);
xnor U22223 (N_22223,N_19207,N_15031);
and U22224 (N_22224,N_15320,N_11333);
or U22225 (N_22225,N_16800,N_14768);
or U22226 (N_22226,N_13690,N_12999);
and U22227 (N_22227,N_16075,N_14382);
xor U22228 (N_22228,N_15760,N_19195);
or U22229 (N_22229,N_16701,N_19243);
xor U22230 (N_22230,N_15319,N_19901);
nor U22231 (N_22231,N_11742,N_14031);
xnor U22232 (N_22232,N_11663,N_16960);
nand U22233 (N_22233,N_16741,N_12908);
xor U22234 (N_22234,N_13527,N_17814);
or U22235 (N_22235,N_12023,N_11618);
xnor U22236 (N_22236,N_13722,N_12120);
and U22237 (N_22237,N_18012,N_17366);
or U22238 (N_22238,N_12231,N_10153);
nand U22239 (N_22239,N_16349,N_12971);
and U22240 (N_22240,N_14092,N_19784);
nor U22241 (N_22241,N_19794,N_19678);
and U22242 (N_22242,N_19149,N_10124);
or U22243 (N_22243,N_15691,N_18933);
nand U22244 (N_22244,N_11546,N_18652);
and U22245 (N_22245,N_10482,N_17358);
nor U22246 (N_22246,N_13934,N_12313);
and U22247 (N_22247,N_12988,N_10692);
xnor U22248 (N_22248,N_19575,N_15340);
nand U22249 (N_22249,N_17043,N_18155);
nor U22250 (N_22250,N_18680,N_11707);
or U22251 (N_22251,N_14436,N_15630);
xnor U22252 (N_22252,N_11313,N_17895);
nand U22253 (N_22253,N_19117,N_15904);
or U22254 (N_22254,N_10432,N_13565);
nand U22255 (N_22255,N_14407,N_16520);
and U22256 (N_22256,N_11127,N_18502);
nor U22257 (N_22257,N_18533,N_14185);
xor U22258 (N_22258,N_19972,N_19352);
xor U22259 (N_22259,N_12393,N_12821);
and U22260 (N_22260,N_18171,N_16443);
and U22261 (N_22261,N_19757,N_10161);
nand U22262 (N_22262,N_12579,N_15208);
xor U22263 (N_22263,N_12438,N_16289);
nand U22264 (N_22264,N_14813,N_19055);
and U22265 (N_22265,N_19476,N_16278);
nor U22266 (N_22266,N_10237,N_15517);
and U22267 (N_22267,N_17843,N_13639);
nor U22268 (N_22268,N_11391,N_18863);
nand U22269 (N_22269,N_10192,N_13331);
and U22270 (N_22270,N_16514,N_18159);
nand U22271 (N_22271,N_12780,N_13508);
xor U22272 (N_22272,N_14422,N_17888);
xor U22273 (N_22273,N_17039,N_19860);
xor U22274 (N_22274,N_10485,N_14689);
nand U22275 (N_22275,N_16038,N_19315);
or U22276 (N_22276,N_16634,N_12102);
nor U22277 (N_22277,N_19606,N_16508);
xor U22278 (N_22278,N_11717,N_14328);
or U22279 (N_22279,N_11045,N_18070);
or U22280 (N_22280,N_15803,N_12914);
xor U22281 (N_22281,N_18746,N_15798);
nand U22282 (N_22282,N_17178,N_15489);
and U22283 (N_22283,N_19985,N_17658);
nand U22284 (N_22284,N_17143,N_11923);
and U22285 (N_22285,N_16357,N_17269);
and U22286 (N_22286,N_10029,N_16885);
nand U22287 (N_22287,N_16112,N_13177);
xnor U22288 (N_22288,N_15486,N_14466);
or U22289 (N_22289,N_13329,N_10299);
nor U22290 (N_22290,N_18288,N_13231);
and U22291 (N_22291,N_16757,N_11420);
nand U22292 (N_22292,N_13671,N_12568);
and U22293 (N_22293,N_18797,N_17425);
nand U22294 (N_22294,N_11326,N_19122);
and U22295 (N_22295,N_13422,N_13259);
nand U22296 (N_22296,N_17946,N_15622);
or U22297 (N_22297,N_17636,N_11972);
xor U22298 (N_22298,N_13546,N_17587);
xor U22299 (N_22299,N_15702,N_10441);
and U22300 (N_22300,N_16256,N_19298);
nor U22301 (N_22301,N_14360,N_16003);
and U22302 (N_22302,N_14423,N_11325);
or U22303 (N_22303,N_19868,N_11573);
and U22304 (N_22304,N_15156,N_18636);
nand U22305 (N_22305,N_15657,N_10690);
nor U22306 (N_22306,N_17485,N_11843);
xor U22307 (N_22307,N_17265,N_19418);
nor U22308 (N_22308,N_11614,N_18285);
nand U22309 (N_22309,N_12758,N_14392);
and U22310 (N_22310,N_12374,N_11583);
nand U22311 (N_22311,N_13768,N_18106);
nand U22312 (N_22312,N_13089,N_18114);
and U22313 (N_22313,N_16350,N_13305);
xnor U22314 (N_22314,N_15813,N_14386);
nor U22315 (N_22315,N_17045,N_17778);
xor U22316 (N_22316,N_14117,N_16816);
nand U22317 (N_22317,N_16782,N_15476);
or U22318 (N_22318,N_10915,N_10602);
nand U22319 (N_22319,N_12972,N_19310);
and U22320 (N_22320,N_11181,N_15570);
nor U22321 (N_22321,N_12680,N_19727);
nor U22322 (N_22322,N_10680,N_17129);
and U22323 (N_22323,N_18616,N_16466);
or U22324 (N_22324,N_16264,N_17053);
xor U22325 (N_22325,N_19015,N_12222);
nand U22326 (N_22326,N_12811,N_10063);
nor U22327 (N_22327,N_16939,N_15081);
nor U22328 (N_22328,N_18539,N_11384);
and U22329 (N_22329,N_17071,N_12318);
or U22330 (N_22330,N_17166,N_10087);
xor U22331 (N_22331,N_18695,N_11310);
or U22332 (N_22332,N_13698,N_17724);
nand U22333 (N_22333,N_18580,N_18698);
and U22334 (N_22334,N_11415,N_15248);
or U22335 (N_22335,N_13801,N_11612);
nor U22336 (N_22336,N_11805,N_10339);
and U22337 (N_22337,N_12926,N_16679);
and U22338 (N_22338,N_17854,N_16236);
or U22339 (N_22339,N_19820,N_16095);
nor U22340 (N_22340,N_10615,N_13418);
nand U22341 (N_22341,N_11459,N_10300);
and U22342 (N_22342,N_13136,N_12573);
xnor U22343 (N_22343,N_15821,N_16995);
or U22344 (N_22344,N_14457,N_14113);
xor U22345 (N_22345,N_10077,N_11315);
nor U22346 (N_22346,N_14590,N_17382);
and U22347 (N_22347,N_17031,N_18453);
or U22348 (N_22348,N_17722,N_15606);
or U22349 (N_22349,N_11001,N_14618);
or U22350 (N_22350,N_13644,N_11630);
xnor U22351 (N_22351,N_19411,N_13033);
nand U22352 (N_22352,N_18801,N_14663);
nor U22353 (N_22353,N_10569,N_14668);
xnor U22354 (N_22354,N_13574,N_14406);
nand U22355 (N_22355,N_10520,N_18220);
nor U22356 (N_22356,N_16060,N_17106);
nand U22357 (N_22357,N_12127,N_17450);
and U22358 (N_22358,N_10760,N_13024);
nand U22359 (N_22359,N_17750,N_19050);
or U22360 (N_22360,N_16881,N_14796);
nand U22361 (N_22361,N_17839,N_11316);
xnor U22362 (N_22362,N_17292,N_14973);
nand U22363 (N_22363,N_18699,N_13531);
or U22364 (N_22364,N_11350,N_16441);
and U22365 (N_22365,N_18060,N_11651);
xor U22366 (N_22366,N_11952,N_19293);
nand U22367 (N_22367,N_17982,N_17623);
xnor U22368 (N_22368,N_19158,N_19183);
nand U22369 (N_22369,N_13770,N_17828);
nand U22370 (N_22370,N_14264,N_15327);
or U22371 (N_22371,N_16838,N_16094);
nand U22372 (N_22372,N_15176,N_11668);
nor U22373 (N_22373,N_12862,N_12781);
or U22374 (N_22374,N_13549,N_19070);
xor U22375 (N_22375,N_11009,N_13529);
or U22376 (N_22376,N_10456,N_10900);
nand U22377 (N_22377,N_19405,N_11272);
nor U22378 (N_22378,N_19577,N_10815);
xnor U22379 (N_22379,N_14778,N_11636);
nand U22380 (N_22380,N_16435,N_18291);
nor U22381 (N_22381,N_11621,N_14069);
xor U22382 (N_22382,N_13759,N_18827);
nor U22383 (N_22383,N_14139,N_18874);
nor U22384 (N_22384,N_17773,N_10665);
or U22385 (N_22385,N_17310,N_14123);
and U22386 (N_22386,N_14806,N_16134);
and U22387 (N_22387,N_14585,N_15952);
xor U22388 (N_22388,N_16813,N_18849);
or U22389 (N_22389,N_14950,N_16322);
and U22390 (N_22390,N_15782,N_12410);
nand U22391 (N_22391,N_15311,N_14308);
and U22392 (N_22392,N_14818,N_11730);
and U22393 (N_22393,N_14144,N_19717);
and U22394 (N_22394,N_18965,N_19766);
or U22395 (N_22395,N_16829,N_11030);
xor U22396 (N_22396,N_13728,N_10060);
and U22397 (N_22397,N_13264,N_13726);
and U22398 (N_22398,N_14208,N_11670);
xor U22399 (N_22399,N_15646,N_13630);
nand U22400 (N_22400,N_17609,N_18022);
nor U22401 (N_22401,N_13598,N_10012);
and U22402 (N_22402,N_17900,N_15773);
xor U22403 (N_22403,N_10253,N_16649);
nand U22404 (N_22404,N_15865,N_15028);
xor U22405 (N_22405,N_11557,N_11606);
xnor U22406 (N_22406,N_11891,N_13964);
nand U22407 (N_22407,N_17802,N_10672);
and U22408 (N_22408,N_10472,N_13749);
or U22409 (N_22409,N_14863,N_15765);
nand U22410 (N_22410,N_10031,N_18062);
nor U22411 (N_22411,N_16148,N_19115);
and U22412 (N_22412,N_10099,N_11874);
nor U22413 (N_22413,N_10151,N_14959);
or U22414 (N_22414,N_18859,N_15088);
or U22415 (N_22415,N_14265,N_16361);
nand U22416 (N_22416,N_15001,N_15712);
xor U22417 (N_22417,N_17964,N_18609);
or U22418 (N_22418,N_12581,N_15721);
nor U22419 (N_22419,N_17663,N_19838);
nor U22420 (N_22420,N_16774,N_19384);
nor U22421 (N_22421,N_14175,N_19116);
nand U22422 (N_22422,N_17473,N_13101);
nand U22423 (N_22423,N_15356,N_16630);
or U22424 (N_22424,N_16008,N_17782);
xnor U22425 (N_22425,N_14732,N_19744);
or U22426 (N_22426,N_18294,N_10600);
xnor U22427 (N_22427,N_15577,N_17014);
or U22428 (N_22428,N_18107,N_11511);
and U22429 (N_22429,N_12283,N_18359);
and U22430 (N_22430,N_14632,N_18351);
xor U22431 (N_22431,N_19643,N_17543);
nor U22432 (N_22432,N_15662,N_16709);
nor U22433 (N_22433,N_12286,N_10475);
or U22434 (N_22434,N_19198,N_14628);
xor U22435 (N_22435,N_19142,N_16564);
nand U22436 (N_22436,N_10517,N_14911);
nand U22437 (N_22437,N_15943,N_14814);
or U22438 (N_22438,N_18945,N_13148);
nor U22439 (N_22439,N_14980,N_10364);
xor U22440 (N_22440,N_14816,N_12028);
or U22441 (N_22441,N_18180,N_10191);
nand U22442 (N_22442,N_10752,N_16865);
xor U22443 (N_22443,N_11578,N_17409);
and U22444 (N_22444,N_14499,N_12307);
xor U22445 (N_22445,N_17111,N_10898);
nand U22446 (N_22446,N_19415,N_15874);
nor U22447 (N_22447,N_16380,N_14898);
xor U22448 (N_22448,N_14836,N_11237);
and U22449 (N_22449,N_14261,N_10347);
nor U22450 (N_22450,N_19099,N_14186);
nand U22451 (N_22451,N_12631,N_10221);
and U22452 (N_22452,N_10799,N_18036);
xor U22453 (N_22453,N_18358,N_17024);
nand U22454 (N_22454,N_11679,N_14447);
xor U22455 (N_22455,N_15159,N_16903);
nand U22456 (N_22456,N_17416,N_12082);
and U22457 (N_22457,N_10363,N_12424);
and U22458 (N_22458,N_10424,N_11561);
xnor U22459 (N_22459,N_10335,N_13300);
nor U22460 (N_22460,N_18189,N_18043);
nand U22461 (N_22461,N_14621,N_14045);
or U22462 (N_22462,N_18457,N_12712);
or U22463 (N_22463,N_18477,N_11494);
or U22464 (N_22464,N_14785,N_11273);
nor U22465 (N_22465,N_13609,N_13137);
and U22466 (N_22466,N_12118,N_10385);
xor U22467 (N_22467,N_17644,N_19280);
nand U22468 (N_22468,N_13285,N_17319);
or U22469 (N_22469,N_13330,N_11044);
or U22470 (N_22470,N_17860,N_12561);
and U22471 (N_22471,N_14892,N_11141);
nand U22472 (N_22472,N_17116,N_14065);
nor U22473 (N_22473,N_16517,N_14993);
nand U22474 (N_22474,N_11171,N_15082);
and U22475 (N_22475,N_15300,N_12319);
nor U22476 (N_22476,N_14497,N_10030);
xnor U22477 (N_22477,N_18744,N_14287);
xor U22478 (N_22478,N_13732,N_19892);
nor U22479 (N_22479,N_15684,N_10501);
or U22480 (N_22480,N_17580,N_17651);
nand U22481 (N_22481,N_18721,N_19879);
nor U22482 (N_22482,N_10552,N_15260);
xnor U22483 (N_22483,N_16543,N_11363);
nand U22484 (N_22484,N_13535,N_14795);
nand U22485 (N_22485,N_13796,N_18072);
or U22486 (N_22486,N_18610,N_13425);
xor U22487 (N_22487,N_19584,N_11035);
or U22488 (N_22488,N_19110,N_16720);
or U22489 (N_22489,N_11980,N_17213);
nor U22490 (N_22490,N_18777,N_17410);
nand U22491 (N_22491,N_16488,N_10534);
and U22492 (N_22492,N_12459,N_12726);
xor U22493 (N_22493,N_14587,N_15624);
or U22494 (N_22494,N_14273,N_10401);
and U22495 (N_22495,N_18325,N_11021);
or U22496 (N_22496,N_15141,N_10497);
xnor U22497 (N_22497,N_14559,N_13509);
or U22498 (N_22498,N_18891,N_18447);
or U22499 (N_22499,N_11288,N_15993);
nand U22500 (N_22500,N_13936,N_13307);
or U22501 (N_22501,N_12330,N_15097);
and U22502 (N_22502,N_14233,N_10135);
nand U22503 (N_22503,N_16578,N_17994);
xor U22504 (N_22504,N_15424,N_12730);
nand U22505 (N_22505,N_16790,N_14280);
or U22506 (N_22506,N_17858,N_14227);
and U22507 (N_22507,N_19688,N_10451);
and U22508 (N_22508,N_19398,N_13492);
and U22509 (N_22509,N_15786,N_19681);
or U22510 (N_22510,N_18743,N_18855);
and U22511 (N_22511,N_12893,N_15432);
nor U22512 (N_22512,N_14916,N_18787);
nor U22513 (N_22513,N_15969,N_15674);
nor U22514 (N_22514,N_16042,N_12368);
and U22515 (N_22515,N_16464,N_12523);
xor U22516 (N_22516,N_10599,N_12375);
and U22517 (N_22517,N_18212,N_13882);
or U22518 (N_22518,N_17848,N_18173);
nand U22519 (N_22519,N_13029,N_18025);
or U22520 (N_22520,N_17577,N_10513);
nand U22521 (N_22521,N_18344,N_15675);
and U22522 (N_22522,N_12360,N_10059);
xor U22523 (N_22523,N_11228,N_13612);
xnor U22524 (N_22524,N_18545,N_17223);
xnor U22525 (N_22525,N_12912,N_18419);
xor U22526 (N_22526,N_11024,N_14129);
or U22527 (N_22527,N_13457,N_16067);
nor U22528 (N_22528,N_19918,N_13528);
or U22529 (N_22529,N_19494,N_15540);
xor U22530 (N_22530,N_16188,N_10532);
nand U22531 (N_22531,N_11808,N_11116);
nor U22532 (N_22532,N_10824,N_18218);
nor U22533 (N_22533,N_14154,N_18972);
or U22534 (N_22534,N_10985,N_12033);
nand U22535 (N_22535,N_15276,N_10845);
and U22536 (N_22536,N_16238,N_18365);
nand U22537 (N_22537,N_16296,N_10706);
nor U22538 (N_22538,N_15823,N_19225);
xor U22539 (N_22539,N_13133,N_15573);
and U22540 (N_22540,N_17602,N_10816);
nand U22541 (N_22541,N_18075,N_16052);
and U22542 (N_22542,N_15032,N_18257);
xnor U22543 (N_22543,N_18284,N_16704);
and U22544 (N_22544,N_10450,N_14502);
nand U22545 (N_22545,N_15520,N_16860);
and U22546 (N_22546,N_13015,N_16697);
xnor U22547 (N_22547,N_13124,N_14516);
xnor U22548 (N_22548,N_18208,N_19595);
or U22549 (N_22549,N_12007,N_19168);
xnor U22550 (N_22550,N_17885,N_15884);
nor U22551 (N_22551,N_11209,N_11924);
or U22552 (N_22552,N_16946,N_11948);
or U22553 (N_22553,N_17481,N_19119);
nand U22554 (N_22554,N_10412,N_16997);
nor U22555 (N_22555,N_11393,N_16416);
xor U22556 (N_22556,N_18663,N_10211);
xnor U22557 (N_22557,N_14991,N_16874);
and U22558 (N_22558,N_11716,N_11545);
nand U22559 (N_22559,N_17648,N_13052);
nor U22560 (N_22560,N_15169,N_10762);
nor U22561 (N_22561,N_11956,N_12605);
or U22562 (N_22562,N_16707,N_17533);
xor U22563 (N_22563,N_16114,N_15378);
nand U22564 (N_22564,N_12184,N_19365);
nor U22565 (N_22565,N_19531,N_15252);
xor U22566 (N_22566,N_19644,N_12110);
or U22567 (N_22567,N_14913,N_11192);
nor U22568 (N_22568,N_15245,N_10897);
xor U22569 (N_22569,N_10543,N_16479);
and U22570 (N_22570,N_19199,N_11260);
nand U22571 (N_22571,N_13417,N_18305);
and U22572 (N_22572,N_17921,N_13629);
nand U22573 (N_22573,N_10362,N_19649);
xor U22574 (N_22574,N_12471,N_13115);
nor U22575 (N_22575,N_16822,N_13458);
or U22576 (N_22576,N_18160,N_12848);
nand U22577 (N_22577,N_11705,N_17284);
xnor U22578 (N_22578,N_17161,N_18977);
or U22579 (N_22579,N_19475,N_16875);
and U22580 (N_22580,N_10916,N_18262);
and U22581 (N_22581,N_12344,N_11906);
nand U22582 (N_22582,N_18524,N_11423);
nor U22583 (N_22583,N_10797,N_13756);
or U22584 (N_22584,N_14767,N_10040);
xnor U22585 (N_22585,N_15105,N_17719);
nor U22586 (N_22586,N_11179,N_12455);
xor U22587 (N_22587,N_18361,N_10186);
xor U22588 (N_22588,N_17928,N_16585);
nor U22589 (N_22589,N_15921,N_15024);
nor U22590 (N_22590,N_10119,N_18791);
and U22591 (N_22591,N_16233,N_14451);
nand U22592 (N_22592,N_15920,N_11331);
nand U22593 (N_22593,N_13131,N_19841);
nand U22594 (N_22594,N_11476,N_18217);
and U22595 (N_22595,N_12868,N_14665);
nand U22596 (N_22596,N_18991,N_10396);
or U22597 (N_22597,N_17917,N_19232);
nand U22598 (N_22598,N_19751,N_18023);
nor U22599 (N_22599,N_19113,N_19760);
or U22600 (N_22600,N_15997,N_16420);
nor U22601 (N_22601,N_11289,N_13073);
nor U22602 (N_22602,N_16728,N_13567);
xor U22603 (N_22603,N_11527,N_17726);
or U22604 (N_22604,N_18999,N_13368);
and U22605 (N_22605,N_14986,N_18630);
nand U22606 (N_22606,N_10791,N_10737);
and U22607 (N_22607,N_15956,N_10003);
xnor U22608 (N_22608,N_11975,N_18967);
and U22609 (N_22609,N_12702,N_19615);
nand U22610 (N_22610,N_15186,N_10354);
xnor U22611 (N_22611,N_13180,N_16397);
xor U22612 (N_22612,N_14792,N_16579);
xnor U22613 (N_22613,N_12937,N_19692);
xor U22614 (N_22614,N_12411,N_11152);
nand U22615 (N_22615,N_19302,N_15427);
and U22616 (N_22616,N_12367,N_15578);
nor U22617 (N_22617,N_12473,N_16612);
and U22618 (N_22618,N_16240,N_15981);
and U22619 (N_22619,N_16762,N_11974);
or U22620 (N_22620,N_10438,N_18307);
and U22621 (N_22621,N_13245,N_11056);
xor U22622 (N_22622,N_16742,N_17313);
xor U22623 (N_22623,N_12720,N_13834);
xnor U22624 (N_22624,N_11785,N_13114);
nand U22625 (N_22625,N_17464,N_19131);
and U22626 (N_22626,N_15600,N_11720);
nor U22627 (N_22627,N_13746,N_13439);
and U22628 (N_22628,N_14320,N_18538);
nand U22629 (N_22629,N_11863,N_11633);
and U22630 (N_22630,N_10743,N_18154);
nand U22631 (N_22631,N_18380,N_16969);
and U22632 (N_22632,N_19925,N_17336);
nand U22633 (N_22633,N_10713,N_10287);
or U22634 (N_22634,N_10002,N_12851);
or U22635 (N_22635,N_13596,N_14627);
or U22636 (N_22636,N_18660,N_19680);
nor U22637 (N_22637,N_11829,N_17786);
and U22638 (N_22638,N_17353,N_17941);
xnor U22639 (N_22639,N_18481,N_18542);
xor U22640 (N_22640,N_15272,N_13076);
xnor U22641 (N_22641,N_11248,N_10911);
xnor U22642 (N_22642,N_16485,N_18817);
and U22643 (N_22643,N_12678,N_17463);
nor U22644 (N_22644,N_11125,N_14192);
or U22645 (N_22645,N_11443,N_12332);
nand U22646 (N_22646,N_11880,N_19716);
and U22647 (N_22647,N_14494,N_15664);
nand U22648 (N_22648,N_18437,N_10295);
nor U22649 (N_22649,N_12017,N_17413);
nand U22650 (N_22650,N_13165,N_15126);
xnor U22651 (N_22651,N_10979,N_18058);
or U22652 (N_22652,N_15561,N_11245);
nor U22653 (N_22653,N_17427,N_19409);
and U22654 (N_22654,N_12364,N_11531);
nand U22655 (N_22655,N_19872,N_15121);
nand U22656 (N_22656,N_10173,N_10961);
xnor U22657 (N_22657,N_19171,N_15422);
nand U22658 (N_22658,N_15344,N_12886);
nand U22659 (N_22659,N_17257,N_15234);
nor U22660 (N_22660,N_12874,N_11596);
nand U22661 (N_22661,N_18033,N_14409);
nor U22662 (N_22662,N_12242,N_12939);
and U22663 (N_22663,N_14193,N_16099);
xnor U22664 (N_22664,N_10521,N_17453);
nand U22665 (N_22665,N_15471,N_18685);
or U22666 (N_22666,N_11337,N_13760);
and U22667 (N_22667,N_11703,N_18420);
or U22668 (N_22668,N_13641,N_11794);
nor U22669 (N_22669,N_18013,N_14743);
nor U22670 (N_22670,N_18670,N_18244);
or U22671 (N_22671,N_19355,N_19346);
xor U22672 (N_22672,N_18256,N_14567);
xnor U22673 (N_22673,N_13831,N_16417);
or U22674 (N_22674,N_19368,N_16582);
nor U22675 (N_22675,N_15644,N_10194);
or U22676 (N_22676,N_14727,N_16667);
xor U22677 (N_22677,N_17320,N_17499);
nand U22678 (N_22678,N_11351,N_14107);
and U22679 (N_22679,N_12268,N_10567);
xor U22680 (N_22680,N_13872,N_16914);
or U22681 (N_22681,N_17666,N_17034);
or U22682 (N_22682,N_19746,N_19563);
nand U22683 (N_22683,N_10216,N_10946);
nand U22684 (N_22684,N_15221,N_11803);
nor U22685 (N_22685,N_10819,N_15538);
nor U22686 (N_22686,N_13714,N_18484);
and U22687 (N_22687,N_13213,N_11689);
or U22688 (N_22688,N_12292,N_11697);
and U22689 (N_22689,N_12302,N_10919);
xor U22690 (N_22690,N_10422,N_12592);
nand U22691 (N_22691,N_13862,N_16522);
nor U22692 (N_22692,N_16695,N_19854);
xnor U22693 (N_22693,N_19851,N_14867);
xnor U22694 (N_22694,N_10149,N_15249);
and U22695 (N_22695,N_19362,N_12249);
and U22696 (N_22696,N_11341,N_14687);
and U22697 (N_22697,N_19822,N_18350);
xnor U22698 (N_22698,N_10428,N_16424);
nor U22699 (N_22699,N_16110,N_10183);
or U22700 (N_22700,N_16542,N_13839);
nand U22701 (N_22701,N_12701,N_15879);
xor U22702 (N_22702,N_19573,N_13146);
and U22703 (N_22703,N_19565,N_14090);
or U22704 (N_22704,N_17770,N_12555);
nor U22705 (N_22705,N_11087,N_16994);
and U22706 (N_22706,N_17454,N_19247);
nand U22707 (N_22707,N_17743,N_17673);
nand U22708 (N_22708,N_14016,N_11429);
and U22709 (N_22709,N_14960,N_10292);
xnor U22710 (N_22710,N_16059,N_16748);
nor U22711 (N_22711,N_12273,N_19980);
nand U22712 (N_22712,N_12495,N_16381);
and U22713 (N_22713,N_15636,N_17415);
and U22714 (N_22714,N_10542,N_16607);
nand U22715 (N_22715,N_12840,N_19535);
nand U22716 (N_22716,N_14918,N_18754);
and U22717 (N_22717,N_14551,N_13919);
nand U22718 (N_22718,N_19834,N_16147);
nor U22719 (N_22719,N_12164,N_12844);
or U22720 (N_22720,N_10836,N_18418);
xnor U22721 (N_22721,N_17616,N_11417);
nor U22722 (N_22722,N_17137,N_17335);
nor U22723 (N_22723,N_15958,N_17503);
nor U22724 (N_22724,N_15546,N_17869);
nor U22725 (N_22725,N_13678,N_15617);
xnor U22726 (N_22726,N_15022,N_18804);
nand U22727 (N_22727,N_10942,N_12532);
xor U22728 (N_22728,N_17321,N_19516);
nand U22729 (N_22729,N_10723,N_13570);
or U22730 (N_22730,N_16796,N_13742);
and U22731 (N_22731,N_17932,N_16193);
xor U22732 (N_22732,N_10020,N_12134);
xor U22733 (N_22733,N_13990,N_19526);
or U22734 (N_22734,N_18061,N_13961);
nor U22735 (N_22735,N_18362,N_15564);
xor U22736 (N_22736,N_10467,N_16493);
and U22737 (N_22737,N_16502,N_14134);
xnor U22738 (N_22738,N_13821,N_11483);
nor U22739 (N_22739,N_14449,N_12048);
nand U22740 (N_22740,N_11153,N_12031);
nor U22741 (N_22741,N_14896,N_11162);
and U22742 (N_22742,N_15550,N_19107);
nor U22743 (N_22743,N_19347,N_14161);
or U22744 (N_22744,N_16414,N_19540);
nand U22745 (N_22745,N_17197,N_17199);
nand U22746 (N_22746,N_12228,N_14637);
nor U22747 (N_22747,N_10766,N_13160);
nor U22748 (N_22748,N_10510,N_18282);
or U22749 (N_22749,N_15792,N_14464);
and U22750 (N_22750,N_13081,N_17397);
nand U22751 (N_22751,N_14468,N_19403);
or U22752 (N_22752,N_18596,N_11724);
and U22753 (N_22753,N_14211,N_13193);
nand U22754 (N_22754,N_16551,N_14615);
nor U22755 (N_22755,N_18548,N_17032);
nand U22756 (N_22756,N_12403,N_13622);
nand U22757 (N_22757,N_18997,N_18528);
nor U22758 (N_22758,N_17916,N_13055);
and U22759 (N_22759,N_10398,N_13271);
or U22760 (N_22760,N_18462,N_15931);
and U22761 (N_22761,N_12266,N_14415);
or U22762 (N_22762,N_13949,N_18654);
and U22763 (N_22763,N_15531,N_17774);
nor U22764 (N_22764,N_11710,N_19221);
xnor U22765 (N_22765,N_18197,N_17471);
or U22766 (N_22766,N_19984,N_15751);
or U22767 (N_22767,N_15322,N_10731);
xor U22768 (N_22768,N_15409,N_15506);
xor U22769 (N_22769,N_19752,N_18497);
and U22770 (N_22770,N_17248,N_11493);
nand U22771 (N_22771,N_17877,N_18301);
nand U22772 (N_22772,N_12470,N_13424);
or U22773 (N_22773,N_18536,N_10155);
and U22774 (N_22774,N_17123,N_10558);
nor U22775 (N_22775,N_11627,N_10581);
xnor U22776 (N_22776,N_19287,N_19433);
nor U22777 (N_22777,N_18204,N_11682);
and U22778 (N_22778,N_18751,N_18657);
nand U22779 (N_22779,N_16140,N_12672);
nand U22780 (N_22780,N_15919,N_12501);
and U22781 (N_22781,N_12234,N_18932);
nor U22782 (N_22782,N_19445,N_12763);
nor U22783 (N_22783,N_17943,N_11734);
nand U22784 (N_22784,N_17268,N_15160);
or U22785 (N_22785,N_15388,N_16367);
nor U22786 (N_22786,N_11292,N_18309);
and U22787 (N_22787,N_18789,N_15758);
nand U22788 (N_22788,N_10414,N_13586);
nand U22789 (N_22789,N_18050,N_18020);
and U22790 (N_22790,N_19437,N_10920);
and U22791 (N_22791,N_17930,N_18078);
xor U22792 (N_22792,N_11381,N_14948);
nor U22793 (N_22793,N_16363,N_18206);
xor U22794 (N_22794,N_16580,N_15152);
nor U22795 (N_22795,N_11655,N_19762);
nand U22796 (N_22796,N_16156,N_13105);
nor U22797 (N_22797,N_18403,N_17333);
nand U22798 (N_22798,N_14921,N_16224);
or U22799 (N_22799,N_16200,N_12634);
nor U22800 (N_22800,N_12080,N_16664);
and U22801 (N_22801,N_18198,N_10195);
and U22802 (N_22802,N_11549,N_17507);
xor U22803 (N_22803,N_15700,N_19147);
nand U22804 (N_22804,N_17914,N_18549);
nor U22805 (N_22805,N_14872,N_19761);
xnor U22806 (N_22806,N_14623,N_17926);
and U22807 (N_22807,N_13989,N_16086);
and U22808 (N_22808,N_10736,N_19326);
or U22809 (N_22809,N_12141,N_17966);
nand U22810 (N_22810,N_11990,N_15255);
or U22811 (N_22811,N_10738,N_16486);
nand U22812 (N_22812,N_10140,N_15037);
or U22813 (N_22813,N_10653,N_12625);
and U22814 (N_22814,N_14448,N_15295);
nand U22815 (N_22815,N_15586,N_10370);
xnor U22816 (N_22816,N_11645,N_11092);
nand U22817 (N_22817,N_16310,N_18037);
or U22818 (N_22818,N_19062,N_11694);
and U22819 (N_22819,N_14954,N_11526);
and U22820 (N_22820,N_18424,N_19429);
or U22821 (N_22821,N_15231,N_10305);
nand U22822 (N_22822,N_19789,N_19428);
nor U22823 (N_22823,N_16736,N_14365);
nor U22824 (N_22824,N_15910,N_19675);
nor U22825 (N_22825,N_16037,N_11361);
nand U22826 (N_22826,N_12960,N_14979);
nand U22827 (N_22827,N_10889,N_12216);
nor U22828 (N_22828,N_10459,N_18192);
nor U22829 (N_22829,N_13658,N_10217);
or U22830 (N_22830,N_19856,N_19422);
nand U22831 (N_22831,N_19667,N_11446);
nand U22832 (N_22832,N_15701,N_15966);
nand U22833 (N_22833,N_13426,N_10934);
xor U22834 (N_22834,N_13943,N_19934);
nor U22835 (N_22835,N_15730,N_14771);
xnor U22836 (N_22836,N_13777,N_13455);
nand U22837 (N_22837,N_11567,N_14729);
xnor U22838 (N_22838,N_10315,N_11071);
nor U22839 (N_22839,N_10065,N_18729);
and U22840 (N_22840,N_12541,N_12594);
xnor U22841 (N_22841,N_10219,N_13526);
nand U22842 (N_22842,N_18300,N_13448);
xor U22843 (N_22843,N_10588,N_12391);
nor U22844 (N_22844,N_12771,N_18360);
or U22845 (N_22845,N_19129,N_14126);
nand U22846 (N_22846,N_11934,N_16556);
xnor U22847 (N_22847,N_13784,N_15455);
nor U22848 (N_22848,N_12841,N_14259);
nand U22849 (N_22849,N_15433,N_16446);
nor U22850 (N_22850,N_19380,N_18161);
xor U22851 (N_22851,N_18237,N_19654);
xnor U22852 (N_22852,N_15418,N_17400);
nor U22853 (N_22853,N_15558,N_18210);
xor U22854 (N_22854,N_13858,N_19523);
nor U22855 (N_22855,N_15029,N_18813);
and U22856 (N_22856,N_13692,N_17510);
and U22857 (N_22857,N_10181,N_16557);
or U22858 (N_22858,N_15780,N_11822);
and U22859 (N_22859,N_15562,N_16377);
xor U22860 (N_22860,N_11873,N_15979);
nor U22861 (N_22861,N_17680,N_14390);
nand U22862 (N_22862,N_13269,N_19277);
nand U22863 (N_22863,N_14076,N_16404);
xor U22864 (N_22864,N_15510,N_14786);
or U22865 (N_22865,N_14219,N_13985);
and U22866 (N_22866,N_11422,N_16399);
xnor U22867 (N_22867,N_12863,N_12211);
and U22868 (N_22868,N_10965,N_14652);
xnor U22869 (N_22869,N_13155,N_14737);
or U22870 (N_22870,N_11239,N_11293);
xnor U22871 (N_22871,N_15971,N_13652);
xor U22872 (N_22872,N_13802,N_13412);
nor U22873 (N_22873,N_15197,N_17714);
and U22874 (N_22874,N_15155,N_11186);
nand U22875 (N_22875,N_18768,N_10058);
and U22876 (N_22876,N_12058,N_13036);
and U22877 (N_22877,N_11890,N_11184);
and U22878 (N_22878,N_13480,N_15505);
nor U22879 (N_22879,N_12179,N_13915);
and U22880 (N_22880,N_18893,N_16973);
nor U22881 (N_22881,N_12138,N_15071);
or U22882 (N_22882,N_11265,N_13469);
nand U22883 (N_22883,N_17497,N_18394);
xor U22884 (N_22884,N_10651,N_17661);
nor U22885 (N_22885,N_11497,N_10212);
or U22886 (N_22886,N_14458,N_19196);
or U22887 (N_22887,N_13993,N_13278);
xor U22888 (N_22888,N_14840,N_16561);
nor U22889 (N_22889,N_12525,N_15783);
and U22890 (N_22890,N_19582,N_17716);
and U22891 (N_22891,N_10559,N_15608);
nand U22892 (N_22892,N_12220,N_16716);
nand U22893 (N_22893,N_16195,N_17302);
or U22894 (N_22894,N_19204,N_19943);
nor U22895 (N_22895,N_19864,N_14481);
or U22896 (N_22896,N_15523,N_10081);
or U22897 (N_22897,N_11367,N_19932);
nand U22898 (N_22898,N_13166,N_19913);
or U22899 (N_22899,N_15677,N_10886);
nand U22900 (N_22900,N_14851,N_15294);
nand U22901 (N_22901,N_16777,N_13957);
and U22902 (N_22902,N_10947,N_10536);
nor U22903 (N_22903,N_15464,N_16886);
or U22904 (N_22904,N_18819,N_13638);
nor U22905 (N_22905,N_10583,N_18314);
or U22906 (N_22906,N_11802,N_16930);
or U22907 (N_22907,N_13243,N_13677);
or U22908 (N_22908,N_13776,N_15944);
and U22909 (N_22909,N_17734,N_19095);
or U22910 (N_22910,N_10079,N_12807);
and U22911 (N_22911,N_15456,N_13800);
xor U22912 (N_22912,N_11595,N_10684);
xor U22913 (N_22913,N_17424,N_12578);
nor U22914 (N_22914,N_16328,N_15707);
nor U22915 (N_22915,N_13450,N_14927);
nor U22916 (N_22916,N_17435,N_11267);
and U22917 (N_22917,N_12564,N_12795);
nor U22918 (N_22918,N_15175,N_14519);
xnor U22919 (N_22919,N_16074,N_18906);
and U22920 (N_22920,N_18831,N_19695);
nand U22921 (N_22921,N_19611,N_15437);
and U22922 (N_22922,N_17984,N_16763);
and U22923 (N_22923,N_12793,N_12343);
or U22924 (N_22924,N_16978,N_11061);
nor U22925 (N_22925,N_11075,N_15830);
or U22926 (N_22926,N_16076,N_11961);
xor U22927 (N_22927,N_15204,N_12903);
nand U22928 (N_22928,N_19169,N_13176);
and U22929 (N_22929,N_14344,N_19732);
xor U22930 (N_22930,N_15411,N_18111);
nor U22931 (N_22931,N_18623,N_10880);
nor U22932 (N_22932,N_11193,N_12537);
or U22933 (N_22933,N_12614,N_12370);
nand U22934 (N_22934,N_16150,N_11327);
xnor U22935 (N_22935,N_18228,N_18522);
nand U22936 (N_22936,N_18955,N_16864);
or U22937 (N_22937,N_18088,N_12311);
and U22938 (N_22938,N_14846,N_12761);
and U22939 (N_22939,N_17572,N_14177);
nand U22940 (N_22940,N_18326,N_11458);
xor U22941 (N_22941,N_13436,N_11468);
or U22942 (N_22942,N_13250,N_10045);
or U22943 (N_22943,N_18658,N_11942);
and U22944 (N_22944,N_10933,N_19958);
and U22945 (N_22945,N_13129,N_11669);
and U22946 (N_22946,N_14333,N_15583);
nor U22947 (N_22947,N_10603,N_14120);
and U22948 (N_22948,N_14437,N_16588);
nand U22949 (N_22949,N_16047,N_19579);
nand U22950 (N_22950,N_10156,N_16287);
nor U22951 (N_22951,N_10932,N_16611);
nor U22952 (N_22952,N_16297,N_18480);
nand U22953 (N_22953,N_15241,N_10590);
nand U22954 (N_22954,N_15124,N_19442);
and U22955 (N_22955,N_17968,N_18701);
xnor U22956 (N_22956,N_14849,N_17906);
and U22957 (N_22957,N_16689,N_10574);
nor U22958 (N_22958,N_19301,N_18135);
and U22959 (N_22959,N_12812,N_11490);
xnor U22960 (N_22960,N_10196,N_13932);
nand U22961 (N_22961,N_15647,N_14717);
nand U22962 (N_22962,N_11308,N_12143);
nand U22963 (N_22963,N_10624,N_19078);
nor U22964 (N_22964,N_15869,N_17694);
nand U22965 (N_22965,N_16722,N_13327);
xor U22966 (N_22966,N_19270,N_12657);
and U22967 (N_22967,N_12392,N_13315);
or U22968 (N_22968,N_16636,N_15195);
and U22969 (N_22969,N_15004,N_10477);
nand U22970 (N_22970,N_11322,N_15699);
and U22971 (N_22971,N_19541,N_18145);
or U22972 (N_22972,N_16009,N_15302);
and U22973 (N_22973,N_19898,N_10994);
xnor U22974 (N_22974,N_19343,N_11943);
xnor U22975 (N_22975,N_13946,N_12703);
or U22976 (N_22976,N_11098,N_14542);
and U22977 (N_22977,N_13584,N_13378);
xnor U22978 (N_22978,N_14317,N_15887);
nand U22979 (N_22979,N_15171,N_16625);
and U22980 (N_22980,N_18684,N_18076);
xnor U22981 (N_22981,N_18550,N_11115);
and U22982 (N_22982,N_13813,N_11708);
and U22983 (N_22983,N_18261,N_16823);
nand U22984 (N_22984,N_15099,N_16309);
or U22985 (N_22985,N_14188,N_17156);
and U22986 (N_22986,N_16243,N_15722);
xor U22987 (N_22987,N_10091,N_13318);
or U22988 (N_22988,N_14661,N_11304);
nand U22989 (N_22989,N_11371,N_18830);
xor U22990 (N_22990,N_13293,N_18834);
and U22991 (N_22991,N_16526,N_17150);
nor U22992 (N_22992,N_17911,N_13737);
xor U22993 (N_22993,N_14812,N_16395);
xnor U22994 (N_22994,N_14411,N_16410);
nor U22995 (N_22995,N_11848,N_17957);
xnor U22996 (N_22996,N_13282,N_19648);
nor U22997 (N_22997,N_18035,N_15643);
xnor U22998 (N_22998,N_10568,N_14683);
and U22999 (N_22999,N_10969,N_12662);
and U23000 (N_23000,N_13688,N_13288);
or U23001 (N_23001,N_10891,N_17929);
and U23002 (N_23002,N_10868,N_14106);
nand U23003 (N_23003,N_14719,N_12600);
nor U23004 (N_23004,N_12209,N_17904);
xnor U23005 (N_23005,N_16892,N_12460);
xnor U23006 (N_23006,N_11871,N_16912);
or U23007 (N_23007,N_18575,N_15724);
xnor U23008 (N_23008,N_16174,N_12878);
or U23009 (N_23009,N_19917,N_12498);
and U23010 (N_23010,N_15283,N_14331);
or U23011 (N_23011,N_13780,N_17548);
or U23012 (N_23012,N_19825,N_10056);
xnor U23013 (N_23013,N_19924,N_15205);
xnor U23014 (N_23014,N_15990,N_13938);
nand U23015 (N_23015,N_12787,N_14002);
or U23016 (N_23016,N_15584,N_10378);
and U23017 (N_23017,N_11416,N_14508);
and U23018 (N_23018,N_12705,N_12717);
nor U23019 (N_23019,N_10068,N_11522);
nor U23020 (N_23020,N_12922,N_15444);
or U23021 (N_23021,N_14939,N_19995);
xor U23022 (N_23022,N_11599,N_16512);
or U23023 (N_23023,N_13689,N_18194);
nor U23024 (N_23024,N_12142,N_18048);
xnor U23025 (N_23025,N_10484,N_15167);
nand U23026 (N_23026,N_10547,N_18631);
nand U23027 (N_23027,N_13135,N_19527);
or U23028 (N_23028,N_12817,N_13020);
xor U23029 (N_23029,N_18461,N_11850);
nand U23030 (N_23030,N_16944,N_17987);
nor U23031 (N_23031,N_15923,N_16321);
and U23032 (N_23032,N_18742,N_16393);
xor U23033 (N_23033,N_13403,N_14606);
or U23034 (N_23034,N_10570,N_14907);
nor U23035 (N_23035,N_14292,N_14766);
and U23036 (N_23036,N_12276,N_10783);
and U23037 (N_23037,N_13423,N_13904);
or U23038 (N_23038,N_11660,N_17430);
and U23039 (N_23039,N_16127,N_14788);
and U23040 (N_23040,N_19305,N_16187);
xor U23041 (N_23041,N_15226,N_17913);
nor U23042 (N_23042,N_12247,N_18740);
nand U23043 (N_23043,N_16452,N_12386);
nor U23044 (N_23044,N_17607,N_19750);
and U23045 (N_23045,N_12230,N_17013);
and U23046 (N_23046,N_17870,N_15868);
and U23047 (N_23047,N_11881,N_18644);
and U23048 (N_23048,N_18207,N_12725);
and U23049 (N_23049,N_10742,N_12842);
and U23050 (N_23050,N_18865,N_15482);
and U23051 (N_23051,N_19057,N_18532);
nor U23052 (N_23052,N_13127,N_15513);
xor U23053 (N_23053,N_12203,N_19317);
nor U23054 (N_23054,N_14631,N_12740);
or U23055 (N_23055,N_18615,N_18531);
and U23056 (N_23056,N_17040,N_13296);
nor U23057 (N_23057,N_17810,N_10025);
and U23058 (N_23058,N_10226,N_14197);
nor U23059 (N_23059,N_15534,N_17242);
xnor U23060 (N_23060,N_10589,N_13906);
nor U23061 (N_23061,N_18992,N_17216);
xor U23062 (N_23062,N_18811,N_16887);
nor U23063 (N_23063,N_17674,N_14334);
or U23064 (N_23064,N_17017,N_19694);
or U23065 (N_23065,N_16386,N_17511);
nor U23066 (N_23066,N_11922,N_17660);
xnor U23067 (N_23067,N_15142,N_13560);
nor U23068 (N_23068,N_17509,N_12435);
nor U23069 (N_23069,N_19815,N_15123);
xor U23070 (N_23070,N_12398,N_17690);
or U23071 (N_23071,N_13797,N_17945);
or U23072 (N_23072,N_17270,N_12980);
nor U23073 (N_23073,N_11303,N_18773);
xor U23074 (N_23074,N_10409,N_15225);
xnor U23075 (N_23075,N_17211,N_17190);
nor U23076 (N_23076,N_17939,N_19340);
nand U23077 (N_23077,N_15806,N_18349);
nor U23078 (N_23078,N_19650,N_14307);
or U23079 (N_23079,N_12457,N_17508);
and U23080 (N_23080,N_17989,N_18008);
and U23081 (N_23081,N_16490,N_10343);
xnor U23082 (N_23082,N_11020,N_19331);
and U23083 (N_23083,N_13167,N_12876);
and U23084 (N_23084,N_17937,N_11194);
nand U23085 (N_23085,N_15772,N_14612);
and U23086 (N_23086,N_16546,N_14213);
and U23087 (N_23087,N_15368,N_15130);
and U23088 (N_23088,N_19264,N_16209);
or U23089 (N_23089,N_19000,N_19862);
or U23090 (N_23090,N_16638,N_14051);
or U23091 (N_23091,N_18491,N_14098);
xor U23092 (N_23092,N_12282,N_14885);
nand U23093 (N_23093,N_19125,N_12935);
or U23094 (N_23094,N_10789,N_19759);
nand U23095 (N_23095,N_14318,N_17407);
nor U23096 (N_23096,N_17569,N_12073);
or U23097 (N_23097,N_14779,N_15314);
nor U23098 (N_23098,N_16032,N_13144);
nor U23099 (N_23099,N_10233,N_11250);
and U23100 (N_23100,N_10493,N_12380);
nand U23101 (N_23101,N_18697,N_15017);
nor U23102 (N_23102,N_18375,N_13258);
nand U23103 (N_23103,N_12196,N_14472);
nand U23104 (N_23104,N_12275,N_14938);
and U23105 (N_23105,N_18329,N_16218);
nor U23106 (N_23106,N_19160,N_11918);
or U23107 (N_23107,N_12824,N_12965);
or U23108 (N_23108,N_12433,N_12452);
nor U23109 (N_23109,N_14617,N_18465);
nor U23110 (N_23110,N_15014,N_11982);
nand U23111 (N_23111,N_17631,N_18903);
nand U23112 (N_23112,N_18275,N_13397);
xnor U23113 (N_23113,N_13578,N_13452);
nor U23114 (N_23114,N_18557,N_19740);
nand U23115 (N_23115,N_17388,N_18181);
nor U23116 (N_23116,N_14773,N_19756);
nor U23117 (N_23117,N_11535,N_15117);
xnor U23118 (N_23118,N_18705,N_13758);
or U23119 (N_23119,N_13899,N_16382);
and U23120 (N_23120,N_11283,N_16802);
nor U23121 (N_23121,N_11712,N_17959);
and U23122 (N_23122,N_10660,N_14148);
nand U23123 (N_23123,N_19745,N_15817);
xor U23124 (N_23124,N_11454,N_10024);
or U23125 (N_23125,N_10776,N_15536);
or U23126 (N_23126,N_14027,N_13324);
nor U23127 (N_23127,N_13445,N_11778);
nor U23128 (N_23128,N_16249,N_18710);
and U23129 (N_23129,N_18521,N_12394);
or U23130 (N_23130,N_13279,N_17456);
or U23131 (N_23131,N_19840,N_10707);
xor U23132 (N_23132,N_11728,N_19817);
nand U23133 (N_23133,N_15380,N_16991);
nand U23134 (N_23134,N_16071,N_15265);
nand U23135 (N_23135,N_17691,N_19051);
and U23136 (N_23136,N_18583,N_10230);
and U23137 (N_23137,N_13750,N_12310);
xor U23138 (N_23138,N_17983,N_14705);
or U23139 (N_23139,N_11065,N_19986);
or U23140 (N_23140,N_13924,N_18451);
or U23141 (N_23141,N_12695,N_10086);
and U23142 (N_23142,N_12015,N_16811);
nor U23143 (N_23143,N_13019,N_10337);
nor U23144 (N_23144,N_16053,N_10375);
and U23145 (N_23145,N_18221,N_19075);
and U23146 (N_23146,N_19471,N_11814);
nand U23147 (N_23147,N_12423,N_13525);
nand U23148 (N_23148,N_12369,N_13583);
nor U23149 (N_23149,N_11438,N_19488);
xnor U23150 (N_23150,N_13338,N_10750);
xor U23151 (N_23151,N_12450,N_13740);
nor U23152 (N_23152,N_14600,N_17350);
and U23153 (N_23153,N_15212,N_18651);
nand U23154 (N_23154,N_15620,N_12032);
or U23155 (N_23155,N_14878,N_13361);
xor U23156 (N_23156,N_16430,N_11727);
or U23157 (N_23157,N_14622,N_12877);
nor U23158 (N_23158,N_11574,N_13037);
and U23159 (N_23159,N_11414,N_18001);
and U23160 (N_23160,N_10046,N_16916);
xor U23161 (N_23161,N_17241,N_10325);
or U23162 (N_23162,N_16998,N_10910);
nor U23163 (N_23163,N_13650,N_12365);
xor U23164 (N_23164,N_19001,N_12598);
xnor U23165 (N_23165,N_18459,N_13202);
xor U23166 (N_23166,N_11649,N_15631);
and U23167 (N_23167,N_14441,N_10921);
nand U23168 (N_23168,N_17504,N_15440);
nand U23169 (N_23169,N_13086,N_18265);
nor U23170 (N_23170,N_16318,N_19936);
nor U23171 (N_23171,N_13440,N_14326);
nand U23172 (N_23172,N_13788,N_14722);
nand U23173 (N_23173,N_11442,N_14515);
and U23174 (N_23174,N_18678,N_15922);
nor U23175 (N_23175,N_14566,N_19172);
nor U23176 (N_23176,N_14270,N_19387);
nor U23177 (N_23177,N_12516,N_16347);
and U23178 (N_23178,N_17995,N_10455);
nand U23179 (N_23179,N_10344,N_14194);
nor U23180 (N_23180,N_12630,N_18499);
xor U23181 (N_23181,N_17938,N_18400);
xnor U23182 (N_23182,N_11865,N_11579);
nor U23183 (N_23183,N_19987,N_11875);
and U23184 (N_23184,N_12215,N_16795);
or U23185 (N_23185,N_10907,N_13206);
nor U23186 (N_23186,N_11366,N_15172);
or U23187 (N_23187,N_10126,N_13241);
nor U23188 (N_23188,N_11739,N_11744);
nor U23189 (N_23189,N_15045,N_15744);
nand U23190 (N_23190,N_12956,N_14919);
xnor U23191 (N_23191,N_13602,N_19604);
nand U23192 (N_23192,N_10548,N_19974);
or U23193 (N_23193,N_18734,N_15449);
and U23194 (N_23194,N_10115,N_10376);
xor U23195 (N_23195,N_10108,N_19482);
nor U23196 (N_23196,N_11300,N_16016);
xnor U23197 (N_23197,N_18952,N_12667);
nor U23198 (N_23198,N_14555,N_19098);
nand U23199 (N_23199,N_19460,N_13600);
nand U23200 (N_23200,N_10284,N_16211);
and U23201 (N_23201,N_13237,N_11036);
xnor U23202 (N_23202,N_12633,N_15860);
or U23203 (N_23203,N_15274,N_15280);
nor U23204 (N_23204,N_18890,N_17324);
nand U23205 (N_23205,N_18219,N_17979);
nand U23206 (N_23206,N_10349,N_13344);
and U23207 (N_23207,N_18836,N_17849);
nand U23208 (N_23208,N_12647,N_10541);
and U23209 (N_23209,N_11256,N_15338);
or U23210 (N_23210,N_10302,N_17646);
nand U23211 (N_23211,N_17781,N_18969);
nand U23212 (N_23212,N_18671,N_11460);
and U23213 (N_23213,N_18704,N_19224);
nand U23214 (N_23214,N_11275,N_17022);
nor U23215 (N_23215,N_15632,N_19162);
or U23216 (N_23216,N_18079,N_16040);
nor U23217 (N_23217,N_13191,N_15287);
nand U23218 (N_23218,N_13208,N_14883);
and U23219 (N_23219,N_15825,N_19855);
and U23220 (N_23220,N_13910,N_18719);
xor U23221 (N_23221,N_17922,N_12707);
xor U23222 (N_23222,N_15667,N_10512);
and U23223 (N_23223,N_14214,N_12737);
xor U23224 (N_23224,N_13587,N_14235);
nand U23225 (N_23225,N_10318,N_19140);
nor U23226 (N_23226,N_10324,N_19574);
and U23227 (N_23227,N_10404,N_16911);
or U23228 (N_23228,N_17593,N_12623);
nand U23229 (N_23229,N_13179,N_18054);
nand U23230 (N_23230,N_18016,N_19905);
and U23231 (N_23231,N_11876,N_14754);
or U23232 (N_23232,N_17701,N_12295);
and U23233 (N_23233,N_17635,N_15417);
nand U23234 (N_23234,N_18306,N_16610);
nor U23235 (N_23235,N_12924,N_15660);
xnor U23236 (N_23236,N_11576,N_18374);
or U23237 (N_23237,N_14005,N_13370);
nor U23238 (N_23238,N_13303,N_17107);
and U23239 (N_23239,N_15739,N_10877);
and U23240 (N_23240,N_18357,N_10681);
xnor U23241 (N_23241,N_17518,N_10248);
nor U23242 (N_23242,N_11959,N_12414);
nor U23243 (N_23243,N_16136,N_11554);
or U23244 (N_23244,N_16718,N_13354);
xor U23245 (N_23245,N_11514,N_19491);
or U23246 (N_23246,N_16809,N_18225);
nand U23247 (N_23247,N_12169,N_13499);
or U23248 (N_23248,N_10270,N_19660);
or U23249 (N_23249,N_13861,N_12181);
xor U23250 (N_23250,N_12792,N_17728);
xor U23251 (N_23251,N_17872,N_12060);
xor U23252 (N_23252,N_13835,N_14841);
nand U23253 (N_23253,N_14630,N_10671);
or U23254 (N_23254,N_15261,N_19959);
and U23255 (N_23255,N_12003,N_17192);
xor U23256 (N_23256,N_17075,N_16315);
nor U23257 (N_23257,N_16964,N_14028);
nand U23258 (N_23258,N_15382,N_17049);
nor U23259 (N_23259,N_18266,N_16251);
xnor U23260 (N_23260,N_17650,N_17985);
nor U23261 (N_23261,N_14750,N_14081);
and U23262 (N_23262,N_14882,N_13066);
nand U23263 (N_23263,N_13716,N_15369);
nor U23264 (N_23264,N_12961,N_19989);
nor U23265 (N_23265,N_18605,N_12437);
nor U23266 (N_23266,N_13211,N_10350);
or U23267 (N_23267,N_11859,N_17101);
or U23268 (N_23268,N_19238,N_19190);
and U23269 (N_23269,N_18295,N_12519);
nor U23270 (N_23270,N_10038,N_14271);
nand U23271 (N_23271,N_11905,N_15292);
nand U23272 (N_23272,N_19167,N_10598);
nor U23273 (N_23273,N_11570,N_12172);
nand U23274 (N_23274,N_16354,N_17383);
or U23275 (N_23275,N_19286,N_16622);
xnor U23276 (N_23276,N_14654,N_14203);
or U23277 (N_23277,N_16876,N_14080);
nor U23278 (N_23278,N_19054,N_13084);
xnor U23279 (N_23279,N_18254,N_17451);
or U23280 (N_23280,N_16167,N_19931);
and U23281 (N_23281,N_11392,N_17671);
xor U23282 (N_23282,N_15232,N_13561);
xnor U23283 (N_23283,N_14173,N_16028);
or U23284 (N_23284,N_19440,N_15652);
nand U23285 (N_23285,N_13545,N_12599);
nor U23286 (N_23286,N_13853,N_19747);
or U23287 (N_23287,N_13254,N_17287);
or U23288 (N_23288,N_13244,N_18454);
nand U23289 (N_23289,N_15410,N_14396);
and U23290 (N_23290,N_13779,N_11768);
nand U23291 (N_23291,N_18002,N_12113);
or U23292 (N_23292,N_11073,N_16686);
xnor U23293 (N_23293,N_11349,N_11354);
nor U23294 (N_23294,N_17224,N_13988);
nor U23295 (N_23295,N_15519,N_13209);
nor U23296 (N_23296,N_19028,N_11406);
xnor U23297 (N_23297,N_10939,N_12602);
and U23298 (N_23298,N_19930,N_12638);
nor U23299 (N_23299,N_14014,N_12094);
nand U23300 (N_23300,N_14068,N_19941);
or U23301 (N_23301,N_12552,N_13734);
and U23302 (N_23302,N_17115,N_14017);
xor U23303 (N_23303,N_19420,N_10064);
or U23304 (N_23304,N_17283,N_10812);
nand U23305 (N_23305,N_16482,N_17112);
xor U23306 (N_23306,N_18283,N_19438);
xnor U23307 (N_23307,N_17258,N_12785);
xnor U23308 (N_23308,N_18717,N_10663);
and U23309 (N_23309,N_19188,N_10779);
nor U23310 (N_23310,N_13017,N_12325);
nor U23311 (N_23311,N_16646,N_17121);
nand U23312 (N_23312,N_14616,N_17030);
nand U23313 (N_23313,N_12356,N_12928);
xnor U23314 (N_23314,N_18553,N_19210);
xnor U23315 (N_23315,N_10103,N_16155);
xor U23316 (N_23316,N_14805,N_15038);
nor U23317 (N_23317,N_16683,N_11418);
nor U23318 (N_23318,N_18317,N_13484);
nor U23319 (N_23319,N_14999,N_16852);
nand U23320 (N_23320,N_17393,N_16519);
and U23321 (N_23321,N_14171,N_12254);
or U23322 (N_23322,N_16798,N_16702);
and U23323 (N_23323,N_19356,N_16248);
xnor U23324 (N_23324,N_17220,N_18530);
xnor U23325 (N_23325,N_18124,N_10048);
or U23326 (N_23326,N_14222,N_18042);
xnor U23327 (N_23327,N_13088,N_18142);
and U23328 (N_23328,N_11129,N_17091);
and U23329 (N_23329,N_12896,N_15364);
nand U23330 (N_23330,N_13523,N_15100);
and U23331 (N_23331,N_10274,N_18515);
or U23332 (N_23332,N_18149,N_16713);
and U23333 (N_23333,N_18723,N_11017);
nor U23334 (N_23334,N_18458,N_15069);
or U23335 (N_23335,N_12093,N_17706);
or U23336 (N_23336,N_11550,N_14125);
nor U23337 (N_23337,N_15793,N_14136);
nand U23338 (N_23338,N_14696,N_19353);
nor U23339 (N_23339,N_11672,N_10561);
or U23340 (N_23340,N_11495,N_14251);
nand U23341 (N_23341,N_11463,N_19137);
and U23342 (N_23342,N_19043,N_10553);
or U23343 (N_23343,N_18203,N_14691);
or U23344 (N_23344,N_14889,N_13553);
nand U23345 (N_23345,N_14474,N_16204);
nand U23346 (N_23346,N_10224,N_16476);
nor U23347 (N_23347,N_19189,N_10826);
and U23348 (N_23348,N_19689,N_13485);
xor U23349 (N_23349,N_16202,N_13263);
and U23350 (N_23350,N_13674,N_12888);
nand U23351 (N_23351,N_10225,N_12265);
and U23352 (N_23352,N_18234,N_16341);
nor U23353 (N_23353,N_13844,N_11505);
nand U23354 (N_23354,N_14383,N_18683);
and U23355 (N_23355,N_16873,N_12175);
nand U23356 (N_23356,N_15285,N_14803);
or U23357 (N_23357,N_19215,N_11502);
xor U23358 (N_23358,N_16812,N_12287);
or U23359 (N_23359,N_12869,N_10835);
xor U23360 (N_23360,N_16453,N_13227);
or U23361 (N_23361,N_11926,N_13222);
nand U23362 (N_23362,N_14327,N_17702);
and U23363 (N_23363,N_10711,N_17482);
nor U23364 (N_23364,N_12651,N_13903);
nand U23365 (N_23365,N_14418,N_17565);
nor U23366 (N_23366,N_16613,N_18620);
nand U23367 (N_23367,N_19489,N_17339);
and U23368 (N_23368,N_15030,N_14229);
or U23369 (N_23369,N_13572,N_19674);
and U23370 (N_23370,N_19585,N_11150);
nor U23371 (N_23371,N_11541,N_11224);
xnor U23372 (N_23372,N_12144,N_17523);
nor U23373 (N_23373,N_18517,N_14049);
xnor U23374 (N_23374,N_12517,N_15332);
nor U23375 (N_23375,N_10346,N_18725);
xor U23376 (N_23376,N_12621,N_12637);
or U23377 (N_23377,N_11804,N_11609);
and U23378 (N_23378,N_11064,N_14225);
nand U23379 (N_23379,N_17301,N_10232);
and U23380 (N_23380,N_17217,N_12496);
nand U23381 (N_23381,N_15727,N_15877);
nor U23382 (N_23382,N_15864,N_14323);
nand U23383 (N_23383,N_17944,N_17844);
and U23384 (N_23384,N_18417,N_16999);
or U23385 (N_23385,N_14692,N_15023);
nand U23386 (N_23386,N_10678,N_11825);
or U23387 (N_23387,N_19915,N_17785);
or U23388 (N_23388,N_14694,N_11247);
nor U23389 (N_23389,N_13446,N_15403);
and U23390 (N_23390,N_16181,N_12813);
xor U23391 (N_23391,N_19944,N_14166);
nand U23392 (N_23392,N_13460,N_18561);
and U23393 (N_23393,N_14131,N_12819);
and U23394 (N_23394,N_12900,N_14777);
nor U23395 (N_23395,N_12704,N_16959);
nor U23396 (N_23396,N_15616,N_11074);
xnor U23397 (N_23397,N_16883,N_11298);
and U23398 (N_23398,N_16659,N_11516);
and U23399 (N_23399,N_17820,N_19049);
nand U23400 (N_23400,N_14429,N_14725);
or U23401 (N_23401,N_19795,N_16122);
xnor U23402 (N_23402,N_11586,N_15383);
and U23403 (N_23403,N_14479,N_19245);
nor U23404 (N_23404,N_11823,N_12068);
nand U23405 (N_23405,N_13068,N_12018);
nor U23406 (N_23406,N_16918,N_19161);
xnor U23407 (N_23407,N_13248,N_14446);
or U23408 (N_23408,N_10565,N_18172);
nand U23409 (N_23409,N_11706,N_10850);
or U23410 (N_23410,N_15115,N_15670);
and U23411 (N_23411,N_14063,N_12968);
and U23412 (N_23412,N_16406,N_18421);
xnor U23413 (N_23413,N_18456,N_14577);
and U23414 (N_23414,N_17462,N_10703);
or U23415 (N_23415,N_17067,N_12419);
xnor U23416 (N_23416,N_15222,N_19539);
and U23417 (N_23417,N_10112,N_14142);
or U23418 (N_23418,N_11940,N_11733);
nand U23419 (N_23419,N_14046,N_10833);
nor U23420 (N_23420,N_17195,N_12833);
and U23421 (N_23421,N_10440,N_13373);
nand U23422 (N_23422,N_16513,N_12889);
nor U23423 (N_23423,N_13859,N_18379);
and U23424 (N_23424,N_13571,N_11199);
xnor U23425 (N_23425,N_12870,N_11662);
and U23426 (N_23426,N_11667,N_14944);
and U23427 (N_23427,N_17652,N_11631);
and U23428 (N_23428,N_19275,N_15715);
xnor U23429 (N_23429,N_19205,N_11945);
nor U23430 (N_23430,N_17803,N_18713);
nand U23431 (N_23431,N_17780,N_18068);
and U23432 (N_23432,N_18441,N_19338);
xnor U23433 (N_23433,N_13323,N_13864);
or U23434 (N_23434,N_11063,N_15678);
nor U23435 (N_23435,N_12269,N_17373);
nor U23436 (N_23436,N_10956,N_16065);
nand U23437 (N_23437,N_15342,N_18726);
or U23438 (N_23438,N_11286,N_12225);
nor U23439 (N_23439,N_19431,N_10419);
or U23440 (N_23440,N_13194,N_12986);
nand U23441 (N_23441,N_19251,N_14302);
nand U23442 (N_23442,N_18131,N_12533);
nor U23443 (N_23443,N_12693,N_14401);
and U23444 (N_23444,N_11147,N_17015);
and U23445 (N_23445,N_10034,N_11693);
or U23446 (N_23446,N_18634,N_10869);
nor U23447 (N_23447,N_14329,N_15438);
nor U23448 (N_23448,N_12773,N_14970);
nand U23449 (N_23449,N_12182,N_18520);
or U23450 (N_23450,N_10758,N_10162);
nor U23451 (N_23451,N_17974,N_14262);
nand U23452 (N_23452,N_16948,N_17479);
nor U23453 (N_23453,N_17841,N_14170);
xnor U23454 (N_23454,N_15826,N_18398);
nor U23455 (N_23455,N_18174,N_19588);
nor U23456 (N_23456,N_14595,N_16468);
nor U23457 (N_23457,N_14255,N_18409);
and U23458 (N_23458,N_11062,N_13164);
nor U23459 (N_23459,N_18988,N_14804);
nor U23460 (N_23460,N_17852,N_14198);
and U23461 (N_23461,N_16866,N_15077);
xnor U23462 (N_23462,N_18199,N_16688);
nand U23463 (N_23463,N_16818,N_15973);
and U23464 (N_23464,N_13063,N_17757);
or U23465 (N_23465,N_11302,N_14298);
xor U23466 (N_23466,N_14371,N_15847);
or U23467 (N_23467,N_15539,N_10504);
xor U23468 (N_23468,N_10279,N_11139);
xnor U23469 (N_23469,N_10257,N_11226);
or U23470 (N_23470,N_14482,N_11334);
nor U23471 (N_23471,N_14311,N_19819);
or U23472 (N_23472,N_11383,N_17285);
or U23473 (N_23473,N_17732,N_19798);
nand U23474 (N_23474,N_17612,N_13937);
nand U23475 (N_23475,N_12871,N_10754);
nand U23476 (N_23476,N_10461,N_19846);
xor U23477 (N_23477,N_15397,N_17235);
or U23478 (N_23478,N_12601,N_19997);
nand U23479 (N_23479,N_17687,N_19888);
nand U23480 (N_23480,N_19046,N_10371);
xor U23481 (N_23481,N_16106,N_14444);
nor U23482 (N_23482,N_10803,N_13091);
and U23483 (N_23483,N_11559,N_14127);
and U23484 (N_23484,N_10096,N_11388);
xnor U23485 (N_23485,N_12062,N_15797);
nand U23486 (N_23486,N_10127,N_11183);
nor U23487 (N_23487,N_15888,N_16528);
nand U23488 (N_23488,N_13270,N_17372);
nand U23489 (N_23489,N_14283,N_13789);
or U23490 (N_23490,N_11430,N_12990);
nand U23491 (N_23491,N_11376,N_15467);
and U23492 (N_23492,N_18635,N_18514);
nand U23493 (N_23493,N_16694,N_14611);
or U23494 (N_23494,N_10645,N_18689);
and U23495 (N_23495,N_14639,N_19444);
or U23496 (N_23496,N_12434,N_14789);
or U23497 (N_23497,N_18501,N_14475);
and U23498 (N_23498,N_11114,N_11725);
and U23499 (N_23499,N_14880,N_17308);
xnor U23500 (N_23500,N_15308,N_14152);
nand U23501 (N_23501,N_13772,N_12244);
xnor U23502 (N_23502,N_19569,N_15119);
nand U23503 (N_23503,N_14610,N_12895);
xor U23504 (N_23504,N_14442,N_17812);
and U23505 (N_23505,N_18523,N_19013);
or U23506 (N_23506,N_13715,N_19141);
nand U23507 (N_23507,N_14581,N_13474);
xnor U23508 (N_23508,N_19194,N_18006);
or U23509 (N_23509,N_10061,N_13051);
or U23510 (N_23510,N_10580,N_12174);
nand U23511 (N_23511,N_12762,N_13360);
xor U23512 (N_23512,N_10687,N_15709);
and U23513 (N_23513,N_16840,N_19309);
or U23514 (N_23514,N_18304,N_18065);
xor U23515 (N_23515,N_17560,N_11424);
xor U23516 (N_23516,N_11128,N_10017);
nor U23517 (N_23517,N_14624,N_13226);
and U23518 (N_23518,N_11882,N_17579);
xnor U23519 (N_23519,N_16749,N_14301);
nor U23520 (N_23520,N_18336,N_16700);
xor U23521 (N_23521,N_15933,N_10862);
nor U23522 (N_23522,N_15927,N_11268);
xor U23523 (N_23523,N_19311,N_14348);
or U23524 (N_23524,N_19914,N_15070);
and U23525 (N_23525,N_16058,N_15463);
and U23526 (N_23526,N_13393,N_13488);
or U23527 (N_23527,N_18137,N_17016);
and U23528 (N_23528,N_19824,N_12835);
and U23529 (N_23529,N_19711,N_15960);
xor U23530 (N_23530,N_19259,N_16438);
or U23531 (N_23531,N_14369,N_17545);
nor U23532 (N_23532,N_10849,N_14282);
xnor U23533 (N_23533,N_10264,N_12348);
nor U23534 (N_23534,N_18041,N_19104);
or U23535 (N_23535,N_19166,N_18308);
nor U23536 (N_23536,N_11699,N_14643);
xnor U23537 (N_23537,N_10235,N_15511);
nor U23538 (N_23538,N_16433,N_18138);
and U23539 (N_23539,N_14048,N_16706);
xnor U23540 (N_23540,N_16870,N_10366);
xnor U23541 (N_23541,N_11691,N_12942);
nand U23542 (N_23542,N_18162,N_17025);
or U23543 (N_23543,N_17468,N_13833);
nand U23544 (N_23544,N_13059,N_17948);
nor U23545 (N_23545,N_14953,N_16603);
nor U23546 (N_23546,N_16316,N_15202);
and U23547 (N_23547,N_10526,N_16623);
xnor U23548 (N_23548,N_10975,N_18428);
xnor U23549 (N_23549,N_17374,N_18214);
or U23550 (N_23550,N_19886,N_13094);
and U23551 (N_23551,N_15496,N_17084);
and U23552 (N_23552,N_13168,N_14108);
or U23553 (N_23553,N_14077,N_18019);
nand U23554 (N_23554,N_12627,N_17942);
or U23555 (N_23555,N_17086,N_18786);
xnor U23556 (N_23556,N_14721,N_16889);
and U23557 (N_23557,N_12683,N_18347);
nand U23558 (N_23558,N_13808,N_16480);
xnor U23559 (N_23559,N_18931,N_11847);
or U23560 (N_23560,N_18608,N_10951);
nor U23561 (N_23561,N_13340,N_15734);
nor U23562 (N_23562,N_13046,N_10792);
nor U23563 (N_23563,N_11404,N_13451);
nand U23564 (N_23564,N_13011,N_15240);
and U23565 (N_23565,N_12644,N_11782);
and U23566 (N_23566,N_18183,N_10145);
nor U23567 (N_23567,N_14541,N_12503);
xor U23568 (N_23568,N_18896,N_11440);
nor U23569 (N_23569,N_13111,N_12260);
or U23570 (N_23570,N_10448,N_10935);
nor U23571 (N_23571,N_14459,N_12531);
nor U23572 (N_23572,N_15009,N_15905);
and U23573 (N_23573,N_10798,N_13337);
xnor U23574 (N_23574,N_13841,N_19176);
xor U23575 (N_23575,N_17449,N_11786);
or U23576 (N_23576,N_14563,N_18170);
xor U23577 (N_23577,N_10488,N_19388);
and U23578 (N_23578,N_15384,N_16429);
nor U23579 (N_23579,N_18298,N_16046);
xnor U23580 (N_23580,N_11229,N_12596);
nor U23581 (N_23581,N_14578,N_16927);
nor U23582 (N_23582,N_18405,N_13413);
nor U23583 (N_23583,N_12281,N_13704);
and U23584 (N_23584,N_12202,N_10654);
nand U23585 (N_23585,N_12191,N_18355);
and U23586 (N_23586,N_16784,N_15861);
and U23587 (N_23587,N_15153,N_10416);
and U23588 (N_23588,N_10962,N_10746);
and U23589 (N_23589,N_11264,N_18368);
or U23590 (N_23590,N_18293,N_16515);
nor U23591 (N_23591,N_13504,N_10874);
nor U23592 (N_23592,N_13582,N_11629);
or U23593 (N_23593,N_19284,N_16033);
xor U23594 (N_23594,N_11291,N_16263);
nor U23595 (N_23595,N_17735,N_18296);
xnor U23596 (N_23596,N_15487,N_14894);
xor U23597 (N_23597,N_19884,N_15233);
nand U23598 (N_23598,N_11086,N_17816);
and U23599 (N_23599,N_19089,N_12301);
nand U23600 (N_23600,N_13954,N_10102);
nor U23601 (N_23601,N_15235,N_10306);
xnor U23602 (N_23602,N_18666,N_18063);
nor U23603 (N_23603,N_16384,N_12923);
nor U23604 (N_23604,N_13421,N_14037);
nand U23605 (N_23605,N_14240,N_19823);
nand U23606 (N_23606,N_17884,N_10355);
and U23607 (N_23607,N_18290,N_14013);
and U23608 (N_23608,N_16376,N_15844);
nor U23609 (N_23609,N_18372,N_19447);
nor U23610 (N_23610,N_19863,N_13428);
nand U23611 (N_23611,N_12324,N_10864);
or U23612 (N_23612,N_18679,N_18909);
or U23613 (N_23613,N_15731,N_14487);
and U23614 (N_23614,N_17000,N_16473);
or U23615 (N_23615,N_16698,N_13693);
nor U23616 (N_23616,N_12736,N_18323);
xor U23617 (N_23617,N_17061,N_12748);
nor U23618 (N_23618,N_10142,N_11969);
xor U23619 (N_23619,N_17273,N_13098);
or U23620 (N_23620,N_17188,N_18716);
xor U23621 (N_23621,N_17901,N_16808);
nand U23622 (N_23622,N_18095,N_12996);
nand U23623 (N_23623,N_12197,N_14674);
nand U23624 (N_23624,N_11013,N_11568);
xor U23625 (N_23625,N_10940,N_14443);
nand U23626 (N_23626,N_15386,N_19239);
xnor U23627 (N_23627,N_10255,N_18763);
nor U23628 (N_23628,N_17119,N_17996);
nand U23629 (N_23629,N_15426,N_18397);
xor U23630 (N_23630,N_10955,N_14035);
and U23631 (N_23631,N_17592,N_16565);
xor U23632 (N_23632,N_15951,N_11078);
xnor U23633 (N_23633,N_14121,N_19413);
and U23634 (N_23634,N_12210,N_18790);
nand U23635 (N_23635,N_18722,N_18242);
nor U23636 (N_23636,N_14640,N_15784);
or U23637 (N_23637,N_16972,N_16177);
nor U23638 (N_23638,N_17887,N_14169);
nand U23639 (N_23639,N_19873,N_19202);
nor U23640 (N_23640,N_14460,N_15013);
or U23641 (N_23641,N_18926,N_13372);
or U23642 (N_23642,N_15048,N_17060);
nand U23643 (N_23643,N_11262,N_16732);
nand U23644 (N_23644,N_19271,N_11998);
nand U23645 (N_23645,N_16745,N_19963);
nand U23646 (N_23646,N_19999,N_16863);
xnor U23647 (N_23647,N_13597,N_18730);
or U23648 (N_23648,N_11026,N_13793);
or U23649 (N_23649,N_14006,N_19081);
nand U23650 (N_23650,N_15251,N_17414);
or U23651 (N_23651,N_12204,N_14345);
or U23652 (N_23652,N_18119,N_10094);
nand U23653 (N_23653,N_14538,N_10489);
xor U23654 (N_23654,N_16599,N_10481);
nand U23655 (N_23655,N_16643,N_13242);
nand U23656 (N_23656,N_18864,N_15060);
and U23657 (N_23657,N_10054,N_12272);
and U23658 (N_23658,N_18479,N_13113);
or U23659 (N_23659,N_11536,N_11210);
nand U23660 (N_23660,N_15469,N_18460);
and U23661 (N_23661,N_10377,N_19703);
nand U23662 (N_23662,N_10380,N_11996);
xnor U23663 (N_23663,N_14708,N_13461);
nand U23664 (N_23664,N_10322,N_16896);
or U23665 (N_23665,N_16092,N_15484);
xor U23666 (N_23666,N_15738,N_18862);
or U23667 (N_23667,N_16168,N_13902);
nor U23668 (N_23668,N_16454,N_16836);
nor U23669 (N_23669,N_18866,N_15102);
or U23670 (N_23670,N_14512,N_14260);
or U23671 (N_23671,N_13648,N_11910);
nand U23672 (N_23672,N_19401,N_12778);
or U23673 (N_23673,N_17246,N_14731);
and U23674 (N_23674,N_16104,N_10262);
xnor U23675 (N_23675,N_16101,N_17317);
nand U23676 (N_23676,N_15230,N_18253);
and U23677 (N_23677,N_13555,N_15936);
or U23678 (N_23678,N_14452,N_10492);
xnor U23679 (N_23679,N_14635,N_17157);
or U23680 (N_23680,N_17077,N_18231);
or U23681 (N_23681,N_19607,N_13909);
nand U23682 (N_23682,N_12921,N_11893);
xor U23683 (N_23683,N_10204,N_18872);
nor U23684 (N_23684,N_18875,N_12122);
or U23685 (N_23685,N_18444,N_11991);
nand U23686 (N_23686,N_10015,N_14243);
xor U23687 (N_23687,N_11448,N_16010);
nand U23688 (N_23688,N_16666,N_11792);
nand U23689 (N_23689,N_19012,N_15832);
and U23690 (N_23690,N_12786,N_14762);
nand U23691 (N_23691,N_12765,N_12453);
nand U23692 (N_23692,N_15549,N_11686);
and U23693 (N_23693,N_12091,N_13214);
nand U23694 (N_23694,N_10830,N_19719);
or U23695 (N_23695,N_10659,N_13257);
nor U23696 (N_23696,N_18388,N_14787);
or U23697 (N_23697,N_14414,N_19465);
xnor U23698 (N_23698,N_10072,N_14408);
nand U23699 (N_23699,N_13260,N_12918);
or U23700 (N_23700,N_15761,N_17201);
or U23701 (N_23701,N_15350,N_14137);
and U23702 (N_23702,N_19971,N_15296);
xnor U23703 (N_23703,N_16090,N_19512);
or U23704 (N_23704,N_14968,N_10392);
xnor U23705 (N_23705,N_14054,N_14588);
xnor U23706 (N_23706,N_12832,N_14912);
xnor U23707 (N_23707,N_18267,N_15284);
nor U23708 (N_23708,N_11213,N_12635);
xor U23709 (N_23709,N_12426,N_15811);
nor U23710 (N_23710,N_16945,N_14653);
or U23711 (N_23711,N_10113,N_13752);
nand U23712 (N_23712,N_10794,N_12154);
xnor U23713 (N_23713,N_13483,N_15889);
and U23714 (N_23714,N_12706,N_15746);
or U23715 (N_23715,N_14367,N_15157);
xor U23716 (N_23716,N_19250,N_14967);
nand U23717 (N_23717,N_14278,N_13027);
and U23718 (N_23718,N_10984,N_11721);
nor U23719 (N_23719,N_11500,N_12808);
and U23720 (N_23720,N_13400,N_18551);
xnor U23721 (N_23721,N_19146,N_17590);
xnor U23722 (N_23722,N_11580,N_10200);
or U23723 (N_23723,N_19474,N_18443);
xor U23724 (N_23724,N_14930,N_11270);
xor U23725 (N_23725,N_13977,N_11137);
nand U23726 (N_23726,N_15892,N_16834);
and U23727 (N_23727,N_11196,N_10443);
xnor U23728 (N_23728,N_17008,N_14535);
nand U23729 (N_23729,N_18669,N_11112);
and U23730 (N_23730,N_12472,N_13931);
nor U23731 (N_23731,N_14032,N_12323);
nand U23732 (N_23732,N_14195,N_19818);
xnor U23733 (N_23733,N_18264,N_15306);
and U23734 (N_23734,N_15216,N_19640);
nor U23735 (N_23735,N_16645,N_11159);
and U23736 (N_23736,N_15548,N_10154);
nor U23737 (N_23737,N_17883,N_16842);
nand U23738 (N_23738,N_15183,N_11378);
xnor U23739 (N_23739,N_13230,N_18995);
xor U23740 (N_23740,N_12927,N_15485);
nand U23741 (N_23741,N_13593,N_17678);
nor U23742 (N_23742,N_12941,N_15668);
or U23743 (N_23743,N_10785,N_10215);
xor U23744 (N_23744,N_19097,N_11701);
nand U23745 (N_23745,N_13626,N_13284);
xnor U23746 (N_23746,N_10890,N_17367);
and U23747 (N_23747,N_15134,N_16208);
xor U23748 (N_23748,N_13850,N_19910);
or U23749 (N_23749,N_19627,N_18812);
nand U23750 (N_23750,N_14056,N_19942);
nor U23751 (N_23751,N_18569,N_13854);
nand U23752 (N_23752,N_15279,N_12949);
and U23753 (N_23753,N_12303,N_12597);
or U23754 (N_23754,N_13384,N_10925);
and U23755 (N_23755,N_10617,N_11968);
nand U23756 (N_23756,N_15103,N_19314);
nand U23757 (N_23757,N_16953,N_11640);
xnor U23758 (N_23758,N_18147,N_19697);
nand U23759 (N_23759,N_13139,N_18956);
or U23760 (N_23760,N_11613,N_12752);
nor U23761 (N_23761,N_15435,N_15580);
and U23762 (N_23762,N_19159,N_13505);
xnor U23763 (N_23763,N_14297,N_16844);
xor U23764 (N_23764,N_11688,N_12721);
or U23765 (N_23765,N_16317,N_15136);
and U23766 (N_23766,N_14347,N_19708);
xor U23767 (N_23767,N_15545,N_11274);
nand U23768 (N_23768,N_17019,N_12540);
xnor U23769 (N_23769,N_17958,N_15146);
or U23770 (N_23770,N_14058,N_10114);
nand U23771 (N_23771,N_17531,N_19258);
xor U23772 (N_23772,N_13863,N_10369);
xor U23773 (N_23773,N_16771,N_15524);
nand U23774 (N_23774,N_11249,N_10282);
xnor U23775 (N_23775,N_18687,N_14379);
xor U23776 (N_23776,N_13074,N_17215);
xor U23777 (N_23777,N_11849,N_14254);
nand U23778 (N_23778,N_18820,N_14416);
and U23779 (N_23779,N_16593,N_11142);
and U23780 (N_23780,N_18920,N_14130);
nand U23781 (N_23781,N_10229,N_11501);
or U23782 (N_23782,N_19551,N_15040);
nand U23783 (N_23783,N_11052,N_17664);
nor U23784 (N_23784,N_17375,N_18472);
nand U23785 (N_23785,N_17371,N_11964);
nor U23786 (N_23786,N_16422,N_11532);
nand U23787 (N_23787,N_13717,N_15638);
and U23788 (N_23788,N_10494,N_18471);
nor U23789 (N_23789,N_19704,N_16164);
or U23790 (N_23790,N_10415,N_18600);
nor U23791 (N_23791,N_10560,N_13374);
nor U23792 (N_23792,N_14711,N_14522);
or U23793 (N_23793,N_10579,N_16820);
and U23794 (N_23794,N_15635,N_18749);
and U23795 (N_23795,N_18739,N_10473);
nor U23796 (N_23796,N_17675,N_19638);
or U23797 (N_23797,N_16773,N_13376);
nor U23798 (N_23798,N_14697,N_14072);
nor U23799 (N_23799,N_16503,N_17840);
nor U23800 (N_23800,N_14044,N_17460);
or U23801 (N_23801,N_12628,N_13817);
nor U23802 (N_23802,N_10372,N_12729);
or U23803 (N_23803,N_18427,N_11524);
nor U23804 (N_23804,N_19557,N_18676);
nand U23805 (N_23805,N_14476,N_16427);
and U23806 (N_23806,N_15361,N_12897);
nor U23807 (N_23807,N_14061,N_16277);
and U23808 (N_23808,N_12826,N_10610);
nor U23809 (N_23809,N_19019,N_15101);
nor U23810 (N_23810,N_16789,N_12338);
or U23811 (N_23811,N_13520,N_14224);
xor U23812 (N_23812,N_18873,N_16926);
or U23813 (N_23813,N_15834,N_12546);
nor U23814 (N_23814,N_15179,N_13653);
and U23815 (N_23815,N_14536,N_15567);
nor U23816 (N_23816,N_15127,N_13983);
nand U23817 (N_23817,N_11625,N_13506);
and U23818 (N_23818,N_13855,N_15374);
nor U23819 (N_23819,N_13547,N_14086);
nor U23820 (N_23820,N_16668,N_18519);
xor U23821 (N_23821,N_18798,N_19292);
xnor U23822 (N_23822,N_17417,N_10527);
nand U23823 (N_23823,N_13266,N_14368);
nand U23824 (N_23824,N_13223,N_11769);
and U23825 (N_23825,N_10786,N_13121);
nand U23826 (N_23826,N_11342,N_16970);
and U23827 (N_23827,N_11528,N_15217);
or U23828 (N_23828,N_12476,N_12947);
nor U23829 (N_23829,N_15824,N_11478);
nand U23830 (N_23830,N_16780,N_11323);
xnor U23831 (N_23831,N_18911,N_18413);
nor U23832 (N_23832,N_11107,N_16364);
and U23833 (N_23833,N_18369,N_13968);
nor U23834 (N_23834,N_14614,N_14833);
nor U23835 (N_23835,N_15776,N_12810);
and U23836 (N_23836,N_12337,N_16663);
or U23837 (N_23837,N_17500,N_13877);
or U23838 (N_23838,N_15425,N_10503);
xor U23839 (N_23839,N_19866,N_18767);
nand U23840 (N_23840,N_18370,N_15977);
or U23841 (N_23841,N_11201,N_11723);
and U23842 (N_23842,N_18564,N_13992);
and U23843 (N_23843,N_14231,N_17799);
and U23844 (N_23844,N_10685,N_15687);
and U23845 (N_23845,N_14477,N_11028);
and U23846 (N_23846,N_17599,N_17288);
and U23847 (N_23847,N_10275,N_19069);
nand U23848 (N_23848,N_18100,N_10673);
or U23849 (N_23849,N_19983,N_15658);
or U23850 (N_23850,N_17603,N_14910);
xnor U23851 (N_23851,N_19230,N_14984);
xnor U23852 (N_23852,N_12731,N_15055);
nor U23853 (N_23853,N_13008,N_16553);
or U23854 (N_23854,N_15881,N_15937);
nand U23855 (N_23855,N_10982,N_19067);
nor U23856 (N_23856,N_13557,N_11637);
nand U23857 (N_23857,N_13325,N_17171);
nand U23858 (N_23858,N_17203,N_10918);
xor U23859 (N_23859,N_12474,N_10436);
or U23860 (N_23860,N_10361,N_10159);
nor U23861 (N_23861,N_15787,N_16690);
nand U23862 (N_23862,N_11131,N_16288);
and U23863 (N_23863,N_17050,N_13878);
or U23864 (N_23864,N_18113,N_14613);
nor U23865 (N_23865,N_10695,N_16574);
nor U23866 (N_23866,N_16339,N_16909);
nor U23867 (N_23867,N_10945,N_19294);
and U23868 (N_23868,N_14799,N_14730);
and U23869 (N_23869,N_13427,N_14471);
nor U23870 (N_23870,N_18962,N_16093);
xnor U23871 (N_23871,N_12746,N_16301);
or U23872 (N_23872,N_18433,N_15006);
nand U23873 (N_23873,N_16197,N_10943);
and U23874 (N_23874,N_11553,N_10390);
nand U23875 (N_23875,N_10635,N_16624);
and U23876 (N_23876,N_19929,N_11540);
xor U23877 (N_23877,N_16281,N_17252);
nand U23878 (N_23878,N_12526,N_10246);
nor U23879 (N_23879,N_11188,N_12803);
nor U23880 (N_23880,N_13070,N_10367);
xor U23881 (N_23881,N_11587,N_18957);
or U23882 (N_23882,N_14257,N_12087);
and U23883 (N_23883,N_17122,N_14427);
nor U23884 (N_23884,N_10620,N_17475);
nand U23885 (N_23885,N_17444,N_11806);
and U23886 (N_23886,N_13128,N_19713);
and U23887 (N_23887,N_15836,N_13604);
nor U23888 (N_23888,N_19560,N_16138);
xnor U23889 (N_23889,N_14609,N_15018);
or U23890 (N_23890,N_16699,N_10134);
xnor U23891 (N_23891,N_10871,N_18255);
and U23892 (N_23892,N_11164,N_15954);
nor U23893 (N_23893,N_12728,N_14118);
nand U23894 (N_23894,N_18195,N_18918);
nand U23895 (N_23895,N_10266,N_15893);
and U23896 (N_23896,N_16910,N_19257);
and U23897 (N_23897,N_12167,N_12603);
and U23898 (N_23898,N_12742,N_15334);
nor U23899 (N_23899,N_14593,N_15775);
xnor U23900 (N_23900,N_13459,N_14770);
or U23901 (N_23901,N_15745,N_10614);
nand U23902 (N_23902,N_12952,N_18239);
nor U23903 (N_23903,N_16496,N_15203);
nor U23904 (N_23904,N_10498,N_19587);
nand U23905 (N_23905,N_19324,N_14823);
xor U23906 (N_23906,N_10693,N_17934);
or U23907 (N_23907,N_14977,N_10359);
nor U23908 (N_23908,N_12991,N_13396);
and U23909 (N_23909,N_17689,N_16437);
nor U23910 (N_23910,N_12890,N_12514);
nand U23911 (N_23911,N_12201,N_14620);
nand U23912 (N_23912,N_18655,N_15515);
nand U23913 (N_23913,N_19621,N_14646);
and U23914 (N_23914,N_12982,N_15759);
or U23915 (N_23915,N_10026,N_17837);
xnor U23916 (N_23916,N_16300,N_11653);
nor U23917 (N_23917,N_18469,N_14350);
or U23918 (N_23918,N_16619,N_16851);
and U23919 (N_23919,N_13538,N_14843);
nor U23920 (N_23920,N_17971,N_16403);
xnor U23921 (N_23921,N_12989,N_11851);
nand U23922 (N_23922,N_11783,N_14995);
xnor U23923 (N_23923,N_15565,N_19453);
xor U23924 (N_23924,N_11869,N_15556);
nor U23925 (N_23925,N_15148,N_17385);
nor U23926 (N_23926,N_17306,N_14997);
and U23927 (N_23927,N_18914,N_10073);
nor U23928 (N_23928,N_15576,N_12671);
or U23929 (N_23929,N_10606,N_13229);
nor U23930 (N_23930,N_13386,N_11504);
and U23931 (N_23931,N_12106,N_13654);
and U23932 (N_23932,N_13151,N_18186);
and U23933 (N_23933,N_16246,N_18860);
nor U23934 (N_23934,N_16928,N_13836);
and U23935 (N_23935,N_10834,N_12417);
nand U23936 (N_23936,N_10313,N_11301);
nand U23937 (N_23937,N_18568,N_11665);
nand U23938 (N_23938,N_11077,N_17492);
and U23939 (N_23939,N_19780,N_18953);
nand U23940 (N_23940,N_11784,N_13849);
nand U23941 (N_23941,N_13754,N_17703);
nand U23942 (N_23942,N_18205,N_11979);
nor U23943 (N_23943,N_12558,N_11548);
nand U23944 (N_23944,N_17764,N_10259);
xnor U23945 (N_23945,N_10732,N_15012);
xor U23946 (N_23946,N_12025,N_18870);
nand U23947 (N_23947,N_11180,N_15206);
nand U23948 (N_23948,N_10811,N_16081);
xnor U23949 (N_23949,N_12372,N_19880);
nor U23950 (N_23950,N_19165,N_18696);
nor U23951 (N_23951,N_11925,N_17556);
nor U23952 (N_23952,N_15692,N_11257);
or U23953 (N_23953,N_11967,N_10701);
and U23954 (N_23954,N_12125,N_18795);
or U23955 (N_23955,N_15434,N_15020);
nor U23956 (N_23956,N_19066,N_12632);
nand U23957 (N_23957,N_14119,N_14988);
nor U23958 (N_23958,N_10626,N_12906);
or U23959 (N_23959,N_12910,N_16308);
or U23960 (N_23960,N_11646,N_14438);
nand U23961 (N_23961,N_19092,N_11575);
nor U23962 (N_23962,N_17165,N_15599);
nand U23963 (N_23963,N_16608,N_13893);
xnor U23964 (N_23964,N_16170,N_12944);
xnor U23965 (N_23965,N_12240,N_18455);
and U23966 (N_23966,N_19500,N_15938);
nor U23967 (N_23967,N_19493,N_14553);
nor U23968 (N_23968,N_15820,N_14655);
xor U23969 (N_23969,N_14675,N_11203);
and U23970 (N_23970,N_18211,N_11666);
or U23971 (N_23971,N_10878,N_15618);
xor U23972 (N_23972,N_13848,N_10276);
xor U23973 (N_23973,N_10537,N_13663);
nor U23974 (N_23974,N_11853,N_13268);
nand U23975 (N_23975,N_19657,N_15084);
and U23976 (N_23976,N_15076,N_15805);
nor U23977 (N_23977,N_14752,N_19278);
or U23978 (N_23978,N_13442,N_14774);
xor U23979 (N_23979,N_17286,N_18141);
nand U23980 (N_23980,N_16113,N_12408);
nand U23981 (N_23981,N_13040,N_14709);
xnor U23982 (N_23982,N_12066,N_15238);
or U23983 (N_23983,N_19926,N_10066);
xnor U23984 (N_23984,N_18772,N_10721);
xor U23985 (N_23985,N_16589,N_12183);
nand U23986 (N_23986,N_12557,N_16212);
and U23987 (N_23987,N_12587,N_19006);
xor U23988 (N_23988,N_16681,N_12802);
xor U23989 (N_23989,N_12591,N_12608);
nand U23990 (N_23990,N_16117,N_16056);
nand U23991 (N_23991,N_15078,N_19008);
and U23992 (N_23992,N_17041,N_12688);
or U23993 (N_23993,N_19448,N_11687);
or U23994 (N_23994,N_19120,N_19764);
nand U23995 (N_23995,N_19743,N_15089);
nor U23996 (N_23996,N_17396,N_12071);
nor U23997 (N_23997,N_15640,N_17114);
nor U23998 (N_23998,N_16456,N_11585);
nand U23999 (N_23999,N_18500,N_11817);
or U24000 (N_24000,N_10070,N_17638);
and U24001 (N_24001,N_17715,N_13201);
and U24002 (N_24002,N_11754,N_17683);
or U24003 (N_24003,N_19237,N_10238);
xnor U24004 (N_24004,N_11167,N_12399);
or U24005 (N_24005,N_12759,N_13012);
or U24006 (N_24006,N_14099,N_11132);
and U24007 (N_24007,N_17309,N_18766);
or U24008 (N_24008,N_17351,N_17047);
and U24009 (N_24009,N_19307,N_11252);
nand U24010 (N_24010,N_18423,N_18319);
nand U24011 (N_24011,N_16015,N_18688);
and U24012 (N_24012,N_11530,N_10929);
and U24013 (N_24013,N_13711,N_14191);
or U24014 (N_24014,N_15321,N_15108);
or U24015 (N_24015,N_13811,N_11777);
nor U24016 (N_24016,N_10334,N_11604);
nand U24017 (N_24017,N_10431,N_19668);
nor U24018 (N_24018,N_15133,N_19133);
and U24019 (N_24019,N_17274,N_10291);
nand U24020 (N_24020,N_11161,N_10832);
or U24021 (N_24021,N_16405,N_13080);
nand U24022 (N_24022,N_17011,N_15655);
and U24023 (N_24023,N_13343,N_14829);
or U24024 (N_24024,N_13388,N_14004);
nand U24025 (N_24025,N_12815,N_13240);
nand U24026 (N_24026,N_18007,N_10914);
and U24027 (N_24027,N_17480,N_19175);
xnor U24028 (N_24028,N_15365,N_13294);
nor U24029 (N_24029,N_19938,N_12208);
xnor U24030 (N_24030,N_17783,N_19715);
nand U24031 (N_24031,N_18348,N_14511);
and U24032 (N_24032,N_14957,N_18632);
or U24033 (N_24033,N_13676,N_11266);
or U24034 (N_24034,N_15856,N_19139);
nor U24035 (N_24035,N_12005,N_18887);
xnor U24036 (N_24036,N_13852,N_14558);
xor U24037 (N_24037,N_19220,N_13486);
and U24038 (N_24038,N_18877,N_19263);
nor U24039 (N_24039,N_16740,N_16767);
and U24040 (N_24040,N_14903,N_16655);
nor U24041 (N_24041,N_11123,N_16100);
nand U24042 (N_24042,N_10903,N_11563);
or U24043 (N_24043,N_13782,N_17394);
and U24044 (N_24044,N_10987,N_11695);
or U24045 (N_24045,N_19416,N_13276);
and U24046 (N_24046,N_10294,N_12285);
and U24047 (N_24047,N_18190,N_17037);
nor U24048 (N_24048,N_12056,N_10243);
and U24049 (N_24049,N_16031,N_13364);
xnor U24050 (N_24050,N_10710,N_10345);
nor U24051 (N_24051,N_16817,N_12341);
nand U24052 (N_24052,N_10121,N_16755);
nand U24053 (N_24053,N_16189,N_15316);
nor U24054 (N_24054,N_13543,N_18781);
and U24055 (N_24055,N_14826,N_17669);
and U24056 (N_24056,N_19087,N_11145);
and U24057 (N_24057,N_14701,N_19458);
or U24058 (N_24058,N_13605,N_15429);
xnor U24059 (N_24059,N_19395,N_14647);
and U24060 (N_24060,N_17586,N_12315);
or U24061 (N_24061,N_12585,N_14817);
and U24062 (N_24062,N_17571,N_10265);
or U24063 (N_24063,N_14284,N_13382);
and U24064 (N_24064,N_14096,N_16378);
and U24065 (N_24065,N_11680,N_18852);
xnor U24066 (N_24066,N_16130,N_19348);
and U24067 (N_24067,N_18005,N_10937);
and U24068 (N_24068,N_11718,N_17857);
xor U24069 (N_24069,N_11324,N_19214);
or U24070 (N_24070,N_15908,N_17772);
nor U24071 (N_24071,N_19371,N_14554);
xnor U24072 (N_24072,N_18384,N_12092);
and U24073 (N_24073,N_13972,N_14641);
nand U24074 (N_24074,N_10978,N_19593);
xnor U24075 (N_24075,N_15049,N_11169);
xnor U24076 (N_24076,N_16869,N_19184);
xor U24077 (N_24077,N_18612,N_18759);
and U24078 (N_24078,N_16351,N_15555);
nand U24079 (N_24079,N_13336,N_15307);
nand U24080 (N_24080,N_18407,N_12131);
or U24081 (N_24081,N_18202,N_13826);
nand U24082 (N_24082,N_18560,N_15569);
nor U24083 (N_24083,N_14218,N_17940);
xnor U24084 (N_24084,N_19791,N_15488);
or U24085 (N_24085,N_11136,N_14850);
nor U24086 (N_24086,N_11937,N_14835);
nand U24087 (N_24087,N_12777,N_14914);
nor U24088 (N_24088,N_18785,N_17515);
xor U24089 (N_24089,N_15065,N_19628);
nand U24090 (N_24090,N_11477,N_12734);
xor U24091 (N_24091,N_13377,N_19265);
nor U24092 (N_24092,N_19454,N_10608);
nor U24093 (N_24093,N_17639,N_17191);
nand U24094 (N_24094,N_19323,N_11675);
nand U24095 (N_24095,N_17169,N_19768);
nand U24096 (N_24096,N_12037,N_12899);
nand U24097 (N_24097,N_12178,N_12583);
or U24098 (N_24098,N_12046,N_12774);
or U24099 (N_24099,N_15257,N_17487);
nor U24100 (N_24100,N_13963,N_17243);
and U24101 (N_24101,N_14340,N_11955);
nor U24102 (N_24102,N_12767,N_14586);
xor U24103 (N_24103,N_19887,N_14332);
and U24104 (N_24104,N_17859,N_17059);
nor U24105 (N_24105,N_13869,N_11437);
nor U24106 (N_24106,N_15390,N_12238);
nor U24107 (N_24107,N_15158,N_17619);
and U24108 (N_24108,N_19378,N_15005);
and U24109 (N_24109,N_18946,N_13723);
and U24110 (N_24110,N_18108,N_19973);
and U24111 (N_24111,N_14941,N_11034);
nor U24112 (N_24112,N_19470,N_11401);
and U24113 (N_24113,N_16677,N_14895);
and U24114 (N_24114,N_11999,N_13892);
and U24115 (N_24115,N_17712,N_17516);
nor U24116 (N_24116,N_17218,N_11671);
xor U24117 (N_24117,N_13026,N_16768);
and U24118 (N_24118,N_13381,N_17653);
or U24119 (N_24119,N_19592,N_13032);
nand U24120 (N_24120,N_14738,N_16563);
xnor U24121 (N_24121,N_12246,N_12849);
xnor U24122 (N_24122,N_12692,N_13706);
nor U24123 (N_24123,N_18395,N_15945);
nor U24124 (N_24124,N_16717,N_16772);
and U24125 (N_24125,N_18764,N_10633);
nand U24126 (N_24126,N_17263,N_19231);
nor U24127 (N_24127,N_19515,N_11983);
xnor U24128 (N_24128,N_11105,N_19342);
and U24129 (N_24129,N_12902,N_16990);
or U24130 (N_24130,N_16935,N_13219);
and U24131 (N_24131,N_17440,N_18778);
or U24132 (N_24132,N_12639,N_19671);
nor U24133 (N_24133,N_17020,N_15063);
or U24134 (N_24134,N_10573,N_11886);
nand U24135 (N_24135,N_17969,N_19480);
and U24136 (N_24136,N_17893,N_13564);
or U24137 (N_24137,N_10111,N_13320);
or U24138 (N_24138,N_15094,N_19867);
or U24139 (N_24139,N_10000,N_17688);
and U24140 (N_24140,N_18425,N_11100);
nor U24141 (N_24141,N_10338,N_11884);
nor U24142 (N_24142,N_12973,N_15994);
or U24143 (N_24143,N_17441,N_16478);
nand U24144 (N_24144,N_17448,N_16185);
and U24145 (N_24145,N_18328,N_18990);
nor U24146 (N_24146,N_10618,N_16036);
xnor U24147 (N_24147,N_13830,N_16055);
nand U24148 (N_24148,N_10182,N_19084);
nand U24149 (N_24149,N_18489,N_16746);
and U24150 (N_24150,N_14759,N_16856);
nand U24151 (N_24151,N_19100,N_13747);
or U24152 (N_24152,N_15716,N_14040);
nor U24153 (N_24153,N_13840,N_17826);
xnor U24154 (N_24154,N_16660,N_11812);
nor U24155 (N_24155,N_12553,N_14042);
and U24156 (N_24156,N_13664,N_10360);
nand U24157 (N_24157,N_13642,N_17076);
xnor U24158 (N_24158,N_15286,N_13234);
nor U24159 (N_24159,N_16559,N_15996);
nor U24160 (N_24160,N_12931,N_10727);
nor U24161 (N_24161,N_12645,N_15201);
nor U24162 (N_24162,N_18182,N_17598);
xnor U24163 (N_24163,N_13071,N_18552);
xnor U24164 (N_24164,N_14376,N_11014);
or U24165 (N_24165,N_16007,N_12019);
and U24166 (N_24166,N_17006,N_12259);
nand U24167 (N_24167,N_18345,N_17634);
and U24168 (N_24168,N_11195,N_17337);
nand U24169 (N_24169,N_13542,N_16956);
nor U24170 (N_24170,N_16680,N_18339);
nand U24171 (N_24171,N_15896,N_19072);
xor U24172 (N_24172,N_15349,N_14242);
xnor U24173 (N_24173,N_17057,N_15907);
nor U24174 (N_24174,N_14925,N_17662);
xor U24175 (N_24175,N_10729,N_18085);
nand U24176 (N_24176,N_13175,N_13548);
nand U24177 (N_24177,N_16540,N_17160);
xnor U24178 (N_24178,N_18122,N_10256);
nand U24179 (N_24179,N_10357,N_15262);
nand U24180 (N_24180,N_10823,N_10715);
xnor U24181 (N_24181,N_11562,N_11544);
and U24182 (N_24182,N_16139,N_10867);
or U24183 (N_24183,N_18748,N_13838);
or U24184 (N_24184,N_16841,N_15711);
nor U24185 (N_24185,N_12528,N_19312);
and U24186 (N_24186,N_18313,N_19613);
nand U24187 (N_24187,N_16535,N_13332);
and U24188 (N_24188,N_17797,N_16011);
or U24189 (N_24189,N_13822,N_19377);
nor U24190 (N_24190,N_13434,N_13416);
or U24191 (N_24191,N_16901,N_19964);
nand U24192 (N_24192,N_13149,N_14781);
nand U24193 (N_24193,N_13030,N_11791);
nand U24194 (N_24194,N_12329,N_10032);
xnor U24195 (N_24195,N_17139,N_17753);
nor U24196 (N_24196,N_15016,N_11355);
nand U24197 (N_24197,N_13775,N_11208);
and U24198 (N_24198,N_19439,N_15348);
nand U24199 (N_24199,N_19871,N_13998);
nand U24200 (N_24200,N_11538,N_14745);
nor U24201 (N_24201,N_13196,N_11813);
nand U24202 (N_24202,N_16049,N_14380);
nor U24203 (N_24203,N_10702,N_15399);
nor U24204 (N_24204,N_12040,N_14322);
nand U24205 (N_24205,N_11510,N_16129);
nand U24206 (N_24206,N_12749,N_18547);
nor U24207 (N_24207,N_13156,N_14933);
and U24208 (N_24208,N_14858,N_10677);
nand U24209 (N_24209,N_16913,N_17829);
xnor U24210 (N_24210,N_13182,N_13348);
or U24211 (N_24211,N_19383,N_13868);
nand U24212 (N_24212,N_11986,N_14079);
xor U24213 (N_24213,N_14607,N_14204);
xor U24214 (N_24214,N_16858,N_19086);
and U24215 (N_24215,N_12137,N_14664);
and U24216 (N_24216,N_12521,N_16652);
and U24217 (N_24217,N_12382,N_17152);
nor U24218 (N_24218,N_18014,N_13409);
nand U24219 (N_24219,N_15848,N_16541);
xor U24220 (N_24220,N_12478,N_14232);
nor U24221 (N_24221,N_16290,N_19599);
nor U24222 (N_24222,N_17421,N_13580);
nand U24223 (N_24223,N_13865,N_16587);
nor U24224 (N_24224,N_15839,N_13890);
and U24225 (N_24225,N_11465,N_12962);
and U24226 (N_24226,N_19485,N_14361);
and U24227 (N_24227,N_17314,N_17698);
and U24228 (N_24228,N_18540,N_15693);
xnor U24229 (N_24229,N_19881,N_10768);
nor U24230 (N_24230,N_14673,N_12751);
nor U24231 (N_24231,N_10544,N_19618);
and U24232 (N_24232,N_17956,N_17771);
nand U24233 (N_24233,N_14780,N_12543);
or U24234 (N_24234,N_10214,N_19921);
nor U24235 (N_24235,N_17465,N_17158);
or U24236 (N_24236,N_16445,N_17021);
nand U24237 (N_24237,N_14104,N_14940);
or U24238 (N_24238,N_11650,N_19562);
or U24239 (N_24239,N_17325,N_19185);
nor U24240 (N_24240,N_17749,N_14575);
nand U24241 (N_24241,N_18566,N_15312);
nor U24242 (N_24242,N_15572,N_17925);
xor U24243 (N_24243,N_13635,N_14714);
or U24244 (N_24244,N_17682,N_14189);
xnor U24245 (N_24245,N_13669,N_11146);
or U24246 (N_24246,N_13235,N_10596);
nor U24247 (N_24247,N_17279,N_19018);
and U24248 (N_24248,N_11091,N_15184);
and U24249 (N_24249,N_12097,N_19336);
or U24250 (N_24250,N_17434,N_14528);
and U24251 (N_24251,N_18450,N_18858);
xnor U24252 (N_24252,N_14716,N_11198);
nor U24253 (N_24253,N_16319,N_18884);
or U24254 (N_24254,N_14306,N_11353);
and U24255 (N_24255,N_16907,N_17657);
and U24256 (N_24256,N_12425,N_10052);
nor U24257 (N_24257,N_13228,N_12756);
xor U24258 (N_24258,N_16390,N_17094);
nand U24259 (N_24259,N_17323,N_17815);
nor U24260 (N_24260,N_13210,N_18839);
or U24261 (N_24261,N_13991,N_13613);
nand U24262 (N_24262,N_10807,N_16692);
nor U24263 (N_24263,N_12128,N_10884);
or U24264 (N_24264,N_15597,N_10290);
or U24265 (N_24265,N_10601,N_19586);
nor U24266 (N_24266,N_13766,N_12083);
nor U24267 (N_24267,N_19103,N_11835);
or U24268 (N_24268,N_11914,N_10486);
nor U24269 (N_24269,N_11282,N_16421);
or U24270 (N_24270,N_18818,N_11400);
and U24271 (N_24271,N_15395,N_19623);
nand U24272 (N_24272,N_14091,N_11591);
nand U24273 (N_24273,N_14463,N_14985);
xor U24274 (N_24274,N_12430,N_15219);
nand U24275 (N_24275,N_14312,N_10875);
and U24276 (N_24276,N_14290,N_12233);
xnor U24277 (N_24277,N_14690,N_18640);
or U24278 (N_24278,N_10098,N_15345);
nor U24279 (N_24279,N_16160,N_19229);
or U24280 (N_24280,N_19402,N_19597);
nand U24281 (N_24281,N_13942,N_12641);
nor U24282 (N_24282,N_10462,N_17074);
nand U24283 (N_24283,N_10533,N_12482);
nor U24284 (N_24284,N_18096,N_14288);
or U24285 (N_24285,N_16714,N_10374);
xnor U24286 (N_24286,N_15180,N_18828);
xnor U24287 (N_24287,N_17566,N_19108);
nand U24288 (N_24288,N_19524,N_11565);
and U24289 (N_24289,N_15500,N_18973);
and U24290 (N_24290,N_12859,N_17120);
nor U24291 (N_24291,N_17792,N_18626);
xnor U24292 (N_24292,N_18761,N_16025);
nor U24293 (N_24293,N_10382,N_10953);
and U24294 (N_24294,N_17079,N_18303);
and U24295 (N_24295,N_17808,N_17151);
or U24296 (N_24296,N_12884,N_18959);
and U24297 (N_24297,N_13106,N_14394);
nand U24298 (N_24298,N_13558,N_15002);
nor U24299 (N_24299,N_18966,N_14712);
or U24300 (N_24300,N_18216,N_13289);
nor U24301 (N_24301,N_19729,N_13697);
or U24302 (N_24302,N_13588,N_18507);
nor U24303 (N_24303,N_11756,N_10519);
xnor U24304 (N_24304,N_13249,N_13971);
and U24305 (N_24305,N_15891,N_12461);
nor U24306 (N_24306,N_18832,N_13042);
nand U24307 (N_24307,N_12293,N_11900);
or U24308 (N_24308,N_16673,N_14868);
or U24309 (N_24309,N_18576,N_14285);
or U24310 (N_24310,N_14253,N_12159);
nor U24311 (N_24311,N_12850,N_12104);
or U24312 (N_24312,N_12126,N_18774);
and U24313 (N_24313,N_11294,N_14256);
nand U24314 (N_24314,N_13958,N_18904);
nor U24315 (N_24315,N_11917,N_11269);
nand U24316 (N_24316,N_13783,N_11771);
and U24317 (N_24317,N_11254,N_13771);
nand U24318 (N_24318,N_17878,N_16215);
and U24319 (N_24319,N_16648,N_14486);
nand U24320 (N_24320,N_10700,N_17118);
nor U24321 (N_24321,N_14915,N_13927);
nor U24322 (N_24322,N_11143,N_15446);
nor U24323 (N_24323,N_12711,N_10604);
and U24324 (N_24324,N_16145,N_18810);
nor U24325 (N_24325,N_18617,N_10297);
xnor U24326 (N_24326,N_15604,N_19802);
nand U24327 (N_24327,N_10698,N_18613);
nand U24328 (N_24328,N_11664,N_10708);
nor U24329 (N_24329,N_19712,N_15057);
and U24330 (N_24330,N_15723,N_15862);
nand U24331 (N_24331,N_10018,N_17960);
nand U24332 (N_24332,N_11170,N_18526);
xor U24333 (N_24333,N_18879,N_17833);
xor U24334 (N_24334,N_17699,N_19706);
or U24335 (N_24335,N_13647,N_16958);
nor U24336 (N_24336,N_12733,N_10787);
nor U24337 (N_24337,N_17056,N_18223);
and U24338 (N_24338,N_11011,N_15275);
and U24339 (N_24339,N_18333,N_19063);
nor U24340 (N_24340,N_15527,N_16078);
nor U24341 (N_24341,N_17204,N_10055);
or U24342 (N_24342,N_18269,N_19134);
and U24343 (N_24343,N_12006,N_11616);
nor U24344 (N_24344,N_13475,N_11901);
and U24345 (N_24345,N_18158,N_16132);
xor U24346 (N_24346,N_13273,N_10619);
and U24347 (N_24347,N_19919,N_11735);
nand U24348 (N_24348,N_12108,N_12801);
and U24349 (N_24349,N_19372,N_18222);
nor U24350 (N_24350,N_17090,N_10201);
or U24351 (N_24351,N_11207,N_14537);
xor U24352 (N_24352,N_18292,N_12669);
and U24353 (N_24353,N_15528,N_12898);
nand U24354 (N_24354,N_14293,N_14483);
or U24355 (N_24355,N_12490,N_11320);
and U24356 (N_24356,N_17105,N_16196);
xnor U24357 (N_24357,N_12270,N_11309);
nor U24358 (N_24358,N_17027,N_16362);
nand U24359 (N_24359,N_11582,N_16191);
or U24360 (N_24360,N_15415,N_12809);
and U24361 (N_24361,N_10298,N_18034);
or U24362 (N_24362,N_12165,N_17767);
and U24363 (N_24363,N_12816,N_12951);
or U24364 (N_24364,N_16151,N_10524);
or U24365 (N_24365,N_10352,N_19456);
xnor U24366 (N_24366,N_16779,N_17426);
nor U24367 (N_24367,N_19832,N_16629);
nor U24368 (N_24368,N_13025,N_14012);
nand U24369 (N_24369,N_17997,N_14389);
and U24370 (N_24370,N_17552,N_14465);
xnor U24371 (N_24371,N_19869,N_14956);
xnor U24372 (N_24372,N_13291,N_16120);
xor U24373 (N_24373,N_11904,N_14095);
nor U24374 (N_24374,N_10566,N_16627);
nor U24375 (N_24375,N_18166,N_14932);
and U24376 (N_24376,N_10021,N_15953);
and U24377 (N_24377,N_18030,N_17931);
xnor U24378 (N_24378,N_16311,N_15163);
and U24379 (N_24379,N_14733,N_17846);
nand U24380 (N_24380,N_16938,N_18639);
nand U24381 (N_24381,N_11253,N_16213);
or U24382 (N_24382,N_18018,N_13205);
nor U24383 (N_24383,N_13633,N_11436);
nand U24384 (N_24384,N_18476,N_19786);
xnor U24385 (N_24385,N_13984,N_13851);
nor U24386 (N_24386,N_16676,N_17100);
xor U24387 (N_24387,N_12016,N_19544);
and U24388 (N_24388,N_12189,N_13408);
or U24389 (N_24389,N_19828,N_11895);
or U24390 (N_24390,N_18143,N_12418);
or U24391 (N_24391,N_13507,N_17149);
xor U24392 (N_24392,N_17711,N_10959);
xor U24393 (N_24393,N_17950,N_10843);
or U24394 (N_24394,N_11788,N_17632);
and U24395 (N_24395,N_12562,N_17398);
or U24396 (N_24396,N_11761,N_19464);
and U24397 (N_24397,N_17898,N_16937);
nor U24398 (N_24398,N_18112,N_19226);
or U24399 (N_24399,N_12385,N_17890);
nor U24400 (N_24400,N_11644,N_11820);
xor U24401 (N_24401,N_10109,N_15034);
nand U24402 (N_24402,N_12770,N_19626);
nand U24403 (N_24403,N_15253,N_18625);
or U24404 (N_24404,N_13404,N_11206);
nor U24405 (N_24405,N_18854,N_12822);
nand U24406 (N_24406,N_17777,N_14124);
nor U24407 (N_24407,N_19981,N_14704);
and U24408 (N_24408,N_14151,N_12036);
nand U24409 (N_24409,N_17787,N_15120);
nor U24410 (N_24410,N_15015,N_13472);
xor U24411 (N_24411,N_17718,N_10852);
nand U24412 (N_24412,N_14397,N_14384);
or U24413 (N_24413,N_12716,N_14413);
nand U24414 (N_24414,N_16586,N_17697);
nor U24415 (N_24415,N_10630,N_13449);
nor U24416 (N_24416,N_18637,N_17563);
nor U24417 (N_24417,N_18392,N_11654);
xor U24418 (N_24418,N_11093,N_10278);
nor U24419 (N_24419,N_11683,N_13601);
xnor U24420 (N_24420,N_17993,N_11402);
nor U24421 (N_24421,N_17005,N_19724);
nor U24422 (N_24422,N_18894,N_18134);
and U24423 (N_24423,N_11958,N_19852);
nand U24424 (N_24424,N_11810,N_14102);
xnor U24425 (N_24425,N_17791,N_19071);
xnor U24426 (N_24426,N_19144,N_15808);
nor U24427 (N_24427,N_19033,N_17422);
or U24428 (N_24428,N_10808,N_14172);
nor U24429 (N_24429,N_17591,N_17547);
or U24430 (N_24430,N_19285,N_16434);
and U24431 (N_24431,N_16815,N_17048);
xor U24432 (N_24432,N_19466,N_10093);
nand U24433 (N_24433,N_13940,N_14110);
and U24434 (N_24434,N_19274,N_14531);
nor U24435 (N_24435,N_16467,N_12076);
nand U24436 (N_24436,N_19186,N_16961);
and U24437 (N_24437,N_10860,N_11907);
nand U24438 (N_24438,N_17537,N_12010);
or U24439 (N_24439,N_15246,N_16124);
nor U24440 (N_24440,N_14946,N_17179);
and U24441 (N_24441,N_18177,N_10949);
or U24442 (N_24442,N_13184,N_13860);
xor U24443 (N_24443,N_12124,N_14228);
or U24444 (N_24444,N_13922,N_11049);
or U24445 (N_24445,N_11243,N_12336);
nor U24446 (N_24446,N_11919,N_12499);
or U24447 (N_24447,N_10636,N_12462);
or U24448 (N_24448,N_12536,N_17228);
or U24449 (N_24449,N_11632,N_11927);
nor U24450 (N_24450,N_12339,N_14038);
nand U24451 (N_24451,N_12277,N_11534);
nand U24452 (N_24452,N_11368,N_16955);
nor U24453 (N_24453,N_14372,N_13713);
nor U24454 (N_24454,N_15785,N_14187);
xnor U24455 (N_24455,N_13965,N_11178);
or U24456 (N_24456,N_15419,N_10202);
nand U24457 (N_24457,N_15726,N_10587);
nand U24458 (N_24458,N_12404,N_10053);
nand U24459 (N_24459,N_19723,N_14140);
and U24460 (N_24460,N_10621,N_10637);
and U24461 (N_24461,N_11838,N_19252);
nand U24462 (N_24462,N_16536,N_17033);
and U24463 (N_24463,N_14488,N_11572);
xnor U24464 (N_24464,N_10788,N_16693);
nand U24465 (N_24465,N_19469,N_17159);
and U24466 (N_24466,N_13349,N_14801);
nand U24467 (N_24467,N_12441,N_18619);
or U24468 (N_24468,N_19492,N_15113);
xnor U24469 (N_24469,N_11512,N_11489);
or U24470 (N_24470,N_17535,N_16661);
and U24471 (N_24471,N_18736,N_17290);
xor U24472 (N_24472,N_18487,N_12352);
nor U24473 (N_24473,N_13753,N_10152);
or U24474 (N_24474,N_17501,N_10623);
nand U24475 (N_24475,N_16231,N_12515);
xor U24476 (N_24476,N_11624,N_19096);
and U24477 (N_24477,N_16925,N_14550);
and U24478 (N_24478,N_15154,N_19933);
xnor U24479 (N_24479,N_10252,N_17873);
or U24480 (N_24480,N_18178,N_13705);
nand U24481 (N_24481,N_17131,N_11278);
or U24482 (N_24482,N_19467,N_14088);
or U24483 (N_24483,N_19755,N_11103);
or U24484 (N_24484,N_13581,N_14761);
nor U24485 (N_24485,N_19337,N_11678);
and U24486 (N_24486,N_10213,N_15735);
nor U24487 (N_24487,N_16786,N_14660);
and U24488 (N_24488,N_15849,N_17521);
nor U24489 (N_24489,N_14965,N_17628);
xor U24490 (N_24490,N_18343,N_13275);
nand U24491 (N_24491,N_12789,N_19911);
nor U24492 (N_24492,N_17790,N_19282);
nand U24493 (N_24493,N_16492,N_17295);
xnor U24494 (N_24494,N_18117,N_19553);
nand U24495 (N_24495,N_15679,N_13681);
nand U24496 (N_24496,N_15431,N_17001);
nor U24497 (N_24497,N_10168,N_13326);
or U24498 (N_24498,N_16190,N_17752);
nor U24499 (N_24499,N_13306,N_19472);
or U24500 (N_24500,N_13769,N_12510);
nor U24501 (N_24501,N_12384,N_16431);
xnor U24502 (N_24502,N_12038,N_11488);
xnor U24503 (N_24503,N_10323,N_19256);
nor U24504 (N_24504,N_11508,N_17489);
xnor U24505 (N_24505,N_13502,N_12464);
nor U24506 (N_24506,N_14736,N_14286);
xor U24507 (N_24507,N_16537,N_10110);
nor U24508 (N_24508,N_16348,N_19836);
nand U24509 (N_24509,N_16986,N_19594);
nor U24510 (N_24510,N_17737,N_17154);
or U24511 (N_24511,N_17068,N_10090);
nor U24512 (N_24512,N_13198,N_11963);
xnor U24513 (N_24513,N_14183,N_11634);
or U24514 (N_24514,N_13552,N_13731);
xnor U24515 (N_24515,N_10793,N_10240);
nand U24516 (N_24516,N_13494,N_13727);
and U24517 (N_24517,N_12616,N_14739);
xor U24518 (N_24518,N_11379,N_15590);
or U24519 (N_24519,N_12825,N_17403);
nand U24520 (N_24520,N_14539,N_11163);
or U24521 (N_24521,N_15086,N_17142);
and U24522 (N_24522,N_11741,N_17247);
xor U24523 (N_24523,N_14033,N_18733);
xor U24524 (N_24524,N_12779,N_17230);
nor U24525 (N_24525,N_10976,N_11475);
and U24526 (N_24526,N_19927,N_19559);
and U24527 (N_24527,N_12864,N_17354);
or U24528 (N_24528,N_10952,N_11877);
xor U24529 (N_24529,N_12387,N_14485);
nor U24530 (N_24530,N_11216,N_11759);
and U24531 (N_24531,N_19390,N_12588);
and U24532 (N_24532,N_15168,N_13763);
xnor U24533 (N_24533,N_12520,N_11729);
and U24534 (N_24534,N_19313,N_19434);
nand U24535 (N_24535,N_17052,N_18097);
or U24536 (N_24536,N_17128,N_10386);
or U24537 (N_24537,N_12449,N_18794);
or U24538 (N_24538,N_11217,N_12243);
nor U24539 (N_24539,N_15946,N_15686);
xor U24540 (N_24540,N_19979,N_14530);
nand U24541 (N_24541,N_18703,N_16684);
nand U24542 (N_24542,N_10944,N_17551);
or U24543 (N_24543,N_12518,N_14146);
nor U24544 (N_24544,N_16824,N_14666);
or U24545 (N_24545,N_12139,N_14507);
and U24546 (N_24546,N_18825,N_12966);
xor U24547 (N_24547,N_19283,N_18986);
nor U24548 (N_24548,N_17532,N_14168);
nand U24549 (N_24549,N_15401,N_10316);
or U24550 (N_24550,N_10870,N_16804);
nand U24551 (N_24551,N_16550,N_19690);
or U24552 (N_24552,N_14923,N_18595);
or U24553 (N_24553,N_15465,N_14021);
nor U24554 (N_24554,N_14604,N_14115);
or U24555 (N_24555,N_17126,N_14453);
xnor U24556 (N_24556,N_19758,N_13627);
nand U24557 (N_24557,N_16919,N_12458);
and U24558 (N_24558,N_16894,N_18233);
nand U24559 (N_24559,N_15147,N_14341);
or U24560 (N_24560,N_11277,N_14811);
and U24561 (N_24561,N_19145,N_11010);
nor U24562 (N_24562,N_13473,N_13391);
and U24563 (N_24563,N_13628,N_13672);
nor U24564 (N_24564,N_15151,N_16299);
nor U24565 (N_24565,N_14981,N_10718);
xor U24566 (N_24566,N_18775,N_14354);
or U24567 (N_24567,N_16302,N_15729);
nand U24568 (N_24568,N_13463,N_14827);
or U24569 (N_24569,N_16504,N_15682);
or U24570 (N_24570,N_10389,N_15358);
nor U24571 (N_24571,N_10067,N_15588);
nand U24572 (N_24572,N_19441,N_15355);
and U24573 (N_24573,N_19691,N_17617);
or U24574 (N_24574,N_13478,N_19135);
or U24575 (N_24575,N_17227,N_13825);
and U24576 (N_24576,N_19665,N_16985);
or U24577 (N_24577,N_16979,N_17108);
nor U24578 (N_24578,N_18287,N_16268);
and U24579 (N_24579,N_14735,N_16725);
or U24580 (N_24580,N_16214,N_13603);
and U24581 (N_24581,N_16387,N_10818);
nor U24582 (N_24582,N_10820,N_12901);
nor U24583 (N_24583,N_18574,N_10465);
nand U24584 (N_24584,N_14128,N_18841);
or U24585 (N_24585,N_19787,N_16073);
nor U24586 (N_24586,N_16102,N_14579);
nand U24587 (N_24587,N_15857,N_14807);
nor U24588 (N_24588,N_11798,N_15499);
nor U24589 (N_24589,N_14337,N_19111);
and U24590 (N_24590,N_14688,N_14886);
nand U24591 (N_24591,N_11902,N_12919);
or U24592 (N_24592,N_10988,N_18021);
nor U24593 (N_24593,N_19109,N_16392);
or U24594 (N_24594,N_13161,N_12534);
xnor U24595 (N_24595,N_19955,N_18936);
and U24596 (N_24596,N_19842,N_17549);
nand U24597 (N_24597,N_10909,N_14533);
nand U24598 (N_24598,N_10458,N_13058);
and U24599 (N_24599,N_11059,N_12527);
xor U24600 (N_24600,N_16303,N_15339);
and U24601 (N_24601,N_16369,N_11395);
and U24602 (N_24602,N_17293,N_12116);
or U24603 (N_24603,N_10917,N_15405);
and U24604 (N_24604,N_13112,N_15211);
nand U24605 (N_24605,N_10088,N_12646);
nand U24606 (N_24606,N_11120,N_17819);
nor U24607 (N_24607,N_10957,N_18389);
or U24608 (N_24608,N_14897,N_11314);
or U24609 (N_24609,N_16734,N_11012);
nor U24610 (N_24610,N_14450,N_17423);
or U24611 (N_24611,N_18445,N_13347);
nand U24612 (N_24612,N_19233,N_10858);
nand U24613 (N_24613,N_11864,N_15683);
and U24614 (N_24614,N_11117,N_13215);
or U24615 (N_24615,N_15942,N_12448);
nand U24616 (N_24616,N_18779,N_17083);
xnor U24617 (N_24617,N_19417,N_15367);
xor U24618 (N_24618,N_16859,N_12611);
and U24619 (N_24619,N_10131,N_18302);
and U24620 (N_24620,N_17088,N_12932);
xor U24621 (N_24621,N_18741,N_13787);
or U24622 (N_24622,N_18816,N_17755);
and U24623 (N_24623,N_15091,N_11790);
or U24624 (N_24624,N_17332,N_15305);
xor U24625 (N_24625,N_18187,N_12700);
nand U24626 (N_24626,N_11482,N_19192);
nand U24627 (N_24627,N_17297,N_19381);
and U24628 (N_24628,N_16687,N_18116);
and U24629 (N_24629,N_10578,N_13456);
xor U24630 (N_24630,N_12456,N_15106);
or U24631 (N_24631,N_12620,N_14402);
or U24632 (N_24632,N_19635,N_18747);
and U24633 (N_24633,N_13792,N_16097);
or U24634 (N_24634,N_19645,N_17109);
and U24635 (N_24635,N_17298,N_19528);
and U24636 (N_24636,N_13729,N_17255);
or U24637 (N_24637,N_18572,N_17835);
nor U24638 (N_24638,N_12823,N_11931);
xor U24639 (N_24639,N_13313,N_12400);
xor U24640 (N_24640,N_11374,N_13093);
xnor U24641 (N_24641,N_13041,N_16837);
or U24642 (N_24642,N_10158,N_19187);
nand U24643 (N_24643,N_11053,N_19328);
or U24644 (N_24644,N_15412,N_17004);
xnor U24645 (N_24645,N_18546,N_18165);
or U24646 (N_24646,N_16733,N_15568);
or U24647 (N_24647,N_12487,N_16656);
nand U24648 (N_24648,N_19300,N_18614);
nand U24649 (N_24649,N_11456,N_16274);
and U24650 (N_24650,N_18850,N_12147);
nor U24651 (N_24651,N_17923,N_11711);
and U24652 (N_24652,N_14928,N_17187);
xnor U24653 (N_24653,N_10169,N_16306);
or U24654 (N_24654,N_15753,N_19455);
nand U24655 (N_24655,N_17469,N_17029);
and U24656 (N_24656,N_11519,N_13395);
nand U24657 (N_24657,N_18633,N_13431);
or U24658 (N_24658,N_19025,N_12107);
xnor U24659 (N_24659,N_10383,N_11796);
xor U24660 (N_24660,N_12978,N_11878);
or U24661 (N_24661,N_11018,N_16283);
and U24662 (N_24662,N_15778,N_12135);
xor U24663 (N_24663,N_14724,N_16616);
and U24664 (N_24664,N_19490,N_14003);
nor U24665 (N_24665,N_19728,N_15854);
nand U24666 (N_24666,N_12617,N_11758);
nand U24667 (N_24667,N_18133,N_12194);
xor U24668 (N_24668,N_19662,N_10332);
nand U24669 (N_24669,N_16971,N_14877);
nand U24670 (N_24670,N_15858,N_19567);
or U24671 (N_24671,N_13916,N_14847);
xor U24672 (N_24672,N_14839,N_16495);
or U24673 (N_24673,N_13419,N_17864);
xnor U24674 (N_24674,N_18807,N_19737);
nor U24675 (N_24675,N_15666,N_15747);
nor U24676 (N_24676,N_11155,N_16475);
and U24677 (N_24677,N_16703,N_14791);
and U24678 (N_24678,N_17433,N_18930);
or U24679 (N_24679,N_15764,N_15061);
or U24680 (N_24680,N_14951,N_11005);
xor U24681 (N_24681,N_18148,N_16461);
and U24682 (N_24682,N_11954,N_19061);
nor U24683 (N_24683,N_15901,N_18978);
nor U24684 (N_24684,N_12566,N_12853);
and U24685 (N_24685,N_10148,N_19625);
xnor U24686 (N_24686,N_14349,N_19949);
nor U24687 (N_24687,N_17525,N_14983);
or U24688 (N_24688,N_10641,N_16861);
xor U24689 (N_24689,N_13007,N_17633);
xor U24690 (N_24690,N_12814,N_17693);
nor U24691 (N_24691,N_17610,N_18404);
nand U24692 (N_24692,N_17405,N_11537);
xnor U24693 (N_24693,N_18601,N_19178);
nor U24694 (N_24694,N_13673,N_19865);
xor U24695 (N_24695,N_10071,N_10406);
and U24696 (N_24696,N_10584,N_15170);
or U24697 (N_24697,N_18835,N_10765);
or U24698 (N_24698,N_11312,N_12267);
or U24699 (N_24699,N_11749,N_15090);
nor U24700 (N_24700,N_13004,N_14926);
nor U24701 (N_24701,N_11622,N_14490);
xor U24702 (N_24702,N_11989,N_18892);
or U24703 (N_24703,N_19885,N_19718);
nand U24704 (N_24704,N_17404,N_18928);
xor U24705 (N_24705,N_13468,N_18700);
and U24706 (N_24706,N_13481,N_15883);
or U24707 (N_24707,N_11158,N_15174);
xnor U24708 (N_24708,N_10656,N_16594);
or U24709 (N_24709,N_14942,N_18929);
xor U24710 (N_24710,N_14055,N_13197);
nor U24711 (N_24711,N_18987,N_16590);
and U24712 (N_24712,N_13126,N_14713);
and U24713 (N_24713,N_12013,N_17278);
nand U24714 (N_24714,N_19240,N_12709);
xnor U24715 (N_24715,N_13683,N_14669);
xnor U24716 (N_24716,N_11287,N_11962);
nand U24717 (N_24717,N_10495,N_10782);
or U24718 (N_24718,N_12613,N_17759);
and U24719 (N_24719,N_11338,N_14974);
xnor U24720 (N_24720,N_13466,N_19361);
and U24721 (N_24721,N_18876,N_15458);
nand U24722 (N_24722,N_12892,N_16229);
nand U24723 (N_24723,N_11138,N_18883);
and U24724 (N_24724,N_13471,N_12668);
nand U24725 (N_24725,N_12907,N_13256);
nand U24726 (N_24726,N_18996,N_18232);
and U24727 (N_24727,N_13283,N_14929);
or U24728 (N_24728,N_19769,N_14245);
nand U24729 (N_24729,N_14212,N_19568);
and U24730 (N_24730,N_10049,N_18960);
xnor U24731 (N_24731,N_12885,N_15708);
or U24732 (N_24732,N_18847,N_18353);
and U24733 (N_24733,N_12111,N_17588);
or U24734 (N_24734,N_11889,N_18869);
and U24735 (N_24735,N_15282,N_14748);
nor U24736 (N_24736,N_19032,N_12933);
and U24737 (N_24737,N_12195,N_12050);
and U24738 (N_24738,N_10446,N_15189);
and U24739 (N_24739,N_12205,N_10859);
nor U24740 (N_24740,N_16715,N_18431);
nor U24741 (N_24741,N_17909,N_14269);
or U24742 (N_24742,N_14678,N_12440);
or U24743 (N_24743,N_11360,N_13736);
nand U24744 (N_24744,N_19148,N_15398);
and U24745 (N_24745,N_19114,N_11953);
nor U24746 (N_24746,N_11452,N_12839);
nor U24747 (N_24747,N_14364,N_17568);
and U24748 (N_24748,N_13702,N_11762);
or U24749 (N_24749,N_13365,N_13371);
nor U24750 (N_24750,N_11602,N_17536);
nor U24751 (N_24751,N_17611,N_16162);
nand U24752 (N_24752,N_16529,N_14526);
nand U24753 (N_24753,N_17546,N_19853);
nand U24754 (N_24754,N_17355,N_16089);
or U24755 (N_24755,N_11408,N_11094);
nand U24756 (N_24756,N_14138,N_15740);
nand U24757 (N_24757,N_16402,N_16678);
nand U24758 (N_24758,N_10205,N_18844);
and U24759 (N_24759,N_16451,N_17458);
xnor U24760 (N_24760,N_19126,N_15035);
xor U24761 (N_24761,N_17627,N_13265);
xor U24762 (N_24762,N_16867,N_18974);
and U24763 (N_24763,N_13921,N_11370);
or U24764 (N_24764,N_18535,N_12576);
xnor U24765 (N_24765,N_10667,N_19666);
xor U24766 (N_24766,N_11271,N_15430);
or U24767 (N_24767,N_13806,N_15846);
or U24768 (N_24768,N_14992,N_14181);
xnor U24769 (N_24769,N_18466,N_18213);
nor U24770 (N_24770,N_16436,N_14749);
and U24771 (N_24771,N_17124,N_12556);
xor U24772 (N_24772,N_18840,N_10080);
nand U24773 (N_24773,N_17334,N_11154);
nand U24774 (N_24774,N_13594,N_18448);
xor U24775 (N_24775,N_15114,N_12484);
or U24776 (N_24776,N_10769,N_15975);
nor U24777 (N_24777,N_10105,N_12917);
xnor U24778 (N_24778,N_16976,N_18563);
xnor U24779 (N_24779,N_19045,N_17836);
xnor U24780 (N_24780,N_14596,N_17276);
xnor U24781 (N_24781,N_18377,N_19622);
xor U24782 (N_24782,N_16223,N_15377);
or U24783 (N_24783,N_10972,N_16352);
nand U24784 (N_24784,N_11070,N_17740);
and U24785 (N_24785,N_19572,N_12163);
xnor U24786 (N_24786,N_10474,N_17162);
xor U24787 (N_24787,N_17442,N_14520);
or U24788 (N_24788,N_19073,N_11681);
nand U24789 (N_24789,N_17234,N_17875);
or U24790 (N_24790,N_17428,N_16675);
nor U24791 (N_24791,N_18387,N_12675);
nor U24792 (N_24792,N_14947,N_18464);
nor U24793 (N_24793,N_16731,N_11753);
xnor U24794 (N_24794,N_15083,N_18064);
and U24795 (N_24795,N_17876,N_12354);
xnor U24796 (N_24796,N_12278,N_19501);
nor U24797 (N_24797,N_17741,N_13725);
and U24798 (N_24798,N_11227,N_16269);
nand U24799 (N_24799,N_12560,N_11067);
or U24800 (N_24800,N_14514,N_15873);
nor U24801 (N_24801,N_13232,N_15794);
or U24802 (N_24802,N_14582,N_19222);
or U24803 (N_24803,N_10271,N_13748);
xnor U24804 (N_24804,N_13798,N_14009);
xor U24805 (N_24805,N_13363,N_16760);
nand U24806 (N_24806,N_13809,N_10470);
xor U24807 (N_24807,N_11605,N_16221);
nor U24808 (N_24808,N_18024,N_12698);
xor U24809 (N_24809,N_15131,N_14071);
xnor U24810 (N_24810,N_12891,N_14230);
and U24811 (N_24811,N_11496,N_14602);
and U24812 (N_24812,N_13684,N_17654);
xnor U24813 (N_24813,N_15628,N_11066);
and U24814 (N_24814,N_18188,N_17756);
nand U24815 (N_24815,N_10753,N_16375);
xor U24816 (N_24816,N_15557,N_18259);
or U24817 (N_24817,N_12162,N_10745);
nand U24818 (N_24818,N_14300,N_15473);
nand U24819 (N_24819,N_14800,N_13309);
nand U24820 (N_24820,N_14094,N_13522);
xnor U24821 (N_24821,N_11080,N_15079);
or U24822 (N_24822,N_10130,N_10774);
and U24823 (N_24823,N_13515,N_17955);
xnor U24824 (N_24824,N_10545,N_16220);
nor U24825 (N_24825,N_12953,N_13023);
or U24826 (N_24826,N_17327,N_11047);
nand U24827 (N_24827,N_16483,N_12121);
and U24828 (N_24828,N_18156,N_13321);
xor U24829 (N_24829,N_17073,N_17905);
nand U24830 (N_24830,N_18099,N_16781);
nor U24831 (N_24831,N_18130,N_18681);
and U24832 (N_24832,N_16054,N_18606);
xor U24833 (N_24833,N_10838,N_19907);
nand U24834 (N_24834,N_17089,N_17222);
nand U24835 (N_24835,N_18031,N_10326);
or U24836 (N_24836,N_16472,N_19969);
and U24837 (N_24837,N_13994,N_12529);
and U24838 (N_24838,N_17751,N_18092);
or U24839 (N_24839,N_11551,N_19682);
and U24840 (N_24840,N_14837,N_19519);
nand U24841 (N_24841,N_11856,N_18624);
or U24842 (N_24842,N_10964,N_11069);
and U24843 (N_24843,N_19005,N_15281);
or U24844 (N_24844,N_14682,N_16307);
nand U24845 (N_24845,N_12467,N_12304);
and U24846 (N_24846,N_12881,N_16014);
nor U24847 (N_24847,N_14574,N_13031);
nand U24848 (N_24848,N_16538,N_19698);
or U24849 (N_24849,N_19039,N_16026);
xor U24850 (N_24850,N_10285,N_17392);
xor U24851 (N_24851,N_11189,N_13945);
and U24852 (N_24852,N_11407,N_14258);
and U24853 (N_24853,N_10837,N_12489);
and U24854 (N_24854,N_11122,N_15354);
nand U24855 (N_24855,N_16439,N_19683);
or U24856 (N_24856,N_17380,N_18948);
xor U24857 (N_24857,N_11057,N_11738);
xor U24858 (N_24858,N_17098,N_19701);
or U24859 (N_24859,N_18650,N_16984);
xor U24860 (N_24860,N_12271,N_13794);
or U24861 (N_24861,N_14473,N_10733);
xor U24862 (N_24862,N_13907,N_10189);
nand U24863 (N_24863,N_13827,N_16333);
xor U24864 (N_24864,N_10341,N_13013);
or U24865 (N_24865,N_14871,N_13735);
nand U24866 (N_24866,N_19748,N_18115);
or U24867 (N_24867,N_17910,N_18245);
nor U24868 (N_24868,N_11929,N_14917);
nor U24869 (N_24869,N_13138,N_10050);
nand U24870 (N_24870,N_17180,N_11007);
nor U24871 (N_24871,N_16831,N_13437);
nand U24872 (N_24872,N_13328,N_18504);
nor U24873 (N_24873,N_13224,N_19396);
or U24874 (N_24874,N_12754,N_17023);
xnor U24875 (N_24875,N_13532,N_19672);
xnor U24876 (N_24876,N_11410,N_19432);
nor U24877 (N_24877,N_15941,N_11412);
or U24878 (N_24878,N_13995,N_16531);
or U24879 (N_24879,N_19578,N_15659);
and U24880 (N_24880,N_16571,N_12035);
xnor U24881 (N_24881,N_14445,N_11950);
and U24882 (N_24882,N_12067,N_10220);
xnor U24883 (N_24883,N_19003,N_12306);
or U24884 (N_24884,N_15406,N_16499);
xor U24885 (N_24885,N_12542,N_11981);
nor U24886 (N_24886,N_11659,N_17102);
and U24887 (N_24887,N_18853,N_13657);
xor U24888 (N_24888,N_12180,N_13002);
nor U24889 (N_24889,N_18737,N_18738);
nand U24890 (N_24890,N_16254,N_19861);
nor U24891 (N_24891,N_11205,N_13519);
or U24892 (N_24892,N_13617,N_14540);
and U24893 (N_24893,N_19583,N_18241);
xnor U24894 (N_24894,N_12830,N_10307);
and U24895 (N_24895,N_16158,N_15968);
xor U24896 (N_24896,N_18511,N_10228);
xor U24897 (N_24897,N_13430,N_12466);
xnor U24898 (N_24898,N_16270,N_17976);
or U24899 (N_24899,N_19216,N_15733);
xor U24900 (N_24900,N_15689,N_12545);
nor U24901 (N_24901,N_18752,N_19673);
and U24902 (N_24902,N_11809,N_19803);
nor U24903 (N_24903,N_11457,N_19767);
nor U24904 (N_24904,N_12088,N_16868);
nor U24905 (N_24905,N_14157,N_11830);
nor U24906 (N_24906,N_18555,N_11050);
and U24907 (N_24907,N_16050,N_14150);
or U24908 (N_24908,N_19733,N_19290);
nand U24909 (N_24909,N_14114,N_19774);
nor U24910 (N_24910,N_15637,N_15254);
xnor U24911 (N_24911,N_15886,N_18565);
nor U24912 (N_24912,N_16180,N_10773);
nor U24913 (N_24913,N_17493,N_17395);
nor U24914 (N_24914,N_10865,N_11746);
and U24915 (N_24915,N_12502,N_10970);
and U24916 (N_24916,N_11547,N_13573);
nor U24917 (N_24917,N_18941,N_18750);
xnor U24918 (N_24918,N_13178,N_15895);
nor U24919 (N_24919,N_10373,N_11377);
nand U24920 (N_24920,N_16063,N_19351);
and U24921 (N_24921,N_19687,N_19571);
or U24922 (N_24922,N_15493,N_14765);
or U24923 (N_24923,N_10904,N_12096);
or U24924 (N_24924,N_13815,N_19614);
and U24925 (N_24925,N_13636,N_12241);
xnor U24926 (N_24926,N_11844,N_11912);
xor U24927 (N_24927,N_11584,N_19130);
xnor U24928 (N_24928,N_19603,N_12381);
and U24929 (N_24929,N_18556,N_18958);
xnor U24930 (N_24930,N_13829,N_15771);
and U24931 (N_24931,N_16987,N_16459);
nand U24932 (N_24932,N_13298,N_10728);
xnor U24933 (N_24933,N_15389,N_11389);
nor U24934 (N_24934,N_11403,N_18878);
xor U24935 (N_24935,N_14330,N_10047);
nand U24936 (N_24936,N_19659,N_14495);
xor U24937 (N_24937,N_18432,N_18248);
nor U24938 (N_24938,N_15598,N_19801);
xnor U24939 (N_24939,N_14700,N_17225);
and U24940 (N_24940,N_16359,N_12256);
and U24941 (N_24941,N_15533,N_19857);
or U24942 (N_24942,N_13569,N_18363);
or U24943 (N_24943,N_15317,N_19320);
and U24944 (N_24944,N_19197,N_12615);
nor U24945 (N_24945,N_12661,N_12974);
and U24946 (N_24946,N_16330,N_19950);
and U24947 (N_24947,N_12024,N_19241);
and U24948 (N_24948,N_17401,N_15591);
and U24949 (N_24949,N_17261,N_14132);
nand U24950 (N_24950,N_13901,N_15696);
xor U24951 (N_24951,N_12465,N_17618);
nor U24952 (N_24952,N_17907,N_15680);
nand U24953 (N_24953,N_15948,N_13804);
nand U24954 (N_24954,N_16061,N_11800);
nand U24955 (N_24955,N_11698,N_13619);
nand U24956 (N_24956,N_18436,N_15695);
nand U24957 (N_24957,N_11658,N_16035);
and U24958 (N_24958,N_19461,N_10658);
nor U24959 (N_24959,N_10177,N_13280);
xnor U24960 (N_24960,N_13286,N_19509);
nand U24961 (N_24961,N_10277,N_17457);
xnor U24962 (N_24962,N_19366,N_12513);
nand U24963 (N_24963,N_13807,N_15074);
or U24964 (N_24964,N_13982,N_16085);
and U24965 (N_24965,N_14848,N_11340);
xor U24966 (N_24966,N_11220,N_19391);
and U24967 (N_24967,N_18077,N_19833);
nor U24968 (N_24968,N_17237,N_10991);
nand U24969 (N_24969,N_14976,N_11709);
or U24970 (N_24970,N_16884,N_19505);
xor U24971 (N_24971,N_18440,N_16783);
or U24972 (N_24972,N_10150,N_19845);
xnor U24973 (N_24973,N_14363,N_15266);
xnor U24974 (N_24974,N_16358,N_10775);
nand U24975 (N_24975,N_16072,N_14419);
nor U24976 (N_24976,N_17484,N_18003);
nor U24977 (N_24977,N_15165,N_18371);
or U24978 (N_24978,N_10311,N_10199);
and U24979 (N_24979,N_19369,N_12934);
and U24980 (N_24980,N_16146,N_12867);
xnor U24981 (N_24981,N_18968,N_17026);
and U24982 (N_24982,N_17483,N_14569);
or U24983 (N_24983,N_16674,N_10913);
and U24984 (N_24984,N_13952,N_14325);
nor U24985 (N_24985,N_15714,N_13544);
nand U24986 (N_24986,N_14556,N_10321);
or U24987 (N_24987,N_19180,N_12245);
nand U24988 (N_24988,N_11797,N_19249);
nand U24989 (N_24989,N_17183,N_18277);
and U24990 (N_24990,N_19812,N_12086);
nor U24991 (N_24991,N_11833,N_14018);
xor U24992 (N_24992,N_10535,N_15774);
or U24993 (N_24993,N_12213,N_15649);
nor U24994 (N_24994,N_19421,N_16000);
nor U24995 (N_24995,N_16477,N_17739);
nand U24996 (N_24996,N_12548,N_17578);
nor U24997 (N_24997,N_10092,N_17051);
xor U24998 (N_24998,N_10950,N_19720);
and U24999 (N_24999,N_13908,N_18649);
and U25000 (N_25000,N_17352,N_14547);
xor U25001 (N_25001,N_15513,N_19920);
nor U25002 (N_25002,N_19364,N_14702);
xor U25003 (N_25003,N_10686,N_13907);
and U25004 (N_25004,N_19832,N_15930);
nand U25005 (N_25005,N_16969,N_10206);
or U25006 (N_25006,N_10723,N_10531);
nor U25007 (N_25007,N_12328,N_14274);
nor U25008 (N_25008,N_11303,N_15312);
or U25009 (N_25009,N_16270,N_17557);
nand U25010 (N_25010,N_10500,N_12025);
or U25011 (N_25011,N_12581,N_11612);
or U25012 (N_25012,N_14059,N_16703);
and U25013 (N_25013,N_18702,N_13063);
nor U25014 (N_25014,N_19607,N_16072);
nor U25015 (N_25015,N_19136,N_11094);
and U25016 (N_25016,N_11480,N_13537);
and U25017 (N_25017,N_12480,N_16712);
and U25018 (N_25018,N_19979,N_12136);
or U25019 (N_25019,N_10342,N_18022);
nor U25020 (N_25020,N_19829,N_19649);
and U25021 (N_25021,N_12915,N_11586);
or U25022 (N_25022,N_15858,N_15814);
or U25023 (N_25023,N_10495,N_12382);
nand U25024 (N_25024,N_19545,N_19934);
xnor U25025 (N_25025,N_19215,N_15505);
xnor U25026 (N_25026,N_17129,N_10755);
xor U25027 (N_25027,N_12995,N_15419);
xnor U25028 (N_25028,N_19728,N_19784);
nand U25029 (N_25029,N_15966,N_13753);
nor U25030 (N_25030,N_19868,N_19998);
nor U25031 (N_25031,N_12220,N_12323);
or U25032 (N_25032,N_10312,N_17573);
and U25033 (N_25033,N_17296,N_13504);
nor U25034 (N_25034,N_18933,N_18912);
and U25035 (N_25035,N_16758,N_14751);
nand U25036 (N_25036,N_10966,N_13828);
nand U25037 (N_25037,N_15553,N_10412);
nor U25038 (N_25038,N_13960,N_13789);
nand U25039 (N_25039,N_13286,N_11423);
and U25040 (N_25040,N_13002,N_14319);
or U25041 (N_25041,N_11188,N_12319);
nor U25042 (N_25042,N_17761,N_11463);
nand U25043 (N_25043,N_16754,N_18070);
nor U25044 (N_25044,N_12367,N_17904);
nand U25045 (N_25045,N_17521,N_19078);
and U25046 (N_25046,N_15582,N_19479);
nand U25047 (N_25047,N_12204,N_16030);
nor U25048 (N_25048,N_10543,N_10520);
and U25049 (N_25049,N_19577,N_16373);
or U25050 (N_25050,N_15744,N_18212);
nor U25051 (N_25051,N_18990,N_18241);
xor U25052 (N_25052,N_12129,N_19962);
xnor U25053 (N_25053,N_11729,N_18878);
or U25054 (N_25054,N_16652,N_18679);
nor U25055 (N_25055,N_14079,N_16077);
or U25056 (N_25056,N_14683,N_10158);
and U25057 (N_25057,N_12091,N_16468);
or U25058 (N_25058,N_13271,N_18187);
nor U25059 (N_25059,N_19526,N_18048);
or U25060 (N_25060,N_16482,N_13016);
nor U25061 (N_25061,N_18548,N_15949);
nand U25062 (N_25062,N_14083,N_11626);
and U25063 (N_25063,N_14831,N_11639);
or U25064 (N_25064,N_11755,N_13773);
xnor U25065 (N_25065,N_11934,N_19120);
nor U25066 (N_25066,N_16034,N_10313);
and U25067 (N_25067,N_13107,N_19609);
xor U25068 (N_25068,N_13621,N_13073);
or U25069 (N_25069,N_10663,N_13870);
or U25070 (N_25070,N_17254,N_18147);
nand U25071 (N_25071,N_18722,N_17910);
or U25072 (N_25072,N_18278,N_14702);
or U25073 (N_25073,N_19141,N_17374);
nor U25074 (N_25074,N_10512,N_12683);
xor U25075 (N_25075,N_18731,N_13847);
and U25076 (N_25076,N_15122,N_19682);
or U25077 (N_25077,N_15551,N_17278);
nand U25078 (N_25078,N_12937,N_13002);
or U25079 (N_25079,N_17667,N_16225);
nand U25080 (N_25080,N_10920,N_19661);
nand U25081 (N_25081,N_12806,N_12228);
xnor U25082 (N_25082,N_12817,N_16260);
and U25083 (N_25083,N_10515,N_16015);
nand U25084 (N_25084,N_16510,N_19123);
or U25085 (N_25085,N_15851,N_13021);
nand U25086 (N_25086,N_18168,N_16406);
or U25087 (N_25087,N_18928,N_19415);
and U25088 (N_25088,N_12692,N_19847);
or U25089 (N_25089,N_12569,N_10720);
or U25090 (N_25090,N_18138,N_17726);
or U25091 (N_25091,N_15490,N_16074);
or U25092 (N_25092,N_17909,N_11025);
nand U25093 (N_25093,N_19236,N_10890);
nor U25094 (N_25094,N_15736,N_15034);
xnor U25095 (N_25095,N_13842,N_19032);
and U25096 (N_25096,N_19344,N_17908);
nand U25097 (N_25097,N_14559,N_19193);
nand U25098 (N_25098,N_17935,N_19511);
xnor U25099 (N_25099,N_16376,N_11482);
or U25100 (N_25100,N_18779,N_11429);
or U25101 (N_25101,N_10112,N_15979);
or U25102 (N_25102,N_17744,N_15441);
xnor U25103 (N_25103,N_15953,N_11556);
and U25104 (N_25104,N_19121,N_14489);
or U25105 (N_25105,N_13790,N_13713);
xnor U25106 (N_25106,N_11605,N_10354);
nor U25107 (N_25107,N_17625,N_16828);
and U25108 (N_25108,N_17883,N_17861);
xnor U25109 (N_25109,N_18268,N_18818);
or U25110 (N_25110,N_10022,N_10351);
nor U25111 (N_25111,N_12276,N_19038);
nor U25112 (N_25112,N_18510,N_19291);
xnor U25113 (N_25113,N_18959,N_16893);
xnor U25114 (N_25114,N_17691,N_17227);
xor U25115 (N_25115,N_19267,N_17369);
nand U25116 (N_25116,N_12579,N_12575);
and U25117 (N_25117,N_14970,N_12259);
nand U25118 (N_25118,N_15461,N_13872);
or U25119 (N_25119,N_10914,N_15586);
nand U25120 (N_25120,N_10768,N_11138);
xor U25121 (N_25121,N_12333,N_19434);
nand U25122 (N_25122,N_13306,N_10595);
nand U25123 (N_25123,N_11912,N_19292);
and U25124 (N_25124,N_19370,N_17331);
and U25125 (N_25125,N_16523,N_11778);
nand U25126 (N_25126,N_17568,N_10397);
xnor U25127 (N_25127,N_18285,N_14909);
nand U25128 (N_25128,N_15913,N_13855);
xnor U25129 (N_25129,N_11193,N_11964);
nor U25130 (N_25130,N_19733,N_11382);
or U25131 (N_25131,N_10411,N_10661);
nor U25132 (N_25132,N_10496,N_13948);
xnor U25133 (N_25133,N_11440,N_16988);
and U25134 (N_25134,N_15830,N_19642);
nor U25135 (N_25135,N_13227,N_11126);
or U25136 (N_25136,N_17839,N_19335);
nand U25137 (N_25137,N_10276,N_16258);
or U25138 (N_25138,N_13020,N_11430);
nand U25139 (N_25139,N_12321,N_11664);
and U25140 (N_25140,N_16762,N_12149);
xor U25141 (N_25141,N_11811,N_16480);
and U25142 (N_25142,N_17855,N_12545);
nor U25143 (N_25143,N_17446,N_12936);
xor U25144 (N_25144,N_16862,N_17411);
xor U25145 (N_25145,N_17186,N_18118);
and U25146 (N_25146,N_19379,N_17143);
xnor U25147 (N_25147,N_18075,N_15318);
or U25148 (N_25148,N_12703,N_15384);
and U25149 (N_25149,N_13611,N_17486);
xnor U25150 (N_25150,N_17841,N_12744);
nor U25151 (N_25151,N_10291,N_17953);
and U25152 (N_25152,N_13833,N_14461);
and U25153 (N_25153,N_14127,N_18806);
nand U25154 (N_25154,N_15323,N_15941);
nand U25155 (N_25155,N_19152,N_16728);
nand U25156 (N_25156,N_14051,N_14026);
nor U25157 (N_25157,N_16852,N_15923);
and U25158 (N_25158,N_18266,N_17706);
and U25159 (N_25159,N_19941,N_14643);
nand U25160 (N_25160,N_15926,N_12679);
xnor U25161 (N_25161,N_12742,N_18154);
and U25162 (N_25162,N_11869,N_19633);
xnor U25163 (N_25163,N_16366,N_12625);
nand U25164 (N_25164,N_10302,N_11357);
nor U25165 (N_25165,N_11425,N_16968);
nor U25166 (N_25166,N_13934,N_10152);
or U25167 (N_25167,N_10877,N_14656);
and U25168 (N_25168,N_18652,N_12178);
nand U25169 (N_25169,N_15712,N_11818);
and U25170 (N_25170,N_19071,N_17619);
or U25171 (N_25171,N_11437,N_10966);
and U25172 (N_25172,N_17659,N_11045);
or U25173 (N_25173,N_12278,N_14156);
and U25174 (N_25174,N_19085,N_10365);
nand U25175 (N_25175,N_13981,N_16399);
nand U25176 (N_25176,N_18373,N_12877);
and U25177 (N_25177,N_14027,N_17362);
nand U25178 (N_25178,N_14190,N_19080);
nor U25179 (N_25179,N_13651,N_10206);
or U25180 (N_25180,N_19910,N_18993);
and U25181 (N_25181,N_17175,N_11911);
nor U25182 (N_25182,N_14342,N_17050);
xnor U25183 (N_25183,N_13803,N_13212);
nor U25184 (N_25184,N_18556,N_16533);
and U25185 (N_25185,N_10337,N_19832);
nor U25186 (N_25186,N_16036,N_17544);
nand U25187 (N_25187,N_12889,N_18566);
nand U25188 (N_25188,N_16778,N_18610);
nor U25189 (N_25189,N_13853,N_13760);
and U25190 (N_25190,N_14302,N_15886);
xor U25191 (N_25191,N_11986,N_16787);
and U25192 (N_25192,N_17705,N_12897);
xnor U25193 (N_25193,N_10169,N_17674);
nand U25194 (N_25194,N_11542,N_17478);
and U25195 (N_25195,N_18822,N_11547);
xor U25196 (N_25196,N_10952,N_10515);
or U25197 (N_25197,N_14794,N_11566);
and U25198 (N_25198,N_10545,N_12269);
xor U25199 (N_25199,N_13259,N_18138);
xnor U25200 (N_25200,N_18625,N_11638);
or U25201 (N_25201,N_14566,N_15336);
or U25202 (N_25202,N_19376,N_17444);
xor U25203 (N_25203,N_11008,N_19049);
and U25204 (N_25204,N_19822,N_18767);
nand U25205 (N_25205,N_14235,N_19603);
nand U25206 (N_25206,N_12579,N_14881);
or U25207 (N_25207,N_18950,N_14774);
nor U25208 (N_25208,N_15188,N_13828);
or U25209 (N_25209,N_15841,N_18220);
nand U25210 (N_25210,N_19645,N_10852);
nor U25211 (N_25211,N_14415,N_16063);
and U25212 (N_25212,N_17789,N_13591);
nand U25213 (N_25213,N_11523,N_15132);
nand U25214 (N_25214,N_13556,N_18682);
xnor U25215 (N_25215,N_15019,N_12176);
xor U25216 (N_25216,N_15332,N_17979);
xor U25217 (N_25217,N_16322,N_17598);
or U25218 (N_25218,N_10841,N_15746);
or U25219 (N_25219,N_11451,N_11714);
nor U25220 (N_25220,N_13438,N_10604);
and U25221 (N_25221,N_13191,N_12619);
and U25222 (N_25222,N_11692,N_13432);
and U25223 (N_25223,N_11360,N_12355);
nand U25224 (N_25224,N_19403,N_14867);
nor U25225 (N_25225,N_15792,N_17547);
xor U25226 (N_25226,N_18739,N_17065);
xor U25227 (N_25227,N_16762,N_13625);
and U25228 (N_25228,N_13883,N_16470);
xnor U25229 (N_25229,N_13655,N_16939);
and U25230 (N_25230,N_15548,N_17567);
or U25231 (N_25231,N_13407,N_18370);
and U25232 (N_25232,N_10558,N_15199);
or U25233 (N_25233,N_12641,N_14952);
and U25234 (N_25234,N_12692,N_12661);
xnor U25235 (N_25235,N_15924,N_13368);
xnor U25236 (N_25236,N_12530,N_11062);
or U25237 (N_25237,N_14959,N_15269);
and U25238 (N_25238,N_13118,N_13184);
xor U25239 (N_25239,N_17256,N_16233);
xor U25240 (N_25240,N_16770,N_17377);
nor U25241 (N_25241,N_13278,N_18291);
xnor U25242 (N_25242,N_12538,N_12720);
and U25243 (N_25243,N_17393,N_15701);
and U25244 (N_25244,N_14007,N_19996);
nor U25245 (N_25245,N_10310,N_13981);
or U25246 (N_25246,N_17584,N_10972);
nor U25247 (N_25247,N_18054,N_18134);
nor U25248 (N_25248,N_10086,N_13221);
nand U25249 (N_25249,N_10897,N_13141);
xor U25250 (N_25250,N_13335,N_14365);
or U25251 (N_25251,N_19204,N_14546);
nor U25252 (N_25252,N_11048,N_17883);
or U25253 (N_25253,N_13224,N_12770);
nor U25254 (N_25254,N_12007,N_19425);
nand U25255 (N_25255,N_14160,N_12378);
or U25256 (N_25256,N_14045,N_19009);
or U25257 (N_25257,N_15223,N_12618);
nor U25258 (N_25258,N_16179,N_12631);
nor U25259 (N_25259,N_15735,N_13349);
or U25260 (N_25260,N_10489,N_15344);
or U25261 (N_25261,N_15701,N_14967);
or U25262 (N_25262,N_17949,N_10529);
xor U25263 (N_25263,N_18779,N_15170);
nand U25264 (N_25264,N_19211,N_19675);
or U25265 (N_25265,N_17026,N_14100);
xor U25266 (N_25266,N_10503,N_15053);
nand U25267 (N_25267,N_10575,N_18489);
and U25268 (N_25268,N_14992,N_19472);
nor U25269 (N_25269,N_19310,N_14705);
nand U25270 (N_25270,N_12626,N_15929);
xnor U25271 (N_25271,N_15173,N_12776);
nand U25272 (N_25272,N_13719,N_10693);
nor U25273 (N_25273,N_12014,N_16986);
xor U25274 (N_25274,N_19264,N_12748);
and U25275 (N_25275,N_11476,N_10429);
and U25276 (N_25276,N_16285,N_17876);
or U25277 (N_25277,N_16832,N_17677);
nor U25278 (N_25278,N_11537,N_16028);
xnor U25279 (N_25279,N_13049,N_10657);
or U25280 (N_25280,N_15071,N_15653);
xnor U25281 (N_25281,N_15058,N_14680);
or U25282 (N_25282,N_18317,N_14151);
and U25283 (N_25283,N_16204,N_17071);
xor U25284 (N_25284,N_17151,N_15665);
and U25285 (N_25285,N_15699,N_13934);
nor U25286 (N_25286,N_19361,N_13950);
nand U25287 (N_25287,N_14921,N_18019);
and U25288 (N_25288,N_10246,N_11912);
xnor U25289 (N_25289,N_14184,N_11031);
xnor U25290 (N_25290,N_16421,N_17437);
and U25291 (N_25291,N_19526,N_10613);
xor U25292 (N_25292,N_13220,N_11432);
xnor U25293 (N_25293,N_13019,N_18971);
and U25294 (N_25294,N_18782,N_12134);
nor U25295 (N_25295,N_19486,N_11409);
nor U25296 (N_25296,N_17964,N_15524);
or U25297 (N_25297,N_19922,N_11288);
xor U25298 (N_25298,N_15227,N_13254);
xor U25299 (N_25299,N_15579,N_14005);
and U25300 (N_25300,N_15988,N_13622);
xor U25301 (N_25301,N_11911,N_11959);
xor U25302 (N_25302,N_10668,N_11045);
and U25303 (N_25303,N_17337,N_14609);
nand U25304 (N_25304,N_14900,N_18014);
or U25305 (N_25305,N_11791,N_12304);
and U25306 (N_25306,N_13769,N_14506);
xnor U25307 (N_25307,N_11237,N_15702);
and U25308 (N_25308,N_18817,N_19589);
and U25309 (N_25309,N_13967,N_18603);
nand U25310 (N_25310,N_15597,N_16367);
or U25311 (N_25311,N_15965,N_14622);
nor U25312 (N_25312,N_10053,N_11467);
xnor U25313 (N_25313,N_10520,N_12114);
nand U25314 (N_25314,N_12019,N_17160);
xor U25315 (N_25315,N_11603,N_16040);
or U25316 (N_25316,N_15994,N_14670);
nand U25317 (N_25317,N_10546,N_14090);
and U25318 (N_25318,N_17472,N_14684);
nor U25319 (N_25319,N_13705,N_15916);
nand U25320 (N_25320,N_12598,N_18733);
and U25321 (N_25321,N_19838,N_16508);
nor U25322 (N_25322,N_12693,N_13622);
xnor U25323 (N_25323,N_14226,N_19845);
nand U25324 (N_25324,N_19924,N_11372);
xnor U25325 (N_25325,N_14349,N_16909);
nor U25326 (N_25326,N_13770,N_14853);
and U25327 (N_25327,N_15909,N_10742);
and U25328 (N_25328,N_13458,N_10507);
or U25329 (N_25329,N_11875,N_16868);
nor U25330 (N_25330,N_12036,N_10333);
and U25331 (N_25331,N_19328,N_13963);
nand U25332 (N_25332,N_10034,N_15109);
or U25333 (N_25333,N_12849,N_13855);
xnor U25334 (N_25334,N_16649,N_15101);
nand U25335 (N_25335,N_15193,N_16641);
nor U25336 (N_25336,N_17765,N_19920);
and U25337 (N_25337,N_12940,N_16406);
xor U25338 (N_25338,N_12618,N_11447);
and U25339 (N_25339,N_11572,N_17679);
and U25340 (N_25340,N_17249,N_16565);
and U25341 (N_25341,N_17324,N_19514);
nor U25342 (N_25342,N_10282,N_18092);
or U25343 (N_25343,N_19103,N_14893);
or U25344 (N_25344,N_15562,N_10880);
and U25345 (N_25345,N_13208,N_10619);
or U25346 (N_25346,N_13961,N_11403);
nand U25347 (N_25347,N_13146,N_19744);
xnor U25348 (N_25348,N_11887,N_13771);
and U25349 (N_25349,N_12926,N_10586);
or U25350 (N_25350,N_10454,N_11860);
nor U25351 (N_25351,N_11821,N_11722);
or U25352 (N_25352,N_12591,N_16143);
nor U25353 (N_25353,N_19383,N_17706);
nor U25354 (N_25354,N_18053,N_15096);
and U25355 (N_25355,N_14001,N_19979);
or U25356 (N_25356,N_13680,N_14470);
xnor U25357 (N_25357,N_11033,N_18560);
nor U25358 (N_25358,N_15196,N_15991);
or U25359 (N_25359,N_12230,N_16285);
nand U25360 (N_25360,N_15183,N_17186);
xor U25361 (N_25361,N_18448,N_17137);
or U25362 (N_25362,N_16452,N_17898);
nand U25363 (N_25363,N_12033,N_18047);
and U25364 (N_25364,N_14076,N_12387);
nor U25365 (N_25365,N_12277,N_11749);
xor U25366 (N_25366,N_10493,N_16871);
or U25367 (N_25367,N_19395,N_19647);
or U25368 (N_25368,N_15216,N_19502);
or U25369 (N_25369,N_12885,N_16828);
xnor U25370 (N_25370,N_17351,N_15588);
nand U25371 (N_25371,N_10344,N_18949);
xnor U25372 (N_25372,N_15647,N_19037);
or U25373 (N_25373,N_14964,N_17356);
nor U25374 (N_25374,N_11908,N_18814);
nor U25375 (N_25375,N_19765,N_10645);
xnor U25376 (N_25376,N_11468,N_18742);
xor U25377 (N_25377,N_19331,N_10281);
nand U25378 (N_25378,N_15676,N_16411);
xor U25379 (N_25379,N_12374,N_17132);
nor U25380 (N_25380,N_14390,N_12879);
nor U25381 (N_25381,N_14431,N_18279);
nand U25382 (N_25382,N_12453,N_16465);
and U25383 (N_25383,N_17933,N_11211);
nand U25384 (N_25384,N_18203,N_17234);
xor U25385 (N_25385,N_10083,N_14818);
xnor U25386 (N_25386,N_16672,N_17313);
and U25387 (N_25387,N_17038,N_10691);
or U25388 (N_25388,N_14390,N_12260);
or U25389 (N_25389,N_11645,N_19183);
nand U25390 (N_25390,N_14781,N_12271);
nor U25391 (N_25391,N_15122,N_17717);
nor U25392 (N_25392,N_18731,N_19137);
and U25393 (N_25393,N_10671,N_14214);
and U25394 (N_25394,N_19439,N_19685);
nor U25395 (N_25395,N_14875,N_14985);
nand U25396 (N_25396,N_15016,N_10473);
nor U25397 (N_25397,N_16234,N_19592);
and U25398 (N_25398,N_19762,N_16254);
nand U25399 (N_25399,N_13630,N_16298);
and U25400 (N_25400,N_10315,N_11650);
or U25401 (N_25401,N_19771,N_19692);
nor U25402 (N_25402,N_15958,N_10712);
and U25403 (N_25403,N_15672,N_11294);
nor U25404 (N_25404,N_14092,N_10830);
or U25405 (N_25405,N_10720,N_18578);
or U25406 (N_25406,N_14369,N_11068);
and U25407 (N_25407,N_13260,N_17416);
or U25408 (N_25408,N_13592,N_17751);
nand U25409 (N_25409,N_13755,N_13763);
nor U25410 (N_25410,N_13830,N_11984);
or U25411 (N_25411,N_18253,N_13902);
and U25412 (N_25412,N_18823,N_11383);
and U25413 (N_25413,N_12521,N_13703);
nor U25414 (N_25414,N_14606,N_16287);
nand U25415 (N_25415,N_10504,N_15679);
or U25416 (N_25416,N_12511,N_14860);
and U25417 (N_25417,N_16998,N_19899);
nor U25418 (N_25418,N_18221,N_14164);
and U25419 (N_25419,N_14199,N_16342);
nor U25420 (N_25420,N_14771,N_11598);
nand U25421 (N_25421,N_19163,N_18959);
nor U25422 (N_25422,N_16910,N_17282);
or U25423 (N_25423,N_16270,N_17567);
nand U25424 (N_25424,N_14599,N_19733);
and U25425 (N_25425,N_12419,N_12393);
nor U25426 (N_25426,N_10664,N_15136);
or U25427 (N_25427,N_10475,N_11583);
and U25428 (N_25428,N_12017,N_15109);
and U25429 (N_25429,N_15851,N_16271);
or U25430 (N_25430,N_16132,N_16552);
nor U25431 (N_25431,N_11149,N_12626);
nor U25432 (N_25432,N_16916,N_13856);
nand U25433 (N_25433,N_18819,N_12149);
and U25434 (N_25434,N_10403,N_13299);
nand U25435 (N_25435,N_11069,N_15854);
or U25436 (N_25436,N_10842,N_15421);
and U25437 (N_25437,N_14416,N_14320);
nand U25438 (N_25438,N_11679,N_14328);
nor U25439 (N_25439,N_16169,N_15409);
xnor U25440 (N_25440,N_18951,N_15782);
xor U25441 (N_25441,N_15484,N_11363);
and U25442 (N_25442,N_18667,N_18897);
or U25443 (N_25443,N_19926,N_17216);
xor U25444 (N_25444,N_10864,N_11990);
or U25445 (N_25445,N_19695,N_11872);
nand U25446 (N_25446,N_18439,N_14277);
xor U25447 (N_25447,N_16245,N_15555);
xnor U25448 (N_25448,N_19081,N_12999);
or U25449 (N_25449,N_16073,N_17550);
and U25450 (N_25450,N_19737,N_16491);
nand U25451 (N_25451,N_14078,N_17931);
or U25452 (N_25452,N_19165,N_19134);
or U25453 (N_25453,N_15850,N_10385);
nand U25454 (N_25454,N_19374,N_15846);
nand U25455 (N_25455,N_12876,N_19144);
xor U25456 (N_25456,N_14910,N_10444);
nand U25457 (N_25457,N_19622,N_16295);
and U25458 (N_25458,N_16331,N_10133);
nor U25459 (N_25459,N_16447,N_13083);
nor U25460 (N_25460,N_13927,N_15569);
xnor U25461 (N_25461,N_11612,N_12379);
nor U25462 (N_25462,N_12798,N_14318);
xnor U25463 (N_25463,N_15647,N_15669);
nand U25464 (N_25464,N_17133,N_16510);
nand U25465 (N_25465,N_15223,N_13275);
and U25466 (N_25466,N_14902,N_13001);
xnor U25467 (N_25467,N_14727,N_17929);
xnor U25468 (N_25468,N_15772,N_19167);
xor U25469 (N_25469,N_10703,N_16890);
xor U25470 (N_25470,N_15041,N_19883);
xnor U25471 (N_25471,N_13618,N_19349);
nor U25472 (N_25472,N_18272,N_17017);
nor U25473 (N_25473,N_12265,N_17803);
and U25474 (N_25474,N_14959,N_11703);
nand U25475 (N_25475,N_18371,N_10563);
and U25476 (N_25476,N_11322,N_14811);
xnor U25477 (N_25477,N_15914,N_12615);
xnor U25478 (N_25478,N_10098,N_19849);
and U25479 (N_25479,N_14822,N_16376);
and U25480 (N_25480,N_17444,N_18175);
and U25481 (N_25481,N_15473,N_13886);
xnor U25482 (N_25482,N_19277,N_14504);
nand U25483 (N_25483,N_14669,N_17686);
nor U25484 (N_25484,N_13665,N_10223);
xor U25485 (N_25485,N_11771,N_19477);
and U25486 (N_25486,N_19963,N_15058);
nand U25487 (N_25487,N_15634,N_12708);
nand U25488 (N_25488,N_15010,N_10523);
xnor U25489 (N_25489,N_18303,N_17380);
and U25490 (N_25490,N_12548,N_12779);
nand U25491 (N_25491,N_16264,N_14399);
and U25492 (N_25492,N_14741,N_15772);
nand U25493 (N_25493,N_11276,N_18289);
and U25494 (N_25494,N_18502,N_13543);
and U25495 (N_25495,N_16932,N_16572);
nand U25496 (N_25496,N_13550,N_13355);
nand U25497 (N_25497,N_19053,N_14245);
nand U25498 (N_25498,N_16609,N_13011);
and U25499 (N_25499,N_13504,N_11419);
nor U25500 (N_25500,N_19468,N_17142);
xnor U25501 (N_25501,N_17322,N_10916);
nor U25502 (N_25502,N_15074,N_16891);
and U25503 (N_25503,N_17339,N_10072);
xor U25504 (N_25504,N_19791,N_11895);
xor U25505 (N_25505,N_16705,N_17500);
and U25506 (N_25506,N_15738,N_11951);
xnor U25507 (N_25507,N_15349,N_15142);
or U25508 (N_25508,N_18810,N_17274);
or U25509 (N_25509,N_16338,N_19949);
nand U25510 (N_25510,N_17112,N_17624);
or U25511 (N_25511,N_19292,N_12103);
nor U25512 (N_25512,N_17224,N_17098);
or U25513 (N_25513,N_13737,N_11507);
or U25514 (N_25514,N_15527,N_13551);
nor U25515 (N_25515,N_12998,N_18311);
and U25516 (N_25516,N_17529,N_14649);
or U25517 (N_25517,N_14511,N_14127);
nand U25518 (N_25518,N_19103,N_10725);
and U25519 (N_25519,N_17704,N_12460);
nand U25520 (N_25520,N_12344,N_17122);
nor U25521 (N_25521,N_11664,N_10311);
and U25522 (N_25522,N_11495,N_13260);
and U25523 (N_25523,N_15691,N_13552);
xnor U25524 (N_25524,N_17441,N_10135);
and U25525 (N_25525,N_18892,N_10743);
or U25526 (N_25526,N_14929,N_15763);
and U25527 (N_25527,N_17599,N_15575);
or U25528 (N_25528,N_16719,N_16873);
and U25529 (N_25529,N_17652,N_10507);
or U25530 (N_25530,N_19627,N_10673);
nor U25531 (N_25531,N_13283,N_14136);
or U25532 (N_25532,N_10619,N_12389);
and U25533 (N_25533,N_15184,N_14321);
xor U25534 (N_25534,N_15858,N_15647);
and U25535 (N_25535,N_13485,N_12380);
xor U25536 (N_25536,N_17038,N_19857);
nor U25537 (N_25537,N_14067,N_19083);
or U25538 (N_25538,N_12454,N_12907);
nand U25539 (N_25539,N_17147,N_13580);
or U25540 (N_25540,N_11063,N_17886);
nor U25541 (N_25541,N_10674,N_19896);
and U25542 (N_25542,N_12924,N_15221);
nand U25543 (N_25543,N_18006,N_17468);
nor U25544 (N_25544,N_17420,N_13428);
and U25545 (N_25545,N_14838,N_18650);
or U25546 (N_25546,N_10943,N_14188);
xnor U25547 (N_25547,N_13601,N_18131);
nor U25548 (N_25548,N_12029,N_17495);
or U25549 (N_25549,N_14247,N_12432);
xor U25550 (N_25550,N_12881,N_13812);
xnor U25551 (N_25551,N_10510,N_10607);
and U25552 (N_25552,N_12082,N_11460);
xnor U25553 (N_25553,N_15555,N_16058);
or U25554 (N_25554,N_17617,N_12250);
and U25555 (N_25555,N_10933,N_14380);
nand U25556 (N_25556,N_18826,N_13592);
and U25557 (N_25557,N_16060,N_10771);
or U25558 (N_25558,N_13491,N_14355);
or U25559 (N_25559,N_10894,N_17319);
xor U25560 (N_25560,N_17840,N_11178);
xor U25561 (N_25561,N_19285,N_11373);
and U25562 (N_25562,N_18445,N_16735);
nand U25563 (N_25563,N_17431,N_15677);
nor U25564 (N_25564,N_14625,N_12268);
or U25565 (N_25565,N_16637,N_17431);
xnor U25566 (N_25566,N_17311,N_11656);
nand U25567 (N_25567,N_12885,N_11051);
nor U25568 (N_25568,N_10175,N_16996);
nor U25569 (N_25569,N_18204,N_16397);
nand U25570 (N_25570,N_18608,N_13052);
and U25571 (N_25571,N_19755,N_17443);
nand U25572 (N_25572,N_18276,N_18247);
or U25573 (N_25573,N_19656,N_17321);
nand U25574 (N_25574,N_16867,N_12236);
nor U25575 (N_25575,N_14515,N_11857);
xnor U25576 (N_25576,N_15738,N_18228);
or U25577 (N_25577,N_17900,N_12727);
nor U25578 (N_25578,N_10955,N_18923);
nor U25579 (N_25579,N_13299,N_14232);
xor U25580 (N_25580,N_17441,N_10713);
and U25581 (N_25581,N_11235,N_19463);
and U25582 (N_25582,N_10357,N_11610);
xnor U25583 (N_25583,N_18813,N_11241);
and U25584 (N_25584,N_12246,N_17132);
nand U25585 (N_25585,N_19737,N_18855);
and U25586 (N_25586,N_14154,N_13232);
and U25587 (N_25587,N_10623,N_15412);
nor U25588 (N_25588,N_11567,N_15375);
nand U25589 (N_25589,N_14121,N_12377);
nor U25590 (N_25590,N_14727,N_11209);
nor U25591 (N_25591,N_18162,N_19725);
and U25592 (N_25592,N_19834,N_19256);
nand U25593 (N_25593,N_12861,N_12860);
nor U25594 (N_25594,N_14337,N_18961);
xor U25595 (N_25595,N_12859,N_10267);
and U25596 (N_25596,N_19801,N_17347);
nor U25597 (N_25597,N_18212,N_13231);
and U25598 (N_25598,N_17525,N_17631);
nor U25599 (N_25599,N_13840,N_12503);
or U25600 (N_25600,N_10737,N_15979);
nor U25601 (N_25601,N_12409,N_15804);
xnor U25602 (N_25602,N_17884,N_11693);
or U25603 (N_25603,N_13123,N_13512);
xnor U25604 (N_25604,N_15292,N_18216);
nand U25605 (N_25605,N_12513,N_18627);
nor U25606 (N_25606,N_12068,N_10907);
xor U25607 (N_25607,N_17662,N_17340);
nor U25608 (N_25608,N_18050,N_13193);
or U25609 (N_25609,N_14145,N_16792);
or U25610 (N_25610,N_16605,N_13055);
nand U25611 (N_25611,N_18404,N_13239);
and U25612 (N_25612,N_16741,N_12605);
and U25613 (N_25613,N_17205,N_18647);
xor U25614 (N_25614,N_11980,N_15300);
xnor U25615 (N_25615,N_11649,N_11626);
or U25616 (N_25616,N_15585,N_19846);
nor U25617 (N_25617,N_17775,N_18660);
and U25618 (N_25618,N_15687,N_17719);
nor U25619 (N_25619,N_12879,N_19918);
nor U25620 (N_25620,N_15940,N_15591);
or U25621 (N_25621,N_12426,N_14066);
nor U25622 (N_25622,N_11879,N_17121);
and U25623 (N_25623,N_15145,N_10878);
and U25624 (N_25624,N_14413,N_18437);
and U25625 (N_25625,N_19144,N_16936);
nor U25626 (N_25626,N_12798,N_11451);
nand U25627 (N_25627,N_11404,N_19064);
or U25628 (N_25628,N_18505,N_14088);
xnor U25629 (N_25629,N_15258,N_15778);
xor U25630 (N_25630,N_16016,N_17180);
or U25631 (N_25631,N_15637,N_13009);
nor U25632 (N_25632,N_18129,N_12715);
or U25633 (N_25633,N_10202,N_12562);
or U25634 (N_25634,N_13585,N_11768);
nor U25635 (N_25635,N_19596,N_14676);
nor U25636 (N_25636,N_13760,N_15569);
nand U25637 (N_25637,N_17853,N_10828);
nor U25638 (N_25638,N_13419,N_16131);
nand U25639 (N_25639,N_15773,N_12651);
or U25640 (N_25640,N_19695,N_12074);
nand U25641 (N_25641,N_10008,N_16535);
and U25642 (N_25642,N_13719,N_15552);
and U25643 (N_25643,N_15071,N_18046);
nor U25644 (N_25644,N_13133,N_12099);
xor U25645 (N_25645,N_12042,N_12246);
nor U25646 (N_25646,N_12950,N_14942);
and U25647 (N_25647,N_15066,N_10524);
nor U25648 (N_25648,N_12691,N_12560);
nor U25649 (N_25649,N_17636,N_18453);
and U25650 (N_25650,N_11922,N_11708);
nand U25651 (N_25651,N_11745,N_13438);
nand U25652 (N_25652,N_13283,N_18325);
xor U25653 (N_25653,N_19975,N_17884);
nor U25654 (N_25654,N_18347,N_10237);
xor U25655 (N_25655,N_16178,N_12170);
and U25656 (N_25656,N_18774,N_11486);
xnor U25657 (N_25657,N_10467,N_14367);
nand U25658 (N_25658,N_15406,N_16891);
or U25659 (N_25659,N_11042,N_10354);
and U25660 (N_25660,N_15847,N_12593);
xnor U25661 (N_25661,N_16875,N_11531);
or U25662 (N_25662,N_12469,N_13482);
nor U25663 (N_25663,N_13104,N_14046);
and U25664 (N_25664,N_16749,N_19103);
nand U25665 (N_25665,N_16419,N_16235);
and U25666 (N_25666,N_19930,N_17630);
xor U25667 (N_25667,N_13324,N_19989);
or U25668 (N_25668,N_10906,N_13346);
xor U25669 (N_25669,N_15070,N_15281);
and U25670 (N_25670,N_16558,N_16255);
or U25671 (N_25671,N_13909,N_13801);
or U25672 (N_25672,N_12441,N_11639);
nand U25673 (N_25673,N_13573,N_10993);
or U25674 (N_25674,N_16095,N_17015);
xnor U25675 (N_25675,N_17056,N_13438);
or U25676 (N_25676,N_11466,N_19701);
and U25677 (N_25677,N_10216,N_15960);
or U25678 (N_25678,N_12550,N_15195);
xnor U25679 (N_25679,N_19816,N_18880);
xnor U25680 (N_25680,N_10049,N_11506);
and U25681 (N_25681,N_10163,N_11940);
nor U25682 (N_25682,N_18353,N_14343);
nand U25683 (N_25683,N_16622,N_11165);
nor U25684 (N_25684,N_15700,N_12194);
and U25685 (N_25685,N_12829,N_10159);
nor U25686 (N_25686,N_13654,N_14629);
and U25687 (N_25687,N_15172,N_12280);
or U25688 (N_25688,N_16825,N_11954);
or U25689 (N_25689,N_13702,N_14552);
and U25690 (N_25690,N_15223,N_17303);
nand U25691 (N_25691,N_12488,N_13550);
xor U25692 (N_25692,N_12281,N_12716);
and U25693 (N_25693,N_17835,N_16600);
or U25694 (N_25694,N_17030,N_16917);
nor U25695 (N_25695,N_13345,N_19698);
nor U25696 (N_25696,N_14598,N_15031);
xor U25697 (N_25697,N_18957,N_15374);
nand U25698 (N_25698,N_19290,N_17779);
and U25699 (N_25699,N_19008,N_19250);
xor U25700 (N_25700,N_10856,N_13348);
and U25701 (N_25701,N_18626,N_14485);
nand U25702 (N_25702,N_17893,N_19792);
or U25703 (N_25703,N_14784,N_14584);
xnor U25704 (N_25704,N_17610,N_12517);
nand U25705 (N_25705,N_14204,N_17939);
nor U25706 (N_25706,N_17978,N_16258);
and U25707 (N_25707,N_15662,N_14751);
and U25708 (N_25708,N_14674,N_14484);
nor U25709 (N_25709,N_15250,N_18809);
and U25710 (N_25710,N_15963,N_11152);
and U25711 (N_25711,N_13744,N_18655);
and U25712 (N_25712,N_19664,N_16360);
and U25713 (N_25713,N_13936,N_14997);
or U25714 (N_25714,N_13650,N_19297);
or U25715 (N_25715,N_18602,N_16163);
nor U25716 (N_25716,N_13699,N_12174);
and U25717 (N_25717,N_13710,N_17573);
nor U25718 (N_25718,N_17547,N_18812);
nand U25719 (N_25719,N_16990,N_11813);
and U25720 (N_25720,N_12167,N_18309);
nand U25721 (N_25721,N_15005,N_19122);
nand U25722 (N_25722,N_12084,N_10995);
and U25723 (N_25723,N_11648,N_18092);
and U25724 (N_25724,N_19882,N_17090);
nor U25725 (N_25725,N_15424,N_10130);
nor U25726 (N_25726,N_11189,N_11599);
and U25727 (N_25727,N_14760,N_15366);
nor U25728 (N_25728,N_12085,N_12949);
nand U25729 (N_25729,N_18635,N_13224);
and U25730 (N_25730,N_17486,N_13191);
and U25731 (N_25731,N_19141,N_10768);
nand U25732 (N_25732,N_18198,N_19599);
or U25733 (N_25733,N_15656,N_15155);
xnor U25734 (N_25734,N_12957,N_10910);
xnor U25735 (N_25735,N_16213,N_17652);
or U25736 (N_25736,N_16888,N_19045);
or U25737 (N_25737,N_18369,N_19802);
or U25738 (N_25738,N_18497,N_19128);
nor U25739 (N_25739,N_17735,N_10371);
nand U25740 (N_25740,N_15955,N_19122);
nand U25741 (N_25741,N_15870,N_17895);
xor U25742 (N_25742,N_13708,N_15671);
or U25743 (N_25743,N_14962,N_15064);
or U25744 (N_25744,N_19488,N_18603);
or U25745 (N_25745,N_18223,N_10903);
nor U25746 (N_25746,N_10910,N_12116);
nor U25747 (N_25747,N_17650,N_11211);
xor U25748 (N_25748,N_16738,N_11740);
or U25749 (N_25749,N_18941,N_19671);
or U25750 (N_25750,N_11951,N_19598);
xor U25751 (N_25751,N_13458,N_10749);
xor U25752 (N_25752,N_10675,N_19909);
and U25753 (N_25753,N_14253,N_13258);
xnor U25754 (N_25754,N_15743,N_17947);
xnor U25755 (N_25755,N_11202,N_14988);
nand U25756 (N_25756,N_16466,N_12978);
xor U25757 (N_25757,N_12421,N_14530);
and U25758 (N_25758,N_18845,N_10010);
nand U25759 (N_25759,N_14311,N_13252);
xnor U25760 (N_25760,N_15983,N_10948);
xnor U25761 (N_25761,N_18430,N_16897);
and U25762 (N_25762,N_16833,N_10600);
xor U25763 (N_25763,N_16011,N_16566);
and U25764 (N_25764,N_17648,N_18324);
xor U25765 (N_25765,N_17040,N_19313);
nor U25766 (N_25766,N_17165,N_16299);
and U25767 (N_25767,N_18855,N_13607);
or U25768 (N_25768,N_11060,N_17179);
nand U25769 (N_25769,N_18106,N_13086);
and U25770 (N_25770,N_11470,N_19147);
nor U25771 (N_25771,N_11841,N_14749);
xor U25772 (N_25772,N_13691,N_11203);
or U25773 (N_25773,N_18143,N_18134);
nor U25774 (N_25774,N_14372,N_10166);
nand U25775 (N_25775,N_10032,N_12437);
xor U25776 (N_25776,N_10747,N_18751);
and U25777 (N_25777,N_19351,N_19024);
nor U25778 (N_25778,N_10803,N_15787);
nand U25779 (N_25779,N_13062,N_11777);
nor U25780 (N_25780,N_17825,N_17660);
or U25781 (N_25781,N_14284,N_14345);
nor U25782 (N_25782,N_14451,N_17357);
nand U25783 (N_25783,N_18277,N_14090);
nand U25784 (N_25784,N_19801,N_10122);
nand U25785 (N_25785,N_12237,N_15717);
nor U25786 (N_25786,N_17180,N_16475);
xnor U25787 (N_25787,N_12655,N_16238);
nand U25788 (N_25788,N_17062,N_17883);
xor U25789 (N_25789,N_11104,N_12318);
xnor U25790 (N_25790,N_15319,N_16852);
nand U25791 (N_25791,N_11100,N_10775);
xnor U25792 (N_25792,N_16858,N_17050);
nor U25793 (N_25793,N_15689,N_12717);
xnor U25794 (N_25794,N_13161,N_12665);
or U25795 (N_25795,N_18734,N_16064);
nand U25796 (N_25796,N_11130,N_15114);
or U25797 (N_25797,N_10319,N_13168);
or U25798 (N_25798,N_10543,N_14645);
xnor U25799 (N_25799,N_16138,N_19602);
nand U25800 (N_25800,N_19701,N_18056);
or U25801 (N_25801,N_19045,N_13123);
or U25802 (N_25802,N_13232,N_10625);
and U25803 (N_25803,N_13827,N_11234);
and U25804 (N_25804,N_16746,N_15789);
nor U25805 (N_25805,N_14021,N_19268);
xor U25806 (N_25806,N_16161,N_19500);
nand U25807 (N_25807,N_15311,N_14230);
and U25808 (N_25808,N_19540,N_17983);
or U25809 (N_25809,N_15685,N_15531);
or U25810 (N_25810,N_12129,N_11111);
nor U25811 (N_25811,N_13107,N_17276);
nand U25812 (N_25812,N_15038,N_18994);
and U25813 (N_25813,N_11345,N_19716);
nor U25814 (N_25814,N_13583,N_16464);
xor U25815 (N_25815,N_17519,N_10182);
nor U25816 (N_25816,N_14339,N_11486);
xor U25817 (N_25817,N_12035,N_17669);
xnor U25818 (N_25818,N_19252,N_17068);
nand U25819 (N_25819,N_18056,N_17643);
nor U25820 (N_25820,N_12002,N_18980);
and U25821 (N_25821,N_19599,N_14200);
nor U25822 (N_25822,N_18296,N_19327);
nor U25823 (N_25823,N_12518,N_19513);
xor U25824 (N_25824,N_11896,N_19992);
and U25825 (N_25825,N_16807,N_16929);
xor U25826 (N_25826,N_15436,N_15664);
nand U25827 (N_25827,N_13136,N_18791);
and U25828 (N_25828,N_19065,N_13363);
nand U25829 (N_25829,N_18539,N_10784);
xnor U25830 (N_25830,N_16663,N_13757);
or U25831 (N_25831,N_19235,N_17515);
and U25832 (N_25832,N_15961,N_12086);
xnor U25833 (N_25833,N_10018,N_10693);
nor U25834 (N_25834,N_11933,N_18030);
nor U25835 (N_25835,N_16632,N_11271);
and U25836 (N_25836,N_16800,N_11551);
or U25837 (N_25837,N_13242,N_15507);
nor U25838 (N_25838,N_19226,N_16619);
and U25839 (N_25839,N_16538,N_13044);
or U25840 (N_25840,N_14693,N_17900);
nor U25841 (N_25841,N_18367,N_19583);
xnor U25842 (N_25842,N_16942,N_14695);
nor U25843 (N_25843,N_15057,N_16012);
and U25844 (N_25844,N_13733,N_19112);
xor U25845 (N_25845,N_19869,N_14487);
nand U25846 (N_25846,N_18476,N_10676);
or U25847 (N_25847,N_19507,N_13502);
xnor U25848 (N_25848,N_19179,N_10936);
or U25849 (N_25849,N_12316,N_16058);
nor U25850 (N_25850,N_14663,N_18978);
nor U25851 (N_25851,N_18371,N_17693);
and U25852 (N_25852,N_10050,N_17554);
xor U25853 (N_25853,N_17580,N_17624);
xor U25854 (N_25854,N_12417,N_19498);
nor U25855 (N_25855,N_12993,N_11362);
xnor U25856 (N_25856,N_14357,N_13119);
xnor U25857 (N_25857,N_15239,N_12729);
or U25858 (N_25858,N_13200,N_18140);
nor U25859 (N_25859,N_19331,N_16198);
xor U25860 (N_25860,N_12478,N_14325);
nor U25861 (N_25861,N_15231,N_19199);
xnor U25862 (N_25862,N_14394,N_18877);
nand U25863 (N_25863,N_12432,N_16432);
xor U25864 (N_25864,N_18679,N_15504);
nor U25865 (N_25865,N_14476,N_12661);
nand U25866 (N_25866,N_13042,N_14980);
xnor U25867 (N_25867,N_14282,N_13929);
nand U25868 (N_25868,N_18385,N_11375);
xor U25869 (N_25869,N_15778,N_14483);
nand U25870 (N_25870,N_15627,N_18030);
nor U25871 (N_25871,N_14251,N_10739);
nor U25872 (N_25872,N_15108,N_18180);
or U25873 (N_25873,N_13845,N_10014);
nor U25874 (N_25874,N_16028,N_10201);
nand U25875 (N_25875,N_16759,N_13475);
xor U25876 (N_25876,N_13572,N_13562);
and U25877 (N_25877,N_10553,N_16987);
nand U25878 (N_25878,N_14350,N_16240);
and U25879 (N_25879,N_10149,N_18351);
nor U25880 (N_25880,N_19588,N_15392);
nand U25881 (N_25881,N_19176,N_11917);
nand U25882 (N_25882,N_12799,N_13932);
xnor U25883 (N_25883,N_12761,N_15295);
nor U25884 (N_25884,N_19834,N_17784);
or U25885 (N_25885,N_13589,N_16342);
xnor U25886 (N_25886,N_12104,N_11147);
xor U25887 (N_25887,N_18984,N_15024);
nor U25888 (N_25888,N_16402,N_13596);
or U25889 (N_25889,N_17291,N_14286);
and U25890 (N_25890,N_10296,N_17944);
or U25891 (N_25891,N_10008,N_10186);
and U25892 (N_25892,N_16625,N_10116);
nor U25893 (N_25893,N_10784,N_13616);
and U25894 (N_25894,N_10303,N_14600);
or U25895 (N_25895,N_10866,N_16584);
nand U25896 (N_25896,N_17965,N_12311);
nor U25897 (N_25897,N_19824,N_15570);
xor U25898 (N_25898,N_13244,N_12577);
nor U25899 (N_25899,N_19498,N_11525);
xnor U25900 (N_25900,N_14295,N_13199);
or U25901 (N_25901,N_18576,N_18023);
nand U25902 (N_25902,N_17878,N_17561);
or U25903 (N_25903,N_15179,N_13007);
and U25904 (N_25904,N_17804,N_18387);
nand U25905 (N_25905,N_11298,N_15761);
or U25906 (N_25906,N_16801,N_17478);
or U25907 (N_25907,N_16990,N_16917);
nor U25908 (N_25908,N_14290,N_15685);
nand U25909 (N_25909,N_14103,N_17648);
and U25910 (N_25910,N_12250,N_16180);
nand U25911 (N_25911,N_19996,N_13289);
nor U25912 (N_25912,N_11590,N_15613);
nor U25913 (N_25913,N_15937,N_13261);
or U25914 (N_25914,N_15504,N_19576);
nor U25915 (N_25915,N_13828,N_16544);
nand U25916 (N_25916,N_12845,N_12097);
nand U25917 (N_25917,N_16228,N_19137);
xor U25918 (N_25918,N_12654,N_12257);
and U25919 (N_25919,N_10107,N_15217);
or U25920 (N_25920,N_15449,N_10822);
or U25921 (N_25921,N_12598,N_19038);
and U25922 (N_25922,N_13266,N_13002);
nor U25923 (N_25923,N_15036,N_16247);
or U25924 (N_25924,N_18962,N_15817);
xnor U25925 (N_25925,N_15042,N_13419);
xor U25926 (N_25926,N_19159,N_16161);
or U25927 (N_25927,N_12852,N_19435);
nor U25928 (N_25928,N_17545,N_11105);
and U25929 (N_25929,N_13370,N_14527);
and U25930 (N_25930,N_13431,N_16262);
nand U25931 (N_25931,N_16901,N_19169);
xnor U25932 (N_25932,N_18846,N_10953);
nor U25933 (N_25933,N_11753,N_12384);
xnor U25934 (N_25934,N_15242,N_13719);
nor U25935 (N_25935,N_11637,N_12891);
and U25936 (N_25936,N_10342,N_15685);
xnor U25937 (N_25937,N_19142,N_19310);
or U25938 (N_25938,N_18725,N_14467);
xor U25939 (N_25939,N_12995,N_13344);
and U25940 (N_25940,N_14617,N_19581);
or U25941 (N_25941,N_10477,N_17366);
or U25942 (N_25942,N_18520,N_10951);
nand U25943 (N_25943,N_13357,N_10995);
nor U25944 (N_25944,N_11818,N_13590);
nand U25945 (N_25945,N_17120,N_11649);
or U25946 (N_25946,N_18540,N_10909);
nand U25947 (N_25947,N_15803,N_10069);
nor U25948 (N_25948,N_11122,N_12655);
and U25949 (N_25949,N_15933,N_14058);
and U25950 (N_25950,N_17921,N_13808);
nand U25951 (N_25951,N_11159,N_10896);
or U25952 (N_25952,N_15056,N_18919);
nor U25953 (N_25953,N_17816,N_10160);
nor U25954 (N_25954,N_14794,N_15988);
and U25955 (N_25955,N_11793,N_12442);
nor U25956 (N_25956,N_10214,N_17450);
nor U25957 (N_25957,N_14577,N_12042);
or U25958 (N_25958,N_17631,N_16517);
nor U25959 (N_25959,N_17545,N_10974);
or U25960 (N_25960,N_16034,N_11550);
or U25961 (N_25961,N_16351,N_17999);
or U25962 (N_25962,N_17008,N_15006);
nor U25963 (N_25963,N_13118,N_15191);
nand U25964 (N_25964,N_13396,N_12174);
and U25965 (N_25965,N_16400,N_11625);
nand U25966 (N_25966,N_18961,N_11023);
and U25967 (N_25967,N_14845,N_18025);
nand U25968 (N_25968,N_19843,N_19855);
or U25969 (N_25969,N_16958,N_11680);
and U25970 (N_25970,N_15837,N_10191);
and U25971 (N_25971,N_12624,N_18234);
and U25972 (N_25972,N_10090,N_15363);
nand U25973 (N_25973,N_12647,N_10343);
and U25974 (N_25974,N_13215,N_16853);
nor U25975 (N_25975,N_10976,N_19976);
nor U25976 (N_25976,N_11526,N_16301);
or U25977 (N_25977,N_12298,N_11802);
nand U25978 (N_25978,N_10710,N_15992);
xnor U25979 (N_25979,N_11099,N_13481);
nand U25980 (N_25980,N_14897,N_13337);
nand U25981 (N_25981,N_12039,N_18240);
xor U25982 (N_25982,N_13131,N_13711);
or U25983 (N_25983,N_15041,N_19188);
nand U25984 (N_25984,N_13521,N_11299);
nor U25985 (N_25985,N_11802,N_11880);
and U25986 (N_25986,N_15097,N_12087);
or U25987 (N_25987,N_10018,N_12203);
or U25988 (N_25988,N_18052,N_10062);
or U25989 (N_25989,N_15656,N_15675);
or U25990 (N_25990,N_13520,N_19654);
xnor U25991 (N_25991,N_11621,N_16599);
nor U25992 (N_25992,N_15274,N_10096);
nor U25993 (N_25993,N_17143,N_12694);
or U25994 (N_25994,N_18892,N_17431);
xor U25995 (N_25995,N_19995,N_11461);
nor U25996 (N_25996,N_13149,N_16266);
and U25997 (N_25997,N_17396,N_11298);
nor U25998 (N_25998,N_18358,N_13242);
xnor U25999 (N_25999,N_18579,N_13906);
or U26000 (N_26000,N_17193,N_18484);
xor U26001 (N_26001,N_15463,N_17563);
xnor U26002 (N_26002,N_17788,N_10168);
nand U26003 (N_26003,N_17159,N_15660);
nor U26004 (N_26004,N_10067,N_11404);
nor U26005 (N_26005,N_12644,N_14912);
nor U26006 (N_26006,N_15361,N_10003);
or U26007 (N_26007,N_14631,N_10514);
nand U26008 (N_26008,N_12952,N_18442);
and U26009 (N_26009,N_11420,N_11963);
nand U26010 (N_26010,N_19821,N_16398);
nor U26011 (N_26011,N_16035,N_14368);
nand U26012 (N_26012,N_11670,N_10933);
and U26013 (N_26013,N_19758,N_16141);
nand U26014 (N_26014,N_19616,N_14251);
nor U26015 (N_26015,N_10020,N_19523);
nor U26016 (N_26016,N_11745,N_19145);
and U26017 (N_26017,N_19368,N_12128);
or U26018 (N_26018,N_17927,N_17030);
nand U26019 (N_26019,N_18645,N_10313);
and U26020 (N_26020,N_10338,N_11994);
nor U26021 (N_26021,N_11324,N_19974);
nor U26022 (N_26022,N_17681,N_16395);
nor U26023 (N_26023,N_19979,N_16071);
xor U26024 (N_26024,N_19500,N_15117);
nand U26025 (N_26025,N_14237,N_13180);
or U26026 (N_26026,N_13691,N_12509);
xnor U26027 (N_26027,N_11945,N_14918);
or U26028 (N_26028,N_17695,N_16796);
and U26029 (N_26029,N_11624,N_11204);
or U26030 (N_26030,N_15655,N_11036);
and U26031 (N_26031,N_10254,N_15331);
and U26032 (N_26032,N_11927,N_14536);
nor U26033 (N_26033,N_16375,N_15860);
xnor U26034 (N_26034,N_15659,N_13560);
and U26035 (N_26035,N_12514,N_19663);
and U26036 (N_26036,N_15883,N_14223);
nand U26037 (N_26037,N_14338,N_16228);
nor U26038 (N_26038,N_16564,N_19504);
and U26039 (N_26039,N_16081,N_16013);
or U26040 (N_26040,N_11103,N_13866);
xor U26041 (N_26041,N_16266,N_14409);
nand U26042 (N_26042,N_17175,N_15465);
nand U26043 (N_26043,N_18544,N_17906);
nor U26044 (N_26044,N_11848,N_15569);
nor U26045 (N_26045,N_19988,N_14809);
xnor U26046 (N_26046,N_14577,N_19937);
or U26047 (N_26047,N_14215,N_15964);
xnor U26048 (N_26048,N_12418,N_18787);
nor U26049 (N_26049,N_10502,N_10237);
nor U26050 (N_26050,N_11564,N_12305);
xor U26051 (N_26051,N_13103,N_18173);
and U26052 (N_26052,N_12228,N_17403);
nand U26053 (N_26053,N_10328,N_12573);
nor U26054 (N_26054,N_16683,N_16085);
or U26055 (N_26055,N_13691,N_10310);
and U26056 (N_26056,N_18015,N_16788);
or U26057 (N_26057,N_13867,N_16821);
xor U26058 (N_26058,N_13346,N_10752);
or U26059 (N_26059,N_16889,N_15163);
and U26060 (N_26060,N_14485,N_19498);
or U26061 (N_26061,N_12704,N_14756);
and U26062 (N_26062,N_12387,N_13612);
and U26063 (N_26063,N_13616,N_12601);
nand U26064 (N_26064,N_13986,N_10803);
nor U26065 (N_26065,N_10062,N_16187);
or U26066 (N_26066,N_14194,N_11747);
and U26067 (N_26067,N_19348,N_16288);
nand U26068 (N_26068,N_12276,N_10103);
and U26069 (N_26069,N_11653,N_14059);
and U26070 (N_26070,N_19035,N_18047);
and U26071 (N_26071,N_14518,N_17220);
nor U26072 (N_26072,N_16738,N_13375);
and U26073 (N_26073,N_14542,N_17640);
xor U26074 (N_26074,N_18854,N_18322);
and U26075 (N_26075,N_17065,N_13660);
nand U26076 (N_26076,N_13209,N_12974);
and U26077 (N_26077,N_12181,N_16284);
nor U26078 (N_26078,N_19613,N_10182);
and U26079 (N_26079,N_19765,N_12809);
xor U26080 (N_26080,N_14809,N_19111);
and U26081 (N_26081,N_13574,N_19353);
nor U26082 (N_26082,N_13627,N_16420);
nor U26083 (N_26083,N_16285,N_13708);
xor U26084 (N_26084,N_17046,N_17168);
xnor U26085 (N_26085,N_16326,N_16236);
xnor U26086 (N_26086,N_14969,N_17633);
or U26087 (N_26087,N_11003,N_15212);
nand U26088 (N_26088,N_14873,N_18526);
xor U26089 (N_26089,N_16606,N_17016);
or U26090 (N_26090,N_15521,N_14798);
or U26091 (N_26091,N_17097,N_19282);
xor U26092 (N_26092,N_15583,N_11033);
and U26093 (N_26093,N_19240,N_10113);
xnor U26094 (N_26094,N_17710,N_13861);
nor U26095 (N_26095,N_18173,N_15839);
xor U26096 (N_26096,N_19084,N_12663);
and U26097 (N_26097,N_18119,N_10216);
or U26098 (N_26098,N_13487,N_13425);
or U26099 (N_26099,N_13040,N_10118);
or U26100 (N_26100,N_18981,N_14031);
nand U26101 (N_26101,N_12583,N_12495);
xnor U26102 (N_26102,N_19517,N_14295);
xor U26103 (N_26103,N_10400,N_18042);
nor U26104 (N_26104,N_12476,N_14122);
nor U26105 (N_26105,N_15722,N_15772);
xor U26106 (N_26106,N_15717,N_11862);
and U26107 (N_26107,N_17993,N_11858);
nand U26108 (N_26108,N_15993,N_14370);
and U26109 (N_26109,N_14526,N_11487);
and U26110 (N_26110,N_10898,N_16235);
or U26111 (N_26111,N_14721,N_15959);
nand U26112 (N_26112,N_17601,N_14388);
or U26113 (N_26113,N_15674,N_16178);
xor U26114 (N_26114,N_19959,N_14341);
xnor U26115 (N_26115,N_16426,N_14777);
nor U26116 (N_26116,N_14788,N_16163);
xor U26117 (N_26117,N_16532,N_12680);
xnor U26118 (N_26118,N_15739,N_19603);
nand U26119 (N_26119,N_10060,N_10943);
and U26120 (N_26120,N_12926,N_10682);
nand U26121 (N_26121,N_12965,N_16331);
nor U26122 (N_26122,N_16019,N_15747);
or U26123 (N_26123,N_17019,N_18343);
nand U26124 (N_26124,N_15474,N_14434);
xnor U26125 (N_26125,N_11385,N_12126);
xnor U26126 (N_26126,N_12330,N_18191);
nor U26127 (N_26127,N_18840,N_19325);
xnor U26128 (N_26128,N_16704,N_16474);
xor U26129 (N_26129,N_17460,N_15540);
nand U26130 (N_26130,N_10648,N_11176);
nor U26131 (N_26131,N_19630,N_16694);
nor U26132 (N_26132,N_11786,N_16071);
and U26133 (N_26133,N_19469,N_13947);
nor U26134 (N_26134,N_10713,N_13611);
nand U26135 (N_26135,N_11696,N_12117);
or U26136 (N_26136,N_10831,N_15727);
nor U26137 (N_26137,N_12288,N_15972);
nand U26138 (N_26138,N_18641,N_18433);
nor U26139 (N_26139,N_13924,N_19174);
or U26140 (N_26140,N_13993,N_11426);
or U26141 (N_26141,N_10305,N_14124);
nor U26142 (N_26142,N_10179,N_11862);
nor U26143 (N_26143,N_12343,N_18234);
and U26144 (N_26144,N_12789,N_16285);
xnor U26145 (N_26145,N_17865,N_14364);
or U26146 (N_26146,N_11549,N_16323);
or U26147 (N_26147,N_16235,N_13334);
or U26148 (N_26148,N_17893,N_16486);
and U26149 (N_26149,N_14335,N_13282);
nand U26150 (N_26150,N_10179,N_10714);
nor U26151 (N_26151,N_19216,N_16323);
nor U26152 (N_26152,N_15224,N_16643);
nand U26153 (N_26153,N_12717,N_11453);
nor U26154 (N_26154,N_13007,N_10304);
xnor U26155 (N_26155,N_10356,N_12093);
or U26156 (N_26156,N_15157,N_18043);
nand U26157 (N_26157,N_16417,N_17981);
nand U26158 (N_26158,N_12081,N_17306);
xnor U26159 (N_26159,N_19389,N_14710);
and U26160 (N_26160,N_11646,N_18586);
or U26161 (N_26161,N_12196,N_12647);
nor U26162 (N_26162,N_15147,N_12380);
or U26163 (N_26163,N_18273,N_15643);
or U26164 (N_26164,N_11196,N_16520);
and U26165 (N_26165,N_12983,N_12313);
nor U26166 (N_26166,N_10176,N_11041);
nor U26167 (N_26167,N_15699,N_13707);
and U26168 (N_26168,N_15337,N_17520);
xor U26169 (N_26169,N_15019,N_10909);
and U26170 (N_26170,N_16898,N_10804);
nand U26171 (N_26171,N_16676,N_19431);
and U26172 (N_26172,N_12669,N_11618);
nor U26173 (N_26173,N_11148,N_12550);
and U26174 (N_26174,N_15615,N_11595);
and U26175 (N_26175,N_13615,N_15515);
nor U26176 (N_26176,N_19847,N_14958);
nand U26177 (N_26177,N_11651,N_12289);
nor U26178 (N_26178,N_12302,N_17012);
nor U26179 (N_26179,N_12367,N_14268);
nand U26180 (N_26180,N_13855,N_19570);
xnor U26181 (N_26181,N_17883,N_19697);
nand U26182 (N_26182,N_11392,N_13362);
nor U26183 (N_26183,N_16600,N_18469);
xnor U26184 (N_26184,N_10524,N_19991);
nand U26185 (N_26185,N_10659,N_18072);
xnor U26186 (N_26186,N_13354,N_10983);
nand U26187 (N_26187,N_14244,N_11194);
nor U26188 (N_26188,N_16074,N_19172);
or U26189 (N_26189,N_13425,N_11778);
xor U26190 (N_26190,N_18811,N_10357);
xnor U26191 (N_26191,N_11349,N_14566);
nand U26192 (N_26192,N_15260,N_14880);
xnor U26193 (N_26193,N_18037,N_11501);
nand U26194 (N_26194,N_15394,N_12575);
and U26195 (N_26195,N_10260,N_10672);
nand U26196 (N_26196,N_17187,N_13375);
and U26197 (N_26197,N_13059,N_18652);
xnor U26198 (N_26198,N_15695,N_19208);
xnor U26199 (N_26199,N_11836,N_17476);
xor U26200 (N_26200,N_14690,N_17979);
nand U26201 (N_26201,N_10595,N_15671);
xnor U26202 (N_26202,N_18466,N_18858);
xnor U26203 (N_26203,N_14628,N_19598);
and U26204 (N_26204,N_11784,N_19963);
xor U26205 (N_26205,N_11867,N_10163);
or U26206 (N_26206,N_13610,N_15336);
xnor U26207 (N_26207,N_10406,N_15456);
nand U26208 (N_26208,N_15665,N_12885);
nor U26209 (N_26209,N_12910,N_13004);
nand U26210 (N_26210,N_17105,N_18241);
nor U26211 (N_26211,N_10420,N_19363);
or U26212 (N_26212,N_15935,N_10595);
and U26213 (N_26213,N_12711,N_11590);
and U26214 (N_26214,N_18261,N_14285);
nor U26215 (N_26215,N_15804,N_17903);
xor U26216 (N_26216,N_17075,N_18254);
and U26217 (N_26217,N_12955,N_15045);
and U26218 (N_26218,N_16623,N_11211);
or U26219 (N_26219,N_12177,N_14906);
or U26220 (N_26220,N_16927,N_15258);
or U26221 (N_26221,N_11623,N_17727);
and U26222 (N_26222,N_16376,N_12891);
nand U26223 (N_26223,N_16109,N_10885);
and U26224 (N_26224,N_16510,N_18310);
nor U26225 (N_26225,N_18400,N_14061);
or U26226 (N_26226,N_10713,N_19618);
nand U26227 (N_26227,N_18175,N_18015);
xnor U26228 (N_26228,N_13785,N_12637);
nor U26229 (N_26229,N_15981,N_16730);
or U26230 (N_26230,N_13951,N_14736);
nand U26231 (N_26231,N_13899,N_13035);
nor U26232 (N_26232,N_15953,N_11150);
nand U26233 (N_26233,N_17299,N_10963);
or U26234 (N_26234,N_13186,N_14859);
xnor U26235 (N_26235,N_11518,N_19283);
or U26236 (N_26236,N_10623,N_12472);
xnor U26237 (N_26237,N_13266,N_10151);
nand U26238 (N_26238,N_19934,N_16240);
nand U26239 (N_26239,N_17569,N_10485);
or U26240 (N_26240,N_18028,N_12385);
and U26241 (N_26241,N_10091,N_19762);
nor U26242 (N_26242,N_15458,N_10405);
nand U26243 (N_26243,N_18324,N_18607);
and U26244 (N_26244,N_18272,N_16274);
xor U26245 (N_26245,N_11766,N_14334);
nand U26246 (N_26246,N_15937,N_19496);
nor U26247 (N_26247,N_11493,N_17794);
and U26248 (N_26248,N_17815,N_12485);
and U26249 (N_26249,N_13394,N_12647);
and U26250 (N_26250,N_10830,N_14847);
nor U26251 (N_26251,N_15662,N_16769);
nand U26252 (N_26252,N_19046,N_16317);
xnor U26253 (N_26253,N_19495,N_18920);
nand U26254 (N_26254,N_18311,N_12048);
or U26255 (N_26255,N_12826,N_14296);
xor U26256 (N_26256,N_11807,N_18860);
nand U26257 (N_26257,N_19061,N_14369);
nor U26258 (N_26258,N_16864,N_10555);
nand U26259 (N_26259,N_13637,N_10778);
nand U26260 (N_26260,N_18060,N_16241);
or U26261 (N_26261,N_12755,N_17312);
nand U26262 (N_26262,N_17965,N_16343);
xnor U26263 (N_26263,N_11750,N_13633);
or U26264 (N_26264,N_14316,N_12215);
nand U26265 (N_26265,N_10975,N_16376);
or U26266 (N_26266,N_15278,N_16267);
xnor U26267 (N_26267,N_17110,N_19243);
nand U26268 (N_26268,N_10907,N_12155);
nor U26269 (N_26269,N_17789,N_18733);
xor U26270 (N_26270,N_19799,N_11184);
nor U26271 (N_26271,N_11426,N_12033);
or U26272 (N_26272,N_15905,N_13011);
or U26273 (N_26273,N_10525,N_17483);
nand U26274 (N_26274,N_13261,N_16771);
xnor U26275 (N_26275,N_13150,N_17825);
and U26276 (N_26276,N_19791,N_10699);
and U26277 (N_26277,N_14507,N_14939);
xor U26278 (N_26278,N_12653,N_18769);
xnor U26279 (N_26279,N_15187,N_18732);
nand U26280 (N_26280,N_14483,N_11347);
nor U26281 (N_26281,N_11750,N_19899);
nor U26282 (N_26282,N_12489,N_10774);
and U26283 (N_26283,N_11000,N_12641);
nor U26284 (N_26284,N_13712,N_10759);
and U26285 (N_26285,N_13726,N_13522);
nor U26286 (N_26286,N_14366,N_12252);
nand U26287 (N_26287,N_12586,N_11228);
or U26288 (N_26288,N_19796,N_13152);
and U26289 (N_26289,N_15222,N_18282);
nand U26290 (N_26290,N_12738,N_11404);
xnor U26291 (N_26291,N_15457,N_14932);
or U26292 (N_26292,N_19111,N_11680);
nand U26293 (N_26293,N_15014,N_17522);
and U26294 (N_26294,N_15285,N_14039);
xor U26295 (N_26295,N_13113,N_18022);
nor U26296 (N_26296,N_15191,N_12586);
and U26297 (N_26297,N_14362,N_16758);
xnor U26298 (N_26298,N_19158,N_18175);
or U26299 (N_26299,N_19236,N_14755);
nand U26300 (N_26300,N_15124,N_18619);
nor U26301 (N_26301,N_14533,N_12102);
and U26302 (N_26302,N_11487,N_14625);
nand U26303 (N_26303,N_15021,N_16637);
nor U26304 (N_26304,N_14238,N_10673);
nor U26305 (N_26305,N_16683,N_14599);
and U26306 (N_26306,N_12056,N_17866);
nand U26307 (N_26307,N_13932,N_19994);
or U26308 (N_26308,N_18861,N_13068);
nand U26309 (N_26309,N_19754,N_18261);
nor U26310 (N_26310,N_16479,N_10427);
xor U26311 (N_26311,N_17109,N_11632);
nand U26312 (N_26312,N_16461,N_17339);
xnor U26313 (N_26313,N_17911,N_10239);
nand U26314 (N_26314,N_19870,N_11924);
and U26315 (N_26315,N_12290,N_17629);
and U26316 (N_26316,N_13716,N_10722);
nor U26317 (N_26317,N_11615,N_19355);
xnor U26318 (N_26318,N_10773,N_14114);
and U26319 (N_26319,N_15944,N_17000);
and U26320 (N_26320,N_19439,N_17445);
and U26321 (N_26321,N_19167,N_16084);
xnor U26322 (N_26322,N_13665,N_15780);
and U26323 (N_26323,N_14979,N_15440);
xnor U26324 (N_26324,N_13304,N_18985);
and U26325 (N_26325,N_18403,N_14110);
xnor U26326 (N_26326,N_17443,N_13036);
xor U26327 (N_26327,N_14245,N_15241);
or U26328 (N_26328,N_18013,N_15226);
and U26329 (N_26329,N_17359,N_14735);
xor U26330 (N_26330,N_16664,N_12177);
and U26331 (N_26331,N_14019,N_13898);
and U26332 (N_26332,N_11943,N_18146);
xor U26333 (N_26333,N_16287,N_18211);
or U26334 (N_26334,N_17742,N_10134);
nand U26335 (N_26335,N_18702,N_19754);
nand U26336 (N_26336,N_13541,N_19243);
nand U26337 (N_26337,N_13611,N_16605);
or U26338 (N_26338,N_15245,N_10421);
and U26339 (N_26339,N_12734,N_13971);
and U26340 (N_26340,N_15374,N_11089);
xnor U26341 (N_26341,N_11466,N_11391);
xnor U26342 (N_26342,N_15910,N_16379);
nand U26343 (N_26343,N_17565,N_18382);
and U26344 (N_26344,N_12982,N_14119);
and U26345 (N_26345,N_11073,N_13087);
and U26346 (N_26346,N_10315,N_19591);
nor U26347 (N_26347,N_15928,N_16773);
nor U26348 (N_26348,N_19405,N_19025);
nand U26349 (N_26349,N_15233,N_18107);
xnor U26350 (N_26350,N_18311,N_13777);
or U26351 (N_26351,N_15525,N_11914);
nand U26352 (N_26352,N_12055,N_14161);
nand U26353 (N_26353,N_16323,N_14905);
and U26354 (N_26354,N_15549,N_13778);
or U26355 (N_26355,N_15322,N_10032);
nor U26356 (N_26356,N_14829,N_15951);
or U26357 (N_26357,N_11138,N_14545);
or U26358 (N_26358,N_14246,N_14569);
and U26359 (N_26359,N_19343,N_16053);
nor U26360 (N_26360,N_13696,N_17374);
or U26361 (N_26361,N_14710,N_15348);
or U26362 (N_26362,N_17812,N_15245);
nor U26363 (N_26363,N_15951,N_18899);
xnor U26364 (N_26364,N_13270,N_16779);
nor U26365 (N_26365,N_10189,N_16275);
or U26366 (N_26366,N_10262,N_16222);
nand U26367 (N_26367,N_19443,N_18542);
and U26368 (N_26368,N_12619,N_13052);
or U26369 (N_26369,N_16710,N_13115);
or U26370 (N_26370,N_13571,N_14290);
or U26371 (N_26371,N_15690,N_12460);
and U26372 (N_26372,N_13304,N_14030);
and U26373 (N_26373,N_17281,N_11331);
nor U26374 (N_26374,N_12276,N_11586);
xnor U26375 (N_26375,N_10609,N_12958);
xnor U26376 (N_26376,N_17624,N_15304);
xor U26377 (N_26377,N_18629,N_17057);
and U26378 (N_26378,N_13438,N_18933);
xor U26379 (N_26379,N_18636,N_14025);
nor U26380 (N_26380,N_18938,N_16564);
xnor U26381 (N_26381,N_10848,N_10816);
and U26382 (N_26382,N_12406,N_19560);
nor U26383 (N_26383,N_14316,N_16114);
or U26384 (N_26384,N_18475,N_16662);
xnor U26385 (N_26385,N_10574,N_17790);
xor U26386 (N_26386,N_13505,N_11236);
xor U26387 (N_26387,N_16776,N_15974);
xor U26388 (N_26388,N_10427,N_10306);
xor U26389 (N_26389,N_17766,N_17629);
or U26390 (N_26390,N_19286,N_16002);
xnor U26391 (N_26391,N_17367,N_19206);
nor U26392 (N_26392,N_16423,N_11533);
or U26393 (N_26393,N_10089,N_12460);
or U26394 (N_26394,N_14679,N_19393);
xnor U26395 (N_26395,N_12197,N_13430);
xor U26396 (N_26396,N_19749,N_16563);
nand U26397 (N_26397,N_11468,N_10230);
xor U26398 (N_26398,N_16750,N_10441);
nor U26399 (N_26399,N_19476,N_19659);
nand U26400 (N_26400,N_17358,N_13632);
or U26401 (N_26401,N_10190,N_13279);
nand U26402 (N_26402,N_15807,N_14014);
xnor U26403 (N_26403,N_15416,N_18068);
and U26404 (N_26404,N_15789,N_13255);
or U26405 (N_26405,N_12001,N_10738);
and U26406 (N_26406,N_15275,N_16129);
nand U26407 (N_26407,N_16782,N_18870);
nor U26408 (N_26408,N_12536,N_14847);
and U26409 (N_26409,N_17918,N_14189);
nand U26410 (N_26410,N_18493,N_15077);
and U26411 (N_26411,N_13427,N_13462);
nand U26412 (N_26412,N_13172,N_15128);
or U26413 (N_26413,N_12353,N_10330);
nor U26414 (N_26414,N_13729,N_16504);
and U26415 (N_26415,N_11178,N_13359);
or U26416 (N_26416,N_19128,N_18321);
or U26417 (N_26417,N_18551,N_16778);
and U26418 (N_26418,N_18690,N_10575);
nand U26419 (N_26419,N_17168,N_10821);
xor U26420 (N_26420,N_18329,N_10888);
and U26421 (N_26421,N_14928,N_10842);
or U26422 (N_26422,N_11822,N_13619);
xnor U26423 (N_26423,N_14594,N_15718);
nand U26424 (N_26424,N_10642,N_18818);
or U26425 (N_26425,N_10982,N_14836);
or U26426 (N_26426,N_15014,N_13888);
nand U26427 (N_26427,N_19107,N_14287);
and U26428 (N_26428,N_13332,N_12382);
nor U26429 (N_26429,N_17073,N_19008);
nand U26430 (N_26430,N_10580,N_18754);
and U26431 (N_26431,N_18679,N_10923);
nand U26432 (N_26432,N_11599,N_19632);
and U26433 (N_26433,N_18375,N_11496);
nor U26434 (N_26434,N_15074,N_14988);
nor U26435 (N_26435,N_18047,N_14547);
nor U26436 (N_26436,N_15050,N_14132);
nand U26437 (N_26437,N_11289,N_14380);
nand U26438 (N_26438,N_16416,N_17930);
or U26439 (N_26439,N_15295,N_14108);
nor U26440 (N_26440,N_19013,N_18882);
or U26441 (N_26441,N_13558,N_17966);
nor U26442 (N_26442,N_19125,N_16830);
nand U26443 (N_26443,N_11798,N_12311);
and U26444 (N_26444,N_14908,N_17915);
xnor U26445 (N_26445,N_13659,N_11882);
and U26446 (N_26446,N_18608,N_17366);
or U26447 (N_26447,N_15439,N_16002);
and U26448 (N_26448,N_12508,N_11766);
xnor U26449 (N_26449,N_14025,N_13289);
xnor U26450 (N_26450,N_17918,N_12423);
and U26451 (N_26451,N_18430,N_19283);
xor U26452 (N_26452,N_17917,N_17194);
and U26453 (N_26453,N_16946,N_15355);
nand U26454 (N_26454,N_18548,N_10731);
nor U26455 (N_26455,N_18926,N_12962);
nor U26456 (N_26456,N_11655,N_12505);
nor U26457 (N_26457,N_16933,N_15972);
or U26458 (N_26458,N_15657,N_12139);
or U26459 (N_26459,N_19820,N_10331);
or U26460 (N_26460,N_15794,N_19932);
nand U26461 (N_26461,N_13885,N_19267);
nand U26462 (N_26462,N_16303,N_17903);
nor U26463 (N_26463,N_12831,N_11688);
and U26464 (N_26464,N_15225,N_12416);
xor U26465 (N_26465,N_16772,N_13002);
and U26466 (N_26466,N_16733,N_19837);
xnor U26467 (N_26467,N_13101,N_11751);
nor U26468 (N_26468,N_18327,N_16348);
and U26469 (N_26469,N_16380,N_12273);
nand U26470 (N_26470,N_12208,N_14619);
nor U26471 (N_26471,N_11731,N_15168);
xnor U26472 (N_26472,N_16337,N_13664);
nor U26473 (N_26473,N_18790,N_13247);
nand U26474 (N_26474,N_12607,N_16456);
or U26475 (N_26475,N_10720,N_12010);
xnor U26476 (N_26476,N_17272,N_11860);
xor U26477 (N_26477,N_18704,N_16259);
xor U26478 (N_26478,N_16734,N_18343);
xor U26479 (N_26479,N_18361,N_11748);
xnor U26480 (N_26480,N_12868,N_19128);
nor U26481 (N_26481,N_13680,N_17781);
or U26482 (N_26482,N_17137,N_12681);
xnor U26483 (N_26483,N_11300,N_14811);
nor U26484 (N_26484,N_19535,N_16752);
or U26485 (N_26485,N_14387,N_12819);
xnor U26486 (N_26486,N_17658,N_14762);
or U26487 (N_26487,N_12944,N_12357);
nor U26488 (N_26488,N_15085,N_18570);
and U26489 (N_26489,N_13513,N_13037);
or U26490 (N_26490,N_17133,N_14813);
xnor U26491 (N_26491,N_16216,N_16127);
xor U26492 (N_26492,N_19532,N_12196);
nand U26493 (N_26493,N_12353,N_10240);
xnor U26494 (N_26494,N_10386,N_15884);
nor U26495 (N_26495,N_17324,N_12135);
or U26496 (N_26496,N_11834,N_15897);
and U26497 (N_26497,N_16917,N_17593);
nor U26498 (N_26498,N_14786,N_15617);
nand U26499 (N_26499,N_18740,N_15051);
or U26500 (N_26500,N_18084,N_12506);
nand U26501 (N_26501,N_16995,N_13555);
or U26502 (N_26502,N_16118,N_11678);
or U26503 (N_26503,N_19452,N_17293);
and U26504 (N_26504,N_10593,N_16978);
xnor U26505 (N_26505,N_19655,N_13791);
or U26506 (N_26506,N_17526,N_18266);
xor U26507 (N_26507,N_17346,N_16927);
nand U26508 (N_26508,N_15963,N_16861);
and U26509 (N_26509,N_11267,N_17697);
nor U26510 (N_26510,N_18955,N_15196);
xnor U26511 (N_26511,N_16798,N_10085);
nand U26512 (N_26512,N_14003,N_12698);
nor U26513 (N_26513,N_18142,N_11508);
xor U26514 (N_26514,N_17030,N_18109);
nor U26515 (N_26515,N_10959,N_16330);
xnor U26516 (N_26516,N_16203,N_10196);
and U26517 (N_26517,N_15654,N_12581);
and U26518 (N_26518,N_18792,N_13148);
or U26519 (N_26519,N_18330,N_12046);
and U26520 (N_26520,N_14117,N_15643);
nand U26521 (N_26521,N_19796,N_15490);
nand U26522 (N_26522,N_17499,N_14740);
nor U26523 (N_26523,N_16457,N_18778);
and U26524 (N_26524,N_19438,N_10415);
nor U26525 (N_26525,N_10108,N_12457);
and U26526 (N_26526,N_17538,N_18532);
nand U26527 (N_26527,N_16334,N_14171);
xnor U26528 (N_26528,N_10773,N_11104);
xor U26529 (N_26529,N_10801,N_17784);
xnor U26530 (N_26530,N_17144,N_10447);
xor U26531 (N_26531,N_18926,N_13406);
or U26532 (N_26532,N_13336,N_11467);
or U26533 (N_26533,N_19059,N_13942);
or U26534 (N_26534,N_19332,N_13468);
nor U26535 (N_26535,N_10761,N_19163);
nand U26536 (N_26536,N_10697,N_11577);
nand U26537 (N_26537,N_10275,N_18383);
xnor U26538 (N_26538,N_13662,N_13158);
nor U26539 (N_26539,N_18968,N_15391);
or U26540 (N_26540,N_16181,N_10730);
nor U26541 (N_26541,N_16133,N_16278);
nor U26542 (N_26542,N_17272,N_14773);
xnor U26543 (N_26543,N_13416,N_18655);
nand U26544 (N_26544,N_15727,N_17199);
nand U26545 (N_26545,N_19314,N_14502);
nand U26546 (N_26546,N_17473,N_16982);
nor U26547 (N_26547,N_17108,N_13135);
nor U26548 (N_26548,N_11494,N_13255);
and U26549 (N_26549,N_11256,N_10178);
xor U26550 (N_26550,N_12094,N_17205);
nor U26551 (N_26551,N_10565,N_11781);
or U26552 (N_26552,N_16901,N_19302);
nor U26553 (N_26553,N_17841,N_15558);
nand U26554 (N_26554,N_19754,N_12701);
or U26555 (N_26555,N_18546,N_13723);
xor U26556 (N_26556,N_18813,N_10733);
or U26557 (N_26557,N_16815,N_10672);
and U26558 (N_26558,N_13505,N_12240);
and U26559 (N_26559,N_11033,N_18388);
nand U26560 (N_26560,N_19117,N_14797);
xor U26561 (N_26561,N_18453,N_11206);
xnor U26562 (N_26562,N_13198,N_10835);
and U26563 (N_26563,N_18620,N_14732);
nor U26564 (N_26564,N_14502,N_14217);
and U26565 (N_26565,N_13689,N_18864);
nand U26566 (N_26566,N_13373,N_11783);
xor U26567 (N_26567,N_18052,N_18037);
xor U26568 (N_26568,N_13466,N_11822);
nand U26569 (N_26569,N_12772,N_18223);
nand U26570 (N_26570,N_16615,N_18380);
and U26571 (N_26571,N_16817,N_10774);
nand U26572 (N_26572,N_14444,N_18764);
nor U26573 (N_26573,N_19007,N_19530);
or U26574 (N_26574,N_18664,N_18508);
and U26575 (N_26575,N_12385,N_17965);
xor U26576 (N_26576,N_13982,N_13699);
and U26577 (N_26577,N_15612,N_11378);
and U26578 (N_26578,N_18137,N_14934);
xnor U26579 (N_26579,N_10139,N_19146);
or U26580 (N_26580,N_19403,N_19672);
nor U26581 (N_26581,N_12565,N_12312);
xnor U26582 (N_26582,N_13877,N_16165);
nand U26583 (N_26583,N_17030,N_13978);
xnor U26584 (N_26584,N_10019,N_15468);
xor U26585 (N_26585,N_18734,N_16813);
nor U26586 (N_26586,N_10928,N_14469);
nand U26587 (N_26587,N_12421,N_11879);
xor U26588 (N_26588,N_15614,N_16171);
nand U26589 (N_26589,N_18544,N_18551);
or U26590 (N_26590,N_16496,N_15802);
nand U26591 (N_26591,N_11852,N_17323);
xnor U26592 (N_26592,N_14179,N_18934);
nand U26593 (N_26593,N_16624,N_16218);
or U26594 (N_26594,N_15760,N_17119);
nand U26595 (N_26595,N_10371,N_14693);
nor U26596 (N_26596,N_16801,N_16954);
and U26597 (N_26597,N_17527,N_15623);
nor U26598 (N_26598,N_13481,N_17537);
or U26599 (N_26599,N_19018,N_16737);
nor U26600 (N_26600,N_12786,N_12592);
xor U26601 (N_26601,N_10756,N_19442);
or U26602 (N_26602,N_17546,N_14365);
or U26603 (N_26603,N_13361,N_13355);
or U26604 (N_26604,N_12649,N_14977);
xor U26605 (N_26605,N_17255,N_19978);
nor U26606 (N_26606,N_12296,N_12991);
nand U26607 (N_26607,N_12657,N_18537);
xor U26608 (N_26608,N_16667,N_15488);
nand U26609 (N_26609,N_18648,N_13279);
nand U26610 (N_26610,N_16017,N_17116);
xor U26611 (N_26611,N_11438,N_17896);
and U26612 (N_26612,N_11143,N_13990);
and U26613 (N_26613,N_18037,N_17256);
nor U26614 (N_26614,N_13706,N_15790);
nand U26615 (N_26615,N_17338,N_18404);
nand U26616 (N_26616,N_18946,N_19546);
xor U26617 (N_26617,N_15285,N_10019);
or U26618 (N_26618,N_18810,N_12631);
and U26619 (N_26619,N_18534,N_15135);
or U26620 (N_26620,N_19556,N_14845);
nand U26621 (N_26621,N_16647,N_15846);
xor U26622 (N_26622,N_11981,N_18213);
or U26623 (N_26623,N_11371,N_18608);
nand U26624 (N_26624,N_17832,N_13096);
and U26625 (N_26625,N_14320,N_19754);
nand U26626 (N_26626,N_18234,N_12151);
and U26627 (N_26627,N_16898,N_14026);
or U26628 (N_26628,N_13331,N_19162);
xor U26629 (N_26629,N_10379,N_15154);
nor U26630 (N_26630,N_18811,N_15165);
nor U26631 (N_26631,N_14576,N_10094);
and U26632 (N_26632,N_12598,N_16670);
xnor U26633 (N_26633,N_11319,N_19142);
xor U26634 (N_26634,N_18290,N_14664);
nand U26635 (N_26635,N_16879,N_10390);
nor U26636 (N_26636,N_17801,N_11196);
xor U26637 (N_26637,N_12549,N_13286);
nand U26638 (N_26638,N_14027,N_13886);
and U26639 (N_26639,N_16579,N_10337);
or U26640 (N_26640,N_13526,N_16335);
xnor U26641 (N_26641,N_14532,N_14680);
or U26642 (N_26642,N_11411,N_12596);
nand U26643 (N_26643,N_12673,N_10352);
nor U26644 (N_26644,N_12470,N_16313);
and U26645 (N_26645,N_15788,N_14964);
nand U26646 (N_26646,N_10276,N_18331);
nor U26647 (N_26647,N_12851,N_15518);
and U26648 (N_26648,N_15073,N_10938);
and U26649 (N_26649,N_10795,N_16724);
xor U26650 (N_26650,N_10396,N_17374);
or U26651 (N_26651,N_10205,N_17137);
or U26652 (N_26652,N_16390,N_12352);
or U26653 (N_26653,N_15700,N_14542);
nor U26654 (N_26654,N_19435,N_17207);
nor U26655 (N_26655,N_15652,N_15606);
and U26656 (N_26656,N_19846,N_15028);
nand U26657 (N_26657,N_17530,N_17544);
xnor U26658 (N_26658,N_11421,N_12143);
xor U26659 (N_26659,N_19064,N_12911);
or U26660 (N_26660,N_11639,N_12397);
xor U26661 (N_26661,N_18179,N_14196);
nor U26662 (N_26662,N_15885,N_11909);
nand U26663 (N_26663,N_15073,N_11377);
or U26664 (N_26664,N_15962,N_14732);
nor U26665 (N_26665,N_18555,N_16683);
and U26666 (N_26666,N_19286,N_18988);
nand U26667 (N_26667,N_11240,N_16365);
or U26668 (N_26668,N_15631,N_14082);
xnor U26669 (N_26669,N_18958,N_16310);
and U26670 (N_26670,N_14392,N_14079);
and U26671 (N_26671,N_10829,N_14730);
xnor U26672 (N_26672,N_16995,N_14387);
and U26673 (N_26673,N_10197,N_10480);
xor U26674 (N_26674,N_13451,N_16513);
xor U26675 (N_26675,N_14300,N_15329);
xnor U26676 (N_26676,N_19452,N_14640);
or U26677 (N_26677,N_15703,N_11421);
or U26678 (N_26678,N_15432,N_10800);
and U26679 (N_26679,N_13301,N_19732);
and U26680 (N_26680,N_18836,N_17382);
xnor U26681 (N_26681,N_10198,N_19847);
xor U26682 (N_26682,N_19105,N_16496);
nand U26683 (N_26683,N_11257,N_19025);
or U26684 (N_26684,N_11473,N_15599);
nand U26685 (N_26685,N_19165,N_15139);
or U26686 (N_26686,N_10854,N_13526);
nand U26687 (N_26687,N_13426,N_16689);
xnor U26688 (N_26688,N_17109,N_15268);
and U26689 (N_26689,N_17525,N_12088);
and U26690 (N_26690,N_16774,N_14361);
and U26691 (N_26691,N_16060,N_19740);
xnor U26692 (N_26692,N_13798,N_15958);
or U26693 (N_26693,N_10097,N_15443);
xnor U26694 (N_26694,N_15234,N_14685);
or U26695 (N_26695,N_16209,N_10414);
nand U26696 (N_26696,N_12935,N_14279);
or U26697 (N_26697,N_19990,N_19744);
nor U26698 (N_26698,N_19034,N_17408);
nand U26699 (N_26699,N_14233,N_10424);
and U26700 (N_26700,N_13254,N_12269);
nand U26701 (N_26701,N_13432,N_10066);
and U26702 (N_26702,N_12889,N_17843);
nor U26703 (N_26703,N_11625,N_16891);
nand U26704 (N_26704,N_15746,N_14967);
nand U26705 (N_26705,N_13082,N_15633);
xor U26706 (N_26706,N_15573,N_12709);
and U26707 (N_26707,N_13563,N_16755);
xnor U26708 (N_26708,N_16171,N_14868);
or U26709 (N_26709,N_13865,N_19708);
nor U26710 (N_26710,N_13922,N_12751);
nor U26711 (N_26711,N_19688,N_19606);
nand U26712 (N_26712,N_15668,N_13403);
or U26713 (N_26713,N_15417,N_18378);
and U26714 (N_26714,N_14640,N_14024);
xor U26715 (N_26715,N_14781,N_11800);
and U26716 (N_26716,N_12175,N_15996);
or U26717 (N_26717,N_19460,N_14088);
nor U26718 (N_26718,N_16957,N_12267);
or U26719 (N_26719,N_19902,N_15107);
or U26720 (N_26720,N_14820,N_14113);
xor U26721 (N_26721,N_15235,N_19178);
and U26722 (N_26722,N_17683,N_17876);
nor U26723 (N_26723,N_19553,N_13526);
or U26724 (N_26724,N_14502,N_11639);
xor U26725 (N_26725,N_19787,N_17353);
nor U26726 (N_26726,N_12282,N_12462);
nor U26727 (N_26727,N_17378,N_17755);
nand U26728 (N_26728,N_13944,N_16702);
or U26729 (N_26729,N_10769,N_13709);
and U26730 (N_26730,N_18999,N_12381);
or U26731 (N_26731,N_14786,N_11648);
nor U26732 (N_26732,N_17624,N_11763);
nor U26733 (N_26733,N_10450,N_14466);
and U26734 (N_26734,N_12113,N_18873);
nor U26735 (N_26735,N_11534,N_19909);
nand U26736 (N_26736,N_18477,N_16733);
nor U26737 (N_26737,N_14231,N_13298);
and U26738 (N_26738,N_19343,N_16642);
xnor U26739 (N_26739,N_17562,N_14989);
nor U26740 (N_26740,N_13040,N_12174);
and U26741 (N_26741,N_15762,N_15855);
nand U26742 (N_26742,N_13104,N_12905);
or U26743 (N_26743,N_15159,N_11270);
xnor U26744 (N_26744,N_16906,N_19802);
and U26745 (N_26745,N_15237,N_13955);
nor U26746 (N_26746,N_17329,N_13980);
or U26747 (N_26747,N_12450,N_19366);
xnor U26748 (N_26748,N_12619,N_10786);
nand U26749 (N_26749,N_19175,N_19543);
nor U26750 (N_26750,N_18840,N_19478);
nor U26751 (N_26751,N_12035,N_17184);
nor U26752 (N_26752,N_19385,N_11691);
xnor U26753 (N_26753,N_15012,N_12155);
nor U26754 (N_26754,N_11205,N_12437);
xor U26755 (N_26755,N_14285,N_14106);
nor U26756 (N_26756,N_16054,N_13512);
or U26757 (N_26757,N_18689,N_12144);
nor U26758 (N_26758,N_17091,N_10397);
nand U26759 (N_26759,N_12075,N_12143);
or U26760 (N_26760,N_15155,N_13679);
and U26761 (N_26761,N_10848,N_15326);
and U26762 (N_26762,N_13464,N_18870);
nor U26763 (N_26763,N_16441,N_13674);
nand U26764 (N_26764,N_12332,N_12621);
or U26765 (N_26765,N_15962,N_15533);
xor U26766 (N_26766,N_16156,N_10077);
nand U26767 (N_26767,N_19020,N_15110);
and U26768 (N_26768,N_14013,N_10671);
xnor U26769 (N_26769,N_15247,N_10319);
xnor U26770 (N_26770,N_16344,N_17890);
or U26771 (N_26771,N_19724,N_13193);
or U26772 (N_26772,N_18823,N_16063);
or U26773 (N_26773,N_16368,N_16143);
nand U26774 (N_26774,N_18416,N_12741);
or U26775 (N_26775,N_16465,N_18078);
nor U26776 (N_26776,N_13047,N_16467);
nor U26777 (N_26777,N_14201,N_10467);
nor U26778 (N_26778,N_13266,N_10852);
nor U26779 (N_26779,N_16287,N_15560);
nor U26780 (N_26780,N_14212,N_11652);
or U26781 (N_26781,N_12144,N_15473);
or U26782 (N_26782,N_11318,N_16382);
xor U26783 (N_26783,N_11688,N_18020);
or U26784 (N_26784,N_18266,N_10080);
nor U26785 (N_26785,N_18069,N_13788);
nand U26786 (N_26786,N_11198,N_10651);
xnor U26787 (N_26787,N_17104,N_19278);
or U26788 (N_26788,N_15221,N_18955);
xnor U26789 (N_26789,N_13549,N_11515);
and U26790 (N_26790,N_16864,N_19862);
nor U26791 (N_26791,N_12508,N_12628);
nor U26792 (N_26792,N_18160,N_18428);
nand U26793 (N_26793,N_13579,N_19746);
nand U26794 (N_26794,N_12769,N_16122);
nand U26795 (N_26795,N_17737,N_14123);
xor U26796 (N_26796,N_11160,N_16805);
xor U26797 (N_26797,N_13340,N_16492);
or U26798 (N_26798,N_12238,N_12929);
xnor U26799 (N_26799,N_11137,N_15068);
xor U26800 (N_26800,N_19244,N_16488);
nand U26801 (N_26801,N_16911,N_12443);
xnor U26802 (N_26802,N_10397,N_13790);
and U26803 (N_26803,N_13048,N_18921);
nand U26804 (N_26804,N_17746,N_11987);
nand U26805 (N_26805,N_18631,N_16550);
xnor U26806 (N_26806,N_13692,N_18369);
or U26807 (N_26807,N_17866,N_11927);
xor U26808 (N_26808,N_17162,N_18466);
nand U26809 (N_26809,N_17667,N_17145);
nor U26810 (N_26810,N_12704,N_16449);
or U26811 (N_26811,N_17982,N_19639);
and U26812 (N_26812,N_11482,N_18630);
nor U26813 (N_26813,N_19123,N_14439);
nor U26814 (N_26814,N_15839,N_11348);
or U26815 (N_26815,N_19575,N_16804);
xnor U26816 (N_26816,N_10641,N_16216);
and U26817 (N_26817,N_12688,N_19976);
and U26818 (N_26818,N_15818,N_19735);
or U26819 (N_26819,N_15747,N_18794);
xnor U26820 (N_26820,N_14472,N_18555);
or U26821 (N_26821,N_18326,N_10599);
and U26822 (N_26822,N_10608,N_18016);
xnor U26823 (N_26823,N_13133,N_15558);
or U26824 (N_26824,N_16491,N_13284);
or U26825 (N_26825,N_17562,N_16072);
nor U26826 (N_26826,N_11882,N_13901);
and U26827 (N_26827,N_12755,N_14808);
and U26828 (N_26828,N_15492,N_16159);
nand U26829 (N_26829,N_17815,N_10608);
and U26830 (N_26830,N_10184,N_16919);
and U26831 (N_26831,N_12435,N_16284);
or U26832 (N_26832,N_19422,N_10403);
xor U26833 (N_26833,N_11676,N_15903);
and U26834 (N_26834,N_10179,N_15552);
and U26835 (N_26835,N_18894,N_17463);
xnor U26836 (N_26836,N_10479,N_14244);
nor U26837 (N_26837,N_13572,N_11693);
and U26838 (N_26838,N_15079,N_11853);
or U26839 (N_26839,N_16009,N_14505);
and U26840 (N_26840,N_15813,N_16172);
nor U26841 (N_26841,N_14494,N_19522);
nor U26842 (N_26842,N_12750,N_10289);
nor U26843 (N_26843,N_19731,N_13051);
and U26844 (N_26844,N_11410,N_14798);
nand U26845 (N_26845,N_19036,N_16389);
or U26846 (N_26846,N_14409,N_15592);
xnor U26847 (N_26847,N_14364,N_16463);
or U26848 (N_26848,N_19599,N_18044);
nand U26849 (N_26849,N_14578,N_15698);
and U26850 (N_26850,N_12693,N_11778);
nor U26851 (N_26851,N_14422,N_15884);
xor U26852 (N_26852,N_10110,N_17796);
xnor U26853 (N_26853,N_18314,N_14836);
or U26854 (N_26854,N_17112,N_12265);
or U26855 (N_26855,N_15157,N_16407);
and U26856 (N_26856,N_12857,N_18213);
and U26857 (N_26857,N_15314,N_17182);
xnor U26858 (N_26858,N_16711,N_19994);
nor U26859 (N_26859,N_16289,N_19371);
or U26860 (N_26860,N_17778,N_10253);
nor U26861 (N_26861,N_19352,N_12397);
or U26862 (N_26862,N_17162,N_12024);
or U26863 (N_26863,N_12349,N_15231);
xor U26864 (N_26864,N_10808,N_17504);
nand U26865 (N_26865,N_19620,N_10508);
nand U26866 (N_26866,N_19051,N_10528);
nor U26867 (N_26867,N_18035,N_12492);
or U26868 (N_26868,N_16320,N_14565);
nand U26869 (N_26869,N_18747,N_11753);
nor U26870 (N_26870,N_19497,N_18622);
or U26871 (N_26871,N_15399,N_19136);
nand U26872 (N_26872,N_18135,N_15059);
xor U26873 (N_26873,N_15378,N_19703);
or U26874 (N_26874,N_15487,N_11002);
nor U26875 (N_26875,N_10838,N_13472);
or U26876 (N_26876,N_18729,N_19091);
xor U26877 (N_26877,N_16834,N_17808);
and U26878 (N_26878,N_16944,N_16283);
nand U26879 (N_26879,N_11173,N_13036);
nand U26880 (N_26880,N_12002,N_10080);
or U26881 (N_26881,N_17078,N_16684);
or U26882 (N_26882,N_18301,N_10831);
xor U26883 (N_26883,N_16091,N_16148);
or U26884 (N_26884,N_12303,N_19738);
and U26885 (N_26885,N_19677,N_14322);
xnor U26886 (N_26886,N_17478,N_18988);
or U26887 (N_26887,N_18998,N_16785);
nor U26888 (N_26888,N_13131,N_14487);
and U26889 (N_26889,N_11448,N_11477);
nor U26890 (N_26890,N_13454,N_10359);
or U26891 (N_26891,N_10013,N_16291);
nand U26892 (N_26892,N_12066,N_19597);
xnor U26893 (N_26893,N_13092,N_17983);
nand U26894 (N_26894,N_16490,N_11547);
or U26895 (N_26895,N_18399,N_18277);
nand U26896 (N_26896,N_11215,N_11756);
nand U26897 (N_26897,N_12660,N_14283);
xnor U26898 (N_26898,N_19401,N_11152);
or U26899 (N_26899,N_16590,N_16638);
nand U26900 (N_26900,N_10929,N_14074);
nand U26901 (N_26901,N_18319,N_14958);
nor U26902 (N_26902,N_12081,N_14554);
nor U26903 (N_26903,N_17931,N_14142);
nor U26904 (N_26904,N_11597,N_14934);
nand U26905 (N_26905,N_10995,N_18611);
and U26906 (N_26906,N_11661,N_15246);
and U26907 (N_26907,N_16764,N_17404);
xor U26908 (N_26908,N_17040,N_11467);
and U26909 (N_26909,N_13432,N_12750);
nand U26910 (N_26910,N_11460,N_12861);
or U26911 (N_26911,N_12173,N_11568);
or U26912 (N_26912,N_11747,N_11398);
xnor U26913 (N_26913,N_19889,N_16862);
nand U26914 (N_26914,N_19354,N_11330);
or U26915 (N_26915,N_15524,N_18063);
and U26916 (N_26916,N_15454,N_13293);
nand U26917 (N_26917,N_10703,N_13657);
nor U26918 (N_26918,N_12658,N_15768);
nor U26919 (N_26919,N_13003,N_17917);
xnor U26920 (N_26920,N_17609,N_19133);
nand U26921 (N_26921,N_17828,N_14112);
and U26922 (N_26922,N_19754,N_12866);
or U26923 (N_26923,N_10626,N_11345);
xor U26924 (N_26924,N_15434,N_10432);
xnor U26925 (N_26925,N_11065,N_13388);
nor U26926 (N_26926,N_19528,N_10707);
or U26927 (N_26927,N_12623,N_12367);
nor U26928 (N_26928,N_15061,N_12673);
or U26929 (N_26929,N_13931,N_16879);
nor U26930 (N_26930,N_12067,N_13271);
and U26931 (N_26931,N_15134,N_19193);
or U26932 (N_26932,N_19326,N_17412);
nor U26933 (N_26933,N_12895,N_16236);
nor U26934 (N_26934,N_18895,N_19952);
nand U26935 (N_26935,N_18557,N_17454);
or U26936 (N_26936,N_19755,N_15551);
nor U26937 (N_26937,N_17406,N_12597);
and U26938 (N_26938,N_13912,N_16372);
xor U26939 (N_26939,N_16897,N_11177);
and U26940 (N_26940,N_16617,N_16432);
xor U26941 (N_26941,N_10030,N_14041);
nor U26942 (N_26942,N_11603,N_10824);
and U26943 (N_26943,N_11362,N_10852);
xnor U26944 (N_26944,N_16326,N_17262);
nor U26945 (N_26945,N_11206,N_14185);
and U26946 (N_26946,N_14689,N_14473);
and U26947 (N_26947,N_19740,N_17344);
or U26948 (N_26948,N_13235,N_18964);
nor U26949 (N_26949,N_16442,N_14655);
xnor U26950 (N_26950,N_16982,N_11208);
nand U26951 (N_26951,N_16800,N_16638);
nand U26952 (N_26952,N_19088,N_14097);
or U26953 (N_26953,N_11732,N_11993);
and U26954 (N_26954,N_17920,N_14885);
nand U26955 (N_26955,N_19373,N_19688);
nand U26956 (N_26956,N_11035,N_10354);
nand U26957 (N_26957,N_15876,N_15327);
or U26958 (N_26958,N_12174,N_18615);
nand U26959 (N_26959,N_12864,N_10897);
nand U26960 (N_26960,N_11075,N_16446);
nor U26961 (N_26961,N_19465,N_15077);
xor U26962 (N_26962,N_14646,N_10513);
and U26963 (N_26963,N_13199,N_14597);
xnor U26964 (N_26964,N_14890,N_14307);
and U26965 (N_26965,N_15710,N_15650);
nor U26966 (N_26966,N_16433,N_10661);
and U26967 (N_26967,N_16982,N_18508);
or U26968 (N_26968,N_16505,N_18675);
xor U26969 (N_26969,N_14567,N_17554);
and U26970 (N_26970,N_19650,N_10389);
nor U26971 (N_26971,N_14228,N_19885);
nand U26972 (N_26972,N_16216,N_19295);
or U26973 (N_26973,N_13889,N_11466);
and U26974 (N_26974,N_14974,N_12757);
nor U26975 (N_26975,N_11211,N_12772);
or U26976 (N_26976,N_15581,N_18157);
and U26977 (N_26977,N_10287,N_10940);
and U26978 (N_26978,N_16515,N_15749);
nor U26979 (N_26979,N_11280,N_18294);
or U26980 (N_26980,N_16566,N_14849);
nand U26981 (N_26981,N_16456,N_17768);
nand U26982 (N_26982,N_18808,N_14041);
nand U26983 (N_26983,N_10905,N_15022);
nor U26984 (N_26984,N_13925,N_14601);
xnor U26985 (N_26985,N_15695,N_12677);
nand U26986 (N_26986,N_16459,N_11416);
xnor U26987 (N_26987,N_10963,N_19413);
xor U26988 (N_26988,N_12671,N_11027);
nand U26989 (N_26989,N_13544,N_15525);
and U26990 (N_26990,N_12951,N_14847);
xnor U26991 (N_26991,N_13448,N_17807);
and U26992 (N_26992,N_15021,N_10129);
nand U26993 (N_26993,N_12748,N_17785);
nor U26994 (N_26994,N_10756,N_10039);
or U26995 (N_26995,N_16739,N_13310);
and U26996 (N_26996,N_16101,N_11756);
or U26997 (N_26997,N_12198,N_11614);
or U26998 (N_26998,N_10863,N_14755);
xor U26999 (N_26999,N_16223,N_13546);
and U27000 (N_27000,N_17287,N_13468);
or U27001 (N_27001,N_12194,N_10319);
or U27002 (N_27002,N_13250,N_17035);
nand U27003 (N_27003,N_11014,N_13019);
xor U27004 (N_27004,N_16935,N_19771);
xor U27005 (N_27005,N_10810,N_14619);
and U27006 (N_27006,N_15555,N_15799);
nor U27007 (N_27007,N_10456,N_17809);
nor U27008 (N_27008,N_11219,N_11804);
or U27009 (N_27009,N_12528,N_12863);
nand U27010 (N_27010,N_19205,N_11825);
nand U27011 (N_27011,N_10459,N_13746);
nand U27012 (N_27012,N_14724,N_14100);
nor U27013 (N_27013,N_13296,N_14280);
or U27014 (N_27014,N_14375,N_15724);
xnor U27015 (N_27015,N_10356,N_11250);
nor U27016 (N_27016,N_13523,N_10967);
nand U27017 (N_27017,N_13481,N_14771);
and U27018 (N_27018,N_12184,N_19974);
nand U27019 (N_27019,N_14681,N_19421);
xnor U27020 (N_27020,N_12623,N_10762);
nor U27021 (N_27021,N_16840,N_14329);
or U27022 (N_27022,N_17900,N_19705);
xor U27023 (N_27023,N_15145,N_12731);
or U27024 (N_27024,N_18439,N_17018);
xor U27025 (N_27025,N_18382,N_13477);
xor U27026 (N_27026,N_11532,N_18223);
nor U27027 (N_27027,N_10787,N_16710);
or U27028 (N_27028,N_10496,N_18504);
nand U27029 (N_27029,N_12849,N_17663);
and U27030 (N_27030,N_16232,N_17240);
and U27031 (N_27031,N_16967,N_17557);
nor U27032 (N_27032,N_10529,N_19942);
nand U27033 (N_27033,N_16995,N_15805);
xnor U27034 (N_27034,N_19403,N_18548);
or U27035 (N_27035,N_12107,N_15977);
nand U27036 (N_27036,N_17032,N_15007);
xnor U27037 (N_27037,N_12375,N_11606);
and U27038 (N_27038,N_16866,N_10561);
xor U27039 (N_27039,N_12131,N_18861);
nor U27040 (N_27040,N_17372,N_16625);
xor U27041 (N_27041,N_10059,N_10246);
nand U27042 (N_27042,N_10440,N_16464);
or U27043 (N_27043,N_17051,N_10286);
nor U27044 (N_27044,N_10299,N_19026);
nor U27045 (N_27045,N_13493,N_11266);
xor U27046 (N_27046,N_17052,N_13850);
nand U27047 (N_27047,N_15797,N_19987);
nor U27048 (N_27048,N_11082,N_16647);
xnor U27049 (N_27049,N_16127,N_12975);
or U27050 (N_27050,N_14041,N_10822);
nand U27051 (N_27051,N_19336,N_11117);
nor U27052 (N_27052,N_19971,N_16450);
xnor U27053 (N_27053,N_19839,N_15164);
and U27054 (N_27054,N_19989,N_14526);
and U27055 (N_27055,N_13544,N_16256);
nand U27056 (N_27056,N_19968,N_11794);
nor U27057 (N_27057,N_18193,N_11223);
and U27058 (N_27058,N_19202,N_10709);
or U27059 (N_27059,N_19363,N_10018);
xnor U27060 (N_27060,N_18902,N_16591);
and U27061 (N_27061,N_10146,N_18685);
xor U27062 (N_27062,N_15268,N_17408);
and U27063 (N_27063,N_18158,N_17181);
nand U27064 (N_27064,N_19058,N_13537);
or U27065 (N_27065,N_10730,N_17049);
nor U27066 (N_27066,N_15971,N_10554);
and U27067 (N_27067,N_13387,N_19370);
nor U27068 (N_27068,N_10999,N_13606);
nand U27069 (N_27069,N_13151,N_19731);
nor U27070 (N_27070,N_13606,N_10074);
and U27071 (N_27071,N_18690,N_16367);
xor U27072 (N_27072,N_18860,N_12225);
or U27073 (N_27073,N_17519,N_11030);
nand U27074 (N_27074,N_17399,N_18220);
xnor U27075 (N_27075,N_16202,N_19265);
xor U27076 (N_27076,N_15444,N_18384);
and U27077 (N_27077,N_14601,N_15641);
nand U27078 (N_27078,N_16453,N_14435);
and U27079 (N_27079,N_14891,N_16926);
nor U27080 (N_27080,N_16457,N_17427);
or U27081 (N_27081,N_19949,N_13712);
nor U27082 (N_27082,N_17066,N_10046);
nand U27083 (N_27083,N_12173,N_11274);
nand U27084 (N_27084,N_11374,N_19998);
nand U27085 (N_27085,N_10685,N_16269);
or U27086 (N_27086,N_16901,N_14279);
and U27087 (N_27087,N_17505,N_12008);
xor U27088 (N_27088,N_10211,N_15945);
nand U27089 (N_27089,N_14914,N_19866);
xnor U27090 (N_27090,N_14122,N_11233);
and U27091 (N_27091,N_19118,N_18353);
or U27092 (N_27092,N_11252,N_17453);
or U27093 (N_27093,N_11901,N_14859);
and U27094 (N_27094,N_10689,N_15814);
xor U27095 (N_27095,N_14620,N_18714);
xnor U27096 (N_27096,N_16767,N_18679);
nand U27097 (N_27097,N_11757,N_13609);
nand U27098 (N_27098,N_17622,N_13160);
nor U27099 (N_27099,N_10548,N_16496);
and U27100 (N_27100,N_14519,N_17222);
or U27101 (N_27101,N_11076,N_11277);
nand U27102 (N_27102,N_10447,N_13078);
nor U27103 (N_27103,N_10713,N_10202);
xor U27104 (N_27104,N_16378,N_18777);
xnor U27105 (N_27105,N_16864,N_12653);
and U27106 (N_27106,N_19638,N_13682);
xnor U27107 (N_27107,N_12632,N_16720);
and U27108 (N_27108,N_18279,N_15175);
nor U27109 (N_27109,N_15453,N_10412);
xnor U27110 (N_27110,N_16544,N_15529);
xnor U27111 (N_27111,N_12554,N_14807);
or U27112 (N_27112,N_12436,N_16006);
xor U27113 (N_27113,N_16412,N_19632);
nor U27114 (N_27114,N_12510,N_11655);
and U27115 (N_27115,N_18466,N_13915);
nor U27116 (N_27116,N_14453,N_15854);
nand U27117 (N_27117,N_12293,N_15541);
and U27118 (N_27118,N_19933,N_15847);
xnor U27119 (N_27119,N_15676,N_12946);
xor U27120 (N_27120,N_17824,N_10519);
xnor U27121 (N_27121,N_14224,N_10865);
or U27122 (N_27122,N_18011,N_12370);
nor U27123 (N_27123,N_14400,N_12958);
xor U27124 (N_27124,N_16260,N_14852);
nand U27125 (N_27125,N_13104,N_15719);
and U27126 (N_27126,N_15601,N_13978);
xor U27127 (N_27127,N_11061,N_10579);
or U27128 (N_27128,N_19203,N_13921);
nor U27129 (N_27129,N_12408,N_18360);
nor U27130 (N_27130,N_14265,N_17000);
nand U27131 (N_27131,N_16155,N_12187);
nand U27132 (N_27132,N_11490,N_12321);
xnor U27133 (N_27133,N_18571,N_17165);
nand U27134 (N_27134,N_18229,N_14887);
nand U27135 (N_27135,N_12692,N_12177);
and U27136 (N_27136,N_19812,N_11603);
xnor U27137 (N_27137,N_17148,N_15991);
nand U27138 (N_27138,N_11173,N_17456);
nor U27139 (N_27139,N_14035,N_13676);
nor U27140 (N_27140,N_14740,N_16779);
nand U27141 (N_27141,N_17369,N_17957);
nand U27142 (N_27142,N_18549,N_11521);
nor U27143 (N_27143,N_19142,N_10185);
xnor U27144 (N_27144,N_14054,N_10153);
nand U27145 (N_27145,N_14834,N_13521);
and U27146 (N_27146,N_10561,N_19696);
nand U27147 (N_27147,N_17678,N_16394);
nor U27148 (N_27148,N_14042,N_16888);
xor U27149 (N_27149,N_11265,N_16374);
nor U27150 (N_27150,N_11717,N_19319);
and U27151 (N_27151,N_11417,N_10150);
nor U27152 (N_27152,N_14697,N_18005);
and U27153 (N_27153,N_10316,N_10335);
nor U27154 (N_27154,N_11500,N_18057);
nor U27155 (N_27155,N_18064,N_10034);
nand U27156 (N_27156,N_12888,N_12133);
and U27157 (N_27157,N_17599,N_18732);
or U27158 (N_27158,N_16872,N_16018);
nor U27159 (N_27159,N_12433,N_12767);
xnor U27160 (N_27160,N_13666,N_14064);
nor U27161 (N_27161,N_15396,N_16373);
or U27162 (N_27162,N_16649,N_11759);
and U27163 (N_27163,N_11622,N_11909);
nor U27164 (N_27164,N_19348,N_13845);
nor U27165 (N_27165,N_14162,N_13975);
nand U27166 (N_27166,N_18428,N_11627);
nor U27167 (N_27167,N_12043,N_11859);
and U27168 (N_27168,N_15580,N_13460);
nand U27169 (N_27169,N_15824,N_13703);
nand U27170 (N_27170,N_11007,N_19201);
nand U27171 (N_27171,N_18473,N_12007);
xor U27172 (N_27172,N_18164,N_13339);
nor U27173 (N_27173,N_12714,N_16740);
nand U27174 (N_27174,N_19364,N_12655);
nor U27175 (N_27175,N_10044,N_10905);
nor U27176 (N_27176,N_12432,N_13986);
and U27177 (N_27177,N_17556,N_18042);
xnor U27178 (N_27178,N_19048,N_10542);
xnor U27179 (N_27179,N_17754,N_12065);
nor U27180 (N_27180,N_17134,N_12665);
nor U27181 (N_27181,N_14789,N_11694);
and U27182 (N_27182,N_13563,N_11131);
xnor U27183 (N_27183,N_10475,N_10994);
nor U27184 (N_27184,N_10981,N_17312);
and U27185 (N_27185,N_14894,N_12368);
nand U27186 (N_27186,N_14610,N_13196);
or U27187 (N_27187,N_13798,N_14889);
xnor U27188 (N_27188,N_12805,N_18823);
xnor U27189 (N_27189,N_15182,N_10670);
nand U27190 (N_27190,N_19209,N_15856);
xor U27191 (N_27191,N_17270,N_10250);
and U27192 (N_27192,N_10079,N_11115);
or U27193 (N_27193,N_13486,N_13803);
and U27194 (N_27194,N_18682,N_18356);
or U27195 (N_27195,N_14623,N_16263);
and U27196 (N_27196,N_16044,N_11327);
and U27197 (N_27197,N_15252,N_10800);
and U27198 (N_27198,N_14797,N_17592);
nand U27199 (N_27199,N_19880,N_14522);
or U27200 (N_27200,N_18010,N_10105);
and U27201 (N_27201,N_18377,N_12356);
and U27202 (N_27202,N_15093,N_14958);
or U27203 (N_27203,N_14806,N_15821);
or U27204 (N_27204,N_10022,N_12550);
or U27205 (N_27205,N_10469,N_12550);
nand U27206 (N_27206,N_10961,N_15770);
xor U27207 (N_27207,N_18264,N_18105);
nor U27208 (N_27208,N_11605,N_12381);
or U27209 (N_27209,N_19403,N_11600);
xnor U27210 (N_27210,N_14001,N_14883);
or U27211 (N_27211,N_11712,N_15827);
or U27212 (N_27212,N_19633,N_17688);
nor U27213 (N_27213,N_10723,N_19513);
nand U27214 (N_27214,N_13032,N_10742);
or U27215 (N_27215,N_12406,N_17084);
nor U27216 (N_27216,N_10498,N_10104);
nand U27217 (N_27217,N_18686,N_18532);
nor U27218 (N_27218,N_15638,N_11134);
or U27219 (N_27219,N_14996,N_12099);
xor U27220 (N_27220,N_18838,N_10536);
nand U27221 (N_27221,N_12911,N_11339);
or U27222 (N_27222,N_16420,N_16322);
xnor U27223 (N_27223,N_10768,N_12630);
and U27224 (N_27224,N_19566,N_12654);
or U27225 (N_27225,N_17974,N_12335);
nand U27226 (N_27226,N_18723,N_11609);
and U27227 (N_27227,N_14327,N_16869);
nand U27228 (N_27228,N_19249,N_15890);
or U27229 (N_27229,N_16429,N_17454);
or U27230 (N_27230,N_15010,N_16834);
nand U27231 (N_27231,N_12196,N_17954);
and U27232 (N_27232,N_18379,N_14815);
and U27233 (N_27233,N_10207,N_17235);
nor U27234 (N_27234,N_14151,N_12213);
nand U27235 (N_27235,N_17863,N_12934);
and U27236 (N_27236,N_11384,N_18248);
and U27237 (N_27237,N_16117,N_14996);
nand U27238 (N_27238,N_13040,N_15059);
nor U27239 (N_27239,N_16561,N_12902);
nand U27240 (N_27240,N_13005,N_12643);
nand U27241 (N_27241,N_10522,N_13132);
nor U27242 (N_27242,N_14571,N_17935);
nor U27243 (N_27243,N_15479,N_10363);
nor U27244 (N_27244,N_17342,N_10124);
and U27245 (N_27245,N_16076,N_19365);
nand U27246 (N_27246,N_12405,N_14569);
nand U27247 (N_27247,N_15386,N_14814);
and U27248 (N_27248,N_15461,N_13491);
nor U27249 (N_27249,N_16570,N_16833);
nor U27250 (N_27250,N_15788,N_16181);
nor U27251 (N_27251,N_15192,N_19348);
xor U27252 (N_27252,N_19921,N_19517);
or U27253 (N_27253,N_18427,N_14618);
nor U27254 (N_27254,N_13031,N_15910);
nor U27255 (N_27255,N_18020,N_18581);
nor U27256 (N_27256,N_14788,N_15173);
and U27257 (N_27257,N_17004,N_12507);
nand U27258 (N_27258,N_17951,N_11314);
nand U27259 (N_27259,N_11043,N_17112);
nand U27260 (N_27260,N_15552,N_10374);
nand U27261 (N_27261,N_10679,N_16669);
xnor U27262 (N_27262,N_19112,N_16907);
nand U27263 (N_27263,N_15352,N_19268);
or U27264 (N_27264,N_19403,N_18444);
and U27265 (N_27265,N_10929,N_11490);
or U27266 (N_27266,N_11556,N_15292);
or U27267 (N_27267,N_12538,N_16652);
or U27268 (N_27268,N_10082,N_10409);
nor U27269 (N_27269,N_19494,N_18210);
or U27270 (N_27270,N_16307,N_12933);
or U27271 (N_27271,N_11583,N_17609);
nor U27272 (N_27272,N_18037,N_19809);
and U27273 (N_27273,N_18605,N_12598);
nor U27274 (N_27274,N_15338,N_15917);
nor U27275 (N_27275,N_17984,N_16621);
xor U27276 (N_27276,N_16615,N_12974);
xor U27277 (N_27277,N_19509,N_18133);
nor U27278 (N_27278,N_11652,N_16874);
or U27279 (N_27279,N_13990,N_12466);
nor U27280 (N_27280,N_19365,N_16070);
nor U27281 (N_27281,N_18035,N_14470);
nor U27282 (N_27282,N_10811,N_16086);
or U27283 (N_27283,N_16310,N_17684);
nor U27284 (N_27284,N_15383,N_18611);
xnor U27285 (N_27285,N_18172,N_19579);
xnor U27286 (N_27286,N_11263,N_14276);
nor U27287 (N_27287,N_19521,N_16186);
or U27288 (N_27288,N_15602,N_16120);
xor U27289 (N_27289,N_19705,N_10295);
or U27290 (N_27290,N_19813,N_19281);
and U27291 (N_27291,N_12208,N_18086);
or U27292 (N_27292,N_12381,N_10256);
nand U27293 (N_27293,N_12920,N_11769);
nor U27294 (N_27294,N_18141,N_18740);
nor U27295 (N_27295,N_17703,N_17281);
nor U27296 (N_27296,N_19761,N_10793);
and U27297 (N_27297,N_11905,N_10537);
and U27298 (N_27298,N_16923,N_14849);
or U27299 (N_27299,N_11906,N_15186);
xor U27300 (N_27300,N_18289,N_10208);
and U27301 (N_27301,N_15121,N_16117);
nand U27302 (N_27302,N_14347,N_17421);
nand U27303 (N_27303,N_11057,N_11449);
and U27304 (N_27304,N_19324,N_13351);
nor U27305 (N_27305,N_17254,N_14538);
or U27306 (N_27306,N_12113,N_18309);
nor U27307 (N_27307,N_17015,N_16235);
and U27308 (N_27308,N_17204,N_10137);
xnor U27309 (N_27309,N_16476,N_18854);
xnor U27310 (N_27310,N_16558,N_14529);
or U27311 (N_27311,N_18438,N_15157);
and U27312 (N_27312,N_17871,N_11365);
xor U27313 (N_27313,N_13234,N_17617);
and U27314 (N_27314,N_14819,N_18403);
nor U27315 (N_27315,N_18499,N_17964);
nand U27316 (N_27316,N_10622,N_12025);
and U27317 (N_27317,N_15339,N_13279);
nand U27318 (N_27318,N_12411,N_11473);
xor U27319 (N_27319,N_12356,N_15284);
and U27320 (N_27320,N_17046,N_17383);
xnor U27321 (N_27321,N_15241,N_11075);
and U27322 (N_27322,N_19446,N_15532);
xnor U27323 (N_27323,N_10598,N_12537);
nand U27324 (N_27324,N_16491,N_12071);
nand U27325 (N_27325,N_19288,N_16441);
and U27326 (N_27326,N_11750,N_12191);
and U27327 (N_27327,N_17485,N_14725);
or U27328 (N_27328,N_16864,N_12759);
nand U27329 (N_27329,N_10623,N_10045);
nand U27330 (N_27330,N_16274,N_11563);
nand U27331 (N_27331,N_17834,N_14328);
xor U27332 (N_27332,N_19535,N_16571);
nand U27333 (N_27333,N_18768,N_18611);
or U27334 (N_27334,N_13778,N_10601);
and U27335 (N_27335,N_15254,N_11293);
or U27336 (N_27336,N_16072,N_14778);
nand U27337 (N_27337,N_19545,N_17782);
and U27338 (N_27338,N_19447,N_18149);
or U27339 (N_27339,N_10448,N_15373);
or U27340 (N_27340,N_17613,N_12829);
nand U27341 (N_27341,N_12130,N_10057);
or U27342 (N_27342,N_10091,N_17943);
or U27343 (N_27343,N_11417,N_13184);
nand U27344 (N_27344,N_12862,N_19814);
xor U27345 (N_27345,N_16946,N_15130);
and U27346 (N_27346,N_11389,N_14447);
or U27347 (N_27347,N_11799,N_11038);
nand U27348 (N_27348,N_16871,N_11397);
nand U27349 (N_27349,N_16758,N_13771);
xnor U27350 (N_27350,N_15739,N_18348);
xnor U27351 (N_27351,N_19483,N_19407);
nand U27352 (N_27352,N_12117,N_17375);
or U27353 (N_27353,N_16842,N_15522);
nor U27354 (N_27354,N_18817,N_10137);
or U27355 (N_27355,N_16764,N_14774);
and U27356 (N_27356,N_15729,N_10257);
nand U27357 (N_27357,N_12799,N_10199);
or U27358 (N_27358,N_17689,N_13088);
and U27359 (N_27359,N_18529,N_16721);
nor U27360 (N_27360,N_12023,N_19995);
nor U27361 (N_27361,N_10449,N_15434);
xnor U27362 (N_27362,N_19732,N_18245);
nor U27363 (N_27363,N_16320,N_15490);
or U27364 (N_27364,N_16003,N_14826);
and U27365 (N_27365,N_12164,N_11573);
xor U27366 (N_27366,N_13905,N_18730);
and U27367 (N_27367,N_10956,N_11148);
nand U27368 (N_27368,N_13391,N_17647);
or U27369 (N_27369,N_13675,N_10957);
nor U27370 (N_27370,N_12089,N_14803);
or U27371 (N_27371,N_19524,N_14715);
xnor U27372 (N_27372,N_10552,N_17957);
or U27373 (N_27373,N_18984,N_18206);
or U27374 (N_27374,N_13652,N_15466);
xor U27375 (N_27375,N_19544,N_13991);
nor U27376 (N_27376,N_13939,N_11226);
or U27377 (N_27377,N_14793,N_13963);
nor U27378 (N_27378,N_19292,N_11699);
nand U27379 (N_27379,N_11055,N_12886);
or U27380 (N_27380,N_12620,N_17423);
or U27381 (N_27381,N_17266,N_18511);
nand U27382 (N_27382,N_12961,N_19428);
or U27383 (N_27383,N_19992,N_13113);
or U27384 (N_27384,N_14322,N_15833);
xor U27385 (N_27385,N_12389,N_15585);
and U27386 (N_27386,N_11638,N_15209);
nor U27387 (N_27387,N_10953,N_16622);
nor U27388 (N_27388,N_18083,N_14135);
xor U27389 (N_27389,N_10322,N_10017);
nor U27390 (N_27390,N_19696,N_11761);
nor U27391 (N_27391,N_17836,N_18213);
and U27392 (N_27392,N_11836,N_10715);
and U27393 (N_27393,N_17817,N_12978);
nand U27394 (N_27394,N_11917,N_12668);
xor U27395 (N_27395,N_13847,N_11479);
nand U27396 (N_27396,N_19913,N_12445);
or U27397 (N_27397,N_15796,N_16226);
nand U27398 (N_27398,N_11497,N_12122);
and U27399 (N_27399,N_11628,N_11888);
nand U27400 (N_27400,N_10119,N_18578);
xnor U27401 (N_27401,N_12373,N_11619);
or U27402 (N_27402,N_13775,N_12402);
and U27403 (N_27403,N_10423,N_19741);
xor U27404 (N_27404,N_15081,N_14959);
or U27405 (N_27405,N_10729,N_19340);
or U27406 (N_27406,N_19796,N_18858);
or U27407 (N_27407,N_15199,N_14417);
and U27408 (N_27408,N_17095,N_12952);
or U27409 (N_27409,N_13323,N_13148);
nor U27410 (N_27410,N_13691,N_16850);
and U27411 (N_27411,N_12234,N_13699);
and U27412 (N_27412,N_14714,N_13616);
xnor U27413 (N_27413,N_18053,N_12345);
and U27414 (N_27414,N_18251,N_19850);
or U27415 (N_27415,N_16260,N_13075);
nand U27416 (N_27416,N_15488,N_17951);
xnor U27417 (N_27417,N_15886,N_15313);
or U27418 (N_27418,N_12836,N_17731);
nor U27419 (N_27419,N_13271,N_15725);
nor U27420 (N_27420,N_15401,N_15417);
or U27421 (N_27421,N_16626,N_14740);
nor U27422 (N_27422,N_16142,N_18879);
or U27423 (N_27423,N_18443,N_14064);
and U27424 (N_27424,N_17354,N_18135);
nor U27425 (N_27425,N_17915,N_14141);
nand U27426 (N_27426,N_17435,N_18070);
xor U27427 (N_27427,N_19268,N_15671);
and U27428 (N_27428,N_14621,N_11201);
nand U27429 (N_27429,N_16144,N_16562);
xnor U27430 (N_27430,N_11755,N_15219);
nor U27431 (N_27431,N_14418,N_12898);
and U27432 (N_27432,N_10169,N_18531);
and U27433 (N_27433,N_19319,N_17207);
nor U27434 (N_27434,N_16464,N_11326);
nand U27435 (N_27435,N_11001,N_19936);
or U27436 (N_27436,N_15250,N_15084);
xnor U27437 (N_27437,N_17551,N_12488);
and U27438 (N_27438,N_19162,N_14098);
nor U27439 (N_27439,N_10457,N_15432);
or U27440 (N_27440,N_18017,N_11954);
nor U27441 (N_27441,N_15322,N_19228);
nand U27442 (N_27442,N_11898,N_18888);
xnor U27443 (N_27443,N_17742,N_16934);
nor U27444 (N_27444,N_13666,N_16308);
nand U27445 (N_27445,N_19792,N_10342);
xnor U27446 (N_27446,N_16932,N_18924);
nor U27447 (N_27447,N_16768,N_15269);
and U27448 (N_27448,N_15634,N_11030);
nand U27449 (N_27449,N_19249,N_10413);
nor U27450 (N_27450,N_13431,N_16319);
xor U27451 (N_27451,N_14592,N_17603);
and U27452 (N_27452,N_16663,N_12553);
nand U27453 (N_27453,N_11519,N_17560);
and U27454 (N_27454,N_18829,N_14597);
and U27455 (N_27455,N_11749,N_13161);
xnor U27456 (N_27456,N_13738,N_10901);
and U27457 (N_27457,N_13084,N_14780);
nor U27458 (N_27458,N_13084,N_15877);
nor U27459 (N_27459,N_17908,N_17415);
and U27460 (N_27460,N_18185,N_15272);
nand U27461 (N_27461,N_16400,N_14334);
nand U27462 (N_27462,N_18442,N_11063);
nor U27463 (N_27463,N_10888,N_12108);
nand U27464 (N_27464,N_14757,N_15718);
or U27465 (N_27465,N_10353,N_12229);
and U27466 (N_27466,N_10583,N_10353);
or U27467 (N_27467,N_19713,N_15888);
nand U27468 (N_27468,N_15612,N_18057);
or U27469 (N_27469,N_10020,N_11297);
xnor U27470 (N_27470,N_14889,N_13105);
and U27471 (N_27471,N_10126,N_14384);
or U27472 (N_27472,N_18170,N_13636);
nand U27473 (N_27473,N_17146,N_14996);
or U27474 (N_27474,N_18970,N_11895);
nand U27475 (N_27475,N_15792,N_16585);
and U27476 (N_27476,N_14779,N_14044);
nand U27477 (N_27477,N_12119,N_16881);
nand U27478 (N_27478,N_14784,N_10272);
and U27479 (N_27479,N_19891,N_12591);
nor U27480 (N_27480,N_14071,N_13951);
xnor U27481 (N_27481,N_18397,N_12626);
or U27482 (N_27482,N_15415,N_15094);
nor U27483 (N_27483,N_12710,N_14481);
xnor U27484 (N_27484,N_12172,N_11789);
nor U27485 (N_27485,N_17379,N_14725);
nand U27486 (N_27486,N_16834,N_17832);
xor U27487 (N_27487,N_10538,N_13966);
and U27488 (N_27488,N_17819,N_12920);
and U27489 (N_27489,N_13145,N_16367);
nand U27490 (N_27490,N_11419,N_10610);
nand U27491 (N_27491,N_14488,N_17535);
xnor U27492 (N_27492,N_18635,N_11954);
or U27493 (N_27493,N_10034,N_18594);
nand U27494 (N_27494,N_15931,N_16783);
or U27495 (N_27495,N_16021,N_14614);
nand U27496 (N_27496,N_17113,N_14234);
or U27497 (N_27497,N_17258,N_10645);
and U27498 (N_27498,N_14898,N_11538);
and U27499 (N_27499,N_16352,N_19768);
xor U27500 (N_27500,N_11886,N_11734);
nor U27501 (N_27501,N_15252,N_15374);
xor U27502 (N_27502,N_15141,N_12966);
nand U27503 (N_27503,N_15528,N_15684);
xnor U27504 (N_27504,N_17401,N_10039);
nand U27505 (N_27505,N_19772,N_18162);
and U27506 (N_27506,N_15819,N_18765);
xor U27507 (N_27507,N_18255,N_15430);
nor U27508 (N_27508,N_17966,N_18864);
nand U27509 (N_27509,N_10927,N_12027);
xor U27510 (N_27510,N_11284,N_15746);
and U27511 (N_27511,N_19926,N_12486);
nand U27512 (N_27512,N_19559,N_15640);
xor U27513 (N_27513,N_15636,N_16830);
or U27514 (N_27514,N_10765,N_18380);
nor U27515 (N_27515,N_10999,N_19692);
and U27516 (N_27516,N_12615,N_11000);
nor U27517 (N_27517,N_11852,N_16498);
or U27518 (N_27518,N_15984,N_14773);
nor U27519 (N_27519,N_18218,N_10767);
or U27520 (N_27520,N_17891,N_13161);
and U27521 (N_27521,N_14730,N_12538);
nand U27522 (N_27522,N_13506,N_14847);
nand U27523 (N_27523,N_18143,N_14024);
nor U27524 (N_27524,N_18134,N_10556);
xnor U27525 (N_27525,N_16002,N_15705);
nor U27526 (N_27526,N_10195,N_16979);
nand U27527 (N_27527,N_12638,N_11769);
xnor U27528 (N_27528,N_14166,N_15974);
nor U27529 (N_27529,N_16921,N_14545);
nand U27530 (N_27530,N_18913,N_15487);
and U27531 (N_27531,N_18854,N_19426);
or U27532 (N_27532,N_10627,N_14694);
and U27533 (N_27533,N_16000,N_12830);
and U27534 (N_27534,N_15340,N_12737);
and U27535 (N_27535,N_16881,N_10644);
nand U27536 (N_27536,N_13010,N_17727);
nor U27537 (N_27537,N_11485,N_13821);
xnor U27538 (N_27538,N_14941,N_18528);
nor U27539 (N_27539,N_17816,N_18087);
nand U27540 (N_27540,N_14669,N_16029);
xnor U27541 (N_27541,N_18804,N_12968);
or U27542 (N_27542,N_14084,N_15930);
and U27543 (N_27543,N_14411,N_19216);
and U27544 (N_27544,N_11524,N_10396);
nor U27545 (N_27545,N_14554,N_10000);
nor U27546 (N_27546,N_13775,N_12386);
xnor U27547 (N_27547,N_19881,N_16899);
or U27548 (N_27548,N_10710,N_12812);
nor U27549 (N_27549,N_19956,N_12549);
or U27550 (N_27550,N_16702,N_17725);
and U27551 (N_27551,N_11785,N_11711);
or U27552 (N_27552,N_12107,N_17013);
and U27553 (N_27553,N_17706,N_15186);
nor U27554 (N_27554,N_15162,N_13011);
xor U27555 (N_27555,N_19977,N_11534);
nor U27556 (N_27556,N_15531,N_15130);
nand U27557 (N_27557,N_17998,N_10524);
nand U27558 (N_27558,N_17517,N_16213);
nand U27559 (N_27559,N_15335,N_19331);
and U27560 (N_27560,N_19490,N_11325);
or U27561 (N_27561,N_18554,N_10143);
xor U27562 (N_27562,N_17714,N_14132);
nor U27563 (N_27563,N_10606,N_18528);
and U27564 (N_27564,N_12311,N_13730);
nand U27565 (N_27565,N_19171,N_13694);
nor U27566 (N_27566,N_14820,N_14433);
xnor U27567 (N_27567,N_13124,N_15262);
or U27568 (N_27568,N_12856,N_16558);
nor U27569 (N_27569,N_12499,N_18611);
nor U27570 (N_27570,N_14081,N_10717);
or U27571 (N_27571,N_11004,N_15507);
nand U27572 (N_27572,N_16943,N_19945);
and U27573 (N_27573,N_17315,N_14785);
or U27574 (N_27574,N_19005,N_19032);
nor U27575 (N_27575,N_11816,N_12061);
and U27576 (N_27576,N_17671,N_19678);
xor U27577 (N_27577,N_13452,N_15153);
and U27578 (N_27578,N_15298,N_18609);
xnor U27579 (N_27579,N_13998,N_19703);
and U27580 (N_27580,N_16046,N_15665);
and U27581 (N_27581,N_11612,N_19203);
or U27582 (N_27582,N_17585,N_16734);
and U27583 (N_27583,N_18464,N_11826);
and U27584 (N_27584,N_19897,N_12083);
or U27585 (N_27585,N_10141,N_18562);
xor U27586 (N_27586,N_12356,N_10387);
nor U27587 (N_27587,N_18508,N_15053);
nor U27588 (N_27588,N_11315,N_14747);
nand U27589 (N_27589,N_19138,N_17714);
nor U27590 (N_27590,N_18261,N_10514);
nor U27591 (N_27591,N_11789,N_19140);
nor U27592 (N_27592,N_18869,N_16795);
nand U27593 (N_27593,N_11549,N_13690);
nand U27594 (N_27594,N_17544,N_11140);
or U27595 (N_27595,N_12123,N_17050);
or U27596 (N_27596,N_19596,N_12165);
nor U27597 (N_27597,N_19648,N_19622);
or U27598 (N_27598,N_19755,N_17885);
xor U27599 (N_27599,N_15929,N_15767);
nor U27600 (N_27600,N_11532,N_11567);
nor U27601 (N_27601,N_14502,N_16615);
and U27602 (N_27602,N_13193,N_14516);
nand U27603 (N_27603,N_17205,N_14448);
and U27604 (N_27604,N_18800,N_14163);
xor U27605 (N_27605,N_10887,N_13625);
and U27606 (N_27606,N_19793,N_13940);
or U27607 (N_27607,N_17353,N_12464);
xnor U27608 (N_27608,N_17020,N_13867);
xnor U27609 (N_27609,N_19788,N_14650);
xnor U27610 (N_27610,N_15369,N_19276);
or U27611 (N_27611,N_14789,N_19879);
nand U27612 (N_27612,N_11544,N_12822);
nand U27613 (N_27613,N_11840,N_14526);
nor U27614 (N_27614,N_19410,N_19351);
nor U27615 (N_27615,N_18635,N_15140);
and U27616 (N_27616,N_10836,N_16261);
xor U27617 (N_27617,N_11955,N_18816);
nor U27618 (N_27618,N_12351,N_12692);
nor U27619 (N_27619,N_14572,N_18089);
nor U27620 (N_27620,N_15497,N_18262);
nand U27621 (N_27621,N_10555,N_14618);
and U27622 (N_27622,N_10257,N_10012);
and U27623 (N_27623,N_11339,N_13843);
nand U27624 (N_27624,N_12759,N_18685);
and U27625 (N_27625,N_17224,N_15221);
xnor U27626 (N_27626,N_13113,N_13547);
nor U27627 (N_27627,N_15118,N_13032);
nand U27628 (N_27628,N_19757,N_13039);
and U27629 (N_27629,N_13181,N_14216);
xor U27630 (N_27630,N_13458,N_12579);
nor U27631 (N_27631,N_18711,N_14016);
or U27632 (N_27632,N_10643,N_17155);
and U27633 (N_27633,N_14240,N_17628);
and U27634 (N_27634,N_14159,N_13164);
nand U27635 (N_27635,N_14331,N_15651);
and U27636 (N_27636,N_10959,N_14159);
or U27637 (N_27637,N_12009,N_15958);
and U27638 (N_27638,N_15312,N_19040);
and U27639 (N_27639,N_10769,N_16463);
and U27640 (N_27640,N_18490,N_15626);
or U27641 (N_27641,N_11420,N_11533);
nand U27642 (N_27642,N_14372,N_14445);
xnor U27643 (N_27643,N_12116,N_13960);
nor U27644 (N_27644,N_16836,N_12959);
and U27645 (N_27645,N_13803,N_18657);
or U27646 (N_27646,N_15804,N_10589);
and U27647 (N_27647,N_16153,N_18315);
or U27648 (N_27648,N_16039,N_14830);
and U27649 (N_27649,N_11518,N_18669);
nand U27650 (N_27650,N_14501,N_10308);
xnor U27651 (N_27651,N_19322,N_13112);
nand U27652 (N_27652,N_11659,N_10627);
or U27653 (N_27653,N_12388,N_12724);
or U27654 (N_27654,N_18442,N_10800);
xnor U27655 (N_27655,N_17915,N_13452);
nand U27656 (N_27656,N_13871,N_18341);
or U27657 (N_27657,N_17753,N_19918);
or U27658 (N_27658,N_19833,N_13577);
xor U27659 (N_27659,N_18001,N_10754);
or U27660 (N_27660,N_13604,N_10939);
or U27661 (N_27661,N_12268,N_16231);
xnor U27662 (N_27662,N_15937,N_11997);
nand U27663 (N_27663,N_14680,N_16551);
nor U27664 (N_27664,N_13924,N_10296);
or U27665 (N_27665,N_11316,N_17554);
and U27666 (N_27666,N_14070,N_11662);
nor U27667 (N_27667,N_10479,N_13321);
and U27668 (N_27668,N_15803,N_15789);
or U27669 (N_27669,N_12323,N_13645);
and U27670 (N_27670,N_19259,N_10770);
xor U27671 (N_27671,N_12297,N_14399);
xnor U27672 (N_27672,N_15459,N_18237);
or U27673 (N_27673,N_16533,N_10055);
xnor U27674 (N_27674,N_16286,N_10749);
nor U27675 (N_27675,N_13156,N_19597);
nand U27676 (N_27676,N_12900,N_18395);
and U27677 (N_27677,N_14042,N_18805);
nor U27678 (N_27678,N_11681,N_11075);
xnor U27679 (N_27679,N_10029,N_19351);
and U27680 (N_27680,N_19343,N_13804);
nor U27681 (N_27681,N_15126,N_18705);
and U27682 (N_27682,N_13885,N_11430);
nand U27683 (N_27683,N_10537,N_16256);
nor U27684 (N_27684,N_10050,N_19923);
or U27685 (N_27685,N_18567,N_13836);
xnor U27686 (N_27686,N_17775,N_11485);
xnor U27687 (N_27687,N_17692,N_16878);
or U27688 (N_27688,N_12689,N_18669);
xor U27689 (N_27689,N_16754,N_11640);
or U27690 (N_27690,N_14613,N_18965);
xor U27691 (N_27691,N_14282,N_10245);
xnor U27692 (N_27692,N_16495,N_14314);
or U27693 (N_27693,N_16792,N_18745);
or U27694 (N_27694,N_10781,N_13676);
or U27695 (N_27695,N_17588,N_16135);
nor U27696 (N_27696,N_16110,N_10444);
nor U27697 (N_27697,N_17606,N_11401);
xnor U27698 (N_27698,N_10653,N_15859);
xor U27699 (N_27699,N_10073,N_10298);
xnor U27700 (N_27700,N_19881,N_19265);
nand U27701 (N_27701,N_10324,N_12818);
xor U27702 (N_27702,N_19079,N_16708);
nand U27703 (N_27703,N_15537,N_12751);
nor U27704 (N_27704,N_17727,N_13762);
and U27705 (N_27705,N_16055,N_13941);
nand U27706 (N_27706,N_15788,N_14530);
xnor U27707 (N_27707,N_11793,N_16162);
xor U27708 (N_27708,N_13048,N_12792);
nand U27709 (N_27709,N_15267,N_19795);
xnor U27710 (N_27710,N_11110,N_10053);
or U27711 (N_27711,N_17134,N_17858);
or U27712 (N_27712,N_14167,N_18692);
or U27713 (N_27713,N_15524,N_12041);
nand U27714 (N_27714,N_18092,N_19828);
or U27715 (N_27715,N_10769,N_11013);
or U27716 (N_27716,N_16738,N_14803);
and U27717 (N_27717,N_15341,N_15310);
xor U27718 (N_27718,N_15891,N_13004);
xor U27719 (N_27719,N_13459,N_12757);
nand U27720 (N_27720,N_19045,N_16441);
and U27721 (N_27721,N_15836,N_12912);
and U27722 (N_27722,N_14350,N_19228);
xnor U27723 (N_27723,N_19453,N_13357);
xor U27724 (N_27724,N_18398,N_15270);
xor U27725 (N_27725,N_15108,N_11073);
or U27726 (N_27726,N_19813,N_15657);
nand U27727 (N_27727,N_19746,N_10373);
xnor U27728 (N_27728,N_10253,N_18688);
nor U27729 (N_27729,N_15276,N_16911);
nor U27730 (N_27730,N_11683,N_17227);
nor U27731 (N_27731,N_15727,N_15520);
nand U27732 (N_27732,N_11034,N_10541);
nor U27733 (N_27733,N_13537,N_13479);
nand U27734 (N_27734,N_14627,N_18863);
or U27735 (N_27735,N_12594,N_19668);
and U27736 (N_27736,N_16434,N_18428);
nor U27737 (N_27737,N_18779,N_12344);
xnor U27738 (N_27738,N_19208,N_15466);
or U27739 (N_27739,N_18214,N_11551);
nand U27740 (N_27740,N_11708,N_11914);
nor U27741 (N_27741,N_15394,N_11895);
xnor U27742 (N_27742,N_12888,N_14693);
xnor U27743 (N_27743,N_10771,N_17213);
xnor U27744 (N_27744,N_14066,N_13060);
and U27745 (N_27745,N_12633,N_14921);
or U27746 (N_27746,N_18422,N_16180);
nand U27747 (N_27747,N_16064,N_19828);
xnor U27748 (N_27748,N_10308,N_12087);
xor U27749 (N_27749,N_15978,N_11132);
and U27750 (N_27750,N_14884,N_13058);
nor U27751 (N_27751,N_12707,N_17839);
or U27752 (N_27752,N_14534,N_18192);
and U27753 (N_27753,N_17052,N_11532);
and U27754 (N_27754,N_18982,N_14252);
or U27755 (N_27755,N_10582,N_11262);
nor U27756 (N_27756,N_17689,N_14022);
nand U27757 (N_27757,N_14548,N_14338);
xor U27758 (N_27758,N_15860,N_16271);
nand U27759 (N_27759,N_12481,N_16860);
or U27760 (N_27760,N_19921,N_14745);
or U27761 (N_27761,N_18543,N_17623);
nand U27762 (N_27762,N_13456,N_13976);
or U27763 (N_27763,N_17146,N_11890);
or U27764 (N_27764,N_16584,N_12883);
xnor U27765 (N_27765,N_16551,N_19564);
xnor U27766 (N_27766,N_14301,N_13040);
and U27767 (N_27767,N_18766,N_16308);
xor U27768 (N_27768,N_10677,N_15667);
nor U27769 (N_27769,N_14775,N_12891);
nor U27770 (N_27770,N_18685,N_17614);
nand U27771 (N_27771,N_17314,N_12062);
nor U27772 (N_27772,N_16868,N_15683);
nor U27773 (N_27773,N_18340,N_18435);
or U27774 (N_27774,N_13493,N_15481);
nand U27775 (N_27775,N_13064,N_18499);
xnor U27776 (N_27776,N_17759,N_11551);
nand U27777 (N_27777,N_17006,N_11144);
xnor U27778 (N_27778,N_13929,N_11485);
nor U27779 (N_27779,N_14389,N_14174);
nand U27780 (N_27780,N_19572,N_18304);
or U27781 (N_27781,N_17722,N_11022);
nor U27782 (N_27782,N_12557,N_16329);
or U27783 (N_27783,N_13565,N_17088);
nor U27784 (N_27784,N_19470,N_17907);
nor U27785 (N_27785,N_12108,N_11078);
or U27786 (N_27786,N_18274,N_12668);
or U27787 (N_27787,N_16022,N_16724);
or U27788 (N_27788,N_19201,N_18250);
xnor U27789 (N_27789,N_11465,N_16632);
nand U27790 (N_27790,N_10502,N_16003);
nor U27791 (N_27791,N_15195,N_14797);
and U27792 (N_27792,N_16599,N_18991);
or U27793 (N_27793,N_13244,N_11343);
and U27794 (N_27794,N_16722,N_10596);
xnor U27795 (N_27795,N_12203,N_13452);
or U27796 (N_27796,N_14847,N_12913);
nand U27797 (N_27797,N_16050,N_15509);
xnor U27798 (N_27798,N_18256,N_16062);
and U27799 (N_27799,N_15527,N_10171);
and U27800 (N_27800,N_14368,N_15810);
nor U27801 (N_27801,N_19635,N_18572);
or U27802 (N_27802,N_16580,N_19601);
nor U27803 (N_27803,N_14308,N_12475);
nor U27804 (N_27804,N_14106,N_17483);
or U27805 (N_27805,N_14819,N_18903);
and U27806 (N_27806,N_11857,N_13152);
nor U27807 (N_27807,N_14755,N_17214);
nand U27808 (N_27808,N_11537,N_11342);
or U27809 (N_27809,N_14020,N_14706);
nand U27810 (N_27810,N_15673,N_17929);
and U27811 (N_27811,N_17205,N_15827);
or U27812 (N_27812,N_17904,N_14535);
or U27813 (N_27813,N_12759,N_16972);
nand U27814 (N_27814,N_13015,N_11064);
or U27815 (N_27815,N_16808,N_11508);
xnor U27816 (N_27816,N_17799,N_13514);
xor U27817 (N_27817,N_13730,N_19972);
and U27818 (N_27818,N_19562,N_17189);
or U27819 (N_27819,N_12677,N_14581);
nand U27820 (N_27820,N_17599,N_13880);
and U27821 (N_27821,N_11037,N_19044);
and U27822 (N_27822,N_17930,N_15986);
nand U27823 (N_27823,N_13134,N_11677);
nand U27824 (N_27824,N_18271,N_16756);
nand U27825 (N_27825,N_14098,N_18833);
nand U27826 (N_27826,N_15134,N_16435);
or U27827 (N_27827,N_10952,N_16725);
and U27828 (N_27828,N_15335,N_15979);
and U27829 (N_27829,N_18992,N_10534);
nor U27830 (N_27830,N_12167,N_15271);
nor U27831 (N_27831,N_11312,N_13605);
xnor U27832 (N_27832,N_17606,N_19445);
or U27833 (N_27833,N_10853,N_14822);
nand U27834 (N_27834,N_10785,N_18515);
nand U27835 (N_27835,N_17062,N_19712);
or U27836 (N_27836,N_16491,N_10773);
and U27837 (N_27837,N_16528,N_10999);
or U27838 (N_27838,N_17792,N_14902);
xnor U27839 (N_27839,N_10070,N_11459);
xnor U27840 (N_27840,N_19436,N_17436);
or U27841 (N_27841,N_19162,N_16560);
or U27842 (N_27842,N_10725,N_16959);
and U27843 (N_27843,N_19200,N_15550);
nand U27844 (N_27844,N_13242,N_13777);
xnor U27845 (N_27845,N_13194,N_12774);
or U27846 (N_27846,N_18209,N_12850);
xnor U27847 (N_27847,N_18907,N_15803);
or U27848 (N_27848,N_14354,N_14264);
xnor U27849 (N_27849,N_11327,N_17265);
xnor U27850 (N_27850,N_17826,N_15066);
nand U27851 (N_27851,N_10739,N_12509);
nor U27852 (N_27852,N_16929,N_15473);
nand U27853 (N_27853,N_11467,N_10638);
nor U27854 (N_27854,N_17046,N_11952);
and U27855 (N_27855,N_12990,N_14452);
nor U27856 (N_27856,N_17040,N_18807);
nand U27857 (N_27857,N_14083,N_13464);
and U27858 (N_27858,N_12747,N_17202);
xnor U27859 (N_27859,N_10759,N_12170);
nor U27860 (N_27860,N_14010,N_16722);
nand U27861 (N_27861,N_17622,N_11487);
or U27862 (N_27862,N_10751,N_13389);
nand U27863 (N_27863,N_11282,N_16634);
nand U27864 (N_27864,N_10584,N_10312);
or U27865 (N_27865,N_12781,N_18697);
and U27866 (N_27866,N_12945,N_19992);
and U27867 (N_27867,N_16948,N_15037);
or U27868 (N_27868,N_18029,N_18014);
xnor U27869 (N_27869,N_15968,N_12911);
or U27870 (N_27870,N_19782,N_14997);
and U27871 (N_27871,N_16744,N_16254);
or U27872 (N_27872,N_11542,N_16516);
and U27873 (N_27873,N_18508,N_11028);
or U27874 (N_27874,N_17663,N_12253);
nand U27875 (N_27875,N_10545,N_14179);
nand U27876 (N_27876,N_18345,N_11378);
or U27877 (N_27877,N_13632,N_19578);
nand U27878 (N_27878,N_18226,N_17058);
and U27879 (N_27879,N_12030,N_11919);
xor U27880 (N_27880,N_17786,N_12397);
nand U27881 (N_27881,N_14276,N_15210);
and U27882 (N_27882,N_16404,N_11462);
nand U27883 (N_27883,N_19990,N_12871);
nand U27884 (N_27884,N_11687,N_10022);
nor U27885 (N_27885,N_11410,N_16493);
xnor U27886 (N_27886,N_10285,N_19437);
nand U27887 (N_27887,N_15989,N_10243);
xnor U27888 (N_27888,N_16594,N_15728);
nand U27889 (N_27889,N_19543,N_14906);
nand U27890 (N_27890,N_17208,N_15522);
nand U27891 (N_27891,N_14464,N_18707);
xnor U27892 (N_27892,N_18965,N_15368);
nor U27893 (N_27893,N_16477,N_15402);
and U27894 (N_27894,N_12405,N_16177);
xnor U27895 (N_27895,N_18587,N_17184);
nor U27896 (N_27896,N_13037,N_16735);
nand U27897 (N_27897,N_19961,N_15109);
nand U27898 (N_27898,N_18391,N_12582);
or U27899 (N_27899,N_11696,N_14954);
nand U27900 (N_27900,N_11765,N_17042);
xor U27901 (N_27901,N_19874,N_16468);
nor U27902 (N_27902,N_15678,N_14491);
and U27903 (N_27903,N_17531,N_19007);
xnor U27904 (N_27904,N_10938,N_15096);
xor U27905 (N_27905,N_10777,N_18837);
nor U27906 (N_27906,N_19783,N_13755);
nor U27907 (N_27907,N_18392,N_15706);
nor U27908 (N_27908,N_16525,N_10418);
or U27909 (N_27909,N_12620,N_17167);
or U27910 (N_27910,N_13597,N_10578);
and U27911 (N_27911,N_10867,N_13897);
nand U27912 (N_27912,N_14307,N_18550);
xnor U27913 (N_27913,N_11822,N_15031);
xnor U27914 (N_27914,N_19781,N_12223);
xor U27915 (N_27915,N_10227,N_19152);
nand U27916 (N_27916,N_15262,N_14165);
xor U27917 (N_27917,N_10911,N_11396);
or U27918 (N_27918,N_15561,N_14583);
nor U27919 (N_27919,N_19550,N_15330);
and U27920 (N_27920,N_17633,N_14446);
and U27921 (N_27921,N_12285,N_15212);
or U27922 (N_27922,N_12555,N_13935);
nand U27923 (N_27923,N_18372,N_16880);
nor U27924 (N_27924,N_13704,N_11081);
or U27925 (N_27925,N_10156,N_15378);
or U27926 (N_27926,N_14109,N_14144);
nor U27927 (N_27927,N_18547,N_18666);
nor U27928 (N_27928,N_13771,N_17529);
xnor U27929 (N_27929,N_12460,N_17083);
or U27930 (N_27930,N_16692,N_19796);
or U27931 (N_27931,N_11841,N_13335);
or U27932 (N_27932,N_18275,N_10448);
or U27933 (N_27933,N_12271,N_11401);
and U27934 (N_27934,N_19904,N_11704);
nand U27935 (N_27935,N_14500,N_13797);
nor U27936 (N_27936,N_14100,N_14196);
or U27937 (N_27937,N_19876,N_12757);
or U27938 (N_27938,N_11799,N_13463);
or U27939 (N_27939,N_17676,N_18573);
xor U27940 (N_27940,N_10567,N_11002);
nand U27941 (N_27941,N_10645,N_13740);
and U27942 (N_27942,N_12992,N_12476);
xor U27943 (N_27943,N_10287,N_13815);
xor U27944 (N_27944,N_10070,N_16481);
nor U27945 (N_27945,N_19874,N_15895);
or U27946 (N_27946,N_11362,N_19818);
nand U27947 (N_27947,N_10964,N_14455);
and U27948 (N_27948,N_12576,N_14318);
and U27949 (N_27949,N_16049,N_16932);
xnor U27950 (N_27950,N_11463,N_16071);
and U27951 (N_27951,N_15524,N_10682);
xor U27952 (N_27952,N_13336,N_14396);
nor U27953 (N_27953,N_17372,N_17270);
or U27954 (N_27954,N_16488,N_19818);
nor U27955 (N_27955,N_18593,N_15083);
nor U27956 (N_27956,N_16334,N_17918);
xor U27957 (N_27957,N_18728,N_13027);
xnor U27958 (N_27958,N_19152,N_17130);
nand U27959 (N_27959,N_10472,N_13665);
nand U27960 (N_27960,N_14318,N_17251);
or U27961 (N_27961,N_14995,N_16086);
xnor U27962 (N_27962,N_12176,N_11716);
nand U27963 (N_27963,N_13233,N_17448);
and U27964 (N_27964,N_13100,N_15177);
and U27965 (N_27965,N_15151,N_17308);
and U27966 (N_27966,N_19245,N_16768);
nand U27967 (N_27967,N_15090,N_11836);
nand U27968 (N_27968,N_18032,N_15600);
nand U27969 (N_27969,N_15161,N_16571);
nor U27970 (N_27970,N_11865,N_17507);
and U27971 (N_27971,N_18148,N_16730);
nor U27972 (N_27972,N_15019,N_19832);
xor U27973 (N_27973,N_16370,N_19444);
and U27974 (N_27974,N_18425,N_12921);
nand U27975 (N_27975,N_11159,N_14319);
or U27976 (N_27976,N_14380,N_12126);
or U27977 (N_27977,N_12706,N_16551);
nor U27978 (N_27978,N_11184,N_13914);
and U27979 (N_27979,N_17762,N_12359);
nand U27980 (N_27980,N_11473,N_11967);
xnor U27981 (N_27981,N_15819,N_19287);
and U27982 (N_27982,N_10912,N_18020);
nor U27983 (N_27983,N_13451,N_15992);
nor U27984 (N_27984,N_13069,N_14360);
nand U27985 (N_27985,N_19888,N_11978);
and U27986 (N_27986,N_16478,N_19652);
nand U27987 (N_27987,N_13259,N_16966);
and U27988 (N_27988,N_16648,N_12441);
nand U27989 (N_27989,N_16208,N_14863);
xnor U27990 (N_27990,N_19076,N_16088);
or U27991 (N_27991,N_10530,N_15500);
xor U27992 (N_27992,N_14086,N_11240);
or U27993 (N_27993,N_12894,N_10331);
nor U27994 (N_27994,N_18006,N_13040);
nor U27995 (N_27995,N_17059,N_10522);
xnor U27996 (N_27996,N_16998,N_15440);
nand U27997 (N_27997,N_15113,N_16476);
nand U27998 (N_27998,N_19585,N_16138);
nand U27999 (N_27999,N_14998,N_19359);
nor U28000 (N_28000,N_13875,N_18517);
and U28001 (N_28001,N_18917,N_13035);
nor U28002 (N_28002,N_14791,N_13628);
and U28003 (N_28003,N_11456,N_16339);
nor U28004 (N_28004,N_10964,N_17069);
xnor U28005 (N_28005,N_10982,N_18593);
or U28006 (N_28006,N_17732,N_10809);
nor U28007 (N_28007,N_13338,N_11993);
nand U28008 (N_28008,N_18090,N_15766);
xnor U28009 (N_28009,N_14175,N_13002);
xor U28010 (N_28010,N_19641,N_15277);
nor U28011 (N_28011,N_13786,N_14856);
nor U28012 (N_28012,N_10230,N_13728);
xnor U28013 (N_28013,N_17879,N_14688);
or U28014 (N_28014,N_16037,N_17176);
nor U28015 (N_28015,N_11710,N_12138);
nand U28016 (N_28016,N_14513,N_14034);
or U28017 (N_28017,N_11093,N_11355);
and U28018 (N_28018,N_14014,N_19326);
and U28019 (N_28019,N_16164,N_15851);
xnor U28020 (N_28020,N_15801,N_13792);
or U28021 (N_28021,N_13650,N_19374);
and U28022 (N_28022,N_19729,N_15049);
nand U28023 (N_28023,N_17561,N_14633);
or U28024 (N_28024,N_11686,N_13097);
or U28025 (N_28025,N_11561,N_15243);
nor U28026 (N_28026,N_17564,N_17128);
or U28027 (N_28027,N_17465,N_14454);
and U28028 (N_28028,N_13676,N_10106);
nor U28029 (N_28029,N_16002,N_12551);
or U28030 (N_28030,N_17862,N_17208);
nor U28031 (N_28031,N_11663,N_18743);
xnor U28032 (N_28032,N_17130,N_16725);
nor U28033 (N_28033,N_11814,N_15533);
xnor U28034 (N_28034,N_19203,N_15290);
nand U28035 (N_28035,N_10843,N_18170);
xnor U28036 (N_28036,N_14868,N_16247);
nand U28037 (N_28037,N_17977,N_15494);
xor U28038 (N_28038,N_13008,N_12263);
xnor U28039 (N_28039,N_10554,N_17129);
xor U28040 (N_28040,N_13733,N_14775);
nor U28041 (N_28041,N_16094,N_18004);
nor U28042 (N_28042,N_17674,N_12458);
xnor U28043 (N_28043,N_16597,N_14931);
nor U28044 (N_28044,N_13736,N_12842);
nor U28045 (N_28045,N_10049,N_11180);
nor U28046 (N_28046,N_14017,N_14495);
nand U28047 (N_28047,N_13871,N_15737);
and U28048 (N_28048,N_15247,N_15354);
and U28049 (N_28049,N_12642,N_10381);
nor U28050 (N_28050,N_11851,N_12697);
xor U28051 (N_28051,N_12415,N_16147);
and U28052 (N_28052,N_12085,N_12128);
nand U28053 (N_28053,N_11337,N_11613);
xnor U28054 (N_28054,N_16905,N_17617);
nor U28055 (N_28055,N_14647,N_14878);
nand U28056 (N_28056,N_17399,N_11892);
nor U28057 (N_28057,N_17691,N_13242);
nor U28058 (N_28058,N_18460,N_10921);
nor U28059 (N_28059,N_11283,N_12051);
xnor U28060 (N_28060,N_14219,N_11868);
and U28061 (N_28061,N_10257,N_12070);
and U28062 (N_28062,N_10313,N_12310);
nor U28063 (N_28063,N_19580,N_14330);
nand U28064 (N_28064,N_14972,N_17686);
or U28065 (N_28065,N_12351,N_13727);
xnor U28066 (N_28066,N_10568,N_18456);
nand U28067 (N_28067,N_17213,N_11569);
and U28068 (N_28068,N_14196,N_15744);
xnor U28069 (N_28069,N_11662,N_10629);
nor U28070 (N_28070,N_19631,N_10357);
and U28071 (N_28071,N_12509,N_10595);
nand U28072 (N_28072,N_14771,N_10016);
xor U28073 (N_28073,N_14654,N_18506);
nor U28074 (N_28074,N_13868,N_15452);
nand U28075 (N_28075,N_18966,N_16285);
xor U28076 (N_28076,N_10859,N_14627);
nand U28077 (N_28077,N_18613,N_18800);
nand U28078 (N_28078,N_10806,N_11091);
xnor U28079 (N_28079,N_12453,N_15022);
nor U28080 (N_28080,N_11385,N_15634);
nand U28081 (N_28081,N_16763,N_19437);
and U28082 (N_28082,N_12644,N_14655);
nand U28083 (N_28083,N_12074,N_15942);
or U28084 (N_28084,N_13934,N_13032);
nand U28085 (N_28085,N_15081,N_12634);
and U28086 (N_28086,N_15526,N_12314);
nor U28087 (N_28087,N_18922,N_12508);
nor U28088 (N_28088,N_18204,N_10977);
xnor U28089 (N_28089,N_18315,N_13620);
nand U28090 (N_28090,N_19727,N_12363);
nor U28091 (N_28091,N_12666,N_13841);
xor U28092 (N_28092,N_16428,N_12994);
nor U28093 (N_28093,N_14943,N_16802);
nand U28094 (N_28094,N_12890,N_18362);
xor U28095 (N_28095,N_11109,N_13946);
nor U28096 (N_28096,N_12404,N_17719);
or U28097 (N_28097,N_17939,N_17746);
or U28098 (N_28098,N_12658,N_15750);
or U28099 (N_28099,N_15052,N_13980);
or U28100 (N_28100,N_15992,N_10181);
nand U28101 (N_28101,N_11589,N_16333);
nand U28102 (N_28102,N_16764,N_19802);
or U28103 (N_28103,N_18660,N_15310);
nand U28104 (N_28104,N_18672,N_15438);
xor U28105 (N_28105,N_14904,N_12650);
and U28106 (N_28106,N_12204,N_17801);
xnor U28107 (N_28107,N_11933,N_11602);
and U28108 (N_28108,N_17500,N_19559);
nor U28109 (N_28109,N_14027,N_19363);
or U28110 (N_28110,N_19387,N_15949);
xor U28111 (N_28111,N_18874,N_12729);
nand U28112 (N_28112,N_17896,N_12180);
xor U28113 (N_28113,N_13020,N_10001);
xor U28114 (N_28114,N_12735,N_11257);
and U28115 (N_28115,N_11017,N_10544);
and U28116 (N_28116,N_13931,N_14254);
and U28117 (N_28117,N_16841,N_10562);
nor U28118 (N_28118,N_18076,N_14120);
nand U28119 (N_28119,N_14767,N_14546);
nor U28120 (N_28120,N_18995,N_18444);
or U28121 (N_28121,N_12683,N_17945);
and U28122 (N_28122,N_14546,N_18990);
or U28123 (N_28123,N_11690,N_14318);
and U28124 (N_28124,N_18647,N_15768);
nor U28125 (N_28125,N_19958,N_17744);
xor U28126 (N_28126,N_14765,N_16798);
xnor U28127 (N_28127,N_10162,N_11714);
xnor U28128 (N_28128,N_10572,N_10977);
xnor U28129 (N_28129,N_16039,N_13860);
xnor U28130 (N_28130,N_19355,N_16748);
xnor U28131 (N_28131,N_11388,N_11520);
xor U28132 (N_28132,N_18292,N_13583);
and U28133 (N_28133,N_15391,N_17641);
nor U28134 (N_28134,N_14471,N_19645);
xnor U28135 (N_28135,N_15721,N_11939);
and U28136 (N_28136,N_11947,N_13931);
and U28137 (N_28137,N_19329,N_13158);
or U28138 (N_28138,N_11672,N_11192);
nor U28139 (N_28139,N_10609,N_14404);
nand U28140 (N_28140,N_13217,N_17636);
nand U28141 (N_28141,N_12018,N_13401);
xnor U28142 (N_28142,N_17990,N_19715);
nor U28143 (N_28143,N_14098,N_11965);
and U28144 (N_28144,N_19497,N_14445);
or U28145 (N_28145,N_14428,N_10163);
or U28146 (N_28146,N_19282,N_13696);
xor U28147 (N_28147,N_19426,N_10119);
and U28148 (N_28148,N_16938,N_17932);
and U28149 (N_28149,N_14817,N_12596);
xor U28150 (N_28150,N_13981,N_11115);
xnor U28151 (N_28151,N_15831,N_13863);
nor U28152 (N_28152,N_15067,N_18161);
and U28153 (N_28153,N_14346,N_15041);
nor U28154 (N_28154,N_10493,N_12515);
nand U28155 (N_28155,N_12315,N_14452);
nor U28156 (N_28156,N_18298,N_13595);
nor U28157 (N_28157,N_14497,N_12419);
or U28158 (N_28158,N_16375,N_14073);
or U28159 (N_28159,N_17612,N_15700);
nand U28160 (N_28160,N_19053,N_14696);
or U28161 (N_28161,N_18968,N_11332);
or U28162 (N_28162,N_15870,N_14504);
xor U28163 (N_28163,N_19490,N_15899);
or U28164 (N_28164,N_13423,N_16578);
nor U28165 (N_28165,N_18206,N_13426);
nor U28166 (N_28166,N_17045,N_19553);
nand U28167 (N_28167,N_11504,N_13396);
and U28168 (N_28168,N_17472,N_16565);
or U28169 (N_28169,N_11783,N_19501);
nor U28170 (N_28170,N_11441,N_15757);
and U28171 (N_28171,N_19607,N_13463);
or U28172 (N_28172,N_12888,N_10178);
xor U28173 (N_28173,N_19249,N_18715);
nor U28174 (N_28174,N_12943,N_15378);
xor U28175 (N_28175,N_17335,N_15537);
or U28176 (N_28176,N_19107,N_11278);
and U28177 (N_28177,N_16859,N_15112);
or U28178 (N_28178,N_17218,N_18506);
xor U28179 (N_28179,N_12451,N_17605);
or U28180 (N_28180,N_19470,N_14451);
xor U28181 (N_28181,N_17955,N_17729);
nor U28182 (N_28182,N_15601,N_17278);
xor U28183 (N_28183,N_16733,N_19765);
nor U28184 (N_28184,N_18989,N_10746);
xnor U28185 (N_28185,N_15603,N_13677);
and U28186 (N_28186,N_10853,N_16943);
xnor U28187 (N_28187,N_15283,N_19414);
nor U28188 (N_28188,N_18628,N_14885);
or U28189 (N_28189,N_11191,N_14275);
nor U28190 (N_28190,N_11412,N_11440);
or U28191 (N_28191,N_11071,N_17710);
nor U28192 (N_28192,N_19763,N_12323);
nor U28193 (N_28193,N_11336,N_11413);
or U28194 (N_28194,N_19656,N_10885);
nand U28195 (N_28195,N_12015,N_19911);
and U28196 (N_28196,N_16866,N_16406);
nand U28197 (N_28197,N_13802,N_17615);
nand U28198 (N_28198,N_14328,N_11278);
nand U28199 (N_28199,N_12162,N_15430);
and U28200 (N_28200,N_10092,N_13115);
or U28201 (N_28201,N_18606,N_13018);
nand U28202 (N_28202,N_14432,N_14355);
nand U28203 (N_28203,N_10871,N_18267);
or U28204 (N_28204,N_10307,N_16404);
nand U28205 (N_28205,N_10004,N_11490);
nor U28206 (N_28206,N_17939,N_10973);
nor U28207 (N_28207,N_15278,N_19594);
xnor U28208 (N_28208,N_15289,N_10807);
nand U28209 (N_28209,N_16618,N_12707);
or U28210 (N_28210,N_13043,N_15635);
nor U28211 (N_28211,N_13478,N_13362);
xnor U28212 (N_28212,N_17215,N_17947);
and U28213 (N_28213,N_12776,N_18328);
nor U28214 (N_28214,N_15596,N_16003);
and U28215 (N_28215,N_16257,N_12069);
and U28216 (N_28216,N_13761,N_17299);
xor U28217 (N_28217,N_16979,N_14140);
and U28218 (N_28218,N_15654,N_11808);
or U28219 (N_28219,N_17702,N_11805);
xnor U28220 (N_28220,N_12393,N_14009);
nor U28221 (N_28221,N_12501,N_18976);
or U28222 (N_28222,N_13507,N_13473);
and U28223 (N_28223,N_14269,N_11034);
nor U28224 (N_28224,N_12638,N_18900);
and U28225 (N_28225,N_19982,N_17124);
nor U28226 (N_28226,N_18346,N_15394);
or U28227 (N_28227,N_11744,N_19764);
or U28228 (N_28228,N_15764,N_19379);
nor U28229 (N_28229,N_14941,N_11786);
and U28230 (N_28230,N_15619,N_17441);
or U28231 (N_28231,N_18364,N_19293);
and U28232 (N_28232,N_15756,N_12629);
or U28233 (N_28233,N_10065,N_12352);
xnor U28234 (N_28234,N_12148,N_12660);
or U28235 (N_28235,N_13254,N_19080);
xor U28236 (N_28236,N_12318,N_14524);
nand U28237 (N_28237,N_12005,N_17582);
xor U28238 (N_28238,N_16081,N_15469);
and U28239 (N_28239,N_17521,N_17397);
nand U28240 (N_28240,N_17286,N_11142);
xnor U28241 (N_28241,N_14659,N_12880);
nor U28242 (N_28242,N_14179,N_16596);
and U28243 (N_28243,N_12340,N_10363);
and U28244 (N_28244,N_12366,N_11459);
nor U28245 (N_28245,N_16419,N_18353);
xnor U28246 (N_28246,N_18137,N_17816);
or U28247 (N_28247,N_12087,N_10200);
nor U28248 (N_28248,N_19201,N_13985);
or U28249 (N_28249,N_13451,N_15207);
xor U28250 (N_28250,N_11145,N_16446);
and U28251 (N_28251,N_15789,N_11455);
nor U28252 (N_28252,N_14519,N_11190);
and U28253 (N_28253,N_13577,N_15938);
nor U28254 (N_28254,N_18200,N_19764);
or U28255 (N_28255,N_19606,N_15943);
nor U28256 (N_28256,N_16331,N_12534);
nand U28257 (N_28257,N_15559,N_14806);
xnor U28258 (N_28258,N_16137,N_14869);
nor U28259 (N_28259,N_18392,N_10621);
and U28260 (N_28260,N_13451,N_18205);
nor U28261 (N_28261,N_18238,N_19278);
or U28262 (N_28262,N_16191,N_14988);
and U28263 (N_28263,N_12678,N_13700);
nor U28264 (N_28264,N_19372,N_19003);
nor U28265 (N_28265,N_12862,N_17840);
and U28266 (N_28266,N_12243,N_10174);
nor U28267 (N_28267,N_16585,N_17505);
xnor U28268 (N_28268,N_18204,N_12202);
and U28269 (N_28269,N_18633,N_16722);
nor U28270 (N_28270,N_11979,N_18833);
nor U28271 (N_28271,N_13171,N_16417);
or U28272 (N_28272,N_17469,N_16493);
nand U28273 (N_28273,N_10856,N_16277);
or U28274 (N_28274,N_19544,N_11942);
and U28275 (N_28275,N_16152,N_18967);
xnor U28276 (N_28276,N_15263,N_16867);
nor U28277 (N_28277,N_13920,N_15871);
nand U28278 (N_28278,N_11820,N_18308);
xor U28279 (N_28279,N_14792,N_17155);
and U28280 (N_28280,N_18486,N_10875);
xor U28281 (N_28281,N_10035,N_19208);
or U28282 (N_28282,N_14124,N_19807);
nor U28283 (N_28283,N_19492,N_18150);
xor U28284 (N_28284,N_19865,N_16374);
nor U28285 (N_28285,N_10073,N_10293);
and U28286 (N_28286,N_10878,N_17427);
nand U28287 (N_28287,N_17521,N_13493);
or U28288 (N_28288,N_17087,N_16970);
and U28289 (N_28289,N_10777,N_12590);
or U28290 (N_28290,N_10640,N_11426);
nor U28291 (N_28291,N_10879,N_16137);
nand U28292 (N_28292,N_15966,N_10313);
nor U28293 (N_28293,N_16558,N_17155);
and U28294 (N_28294,N_10764,N_17873);
nor U28295 (N_28295,N_17695,N_13642);
nor U28296 (N_28296,N_11273,N_19987);
nor U28297 (N_28297,N_19760,N_12192);
nand U28298 (N_28298,N_10527,N_16466);
or U28299 (N_28299,N_17638,N_12559);
nor U28300 (N_28300,N_12689,N_17215);
xor U28301 (N_28301,N_10343,N_12759);
xor U28302 (N_28302,N_17554,N_17712);
and U28303 (N_28303,N_19138,N_19651);
xor U28304 (N_28304,N_10977,N_10578);
xnor U28305 (N_28305,N_12255,N_19617);
or U28306 (N_28306,N_19110,N_15295);
nor U28307 (N_28307,N_12957,N_16880);
nor U28308 (N_28308,N_18179,N_13482);
and U28309 (N_28309,N_17581,N_11013);
nand U28310 (N_28310,N_13445,N_15842);
nand U28311 (N_28311,N_13198,N_17009);
xnor U28312 (N_28312,N_11745,N_10536);
nand U28313 (N_28313,N_11041,N_19821);
nor U28314 (N_28314,N_10566,N_16937);
nor U28315 (N_28315,N_17347,N_18439);
nand U28316 (N_28316,N_13113,N_13273);
and U28317 (N_28317,N_13956,N_12606);
nand U28318 (N_28318,N_16961,N_14264);
xor U28319 (N_28319,N_12542,N_10291);
or U28320 (N_28320,N_14254,N_10410);
and U28321 (N_28321,N_12676,N_10833);
and U28322 (N_28322,N_14120,N_13230);
or U28323 (N_28323,N_13876,N_17905);
nand U28324 (N_28324,N_16905,N_10568);
nand U28325 (N_28325,N_10822,N_18379);
and U28326 (N_28326,N_17625,N_13085);
nor U28327 (N_28327,N_11703,N_11595);
nor U28328 (N_28328,N_12832,N_18677);
nand U28329 (N_28329,N_10793,N_19657);
and U28330 (N_28330,N_15532,N_12731);
or U28331 (N_28331,N_15579,N_19171);
and U28332 (N_28332,N_14706,N_14170);
xnor U28333 (N_28333,N_17782,N_18291);
nand U28334 (N_28334,N_10443,N_19513);
xnor U28335 (N_28335,N_19933,N_18185);
and U28336 (N_28336,N_17984,N_15689);
nand U28337 (N_28337,N_18064,N_16062);
xor U28338 (N_28338,N_13114,N_13863);
and U28339 (N_28339,N_12926,N_19159);
and U28340 (N_28340,N_19094,N_13177);
and U28341 (N_28341,N_14396,N_18219);
and U28342 (N_28342,N_15821,N_19807);
nor U28343 (N_28343,N_17937,N_19646);
or U28344 (N_28344,N_10377,N_15414);
nor U28345 (N_28345,N_15858,N_15713);
or U28346 (N_28346,N_13242,N_15954);
and U28347 (N_28347,N_12671,N_18243);
and U28348 (N_28348,N_13816,N_15898);
and U28349 (N_28349,N_18273,N_19070);
nand U28350 (N_28350,N_16997,N_11917);
or U28351 (N_28351,N_12638,N_11100);
or U28352 (N_28352,N_10646,N_11973);
or U28353 (N_28353,N_18712,N_11689);
and U28354 (N_28354,N_13039,N_12029);
nor U28355 (N_28355,N_14887,N_19045);
nor U28356 (N_28356,N_18759,N_19332);
or U28357 (N_28357,N_19738,N_13742);
or U28358 (N_28358,N_12082,N_12712);
xor U28359 (N_28359,N_17399,N_13772);
or U28360 (N_28360,N_19100,N_12917);
or U28361 (N_28361,N_16083,N_10644);
xnor U28362 (N_28362,N_17220,N_10002);
or U28363 (N_28363,N_15703,N_18788);
and U28364 (N_28364,N_10317,N_14891);
or U28365 (N_28365,N_13167,N_18296);
and U28366 (N_28366,N_18775,N_19407);
nor U28367 (N_28367,N_11362,N_14611);
nor U28368 (N_28368,N_19064,N_10084);
nor U28369 (N_28369,N_11845,N_11523);
and U28370 (N_28370,N_15826,N_14023);
nand U28371 (N_28371,N_19959,N_11436);
nand U28372 (N_28372,N_14203,N_15744);
xnor U28373 (N_28373,N_12661,N_11024);
and U28374 (N_28374,N_17443,N_10952);
or U28375 (N_28375,N_16500,N_14844);
nor U28376 (N_28376,N_15157,N_10551);
nand U28377 (N_28377,N_16945,N_13048);
and U28378 (N_28378,N_13891,N_16379);
nand U28379 (N_28379,N_10621,N_12100);
and U28380 (N_28380,N_13197,N_17136);
and U28381 (N_28381,N_11544,N_12674);
nand U28382 (N_28382,N_19824,N_15770);
or U28383 (N_28383,N_14359,N_19264);
xnor U28384 (N_28384,N_11098,N_11815);
nand U28385 (N_28385,N_16342,N_12863);
xor U28386 (N_28386,N_16191,N_15357);
and U28387 (N_28387,N_19349,N_18609);
nand U28388 (N_28388,N_14236,N_13141);
or U28389 (N_28389,N_19307,N_14639);
nand U28390 (N_28390,N_13018,N_17849);
xor U28391 (N_28391,N_19902,N_16725);
nand U28392 (N_28392,N_10741,N_19874);
and U28393 (N_28393,N_17444,N_10700);
nor U28394 (N_28394,N_16236,N_16947);
and U28395 (N_28395,N_14531,N_12070);
and U28396 (N_28396,N_12118,N_16225);
nand U28397 (N_28397,N_12439,N_10149);
nand U28398 (N_28398,N_19879,N_18148);
or U28399 (N_28399,N_17902,N_14826);
xor U28400 (N_28400,N_14957,N_10443);
xnor U28401 (N_28401,N_15366,N_13189);
nor U28402 (N_28402,N_12780,N_11027);
and U28403 (N_28403,N_15559,N_13077);
nor U28404 (N_28404,N_13154,N_13009);
nand U28405 (N_28405,N_19447,N_12745);
or U28406 (N_28406,N_13764,N_15578);
nand U28407 (N_28407,N_15571,N_10763);
xor U28408 (N_28408,N_16017,N_12725);
or U28409 (N_28409,N_18870,N_16366);
xor U28410 (N_28410,N_16062,N_15406);
nor U28411 (N_28411,N_13513,N_13164);
or U28412 (N_28412,N_16445,N_18304);
xor U28413 (N_28413,N_10746,N_15719);
and U28414 (N_28414,N_15372,N_12757);
nand U28415 (N_28415,N_16131,N_14019);
nor U28416 (N_28416,N_18225,N_16656);
nand U28417 (N_28417,N_19308,N_19154);
or U28418 (N_28418,N_10194,N_10682);
or U28419 (N_28419,N_17434,N_16738);
and U28420 (N_28420,N_12339,N_15140);
or U28421 (N_28421,N_13464,N_11312);
nand U28422 (N_28422,N_18708,N_19512);
or U28423 (N_28423,N_18805,N_19518);
xnor U28424 (N_28424,N_12728,N_19100);
or U28425 (N_28425,N_14790,N_19932);
xor U28426 (N_28426,N_13235,N_15588);
or U28427 (N_28427,N_17060,N_18749);
nand U28428 (N_28428,N_12816,N_16526);
and U28429 (N_28429,N_10954,N_15393);
nand U28430 (N_28430,N_11190,N_12659);
xnor U28431 (N_28431,N_11185,N_17584);
xor U28432 (N_28432,N_13702,N_12280);
nand U28433 (N_28433,N_13186,N_14542);
and U28434 (N_28434,N_17283,N_12044);
and U28435 (N_28435,N_16330,N_13223);
nand U28436 (N_28436,N_15072,N_15304);
xnor U28437 (N_28437,N_12194,N_16036);
nor U28438 (N_28438,N_16844,N_18446);
and U28439 (N_28439,N_11120,N_17001);
xor U28440 (N_28440,N_12182,N_10792);
nor U28441 (N_28441,N_16031,N_15516);
nor U28442 (N_28442,N_13503,N_16691);
and U28443 (N_28443,N_12071,N_11017);
and U28444 (N_28444,N_19305,N_13479);
xor U28445 (N_28445,N_17886,N_16443);
xnor U28446 (N_28446,N_19750,N_10062);
xnor U28447 (N_28447,N_11777,N_18550);
nand U28448 (N_28448,N_10973,N_17888);
xnor U28449 (N_28449,N_12342,N_17160);
nor U28450 (N_28450,N_19901,N_13892);
xor U28451 (N_28451,N_10537,N_11052);
nor U28452 (N_28452,N_10593,N_16171);
nor U28453 (N_28453,N_16305,N_15739);
and U28454 (N_28454,N_19711,N_17443);
nand U28455 (N_28455,N_17566,N_11443);
xnor U28456 (N_28456,N_10386,N_15784);
and U28457 (N_28457,N_19234,N_13493);
nor U28458 (N_28458,N_17269,N_10298);
and U28459 (N_28459,N_13887,N_18386);
nor U28460 (N_28460,N_19673,N_15312);
xnor U28461 (N_28461,N_13547,N_13751);
xor U28462 (N_28462,N_19630,N_17004);
or U28463 (N_28463,N_16360,N_11083);
xnor U28464 (N_28464,N_18358,N_11942);
nor U28465 (N_28465,N_16070,N_12464);
nand U28466 (N_28466,N_15206,N_13739);
nand U28467 (N_28467,N_18306,N_12778);
nor U28468 (N_28468,N_14113,N_11736);
xnor U28469 (N_28469,N_17880,N_14158);
xnor U28470 (N_28470,N_17934,N_19239);
and U28471 (N_28471,N_14506,N_19112);
nor U28472 (N_28472,N_18264,N_10075);
or U28473 (N_28473,N_12328,N_16043);
xor U28474 (N_28474,N_18960,N_12399);
nor U28475 (N_28475,N_13272,N_13384);
xnor U28476 (N_28476,N_11242,N_10123);
xnor U28477 (N_28477,N_10420,N_15742);
nor U28478 (N_28478,N_19392,N_10325);
or U28479 (N_28479,N_15491,N_18924);
nand U28480 (N_28480,N_13441,N_19078);
xor U28481 (N_28481,N_13040,N_18297);
and U28482 (N_28482,N_16107,N_12889);
or U28483 (N_28483,N_12523,N_18055);
or U28484 (N_28484,N_16284,N_11637);
or U28485 (N_28485,N_15874,N_12978);
nor U28486 (N_28486,N_14981,N_10912);
nor U28487 (N_28487,N_14339,N_10355);
nor U28488 (N_28488,N_16682,N_19878);
nor U28489 (N_28489,N_15686,N_16725);
nor U28490 (N_28490,N_10264,N_14393);
nor U28491 (N_28491,N_11462,N_10369);
and U28492 (N_28492,N_13421,N_13501);
nor U28493 (N_28493,N_13369,N_10290);
xnor U28494 (N_28494,N_19822,N_14273);
or U28495 (N_28495,N_12450,N_18985);
nor U28496 (N_28496,N_11699,N_10079);
xor U28497 (N_28497,N_18667,N_10723);
nand U28498 (N_28498,N_11322,N_10452);
nor U28499 (N_28499,N_10487,N_11483);
nor U28500 (N_28500,N_15990,N_13771);
nand U28501 (N_28501,N_18199,N_18143);
nor U28502 (N_28502,N_19708,N_14003);
or U28503 (N_28503,N_10651,N_10496);
or U28504 (N_28504,N_11025,N_19822);
nor U28505 (N_28505,N_11132,N_10985);
nand U28506 (N_28506,N_13982,N_15986);
nor U28507 (N_28507,N_11504,N_12086);
nor U28508 (N_28508,N_11412,N_17782);
xor U28509 (N_28509,N_18237,N_19231);
and U28510 (N_28510,N_12059,N_14897);
xnor U28511 (N_28511,N_19031,N_12683);
xnor U28512 (N_28512,N_14072,N_17695);
nand U28513 (N_28513,N_10700,N_14914);
and U28514 (N_28514,N_18232,N_15189);
or U28515 (N_28515,N_14590,N_15305);
nor U28516 (N_28516,N_12233,N_11219);
nor U28517 (N_28517,N_14272,N_16285);
or U28518 (N_28518,N_11621,N_14834);
nor U28519 (N_28519,N_15338,N_16406);
and U28520 (N_28520,N_13514,N_19433);
xor U28521 (N_28521,N_10060,N_14397);
xor U28522 (N_28522,N_15875,N_18894);
xor U28523 (N_28523,N_14694,N_19152);
xnor U28524 (N_28524,N_15272,N_14440);
or U28525 (N_28525,N_18752,N_14289);
and U28526 (N_28526,N_10282,N_12725);
nor U28527 (N_28527,N_12393,N_14929);
xor U28528 (N_28528,N_17589,N_16109);
and U28529 (N_28529,N_14278,N_14627);
xor U28530 (N_28530,N_11924,N_15906);
or U28531 (N_28531,N_14947,N_16689);
and U28532 (N_28532,N_11484,N_14975);
and U28533 (N_28533,N_13472,N_14026);
nand U28534 (N_28534,N_14941,N_15683);
nand U28535 (N_28535,N_19530,N_14235);
and U28536 (N_28536,N_14937,N_18939);
nor U28537 (N_28537,N_11670,N_18693);
nor U28538 (N_28538,N_19829,N_12589);
and U28539 (N_28539,N_14256,N_14912);
or U28540 (N_28540,N_15279,N_15110);
nand U28541 (N_28541,N_10539,N_14955);
nand U28542 (N_28542,N_16868,N_13652);
and U28543 (N_28543,N_17443,N_13632);
and U28544 (N_28544,N_19642,N_10273);
nand U28545 (N_28545,N_16680,N_18380);
nor U28546 (N_28546,N_18319,N_16618);
and U28547 (N_28547,N_12020,N_19496);
nand U28548 (N_28548,N_16874,N_13746);
and U28549 (N_28549,N_15918,N_19550);
nor U28550 (N_28550,N_11334,N_13908);
xnor U28551 (N_28551,N_15245,N_19327);
nor U28552 (N_28552,N_11146,N_15167);
xnor U28553 (N_28553,N_15078,N_14834);
xnor U28554 (N_28554,N_14122,N_15270);
nand U28555 (N_28555,N_19314,N_17063);
and U28556 (N_28556,N_12687,N_17099);
nor U28557 (N_28557,N_18983,N_17498);
xor U28558 (N_28558,N_12052,N_16063);
nand U28559 (N_28559,N_17132,N_11056);
nand U28560 (N_28560,N_10980,N_14471);
nor U28561 (N_28561,N_16012,N_15648);
and U28562 (N_28562,N_12766,N_17179);
nor U28563 (N_28563,N_10258,N_16637);
nand U28564 (N_28564,N_13183,N_10376);
xnor U28565 (N_28565,N_11989,N_16874);
nor U28566 (N_28566,N_18071,N_18245);
xor U28567 (N_28567,N_13419,N_10136);
xor U28568 (N_28568,N_17329,N_15278);
and U28569 (N_28569,N_13006,N_11916);
nor U28570 (N_28570,N_10283,N_13240);
and U28571 (N_28571,N_14085,N_18724);
xor U28572 (N_28572,N_13743,N_17760);
xnor U28573 (N_28573,N_18203,N_15429);
xnor U28574 (N_28574,N_19375,N_17677);
xnor U28575 (N_28575,N_18690,N_17109);
nand U28576 (N_28576,N_13231,N_19265);
and U28577 (N_28577,N_17962,N_12912);
nor U28578 (N_28578,N_11904,N_19724);
and U28579 (N_28579,N_12875,N_12836);
or U28580 (N_28580,N_14868,N_10284);
xnor U28581 (N_28581,N_18102,N_10476);
and U28582 (N_28582,N_16822,N_16418);
or U28583 (N_28583,N_13827,N_15156);
nor U28584 (N_28584,N_16708,N_12704);
or U28585 (N_28585,N_18490,N_12184);
or U28586 (N_28586,N_19505,N_11906);
nor U28587 (N_28587,N_19961,N_15280);
nand U28588 (N_28588,N_10665,N_11646);
nand U28589 (N_28589,N_15418,N_15751);
or U28590 (N_28590,N_17215,N_10631);
and U28591 (N_28591,N_18091,N_19259);
nor U28592 (N_28592,N_12952,N_12072);
nand U28593 (N_28593,N_17085,N_15688);
and U28594 (N_28594,N_10871,N_15424);
nand U28595 (N_28595,N_14377,N_13517);
nand U28596 (N_28596,N_10199,N_19642);
nor U28597 (N_28597,N_11993,N_18041);
or U28598 (N_28598,N_14009,N_11171);
or U28599 (N_28599,N_14720,N_19591);
or U28600 (N_28600,N_19410,N_11524);
nand U28601 (N_28601,N_16860,N_15724);
xor U28602 (N_28602,N_16732,N_16601);
and U28603 (N_28603,N_10368,N_17224);
nand U28604 (N_28604,N_10731,N_16519);
xnor U28605 (N_28605,N_15858,N_19656);
or U28606 (N_28606,N_10422,N_17880);
or U28607 (N_28607,N_17262,N_12286);
or U28608 (N_28608,N_13749,N_10117);
or U28609 (N_28609,N_11564,N_11409);
and U28610 (N_28610,N_17528,N_16172);
nand U28611 (N_28611,N_14596,N_10705);
nor U28612 (N_28612,N_12355,N_10394);
or U28613 (N_28613,N_15745,N_17701);
nand U28614 (N_28614,N_11928,N_11743);
and U28615 (N_28615,N_13525,N_18914);
and U28616 (N_28616,N_18584,N_18435);
and U28617 (N_28617,N_19356,N_11189);
and U28618 (N_28618,N_18016,N_16834);
nor U28619 (N_28619,N_18550,N_18313);
or U28620 (N_28620,N_19670,N_17214);
or U28621 (N_28621,N_14158,N_12516);
xnor U28622 (N_28622,N_16516,N_12896);
and U28623 (N_28623,N_12679,N_19715);
nand U28624 (N_28624,N_13793,N_10678);
and U28625 (N_28625,N_17780,N_15721);
and U28626 (N_28626,N_10898,N_13965);
and U28627 (N_28627,N_15010,N_19843);
xor U28628 (N_28628,N_19446,N_16982);
nor U28629 (N_28629,N_11275,N_18912);
nand U28630 (N_28630,N_14301,N_13030);
nor U28631 (N_28631,N_17865,N_17363);
nor U28632 (N_28632,N_11467,N_11381);
nand U28633 (N_28633,N_15987,N_18488);
nor U28634 (N_28634,N_12726,N_17084);
nand U28635 (N_28635,N_19742,N_10430);
xor U28636 (N_28636,N_10711,N_18717);
nand U28637 (N_28637,N_10376,N_16987);
or U28638 (N_28638,N_10933,N_17547);
or U28639 (N_28639,N_16322,N_13556);
or U28640 (N_28640,N_19779,N_11139);
nor U28641 (N_28641,N_10204,N_15501);
xor U28642 (N_28642,N_18982,N_15764);
nor U28643 (N_28643,N_14502,N_18466);
nand U28644 (N_28644,N_12677,N_17103);
xor U28645 (N_28645,N_16426,N_13500);
or U28646 (N_28646,N_10756,N_18084);
nand U28647 (N_28647,N_16047,N_19332);
nor U28648 (N_28648,N_19738,N_10100);
or U28649 (N_28649,N_19041,N_10725);
nand U28650 (N_28650,N_13548,N_15751);
or U28651 (N_28651,N_10104,N_10696);
nand U28652 (N_28652,N_12313,N_15722);
nor U28653 (N_28653,N_10498,N_12864);
and U28654 (N_28654,N_16702,N_13216);
xor U28655 (N_28655,N_13225,N_17846);
nand U28656 (N_28656,N_11222,N_17301);
nand U28657 (N_28657,N_17865,N_17068);
or U28658 (N_28658,N_19730,N_10278);
and U28659 (N_28659,N_11955,N_10394);
nor U28660 (N_28660,N_18526,N_15633);
and U28661 (N_28661,N_17968,N_11438);
xnor U28662 (N_28662,N_11486,N_19566);
nor U28663 (N_28663,N_18721,N_16151);
nand U28664 (N_28664,N_11810,N_10220);
and U28665 (N_28665,N_17454,N_15122);
xor U28666 (N_28666,N_14588,N_10201);
and U28667 (N_28667,N_18287,N_13562);
nor U28668 (N_28668,N_16454,N_11872);
or U28669 (N_28669,N_17911,N_17039);
nand U28670 (N_28670,N_10921,N_12555);
nand U28671 (N_28671,N_14731,N_14510);
nand U28672 (N_28672,N_19604,N_11545);
xor U28673 (N_28673,N_13111,N_12897);
nand U28674 (N_28674,N_16852,N_15141);
and U28675 (N_28675,N_16062,N_13561);
or U28676 (N_28676,N_15248,N_19898);
or U28677 (N_28677,N_19012,N_16042);
xnor U28678 (N_28678,N_16367,N_15393);
nand U28679 (N_28679,N_13526,N_13660);
nor U28680 (N_28680,N_13468,N_10522);
xnor U28681 (N_28681,N_14482,N_10483);
nand U28682 (N_28682,N_12628,N_18672);
and U28683 (N_28683,N_19023,N_13924);
and U28684 (N_28684,N_15068,N_10196);
or U28685 (N_28685,N_10574,N_13969);
or U28686 (N_28686,N_16392,N_14466);
xor U28687 (N_28687,N_11536,N_16387);
nor U28688 (N_28688,N_12401,N_11597);
or U28689 (N_28689,N_16808,N_19997);
nand U28690 (N_28690,N_17299,N_16152);
or U28691 (N_28691,N_15542,N_19830);
nor U28692 (N_28692,N_12423,N_16608);
nand U28693 (N_28693,N_17386,N_16291);
and U28694 (N_28694,N_17868,N_12850);
nand U28695 (N_28695,N_15528,N_14438);
and U28696 (N_28696,N_15756,N_10768);
nor U28697 (N_28697,N_10873,N_10054);
nor U28698 (N_28698,N_11729,N_10455);
xnor U28699 (N_28699,N_15604,N_11998);
and U28700 (N_28700,N_10265,N_16514);
nand U28701 (N_28701,N_19481,N_16914);
nand U28702 (N_28702,N_12698,N_12030);
xnor U28703 (N_28703,N_11101,N_15315);
and U28704 (N_28704,N_13491,N_12234);
nand U28705 (N_28705,N_17093,N_11030);
nor U28706 (N_28706,N_11279,N_16317);
xnor U28707 (N_28707,N_14615,N_11733);
or U28708 (N_28708,N_11254,N_13624);
or U28709 (N_28709,N_19868,N_16407);
xor U28710 (N_28710,N_15553,N_19939);
and U28711 (N_28711,N_16492,N_16001);
nand U28712 (N_28712,N_19058,N_10578);
and U28713 (N_28713,N_16397,N_13602);
xnor U28714 (N_28714,N_12710,N_16116);
xnor U28715 (N_28715,N_17287,N_10438);
and U28716 (N_28716,N_16390,N_15700);
nand U28717 (N_28717,N_10240,N_10811);
or U28718 (N_28718,N_17319,N_11602);
or U28719 (N_28719,N_13372,N_13722);
nor U28720 (N_28720,N_12235,N_12294);
xor U28721 (N_28721,N_14048,N_19768);
nor U28722 (N_28722,N_12378,N_15844);
and U28723 (N_28723,N_11385,N_14279);
xor U28724 (N_28724,N_13091,N_15772);
or U28725 (N_28725,N_13066,N_16774);
xnor U28726 (N_28726,N_16565,N_12142);
or U28727 (N_28727,N_13284,N_15354);
nand U28728 (N_28728,N_19823,N_18309);
nor U28729 (N_28729,N_11756,N_14060);
and U28730 (N_28730,N_13085,N_11703);
and U28731 (N_28731,N_14699,N_10657);
and U28732 (N_28732,N_19798,N_11419);
nand U28733 (N_28733,N_10994,N_13338);
nor U28734 (N_28734,N_12248,N_16787);
and U28735 (N_28735,N_10096,N_16257);
nor U28736 (N_28736,N_16954,N_12961);
and U28737 (N_28737,N_14884,N_17912);
or U28738 (N_28738,N_11379,N_17801);
xnor U28739 (N_28739,N_17767,N_15673);
nand U28740 (N_28740,N_13698,N_17415);
and U28741 (N_28741,N_19747,N_19791);
nor U28742 (N_28742,N_12290,N_13325);
or U28743 (N_28743,N_17277,N_14899);
and U28744 (N_28744,N_14833,N_15807);
and U28745 (N_28745,N_11607,N_17230);
or U28746 (N_28746,N_12603,N_18161);
nor U28747 (N_28747,N_16172,N_10659);
xor U28748 (N_28748,N_13944,N_13316);
nor U28749 (N_28749,N_19486,N_11679);
nor U28750 (N_28750,N_17620,N_19655);
xnor U28751 (N_28751,N_19804,N_14422);
nor U28752 (N_28752,N_17373,N_18910);
or U28753 (N_28753,N_10151,N_10404);
xnor U28754 (N_28754,N_17520,N_14369);
xor U28755 (N_28755,N_19492,N_12870);
xnor U28756 (N_28756,N_11837,N_10555);
nor U28757 (N_28757,N_14311,N_15062);
and U28758 (N_28758,N_11453,N_17272);
and U28759 (N_28759,N_13288,N_12102);
nor U28760 (N_28760,N_18399,N_18034);
and U28761 (N_28761,N_12525,N_19116);
nor U28762 (N_28762,N_19144,N_15435);
or U28763 (N_28763,N_18352,N_18417);
nand U28764 (N_28764,N_10957,N_17419);
xor U28765 (N_28765,N_14145,N_19355);
xnor U28766 (N_28766,N_19130,N_10957);
nand U28767 (N_28767,N_16932,N_14497);
and U28768 (N_28768,N_13959,N_15889);
nand U28769 (N_28769,N_13999,N_15965);
xnor U28770 (N_28770,N_16482,N_16933);
and U28771 (N_28771,N_16787,N_10839);
xnor U28772 (N_28772,N_14936,N_15995);
xnor U28773 (N_28773,N_11897,N_16344);
nor U28774 (N_28774,N_16063,N_15577);
nand U28775 (N_28775,N_15341,N_12643);
xor U28776 (N_28776,N_19481,N_16288);
xnor U28777 (N_28777,N_19549,N_15315);
and U28778 (N_28778,N_15959,N_12692);
xor U28779 (N_28779,N_17145,N_19232);
nor U28780 (N_28780,N_10436,N_15477);
or U28781 (N_28781,N_13259,N_17978);
or U28782 (N_28782,N_18790,N_11638);
xor U28783 (N_28783,N_11688,N_11898);
or U28784 (N_28784,N_10782,N_14000);
nand U28785 (N_28785,N_17852,N_19717);
nor U28786 (N_28786,N_17385,N_10188);
and U28787 (N_28787,N_17907,N_10266);
or U28788 (N_28788,N_16941,N_12746);
nor U28789 (N_28789,N_14287,N_10010);
nor U28790 (N_28790,N_11303,N_11163);
and U28791 (N_28791,N_13288,N_14910);
nand U28792 (N_28792,N_18542,N_10018);
xnor U28793 (N_28793,N_13050,N_12824);
nor U28794 (N_28794,N_15017,N_12333);
xor U28795 (N_28795,N_15760,N_10981);
nand U28796 (N_28796,N_15585,N_18612);
or U28797 (N_28797,N_13187,N_14965);
nor U28798 (N_28798,N_16664,N_10507);
nand U28799 (N_28799,N_18057,N_11909);
nor U28800 (N_28800,N_10073,N_15539);
or U28801 (N_28801,N_17733,N_10798);
or U28802 (N_28802,N_12375,N_16565);
nand U28803 (N_28803,N_18317,N_15917);
xnor U28804 (N_28804,N_17516,N_13837);
or U28805 (N_28805,N_11056,N_15889);
or U28806 (N_28806,N_13631,N_15543);
or U28807 (N_28807,N_10440,N_18492);
and U28808 (N_28808,N_18700,N_18406);
or U28809 (N_28809,N_17325,N_15644);
or U28810 (N_28810,N_14764,N_12188);
and U28811 (N_28811,N_15278,N_18692);
nor U28812 (N_28812,N_12416,N_14291);
xnor U28813 (N_28813,N_15236,N_19072);
and U28814 (N_28814,N_18605,N_15925);
nor U28815 (N_28815,N_18199,N_19388);
xor U28816 (N_28816,N_10626,N_14885);
and U28817 (N_28817,N_11692,N_15626);
xnor U28818 (N_28818,N_14692,N_13748);
nor U28819 (N_28819,N_10023,N_12690);
nand U28820 (N_28820,N_18318,N_16373);
and U28821 (N_28821,N_16624,N_19375);
and U28822 (N_28822,N_19206,N_19174);
nor U28823 (N_28823,N_10554,N_17342);
xnor U28824 (N_28824,N_18705,N_19403);
and U28825 (N_28825,N_13331,N_10850);
or U28826 (N_28826,N_11762,N_15446);
nor U28827 (N_28827,N_12909,N_19727);
and U28828 (N_28828,N_18730,N_18527);
nand U28829 (N_28829,N_15668,N_13185);
nand U28830 (N_28830,N_11186,N_18034);
nand U28831 (N_28831,N_14972,N_12343);
and U28832 (N_28832,N_10394,N_12801);
xnor U28833 (N_28833,N_10517,N_10999);
or U28834 (N_28834,N_11852,N_18193);
nand U28835 (N_28835,N_14558,N_14298);
xnor U28836 (N_28836,N_18016,N_12047);
xor U28837 (N_28837,N_17655,N_12213);
xnor U28838 (N_28838,N_10152,N_13316);
or U28839 (N_28839,N_13970,N_11101);
xnor U28840 (N_28840,N_13952,N_12525);
and U28841 (N_28841,N_19268,N_11779);
and U28842 (N_28842,N_15503,N_19199);
nand U28843 (N_28843,N_12038,N_18384);
and U28844 (N_28844,N_14389,N_17014);
and U28845 (N_28845,N_19638,N_18044);
nor U28846 (N_28846,N_11182,N_19142);
and U28847 (N_28847,N_12957,N_14611);
xnor U28848 (N_28848,N_12163,N_15295);
xor U28849 (N_28849,N_15749,N_12407);
nand U28850 (N_28850,N_10321,N_13789);
and U28851 (N_28851,N_19669,N_15239);
and U28852 (N_28852,N_18624,N_12043);
nor U28853 (N_28853,N_13381,N_13485);
xnor U28854 (N_28854,N_13838,N_13529);
xnor U28855 (N_28855,N_18037,N_10960);
or U28856 (N_28856,N_12721,N_16129);
and U28857 (N_28857,N_16892,N_12590);
or U28858 (N_28858,N_11056,N_11555);
nor U28859 (N_28859,N_18545,N_19480);
or U28860 (N_28860,N_17371,N_11345);
and U28861 (N_28861,N_18777,N_19668);
nor U28862 (N_28862,N_19662,N_16612);
nor U28863 (N_28863,N_19703,N_11798);
or U28864 (N_28864,N_19917,N_12444);
and U28865 (N_28865,N_19857,N_18253);
xor U28866 (N_28866,N_17733,N_16765);
nand U28867 (N_28867,N_11784,N_17827);
or U28868 (N_28868,N_17698,N_12694);
nand U28869 (N_28869,N_10518,N_18000);
and U28870 (N_28870,N_17012,N_18202);
xnor U28871 (N_28871,N_12253,N_18207);
nand U28872 (N_28872,N_10093,N_10555);
and U28873 (N_28873,N_15469,N_18970);
nor U28874 (N_28874,N_13116,N_11108);
nor U28875 (N_28875,N_19774,N_10084);
or U28876 (N_28876,N_14337,N_19044);
or U28877 (N_28877,N_13998,N_15328);
and U28878 (N_28878,N_13425,N_12663);
and U28879 (N_28879,N_15948,N_16027);
nand U28880 (N_28880,N_13918,N_13525);
or U28881 (N_28881,N_12267,N_19506);
xnor U28882 (N_28882,N_11672,N_16628);
xor U28883 (N_28883,N_15035,N_12482);
or U28884 (N_28884,N_19210,N_11699);
nand U28885 (N_28885,N_16961,N_17775);
nand U28886 (N_28886,N_12861,N_12068);
or U28887 (N_28887,N_14636,N_19262);
xnor U28888 (N_28888,N_13917,N_18022);
and U28889 (N_28889,N_18907,N_11693);
xnor U28890 (N_28890,N_11543,N_10678);
and U28891 (N_28891,N_16673,N_12394);
and U28892 (N_28892,N_13603,N_11752);
nor U28893 (N_28893,N_12405,N_14319);
and U28894 (N_28894,N_14224,N_11152);
nor U28895 (N_28895,N_14055,N_13987);
xnor U28896 (N_28896,N_13020,N_11811);
or U28897 (N_28897,N_13809,N_12453);
nand U28898 (N_28898,N_15290,N_17460);
nand U28899 (N_28899,N_17452,N_17638);
or U28900 (N_28900,N_12976,N_18952);
nor U28901 (N_28901,N_10003,N_14644);
or U28902 (N_28902,N_12395,N_10411);
xnor U28903 (N_28903,N_10204,N_11435);
or U28904 (N_28904,N_12245,N_16439);
or U28905 (N_28905,N_15289,N_17835);
nand U28906 (N_28906,N_12026,N_14003);
nor U28907 (N_28907,N_15239,N_18580);
xnor U28908 (N_28908,N_19820,N_19813);
or U28909 (N_28909,N_11898,N_19662);
nand U28910 (N_28910,N_16368,N_15571);
or U28911 (N_28911,N_17482,N_11884);
and U28912 (N_28912,N_15646,N_12163);
or U28913 (N_28913,N_16823,N_13198);
nor U28914 (N_28914,N_15011,N_12704);
or U28915 (N_28915,N_15717,N_14725);
and U28916 (N_28916,N_17266,N_12450);
nand U28917 (N_28917,N_14491,N_13450);
nor U28918 (N_28918,N_13712,N_15525);
nand U28919 (N_28919,N_13599,N_17583);
xor U28920 (N_28920,N_16847,N_11514);
and U28921 (N_28921,N_14950,N_10361);
or U28922 (N_28922,N_19250,N_15743);
and U28923 (N_28923,N_18348,N_18958);
xnor U28924 (N_28924,N_16105,N_13392);
nor U28925 (N_28925,N_18930,N_13492);
nor U28926 (N_28926,N_14883,N_17520);
or U28927 (N_28927,N_11615,N_12075);
nor U28928 (N_28928,N_14728,N_19843);
or U28929 (N_28929,N_10978,N_19018);
or U28930 (N_28930,N_14278,N_10995);
or U28931 (N_28931,N_12924,N_15368);
nor U28932 (N_28932,N_11948,N_10395);
and U28933 (N_28933,N_18843,N_11756);
nand U28934 (N_28934,N_10327,N_11358);
nor U28935 (N_28935,N_17069,N_19874);
or U28936 (N_28936,N_13465,N_13252);
xor U28937 (N_28937,N_17874,N_19880);
xnor U28938 (N_28938,N_12052,N_15511);
and U28939 (N_28939,N_11622,N_10852);
and U28940 (N_28940,N_18970,N_15024);
or U28941 (N_28941,N_16044,N_17814);
nor U28942 (N_28942,N_14377,N_15505);
nor U28943 (N_28943,N_12557,N_17139);
or U28944 (N_28944,N_14151,N_13317);
or U28945 (N_28945,N_10694,N_11195);
nor U28946 (N_28946,N_10956,N_14511);
xor U28947 (N_28947,N_10650,N_17277);
xnor U28948 (N_28948,N_17036,N_18742);
nor U28949 (N_28949,N_15786,N_15007);
xor U28950 (N_28950,N_17057,N_15408);
or U28951 (N_28951,N_18430,N_16176);
or U28952 (N_28952,N_16069,N_18214);
nor U28953 (N_28953,N_16373,N_16362);
xor U28954 (N_28954,N_12808,N_17667);
nor U28955 (N_28955,N_17921,N_15706);
xnor U28956 (N_28956,N_10748,N_11572);
or U28957 (N_28957,N_19605,N_16253);
nor U28958 (N_28958,N_16642,N_10395);
nor U28959 (N_28959,N_18035,N_13761);
nor U28960 (N_28960,N_16044,N_17728);
xor U28961 (N_28961,N_16261,N_14523);
and U28962 (N_28962,N_10941,N_11637);
and U28963 (N_28963,N_12896,N_10653);
or U28964 (N_28964,N_18312,N_13094);
nand U28965 (N_28965,N_19132,N_16383);
xor U28966 (N_28966,N_12198,N_13085);
nand U28967 (N_28967,N_14807,N_13592);
nand U28968 (N_28968,N_16144,N_13019);
or U28969 (N_28969,N_19233,N_16188);
xnor U28970 (N_28970,N_14835,N_12535);
and U28971 (N_28971,N_13314,N_13556);
or U28972 (N_28972,N_14301,N_14055);
and U28973 (N_28973,N_13451,N_18353);
nor U28974 (N_28974,N_18156,N_19924);
nor U28975 (N_28975,N_16809,N_16987);
xnor U28976 (N_28976,N_15751,N_13611);
nand U28977 (N_28977,N_13674,N_12318);
nor U28978 (N_28978,N_16048,N_12888);
nor U28979 (N_28979,N_15413,N_16377);
xor U28980 (N_28980,N_10366,N_12010);
and U28981 (N_28981,N_19219,N_12533);
and U28982 (N_28982,N_18158,N_18428);
nor U28983 (N_28983,N_16395,N_15888);
and U28984 (N_28984,N_16413,N_17592);
nor U28985 (N_28985,N_11273,N_18453);
and U28986 (N_28986,N_14217,N_16812);
and U28987 (N_28987,N_16757,N_19482);
and U28988 (N_28988,N_16301,N_18687);
nor U28989 (N_28989,N_17849,N_12196);
nor U28990 (N_28990,N_16300,N_18271);
or U28991 (N_28991,N_10949,N_17143);
nand U28992 (N_28992,N_16655,N_13800);
or U28993 (N_28993,N_14476,N_17602);
or U28994 (N_28994,N_13168,N_11580);
nor U28995 (N_28995,N_10763,N_19314);
xnor U28996 (N_28996,N_12542,N_14014);
or U28997 (N_28997,N_10623,N_16441);
or U28998 (N_28998,N_13054,N_18897);
nor U28999 (N_28999,N_10460,N_12796);
nor U29000 (N_29000,N_10438,N_16019);
xnor U29001 (N_29001,N_18831,N_10557);
or U29002 (N_29002,N_19602,N_13505);
or U29003 (N_29003,N_17556,N_12756);
xnor U29004 (N_29004,N_11111,N_18752);
and U29005 (N_29005,N_17865,N_12545);
or U29006 (N_29006,N_15532,N_12750);
xnor U29007 (N_29007,N_12512,N_18687);
nand U29008 (N_29008,N_11250,N_19742);
nand U29009 (N_29009,N_10183,N_18095);
or U29010 (N_29010,N_11859,N_10094);
nor U29011 (N_29011,N_19798,N_19151);
nand U29012 (N_29012,N_17601,N_17642);
xnor U29013 (N_29013,N_10754,N_12846);
and U29014 (N_29014,N_17450,N_11626);
or U29015 (N_29015,N_15966,N_10370);
nand U29016 (N_29016,N_17551,N_19295);
or U29017 (N_29017,N_10347,N_15528);
or U29018 (N_29018,N_15122,N_18826);
xor U29019 (N_29019,N_13304,N_16766);
nor U29020 (N_29020,N_13004,N_11795);
xor U29021 (N_29021,N_15899,N_13816);
nand U29022 (N_29022,N_14752,N_17304);
nand U29023 (N_29023,N_15572,N_12625);
xnor U29024 (N_29024,N_17401,N_16485);
nand U29025 (N_29025,N_12775,N_17493);
nor U29026 (N_29026,N_18154,N_13738);
nor U29027 (N_29027,N_11100,N_13201);
and U29028 (N_29028,N_11913,N_17537);
or U29029 (N_29029,N_11452,N_17210);
xnor U29030 (N_29030,N_14579,N_14362);
nand U29031 (N_29031,N_18611,N_15758);
and U29032 (N_29032,N_13983,N_11668);
and U29033 (N_29033,N_12069,N_17627);
xor U29034 (N_29034,N_11505,N_17487);
or U29035 (N_29035,N_10110,N_12650);
or U29036 (N_29036,N_19310,N_16607);
and U29037 (N_29037,N_16344,N_19473);
nand U29038 (N_29038,N_17668,N_11656);
or U29039 (N_29039,N_12654,N_12016);
xor U29040 (N_29040,N_12692,N_13964);
nor U29041 (N_29041,N_19385,N_16399);
nor U29042 (N_29042,N_18989,N_15181);
and U29043 (N_29043,N_18744,N_10680);
xor U29044 (N_29044,N_13062,N_17095);
nand U29045 (N_29045,N_11293,N_10908);
nor U29046 (N_29046,N_17822,N_10443);
or U29047 (N_29047,N_10676,N_11957);
or U29048 (N_29048,N_14070,N_10564);
or U29049 (N_29049,N_13382,N_10310);
and U29050 (N_29050,N_13940,N_17013);
nor U29051 (N_29051,N_11103,N_10955);
nand U29052 (N_29052,N_18091,N_12221);
nand U29053 (N_29053,N_17488,N_13687);
xnor U29054 (N_29054,N_16883,N_19682);
or U29055 (N_29055,N_12319,N_10162);
or U29056 (N_29056,N_12695,N_12789);
or U29057 (N_29057,N_17663,N_10620);
nand U29058 (N_29058,N_11410,N_10390);
and U29059 (N_29059,N_17854,N_14042);
nor U29060 (N_29060,N_15938,N_10160);
or U29061 (N_29061,N_18630,N_19907);
nor U29062 (N_29062,N_16679,N_15509);
nand U29063 (N_29063,N_19372,N_19912);
or U29064 (N_29064,N_16627,N_16716);
xor U29065 (N_29065,N_10096,N_14655);
nor U29066 (N_29066,N_17581,N_11259);
xnor U29067 (N_29067,N_12229,N_14142);
nor U29068 (N_29068,N_15590,N_11999);
or U29069 (N_29069,N_13758,N_10097);
xnor U29070 (N_29070,N_10133,N_10226);
and U29071 (N_29071,N_17794,N_19923);
or U29072 (N_29072,N_16911,N_15680);
or U29073 (N_29073,N_13983,N_10241);
nor U29074 (N_29074,N_14225,N_15320);
nor U29075 (N_29075,N_16824,N_16722);
xor U29076 (N_29076,N_19808,N_16934);
and U29077 (N_29077,N_17799,N_14306);
or U29078 (N_29078,N_13297,N_19015);
or U29079 (N_29079,N_16262,N_14959);
xor U29080 (N_29080,N_10630,N_16128);
nand U29081 (N_29081,N_14363,N_14468);
xor U29082 (N_29082,N_17637,N_16829);
nand U29083 (N_29083,N_16017,N_18710);
nor U29084 (N_29084,N_18224,N_13135);
and U29085 (N_29085,N_17032,N_18627);
and U29086 (N_29086,N_17528,N_15075);
nor U29087 (N_29087,N_11701,N_14074);
nand U29088 (N_29088,N_11701,N_11587);
or U29089 (N_29089,N_14730,N_15313);
and U29090 (N_29090,N_12715,N_15058);
or U29091 (N_29091,N_14466,N_18674);
nor U29092 (N_29092,N_14049,N_11844);
xor U29093 (N_29093,N_12741,N_10442);
xnor U29094 (N_29094,N_15933,N_12033);
xnor U29095 (N_29095,N_15502,N_15983);
nor U29096 (N_29096,N_14147,N_17533);
nor U29097 (N_29097,N_13495,N_19279);
xor U29098 (N_29098,N_17675,N_12522);
xnor U29099 (N_29099,N_13835,N_17431);
and U29100 (N_29100,N_10058,N_12929);
xor U29101 (N_29101,N_10454,N_19029);
xor U29102 (N_29102,N_10528,N_11949);
xor U29103 (N_29103,N_15291,N_11619);
or U29104 (N_29104,N_10328,N_12172);
or U29105 (N_29105,N_11050,N_11429);
nand U29106 (N_29106,N_15381,N_13318);
and U29107 (N_29107,N_15003,N_13633);
and U29108 (N_29108,N_19429,N_14649);
or U29109 (N_29109,N_11686,N_13474);
nor U29110 (N_29110,N_18956,N_17395);
or U29111 (N_29111,N_18211,N_17944);
nand U29112 (N_29112,N_14701,N_13629);
xor U29113 (N_29113,N_11036,N_18625);
nand U29114 (N_29114,N_11273,N_14544);
xnor U29115 (N_29115,N_17766,N_19262);
nand U29116 (N_29116,N_19845,N_17699);
and U29117 (N_29117,N_16985,N_15920);
and U29118 (N_29118,N_18507,N_10942);
and U29119 (N_29119,N_18543,N_17909);
nor U29120 (N_29120,N_15197,N_11015);
nand U29121 (N_29121,N_19791,N_14068);
nor U29122 (N_29122,N_16924,N_10659);
nor U29123 (N_29123,N_12605,N_14780);
nor U29124 (N_29124,N_15858,N_15259);
or U29125 (N_29125,N_12923,N_14108);
nor U29126 (N_29126,N_12425,N_15305);
and U29127 (N_29127,N_15954,N_18645);
nor U29128 (N_29128,N_11580,N_11818);
nor U29129 (N_29129,N_19929,N_14462);
xnor U29130 (N_29130,N_13150,N_11555);
xnor U29131 (N_29131,N_13057,N_16314);
nand U29132 (N_29132,N_19381,N_13272);
and U29133 (N_29133,N_10778,N_14993);
and U29134 (N_29134,N_19766,N_15704);
and U29135 (N_29135,N_16432,N_16221);
nor U29136 (N_29136,N_10790,N_10921);
nand U29137 (N_29137,N_19268,N_13686);
nand U29138 (N_29138,N_19359,N_16187);
or U29139 (N_29139,N_11222,N_11289);
nor U29140 (N_29140,N_13888,N_16975);
or U29141 (N_29141,N_19249,N_12665);
xnor U29142 (N_29142,N_17861,N_14699);
and U29143 (N_29143,N_11493,N_11311);
nand U29144 (N_29144,N_11921,N_19168);
nand U29145 (N_29145,N_13193,N_14216);
and U29146 (N_29146,N_10704,N_10811);
or U29147 (N_29147,N_17814,N_13379);
and U29148 (N_29148,N_14871,N_10426);
and U29149 (N_29149,N_11096,N_15884);
nand U29150 (N_29150,N_15972,N_15552);
xnor U29151 (N_29151,N_11432,N_15145);
and U29152 (N_29152,N_16651,N_11929);
xor U29153 (N_29153,N_17615,N_17219);
xor U29154 (N_29154,N_15021,N_10361);
nand U29155 (N_29155,N_16541,N_12266);
nand U29156 (N_29156,N_18378,N_15863);
nand U29157 (N_29157,N_10864,N_16818);
nand U29158 (N_29158,N_14027,N_12791);
nand U29159 (N_29159,N_16594,N_12534);
and U29160 (N_29160,N_16585,N_19037);
nand U29161 (N_29161,N_11073,N_18617);
xnor U29162 (N_29162,N_12242,N_10181);
and U29163 (N_29163,N_16182,N_16567);
and U29164 (N_29164,N_16665,N_12381);
xor U29165 (N_29165,N_10673,N_17358);
and U29166 (N_29166,N_12603,N_10375);
nor U29167 (N_29167,N_19608,N_16856);
and U29168 (N_29168,N_13373,N_12043);
and U29169 (N_29169,N_12705,N_13473);
or U29170 (N_29170,N_15813,N_11395);
nand U29171 (N_29171,N_15055,N_12750);
nand U29172 (N_29172,N_11789,N_12561);
and U29173 (N_29173,N_18528,N_14862);
nor U29174 (N_29174,N_12908,N_14530);
nand U29175 (N_29175,N_13190,N_18875);
and U29176 (N_29176,N_14334,N_13779);
and U29177 (N_29177,N_13101,N_18082);
and U29178 (N_29178,N_19149,N_17314);
xnor U29179 (N_29179,N_16233,N_13526);
xnor U29180 (N_29180,N_10571,N_17981);
nor U29181 (N_29181,N_18556,N_12340);
or U29182 (N_29182,N_10758,N_16684);
nor U29183 (N_29183,N_15948,N_12337);
nor U29184 (N_29184,N_12894,N_15118);
and U29185 (N_29185,N_17488,N_17450);
and U29186 (N_29186,N_17031,N_15309);
or U29187 (N_29187,N_17627,N_11683);
nand U29188 (N_29188,N_15272,N_17193);
nor U29189 (N_29189,N_10107,N_12201);
or U29190 (N_29190,N_15458,N_12101);
and U29191 (N_29191,N_19587,N_10129);
and U29192 (N_29192,N_12700,N_17972);
nor U29193 (N_29193,N_13586,N_11201);
nor U29194 (N_29194,N_16059,N_18888);
or U29195 (N_29195,N_13138,N_15549);
or U29196 (N_29196,N_17727,N_13617);
or U29197 (N_29197,N_11310,N_11613);
xnor U29198 (N_29198,N_15671,N_14612);
or U29199 (N_29199,N_11842,N_16382);
nand U29200 (N_29200,N_11683,N_14100);
nor U29201 (N_29201,N_15817,N_15077);
and U29202 (N_29202,N_13943,N_18047);
and U29203 (N_29203,N_13699,N_16600);
xnor U29204 (N_29204,N_11743,N_14691);
and U29205 (N_29205,N_15702,N_17378);
nor U29206 (N_29206,N_16063,N_18158);
or U29207 (N_29207,N_13259,N_19095);
or U29208 (N_29208,N_11027,N_13629);
or U29209 (N_29209,N_18258,N_14426);
nor U29210 (N_29210,N_16712,N_10310);
nor U29211 (N_29211,N_12964,N_15911);
and U29212 (N_29212,N_19867,N_14676);
xor U29213 (N_29213,N_14438,N_15001);
or U29214 (N_29214,N_19002,N_11037);
or U29215 (N_29215,N_14786,N_13394);
or U29216 (N_29216,N_11212,N_13924);
or U29217 (N_29217,N_12983,N_19821);
and U29218 (N_29218,N_17328,N_13353);
and U29219 (N_29219,N_16469,N_13233);
and U29220 (N_29220,N_14075,N_17623);
and U29221 (N_29221,N_19638,N_16351);
or U29222 (N_29222,N_12617,N_17590);
and U29223 (N_29223,N_15644,N_19542);
xor U29224 (N_29224,N_16878,N_15059);
or U29225 (N_29225,N_14999,N_15535);
and U29226 (N_29226,N_11478,N_18332);
xor U29227 (N_29227,N_14914,N_13872);
or U29228 (N_29228,N_10378,N_13990);
or U29229 (N_29229,N_19350,N_14088);
nand U29230 (N_29230,N_14805,N_19336);
or U29231 (N_29231,N_18850,N_15379);
xor U29232 (N_29232,N_19855,N_18009);
nand U29233 (N_29233,N_11732,N_11709);
and U29234 (N_29234,N_18460,N_11763);
xor U29235 (N_29235,N_10527,N_10951);
xor U29236 (N_29236,N_12824,N_18079);
and U29237 (N_29237,N_19810,N_17898);
and U29238 (N_29238,N_11548,N_19146);
or U29239 (N_29239,N_15590,N_16318);
xor U29240 (N_29240,N_18209,N_18042);
nand U29241 (N_29241,N_10116,N_15056);
or U29242 (N_29242,N_12971,N_16605);
nand U29243 (N_29243,N_15266,N_14021);
and U29244 (N_29244,N_11965,N_12163);
and U29245 (N_29245,N_19829,N_19648);
or U29246 (N_29246,N_15314,N_12841);
nand U29247 (N_29247,N_10387,N_13115);
nand U29248 (N_29248,N_13675,N_16445);
nand U29249 (N_29249,N_11111,N_19630);
nor U29250 (N_29250,N_15131,N_14944);
and U29251 (N_29251,N_17654,N_16729);
nor U29252 (N_29252,N_14579,N_15038);
nand U29253 (N_29253,N_12559,N_18869);
xor U29254 (N_29254,N_10353,N_13161);
or U29255 (N_29255,N_18790,N_13480);
nor U29256 (N_29256,N_11641,N_18221);
or U29257 (N_29257,N_12523,N_12365);
nor U29258 (N_29258,N_16481,N_13123);
and U29259 (N_29259,N_10106,N_19298);
xor U29260 (N_29260,N_15207,N_10165);
nor U29261 (N_29261,N_12731,N_18511);
or U29262 (N_29262,N_19689,N_16251);
and U29263 (N_29263,N_17337,N_19316);
xor U29264 (N_29264,N_14844,N_18068);
and U29265 (N_29265,N_12775,N_14437);
xor U29266 (N_29266,N_13743,N_19283);
nor U29267 (N_29267,N_14492,N_11252);
nor U29268 (N_29268,N_18824,N_17983);
nor U29269 (N_29269,N_17648,N_12953);
nor U29270 (N_29270,N_10691,N_18175);
xnor U29271 (N_29271,N_12205,N_12732);
xor U29272 (N_29272,N_18333,N_15894);
nor U29273 (N_29273,N_15318,N_12923);
or U29274 (N_29274,N_11824,N_11838);
or U29275 (N_29275,N_17579,N_18172);
or U29276 (N_29276,N_15866,N_19359);
nand U29277 (N_29277,N_19991,N_18073);
and U29278 (N_29278,N_14138,N_13444);
nor U29279 (N_29279,N_14999,N_12785);
nor U29280 (N_29280,N_14709,N_10254);
or U29281 (N_29281,N_19063,N_12135);
nor U29282 (N_29282,N_16913,N_11271);
and U29283 (N_29283,N_11498,N_10265);
nand U29284 (N_29284,N_16689,N_13989);
xor U29285 (N_29285,N_17175,N_19418);
nor U29286 (N_29286,N_19517,N_10227);
or U29287 (N_29287,N_17348,N_12647);
and U29288 (N_29288,N_10075,N_10449);
nand U29289 (N_29289,N_13465,N_19240);
and U29290 (N_29290,N_19034,N_11685);
and U29291 (N_29291,N_11082,N_13581);
nor U29292 (N_29292,N_19224,N_19211);
nor U29293 (N_29293,N_19091,N_14387);
or U29294 (N_29294,N_11775,N_17465);
and U29295 (N_29295,N_10116,N_16773);
or U29296 (N_29296,N_13842,N_18070);
nor U29297 (N_29297,N_17943,N_16259);
nand U29298 (N_29298,N_19741,N_10367);
and U29299 (N_29299,N_10663,N_14667);
or U29300 (N_29300,N_11318,N_14895);
and U29301 (N_29301,N_11657,N_11120);
or U29302 (N_29302,N_14632,N_13010);
nor U29303 (N_29303,N_15937,N_11217);
nor U29304 (N_29304,N_10013,N_17613);
nand U29305 (N_29305,N_11366,N_11544);
or U29306 (N_29306,N_12527,N_11177);
xor U29307 (N_29307,N_16935,N_18568);
nor U29308 (N_29308,N_16347,N_16861);
or U29309 (N_29309,N_11062,N_16788);
and U29310 (N_29310,N_12186,N_15506);
nand U29311 (N_29311,N_12904,N_11488);
xnor U29312 (N_29312,N_16513,N_13743);
nand U29313 (N_29313,N_15540,N_10978);
xnor U29314 (N_29314,N_15447,N_14314);
and U29315 (N_29315,N_16904,N_16995);
and U29316 (N_29316,N_18331,N_12652);
or U29317 (N_29317,N_17883,N_16154);
nand U29318 (N_29318,N_19212,N_18948);
or U29319 (N_29319,N_19209,N_12118);
nor U29320 (N_29320,N_15176,N_17843);
xnor U29321 (N_29321,N_15854,N_14900);
or U29322 (N_29322,N_18722,N_17204);
and U29323 (N_29323,N_10178,N_13366);
or U29324 (N_29324,N_16947,N_18682);
or U29325 (N_29325,N_14030,N_15514);
nor U29326 (N_29326,N_10625,N_19124);
xnor U29327 (N_29327,N_10417,N_11089);
or U29328 (N_29328,N_15768,N_12102);
nand U29329 (N_29329,N_10915,N_11782);
nor U29330 (N_29330,N_18258,N_18848);
nand U29331 (N_29331,N_18698,N_10280);
xnor U29332 (N_29332,N_12415,N_10834);
xor U29333 (N_29333,N_11788,N_14708);
and U29334 (N_29334,N_14952,N_19531);
or U29335 (N_29335,N_19461,N_12379);
xnor U29336 (N_29336,N_18510,N_19056);
nand U29337 (N_29337,N_16226,N_13731);
nor U29338 (N_29338,N_10370,N_16677);
nand U29339 (N_29339,N_19750,N_10315);
or U29340 (N_29340,N_15504,N_19422);
nor U29341 (N_29341,N_17665,N_19273);
or U29342 (N_29342,N_14196,N_16812);
nor U29343 (N_29343,N_14694,N_15246);
or U29344 (N_29344,N_18413,N_18712);
nor U29345 (N_29345,N_11989,N_13041);
and U29346 (N_29346,N_12347,N_15678);
and U29347 (N_29347,N_13924,N_17679);
nor U29348 (N_29348,N_15719,N_11893);
xnor U29349 (N_29349,N_16582,N_14763);
and U29350 (N_29350,N_14539,N_13314);
nand U29351 (N_29351,N_11478,N_17889);
and U29352 (N_29352,N_19380,N_14722);
and U29353 (N_29353,N_17775,N_16941);
nand U29354 (N_29354,N_17968,N_10463);
nor U29355 (N_29355,N_15936,N_18968);
nand U29356 (N_29356,N_18344,N_13903);
and U29357 (N_29357,N_14112,N_17433);
nor U29358 (N_29358,N_19734,N_12379);
nor U29359 (N_29359,N_11071,N_13513);
nand U29360 (N_29360,N_16767,N_16047);
nand U29361 (N_29361,N_18071,N_13121);
and U29362 (N_29362,N_19982,N_13185);
xor U29363 (N_29363,N_19270,N_19229);
xnor U29364 (N_29364,N_16327,N_12046);
xnor U29365 (N_29365,N_18786,N_19376);
and U29366 (N_29366,N_16600,N_16793);
and U29367 (N_29367,N_11482,N_15004);
xor U29368 (N_29368,N_14686,N_14875);
xor U29369 (N_29369,N_19382,N_18127);
nand U29370 (N_29370,N_19448,N_11588);
or U29371 (N_29371,N_16243,N_12915);
nor U29372 (N_29372,N_17042,N_16951);
or U29373 (N_29373,N_15763,N_12728);
xnor U29374 (N_29374,N_15552,N_10612);
xor U29375 (N_29375,N_10241,N_18331);
and U29376 (N_29376,N_10204,N_14770);
nor U29377 (N_29377,N_18198,N_16277);
nand U29378 (N_29378,N_14650,N_17192);
nand U29379 (N_29379,N_12012,N_19541);
or U29380 (N_29380,N_11091,N_15351);
or U29381 (N_29381,N_15388,N_12144);
or U29382 (N_29382,N_12560,N_13385);
nand U29383 (N_29383,N_14821,N_18331);
and U29384 (N_29384,N_16276,N_13304);
xnor U29385 (N_29385,N_15204,N_17593);
or U29386 (N_29386,N_13680,N_18287);
xor U29387 (N_29387,N_15087,N_10936);
or U29388 (N_29388,N_15416,N_12337);
nor U29389 (N_29389,N_19323,N_19320);
or U29390 (N_29390,N_14766,N_11840);
xnor U29391 (N_29391,N_17122,N_13480);
or U29392 (N_29392,N_15306,N_13654);
and U29393 (N_29393,N_14791,N_15472);
nand U29394 (N_29394,N_10741,N_17146);
nand U29395 (N_29395,N_14909,N_11129);
and U29396 (N_29396,N_10270,N_17850);
nand U29397 (N_29397,N_19069,N_14669);
nor U29398 (N_29398,N_11204,N_15013);
and U29399 (N_29399,N_11348,N_13416);
xnor U29400 (N_29400,N_14536,N_17338);
or U29401 (N_29401,N_10536,N_17727);
and U29402 (N_29402,N_12075,N_19511);
and U29403 (N_29403,N_17224,N_18929);
and U29404 (N_29404,N_13805,N_17459);
nand U29405 (N_29405,N_14025,N_18590);
nor U29406 (N_29406,N_12986,N_13855);
xnor U29407 (N_29407,N_14495,N_15445);
nand U29408 (N_29408,N_13849,N_15292);
xor U29409 (N_29409,N_13815,N_17976);
and U29410 (N_29410,N_16113,N_10774);
and U29411 (N_29411,N_12086,N_16652);
xnor U29412 (N_29412,N_11433,N_11066);
xnor U29413 (N_29413,N_11067,N_12657);
xor U29414 (N_29414,N_13492,N_10266);
nand U29415 (N_29415,N_11878,N_14751);
and U29416 (N_29416,N_10901,N_14250);
nor U29417 (N_29417,N_11648,N_16139);
nand U29418 (N_29418,N_11049,N_16689);
nand U29419 (N_29419,N_17961,N_17323);
xnor U29420 (N_29420,N_16337,N_12886);
nand U29421 (N_29421,N_12367,N_13921);
nand U29422 (N_29422,N_15984,N_11398);
and U29423 (N_29423,N_13352,N_18723);
nor U29424 (N_29424,N_11973,N_14047);
and U29425 (N_29425,N_13904,N_11742);
and U29426 (N_29426,N_11598,N_12957);
and U29427 (N_29427,N_10515,N_12678);
xnor U29428 (N_29428,N_13834,N_19310);
or U29429 (N_29429,N_16316,N_11633);
or U29430 (N_29430,N_10608,N_10783);
and U29431 (N_29431,N_15332,N_11785);
or U29432 (N_29432,N_15333,N_11795);
nor U29433 (N_29433,N_17855,N_18493);
and U29434 (N_29434,N_18620,N_14764);
or U29435 (N_29435,N_16540,N_14312);
or U29436 (N_29436,N_17060,N_18209);
or U29437 (N_29437,N_19480,N_17745);
nor U29438 (N_29438,N_14592,N_14884);
nor U29439 (N_29439,N_18614,N_15256);
xor U29440 (N_29440,N_11872,N_10018);
or U29441 (N_29441,N_12106,N_16276);
nand U29442 (N_29442,N_14624,N_17821);
nor U29443 (N_29443,N_14808,N_17824);
xor U29444 (N_29444,N_12991,N_13906);
or U29445 (N_29445,N_14923,N_17833);
xor U29446 (N_29446,N_13225,N_14936);
or U29447 (N_29447,N_11342,N_14161);
nor U29448 (N_29448,N_11299,N_13296);
and U29449 (N_29449,N_15349,N_12947);
nor U29450 (N_29450,N_18416,N_11686);
nand U29451 (N_29451,N_18680,N_14102);
nor U29452 (N_29452,N_13363,N_15155);
nor U29453 (N_29453,N_14059,N_19786);
nand U29454 (N_29454,N_10708,N_11722);
and U29455 (N_29455,N_14445,N_19575);
nand U29456 (N_29456,N_14368,N_12252);
or U29457 (N_29457,N_10192,N_18199);
or U29458 (N_29458,N_15761,N_14182);
nor U29459 (N_29459,N_18533,N_14623);
xor U29460 (N_29460,N_19734,N_16414);
and U29461 (N_29461,N_17292,N_17719);
or U29462 (N_29462,N_11833,N_13748);
or U29463 (N_29463,N_17719,N_17396);
or U29464 (N_29464,N_16249,N_15746);
nor U29465 (N_29465,N_17436,N_10001);
nand U29466 (N_29466,N_17532,N_14947);
nor U29467 (N_29467,N_11106,N_19323);
or U29468 (N_29468,N_15261,N_19472);
or U29469 (N_29469,N_14498,N_19000);
and U29470 (N_29470,N_11555,N_16643);
nor U29471 (N_29471,N_18793,N_11040);
nand U29472 (N_29472,N_14299,N_18454);
nand U29473 (N_29473,N_13796,N_15982);
xnor U29474 (N_29474,N_17801,N_11661);
or U29475 (N_29475,N_14138,N_17612);
xor U29476 (N_29476,N_19657,N_10217);
xor U29477 (N_29477,N_15909,N_12102);
nor U29478 (N_29478,N_19385,N_16743);
or U29479 (N_29479,N_14200,N_10048);
xor U29480 (N_29480,N_18051,N_14976);
or U29481 (N_29481,N_10174,N_13280);
nor U29482 (N_29482,N_11660,N_13985);
and U29483 (N_29483,N_13922,N_17826);
or U29484 (N_29484,N_13686,N_13146);
and U29485 (N_29485,N_15694,N_19379);
and U29486 (N_29486,N_19484,N_10502);
nand U29487 (N_29487,N_17328,N_19420);
and U29488 (N_29488,N_14236,N_16997);
or U29489 (N_29489,N_13926,N_18674);
or U29490 (N_29490,N_17626,N_19120);
nor U29491 (N_29491,N_13517,N_16314);
xor U29492 (N_29492,N_18554,N_19979);
or U29493 (N_29493,N_19078,N_17007);
nor U29494 (N_29494,N_13495,N_16248);
nor U29495 (N_29495,N_11120,N_10510);
nand U29496 (N_29496,N_17002,N_14488);
xor U29497 (N_29497,N_14322,N_12025);
nor U29498 (N_29498,N_10756,N_19689);
and U29499 (N_29499,N_11831,N_17219);
or U29500 (N_29500,N_13417,N_18746);
and U29501 (N_29501,N_19576,N_15779);
or U29502 (N_29502,N_16526,N_14121);
and U29503 (N_29503,N_19203,N_19987);
nor U29504 (N_29504,N_13562,N_14937);
nand U29505 (N_29505,N_10956,N_13589);
nand U29506 (N_29506,N_16310,N_15754);
nor U29507 (N_29507,N_16855,N_10086);
nand U29508 (N_29508,N_11942,N_11278);
or U29509 (N_29509,N_13794,N_10786);
nand U29510 (N_29510,N_16870,N_12650);
and U29511 (N_29511,N_17447,N_10086);
xnor U29512 (N_29512,N_11249,N_17283);
and U29513 (N_29513,N_17403,N_12040);
xor U29514 (N_29514,N_10283,N_11423);
xnor U29515 (N_29515,N_17488,N_13758);
and U29516 (N_29516,N_14969,N_13573);
and U29517 (N_29517,N_12905,N_10374);
and U29518 (N_29518,N_14280,N_15491);
nand U29519 (N_29519,N_10205,N_12873);
and U29520 (N_29520,N_18022,N_13167);
nand U29521 (N_29521,N_11209,N_12930);
xor U29522 (N_29522,N_18029,N_10349);
and U29523 (N_29523,N_11736,N_13425);
xor U29524 (N_29524,N_11384,N_10872);
nand U29525 (N_29525,N_15503,N_18060);
nand U29526 (N_29526,N_17866,N_17461);
xnor U29527 (N_29527,N_14043,N_18497);
and U29528 (N_29528,N_19523,N_14122);
or U29529 (N_29529,N_15531,N_17677);
or U29530 (N_29530,N_15333,N_17959);
xnor U29531 (N_29531,N_11443,N_17350);
or U29532 (N_29532,N_13318,N_10120);
or U29533 (N_29533,N_19456,N_17332);
and U29534 (N_29534,N_18063,N_10480);
xor U29535 (N_29535,N_19588,N_11438);
or U29536 (N_29536,N_13081,N_10964);
nand U29537 (N_29537,N_16544,N_16744);
nand U29538 (N_29538,N_12784,N_11200);
nand U29539 (N_29539,N_17931,N_17660);
nor U29540 (N_29540,N_17117,N_12035);
or U29541 (N_29541,N_16455,N_10470);
xnor U29542 (N_29542,N_18344,N_19055);
or U29543 (N_29543,N_19882,N_12272);
xor U29544 (N_29544,N_16008,N_15447);
xnor U29545 (N_29545,N_17089,N_17837);
or U29546 (N_29546,N_18349,N_13622);
nand U29547 (N_29547,N_13604,N_11657);
nand U29548 (N_29548,N_12469,N_10767);
xnor U29549 (N_29549,N_15908,N_16260);
xor U29550 (N_29550,N_17277,N_17615);
nand U29551 (N_29551,N_11821,N_17467);
nor U29552 (N_29552,N_16729,N_10760);
and U29553 (N_29553,N_10474,N_17878);
nand U29554 (N_29554,N_18641,N_11516);
nor U29555 (N_29555,N_12108,N_15667);
nand U29556 (N_29556,N_14636,N_19496);
nand U29557 (N_29557,N_15127,N_19218);
xor U29558 (N_29558,N_17377,N_16981);
or U29559 (N_29559,N_16149,N_14327);
nor U29560 (N_29560,N_16162,N_17133);
or U29561 (N_29561,N_14247,N_19468);
xnor U29562 (N_29562,N_12089,N_11055);
or U29563 (N_29563,N_14917,N_12361);
xor U29564 (N_29564,N_18285,N_17618);
nand U29565 (N_29565,N_18990,N_15913);
and U29566 (N_29566,N_18706,N_15347);
nand U29567 (N_29567,N_12552,N_15707);
and U29568 (N_29568,N_13626,N_14654);
and U29569 (N_29569,N_15397,N_13866);
nor U29570 (N_29570,N_11216,N_10422);
nor U29571 (N_29571,N_11283,N_13905);
nor U29572 (N_29572,N_11200,N_13596);
nor U29573 (N_29573,N_15775,N_19953);
and U29574 (N_29574,N_17401,N_18340);
and U29575 (N_29575,N_16464,N_16777);
or U29576 (N_29576,N_17178,N_10494);
xor U29577 (N_29577,N_18314,N_13011);
and U29578 (N_29578,N_12220,N_13414);
nand U29579 (N_29579,N_19894,N_15979);
or U29580 (N_29580,N_11187,N_19144);
and U29581 (N_29581,N_18086,N_13129);
or U29582 (N_29582,N_13945,N_10175);
nand U29583 (N_29583,N_16057,N_19314);
and U29584 (N_29584,N_16760,N_18285);
xor U29585 (N_29585,N_16405,N_13791);
and U29586 (N_29586,N_13784,N_10541);
nand U29587 (N_29587,N_16734,N_12364);
xnor U29588 (N_29588,N_16038,N_18018);
xor U29589 (N_29589,N_16442,N_18520);
xnor U29590 (N_29590,N_15424,N_14858);
and U29591 (N_29591,N_13939,N_11516);
xnor U29592 (N_29592,N_12927,N_14096);
nor U29593 (N_29593,N_18188,N_13383);
or U29594 (N_29594,N_18315,N_11431);
nor U29595 (N_29595,N_11482,N_11882);
nor U29596 (N_29596,N_18073,N_17335);
xor U29597 (N_29597,N_13584,N_15355);
and U29598 (N_29598,N_16024,N_16847);
or U29599 (N_29599,N_13308,N_17464);
or U29600 (N_29600,N_12473,N_15918);
or U29601 (N_29601,N_14616,N_19996);
nand U29602 (N_29602,N_18111,N_12536);
nor U29603 (N_29603,N_14235,N_13015);
and U29604 (N_29604,N_14564,N_16708);
or U29605 (N_29605,N_19927,N_13611);
nand U29606 (N_29606,N_14131,N_14943);
and U29607 (N_29607,N_11788,N_10593);
xor U29608 (N_29608,N_16910,N_13472);
nor U29609 (N_29609,N_12334,N_11302);
or U29610 (N_29610,N_16000,N_14752);
nor U29611 (N_29611,N_13119,N_17253);
nor U29612 (N_29612,N_12125,N_19861);
nand U29613 (N_29613,N_16176,N_10210);
or U29614 (N_29614,N_13251,N_11528);
nand U29615 (N_29615,N_17843,N_10647);
nand U29616 (N_29616,N_18862,N_11518);
xnor U29617 (N_29617,N_15495,N_14634);
and U29618 (N_29618,N_15696,N_18319);
nor U29619 (N_29619,N_19583,N_10849);
nor U29620 (N_29620,N_10670,N_18651);
nand U29621 (N_29621,N_10599,N_16633);
and U29622 (N_29622,N_19117,N_13317);
and U29623 (N_29623,N_11671,N_17997);
nand U29624 (N_29624,N_10857,N_16159);
xnor U29625 (N_29625,N_17068,N_12831);
nor U29626 (N_29626,N_14991,N_13036);
xor U29627 (N_29627,N_12318,N_19832);
and U29628 (N_29628,N_16180,N_13238);
nand U29629 (N_29629,N_13515,N_13166);
nor U29630 (N_29630,N_19713,N_12532);
or U29631 (N_29631,N_17533,N_19241);
or U29632 (N_29632,N_19110,N_17231);
xor U29633 (N_29633,N_14553,N_17029);
and U29634 (N_29634,N_11643,N_15715);
nor U29635 (N_29635,N_13246,N_14066);
xnor U29636 (N_29636,N_14668,N_19225);
nand U29637 (N_29637,N_12000,N_11678);
or U29638 (N_29638,N_15250,N_13600);
or U29639 (N_29639,N_18651,N_16484);
and U29640 (N_29640,N_13504,N_19118);
nand U29641 (N_29641,N_10739,N_12445);
xnor U29642 (N_29642,N_10418,N_11249);
nand U29643 (N_29643,N_13174,N_19207);
or U29644 (N_29644,N_10952,N_16161);
and U29645 (N_29645,N_14335,N_18723);
nor U29646 (N_29646,N_12599,N_15196);
or U29647 (N_29647,N_19732,N_17810);
and U29648 (N_29648,N_18053,N_13023);
nand U29649 (N_29649,N_12477,N_15889);
and U29650 (N_29650,N_11443,N_11212);
or U29651 (N_29651,N_12862,N_17686);
nor U29652 (N_29652,N_16955,N_17427);
xnor U29653 (N_29653,N_11194,N_13581);
nor U29654 (N_29654,N_18499,N_14001);
or U29655 (N_29655,N_10292,N_11793);
xor U29656 (N_29656,N_16469,N_11579);
and U29657 (N_29657,N_17305,N_17683);
nand U29658 (N_29658,N_16765,N_17337);
nand U29659 (N_29659,N_16307,N_12747);
xnor U29660 (N_29660,N_14904,N_12609);
nand U29661 (N_29661,N_11107,N_18496);
nand U29662 (N_29662,N_12135,N_10207);
and U29663 (N_29663,N_14425,N_13403);
and U29664 (N_29664,N_12376,N_13265);
nor U29665 (N_29665,N_15511,N_12232);
and U29666 (N_29666,N_17477,N_17587);
nor U29667 (N_29667,N_17898,N_13351);
nand U29668 (N_29668,N_15435,N_18103);
or U29669 (N_29669,N_14808,N_14484);
and U29670 (N_29670,N_11750,N_18695);
or U29671 (N_29671,N_15191,N_16474);
nand U29672 (N_29672,N_18871,N_15834);
or U29673 (N_29673,N_10547,N_12540);
xor U29674 (N_29674,N_17659,N_13087);
nand U29675 (N_29675,N_10324,N_17429);
nor U29676 (N_29676,N_12657,N_16096);
nor U29677 (N_29677,N_16511,N_11471);
and U29678 (N_29678,N_11288,N_12941);
or U29679 (N_29679,N_14922,N_14428);
xnor U29680 (N_29680,N_10083,N_19251);
nand U29681 (N_29681,N_18028,N_19184);
nand U29682 (N_29682,N_10702,N_19834);
and U29683 (N_29683,N_15019,N_16111);
nand U29684 (N_29684,N_10161,N_11091);
or U29685 (N_29685,N_19268,N_14256);
nand U29686 (N_29686,N_18771,N_10436);
xnor U29687 (N_29687,N_18368,N_12380);
nor U29688 (N_29688,N_14685,N_14686);
nor U29689 (N_29689,N_15154,N_13295);
and U29690 (N_29690,N_11164,N_11815);
or U29691 (N_29691,N_13692,N_13800);
and U29692 (N_29692,N_13344,N_10105);
and U29693 (N_29693,N_11883,N_18468);
or U29694 (N_29694,N_15850,N_16372);
nor U29695 (N_29695,N_16405,N_19711);
and U29696 (N_29696,N_14052,N_15623);
or U29697 (N_29697,N_16891,N_17599);
or U29698 (N_29698,N_18112,N_10136);
or U29699 (N_29699,N_13992,N_10752);
and U29700 (N_29700,N_19746,N_15590);
or U29701 (N_29701,N_16964,N_17984);
xnor U29702 (N_29702,N_17023,N_14195);
xnor U29703 (N_29703,N_10900,N_13765);
nor U29704 (N_29704,N_14111,N_10928);
xor U29705 (N_29705,N_16193,N_18755);
nand U29706 (N_29706,N_10571,N_10738);
nand U29707 (N_29707,N_10824,N_11935);
xor U29708 (N_29708,N_13543,N_14750);
nor U29709 (N_29709,N_15057,N_16832);
and U29710 (N_29710,N_18973,N_16850);
and U29711 (N_29711,N_10660,N_16222);
or U29712 (N_29712,N_19473,N_13085);
nor U29713 (N_29713,N_18533,N_16345);
or U29714 (N_29714,N_18206,N_10650);
nand U29715 (N_29715,N_19020,N_18105);
or U29716 (N_29716,N_12556,N_15953);
nand U29717 (N_29717,N_19310,N_14244);
nor U29718 (N_29718,N_17767,N_14478);
nor U29719 (N_29719,N_15796,N_13916);
or U29720 (N_29720,N_16637,N_11435);
or U29721 (N_29721,N_16167,N_11009);
xnor U29722 (N_29722,N_18532,N_18124);
nor U29723 (N_29723,N_18733,N_12558);
nand U29724 (N_29724,N_19372,N_14677);
nand U29725 (N_29725,N_13907,N_16839);
or U29726 (N_29726,N_11466,N_15277);
nand U29727 (N_29727,N_15663,N_19559);
xor U29728 (N_29728,N_18813,N_11726);
and U29729 (N_29729,N_16740,N_19356);
nand U29730 (N_29730,N_19076,N_16958);
nand U29731 (N_29731,N_10311,N_16315);
xor U29732 (N_29732,N_10760,N_14236);
nand U29733 (N_29733,N_16047,N_19658);
and U29734 (N_29734,N_18672,N_11416);
or U29735 (N_29735,N_12809,N_12711);
nand U29736 (N_29736,N_13067,N_11219);
and U29737 (N_29737,N_10209,N_12574);
nand U29738 (N_29738,N_19680,N_14060);
and U29739 (N_29739,N_19198,N_11570);
and U29740 (N_29740,N_16182,N_17263);
nand U29741 (N_29741,N_15633,N_16397);
and U29742 (N_29742,N_14281,N_10547);
or U29743 (N_29743,N_17406,N_15692);
xor U29744 (N_29744,N_11650,N_18400);
and U29745 (N_29745,N_10768,N_12741);
nand U29746 (N_29746,N_13308,N_19576);
xnor U29747 (N_29747,N_14114,N_15081);
and U29748 (N_29748,N_13469,N_11674);
nand U29749 (N_29749,N_14179,N_18014);
nand U29750 (N_29750,N_16141,N_14245);
or U29751 (N_29751,N_12875,N_11618);
nor U29752 (N_29752,N_19752,N_17217);
xnor U29753 (N_29753,N_14925,N_11927);
or U29754 (N_29754,N_18440,N_15596);
and U29755 (N_29755,N_10588,N_17018);
nor U29756 (N_29756,N_14372,N_18032);
and U29757 (N_29757,N_10041,N_11340);
nand U29758 (N_29758,N_19182,N_15013);
and U29759 (N_29759,N_14417,N_12418);
nand U29760 (N_29760,N_16799,N_17582);
nor U29761 (N_29761,N_12035,N_13742);
or U29762 (N_29762,N_16545,N_11626);
nand U29763 (N_29763,N_11578,N_17979);
or U29764 (N_29764,N_17379,N_13125);
or U29765 (N_29765,N_17413,N_15278);
xnor U29766 (N_29766,N_19049,N_10238);
xor U29767 (N_29767,N_16331,N_13786);
and U29768 (N_29768,N_15093,N_19951);
nand U29769 (N_29769,N_11957,N_18433);
and U29770 (N_29770,N_17570,N_12456);
and U29771 (N_29771,N_18410,N_10819);
and U29772 (N_29772,N_10538,N_13878);
and U29773 (N_29773,N_12398,N_13108);
or U29774 (N_29774,N_12918,N_16418);
and U29775 (N_29775,N_13971,N_11250);
or U29776 (N_29776,N_16358,N_14549);
or U29777 (N_29777,N_12431,N_18878);
nand U29778 (N_29778,N_19541,N_18689);
and U29779 (N_29779,N_10826,N_10208);
nand U29780 (N_29780,N_18499,N_10416);
nor U29781 (N_29781,N_17424,N_13403);
and U29782 (N_29782,N_10622,N_17222);
xnor U29783 (N_29783,N_17724,N_11267);
nor U29784 (N_29784,N_16339,N_10439);
and U29785 (N_29785,N_13799,N_15202);
xor U29786 (N_29786,N_15655,N_12483);
nor U29787 (N_29787,N_11604,N_12754);
and U29788 (N_29788,N_14131,N_19416);
xnor U29789 (N_29789,N_19792,N_16424);
nand U29790 (N_29790,N_16050,N_10073);
xnor U29791 (N_29791,N_10840,N_10549);
and U29792 (N_29792,N_15560,N_15072);
nand U29793 (N_29793,N_18646,N_12727);
or U29794 (N_29794,N_12776,N_19765);
xnor U29795 (N_29795,N_14455,N_19748);
or U29796 (N_29796,N_19588,N_16584);
nand U29797 (N_29797,N_13063,N_19307);
and U29798 (N_29798,N_16342,N_19197);
and U29799 (N_29799,N_17295,N_13605);
nor U29800 (N_29800,N_19911,N_13374);
nand U29801 (N_29801,N_18882,N_11965);
nor U29802 (N_29802,N_14443,N_16183);
xor U29803 (N_29803,N_14459,N_11580);
and U29804 (N_29804,N_17640,N_12144);
or U29805 (N_29805,N_18415,N_12681);
and U29806 (N_29806,N_14666,N_13544);
and U29807 (N_29807,N_14830,N_17563);
nand U29808 (N_29808,N_17403,N_19729);
nor U29809 (N_29809,N_15883,N_15591);
nor U29810 (N_29810,N_19637,N_18338);
and U29811 (N_29811,N_12316,N_19607);
and U29812 (N_29812,N_19064,N_15757);
xnor U29813 (N_29813,N_19555,N_11328);
nor U29814 (N_29814,N_10008,N_11226);
or U29815 (N_29815,N_16431,N_19246);
xor U29816 (N_29816,N_13666,N_19280);
and U29817 (N_29817,N_19311,N_17255);
or U29818 (N_29818,N_14182,N_16009);
xor U29819 (N_29819,N_14474,N_18765);
nand U29820 (N_29820,N_16414,N_15083);
nand U29821 (N_29821,N_14206,N_13187);
and U29822 (N_29822,N_10446,N_12337);
and U29823 (N_29823,N_19504,N_18276);
nor U29824 (N_29824,N_13696,N_19056);
and U29825 (N_29825,N_16519,N_17279);
nor U29826 (N_29826,N_16772,N_10986);
nor U29827 (N_29827,N_11732,N_17119);
and U29828 (N_29828,N_17410,N_18505);
or U29829 (N_29829,N_19797,N_18183);
xnor U29830 (N_29830,N_17566,N_10068);
or U29831 (N_29831,N_19564,N_17635);
or U29832 (N_29832,N_11377,N_15709);
xnor U29833 (N_29833,N_19872,N_10731);
and U29834 (N_29834,N_19458,N_15334);
nor U29835 (N_29835,N_16880,N_12825);
xor U29836 (N_29836,N_16775,N_18253);
or U29837 (N_29837,N_10567,N_18914);
and U29838 (N_29838,N_18092,N_13383);
xnor U29839 (N_29839,N_13000,N_15189);
and U29840 (N_29840,N_18563,N_16991);
or U29841 (N_29841,N_17945,N_13933);
xor U29842 (N_29842,N_18025,N_10550);
or U29843 (N_29843,N_19860,N_19487);
nor U29844 (N_29844,N_16988,N_15918);
xnor U29845 (N_29845,N_16511,N_14097);
nor U29846 (N_29846,N_14935,N_10430);
and U29847 (N_29847,N_17581,N_10014);
nand U29848 (N_29848,N_18765,N_13903);
or U29849 (N_29849,N_12640,N_15175);
and U29850 (N_29850,N_14211,N_13444);
and U29851 (N_29851,N_10990,N_10918);
and U29852 (N_29852,N_14949,N_15769);
nor U29853 (N_29853,N_10309,N_14467);
nand U29854 (N_29854,N_18366,N_18873);
nand U29855 (N_29855,N_10159,N_13164);
xnor U29856 (N_29856,N_19027,N_18826);
nand U29857 (N_29857,N_15818,N_16958);
xnor U29858 (N_29858,N_11986,N_14364);
nand U29859 (N_29859,N_13442,N_16829);
xnor U29860 (N_29860,N_16796,N_12120);
nor U29861 (N_29861,N_15624,N_17359);
and U29862 (N_29862,N_14690,N_16371);
nor U29863 (N_29863,N_11145,N_10410);
and U29864 (N_29864,N_18254,N_10399);
xor U29865 (N_29865,N_18924,N_12394);
xnor U29866 (N_29866,N_16077,N_17886);
xnor U29867 (N_29867,N_17223,N_17248);
nand U29868 (N_29868,N_17682,N_10625);
nand U29869 (N_29869,N_10671,N_18395);
nor U29870 (N_29870,N_14211,N_19853);
or U29871 (N_29871,N_17859,N_15144);
nor U29872 (N_29872,N_12677,N_10298);
or U29873 (N_29873,N_11179,N_13619);
nor U29874 (N_29874,N_19642,N_18574);
nand U29875 (N_29875,N_13257,N_16364);
nand U29876 (N_29876,N_19907,N_16816);
nand U29877 (N_29877,N_19564,N_11630);
and U29878 (N_29878,N_12179,N_11841);
and U29879 (N_29879,N_19318,N_12367);
and U29880 (N_29880,N_15260,N_11157);
or U29881 (N_29881,N_16354,N_10206);
and U29882 (N_29882,N_16686,N_16238);
or U29883 (N_29883,N_18217,N_12439);
xor U29884 (N_29884,N_10633,N_13530);
and U29885 (N_29885,N_10015,N_14600);
or U29886 (N_29886,N_12400,N_11644);
nand U29887 (N_29887,N_15987,N_18254);
nor U29888 (N_29888,N_18119,N_11544);
or U29889 (N_29889,N_12012,N_18464);
nand U29890 (N_29890,N_18928,N_15747);
nor U29891 (N_29891,N_13877,N_14270);
and U29892 (N_29892,N_15967,N_14925);
nand U29893 (N_29893,N_19451,N_17782);
nand U29894 (N_29894,N_15969,N_13148);
and U29895 (N_29895,N_13846,N_18219);
xnor U29896 (N_29896,N_13511,N_19322);
and U29897 (N_29897,N_10468,N_14426);
nor U29898 (N_29898,N_14924,N_17557);
or U29899 (N_29899,N_13495,N_18189);
xnor U29900 (N_29900,N_11590,N_10813);
nand U29901 (N_29901,N_12868,N_14607);
nor U29902 (N_29902,N_13374,N_19552);
xnor U29903 (N_29903,N_11504,N_10168);
xor U29904 (N_29904,N_18832,N_11067);
nand U29905 (N_29905,N_12241,N_17992);
nand U29906 (N_29906,N_18276,N_13782);
nor U29907 (N_29907,N_10045,N_11001);
xnor U29908 (N_29908,N_15873,N_13900);
nor U29909 (N_29909,N_19036,N_10217);
nor U29910 (N_29910,N_10880,N_13589);
nor U29911 (N_29911,N_10934,N_13012);
xnor U29912 (N_29912,N_11171,N_11476);
or U29913 (N_29913,N_13606,N_17298);
or U29914 (N_29914,N_19047,N_18193);
xnor U29915 (N_29915,N_10072,N_11556);
xor U29916 (N_29916,N_16539,N_17187);
or U29917 (N_29917,N_12789,N_14659);
nor U29918 (N_29918,N_15017,N_14522);
nand U29919 (N_29919,N_10718,N_15881);
nor U29920 (N_29920,N_17198,N_15414);
xnor U29921 (N_29921,N_13060,N_19521);
or U29922 (N_29922,N_10174,N_11542);
nand U29923 (N_29923,N_10909,N_14665);
nand U29924 (N_29924,N_18389,N_15523);
nand U29925 (N_29925,N_15352,N_14008);
xnor U29926 (N_29926,N_11655,N_12478);
nand U29927 (N_29927,N_12765,N_10409);
nand U29928 (N_29928,N_10298,N_19930);
nor U29929 (N_29929,N_14407,N_17646);
nand U29930 (N_29930,N_19809,N_13847);
and U29931 (N_29931,N_12798,N_15521);
nor U29932 (N_29932,N_10541,N_18489);
nor U29933 (N_29933,N_14883,N_11427);
nand U29934 (N_29934,N_19228,N_10213);
nand U29935 (N_29935,N_10323,N_15336);
or U29936 (N_29936,N_10624,N_15182);
and U29937 (N_29937,N_12384,N_13756);
nand U29938 (N_29938,N_14628,N_19332);
xor U29939 (N_29939,N_17733,N_15664);
xor U29940 (N_29940,N_17482,N_18704);
and U29941 (N_29941,N_11044,N_14708);
nor U29942 (N_29942,N_18835,N_13049);
and U29943 (N_29943,N_15017,N_11383);
or U29944 (N_29944,N_11041,N_13558);
nand U29945 (N_29945,N_12328,N_17300);
nand U29946 (N_29946,N_11945,N_18203);
or U29947 (N_29947,N_19577,N_12553);
nand U29948 (N_29948,N_12965,N_19496);
xnor U29949 (N_29949,N_11676,N_17086);
or U29950 (N_29950,N_12314,N_15798);
xor U29951 (N_29951,N_11495,N_18251);
xnor U29952 (N_29952,N_11471,N_18666);
or U29953 (N_29953,N_19629,N_12584);
or U29954 (N_29954,N_11463,N_17432);
nand U29955 (N_29955,N_19759,N_11824);
nand U29956 (N_29956,N_10788,N_11282);
xor U29957 (N_29957,N_10625,N_11145);
nand U29958 (N_29958,N_11495,N_14167);
nand U29959 (N_29959,N_14971,N_12546);
xnor U29960 (N_29960,N_19878,N_14309);
xor U29961 (N_29961,N_14264,N_19063);
and U29962 (N_29962,N_12944,N_17378);
or U29963 (N_29963,N_13318,N_19530);
nor U29964 (N_29964,N_19788,N_11377);
nor U29965 (N_29965,N_16509,N_15245);
nor U29966 (N_29966,N_10473,N_15510);
and U29967 (N_29967,N_18985,N_12446);
and U29968 (N_29968,N_11942,N_15117);
nor U29969 (N_29969,N_14650,N_10171);
or U29970 (N_29970,N_12085,N_11442);
and U29971 (N_29971,N_10575,N_16855);
and U29972 (N_29972,N_10254,N_11827);
nor U29973 (N_29973,N_10108,N_16503);
nor U29974 (N_29974,N_19295,N_17807);
and U29975 (N_29975,N_13624,N_16454);
xor U29976 (N_29976,N_16882,N_15541);
xor U29977 (N_29977,N_14198,N_16373);
and U29978 (N_29978,N_15583,N_19889);
and U29979 (N_29979,N_12063,N_16180);
nand U29980 (N_29980,N_13122,N_18484);
nand U29981 (N_29981,N_19710,N_17732);
xnor U29982 (N_29982,N_18331,N_13207);
nor U29983 (N_29983,N_15578,N_16518);
and U29984 (N_29984,N_12230,N_14900);
nor U29985 (N_29985,N_19467,N_15349);
nand U29986 (N_29986,N_13214,N_13322);
nor U29987 (N_29987,N_13527,N_12039);
and U29988 (N_29988,N_10385,N_15306);
nor U29989 (N_29989,N_11855,N_19695);
xnor U29990 (N_29990,N_11049,N_18917);
nand U29991 (N_29991,N_12023,N_14634);
and U29992 (N_29992,N_17338,N_15848);
or U29993 (N_29993,N_11236,N_13365);
or U29994 (N_29994,N_14911,N_19453);
and U29995 (N_29995,N_14517,N_13270);
or U29996 (N_29996,N_14711,N_18429);
xor U29997 (N_29997,N_17916,N_15694);
and U29998 (N_29998,N_11265,N_14246);
xor U29999 (N_29999,N_14142,N_13619);
and U30000 (N_30000,N_25507,N_27843);
and U30001 (N_30001,N_22770,N_24875);
and U30002 (N_30002,N_22759,N_26222);
or U30003 (N_30003,N_24000,N_20485);
nor U30004 (N_30004,N_29782,N_27616);
or U30005 (N_30005,N_23938,N_24506);
nand U30006 (N_30006,N_28309,N_28030);
or U30007 (N_30007,N_27367,N_22542);
nand U30008 (N_30008,N_26914,N_29692);
and U30009 (N_30009,N_20161,N_27278);
and U30010 (N_30010,N_23445,N_23302);
or U30011 (N_30011,N_28067,N_23928);
xor U30012 (N_30012,N_27076,N_26989);
nor U30013 (N_30013,N_21586,N_22794);
nand U30014 (N_30014,N_23325,N_22048);
nor U30015 (N_30015,N_26050,N_27964);
or U30016 (N_30016,N_22516,N_29390);
or U30017 (N_30017,N_23007,N_24704);
or U30018 (N_30018,N_25500,N_29015);
and U30019 (N_30019,N_28549,N_21344);
or U30020 (N_30020,N_20770,N_24102);
and U30021 (N_30021,N_27928,N_24291);
xnor U30022 (N_30022,N_25276,N_22891);
nand U30023 (N_30023,N_21773,N_26065);
nor U30024 (N_30024,N_29245,N_26161);
nand U30025 (N_30025,N_28459,N_22472);
nor U30026 (N_30026,N_23461,N_29543);
nand U30027 (N_30027,N_29274,N_26345);
or U30028 (N_30028,N_22817,N_24959);
xor U30029 (N_30029,N_20557,N_23969);
nor U30030 (N_30030,N_26575,N_29779);
xnor U30031 (N_30031,N_24748,N_23207);
or U30032 (N_30032,N_25737,N_20228);
nand U30033 (N_30033,N_20958,N_20178);
or U30034 (N_30034,N_20482,N_20848);
nand U30035 (N_30035,N_27041,N_21516);
xor U30036 (N_30036,N_22800,N_23821);
nand U30037 (N_30037,N_24861,N_22624);
and U30038 (N_30038,N_20144,N_20158);
nand U30039 (N_30039,N_24872,N_26362);
xnor U30040 (N_30040,N_25562,N_26460);
nand U30041 (N_30041,N_27286,N_28970);
xor U30042 (N_30042,N_22562,N_22417);
xnor U30043 (N_30043,N_28454,N_26687);
xor U30044 (N_30044,N_24715,N_26878);
nor U30045 (N_30045,N_29127,N_29568);
or U30046 (N_30046,N_20563,N_25846);
xor U30047 (N_30047,N_21665,N_29485);
nor U30048 (N_30048,N_24422,N_27776);
nand U30049 (N_30049,N_20494,N_26517);
nor U30050 (N_30050,N_27812,N_20465);
or U30051 (N_30051,N_20369,N_26885);
or U30052 (N_30052,N_29511,N_28987);
xnor U30053 (N_30053,N_21270,N_24595);
nand U30054 (N_30054,N_29350,N_26537);
and U30055 (N_30055,N_22169,N_26074);
nor U30056 (N_30056,N_27628,N_23499);
nand U30057 (N_30057,N_26711,N_21560);
nand U30058 (N_30058,N_29554,N_25682);
nor U30059 (N_30059,N_27137,N_25528);
nand U30060 (N_30060,N_23882,N_25952);
and U30061 (N_30061,N_27969,N_29675);
nand U30062 (N_30062,N_21712,N_29225);
and U30063 (N_30063,N_25373,N_28321);
nor U30064 (N_30064,N_27291,N_29179);
nand U30065 (N_30065,N_26151,N_23567);
and U30066 (N_30066,N_20608,N_20022);
xor U30067 (N_30067,N_24464,N_21785);
nor U30068 (N_30068,N_21535,N_23684);
and U30069 (N_30069,N_25961,N_27045);
nand U30070 (N_30070,N_21320,N_25463);
xor U30071 (N_30071,N_25999,N_24455);
nor U30072 (N_30072,N_23787,N_23392);
or U30073 (N_30073,N_25142,N_20857);
nor U30074 (N_30074,N_20719,N_22005);
nor U30075 (N_30075,N_29973,N_29519);
xnor U30076 (N_30076,N_28134,N_28529);
or U30077 (N_30077,N_23604,N_26128);
nand U30078 (N_30078,N_21779,N_23805);
nor U30079 (N_30079,N_23597,N_23330);
xnor U30080 (N_30080,N_22211,N_23878);
or U30081 (N_30081,N_29959,N_29659);
nand U30082 (N_30082,N_24233,N_26674);
xor U30083 (N_30083,N_28364,N_26634);
nor U30084 (N_30084,N_25460,N_21225);
or U30085 (N_30085,N_29770,N_28770);
and U30086 (N_30086,N_24254,N_23415);
xnor U30087 (N_30087,N_23926,N_20860);
xor U30088 (N_30088,N_22635,N_22029);
or U30089 (N_30089,N_22411,N_22805);
or U30090 (N_30090,N_29385,N_25055);
xor U30091 (N_30091,N_21108,N_28943);
nor U30092 (N_30092,N_20548,N_29792);
nand U30093 (N_30093,N_25187,N_24386);
or U30094 (N_30094,N_22359,N_24321);
nor U30095 (N_30095,N_25036,N_28090);
xor U30096 (N_30096,N_28887,N_23923);
and U30097 (N_30097,N_24678,N_23861);
nor U30098 (N_30098,N_28316,N_20835);
xnor U30099 (N_30099,N_27968,N_29491);
nand U30100 (N_30100,N_20297,N_28594);
nor U30101 (N_30101,N_22612,N_23212);
and U30102 (N_30102,N_28659,N_27111);
and U30103 (N_30103,N_29832,N_26646);
xnor U30104 (N_30104,N_22843,N_20493);
and U30105 (N_30105,N_21121,N_23864);
or U30106 (N_30106,N_28170,N_28033);
or U30107 (N_30107,N_20527,N_26941);
and U30108 (N_30108,N_28655,N_22526);
nor U30109 (N_30109,N_25315,N_21130);
nand U30110 (N_30110,N_22969,N_25414);
and U30111 (N_30111,N_24919,N_23956);
nor U30112 (N_30112,N_26335,N_26834);
and U30113 (N_30113,N_22815,N_23135);
nand U30114 (N_30114,N_25242,N_25447);
and U30115 (N_30115,N_27477,N_28968);
xor U30116 (N_30116,N_22754,N_20047);
nand U30117 (N_30117,N_25720,N_24206);
and U30118 (N_30118,N_28455,N_29334);
nand U30119 (N_30119,N_28308,N_26666);
or U30120 (N_30120,N_22210,N_22545);
xor U30121 (N_30121,N_22024,N_25780);
nor U30122 (N_30122,N_27324,N_26645);
and U30123 (N_30123,N_29540,N_25683);
xnor U30124 (N_30124,N_20345,N_23924);
or U30125 (N_30125,N_25743,N_23335);
or U30126 (N_30126,N_28388,N_27813);
nor U30127 (N_30127,N_21182,N_28115);
or U30128 (N_30128,N_25084,N_26073);
or U30129 (N_30129,N_29261,N_24469);
xnor U30130 (N_30130,N_26112,N_25611);
nand U30131 (N_30131,N_25863,N_25858);
xnor U30132 (N_30132,N_25081,N_21633);
nand U30133 (N_30133,N_22599,N_28962);
and U30134 (N_30134,N_23568,N_29430);
or U30135 (N_30135,N_22954,N_27900);
or U30136 (N_30136,N_27890,N_22106);
nor U30137 (N_30137,N_25432,N_26173);
nand U30138 (N_30138,N_20112,N_27453);
nand U30139 (N_30139,N_29913,N_20124);
or U30140 (N_30140,N_24801,N_21596);
nor U30141 (N_30141,N_24251,N_22603);
or U30142 (N_30142,N_27793,N_21036);
or U30143 (N_30143,N_28573,N_20535);
nor U30144 (N_30144,N_29871,N_25016);
or U30145 (N_30145,N_27904,N_20694);
xor U30146 (N_30146,N_29570,N_29704);
and U30147 (N_30147,N_21867,N_20425);
xnor U30148 (N_30148,N_22042,N_27195);
nand U30149 (N_30149,N_22026,N_20564);
and U30150 (N_30150,N_28158,N_26054);
and U30151 (N_30151,N_28286,N_26794);
and U30152 (N_30152,N_25206,N_22136);
nand U30153 (N_30153,N_29373,N_28534);
nor U30154 (N_30154,N_25174,N_20496);
nand U30155 (N_30155,N_29918,N_24557);
nand U30156 (N_30156,N_28692,N_26308);
or U30157 (N_30157,N_22822,N_28038);
nand U30158 (N_30158,N_20332,N_24732);
nor U30159 (N_30159,N_23714,N_29229);
and U30160 (N_30160,N_26313,N_25211);
and U30161 (N_30161,N_23594,N_24038);
nand U30162 (N_30162,N_26531,N_28965);
and U30163 (N_30163,N_27850,N_21025);
nor U30164 (N_30164,N_22880,N_28404);
or U30165 (N_30165,N_22144,N_29369);
nor U30166 (N_30166,N_21663,N_25191);
xor U30167 (N_30167,N_23671,N_26767);
nand U30168 (N_30168,N_27482,N_23528);
nand U30169 (N_30169,N_23009,N_28992);
xor U30170 (N_30170,N_24138,N_20976);
nor U30171 (N_30171,N_27436,N_22115);
nor U30172 (N_30172,N_26657,N_22747);
xor U30173 (N_30173,N_23770,N_20367);
and U30174 (N_30174,N_26723,N_26579);
xnor U30175 (N_30175,N_22512,N_24515);
or U30176 (N_30176,N_22320,N_25976);
xor U30177 (N_30177,N_26326,N_29510);
nand U30178 (N_30178,N_24825,N_22586);
xnor U30179 (N_30179,N_21731,N_22648);
or U30180 (N_30180,N_22540,N_28941);
xnor U30181 (N_30181,N_22498,N_24454);
or U30182 (N_30182,N_23658,N_28403);
or U30183 (N_30183,N_29977,N_20680);
or U30184 (N_30184,N_26338,N_20206);
and U30185 (N_30185,N_28359,N_28409);
or U30186 (N_30186,N_23583,N_25089);
nor U30187 (N_30187,N_26716,N_23044);
or U30188 (N_30188,N_28051,N_25994);
and U30189 (N_30189,N_27199,N_28123);
nand U30190 (N_30190,N_24002,N_21748);
xnor U30191 (N_30191,N_23911,N_27781);
xnor U30192 (N_30192,N_24978,N_29557);
xor U30193 (N_30193,N_26484,N_26061);
or U30194 (N_30194,N_28589,N_24935);
or U30195 (N_30195,N_26009,N_25180);
and U30196 (N_30196,N_24501,N_24562);
or U30197 (N_30197,N_20454,N_25263);
and U30198 (N_30198,N_29997,N_25969);
nand U30199 (N_30199,N_26439,N_26120);
nand U30200 (N_30200,N_23160,N_24886);
and U30201 (N_30201,N_24315,N_23256);
nor U30202 (N_30202,N_24123,N_20745);
and U30203 (N_30203,N_21510,N_22619);
nand U30204 (N_30204,N_27605,N_24186);
and U30205 (N_30205,N_23737,N_27670);
nand U30206 (N_30206,N_23879,N_24112);
or U30207 (N_30207,N_28397,N_24311);
xor U30208 (N_30208,N_25702,N_21038);
and U30209 (N_30209,N_26524,N_24312);
nor U30210 (N_30210,N_25270,N_25295);
nor U30211 (N_30211,N_25599,N_23785);
nor U30212 (N_30212,N_27282,N_23535);
nand U30213 (N_30213,N_24973,N_28978);
or U30214 (N_30214,N_29100,N_24227);
or U30215 (N_30215,N_20852,N_24793);
xor U30216 (N_30216,N_26650,N_23366);
nand U30217 (N_30217,N_23937,N_25024);
xnor U30218 (N_30218,N_25827,N_22507);
nor U30219 (N_30219,N_28559,N_23820);
xnor U30220 (N_30220,N_27791,N_26185);
xnor U30221 (N_30221,N_29115,N_24906);
or U30222 (N_30222,N_21446,N_27224);
and U30223 (N_30223,N_21639,N_29084);
nand U30224 (N_30224,N_28838,N_23317);
nor U30225 (N_30225,N_29874,N_26670);
and U30226 (N_30226,N_28765,N_28742);
nor U30227 (N_30227,N_24272,N_20632);
nand U30228 (N_30228,N_22228,N_20896);
xnor U30229 (N_30229,N_29055,N_29074);
or U30230 (N_30230,N_24583,N_29861);
nand U30231 (N_30231,N_27365,N_29147);
nand U30232 (N_30232,N_25155,N_28752);
xnor U30233 (N_30233,N_22397,N_26370);
and U30234 (N_30234,N_24399,N_27594);
and U30235 (N_30235,N_29988,N_27552);
nor U30236 (N_30236,N_28577,N_29043);
xnor U30237 (N_30237,N_21355,N_20111);
and U30238 (N_30238,N_22157,N_24231);
and U30239 (N_30239,N_29751,N_22022);
or U30240 (N_30240,N_24199,N_20371);
xor U30241 (N_30241,N_23780,N_20524);
xor U30242 (N_30242,N_21627,N_22351);
nor U30243 (N_30243,N_21314,N_23484);
and U30244 (N_30244,N_20409,N_22192);
nand U30245 (N_30245,N_24120,N_22847);
xor U30246 (N_30246,N_20590,N_26259);
or U30247 (N_30247,N_25095,N_25760);
nor U30248 (N_30248,N_21259,N_21859);
xor U30249 (N_30249,N_24617,N_24512);
xor U30250 (N_30250,N_26888,N_27357);
or U30251 (N_30251,N_26561,N_22717);
or U30252 (N_30252,N_21765,N_25797);
xor U30253 (N_30253,N_28291,N_26964);
or U30254 (N_30254,N_20318,N_25007);
nand U30255 (N_30255,N_21189,N_28855);
nor U30256 (N_30256,N_23572,N_24525);
nand U30257 (N_30257,N_22419,N_20227);
nor U30258 (N_30258,N_25604,N_20659);
and U30259 (N_30259,N_21611,N_29531);
xor U30260 (N_30260,N_28236,N_21767);
nor U30261 (N_30261,N_28405,N_21808);
nor U30262 (N_30262,N_23563,N_24083);
or U30263 (N_30263,N_29916,N_26424);
and U30264 (N_30264,N_27898,N_26129);
xor U30265 (N_30265,N_24949,N_29807);
nor U30266 (N_30266,N_29159,N_25813);
and U30267 (N_30267,N_20872,N_27430);
and U30268 (N_30268,N_22914,N_22386);
or U30269 (N_30269,N_20339,N_20569);
and U30270 (N_30270,N_27509,N_21974);
and U30271 (N_30271,N_24461,N_20440);
nand U30272 (N_30272,N_20283,N_20667);
nor U30273 (N_30273,N_27604,N_25681);
nor U30274 (N_30274,N_23197,N_21012);
and U30275 (N_30275,N_21337,N_25750);
nand U30276 (N_30276,N_24362,N_23955);
nand U30277 (N_30277,N_24705,N_25066);
nand U30278 (N_30278,N_24944,N_21333);
or U30279 (N_30279,N_23177,N_24348);
or U30280 (N_30280,N_21832,N_25879);
and U30281 (N_30281,N_21143,N_24534);
nand U30282 (N_30282,N_26633,N_21235);
and U30283 (N_30283,N_21255,N_25882);
and U30284 (N_30284,N_26631,N_26843);
nor U30285 (N_30285,N_29266,N_23965);
nand U30286 (N_30286,N_26215,N_24989);
xor U30287 (N_30287,N_24789,N_25345);
xor U30288 (N_30288,N_23018,N_29493);
and U30289 (N_30289,N_21951,N_23099);
or U30290 (N_30290,N_25204,N_25217);
and U30291 (N_30291,N_27209,N_23818);
nand U30292 (N_30292,N_25859,N_27826);
nand U30293 (N_30293,N_26691,N_28628);
nand U30294 (N_30294,N_21340,N_26139);
and U30295 (N_30295,N_20814,N_26555);
and U30296 (N_30296,N_26642,N_26873);
nand U30297 (N_30297,N_20974,N_27026);
and U30298 (N_30298,N_21232,N_25421);
and U30299 (N_30299,N_25579,N_23114);
xnor U30300 (N_30300,N_25301,N_22559);
nand U30301 (N_30301,N_21881,N_24001);
or U30302 (N_30302,N_28570,N_21917);
and U30303 (N_30303,N_25435,N_20583);
xor U30304 (N_30304,N_21145,N_29424);
xnor U30305 (N_30305,N_27254,N_23659);
nor U30306 (N_30306,N_29780,N_23467);
and U30307 (N_30307,N_29263,N_23623);
or U30308 (N_30308,N_29135,N_25143);
or U30309 (N_30309,N_24594,N_29593);
and U30310 (N_30310,N_21275,N_27390);
nand U30311 (N_30311,N_24868,N_26945);
and U30312 (N_30312,N_22071,N_28325);
xnor U30313 (N_30313,N_26665,N_28937);
or U30314 (N_30314,N_28907,N_28063);
or U30315 (N_30315,N_27483,N_23863);
and U30316 (N_30316,N_26203,N_27473);
and U30317 (N_30317,N_21251,N_24864);
nor U30318 (N_30318,N_28082,N_23799);
nor U30319 (N_30319,N_27516,N_24076);
xor U30320 (N_30320,N_24597,N_28254);
or U30321 (N_30321,N_20592,N_24485);
nor U30322 (N_30322,N_21531,N_29085);
xor U30323 (N_30323,N_28521,N_22433);
nor U30324 (N_30324,N_21517,N_24679);
xnor U30325 (N_30325,N_28536,N_20834);
or U30326 (N_30326,N_29863,N_21511);
nor U30327 (N_30327,N_27093,N_26292);
nor U30328 (N_30328,N_26381,N_25451);
nor U30329 (N_30329,N_26392,N_26934);
xor U30330 (N_30330,N_29439,N_24818);
nor U30331 (N_30331,N_29758,N_28207);
and U30332 (N_30332,N_29258,N_22947);
nand U30333 (N_30333,N_21730,N_23049);
or U30334 (N_30334,N_22148,N_26467);
or U30335 (N_30335,N_27593,N_25352);
and U30336 (N_30336,N_29708,N_23793);
or U30337 (N_30337,N_28955,N_20384);
xor U30338 (N_30338,N_29487,N_22164);
xor U30339 (N_30339,N_25141,N_28342);
nor U30340 (N_30340,N_25782,N_23696);
xnor U30341 (N_30341,N_21863,N_24160);
xor U30342 (N_30342,N_20221,N_20750);
or U30343 (N_30343,N_25057,N_20619);
nor U30344 (N_30344,N_22045,N_27157);
or U30345 (N_30345,N_20438,N_20598);
xor U30346 (N_30346,N_22755,N_28129);
and U30347 (N_30347,N_26440,N_20850);
nand U30348 (N_30348,N_29587,N_27891);
and U30349 (N_30349,N_28212,N_22259);
and U30350 (N_30350,N_26454,N_29940);
nor U30351 (N_30351,N_22182,N_26419);
or U30352 (N_30352,N_23574,N_22667);
nand U30353 (N_30353,N_28776,N_22499);
nor U30354 (N_30354,N_20980,N_22502);
xnor U30355 (N_30355,N_27912,N_27472);
and U30356 (N_30356,N_24330,N_29872);
nand U30357 (N_30357,N_20558,N_23688);
nor U30358 (N_30358,N_28947,N_26833);
and U30359 (N_30359,N_29528,N_25715);
nor U30360 (N_30360,N_26726,N_28015);
nor U30361 (N_30361,N_29244,N_29448);
or U30362 (N_30362,N_21667,N_28340);
nor U30363 (N_30363,N_26137,N_21911);
xnor U30364 (N_30364,N_29887,N_26189);
nor U30365 (N_30365,N_28036,N_20919);
or U30366 (N_30366,N_27457,N_23619);
and U30367 (N_30367,N_28406,N_22319);
nand U30368 (N_30368,N_28348,N_22997);
nand U30369 (N_30369,N_28491,N_21772);
nand U30370 (N_30370,N_26625,N_25525);
xor U30371 (N_30371,N_23599,N_20546);
nor U30372 (N_30372,N_27824,N_25615);
xnor U30373 (N_30373,N_22367,N_20586);
nand U30374 (N_30374,N_27314,N_25706);
nand U30375 (N_30375,N_23062,N_21410);
nor U30376 (N_30376,N_23393,N_25179);
xnor U30377 (N_30377,N_22868,N_22820);
nand U30378 (N_30378,N_21434,N_29743);
nand U30379 (N_30379,N_23096,N_27562);
and U30380 (N_30380,N_21552,N_25202);
and U30381 (N_30381,N_24577,N_26164);
or U30382 (N_30382,N_24470,N_27788);
xnor U30383 (N_30383,N_21977,N_23052);
nand U30384 (N_30384,N_22373,N_21770);
or U30385 (N_30385,N_28166,N_21814);
nand U30386 (N_30386,N_26298,N_22462);
and U30387 (N_30387,N_26821,N_24088);
nor U30388 (N_30388,N_27198,N_24027);
nor U30389 (N_30389,N_22650,N_26731);
nand U30390 (N_30390,N_23839,N_27097);
nand U30391 (N_30391,N_21934,N_22423);
or U30392 (N_30392,N_21339,N_26861);
xnor U30393 (N_30393,N_22834,N_22322);
nand U30394 (N_30394,N_24317,N_25612);
nor U30395 (N_30395,N_25186,N_24073);
xnor U30396 (N_30396,N_23159,N_28535);
xnor U30397 (N_30397,N_26719,N_25934);
and U30398 (N_30398,N_25469,N_20344);
xnor U30399 (N_30399,N_20249,N_24026);
and U30400 (N_30400,N_29597,N_27351);
or U30401 (N_30401,N_21008,N_20254);
nand U30402 (N_30402,N_29262,N_27029);
xor U30403 (N_30403,N_26287,N_26455);
and U30404 (N_30404,N_23038,N_26435);
and U30405 (N_30405,N_23102,N_29711);
and U30406 (N_30406,N_25950,N_25617);
xnor U30407 (N_30407,N_21836,N_27235);
nor U30408 (N_30408,N_24756,N_22356);
nand U30409 (N_30409,N_24293,N_29213);
xnor U30410 (N_30410,N_26700,N_28664);
and U30411 (N_30411,N_24058,N_29333);
and U30412 (N_30412,N_29968,N_20818);
xnor U30413 (N_30413,N_22899,N_26380);
or U30414 (N_30414,N_20908,N_24922);
nand U30415 (N_30415,N_29680,N_23988);
and U30416 (N_30416,N_27775,N_20873);
or U30417 (N_30417,N_28045,N_28605);
nand U30418 (N_30418,N_25896,N_24628);
or U30419 (N_30419,N_26002,N_22907);
nor U30420 (N_30420,N_23061,N_25014);
xnor U30421 (N_30421,N_26224,N_27252);
and U30422 (N_30422,N_24531,N_21868);
xor U30423 (N_30423,N_26079,N_21597);
nor U30424 (N_30424,N_25505,N_22987);
and U30425 (N_30425,N_20754,N_24420);
or U30426 (N_30426,N_24857,N_26567);
or U30427 (N_30427,N_22227,N_22337);
xnor U30428 (N_30428,N_21901,N_20204);
xnor U30429 (N_30429,N_23111,N_29336);
xor U30430 (N_30430,N_21645,N_21690);
nand U30431 (N_30431,N_26456,N_29748);
and U30432 (N_30432,N_22044,N_25798);
xor U30433 (N_30433,N_24842,N_25954);
nand U30434 (N_30434,N_24042,N_20932);
xor U30435 (N_30435,N_21354,N_22034);
nand U30436 (N_30436,N_29435,N_29480);
or U30437 (N_30437,N_20314,N_27372);
nand U30438 (N_30438,N_25508,N_23048);
or U30439 (N_30439,N_27606,N_20728);
xnor U30440 (N_30440,N_27799,N_28415);
xor U30441 (N_30441,N_24914,N_21473);
xnor U30442 (N_30442,N_25719,N_21580);
xor U30443 (N_30443,N_22989,N_20205);
nand U30444 (N_30444,N_21570,N_29267);
or U30445 (N_30445,N_23266,N_28571);
and U30446 (N_30446,N_29744,N_20142);
or U30447 (N_30447,N_20395,N_20963);
xnor U30448 (N_30448,N_22844,N_20135);
and U30449 (N_30449,N_26344,N_28539);
and U30450 (N_30450,N_26149,N_27106);
nand U30451 (N_30451,N_27385,N_20009);
nor U30452 (N_30452,N_29384,N_21579);
xnor U30453 (N_30453,N_25801,N_27712);
and U30454 (N_30454,N_25970,N_29605);
nand U30455 (N_30455,N_25660,N_25958);
and U30456 (N_30456,N_22258,N_29381);
nor U30457 (N_30457,N_27036,N_28394);
and U30458 (N_30458,N_20979,N_24095);
xor U30459 (N_30459,N_23960,N_24113);
nand U30460 (N_30460,N_26959,N_21106);
and U30461 (N_30461,N_28202,N_23475);
or U30462 (N_30462,N_25860,N_24237);
nor U30463 (N_30463,N_20363,N_27767);
or U30464 (N_30464,N_25058,N_28412);
or U30465 (N_30465,N_26486,N_24900);
and U30466 (N_30466,N_24606,N_27249);
xor U30467 (N_30467,N_27088,N_28178);
xnor U30468 (N_30468,N_28502,N_29101);
nand U30469 (N_30469,N_21986,N_26754);
nor U30470 (N_30470,N_27347,N_29892);
and U30471 (N_30471,N_22566,N_28717);
or U30472 (N_30472,N_20515,N_25603);
nand U30473 (N_30473,N_22437,N_26501);
xor U30474 (N_30474,N_29169,N_27227);
nor U30475 (N_30475,N_20916,N_28611);
or U30476 (N_30476,N_22274,N_26141);
and U30477 (N_30477,N_24713,N_21180);
and U30478 (N_30478,N_20336,N_22307);
xnor U30479 (N_30479,N_25668,N_23661);
xnor U30480 (N_30480,N_29466,N_20241);
xor U30481 (N_30481,N_21268,N_28500);
and U30482 (N_30482,N_23981,N_29081);
nor U30483 (N_30483,N_20076,N_29847);
nor U30484 (N_30484,N_28727,N_22435);
and U30485 (N_30485,N_21176,N_20008);
nand U30486 (N_30486,N_25026,N_21966);
or U30487 (N_30487,N_27167,N_25808);
nand U30488 (N_30488,N_21961,N_23005);
or U30489 (N_30489,N_23452,N_29926);
nor U30490 (N_30490,N_23985,N_29732);
xnor U30491 (N_30491,N_27031,N_21278);
nor U30492 (N_30492,N_27066,N_29034);
or U30493 (N_30493,N_21140,N_28738);
nand U30494 (N_30494,N_22855,N_20679);
or U30495 (N_30495,N_24687,N_22230);
or U30496 (N_30496,N_24331,N_28783);
nor U30497 (N_30497,N_22919,N_22364);
or U30498 (N_30498,N_24968,N_27129);
nor U30499 (N_30499,N_23512,N_21385);
xor U30500 (N_30500,N_22078,N_28290);
and U30501 (N_30501,N_24953,N_27825);
and U30502 (N_30502,N_26892,N_25063);
xnor U30503 (N_30503,N_22116,N_28774);
nand U30504 (N_30504,N_28657,N_27926);
xnor U30505 (N_30505,N_29467,N_27865);
or U30506 (N_30506,N_23108,N_26673);
and U30507 (N_30507,N_20714,N_29407);
xor U30508 (N_30508,N_22904,N_24714);
nand U30509 (N_30509,N_23683,N_29265);
and U30510 (N_30510,N_25769,N_27906);
and U30511 (N_30511,N_26289,N_22570);
or U30512 (N_30512,N_20421,N_20543);
nor U30513 (N_30513,N_28851,N_27193);
nor U30514 (N_30514,N_27265,N_21889);
nor U30515 (N_30515,N_21222,N_27676);
nor U30516 (N_30516,N_21835,N_29709);
or U30517 (N_30517,N_23707,N_23933);
nor U30518 (N_30518,N_29446,N_28820);
nor U30519 (N_30519,N_23980,N_26573);
and U30520 (N_30520,N_25369,N_26741);
or U30521 (N_30521,N_24712,N_26418);
nor U30522 (N_30522,N_23476,N_26049);
and U30523 (N_30523,N_24242,N_28383);
nor U30524 (N_30524,N_22114,N_22783);
or U30525 (N_30525,N_26374,N_26369);
or U30526 (N_30526,N_20623,N_23629);
or U30527 (N_30527,N_26494,N_29719);
nor U30528 (N_30528,N_23872,N_24673);
or U30529 (N_30529,N_26428,N_25132);
nand U30530 (N_30530,N_29508,N_23354);
nor U30531 (N_30531,N_28833,N_24623);
nor U30532 (N_30532,N_23122,N_29226);
nand U30533 (N_30533,N_29064,N_28639);
or U30534 (N_30534,N_29613,N_26150);
nand U30535 (N_30535,N_26509,N_25243);
and U30536 (N_30536,N_24390,N_26204);
xor U30537 (N_30537,N_20882,N_20936);
or U30538 (N_30538,N_27887,N_26668);
xor U30539 (N_30539,N_24795,N_26293);
xnor U30540 (N_30540,N_28874,N_24884);
or U30541 (N_30541,N_21306,N_27264);
or U30542 (N_30542,N_26116,N_23527);
xor U30543 (N_30543,N_25527,N_29361);
xor U30544 (N_30544,N_20624,N_22421);
xor U30545 (N_30545,N_23795,N_22239);
and U30546 (N_30546,N_26637,N_21096);
xnor U30547 (N_30547,N_23966,N_28130);
xor U30548 (N_30548,N_27678,N_21753);
and U30549 (N_30549,N_24308,N_23833);
nor U30550 (N_30550,N_26960,N_29498);
xor U30551 (N_30551,N_22235,N_27152);
and U30552 (N_30552,N_23310,N_27624);
nor U30553 (N_30553,N_27187,N_29880);
xnor U30554 (N_30554,N_29614,N_26044);
nor U30555 (N_30555,N_29248,N_25914);
nor U30556 (N_30556,N_25034,N_20035);
nor U30557 (N_30557,N_27735,N_21046);
and U30558 (N_30558,N_25436,N_26426);
nand U30559 (N_30559,N_23334,N_21624);
xnor U30560 (N_30560,N_27188,N_29345);
nor U30561 (N_30561,N_23951,N_25776);
nor U30562 (N_30562,N_27319,N_26588);
nand U30563 (N_30563,N_27397,N_23625);
nor U30564 (N_30564,N_28251,N_29315);
xor U30565 (N_30565,N_20105,N_24119);
and U30566 (N_30566,N_24285,N_20004);
nor U30567 (N_30567,N_21789,N_23262);
xnor U30568 (N_30568,N_20264,N_24249);
nand U30569 (N_30569,N_23501,N_23339);
nor U30570 (N_30570,N_26165,N_28370);
xor U30571 (N_30571,N_25227,N_22272);
nor U30572 (N_30572,N_23559,N_23942);
and U30573 (N_30573,N_29395,N_21377);
xnor U30574 (N_30574,N_27937,N_25059);
and U30575 (N_30575,N_20698,N_20128);
or U30576 (N_30576,N_26286,N_28020);
xor U30577 (N_30577,N_29046,N_24690);
nand U30578 (N_30578,N_25306,N_26263);
nand U30579 (N_30579,N_25150,N_23544);
xor U30580 (N_30580,N_29991,N_24046);
and U30581 (N_30581,N_22434,N_21542);
nand U30582 (N_30582,N_26483,N_27922);
and U30583 (N_30583,N_23973,N_24903);
nor U30584 (N_30584,N_22326,N_25805);
nor U30585 (N_30585,N_25581,N_22590);
xnor U30586 (N_30586,N_23609,N_28220);
nor U30587 (N_30587,N_21382,N_28988);
and U30588 (N_30588,N_27266,N_22517);
nand U30589 (N_30589,N_22934,N_25249);
xnor U30590 (N_30590,N_22951,N_23386);
nor U30591 (N_30591,N_27782,N_20502);
nand U30592 (N_30592,N_29260,N_20731);
or U30593 (N_30593,N_26282,N_24622);
xnor U30594 (N_30594,N_28799,N_27795);
or U30595 (N_30595,N_24588,N_29817);
xor U30596 (N_30596,N_28449,N_29596);
xor U30597 (N_30597,N_20379,N_28352);
nor U30598 (N_30598,N_23307,N_21183);
xor U30599 (N_30599,N_21016,N_24077);
xor U30600 (N_30600,N_28304,N_27728);
nor U30601 (N_30601,N_22712,N_21718);
nand U30602 (N_30602,N_22702,N_22174);
and U30603 (N_30603,N_29496,N_21878);
nor U30604 (N_30604,N_20704,N_28695);
or U30605 (N_30605,N_20029,N_21196);
xor U30606 (N_30606,N_28550,N_20239);
xor U30607 (N_30607,N_24981,N_23054);
xnor U30608 (N_30608,N_22371,N_29921);
nor U30609 (N_30609,N_25284,N_27770);
nand U30610 (N_30610,N_21206,N_24491);
and U30611 (N_30611,N_26544,N_20373);
nand U30612 (N_30612,N_24126,N_23066);
nand U30613 (N_30613,N_22302,N_24725);
xor U30614 (N_30614,N_24010,N_20377);
xor U30615 (N_30615,N_23079,N_22807);
nand U30616 (N_30616,N_27729,N_27827);
xnor U30617 (N_30617,N_25234,N_25758);
nor U30618 (N_30618,N_21087,N_23149);
and U30619 (N_30619,N_27244,N_28533);
nand U30620 (N_30620,N_27480,N_24271);
xor U30621 (N_30621,N_24974,N_20837);
and U30622 (N_30622,N_20999,N_26751);
nand U30623 (N_30623,N_26968,N_26091);
nand U30624 (N_30624,N_22678,N_25433);
xor U30625 (N_30625,N_29812,N_21302);
and U30626 (N_30626,N_26133,N_21364);
and U30627 (N_30627,N_28001,N_27146);
or U30628 (N_30628,N_22335,N_27038);
or U30629 (N_30629,N_21949,N_27095);
and U30630 (N_30630,N_27931,N_21469);
nand U30631 (N_30631,N_29460,N_29177);
nand U30632 (N_30632,N_25319,N_26558);
xnor U30633 (N_30633,N_25031,N_23080);
nor U30634 (N_30634,N_20462,N_21486);
or U30635 (N_30635,N_22952,N_21250);
xor U30636 (N_30636,N_28508,N_23237);
and U30637 (N_30637,N_26318,N_29080);
xor U30638 (N_30638,N_24860,N_27330);
and U30639 (N_30639,N_21203,N_21168);
xor U30640 (N_30640,N_26745,N_23324);
nor U30641 (N_30641,N_20939,N_26411);
nor U30642 (N_30642,N_22185,N_23704);
xor U30643 (N_30643,N_24326,N_26771);
xor U30644 (N_30644,N_29949,N_26748);
or U30645 (N_30645,N_20459,N_28294);
nor U30646 (N_30646,N_26860,N_27673);
or U30647 (N_30647,N_27543,N_21637);
and U30648 (N_30648,N_23552,N_22278);
nand U30649 (N_30649,N_23890,N_23945);
nand U30650 (N_30650,N_26267,N_28532);
nand U30651 (N_30651,N_22571,N_20989);
xor U30652 (N_30652,N_27343,N_27840);
nor U30653 (N_30653,N_27274,N_27707);
nor U30654 (N_30654,N_27484,N_29985);
or U30655 (N_30655,N_22204,N_23417);
xnor U30656 (N_30656,N_24252,N_29954);
and U30657 (N_30657,N_29388,N_20247);
or U30658 (N_30658,N_21361,N_25134);
xor U30659 (N_30659,N_29239,N_23944);
nand U30660 (N_30660,N_25621,N_25003);
or U30661 (N_30661,N_29037,N_29130);
or U30662 (N_30662,N_26361,N_25476);
and U30663 (N_30663,N_28441,N_28054);
xnor U30664 (N_30664,N_28237,N_28740);
nand U30665 (N_30665,N_28852,N_22611);
xnor U30666 (N_30666,N_28418,N_24529);
or U30667 (N_30667,N_20298,N_28486);
nand U30668 (N_30668,N_27718,N_26760);
nand U30669 (N_30669,N_29622,N_24314);
nand U30670 (N_30670,N_29344,N_27040);
or U30671 (N_30671,N_29547,N_21621);
nand U30672 (N_30672,N_21640,N_24462);
xor U30673 (N_30673,N_20222,N_25937);
nand U30674 (N_30674,N_29289,N_28823);
or U30675 (N_30675,N_26566,N_27460);
or U30676 (N_30676,N_26226,N_23202);
and U30677 (N_30677,N_21561,N_28856);
or U30678 (N_30678,N_22265,N_26337);
xor U30679 (N_30679,N_27124,N_23626);
and U30680 (N_30680,N_20027,N_23925);
nand U30681 (N_30681,N_21215,N_24294);
nand U30682 (N_30682,N_23595,N_22445);
and U30683 (N_30683,N_23063,N_24425);
and U30684 (N_30684,N_20032,N_22999);
xnor U30685 (N_30685,N_27464,N_21506);
or U30686 (N_30686,N_20305,N_29562);
xor U30687 (N_30687,N_23729,N_29914);
or U30688 (N_30688,N_29324,N_24576);
nor U30689 (N_30689,N_25366,N_25042);
and U30690 (N_30690,N_23687,N_24437);
nor U30691 (N_30691,N_22122,N_20923);
nand U30692 (N_30692,N_23835,N_23251);
nand U30693 (N_30693,N_28591,N_28199);
or U30694 (N_30694,N_26258,N_21631);
xnor U30695 (N_30695,N_21272,N_23390);
nor U30696 (N_30696,N_26097,N_27440);
nor U30697 (N_30697,N_20321,N_24267);
and U30698 (N_30698,N_28873,N_27518);
or U30699 (N_30699,N_24148,N_26417);
nand U30700 (N_30700,N_23423,N_25183);
xnor U30701 (N_30701,N_25300,N_21670);
or U30702 (N_30702,N_28527,N_21829);
nor U30703 (N_30703,N_23889,N_29560);
nand U30704 (N_30704,N_28763,N_28844);
xnor U30705 (N_30705,N_24329,N_23196);
or U30706 (N_30706,N_28623,N_22486);
nand U30707 (N_30707,N_23996,N_28277);
or U30708 (N_30708,N_27541,N_27339);
nor U30709 (N_30709,N_25147,N_27590);
and U30710 (N_30710,N_21649,N_28546);
xor U30711 (N_30711,N_20699,N_29969);
nor U30712 (N_30712,N_22070,N_28160);
xnor U30713 (N_30713,N_29403,N_29561);
or U30714 (N_30714,N_29158,N_21940);
xor U30715 (N_30715,N_27371,N_23125);
or U30716 (N_30716,N_24572,N_21238);
xor U30717 (N_30717,N_21964,N_25391);
and U30718 (N_30718,N_24091,N_21546);
xnor U30719 (N_30719,N_29903,N_25502);
xor U30720 (N_30720,N_26632,N_26448);
or U30721 (N_30721,N_29053,N_22589);
or U30722 (N_30722,N_28337,N_21816);
or U30723 (N_30723,N_24023,N_26855);
nor U30724 (N_30724,N_28641,N_20646);
nand U30725 (N_30725,N_29944,N_24133);
xor U30726 (N_30726,N_29362,N_26651);
and U30727 (N_30727,N_29272,N_26170);
nand U30728 (N_30728,N_20877,N_27363);
or U30729 (N_30729,N_21501,N_26827);
and U30730 (N_30730,N_26675,N_24599);
or U30731 (N_30731,N_28673,N_28126);
nor U30732 (N_30732,N_22867,N_21701);
nor U30733 (N_30733,N_22393,N_22975);
and U30734 (N_30734,N_26750,N_28520);
or U30735 (N_30735,N_23650,N_27467);
or U30736 (N_30736,N_22330,N_22313);
nor U30737 (N_30737,N_29402,N_24009);
nor U30738 (N_30738,N_24080,N_26474);
nor U30739 (N_30739,N_27854,N_24569);
xor U30740 (N_30740,N_23621,N_25845);
or U30741 (N_30741,N_28132,N_25658);
and U30742 (N_30742,N_21378,N_25926);
or U30743 (N_30743,N_23811,N_28003);
and U30744 (N_30744,N_21946,N_20744);
or U30745 (N_30745,N_25645,N_28420);
and U30746 (N_30746,N_22565,N_24648);
nor U30747 (N_30747,N_25756,N_24570);
and U30748 (N_30748,N_28163,N_21558);
or U30749 (N_30749,N_28881,N_28227);
xor U30750 (N_30750,N_24555,N_22720);
xor U30751 (N_30751,N_25559,N_27165);
nor U30752 (N_30752,N_23908,N_28283);
and U30753 (N_30753,N_21984,N_24739);
xnor U30754 (N_30754,N_20831,N_29958);
or U30755 (N_30755,N_20015,N_29018);
nand U30756 (N_30756,N_27632,N_29172);
xor U30757 (N_30757,N_24365,N_20912);
or U30758 (N_30758,N_25996,N_22615);
nand U30759 (N_30759,N_22646,N_21959);
xnor U30760 (N_30760,N_27113,N_21729);
nor U30761 (N_30761,N_20952,N_25745);
or U30762 (N_30762,N_24368,N_29112);
xor U30763 (N_30763,N_28087,N_23772);
and U30764 (N_30764,N_21178,N_20996);
or U30765 (N_30765,N_24201,N_28164);
nand U30766 (N_30766,N_26319,N_21458);
xor U30767 (N_30767,N_22067,N_27568);
nand U30768 (N_30768,N_28575,N_29616);
and U30769 (N_30769,N_21860,N_29856);
nor U30770 (N_30770,N_26903,N_29741);
xnor U30771 (N_30771,N_26911,N_25552);
and U30772 (N_30772,N_27323,N_20568);
nor U30773 (N_30773,N_24680,N_21027);
nor U30774 (N_30774,N_27099,N_29848);
and U30775 (N_30775,N_29876,N_25566);
xor U30776 (N_30776,N_24828,N_27257);
nand U30777 (N_30777,N_24067,N_21983);
nor U30778 (N_30778,N_23505,N_25631);
nand U30779 (N_30779,N_22375,N_24419);
xor U30780 (N_30780,N_28416,N_27919);
and U30781 (N_30781,N_24574,N_26970);
nand U30782 (N_30782,N_20982,N_29217);
or U30783 (N_30783,N_24367,N_23064);
or U30784 (N_30784,N_23253,N_28530);
or U30785 (N_30785,N_21551,N_28946);
or U30786 (N_30786,N_26415,N_26824);
or U30787 (N_30787,N_29246,N_28173);
nand U30788 (N_30788,N_21045,N_24548);
nor U30789 (N_30789,N_22196,N_24778);
xor U30790 (N_30790,N_23469,N_25815);
nand U30791 (N_30791,N_26399,N_21461);
and U30792 (N_30792,N_23245,N_21660);
and U30793 (N_30793,N_26042,N_20510);
nand U30794 (N_30794,N_21919,N_25348);
nand U30795 (N_30795,N_23078,N_29302);
and U30796 (N_30796,N_25911,N_25431);
nor U30797 (N_30797,N_26146,N_24356);
nor U30798 (N_30798,N_27741,N_24079);
nand U30799 (N_30799,N_29559,N_24636);
nor U30800 (N_30800,N_28219,N_25235);
or U30801 (N_30801,N_25323,N_22529);
nand U30802 (N_30802,N_22708,N_21749);
nand U30803 (N_30803,N_22766,N_28438);
and U30804 (N_30804,N_26610,N_25201);
nor U30805 (N_30805,N_29481,N_27080);
nand U30806 (N_30806,N_26505,N_28414);
nor U30807 (N_30807,N_21602,N_28603);
or U30808 (N_30808,N_20553,N_25596);
nand U30809 (N_30809,N_21015,N_25574);
xor U30810 (N_30810,N_23297,N_24938);
nor U30811 (N_30811,N_26121,N_23947);
or U30812 (N_30812,N_24025,N_22595);
nand U30813 (N_30813,N_24736,N_21450);
xnor U30814 (N_30814,N_25877,N_22018);
nor U30815 (N_30815,N_22218,N_25704);
nand U30816 (N_30816,N_24277,N_26788);
and U30817 (N_30817,N_22779,N_29288);
or U30818 (N_30818,N_20784,N_29690);
nand U30819 (N_30819,N_22814,N_28146);
or U30820 (N_30820,N_20966,N_27626);
nand U30821 (N_30821,N_23550,N_21894);
xor U30822 (N_30822,N_26240,N_23466);
or U30823 (N_30823,N_23332,N_22402);
and U30824 (N_30824,N_22273,N_20602);
or U30825 (N_30825,N_26227,N_29546);
xor U30826 (N_30826,N_29992,N_21857);
xnor U30827 (N_30827,N_29618,N_22483);
or U30828 (N_30828,N_24563,N_25679);
or U30829 (N_30829,N_23384,N_20474);
xor U30830 (N_30830,N_23259,N_23598);
or U30831 (N_30831,N_23184,N_22300);
xnor U30832 (N_30832,N_22731,N_25844);
xnor U30833 (N_30833,N_29307,N_24658);
nor U30834 (N_30834,N_21941,N_20701);
xnor U30835 (N_30835,N_23622,N_22465);
or U30836 (N_30836,N_29401,N_22922);
or U30837 (N_30837,N_29620,N_26813);
and U30838 (N_30838,N_27834,N_26111);
nand U30839 (N_30839,N_22285,N_28137);
nand U30840 (N_30840,N_28124,N_20091);
xnor U30841 (N_30841,N_20172,N_24589);
and U30842 (N_30842,N_23620,N_28501);
nand U30843 (N_30843,N_28723,N_23646);
or U30844 (N_30844,N_24433,N_28471);
xor U30845 (N_30845,N_23668,N_22461);
or U30846 (N_30846,N_26174,N_27119);
or U30847 (N_30847,N_23551,N_28159);
nand U30848 (N_30848,N_20636,N_25347);
xor U30849 (N_30849,N_26902,N_26391);
and U30850 (N_30850,N_28726,N_22111);
nor U30851 (N_30851,N_29774,N_29041);
or U30852 (N_30852,N_23329,N_29655);
xor U30853 (N_30853,N_25597,N_28216);
or U30854 (N_30854,N_22244,N_20077);
nand U30855 (N_30855,N_22138,N_29507);
nor U30856 (N_30856,N_26772,N_23794);
or U30857 (N_30857,N_25639,N_22059);
nand U30858 (N_30858,N_29327,N_23657);
or U30859 (N_30859,N_27288,N_28208);
nand U30860 (N_30860,N_24416,N_22796);
and U30861 (N_30861,N_21489,N_29803);
nor U30862 (N_30862,N_21766,N_24645);
nor U30863 (N_30863,N_25136,N_22058);
or U30864 (N_30864,N_27588,N_26661);
xnor U30865 (N_30865,N_27655,N_21467);
nor U30866 (N_30866,N_20910,N_29086);
nor U30867 (N_30867,N_26277,N_28086);
xnor U30868 (N_30868,N_27130,N_25537);
nand U30869 (N_30869,N_29626,N_27643);
and U30870 (N_30870,N_20726,N_21000);
or U30871 (N_30871,N_20393,N_22818);
nor U30872 (N_30872,N_29627,N_20503);
or U30873 (N_30873,N_25404,N_21041);
and U30874 (N_30874,N_29716,N_23385);
xnor U30875 (N_30875,N_28654,N_21853);
nor U30876 (N_30876,N_28958,N_27222);
nor U30877 (N_30877,N_24954,N_29163);
and U30878 (N_30878,N_28041,N_28391);
nand U30879 (N_30879,N_28377,N_27984);
xnor U30880 (N_30880,N_27219,N_27013);
xnor U30881 (N_30881,N_27074,N_25640);
and U30882 (N_30882,N_20085,N_22887);
or U30883 (N_30883,N_20131,N_20573);
and U30884 (N_30884,N_26015,N_24408);
nand U30885 (N_30885,N_20763,N_22120);
and U30886 (N_30886,N_20517,N_20964);
nor U30887 (N_30887,N_28901,N_20868);
nor U30888 (N_30888,N_23059,N_25448);
and U30889 (N_30889,N_26358,N_26652);
or U30890 (N_30890,N_21734,N_27710);
nor U30891 (N_30891,N_22401,N_29866);
nand U30892 (N_30892,N_26271,N_26306);
xnor U30893 (N_30893,N_25304,N_28301);
nand U30894 (N_30894,N_24890,N_25402);
or U30895 (N_30895,N_22664,N_27148);
or U30896 (N_30896,N_20294,N_26924);
xnor U30897 (N_30897,N_23376,N_26034);
nand U30898 (N_30898,N_21751,N_28850);
and U30899 (N_30899,N_24166,N_29413);
nor U30900 (N_30900,N_28407,N_22458);
xor U30901 (N_30901,N_20490,N_20053);
nand U30902 (N_30902,N_28879,N_29022);
nor U30903 (N_30903,N_29504,N_29123);
xor U30904 (N_30904,N_28810,N_20473);
nor U30905 (N_30905,N_20260,N_20519);
nor U30906 (N_30906,N_28653,N_28050);
and U30907 (N_30907,N_21654,N_24702);
nand U30908 (N_30908,N_22756,N_20168);
or U30909 (N_30909,N_25011,N_20956);
nand U30910 (N_30910,N_20070,N_21350);
or U30911 (N_30911,N_23892,N_29122);
xor U30912 (N_30912,N_28506,N_26387);
nor U30913 (N_30913,N_25223,N_23363);
or U30914 (N_30914,N_27158,N_20181);
xor U30915 (N_30915,N_21852,N_23301);
xnor U30916 (N_30916,N_21440,N_27719);
nand U30917 (N_30917,N_23689,N_25558);
nor U30918 (N_30918,N_28460,N_25158);
nand U30919 (N_30919,N_25149,N_29957);
nand U30920 (N_30920,N_21249,N_23015);
nand U30921 (N_30921,N_20182,N_27486);
nor U30922 (N_30922,N_24423,N_28691);
nand U30923 (N_30923,N_20954,N_20280);
or U30924 (N_30924,N_24893,N_23666);
nand U30925 (N_30925,N_26294,N_22964);
nand U30926 (N_30926,N_26956,N_22443);
and U30927 (N_30927,N_25357,N_27794);
xnor U30928 (N_30928,N_24492,N_28176);
and U30929 (N_30929,N_22123,N_29092);
xnor U30930 (N_30930,N_23819,N_22057);
and U30931 (N_30931,N_26512,N_27849);
nor U30932 (N_30932,N_23103,N_20410);
and U30933 (N_30933,N_24450,N_27120);
nand U30934 (N_30934,N_27230,N_28140);
and U30935 (N_30935,N_21846,N_22232);
nor U30936 (N_30936,N_21768,N_22670);
nor U30937 (N_30937,N_26490,N_25998);
xor U30938 (N_30938,N_28600,N_24276);
or U30939 (N_30939,N_27225,N_26210);
or U30940 (N_30940,N_28974,N_26639);
and U30941 (N_30941,N_22669,N_24915);
nand U30942 (N_30942,N_28221,N_22798);
or U30943 (N_30943,N_20962,N_27162);
and U30944 (N_30944,N_28809,N_23728);
nor U30945 (N_30945,N_28883,N_23487);
xnor U30946 (N_30946,N_26143,N_20780);
or U30947 (N_30947,N_20904,N_29686);
or U30948 (N_30948,N_29077,N_22075);
nand U30949 (N_30949,N_21280,N_22519);
nor U30950 (N_30950,N_23034,N_21011);
nor U30951 (N_30951,N_24436,N_29078);
xor U30952 (N_30952,N_21316,N_20362);
or U30953 (N_30953,N_22154,N_23648);
nand U30954 (N_30954,N_25342,N_29963);
and U30955 (N_30955,N_24780,N_24808);
nand U30956 (N_30956,N_24243,N_23283);
nor U30957 (N_30957,N_23876,N_28194);
or U30958 (N_30958,N_27369,N_22055);
nor U30959 (N_30959,N_25240,N_23843);
and U30960 (N_30960,N_26963,N_26323);
or U30961 (N_30961,N_28453,N_21876);
or U30962 (N_30962,N_27730,N_26342);
xnor U30963 (N_30963,N_29421,N_26950);
nor U30964 (N_30964,N_29422,N_29296);
nand U30965 (N_30965,N_20277,N_24976);
or U30966 (N_30966,N_25985,N_24473);
or U30967 (N_30967,N_29156,N_27005);
nand U30968 (N_30968,N_23978,N_29231);
or U30969 (N_30969,N_28127,N_20516);
xnor U30970 (N_30970,N_20844,N_27862);
nand U30971 (N_30971,N_26067,N_26191);
nand U30972 (N_30972,N_25140,N_20445);
or U30973 (N_30973,N_23888,N_21883);
nand U30974 (N_30974,N_23531,N_29451);
or U30975 (N_30975,N_23398,N_22527);
or U30976 (N_30976,N_22673,N_21435);
xnor U30977 (N_30977,N_25438,N_27246);
nand U30978 (N_30978,N_27658,N_23961);
or U30979 (N_30979,N_21125,N_20867);
nand U30980 (N_30980,N_21136,N_21167);
nand U30981 (N_30981,N_28021,N_20196);
or U30982 (N_30982,N_27948,N_28476);
nand U30983 (N_30983,N_27537,N_24007);
xor U30984 (N_30984,N_21040,N_29826);
xor U30985 (N_30985,N_23083,N_23458);
or U30986 (N_30986,N_21804,N_26171);
nor U30987 (N_30987,N_21674,N_28758);
xnor U30988 (N_30988,N_21741,N_20235);
nand U30989 (N_30989,N_26013,N_29955);
and U30990 (N_30990,N_23472,N_20588);
and U30991 (N_30991,N_25610,N_27991);
nor U30992 (N_30992,N_26893,N_26249);
xor U30993 (N_30993,N_29523,N_28853);
or U30994 (N_30994,N_23806,N_21014);
xor U30995 (N_30995,N_26069,N_28885);
and U30996 (N_30996,N_28519,N_20571);
nor U30997 (N_30997,N_29933,N_21279);
or U30998 (N_30998,N_23643,N_24800);
and U30999 (N_30999,N_28466,N_20040);
xnor U31000 (N_31000,N_21777,N_27725);
nand U31001 (N_31001,N_26952,N_28223);
or U31002 (N_31002,N_27745,N_26403);
nand U31003 (N_31003,N_29406,N_24991);
or U31004 (N_31004,N_23760,N_21420);
nand U31005 (N_31005,N_20734,N_25689);
xor U31006 (N_31006,N_29990,N_28271);
nor U31007 (N_31007,N_26869,N_22098);
xnor U31008 (N_31008,N_28093,N_24523);
nor U31009 (N_31009,N_26409,N_27171);
nor U31010 (N_31010,N_20906,N_28296);
or U31011 (N_31011,N_29321,N_26167);
nand U31012 (N_31012,N_24851,N_26817);
and U31013 (N_31013,N_23396,N_20600);
nor U31014 (N_31014,N_27979,N_26724);
nand U31015 (N_31015,N_21837,N_24719);
nand U31016 (N_31016,N_24682,N_29697);
nand U31017 (N_31017,N_25355,N_21408);
nand U31018 (N_31018,N_26269,N_26030);
or U31019 (N_31019,N_28599,N_28593);
nand U31020 (N_31020,N_26744,N_24475);
nand U31021 (N_31021,N_23172,N_21069);
nand U31022 (N_31022,N_27961,N_29347);
nor U31023 (N_31023,N_28165,N_26729);
and U31024 (N_31024,N_25416,N_23718);
nor U31025 (N_31025,N_25648,N_20050);
or U31026 (N_31026,N_28669,N_25486);
nand U31027 (N_31027,N_29656,N_28979);
or U31028 (N_31028,N_25297,N_26348);
nand U31029 (N_31029,N_29815,N_21508);
and U31030 (N_31030,N_27934,N_28566);
nand U31031 (N_31031,N_24164,N_28934);
xnor U31032 (N_31032,N_21956,N_28555);
nand U31033 (N_31033,N_25004,N_28779);
nor U31034 (N_31034,N_21459,N_22931);
xnor U31035 (N_31035,N_26055,N_24352);
or U31036 (N_31036,N_20753,N_28537);
nand U31037 (N_31037,N_29566,N_29370);
nand U31038 (N_31038,N_23263,N_28930);
xor U31039 (N_31039,N_27927,N_25923);
nor U31040 (N_31040,N_23173,N_29644);
nand U31041 (N_31041,N_27662,N_24114);
xnor U31042 (N_31042,N_24706,N_27179);
or U31043 (N_31043,N_27805,N_20175);
and U31044 (N_31044,N_20096,N_23247);
xor U31045 (N_31045,N_21782,N_20296);
and U31046 (N_31046,N_25909,N_24927);
or U31047 (N_31047,N_28993,N_21074);
and U31048 (N_31048,N_20990,N_20234);
and U31049 (N_31049,N_21433,N_23092);
nand U31050 (N_31050,N_28138,N_22890);
nand U31051 (N_31051,N_22194,N_27259);
nand U31052 (N_31052,N_29417,N_29745);
and U31053 (N_31053,N_20655,N_27387);
nor U31054 (N_31054,N_23548,N_24260);
nor U31055 (N_31055,N_21643,N_27004);
xnor U31056 (N_31056,N_26582,N_24558);
nand U31057 (N_31057,N_23300,N_27600);
nand U31058 (N_31058,N_29565,N_27656);
xor U31059 (N_31059,N_20415,N_29801);
nor U31060 (N_31060,N_28703,N_29429);
or U31061 (N_31061,N_20017,N_24295);
xor U31062 (N_31062,N_25580,N_26493);
and U31063 (N_31063,N_21904,N_29356);
and U31064 (N_31064,N_29173,N_23145);
nor U31065 (N_31065,N_27042,N_29800);
or U31066 (N_31066,N_20039,N_28634);
xor U31067 (N_31067,N_26804,N_21075);
and U31068 (N_31068,N_24106,N_29294);
nor U31069 (N_31069,N_24787,N_23917);
or U31070 (N_31070,N_25832,N_28195);
and U31071 (N_31071,N_28764,N_20309);
xor U31072 (N_31072,N_27450,N_24971);
nor U31073 (N_31073,N_21109,N_25557);
xnor U31074 (N_31074,N_29563,N_27141);
nor U31075 (N_31075,N_21453,N_29023);
or U31076 (N_31076,N_20268,N_25560);
and U31077 (N_31077,N_25705,N_22004);
nor U31078 (N_31078,N_25102,N_26373);
nor U31079 (N_31079,N_27342,N_25429);
nor U31080 (N_31080,N_22656,N_24551);
or U31081 (N_31081,N_24983,N_28780);
and U31082 (N_31082,N_28196,N_25494);
nor U31083 (N_31083,N_27231,N_20909);
nand U31084 (N_31084,N_23724,N_28720);
or U31085 (N_31085,N_20711,N_28540);
and U31086 (N_31086,N_21285,N_23107);
nor U31087 (N_31087,N_21405,N_21813);
nor U31088 (N_31088,N_29447,N_25440);
or U31089 (N_31089,N_27601,N_28074);
or U31090 (N_31090,N_24819,N_25995);
or U31091 (N_31091,N_24456,N_27181);
nand U31092 (N_31092,N_26106,N_21054);
xnor U31093 (N_31093,N_28592,N_21169);
xor U31094 (N_31094,N_23422,N_27696);
xor U31095 (N_31095,N_25354,N_24034);
xor U31096 (N_31096,N_27247,N_26363);
or U31097 (N_31097,N_25659,N_29558);
nand U31098 (N_31098,N_27530,N_24131);
and U31099 (N_31099,N_27558,N_21990);
nor U31100 (N_31100,N_27693,N_27785);
and U31101 (N_31101,N_27462,N_26156);
and U31102 (N_31102,N_26243,N_25229);
or U31103 (N_31103,N_28572,N_24383);
nor U31104 (N_31104,N_22084,N_22900);
nor U31105 (N_31105,N_21666,N_26792);
nand U31106 (N_31106,N_28363,N_25618);
xnor U31107 (N_31107,N_22014,N_23088);
xnor U31108 (N_31108,N_27697,N_24699);
or U31109 (N_31109,N_27642,N_22723);
nand U31110 (N_31110,N_22955,N_21362);
or U31111 (N_31111,N_24998,N_28498);
nor U31112 (N_31112,N_24987,N_29971);
nor U31113 (N_31113,N_27997,N_29956);
nand U31114 (N_31114,N_22788,N_22538);
and U31115 (N_31115,N_29651,N_25748);
and U31116 (N_31116,N_22179,N_24306);
and U31117 (N_31117,N_29853,N_24798);
nor U31118 (N_31118,N_29527,N_20266);
or U31119 (N_31119,N_27603,N_26818);
nor U31120 (N_31120,N_26178,N_22159);
or U31121 (N_31121,N_20561,N_28788);
xnor U31122 (N_31122,N_21090,N_24664);
nor U31123 (N_31123,N_22270,N_27318);
or U31124 (N_31124,N_20597,N_29374);
xnor U31125 (N_31125,N_28753,N_26705);
nor U31126 (N_31126,N_24540,N_22530);
xnor U31127 (N_31127,N_29855,N_29339);
or U31128 (N_31128,N_24651,N_23462);
nand U31129 (N_31129,N_21698,N_20287);
nor U31130 (N_31130,N_22345,N_20153);
or U31131 (N_31131,N_23209,N_26388);
xor U31132 (N_31132,N_24493,N_25250);
xnor U31133 (N_31133,N_22738,N_27197);
or U31134 (N_31134,N_21317,N_26229);
or U31135 (N_31135,N_25037,N_29660);
xor U31136 (N_31136,N_25729,N_29428);
or U31137 (N_31137,N_25075,N_26256);
and U31138 (N_31138,N_23750,N_24354);
xnor U31139 (N_31139,N_21071,N_21035);
and U31140 (N_31140,N_21479,N_21211);
or U31141 (N_31141,N_21697,N_23201);
or U31142 (N_31142,N_27159,N_23129);
and U31143 (N_31143,N_24229,N_29103);
or U31144 (N_31144,N_27060,N_26349);
or U31145 (N_31145,N_29426,N_24518);
nor U31146 (N_31146,N_24274,N_21482);
nor U31147 (N_31147,N_23500,N_26876);
xor U31148 (N_31148,N_21705,N_27079);
xor U31149 (N_31149,N_26477,N_20767);
xor U31150 (N_31150,N_21295,N_25726);
nor U31151 (N_31151,N_20661,N_23979);
xnor U31152 (N_31152,N_29184,N_28315);
nor U31153 (N_31153,N_25262,N_25717);
nand U31154 (N_31154,N_27974,N_27571);
or U31155 (N_31155,N_23192,N_22339);
or U31156 (N_31156,N_21438,N_22932);
nor U31157 (N_31157,N_28487,N_20554);
and U31158 (N_31158,N_25218,N_20660);
nor U31159 (N_31159,N_23592,N_27153);
nand U31160 (N_31160,N_24805,N_21431);
or U31161 (N_31161,N_25613,N_22698);
nand U31162 (N_31162,N_28255,N_21659);
nor U31163 (N_31163,N_23383,N_21017);
xor U31164 (N_31164,N_29689,N_24554);
and U31165 (N_31165,N_27570,N_20710);
nor U31166 (N_31166,N_20073,N_21147);
nor U31167 (N_31167,N_20329,N_20833);
or U31168 (N_31168,N_23610,N_23348);
and U31169 (N_31169,N_28339,N_23733);
xor U31170 (N_31170,N_28457,N_29167);
or U31171 (N_31171,N_24946,N_22849);
or U31172 (N_31172,N_22515,N_24735);
or U31173 (N_31173,N_20436,N_26900);
or U31174 (N_31174,N_23132,N_23012);
nor U31175 (N_31175,N_20291,N_28522);
xnor U31176 (N_31176,N_22468,N_27855);
nand U31177 (N_31177,N_28541,N_28181);
nor U31178 (N_31178,N_29032,N_24899);
nand U31179 (N_31179,N_26004,N_29664);
xnor U31180 (N_31180,N_29594,N_28647);
nand U31181 (N_31181,N_25565,N_20565);
nor U31182 (N_31182,N_28239,N_22487);
xnor U31183 (N_31183,N_29071,N_22132);
or U31184 (N_31184,N_27838,N_24340);
or U31185 (N_31185,N_26208,N_24997);
nor U31186 (N_31186,N_25340,N_29222);
nor U31187 (N_31187,N_27663,N_21216);
xnor U31188 (N_31188,N_23408,N_26351);
nor U31189 (N_31189,N_24912,N_24448);
xnor U31190 (N_31190,N_28849,N_21491);
or U31191 (N_31191,N_25088,N_20514);
or U31192 (N_31192,N_22217,N_20878);
xnor U31193 (N_31193,N_25176,N_24441);
xnor U31194 (N_31194,N_29673,N_26936);
and U31195 (N_31195,N_21064,N_28953);
nand U31196 (N_31196,N_25843,N_28619);
nand U31197 (N_31197,N_24641,N_28627);
xnor U31198 (N_31198,N_25474,N_24353);
xor U31199 (N_31199,N_24302,N_29541);
xor U31200 (N_31200,N_27847,N_22477);
nor U31201 (N_31201,N_26874,N_26820);
or U31202 (N_31202,N_29154,N_28642);
xnor U31203 (N_31203,N_26655,N_24763);
nor U31204 (N_31204,N_26879,N_27686);
nand U31205 (N_31205,N_26839,N_27296);
xnor U31206 (N_31206,N_29026,N_27649);
and U31207 (N_31207,N_27631,N_29625);
nor U31208 (N_31208,N_21656,N_28013);
xnor U31209 (N_31209,N_24761,N_29619);
xnor U31210 (N_31210,N_23722,N_22958);
xor U31211 (N_31211,N_23777,N_21323);
or U31212 (N_31212,N_21842,N_25387);
and U31213 (N_31213,N_28474,N_26475);
or U31214 (N_31214,N_21343,N_23801);
nor U31215 (N_31215,N_25241,N_26733);
or U31216 (N_31216,N_21368,N_22617);
nor U31217 (N_31217,N_27551,N_22579);
xnor U31218 (N_31218,N_28542,N_25945);
and U31219 (N_31219,N_26842,N_24351);
and U31220 (N_31220,N_29210,N_29966);
or U31221 (N_31221,N_20238,N_25786);
and U31222 (N_31222,N_23327,N_24122);
and U31223 (N_31223,N_25030,N_21830);
or U31224 (N_31224,N_21365,N_25956);
xor U31225 (N_31225,N_26718,N_24607);
nand U31226 (N_31226,N_28310,N_27874);
xnor U31227 (N_31227,N_26478,N_25733);
and U31228 (N_31228,N_23120,N_29750);
nand U31229 (N_31229,N_27072,N_21192);
xor U31230 (N_31230,N_29806,N_22903);
nor U31231 (N_31231,N_26246,N_23379);
or U31232 (N_31232,N_27790,N_23219);
and U31233 (N_31233,N_21958,N_26795);
and U31234 (N_31234,N_28341,N_22663);
or U31235 (N_31235,N_27910,N_24054);
nor U31236 (N_31236,N_21443,N_26017);
xor U31237 (N_31237,N_22739,N_24952);
xor U31238 (N_31238,N_24587,N_21715);
or U31239 (N_31239,N_28489,N_24962);
nand U31240 (N_31240,N_24239,N_27623);
and U31241 (N_31241,N_25443,N_26423);
xor U31242 (N_31242,N_25427,N_23526);
or U31243 (N_31243,N_27836,N_21575);
and U31244 (N_31244,N_27277,N_24240);
or U31245 (N_31245,N_24020,N_29753);
nand U31246 (N_31246,N_21321,N_21781);
xor U31247 (N_31247,N_20253,N_27442);
nor U31248 (N_31248,N_25731,N_23943);
nand U31249 (N_31249,N_29900,N_23016);
nand U31250 (N_31250,N_22986,N_26618);
nand U31251 (N_31251,N_25383,N_24085);
nand U31252 (N_31252,N_24109,N_23909);
or U31253 (N_31253,N_22222,N_23403);
nor U31254 (N_31254,N_27683,N_27236);
nor U31255 (N_31255,N_20827,N_27382);
nand U31256 (N_31256,N_27391,N_27470);
xor U31257 (N_31257,N_28300,N_22348);
nor U31258 (N_31258,N_22452,N_26207);
xor U31259 (N_31259,N_27768,N_22476);
xor U31260 (N_31260,N_29537,N_23045);
nand U31261 (N_31261,N_28046,N_21600);
nand U31262 (N_31262,N_21625,N_28444);
or U31263 (N_31263,N_23975,N_24269);
nor U31264 (N_31264,N_24221,N_24374);
xor U31265 (N_31265,N_25696,N_21048);
nand U31266 (N_31266,N_22128,N_29070);
xnor U31267 (N_31267,N_21931,N_21995);
or U31268 (N_31268,N_27645,N_24788);
and U31269 (N_31269,N_28096,N_21172);
or U31270 (N_31270,N_22662,N_27313);
nand U31271 (N_31271,N_21126,N_21175);
and U31272 (N_31272,N_26228,N_29831);
xor U31273 (N_31273,N_26695,N_23607);
nand U31274 (N_31274,N_26176,N_22039);
xor U31275 (N_31275,N_21150,N_24729);
xor U31276 (N_31276,N_22201,N_26096);
and U31277 (N_31277,N_28790,N_23929);
xor U31278 (N_31278,N_29016,N_22406);
xnor U31279 (N_31279,N_29012,N_20897);
nand U31280 (N_31280,N_25963,N_23357);
and U31281 (N_31281,N_24140,N_23883);
nand U31282 (N_31282,N_21073,N_29357);
xor U31283 (N_31283,N_24759,N_27868);
xor U31284 (N_31284,N_26487,N_24750);
nand U31285 (N_31285,N_20823,N_26770);
nor U31286 (N_31286,N_29984,N_29379);
and U31287 (N_31287,N_26836,N_22626);
nor U31288 (N_31288,N_27350,N_22379);
and U31289 (N_31289,N_24615,N_23240);
and U31290 (N_31290,N_29326,N_28719);
nand U31291 (N_31291,N_24447,N_25931);
nor U31292 (N_31292,N_29897,N_28231);
xnor U31293 (N_31293,N_25045,N_22309);
nor U31294 (N_31294,N_29785,N_26988);
nor U31295 (N_31295,N_29608,N_27957);
or U31296 (N_31296,N_25680,N_23449);
or U31297 (N_31297,N_27752,N_20441);
nand U31298 (N_31298,N_26504,N_29910);
xnor U31299 (N_31299,N_28249,N_25892);
nor U31300 (N_31300,N_25908,N_22675);
or U31301 (N_31301,N_26280,N_26600);
or U31302 (N_31302,N_21033,N_23014);
xnor U31303 (N_31303,N_22640,N_23884);
and U31304 (N_31304,N_25987,N_20849);
nand U31305 (N_31305,N_27939,N_25761);
nand U31306 (N_31306,N_22400,N_20046);
xor U31307 (N_31307,N_21483,N_24062);
or U31308 (N_31308,N_21818,N_25905);
nor U31309 (N_31309,N_20385,N_29445);
nand U31310 (N_31310,N_23395,N_26062);
and U31311 (N_31311,N_27492,N_22277);
nor U31312 (N_31312,N_27739,N_25074);
xor U31313 (N_31313,N_21744,N_27086);
or U31314 (N_31314,N_25009,N_27358);
xor U31315 (N_31315,N_21191,N_21208);
or U31316 (N_31316,N_22767,N_27216);
or U31317 (N_31317,N_26182,N_20023);
nor U31318 (N_31318,N_29279,N_20690);
and U31319 (N_31319,N_22035,N_27142);
xor U31320 (N_31320,N_25619,N_21655);
and U31321 (N_31321,N_26603,N_25309);
and U31322 (N_31322,N_23121,N_27689);
nand U31323 (N_31323,N_21686,N_21502);
or U31324 (N_31324,N_27128,N_20498);
or U31325 (N_31325,N_28565,N_23391);
or U31326 (N_31326,N_25472,N_21996);
nand U31327 (N_31327,N_24916,N_23971);
or U31328 (N_31328,N_26814,N_22699);
and U31329 (N_31329,N_24084,N_28387);
or U31330 (N_31330,N_27945,N_26680);
nand U31331 (N_31331,N_29638,N_20145);
xnor U31332 (N_31332,N_27191,N_22614);
nor U31333 (N_31333,N_20180,N_28808);
or U31334 (N_31334,N_23653,N_22833);
or U31335 (N_31335,N_20512,N_26432);
and U31336 (N_31336,N_29586,N_24188);
and U31337 (N_31337,N_23603,N_28122);
and U31338 (N_31338,N_21310,N_23781);
and U31339 (N_31339,N_27629,N_20130);
nand U31340 (N_31340,N_22711,N_22769);
nand U31341 (N_31341,N_25492,N_28478);
nand U31342 (N_31342,N_23258,N_29040);
or U31343 (N_31343,N_22621,N_24535);
xnor U31344 (N_31344,N_22426,N_27107);
and U31345 (N_31345,N_29724,N_20279);
or U31346 (N_31346,N_20043,N_23682);
and U31347 (N_31347,N_29240,N_28556);
and U31348 (N_31348,N_23418,N_20317);
xnor U31349 (N_31349,N_21227,N_23436);
and U31350 (N_31350,N_24458,N_28638);
and U31351 (N_31351,N_29349,N_27138);
nand U31352 (N_31352,N_23962,N_21301);
and U31353 (N_31353,N_25800,N_29468);
or U31354 (N_31354,N_26420,N_24404);
xnor U31355 (N_31355,N_21313,N_20985);
xnor U31356 (N_31356,N_23851,N_26608);
xnor U31357 (N_31357,N_28926,N_23239);
and U31358 (N_31358,N_23275,N_27368);
and U31359 (N_31359,N_27303,N_20949);
or U31360 (N_31360,N_24591,N_20188);
or U31361 (N_31361,N_20098,N_27050);
xnor U31362 (N_31362,N_26683,N_25662);
or U31363 (N_31363,N_27127,N_22832);
xnor U31364 (N_31364,N_25266,N_25163);
nor U31365 (N_31365,N_25606,N_25978);
or U31366 (N_31366,N_20634,N_23556);
nor U31367 (N_31367,N_26764,N_24786);
and U31368 (N_31368,N_22852,N_22008);
nor U31369 (N_31369,N_20148,N_20997);
or U31370 (N_31370,N_27186,N_27292);
or U31371 (N_31371,N_22691,N_28960);
nor U31372 (N_31372,N_26355,N_25459);
and U31373 (N_31373,N_24434,N_24045);
or U31374 (N_31374,N_22804,N_25774);
xor U31375 (N_31375,N_25182,N_29529);
nand U31376 (N_31376,N_29723,N_28006);
nor U31377 (N_31377,N_25856,N_27234);
xor U31378 (N_31378,N_20797,N_25842);
nand U31379 (N_31379,N_24313,N_24412);
and U31380 (N_31380,N_29045,N_23229);
or U31381 (N_31381,N_27875,N_21326);
nand U31382 (N_31382,N_24154,N_24742);
nand U31383 (N_31383,N_29942,N_29058);
nand U31384 (N_31384,N_21566,N_22693);
or U31385 (N_31385,N_29677,N_21615);
xnor U31386 (N_31386,N_21403,N_24539);
or U31387 (N_31387,N_20293,N_22647);
nand U31388 (N_31388,N_20094,N_24579);
and U31389 (N_31389,N_21084,N_29702);
xor U31390 (N_31390,N_28443,N_28252);
or U31391 (N_31391,N_20792,N_28389);
and U31392 (N_31392,N_29516,N_26867);
nor U31393 (N_31393,N_21128,N_23426);
nand U31394 (N_31394,N_26866,N_27701);
and U31395 (N_31395,N_21423,N_28481);
xor U31396 (N_31396,N_21315,N_20495);
and U31397 (N_31397,N_20216,N_24698);
and U31398 (N_31398,N_28103,N_28708);
nor U31399 (N_31399,N_26321,N_21070);
and U31400 (N_31400,N_28281,N_27526);
or U31401 (N_31401,N_23509,N_21262);
xor U31402 (N_31402,N_21568,N_25992);
xnor U31403 (N_31403,N_27220,N_22940);
nand U31404 (N_31404,N_27022,N_25194);
or U31405 (N_31405,N_21850,N_25724);
nor U31406 (N_31406,N_20413,N_25423);
or U31407 (N_31407,N_24015,N_21548);
nand U31408 (N_31408,N_28773,N_23800);
nand U31409 (N_31409,N_24545,N_21545);
nand U31410 (N_31410,N_27929,N_25901);
nor U31411 (N_31411,N_23679,N_28136);
or U31412 (N_31412,N_28125,N_22187);
nor U31413 (N_31413,N_21939,N_27839);
or U31414 (N_31414,N_25390,N_20742);
xor U31415 (N_31415,N_28626,N_26407);
or U31416 (N_31416,N_25871,N_26552);
xor U31417 (N_31417,N_26584,N_20859);
or U31418 (N_31418,N_24135,N_24733);
xnor U31419 (N_31419,N_23789,N_22173);
and U31420 (N_31420,N_29431,N_20491);
nor U31421 (N_31421,N_21963,N_24754);
nor U31422 (N_31422,N_21138,N_28303);
and U31423 (N_31423,N_24760,N_21519);
nand U31424 (N_31424,N_20993,N_21861);
xor U31425 (N_31425,N_26871,N_24649);
or U31426 (N_31426,N_25922,N_21711);
nand U31427 (N_31427,N_21967,N_25195);
xnor U31428 (N_31428,N_27052,N_22518);
nor U31429 (N_31429,N_21352,N_20751);
and U31430 (N_31430,N_20481,N_23997);
and U31431 (N_31431,N_21324,N_21839);
and U31432 (N_31432,N_24005,N_20237);
xor U31433 (N_31433,N_24681,N_23017);
or U31434 (N_31434,N_25607,N_27627);
and U31435 (N_31435,N_22676,N_28514);
nor U31436 (N_31436,N_29170,N_24999);
xnor U31437 (N_31437,N_21026,N_20830);
nor U31438 (N_31438,N_27608,N_28661);
nand U31439 (N_31439,N_23186,N_22430);
nor U31440 (N_31440,N_23039,N_25019);
and U31441 (N_31441,N_20893,N_20358);
and U31442 (N_31442,N_21848,N_22152);
xor U31443 (N_31443,N_27455,N_22193);
xor U31444 (N_31444,N_20270,N_25317);
xnor U31445 (N_31445,N_25793,N_25829);
xnor U31446 (N_31446,N_23731,N_29433);
nand U31447 (N_31447,N_25286,N_20092);
nand U31448 (N_31448,N_24337,N_28261);
xnor U31449 (N_31449,N_21290,N_22684);
xor U31450 (N_31450,N_27253,N_20645);
nand U31451 (N_31451,N_28803,N_25000);
nand U31452 (N_31452,N_28177,N_25869);
nand U31453 (N_31453,N_24653,N_26746);
and U31454 (N_31454,N_20732,N_24216);
nor U31455 (N_31455,N_25189,N_28298);
and U31456 (N_31456,N_23136,N_26703);
and U31457 (N_31457,N_23468,N_26925);
nor U31458 (N_31458,N_25672,N_22389);
and U31459 (N_31459,N_28913,N_26135);
nand U31460 (N_31460,N_22219,N_23776);
or U31461 (N_31461,N_27533,N_29304);
xnor U31462 (N_31462,N_23291,N_26371);
nor U31463 (N_31463,N_23511,N_29868);
and U31464 (N_31464,N_22930,N_20793);
or U31465 (N_31465,N_23148,N_28805);
nand U31466 (N_31466,N_25757,N_26404);
or U31467 (N_31467,N_21274,N_25764);
nor U31468 (N_31468,N_20689,N_26534);
and U31469 (N_31469,N_20312,N_24937);
nor U31470 (N_31470,N_29764,N_21422);
nor U31471 (N_31471,N_20526,N_20585);
xnor U31472 (N_31472,N_29802,N_26800);
and U31473 (N_31473,N_29717,N_26375);
nor U31474 (N_31474,N_24487,N_25039);
xor U31475 (N_31475,N_26672,N_24633);
nor U31476 (N_31476,N_20368,N_27210);
nor U31477 (N_31477,N_26219,N_27985);
xor U31478 (N_31478,N_22729,N_23210);
nor U31479 (N_31479,N_24643,N_22214);
nand U31480 (N_31480,N_26641,N_27923);
and U31481 (N_31481,N_29450,N_24776);
nor U31482 (N_31482,N_24098,N_26725);
or U31483 (N_31483,N_29886,N_28648);
or U31484 (N_31484,N_24366,N_29599);
or U31485 (N_31485,N_27355,N_24344);
and U31486 (N_31486,N_23651,N_20713);
or U31487 (N_31487,N_25302,N_22799);
or U31488 (N_31488,N_22065,N_27208);
and U31489 (N_31489,N_27084,N_20649);
xor U31490 (N_31490,N_22394,N_27376);
xor U31491 (N_31491,N_24564,N_23830);
xor U31492 (N_31492,N_22052,N_28169);
nand U31493 (N_31493,N_25601,N_27733);
nor U31494 (N_31494,N_24524,N_29146);
xnor U31495 (N_31495,N_25938,N_24602);
nor U31496 (N_31496,N_22233,N_29117);
xnor U31497 (N_31497,N_25665,N_25990);
nor U31498 (N_31498,N_25047,N_25236);
and U31499 (N_31499,N_28234,N_26320);
nand U31500 (N_31500,N_22998,N_20010);
nor U31501 (N_31501,N_23699,N_26291);
and U31502 (N_31502,N_27061,N_26436);
xnor U31503 (N_31503,N_22763,N_28156);
or U31504 (N_31504,N_20056,N_20817);
xor U31505 (N_31505,N_21933,N_22889);
and U31506 (N_31506,N_27412,N_29136);
and U31507 (N_31507,N_20507,N_20594);
nand U31508 (N_31508,N_23514,N_26858);
xnor U31509 (N_31509,N_28509,N_28328);
nand U31510 (N_31510,N_28584,N_21112);
or U31511 (N_31511,N_27431,N_20541);
nand U31512 (N_31512,N_22732,N_21726);
nand U31513 (N_31513,N_26253,N_21563);
nor U31514 (N_31514,N_20408,N_25513);
xor U31515 (N_31515,N_22909,N_22826);
and U31516 (N_31516,N_25210,N_26162);
or U31517 (N_31517,N_22427,N_25071);
xor U31518 (N_31518,N_25425,N_26710);
or U31519 (N_31519,N_26312,N_23692);
and U31520 (N_31520,N_23225,N_21617);
or U31521 (N_31521,N_21481,N_20533);
or U31522 (N_31522,N_24182,N_23072);
or U31523 (N_31523,N_24268,N_21221);
xor U31524 (N_31524,N_25907,N_26130);
xnor U31525 (N_31525,N_20136,N_27560);
nand U31526 (N_31526,N_26536,N_26681);
xor U31527 (N_31527,N_26734,N_23675);
or U31528 (N_31528,N_21244,N_24205);
nand U31529 (N_31529,N_27035,N_27089);
nor U31530 (N_31530,N_28270,N_22242);
or U31531 (N_31531,N_20086,N_26288);
nand U31532 (N_31532,N_21590,N_26408);
nand U31533 (N_31533,N_23370,N_20347);
nand U31534 (N_31534,N_23870,N_25175);
or U31535 (N_31535,N_26168,N_26147);
nor U31536 (N_31536,N_26981,N_29232);
nand U31537 (N_31537,N_28585,N_22331);
or U31538 (N_31538,N_27545,N_22979);
xnor U31539 (N_31539,N_26001,N_24381);
and U31540 (N_31540,N_27444,N_21877);
xor U31541 (N_31541,N_28411,N_27156);
nor U31542 (N_31542,N_26072,N_21442);
nor U31543 (N_31543,N_25126,N_27182);
nor U31544 (N_31544,N_29323,N_23560);
nor U31545 (N_31545,N_24642,N_21263);
and U31546 (N_31546,N_20528,N_28347);
xnor U31547 (N_31547,N_28967,N_22726);
xor U31548 (N_31548,N_23218,N_21806);
or U31549 (N_31549,N_29827,N_25310);
nor U31550 (N_31550,N_22638,N_20460);
nor U31551 (N_31551,N_29256,N_20947);
and U31552 (N_31552,N_20390,N_27932);
nand U31553 (N_31553,N_23974,N_20209);
and U31554 (N_31554,N_23152,N_20928);
nand U31555 (N_31555,N_20310,N_23287);
and U31556 (N_31556,N_20851,N_21797);
xnor U31557 (N_31557,N_21891,N_20675);
nor U31558 (N_31558,N_24846,N_25094);
nand U31559 (N_31559,N_21462,N_22694);
and U31560 (N_31560,N_23887,N_25830);
xnor U31561 (N_31561,N_29000,N_21630);
nand U31562 (N_31562,N_20687,N_27829);
or U31563 (N_31563,N_23706,N_21943);
xor U31564 (N_31564,N_29824,N_21055);
nand U31565 (N_31565,N_25455,N_23488);
nand U31566 (N_31566,N_27469,N_27023);
xnor U31567 (N_31567,N_28759,N_24245);
nand U31568 (N_31568,N_23085,N_21534);
nor U31569 (N_31569,N_20122,N_20748);
and U31570 (N_31570,N_28952,N_25602);
and U31571 (N_31571,N_24479,N_25116);
nand U31572 (N_31572,N_26213,N_25053);
nor U31573 (N_31573,N_29754,N_25944);
and U31574 (N_31574,N_20538,N_24508);
xor U31575 (N_31575,N_29628,N_21439);
and U31576 (N_31576,N_21269,N_20532);
and U31577 (N_31577,N_28892,N_24347);
nor U31578 (N_31578,N_29368,N_21792);
nor U31579 (N_31579,N_20693,N_20141);
xor U31580 (N_31580,N_21013,N_27528);
nand U31581 (N_31581,N_26577,N_24686);
nand U31582 (N_31582,N_21978,N_20374);
xor U31583 (N_31583,N_25655,N_29882);
xnor U31584 (N_31584,N_26939,N_28912);
and U31585 (N_31585,N_21417,N_23027);
nor U31586 (N_31586,N_22811,N_26445);
or U31587 (N_31587,N_27386,N_29783);
or U31588 (N_31588,N_23298,N_20920);
xnor U31589 (N_31589,N_25341,N_25291);
or U31590 (N_31590,N_29317,N_24373);
nand U31591 (N_31591,N_29483,N_29457);
and U31592 (N_31592,N_23100,N_27520);
nor U31593 (N_31593,N_26068,N_25115);
xor U31594 (N_31594,N_28047,N_29098);
and U31595 (N_31595,N_23916,N_24089);
and U31596 (N_31596,N_25975,N_21703);
xor U31597 (N_31597,N_27610,N_29301);
or U31598 (N_31598,N_27122,N_20123);
nand U31599 (N_31599,N_25685,N_23046);
nand U31600 (N_31600,N_22360,N_27333);
nor U31601 (N_31601,N_23430,N_25496);
and U31602 (N_31602,N_25093,N_28734);
nor U31603 (N_31603,N_22791,N_25072);
or U31604 (N_31604,N_26131,N_24665);
and U31605 (N_31605,N_26545,N_29941);
nand U31606 (N_31606,N_20051,N_27613);
xnor U31607 (N_31607,N_26730,N_27315);
or U31608 (N_31608,N_28435,N_26383);
nand U31609 (N_31609,N_28079,N_23322);
or U31610 (N_31610,N_27479,N_22746);
and U31611 (N_31611,N_20449,N_20749);
nor U31612 (N_31612,N_25099,N_20370);
nand U31613 (N_31613,N_25884,N_26134);
and U31614 (N_31614,N_23669,N_25520);
or U31615 (N_31615,N_23435,N_20556);
and U31616 (N_31616,N_25541,N_22246);
nand U31617 (N_31617,N_29591,N_27049);
xnor U31618 (N_31618,N_23165,N_20708);
nor U31619 (N_31619,N_22013,N_25997);
and U31620 (N_31620,N_26109,N_20777);
and U31621 (N_31621,N_28903,N_20812);
nand U31622 (N_31622,N_28998,N_25068);
nor U31623 (N_31623,N_29495,N_28098);
or U31624 (N_31624,N_28841,N_27584);
xor U31625 (N_31625,N_22292,N_27955);
nand U31626 (N_31626,N_27515,N_21879);
xnor U31627 (N_31627,N_25162,N_21199);
and U31628 (N_31628,N_20334,N_28368);
and U31629 (N_31629,N_23824,N_20416);
and U31630 (N_31630,N_25272,N_26987);
nor U31631 (N_31631,N_22162,N_20213);
xnor U31632 (N_31632,N_22750,N_26480);
and U31633 (N_31633,N_23359,N_26305);
and U31634 (N_31634,N_29290,N_24947);
nand U31635 (N_31635,N_29987,N_25823);
nand U31636 (N_31636,N_26589,N_25841);
xor U31637 (N_31637,N_29335,N_29577);
nand U31638 (N_31638,N_20045,N_25020);
or U31639 (N_31639,N_22771,N_26384);
and U31640 (N_31640,N_28745,N_24208);
nor U31641 (N_31641,N_24477,N_28706);
nor U31642 (N_31642,N_27190,N_25529);
xnor U31643 (N_31643,N_29895,N_26016);
nand U31644 (N_31644,N_21760,N_25033);
nor U31645 (N_31645,N_20276,N_21230);
nor U31646 (N_31646,N_22245,N_29219);
or U31647 (N_31647,N_26314,N_28684);
nand U31648 (N_31648,N_23873,N_22262);
and U31649 (N_31649,N_23112,N_27857);
nor U31650 (N_31650,N_29160,N_26434);
or U31651 (N_31651,N_21750,N_29720);
nor U31652 (N_31652,N_22112,N_29666);
xor U31653 (N_31653,N_28218,N_20244);
and U31654 (N_31654,N_25049,N_26169);
nand U31655 (N_31655,N_25765,N_26266);
nand U31656 (N_31656,N_20324,N_29056);
or U31657 (N_31657,N_29653,N_29196);
xor U31658 (N_31658,N_25395,N_25521);
nand U31659 (N_31659,N_24298,N_21476);
nand U31660 (N_31660,N_22654,N_23998);
xnor U31661 (N_31661,N_20113,N_23957);
xnor U31662 (N_31662,N_23739,N_23749);
xnor U31663 (N_31663,N_28631,N_23273);
nand U31664 (N_31664,N_29881,N_25292);
nor U31665 (N_31665,N_20733,N_26295);
xor U31666 (N_31666,N_26107,N_26862);
nor U31667 (N_31667,N_29488,N_24049);
nand U31668 (N_31668,N_20165,N_23169);
or U31669 (N_31669,N_23494,N_25891);
xnor U31670 (N_31670,N_24667,N_22225);
nor U31671 (N_31671,N_25105,N_29712);
xnor U31672 (N_31672,N_24191,N_26699);
nor U31673 (N_31673,N_22081,N_27796);
and U31674 (N_31674,N_20062,N_23761);
nand U31675 (N_31675,N_22649,N_26973);
and U31676 (N_31676,N_22881,N_21258);
nor U31677 (N_31677,N_26234,N_25337);
nor U31678 (N_31678,N_22032,N_24167);
nor U31679 (N_31679,N_27844,N_28543);
xnor U31680 (N_31680,N_20120,N_26163);
and U31681 (N_31681,N_21085,N_22706);
or U31682 (N_31682,N_20338,N_22894);
xnor U31683 (N_31683,N_23717,N_22090);
nand U31684 (N_31684,N_28700,N_28899);
xor U31685 (N_31685,N_27085,N_28564);
xnor U31686 (N_31686,N_24323,N_26330);
nand U31687 (N_31687,N_27691,N_28269);
nor U31688 (N_31688,N_23491,N_22564);
xor U31689 (N_31689,N_20179,N_21843);
xor U31690 (N_31690,N_28367,N_21985);
and U31691 (N_31691,N_29678,N_26010);
nor U31692 (N_31692,N_29042,N_22924);
or U31693 (N_31693,N_27763,N_22027);
xnor U31694 (N_31694,N_26961,N_23004);
nand U31695 (N_31695,N_26916,N_24047);
nand U31696 (N_31696,N_27306,N_27105);
and U31697 (N_31697,N_20723,N_25870);
nor U31698 (N_31698,N_23834,N_27435);
nor U31699 (N_31699,N_25349,N_23859);
or U31700 (N_31700,N_28679,N_24905);
nand U31701 (N_31701,N_29097,N_20825);
or U31702 (N_31702,N_27329,N_29380);
and U31703 (N_31703,N_24940,N_25903);
xnor U31704 (N_31704,N_28424,N_28578);
xor U31705 (N_31705,N_22556,N_23557);
xnor U31706 (N_31706,N_27349,N_26272);
or U31707 (N_31707,N_29676,N_22741);
nand U31708 (N_31708,N_23087,N_22622);
and U31709 (N_31709,N_21347,N_27682);
nand U31710 (N_31710,N_22988,N_24746);
nand U31711 (N_31711,N_23098,N_26086);
or U31712 (N_31712,N_22234,N_20705);
xnor U31713 (N_31713,N_27737,N_22497);
nand U31714 (N_31714,N_28306,N_24561);
nand U31715 (N_31715,N_21179,N_26088);
or U31716 (N_31716,N_25197,N_29047);
xor U31717 (N_31717,N_27201,N_22572);
xor U31718 (N_31718,N_22485,N_25692);
or U31719 (N_31719,N_20935,N_22876);
nor U31720 (N_31720,N_28445,N_22133);
xor U31721 (N_31721,N_22596,N_22850);
nor U31722 (N_31722,N_26789,N_26895);
and U31723 (N_31723,N_28650,N_25177);
xnor U31724 (N_31724,N_28266,N_23288);
nor U31725 (N_31725,N_29756,N_25015);
and U31726 (N_31726,N_25740,N_21518);
nor U31727 (N_31727,N_20079,N_26738);
and U31728 (N_31728,N_21201,N_25570);
nand U31729 (N_31729,N_28065,N_25325);
nand U31730 (N_31730,N_26533,N_22709);
nor U31731 (N_31731,N_29947,N_23179);
or U31732 (N_31732,N_20717,N_25866);
xor U31733 (N_31733,N_29821,N_26776);
and U31734 (N_31734,N_21771,N_27895);
nor U31735 (N_31735,N_23342,N_28662);
and U31736 (N_31736,N_26154,N_22573);
nor U31737 (N_31737,N_26690,N_22990);
xor U31738 (N_31738,N_25708,N_26774);
and U31739 (N_31739,N_28446,N_29760);
xor U31740 (N_31740,N_21197,N_29534);
xnor U31741 (N_31741,N_29013,N_24797);
or U31742 (N_31742,N_29503,N_21161);
nand U31743 (N_31743,N_21163,N_22974);
nand U31744 (N_31744,N_26883,N_27810);
and U31745 (N_31745,N_26578,N_20396);
and U31746 (N_31746,N_20177,N_20589);
or U31747 (N_31747,N_21844,N_27980);
xnor U31748 (N_31748,N_20169,N_26469);
nor U31749 (N_31749,N_22037,N_29514);
xnor U31750 (N_31750,N_26212,N_22205);
nor U31751 (N_31751,N_29337,N_27967);
or U31752 (N_31752,N_22066,N_29662);
nor U31753 (N_31753,N_27499,N_23208);
xor U31754 (N_31754,N_28229,N_22163);
and U31755 (N_31755,N_28503,N_24281);
or U31756 (N_31756,N_25787,N_20782);
and U31757 (N_31757,N_20355,N_24553);
xnor U31758 (N_31758,N_27071,N_20233);
nand U31759 (N_31759,N_23516,N_22535);
and U31760 (N_31760,N_26543,N_29864);
and U31761 (N_31761,N_21402,N_25553);
and U31762 (N_31762,N_26022,N_28267);
nor U31763 (N_31763,N_25371,N_21477);
xnor U31764 (N_31764,N_23773,N_23429);
nor U31765 (N_31765,N_20626,N_27746);
and U31766 (N_31766,N_23815,N_24758);
nor U31767 (N_31767,N_21341,N_22968);
nor U31768 (N_31768,N_20000,N_29120);
xnor U31769 (N_31769,N_26812,N_29208);
and U31770 (N_31770,N_20478,N_27920);
nor U31771 (N_31771,N_22701,N_27461);
nand U31772 (N_31772,N_21578,N_27687);
xnor U31773 (N_31773,N_20461,N_28451);
xnor U31774 (N_31774,N_24734,N_22681);
xnor U31775 (N_31775,N_28382,N_29950);
and U31776 (N_31776,N_28938,N_29093);
or U31777 (N_31777,N_20110,N_20559);
nand U31778 (N_31778,N_26037,N_24151);
or U31779 (N_31779,N_20858,N_24248);
nand U31780 (N_31780,N_28675,N_20946);
nand U31781 (N_31781,N_29143,N_20644);
or U31782 (N_31782,N_24165,N_28263);
nand U31783 (N_31783,N_27724,N_27595);
and U31784 (N_31784,N_29549,N_27373);
nor U31785 (N_31785,N_27952,N_22869);
and U31786 (N_31786,N_20819,N_22831);
and U31787 (N_31787,N_27808,N_24094);
xnor U31788 (N_31788,N_24519,N_24782);
xnor U31789 (N_31789,N_28327,N_23520);
nand U31790 (N_31790,N_22387,N_21009);
and U31791 (N_31791,N_25636,N_24339);
and U31792 (N_31792,N_29221,N_22074);
nand U31793 (N_31793,N_20838,N_28061);
nand U31794 (N_31794,N_22466,N_28826);
nand U31795 (N_31795,N_21786,N_25649);
and U31796 (N_31796,N_24869,N_21743);
nor U31797 (N_31797,N_28447,N_28395);
or U31798 (N_31798,N_26366,N_26514);
and U31799 (N_31799,N_28908,N_29929);
nand U31800 (N_31800,N_24810,N_29346);
or U31801 (N_31801,N_29073,N_28257);
and U31802 (N_31802,N_22661,N_24755);
xor U31803 (N_31803,N_20420,N_29178);
nand U31804 (N_31804,N_20242,N_23791);
and U31805 (N_31805,N_28485,N_27418);
and U31806 (N_31806,N_20210,N_20525);
nor U31807 (N_31807,N_22446,N_27660);
nand U31808 (N_31808,N_24779,N_24086);
or U31809 (N_31809,N_28028,N_28696);
and U31810 (N_31810,N_27908,N_23281);
xnor U31811 (N_31811,N_24172,N_21104);
nand U31812 (N_31812,N_26303,N_26541);
xor U31813 (N_31813,N_25600,N_27881);
nor U31814 (N_31814,N_24744,N_28630);
nor U31815 (N_31815,N_21565,N_20898);
nor U31816 (N_31816,N_27784,N_22753);
nor U31817 (N_31817,N_28259,N_27765);
xnor U31818 (N_31818,N_22581,N_24255);
or U31819 (N_31819,N_21668,N_27894);
nor U31820 (N_31820,N_29939,N_25852);
and U31821 (N_31821,N_27016,N_24143);
nand U31822 (N_31822,N_29612,N_21700);
nor U31823 (N_31823,N_22420,N_23605);
nor U31824 (N_31824,N_24666,N_24630);
nor U31825 (N_31825,N_27215,N_24071);
xnor U31826 (N_31826,N_26027,N_26051);
nand U31827 (N_31827,N_22145,N_20054);
and U31828 (N_31828,N_26100,N_28361);
or U31829 (N_31829,N_25512,N_20383);
xor U31830 (N_31830,N_21930,N_23498);
and U31831 (N_31831,N_26819,N_21831);
nor U31832 (N_31832,N_23187,N_21386);
nand U31833 (N_31833,N_20977,N_28761);
nand U31834 (N_31834,N_26845,N_25453);
nor U31835 (N_31835,N_26063,N_25196);
nand U31836 (N_31836,N_28353,N_24149);
or U31837 (N_31837,N_29553,N_23074);
xor U31838 (N_31838,N_21723,N_27151);
and U31839 (N_31839,N_28073,N_29588);
or U31840 (N_31840,N_27787,N_25556);
xor U31841 (N_31841,N_21053,N_21374);
xor U31842 (N_31842,N_23553,N_25498);
or U31843 (N_31843,N_25044,N_25778);
and U31844 (N_31844,N_27574,N_22299);
nor U31845 (N_31845,N_25736,N_23681);
xnor U31846 (N_31846,N_28876,N_22248);
nand U31847 (N_31847,N_25752,N_26251);
and U31848 (N_31848,N_29589,N_23311);
and U31849 (N_31849,N_26270,N_23885);
xnor U31850 (N_31850,N_22506,N_21833);
nor U31851 (N_31851,N_22385,N_23741);
and U31852 (N_31852,N_21576,N_22202);
nor U31853 (N_31853,N_26012,N_25771);
nor U31854 (N_31854,N_28284,N_24835);
or U31855 (N_31855,N_23188,N_21267);
or U31856 (N_31856,N_29075,N_21050);
nand U31857 (N_31857,N_23542,N_20677);
nand U31858 (N_31858,N_27175,N_22665);
xnor U31859 (N_31859,N_21426,N_29332);
or U31860 (N_31860,N_24559,N_21993);
nand U31861 (N_31861,N_22368,N_27648);
and U31862 (N_31862,N_23638,N_27098);
xor U31863 (N_31863,N_21713,N_21735);
nand U31864 (N_31864,N_21427,N_29298);
and U31865 (N_31865,N_25688,N_28601);
and U31866 (N_31866,N_24301,N_21896);
or U31867 (N_31867,N_23460,N_27636);
nor U31868 (N_31868,N_29325,N_21855);
nor U31869 (N_31869,N_20208,N_22505);
nand U31870 (N_31870,N_21866,N_28419);
and U31871 (N_31871,N_21739,N_21970);
nor U31872 (N_31872,N_25215,N_27547);
or U31873 (N_31873,N_29648,N_27020);
and U31874 (N_31874,N_24964,N_21099);
nand U31875 (N_31875,N_22069,N_23213);
xnor U31876 (N_31876,N_21541,N_23628);
xnor U31877 (N_31877,N_29629,N_29312);
xor U31878 (N_31878,N_28064,N_27935);
nor U31879 (N_31879,N_23589,N_25415);
xor U31880 (N_31880,N_27192,N_24033);
or U31881 (N_31881,N_20521,N_27777);
and U31882 (N_31882,N_20203,N_29791);
or U31883 (N_31883,N_20302,N_20930);
or U31884 (N_31884,N_20226,N_24850);
or U31885 (N_31885,N_23025,N_27513);
nor U31886 (N_31886,N_29849,N_21348);
xnor U31887 (N_31887,N_23021,N_23361);
and U31888 (N_31888,N_24259,N_20580);
and U31889 (N_31889,N_26214,N_23131);
and U31890 (N_31890,N_25885,N_29811);
or U31891 (N_31891,N_24822,N_20752);
nor U31892 (N_31892,N_25398,N_26000);
or U31893 (N_31893,N_28230,N_21820);
nand U31894 (N_31894,N_23267,N_27572);
or U31895 (N_31895,N_26211,N_25861);
or U31896 (N_31896,N_25878,N_28437);
or U31897 (N_31897,N_29162,N_23420);
nand U31898 (N_31898,N_21376,N_25930);
nand U31899 (N_31899,N_23473,N_24858);
or U31900 (N_31900,N_24110,N_20880);
nand U31901 (N_31901,N_22028,N_23413);
or U31902 (N_31902,N_21828,N_24659);
and U31903 (N_31903,N_29706,N_28345);
nor U31904 (N_31904,N_24431,N_20534);
or U31905 (N_31905,N_28413,N_29790);
nor U31906 (N_31906,N_29615,N_22938);
nand U31907 (N_31907,N_20160,N_26890);
nor U31908 (N_31908,N_21710,N_29999);
or U31909 (N_31909,N_22631,N_25713);
or U31910 (N_31910,N_27820,N_23123);
nor U31911 (N_31911,N_24108,N_25442);
xor U31912 (N_31912,N_28583,N_29757);
and U31913 (N_31913,N_26520,N_21719);
nand U31914 (N_31914,N_20201,N_23365);
nand U31915 (N_31915,N_26602,N_25714);
or U31916 (N_31916,N_29768,N_20116);
and U31917 (N_31917,N_23503,N_28024);
xor U31918 (N_31918,N_24537,N_27615);
and U31919 (N_31919,N_23060,N_27877);
or U31920 (N_31920,N_23987,N_24613);
and U31921 (N_31921,N_25889,N_28768);
and U31922 (N_31922,N_27899,N_21612);
and U31923 (N_31923,N_23855,N_28288);
nand U31924 (N_31924,N_25046,N_21914);
nand U31925 (N_31925,N_29923,N_25213);
nand U31926 (N_31926,N_24834,N_22412);
and U31927 (N_31927,N_20800,N_23183);
or U31928 (N_31928,N_28032,N_25755);
or U31929 (N_31929,N_20154,N_28801);
and U31930 (N_31930,N_27155,N_24187);
nor U31931 (N_31931,N_20725,N_29696);
nor U31932 (N_31932,N_28915,N_26302);
or U31933 (N_31933,N_25129,N_20505);
nand U31934 (N_31934,N_27396,N_20212);
and U31935 (N_31935,N_29579,N_26463);
and U31936 (N_31936,N_22021,N_23912);
or U31937 (N_31937,N_25890,N_20610);
nor U31938 (N_31938,N_28448,N_27147);
and U31939 (N_31939,N_26278,N_24833);
nand U31940 (N_31940,N_28793,N_28279);
or U31941 (N_31941,N_24061,N_29952);
xnor U31942 (N_31942,N_21745,N_25475);
xor U31943 (N_31943,N_26737,N_21119);
xnor U31944 (N_31944,N_22933,N_28493);
or U31945 (N_31945,N_23865,N_28116);
and U31946 (N_31946,N_25767,N_23451);
or U31947 (N_31947,N_20450,N_27657);
or U31948 (N_31948,N_23639,N_24770);
nand U31949 (N_31949,N_20961,N_25912);
and U31950 (N_31950,N_29621,N_23086);
and U31951 (N_31951,N_29116,N_24963);
xor U31952 (N_31952,N_28985,N_29155);
and U31953 (N_31953,N_20133,N_29187);
or U31954 (N_31954,N_21738,N_28282);
xnor U31955 (N_31955,N_20729,N_26367);
xor U31956 (N_31956,N_29157,N_28900);
and U31957 (N_31957,N_23241,N_20575);
and U31958 (N_31958,N_29600,N_25445);
nand U31959 (N_31959,N_20504,N_24507);
or U31960 (N_31960,N_26708,N_28344);
nand U31961 (N_31961,N_29818,N_23249);
or U31962 (N_31962,N_26449,N_25237);
and U31963 (N_31963,N_28014,N_20769);
and U31964 (N_31964,N_25370,N_24236);
nor U31965 (N_31965,N_29573,N_21581);
or U31966 (N_31966,N_22310,N_29292);
or U31967 (N_31967,N_28280,N_22281);
nand U31968 (N_31968,N_24924,N_20540);
nor U31969 (N_31969,N_29731,N_23115);
nor U31970 (N_31970,N_28128,N_22264);
xnor U31971 (N_31971,N_26115,N_21052);
nand U31972 (N_31972,N_26114,N_25626);
and U31973 (N_31973,N_27704,N_28378);
and U31974 (N_31974,N_28053,N_25536);
and U31975 (N_31975,N_28766,N_29603);
and U31976 (N_31976,N_21592,N_28135);
nand U31977 (N_31977,N_21338,N_25364);
or U31978 (N_31978,N_29551,N_26965);
nor U31979 (N_31979,N_28891,N_29685);
and U31980 (N_31980,N_29982,N_20804);
or U31981 (N_31981,N_20618,N_29898);
xor U31982 (N_31982,N_24985,N_24826);
nor U31983 (N_31983,N_25799,N_20724);
or U31984 (N_31984,N_28183,N_24325);
or U31985 (N_31985,N_28646,N_22690);
and U31986 (N_31986,N_22363,N_26978);
nand U31987 (N_31987,N_20275,N_22728);
or U31988 (N_31988,N_22585,N_29138);
and U31989 (N_31989,N_25273,N_25836);
nor U31990 (N_31990,N_24881,N_26175);
nor U31991 (N_31991,N_23999,N_21897);
or U31992 (N_31992,N_29133,N_26444);
nor U31993 (N_31993,N_20095,N_23713);
nand U31994 (N_31994,N_22707,N_21452);
xor U31995 (N_31995,N_25485,N_28152);
xor U31996 (N_31996,N_29931,N_25258);
nor U31997 (N_31997,N_27394,N_21478);
nand U31998 (N_31998,N_25646,N_29823);
nand U31999 (N_31999,N_26264,N_25493);
xnor U32000 (N_32000,N_22513,N_23758);
xnor U32001 (N_32001,N_26032,N_26758);
and U32002 (N_32002,N_28515,N_28712);
and U32003 (N_32003,N_22514,N_25906);
xor U32004 (N_32004,N_24961,N_28355);
nor U32005 (N_32005,N_23268,N_24453);
or U32006 (N_32006,N_25330,N_28531);
and U32007 (N_32007,N_22023,N_28538);
xor U32008 (N_32008,N_23032,N_22978);
nand U32009 (N_32009,N_29544,N_23134);
and U32010 (N_32010,N_27994,N_29569);
and U32011 (N_32011,N_25188,N_21594);
nor U32012 (N_32012,N_29899,N_21694);
nand U32013 (N_32013,N_24852,N_24069);
xor U32014 (N_32014,N_22287,N_21472);
xor U32015 (N_32015,N_22533,N_24762);
xor U32016 (N_32016,N_23133,N_29574);
nand U32017 (N_32017,N_25305,N_20630);
nand U32018 (N_32018,N_25898,N_23850);
nand U32019 (N_32019,N_21550,N_28285);
nor U32020 (N_32020,N_21913,N_21308);
nand U32021 (N_32021,N_22531,N_26721);
nand U32022 (N_32022,N_24178,N_29228);
nand U32023 (N_32023,N_20567,N_24741);
and U32024 (N_32024,N_24995,N_29223);
nor U32025 (N_32025,N_20263,N_25772);
xnor U32026 (N_32026,N_27553,N_23860);
or U32027 (N_32027,N_29250,N_24224);
nor U32028 (N_32028,N_28426,N_25568);
nand U32029 (N_32029,N_26274,N_22296);
xor U32030 (N_32030,N_26765,N_29009);
nand U32031 (N_32031,N_24960,N_21309);
nand U32032 (N_32032,N_28307,N_28260);
nor U32033 (N_32033,N_29010,N_22213);
or U32034 (N_32034,N_23316,N_22494);
and U32035 (N_32035,N_28858,N_23745);
xnor U32036 (N_32036,N_21190,N_22558);
nand U32037 (N_32037,N_28217,N_23842);
xnor U32038 (N_32038,N_28562,N_24796);
nor U32039 (N_32039,N_29512,N_24036);
xnor U32040 (N_32040,N_26364,N_24153);
or U32041 (N_32041,N_20360,N_20791);
and U32042 (N_32042,N_25418,N_25809);
xor U32043 (N_32043,N_25647,N_25763);
nor U32044 (N_32044,N_21247,N_20720);
or U32045 (N_32045,N_22209,N_22737);
nor U32046 (N_32046,N_25533,N_25380);
nand U32047 (N_32047,N_24567,N_27497);
and U32048 (N_32048,N_24044,N_20246);
or U32049 (N_32049,N_21851,N_24730);
nand U32050 (N_32050,N_29695,N_27821);
nand U32051 (N_32051,N_25819,N_23862);
nor U32052 (N_32052,N_22323,N_27163);
nor U32053 (N_32053,N_22456,N_22671);
xor U32054 (N_32054,N_25849,N_23020);
and U32055 (N_32055,N_20929,N_23765);
nor U32056 (N_32056,N_21882,N_27048);
or U32057 (N_32057,N_27341,N_21652);
nand U32058 (N_32058,N_23282,N_29953);
or U32059 (N_32059,N_29418,N_27294);
xor U32060 (N_32060,N_22966,N_28113);
xor U32061 (N_32061,N_25939,N_22170);
nand U32062 (N_32062,N_25296,N_27118);
and U32063 (N_32063,N_21812,N_23194);
and U32064 (N_32064,N_26118,N_21972);
xnor U32065 (N_32065,N_25392,N_28581);
nand U32066 (N_32066,N_21892,N_26393);
nor U32067 (N_32067,N_22409,N_20171);
or U32068 (N_32068,N_26857,N_23051);
xor U32069 (N_32069,N_20549,N_29836);
and U32070 (N_32070,N_23446,N_29454);
or U32071 (N_32071,N_25428,N_25203);
nor U32072 (N_32072,N_24299,N_20083);
nand U32073 (N_32073,N_22113,N_20652);
or U32074 (N_32074,N_29584,N_28721);
nand U32075 (N_32075,N_20536,N_26728);
nor U32076 (N_32076,N_26179,N_22927);
and U32077 (N_32077,N_20065,N_25231);
nor U32078 (N_32078,N_22724,N_28701);
nand U32079 (N_32079,N_24928,N_26087);
xnor U32080 (N_32080,N_25167,N_24499);
nand U32081 (N_32081,N_21357,N_22266);
nand U32082 (N_32082,N_28392,N_22816);
xor U32083 (N_32083,N_27998,N_25594);
nor U32084 (N_32084,N_24625,N_26752);
xor U32085 (N_32085,N_23170,N_24883);
or U32086 (N_32086,N_27856,N_29919);
or U32087 (N_32087,N_23941,N_27485);
nand U32088 (N_32088,N_25230,N_29781);
xnor U32089 (N_32089,N_22380,N_22865);
or U32090 (N_32090,N_23946,N_26029);
nand U32091 (N_32091,N_29033,N_28702);
xnor U32092 (N_32092,N_20599,N_22349);
nor U32093 (N_32093,N_25479,N_22547);
xor U32094 (N_32094,N_21142,N_28408);
or U32095 (N_32095,N_29759,N_21736);
and U32096 (N_32096,N_26429,N_28121);
nand U32097 (N_32097,N_23763,N_27769);
nand U32098 (N_32098,N_26390,N_21155);
xnor U32099 (N_32099,N_21819,N_27667);
and U32100 (N_32100,N_22119,N_24511);
xor U32101 (N_32101,N_22856,N_20950);
xor U32102 (N_32102,N_23596,N_24496);
or U32103 (N_32103,N_26462,N_27529);
nor U32104 (N_32104,N_29198,N_28265);
or U32105 (N_32105,N_26735,N_25073);
nor U32106 (N_32106,N_25651,N_26835);
nor U32107 (N_32107,N_25661,N_26628);
nand U32108 (N_32108,N_26894,N_29486);
nor U32109 (N_32109,N_28843,N_20057);
nor U32110 (N_32110,N_21360,N_20934);
nor U32111 (N_32111,N_23543,N_28613);
xor U32112 (N_32112,N_26018,N_22679);
xnor U32113 (N_32113,N_20937,N_25232);
nor U32114 (N_32114,N_27284,N_28186);
nor U32115 (N_32115,N_21838,N_20326);
nand U32116 (N_32116,N_29017,N_23845);
nand U32117 (N_32117,N_26954,N_29441);
xor U32118 (N_32118,N_22315,N_24765);
nand U32119 (N_32119,N_26849,N_25121);
or U32120 (N_32120,N_29610,N_23810);
and U32121 (N_32121,N_23913,N_25239);
or U32122 (N_32122,N_22469,N_21174);
nor U32123 (N_32123,N_26757,N_22637);
or U32124 (N_32124,N_27986,N_22719);
xor U32125 (N_32125,N_20356,N_21373);
and U32126 (N_32126,N_23181,N_23984);
nand U32127 (N_32127,N_26262,N_26997);
or U32128 (N_32128,N_29960,N_20475);
nand U32129 (N_32129,N_28244,N_29237);
nor U32130 (N_32130,N_21707,N_26601);
nor U32131 (N_32131,N_25549,N_22369);
xor U32132 (N_32132,N_24626,N_25506);
nand U32133 (N_32133,N_23185,N_29482);
xor U32134 (N_32134,N_22150,N_20090);
nand U32135 (N_32135,N_24345,N_21393);
nor U32136 (N_32136,N_25550,N_24894);
or U32137 (N_32137,N_29844,N_28997);
and U32138 (N_32138,N_21103,N_21336);
xnor U32139 (N_32139,N_26110,N_29168);
and U32140 (N_32140,N_26976,N_24136);
xnor U32141 (N_32141,N_27432,N_28842);
xor U32142 (N_32142,N_29099,N_28683);
and U32143 (N_32143,N_28505,N_21799);
or U32144 (N_32144,N_21764,N_29478);
or U32145 (N_32145,N_20654,N_23232);
nor U32146 (N_32146,N_26574,N_29993);
xor U32147 (N_32147,N_20307,N_22301);
nor U32148 (N_32148,N_29191,N_20429);
xor U32149 (N_32149,N_29970,N_20683);
or U32150 (N_32150,N_27375,N_23521);
nand U32151 (N_32151,N_26014,N_21909);
nor U32152 (N_32152,N_29474,N_27749);
nand U32153 (N_32153,N_26643,N_29555);
xor U32154 (N_32154,N_23529,N_21394);
nor U32155 (N_32155,N_29306,N_24202);
or U32156 (N_32156,N_20121,N_23360);
and U32157 (N_32157,N_28942,N_24198);
nor U32158 (N_32158,N_25988,N_25785);
nand U32159 (N_32159,N_24514,N_28863);
and U32160 (N_32160,N_29667,N_24996);
nor U32161 (N_32161,N_25372,N_26413);
nor U32162 (N_32162,N_24830,N_26547);
or U32163 (N_32163,N_29896,N_20718);
nor U32164 (N_32164,N_24068,N_24290);
nor U32165 (N_32165,N_22009,N_21626);
nor U32166 (N_32166,N_23139,N_23848);
xor U32167 (N_32167,N_29238,N_23155);
nor U32168 (N_32168,N_23725,N_27101);
nor U32169 (N_32169,N_26951,N_23788);
xnor U32170 (N_32170,N_23504,N_20570);
and U32171 (N_32171,N_24849,N_21380);
xnor U32172 (N_32172,N_26005,N_26260);
or U32173 (N_32173,N_20397,N_24361);
xnor U32174 (N_32174,N_20273,N_20785);
nand U32175 (N_32175,N_29111,N_24620);
or U32176 (N_32176,N_29670,N_27963);
and U32177 (N_32177,N_22552,N_26186);
nor U32178 (N_32178,N_26113,N_21091);
or U32179 (N_32179,N_27240,N_25501);
or U32180 (N_32180,N_20741,N_21289);
and U32181 (N_32181,N_25590,N_23011);
or U32182 (N_32182,N_29366,N_23910);
xor U32183 (N_32183,N_26949,N_29270);
nand U32184 (N_32184,N_20471,N_26199);
nand U32185 (N_32185,N_28616,N_22001);
xor U32186 (N_32186,N_26931,N_29469);
xor U32187 (N_32187,N_26896,N_21646);
nand U32188 (N_32188,N_22060,N_26235);
nor U32189 (N_32189,N_27327,N_26591);
xor U32190 (N_32190,N_23636,N_27901);
xnor U32191 (N_32191,N_24410,N_21540);
nor U32192 (N_32192,N_25540,N_21164);
nand U32193 (N_32193,N_22634,N_23948);
or U32194 (N_32194,N_25587,N_21938);
nand U32195 (N_32195,N_20591,N_25368);
nand U32196 (N_32196,N_24745,N_28640);
xor U32197 (N_32197,N_25499,N_29164);
nand U32198 (N_32198,N_24004,N_27959);
nand U32199 (N_32199,N_28456,N_21092);
xnor U32200 (N_32200,N_28289,N_26108);
and U32201 (N_32201,N_28022,N_25569);
nand U32202 (N_32202,N_29364,N_21253);
xnor U32203 (N_32203,N_28618,N_27717);
or U32204 (N_32204,N_20376,N_27757);
nor U32205 (N_32205,N_24832,N_28894);
or U32206 (N_32206,N_20845,N_27228);
or U32207 (N_32207,N_29515,N_22991);
xnor U32208 (N_32208,N_20737,N_27104);
nand U32209 (N_32209,N_23290,N_27705);
xor U32210 (N_32210,N_28336,N_21460);
nand U32211 (N_32211,N_24011,N_29484);
or U32212 (N_32212,N_22778,N_24401);
nor U32213 (N_32213,N_25902,N_28463);
or U32214 (N_32214,N_23444,N_22687);
nor U32215 (N_32215,N_27073,N_29842);
or U32216 (N_32216,N_24030,N_25343);
nand U32217 (N_32217,N_29280,N_21277);
xnor U32218 (N_32218,N_24656,N_22424);
nor U32219 (N_32219,N_25209,N_27766);
or U32220 (N_32220,N_24389,N_26779);
nand U32221 (N_32221,N_26958,N_27117);
and U32222 (N_32222,N_20372,N_25166);
nand U32223 (N_32223,N_24743,N_26922);
xor U32224 (N_32224,N_21032,N_29979);
nor U32225 (N_32225,N_21351,N_29465);
xnor U32226 (N_32226,N_24814,N_21037);
or U32227 (N_32227,N_28963,N_24598);
or U32228 (N_32228,N_20633,N_23270);
and U32229 (N_32229,N_22460,N_22155);
nand U32230 (N_32230,N_29185,N_21609);
nand U32231 (N_32231,N_27194,N_27173);
xor U32232 (N_32232,N_23222,N_28331);
nand U32233 (N_32233,N_29705,N_27680);
xnor U32234 (N_32234,N_24090,N_23936);
xor U32235 (N_32235,N_25096,N_21969);
and U32236 (N_32236,N_25697,N_21870);
xnor U32237 (N_32237,N_29749,N_24777);
xor U32238 (N_32238,N_21810,N_21401);
nand U32239 (N_32239,N_28151,N_29497);
or U32240 (N_32240,N_20444,N_29432);
and U32241 (N_32241,N_26333,N_20712);
xor U32242 (N_32242,N_22971,N_22306);
xor U32243 (N_32243,N_26457,N_26529);
nor U32244 (N_32244,N_21188,N_28620);
nand U32245 (N_32245,N_26678,N_26236);
xor U32246 (N_32246,N_27344,N_29804);
nand U32247 (N_32247,N_22491,N_20764);
nand U32248 (N_32248,N_25820,N_20927);
or U32249 (N_32249,N_21372,N_22238);
xor U32250 (N_32250,N_20071,N_23880);
or U32251 (N_32251,N_26790,N_27140);
nor U32252 (N_32252,N_29814,N_25153);
or U32253 (N_32253,N_29068,N_25921);
or U32254 (N_32254,N_22762,N_24429);
nor U32255 (N_32255,N_23419,N_25893);
nor U32256 (N_32256,N_20290,N_21787);
xnor U32257 (N_32257,N_22429,N_21802);
or U32258 (N_32258,N_24901,N_27764);
or U32259 (N_32259,N_25441,N_27633);
nor U32260 (N_32260,N_21379,N_29106);
nand U32261 (N_32261,N_22582,N_24161);
nor U32262 (N_32262,N_22953,N_23105);
or U32263 (N_32263,N_22632,N_22819);
nand U32264 (N_32264,N_23180,N_23220);
or U32265 (N_32265,N_26400,N_21503);
nand U32266 (N_32266,N_24316,N_20455);
and U32267 (N_32267,N_24214,N_23042);
and U32268 (N_32268,N_25388,N_23738);
nor U32269 (N_32269,N_25735,N_24652);
xnor U32270 (N_32270,N_29767,N_20005);
nor U32271 (N_32271,N_22276,N_22492);
xor U32272 (N_32272,N_21823,N_20760);
xnor U32273 (N_32273,N_21237,N_29739);
nor U32274 (N_32274,N_27635,N_24318);
nor U32275 (N_32275,N_26615,N_26769);
or U32276 (N_32276,N_25847,N_24392);
nor U32277 (N_32277,N_26125,N_28452);
nand U32278 (N_32278,N_28775,N_23071);
nor U32279 (N_32279,N_22970,N_24550);
or U32280 (N_32280,N_22888,N_21613);
or U32281 (N_32281,N_25152,N_22178);
nor U32282 (N_32282,N_22641,N_24867);
nor U32283 (N_32283,N_26232,N_24204);
and U32284 (N_32284,N_29859,N_23507);
nor U32285 (N_32285,N_23591,N_24253);
or U32286 (N_32286,N_25331,N_23030);
nand U32287 (N_32287,N_27883,N_23226);
xnor U32288 (N_32288,N_27815,N_28465);
and U32289 (N_32289,N_28083,N_25271);
and U32290 (N_32290,N_24640,N_24967);
and U32291 (N_32291,N_23203,N_27936);
xnor U32292 (N_32292,N_22134,N_24418);
nand U32293 (N_32293,N_21529,N_24847);
nand U32294 (N_32294,N_22827,N_28480);
nor U32295 (N_32295,N_26093,N_28557);
nor U32296 (N_32296,N_23617,N_27398);
and U32297 (N_32297,N_24129,N_29003);
xnor U32298 (N_32298,N_20489,N_26028);
nor U32299 (N_32299,N_22056,N_26937);
nor U32300 (N_32300,N_20740,N_21759);
or U32301 (N_32301,N_21363,N_23896);
or U32302 (N_32302,N_21242,N_21466);
xor U32303 (N_32303,N_21888,N_20151);
xnor U32304 (N_32304,N_29341,N_28417);
nand U32305 (N_32305,N_26515,N_28665);
nand U32306 (N_32306,N_23755,N_21198);
nor U32307 (N_32307,N_21928,N_23685);
xnor U32308 (N_32308,N_26607,N_29550);
xor U32309 (N_32309,N_22537,N_25008);
or U32310 (N_32310,N_21051,N_29761);
nor U32311 (N_32311,N_26694,N_21549);
nand U32312 (N_32312,N_28749,N_29917);
xor U32313 (N_32313,N_26676,N_24879);
and U32314 (N_32314,N_24355,N_22195);
or U32315 (N_32315,N_21284,N_28299);
or U32316 (N_32316,N_20539,N_24284);
nand U32317 (N_32317,N_20285,N_29691);
nand U32318 (N_32318,N_26430,N_29423);
xor U32319 (N_32319,N_25444,N_24428);
xor U32320 (N_32320,N_26496,N_20183);
nor U32321 (N_32321,N_20446,N_26780);
or U32322 (N_32322,N_27451,N_25701);
or U32323 (N_32323,N_29862,N_28680);
and U32324 (N_32324,N_23877,N_28928);
or U32325 (N_32325,N_25001,N_26148);
xnor U32326 (N_32326,N_23260,N_22215);
and U32327 (N_32327,N_23068,N_25131);
or U32328 (N_32328,N_23457,N_28829);
or U32329 (N_32329,N_27748,N_20971);
or U32330 (N_32330,N_22813,N_25339);
nand U32331 (N_32331,N_26081,N_27965);
nor U32332 (N_32332,N_26482,N_21131);
nand U32333 (N_32333,N_25378,N_24549);
or U32334 (N_32334,N_27990,N_29227);
xnor U32335 (N_32335,N_23816,N_29102);
nand U32336 (N_32336,N_20328,N_24261);
nand U32337 (N_32337,N_29873,N_29522);
xor U32338 (N_32338,N_28101,N_26720);
or U32339 (N_32339,N_28235,N_28645);
and U32340 (N_32340,N_27289,N_23477);
nor U32341 (N_32341,N_21962,N_25200);
nand U32342 (N_32342,N_25495,N_26940);
nor U32343 (N_32343,N_27312,N_21265);
and U32344 (N_32344,N_28400,N_23441);
and U32345 (N_32345,N_24376,N_20587);
nor U32346 (N_32346,N_27519,N_24266);
nor U32347 (N_32347,N_24752,N_22099);
xnor U32348 (N_32348,N_20781,N_27914);
xnor U32349 (N_32349,N_25620,N_21526);
nor U32350 (N_32350,N_20642,N_29996);
or U32351 (N_32351,N_28929,N_24874);
or U32352 (N_32352,N_22346,N_20479);
and U32353 (N_32353,N_27995,N_21960);
nand U32354 (N_32354,N_28276,N_27338);
or U32355 (N_32355,N_26689,N_22061);
or U32356 (N_32356,N_29682,N_22660);
xor U32357 (N_32357,N_29352,N_21587);
and U32358 (N_32358,N_22846,N_22064);
or U32359 (N_32359,N_24176,N_25919);
and U32360 (N_32360,N_26101,N_22842);
and U32361 (N_32361,N_27139,N_26805);
xor U32362 (N_32362,N_20809,N_29679);
and U32363 (N_32363,N_29517,N_25973);
xnor U32364 (N_32364,N_23840,N_27893);
and U32365 (N_32365,N_23109,N_25468);
or U32366 (N_32366,N_22828,N_24917);
and U32367 (N_32367,N_25838,N_22957);
nand U32368 (N_32368,N_20551,N_23537);
nand U32369 (N_32369,N_25628,N_23428);
and U32370 (N_32370,N_21057,N_29808);
or U32371 (N_32371,N_26094,N_22156);
or U32372 (N_32372,N_28840,N_28994);
nor U32373 (N_32373,N_25281,N_22102);
nand U32374 (N_32374,N_27019,N_27150);
nand U32375 (N_32375,N_27017,N_29249);
nor U32376 (N_32376,N_28604,N_29188);
xnor U32377 (N_32377,N_21793,N_29813);
nor U32378 (N_32378,N_27550,N_24585);
nor U32379 (N_32379,N_21982,N_27067);
xnor U32380 (N_32380,N_28602,N_29624);
nor U32381 (N_32381,N_28131,N_27756);
xor U32382 (N_32382,N_28314,N_20451);
and U32383 (N_32383,N_22569,N_22618);
nand U32384 (N_32384,N_23406,N_22083);
xnor U32385 (N_32385,N_22062,N_20981);
nand U32386 (N_32386,N_29255,N_29458);
nand U32387 (N_32387,N_28729,N_23217);
or U32388 (N_32388,N_28687,N_20366);
and U32389 (N_32389,N_23214,N_29607);
xor U32390 (N_32390,N_22482,N_29595);
xor U32391 (N_32391,N_24711,N_20100);
and U32392 (N_32392,N_20951,N_22457);
xor U32393 (N_32393,N_28150,N_28710);
or U32394 (N_32394,N_24663,N_27759);
and U32395 (N_32395,N_22372,N_20953);
and U32396 (N_32396,N_29453,N_22594);
nor U32397 (N_32397,N_29883,N_24190);
nand U32398 (N_32398,N_26311,N_26443);
nand U32399 (N_32399,N_24125,N_29611);
nor U32400 (N_32400,N_23117,N_21513);
nand U32401 (N_32401,N_24031,N_21757);
nand U32402 (N_32402,N_29552,N_29273);
and U32403 (N_32403,N_20243,N_22981);
xor U32404 (N_32404,N_26035,N_25790);
xor U32405 (N_32405,N_23593,N_28402);
nand U32406 (N_32406,N_25503,N_28746);
and U32407 (N_32407,N_26476,N_25888);
xnor U32408 (N_32408,N_26389,N_29797);
xnor U32409 (N_32409,N_20002,N_22780);
nor U32410 (N_32410,N_21381,N_23502);
nor U32411 (N_32411,N_22652,N_24977);
and U32412 (N_32412,N_25684,N_25289);
or U32413 (N_32413,N_24740,N_26056);
xor U32414 (N_32414,N_28428,N_26859);
and U32415 (N_32415,N_26499,N_27506);
nor U32416 (N_32416,N_21413,N_23673);
xor U32417 (N_32417,N_22532,N_24877);
or U32418 (N_32418,N_27217,N_21601);
xnor U32419 (N_32419,N_29472,N_22168);
nor U32420 (N_32420,N_24701,N_21809);
nor U32421 (N_32421,N_29506,N_20431);
and U32422 (N_32422,N_28200,N_22298);
nand U32423 (N_32423,N_25991,N_29281);
and U32424 (N_32424,N_23852,N_23035);
and U32425 (N_32425,N_26556,N_20902);
xor U32426 (N_32426,N_23036,N_22567);
xor U32427 (N_32427,N_22365,N_20084);
and U32428 (N_32428,N_20905,N_29721);
nor U32429 (N_32429,N_22324,N_22772);
nand U32430 (N_32430,N_29688,N_20223);
and U32431 (N_32431,N_24159,N_28553);
nor U32432 (N_32432,N_27459,N_24048);
and U32433 (N_32433,N_27495,N_22327);
and U32434 (N_32434,N_22961,N_29858);
and U32435 (N_32435,N_24180,N_29530);
nand U32436 (N_32436,N_27114,N_24262);
xor U32437 (N_32437,N_25795,N_28292);
xnor U32438 (N_32438,N_26398,N_26882);
nor U32439 (N_32439,N_29295,N_27407);
or U32440 (N_32440,N_27583,N_21524);
nand U32441 (N_32441,N_20638,N_27798);
nor U32442 (N_32442,N_25732,N_29020);
or U32443 (N_32443,N_21539,N_29427);
or U32444 (N_32444,N_29051,N_21769);
nand U32445 (N_32445,N_22633,N_25214);
or U32446 (N_32446,N_21776,N_23243);
nor U32447 (N_32447,N_21791,N_22503);
nand U32448 (N_32448,N_26630,N_20615);
nand U32449 (N_32449,N_22449,N_22568);
nor U32450 (N_32450,N_24794,N_26953);
or U32451 (N_32451,N_24856,N_23640);
or U32452 (N_32452,N_23093,N_28931);
nor U32453 (N_32453,N_21390,N_24006);
and U32454 (N_32454,N_23033,N_29243);
and U32455 (N_32455,N_22269,N_22600);
nor U32456 (N_32456,N_20715,N_21606);
xor U32457 (N_32457,N_23374,N_25534);
xor U32458 (N_32458,N_26846,N_28365);
nor U32459 (N_32459,N_24593,N_25108);
or U32460 (N_32460,N_23970,N_29908);
or U32461 (N_32461,N_23804,N_24671);
nand U32462 (N_32462,N_20476,N_23404);
and U32463 (N_32463,N_25865,N_23990);
nand U32464 (N_32464,N_27062,N_23904);
or U32465 (N_32465,N_23271,N_22672);
nand U32466 (N_32466,N_21305,N_22554);
nand U32467 (N_32467,N_25935,N_29383);
xnor U32468 (N_32468,N_20663,N_27377);
or U32469 (N_32469,N_24387,N_23935);
and U32470 (N_32470,N_24400,N_20097);
nand U32471 (N_32471,N_29548,N_22551);
nor U32472 (N_32472,N_27611,N_25461);
nor U32473 (N_32473,N_21661,N_29736);
and U32474 (N_32474,N_24363,N_28360);
xnor U32475 (N_32475,N_23215,N_23829);
or U32476 (N_32476,N_22625,N_23744);
or U32477 (N_32477,N_22471,N_25598);
nor U32478 (N_32478,N_24349,N_22802);
nor U32479 (N_32479,N_24130,N_29901);
nor U32480 (N_32480,N_29846,N_29029);
nor U32481 (N_32481,N_21375,N_27125);
xor U32482 (N_32482,N_24451,N_26917);
or U32483 (N_32483,N_28722,N_20671);
nand U32484 (N_32484,N_23868,N_26138);
xnor U32485 (N_32485,N_25119,N_20870);
nor U32486 (N_32486,N_26352,N_23891);
or U32487 (N_32487,N_23664,N_21794);
nand U32488 (N_32488,N_27437,N_21682);
or U32489 (N_32489,N_21132,N_28330);
nand U32490 (N_32490,N_20861,N_28649);
nor U32491 (N_32491,N_28886,N_28781);
xnor U32492 (N_32492,N_25491,N_25854);
nand U32493 (N_32493,N_22079,N_22378);
nand U32494 (N_32494,N_24263,N_27421);
nor U32495 (N_32495,N_24709,N_25716);
nor U32496 (N_32496,N_29415,N_24792);
and U32497 (N_32497,N_27443,N_23875);
and U32498 (N_32498,N_26315,N_24965);
nor U32499 (N_32499,N_28624,N_21980);
nor U32500 (N_32500,N_28811,N_23826);
and U32501 (N_32501,N_23314,N_25489);
or U32502 (N_32502,N_21298,N_24820);
or U32503 (N_32503,N_26386,N_20520);
nor U32504 (N_32504,N_27852,N_21102);
nand U32505 (N_32505,N_27830,N_28211);
xnor U32506 (N_32506,N_25694,N_26909);
or U32507 (N_32507,N_29419,N_22862);
and U32508 (N_32508,N_29834,N_21418);
nor U32509 (N_32509,N_29833,N_29129);
nand U32510 (N_32510,N_22151,N_22257);
and U32511 (N_32511,N_20464,N_24070);
xor U32512 (N_32512,N_27287,N_22321);
or U32513 (N_32513,N_21953,N_24060);
and U32514 (N_32514,N_27598,N_23680);
nand U32515 (N_32515,N_23124,N_22610);
and U32516 (N_32516,N_22362,N_26977);
and U32517 (N_32517,N_29398,N_27954);
and U32518 (N_32518,N_23759,N_20822);
and U32519 (N_32519,N_20572,N_27109);
or U32520 (N_32520,N_22091,N_29242);
nor U32521 (N_32521,N_25079,N_20703);
xnor U32522 (N_32522,N_26994,N_23154);
and U32523 (N_32523,N_29360,N_25171);
xnor U32524 (N_32524,N_25983,N_24484);
nand U32525 (N_32525,N_24019,N_20577);
nand U32526 (N_32526,N_24823,N_27226);
nand U32527 (N_32527,N_25282,N_25650);
nand U32528 (N_32528,N_24582,N_20437);
or U32529 (N_32529,N_22830,N_25283);
nand U32530 (N_32530,N_20417,N_24013);
and U32531 (N_32531,N_29601,N_21406);
nor U32532 (N_32532,N_29755,N_25578);
nor U32533 (N_32533,N_26181,N_28008);
nor U32534 (N_32534,N_29965,N_24043);
or U32535 (N_32535,N_21334,N_23206);
and U32536 (N_32536,N_22628,N_27578);
and U32537 (N_32537,N_29631,N_23375);
or U32538 (N_32538,N_21419,N_24443);
and U32539 (N_32539,N_20207,N_27504);
xor U32540 (N_32540,N_21821,N_21327);
and U32541 (N_32541,N_24196,N_26497);
xor U32542 (N_32542,N_20402,N_23378);
or U32543 (N_32543,N_21864,N_25633);
and U32544 (N_32544,N_22440,N_28637);
and U32545 (N_32545,N_27496,N_24866);
nor U32546 (N_32546,N_24343,N_27726);
or U32547 (N_32547,N_26881,N_21708);
nand U32548 (N_32548,N_24718,N_27126);
nand U32549 (N_32549,N_22553,N_26844);
nand U32550 (N_32550,N_28848,N_22574);
nor U32551 (N_32551,N_20560,N_29714);
nand U32552 (N_32552,N_22334,N_24411);
and U32553 (N_32553,N_27732,N_20185);
and U32554 (N_32554,N_21619,N_25290);
or U32555 (N_32555,N_22093,N_20412);
nand U32556 (N_32556,N_22620,N_24497);
and U32557 (N_32557,N_26996,N_27237);
nand U32558 (N_32558,N_27527,N_22361);
nor U32559 (N_32559,N_24646,N_21088);
nor U32560 (N_32560,N_24992,N_26196);
or U32561 (N_32561,N_22578,N_22441);
nand U32562 (N_32562,N_21239,N_24467);
nor U32563 (N_32563,N_29050,N_29342);
nor U32564 (N_32564,N_25156,N_28713);
or U32565 (N_32565,N_25824,N_21470);
or U32566 (N_32566,N_23147,N_21544);
xor U32567 (N_32567,N_24799,N_20315);
nand U32568 (N_32568,N_26787,N_23364);
nand U32569 (N_32569,N_23899,N_25012);
xnor U32570 (N_32570,N_21603,N_29877);
nor U32571 (N_32571,N_20350,N_24530);
xor U32572 (N_32572,N_29838,N_27466);
and U32573 (N_32573,N_25375,N_27110);
or U32574 (N_32574,N_24769,N_20484);
or U32575 (N_32575,N_20853,N_20682);
nand U32576 (N_32576,N_25065,N_26183);
nand U32577 (N_32577,N_25622,N_25123);
nor U32578 (N_32578,N_29652,N_27010);
nor U32579 (N_32579,N_24482,N_22984);
nor U32580 (N_32580,N_24683,N_27233);
nand U32581 (N_32581,N_24614,N_21706);
or U32582 (N_32582,N_22851,N_24244);
nand U32583 (N_32583,N_21950,N_25178);
xor U32584 (N_32584,N_28789,N_23769);
xor U32585 (N_32585,N_27115,N_27028);
or U32586 (N_32586,N_24865,N_29766);
nor U32587 (N_32587,N_24210,N_25173);
or U32588 (N_32588,N_26756,N_28019);
and U32589 (N_32589,N_20890,N_21758);
and U32590 (N_32590,N_23070,N_28320);
and U32591 (N_32591,N_29132,N_21154);
xnor U32592 (N_32592,N_25168,N_21683);
nand U32593 (N_32593,N_27409,N_21885);
or U32594 (N_32594,N_25344,N_29825);
nor U32595 (N_32595,N_22760,N_24969);
nand U32596 (N_32596,N_28072,N_25928);
nor U32597 (N_32597,N_25207,N_24481);
and U32598 (N_32598,N_24333,N_20020);
nand U32599 (N_32599,N_22450,N_29674);
and U32600 (N_32600,N_25821,N_20447);
and U32601 (N_32601,N_22965,N_27685);
xnor U32602 (N_32602,N_22857,N_26905);
or U32603 (N_32603,N_23141,N_27837);
and U32604 (N_32604,N_20202,N_24427);
nand U32605 (N_32605,N_23515,N_26465);
and U32606 (N_32606,N_25267,N_20574);
or U32607 (N_32607,N_24146,N_28037);
nor U32608 (N_32608,N_23028,N_28625);
xnor U32609 (N_32609,N_21398,N_22896);
nand U32610 (N_32610,N_20048,N_20311);
or U32611 (N_32611,N_28909,N_27930);
or U32612 (N_32612,N_27033,N_20824);
or U32613 (N_32613,N_25165,N_21869);
nand U32614 (N_32614,N_28048,N_29394);
nor U32615 (N_32615,N_25563,N_24222);
nand U32616 (N_32616,N_27675,N_29049);
and U32617 (N_32617,N_22137,N_22935);
or U32618 (N_32618,N_20686,N_25840);
and U32619 (N_32619,N_21233,N_25673);
xor U32620 (N_32620,N_26623,N_29646);
nor U32621 (N_32621,N_26948,N_25867);
or U32622 (N_32622,N_27205,N_25773);
nand U32623 (N_32623,N_26140,N_21862);
or U32624 (N_32624,N_28554,N_22749);
nor U32625 (N_32625,N_20024,N_25212);
xor U32626 (N_32626,N_22046,N_27405);
or U32627 (N_32627,N_21185,N_27328);
or U32628 (N_32628,N_25933,N_28380);
xnor U32629 (N_32629,N_26930,N_25555);
nand U32630 (N_32630,N_29201,N_26142);
nand U32631 (N_32631,N_23116,N_22803);
nor U32632 (N_32632,N_24460,N_21170);
xor U32633 (N_32633,N_29575,N_23900);
or U32634 (N_32634,N_28945,N_28596);
nand U32635 (N_32635,N_27858,N_27422);
nand U32636 (N_32636,N_20468,N_22354);
nor U32637 (N_32637,N_20166,N_21217);
xnor U32638 (N_32638,N_25269,N_21148);
and U32639 (N_32639,N_27214,N_22263);
nand U32640 (N_32640,N_26549,N_27817);
or U32641 (N_32641,N_25420,N_20198);
or U32642 (N_32642,N_25627,N_23265);
xor U32643 (N_32643,N_26838,N_25264);
nor U32644 (N_32644,N_23844,N_20941);
nor U32645 (N_32645,N_23715,N_21412);
nand U32646 (N_32646,N_27851,N_24631);
nand U32647 (N_32647,N_28329,N_21288);
nand U32648 (N_32648,N_20452,N_21922);
nor U32649 (N_32649,N_28660,N_29640);
xor U32650 (N_32650,N_22197,N_22177);
and U32651 (N_32651,N_24300,N_27913);
or U32652 (N_32652,N_26565,N_25220);
nand U32653 (N_32653,N_29035,N_25986);
or U32654 (N_32654,N_27262,N_20722);
xor U32655 (N_32655,N_25576,N_20069);
nor U32656 (N_32656,N_26395,N_26806);
and U32657 (N_32657,N_28185,N_21642);
nor U32658 (N_32658,N_24380,N_22249);
xnor U32659 (N_32659,N_29459,N_27760);
or U32660 (N_32660,N_22715,N_27559);
xnor U32661 (N_32661,N_24197,N_25531);
or U32662 (N_32662,N_24710,N_20150);
nand U32663 (N_32663,N_26985,N_20030);
nand U32664 (N_32664,N_28094,N_20359);
nor U32665 (N_32665,N_23790,N_23006);
xnor U32666 (N_32666,N_24639,N_29190);
nand U32667 (N_32667,N_28787,N_21910);
and U32668 (N_32668,N_28214,N_22942);
or U32669 (N_32669,N_28893,N_22792);
nor U32670 (N_32670,N_23151,N_24731);
nor U32671 (N_32671,N_28293,N_23869);
and U32672 (N_32672,N_21886,N_21156);
and U32673 (N_32673,N_21673,N_23053);
xor U32674 (N_32674,N_25279,N_23906);
nor U32675 (N_32675,N_22131,N_21620);
nor U32676 (N_32676,N_24882,N_23866);
nor U32677 (N_32677,N_23674,N_27389);
nor U32678 (N_32678,N_27579,N_26539);
or U32679 (N_32679,N_24142,N_26360);
xor U32680 (N_32680,N_20862,N_23095);
xnor U32681 (N_32681,N_24541,N_28796);
or U32682 (N_32682,N_24012,N_20991);
xor U32683 (N_32683,N_29609,N_24838);
nor U32684 (N_32684,N_22408,N_27755);
nor U32685 (N_32685,N_29986,N_29320);
or U32686 (N_32686,N_29694,N_28516);
or U32687 (N_32687,N_23686,N_25303);
and U32688 (N_32688,N_20157,N_22191);
or U32689 (N_32689,N_24134,N_29822);
and U32690 (N_32690,N_24848,N_23104);
nand U32691 (N_32691,N_24282,N_28925);
and U32692 (N_32692,N_22216,N_22713);
and U32693 (N_32693,N_25775,N_28504);
or U32694 (N_32694,N_23157,N_26450);
and U32695 (N_32695,N_20003,N_24257);
nor U32696 (N_32696,N_20625,N_20282);
nor U32697 (N_32697,N_29567,N_26898);
nand U32698 (N_32698,N_28609,N_23927);
xnor U32699 (N_32699,N_20865,N_21342);
nor U32700 (N_32700,N_23261,N_24230);
and U32701 (N_32701,N_27975,N_22383);
and U32702 (N_32702,N_23439,N_27896);
xor U32703 (N_32703,N_24169,N_24246);
nor U32704 (N_32704,N_28927,N_27082);
nor U32705 (N_32705,N_21763,N_24510);
nand U32706 (N_32706,N_28975,N_27993);
nor U32707 (N_32707,N_22478,N_21414);
or U32708 (N_32708,N_23930,N_28544);
or U32709 (N_32709,N_23538,N_23670);
and U32710 (N_32710,N_23182,N_28561);
xnor U32711 (N_32711,N_21257,N_26921);
or U32712 (N_32712,N_21658,N_27463);
nor U32713 (N_32713,N_26648,N_29287);
nor U32714 (N_32714,N_25886,N_29643);
or U32715 (N_32715,N_27445,N_22786);
nand U32716 (N_32716,N_21097,N_23372);
nor U32717 (N_32717,N_23110,N_22453);
and U32718 (N_32718,N_29650,N_24057);
nand U32719 (N_32719,N_27488,N_20651);
nor U32720 (N_32720,N_24955,N_22250);
nor U32721 (N_32721,N_23541,N_28936);
xor U32722 (N_32722,N_24421,N_22683);
and U32723 (N_32723,N_23128,N_29639);
nand U32724 (N_32724,N_26992,N_23431);
and U32725 (N_32725,N_23903,N_24672);
and U32726 (N_32726,N_22859,N_25382);
nor U32727 (N_32727,N_29442,N_26328);
xnor U32728 (N_32728,N_24241,N_27637);
nor U32729 (N_32729,N_27272,N_23292);
and U32730 (N_32730,N_25894,N_23939);
xnor U32731 (N_32731,N_28084,N_27143);
xor U32732 (N_32732,N_29502,N_23474);
or U32733 (N_32733,N_27260,N_23678);
and U32734 (N_32734,N_27866,N_29837);
or U32735 (N_32735,N_29816,N_26807);
xnor U32736 (N_32736,N_27030,N_23343);
nand U32737 (N_32737,N_24168,N_27801);
and U32738 (N_32738,N_22451,N_21019);
nor U32739 (N_32739,N_25924,N_28075);
nand U32740 (N_32740,N_28567,N_23693);
and U32741 (N_32741,N_22403,N_25413);
or U32742 (N_32742,N_20987,N_26732);
and U32743 (N_32743,N_26785,N_27576);
nand U32744 (N_32744,N_26160,N_28144);
or U32745 (N_32745,N_20755,N_26864);
xor U32746 (N_32746,N_26071,N_25526);
and U32747 (N_32747,N_22108,N_25544);
and U32748 (N_32748,N_25107,N_25456);
xnor U32749 (N_32749,N_21245,N_27668);
xor U32750 (N_32750,N_27411,N_21647);
or U32751 (N_32751,N_27458,N_23355);
nand U32752 (N_32752,N_22399,N_27711);
and U32753 (N_32753,N_21047,N_23323);
and U32754 (N_32754,N_27096,N_24844);
xnor U32755 (N_32755,N_25363,N_20628);
nor U32756 (N_32756,N_21684,N_21283);
nand U32757 (N_32757,N_22575,N_20025);
and U32758 (N_32758,N_21082,N_29309);
xnor U32759 (N_32759,N_25376,N_29386);
nor U32760 (N_32760,N_21622,N_20921);
nand U32761 (N_32761,N_26080,N_23077);
and U32762 (N_32762,N_22797,N_24571);
or U32763 (N_32763,N_23702,N_29044);
nor U32764 (N_32764,N_24737,N_24596);
xor U32765 (N_32765,N_20901,N_22161);
nor U32766 (N_32766,N_26635,N_29359);
xnor U32767 (N_32767,N_27535,N_22282);
xor U32768 (N_32768,N_22226,N_22352);
or U32769 (N_32769,N_26550,N_27362);
and U32770 (N_32770,N_27490,N_21525);
and U32771 (N_32771,N_23272,N_23570);
nor U32772 (N_32772,N_20320,N_27383);
and U32773 (N_32773,N_20864,N_28168);
or U32774 (N_32774,N_22644,N_27531);
or U32775 (N_32775,N_29994,N_25090);
xor U32776 (N_32776,N_21485,N_23523);
xor U32777 (N_32777,N_26919,N_28012);
and U32778 (N_32778,N_26466,N_22016);
nand U32779 (N_32779,N_28896,N_29907);
nand U32780 (N_32780,N_29703,N_20790);
or U32781 (N_32781,N_25446,N_26872);
xor U32782 (N_32782,N_28756,N_27505);
and U32783 (N_32783,N_25359,N_24902);
nand U32784 (N_32784,N_22184,N_24608);
and U32785 (N_32785,N_27268,N_23813);
or U32786 (N_32786,N_23394,N_25112);
or U32787 (N_32787,N_29109,N_20911);
or U32788 (N_32788,N_28496,N_20779);
xnor U32789 (N_32789,N_26935,N_22992);
xnor U32790 (N_32790,N_29974,N_20093);
nand U32791 (N_32791,N_24727,N_26797);
or U32792 (N_32792,N_28563,N_21573);
xor U32793 (N_32793,N_21415,N_20125);
and U32794 (N_32794,N_23369,N_26177);
xnor U32795 (N_32795,N_29408,N_27491);
and U32796 (N_32796,N_27567,N_23854);
or U32797 (N_32797,N_22425,N_25742);
or U32798 (N_32798,N_21671,N_23023);
or U32799 (N_32799,N_26712,N_22782);
nand U32800 (N_32800,N_28957,N_27043);
xor U32801 (N_32801,N_28705,N_28111);
nor U32802 (N_32802,N_29083,N_27938);
or U32803 (N_32803,N_25246,N_25517);
xnor U32804 (N_32804,N_23464,N_26233);
xnor U32805 (N_32805,N_26223,N_22598);
xnor U32806 (N_32806,N_20631,N_22710);
nor U32807 (N_32807,N_28193,N_28477);
or U32808 (N_32808,N_26437,N_29477);
and U32809 (N_32809,N_29189,N_25802);
or U32810 (N_32810,N_27295,N_27659);
nand U32811 (N_32811,N_24396,N_22467);
xnor U32812 (N_32812,N_22038,N_24270);
nor U32813 (N_32813,N_26811,N_23401);
or U32814 (N_32814,N_28939,N_25721);
nand U32815 (N_32815,N_27860,N_28035);
xnor U32816 (N_32816,N_25546,N_28204);
and U32817 (N_32817,N_25138,N_29025);
nor U32818 (N_32818,N_20406,N_20346);
nor U32819 (N_32819,N_27059,N_20799);
nor U32820 (N_32820,N_27835,N_24209);
and U32821 (N_32821,N_23421,N_25789);
or U32822 (N_32822,N_29471,N_28814);
and U32823 (N_32823,N_28175,N_27087);
and U32824 (N_32824,N_27251,N_21120);
or U32825 (N_32825,N_21162,N_23918);
or U32826 (N_32826,N_26671,N_29061);
xor U32827 (N_32827,N_27083,N_21294);
or U32828 (N_32828,N_28728,N_29456);
or U32829 (N_32829,N_26595,N_29411);
nor U32830 (N_32830,N_27454,N_24050);
and U32831 (N_32831,N_25450,N_23402);
nor U32832 (N_32832,N_26592,N_22314);
nor U32833 (N_32833,N_22730,N_23581);
and U32834 (N_32834,N_20938,N_21444);
nand U32835 (N_32835,N_21297,N_24395);
nor U32836 (N_32836,N_27417,N_20139);
or U32837 (N_32837,N_24279,N_23513);
nand U32838 (N_32838,N_28517,N_27514);
or U32839 (N_32839,N_21391,N_22948);
nor U32840 (N_32840,N_20948,N_28238);
nand U32841 (N_32841,N_29572,N_25887);
nor U32842 (N_32842,N_28102,N_27402);
xnor U32843 (N_32843,N_28857,N_29002);
xnor U32844 (N_32844,N_28897,N_20796);
nor U32845 (N_32845,N_25941,N_24225);
xnor U32846 (N_32846,N_29773,N_29436);
nor U32847 (N_32847,N_23037,N_27779);
nand U32848 (N_32848,N_21923,N_28798);
and U32849 (N_32849,N_28935,N_21981);
xnor U32850 (N_32850,N_28632,N_28017);
xor U32851 (N_32851,N_21716,N_25145);
nand U32852 (N_32852,N_28877,N_28468);
xnor U32853 (N_32853,N_26571,N_23190);
and U32854 (N_32854,N_20099,N_24382);
xnor U32855 (N_32855,N_23497,N_23747);
xnor U32856 (N_32856,N_22043,N_26875);
and U32857 (N_32857,N_20407,N_20140);
nand U32858 (N_32858,N_23130,N_25974);
or U32859 (N_32859,N_25967,N_24203);
nand U32860 (N_32860,N_27399,N_23313);
nor U32861 (N_32861,N_28350,N_25106);
nor U32862 (N_32862,N_21817,N_20665);
nor U32863 (N_32863,N_28757,N_24693);
nand U32864 (N_32864,N_26901,N_20807);
nor U32865 (N_32865,N_22901,N_25738);
xor U32866 (N_32866,N_26340,N_24426);
nor U32867 (N_32867,N_29888,N_20894);
nand U32868 (N_32868,N_24956,N_27609);
and U32869 (N_32869,N_25222,N_20871);
and U32870 (N_32870,N_22025,N_27556);
or U32871 (N_32871,N_20391,N_26928);
xnor U32872 (N_32872,N_29718,N_27831);
and U32873 (N_32873,N_26276,N_22695);
and U32874 (N_32874,N_23952,N_27549);
and U32875 (N_32875,N_20576,N_24024);
nand U32876 (N_32876,N_22012,N_21824);
xnor U32877 (N_32877,N_22284,N_22821);
and U32878 (N_32878,N_27420,N_23284);
nor U32879 (N_32879,N_27621,N_21944);
xor U32880 (N_32880,N_23235,N_22381);
nand U32881 (N_32881,N_28959,N_23554);
or U32882 (N_32882,N_25322,N_21307);
and U32883 (N_32883,N_28431,N_22777);
and U32884 (N_32884,N_23367,N_27434);
nand U32885 (N_32885,N_28071,N_25723);
and U32886 (N_32886,N_25462,N_29095);
nand U32887 (N_32887,N_20404,N_22748);
and U32888 (N_32888,N_25437,N_22068);
xnor U32889 (N_32889,N_20805,N_20892);
xor U32890 (N_32890,N_27242,N_29875);
and U32891 (N_32891,N_20075,N_22721);
nor U32892 (N_32892,N_25114,N_25252);
nand U32893 (N_32893,N_21264,N_27273);
nor U32894 (N_32894,N_24379,N_25321);
nand U32895 (N_32895,N_23649,N_23320);
nand U32896 (N_32896,N_21231,N_27524);
xor U32897 (N_32897,N_25040,N_29354);
nor U32898 (N_32898,N_26472,N_21762);
nand U32899 (N_32899,N_20286,N_26891);
nand U32900 (N_32900,N_26511,N_24674);
or U32901 (N_32901,N_28381,N_22422);
and U32902 (N_32902,N_24391,N_26036);
and U32903 (N_32903,N_22286,N_26488);
or U32904 (N_32904,N_21740,N_25002);
or U32905 (N_32905,N_21081,N_20423);
xor U32906 (N_32906,N_27304,N_25554);
xnor U32907 (N_32907,N_26563,N_25473);
xor U32908 (N_32908,N_29118,N_25412);
xor U32909 (N_32909,N_22105,N_22657);
xnor U32910 (N_32910,N_20426,N_21805);
or U32911 (N_32911,N_26654,N_21669);
and U32912 (N_32912,N_21345,N_28932);
or U32913 (N_32913,N_22110,N_23764);
or U32914 (N_32914,N_21139,N_25254);
nand U32915 (N_32915,N_25643,N_25875);
xnor U32916 (N_32916,N_26538,N_26825);
or U32917 (N_32917,N_28157,N_29829);
or U32918 (N_32918,N_24472,N_29728);
and U32919 (N_32919,N_28667,N_27892);
xor U32920 (N_32920,N_24409,N_29438);
xnor U32921 (N_32921,N_27548,N_22718);
or U32922 (N_32922,N_22875,N_20900);
and U32923 (N_32923,N_22845,N_22316);
nand U32924 (N_32924,N_23983,N_22020);
nor U32925 (N_32925,N_20735,N_26863);
and U32926 (N_32926,N_28155,N_22697);
nor U32927 (N_32927,N_26692,N_20746);
xor U32928 (N_32928,N_22682,N_20957);
and U32929 (N_32929,N_21680,N_22601);
and U32930 (N_32930,N_26200,N_26059);
or U32931 (N_32931,N_24235,N_27134);
or U32932 (N_32932,N_27806,N_28834);
and U32933 (N_32933,N_22166,N_26627);
nand U32934 (N_32934,N_27250,N_21293);
or U32935 (N_32935,N_20252,N_20778);
nor U32936 (N_32936,N_23255,N_22340);
and U32937 (N_32937,N_26495,N_20582);
and U32938 (N_32938,N_22358,N_25329);
or U32939 (N_32939,N_27345,N_25788);
nor U32940 (N_32940,N_26762,N_22464);
and U32941 (N_32941,N_26217,N_21815);
nor U32942 (N_32942,N_20684,N_26535);
and U32943 (N_32943,N_24078,N_20653);
or U32944 (N_32944,N_20637,N_24661);
nor U32945 (N_32945,N_26597,N_21158);
nor U32946 (N_32946,N_22175,N_27544);
nand U32947 (N_32947,N_22885,N_28919);
or U32948 (N_32948,N_20299,N_26502);
nand U32949 (N_32949,N_26912,N_29108);
xor U32950 (N_32950,N_27888,N_25086);
xor U32951 (N_32951,N_22651,N_20973);
nor U32952 (N_32952,N_27269,N_20434);
and U32953 (N_32953,N_20700,N_24590);
nand U32954 (N_32954,N_20508,N_25257);
xor U32955 (N_32955,N_21416,N_20306);
and U32956 (N_32956,N_27727,N_22525);
nand U32957 (N_32957,N_21947,N_20082);
nand U32958 (N_32958,N_25434,N_26677);
xor U32959 (N_32959,N_21567,N_20327);
and U32960 (N_32960,N_23691,N_28918);
nand U32961 (N_32961,N_29924,N_24837);
nor U32962 (N_32962,N_20924,N_20028);
nand U32963 (N_32963,N_23333,N_21202);
and U32964 (N_32964,N_22963,N_27713);
and U32965 (N_32965,N_20622,N_26461);
and U32966 (N_32966,N_28754,N_28317);
and U32967 (N_32967,N_21001,N_25595);
nand U32968 (N_32968,N_24505,N_20118);
and U32969 (N_32969,N_23762,N_20813);
nand U32970 (N_32970,N_29784,N_21193);
and U32971 (N_32971,N_20411,N_20162);
nor U32972 (N_32972,N_26279,N_21807);
and U32973 (N_32973,N_26008,N_22993);
nor U32974 (N_32974,N_23562,N_20108);
nand U32975 (N_32975,N_28816,N_22328);
and U32976 (N_32976,N_27577,N_29224);
nor U32977 (N_32977,N_23665,N_27311);
nor U32978 (N_32978,N_25104,N_27832);
or U32979 (N_32979,N_26786,N_25929);
nand U32980 (N_32980,N_27884,N_26446);
and U32981 (N_32981,N_29236,N_20584);
nand U32982 (N_32982,N_23453,N_22200);
and U32983 (N_32983,N_21021,N_24171);
nor U32984 (N_32984,N_22705,N_27933);
nand U32985 (N_32985,N_29234,N_25399);
nand U32986 (N_32986,N_23438,N_28440);
nor U32987 (N_32987,N_27481,N_27861);
or U32988 (N_32988,N_27956,N_20765);
xnor U32989 (N_32989,N_20448,N_27202);
nand U32990 (N_32990,N_20398,N_28062);
nand U32991 (N_32991,N_26433,N_20888);
and U32992 (N_32992,N_21721,N_26510);
nor U32993 (N_32993,N_21569,N_27915);
nand U32994 (N_32994,N_23113,N_21495);
and U32995 (N_32995,N_29278,N_21498);
nor U32996 (N_32996,N_27263,N_24157);
xor U32997 (N_32997,N_25768,N_22692);
nand U32998 (N_32998,N_29642,N_21224);
xnor U32999 (N_32999,N_24350,N_26047);
xor U33000 (N_33000,N_24305,N_25955);
and U33001 (N_33001,N_22480,N_24584);
nand U33002 (N_33002,N_20994,N_26946);
and U33003 (N_33003,N_26325,N_23662);
nand U33004 (N_33004,N_25216,N_27734);
nand U33005 (N_33005,N_29275,N_24121);
xnor U33006 (N_33006,N_20811,N_20149);
xnor U33007 (N_33007,N_29902,N_27433);
and U33008 (N_33008,N_23705,N_25471);
nand U33009 (N_33009,N_29425,N_27818);
and U33010 (N_33010,N_20184,N_24163);
or U33011 (N_33011,N_27679,N_28354);
xnor U33012 (N_33012,N_22438,N_22076);
nor U33013 (N_33013,N_21900,N_26425);
nand U33014 (N_33014,N_22317,N_27716);
or U33015 (N_33015,N_26119,N_29277);
nand U33016 (N_33016,N_24127,N_28854);
xnor U33017 (N_33017,N_21445,N_29283);
nand U33018 (N_33018,N_24175,N_26414);
and U33019 (N_33019,N_25947,N_23703);
and U33020 (N_33020,N_22135,N_27744);
nor U33021 (N_33021,N_20261,N_27591);
nor U33022 (N_33022,N_26832,N_26559);
nand U33023 (N_33023,N_29793,N_28264);
nand U33024 (N_33024,N_29654,N_22775);
nand U33025 (N_33025,N_27392,N_22976);
xnor U33026 (N_33026,N_21515,N_25582);
nor U33027 (N_33027,N_27438,N_20392);
or U33028 (N_33028,N_24871,N_23140);
nor U33029 (N_33029,N_23832,N_26317);
xor U33030 (N_33030,N_21737,N_27241);
xnor U33031 (N_33031,N_27619,N_25678);
and U33032 (N_33032,N_28318,N_26612);
and U33033 (N_33033,N_23388,N_29220);
nor U33034 (N_33034,N_26144,N_24097);
nand U33035 (N_33035,N_28031,N_26685);
nand U33036 (N_33036,N_26775,N_23143);
xnor U33037 (N_33037,N_24773,N_21653);
nor U33038 (N_33038,N_21086,N_28423);
or U33039 (N_33039,N_25608,N_23934);
or U33040 (N_33040,N_25190,N_21367);
and U33041 (N_33041,N_20975,N_23967);
and U33042 (N_33042,N_29912,N_23318);
or U33043 (N_33043,N_23407,N_29769);
and U33044 (N_33044,N_20191,N_21811);
and U33045 (N_33045,N_27189,N_20013);
and U33046 (N_33046,N_23723,N_27271);
and U33047 (N_33047,N_23295,N_28902);
nor U33048 (N_33048,N_24179,N_22548);
and U33049 (N_33049,N_23029,N_21004);
xnor U33050 (N_33050,N_23150,N_23853);
nand U33051 (N_33051,N_24831,N_24371);
and U33052 (N_33052,N_25806,N_23796);
nand U33053 (N_33053,N_28574,N_23118);
xnor U33054 (N_33054,N_27176,N_25653);
or U33055 (N_33055,N_26083,N_24053);
nor U33056 (N_33056,N_28174,N_24035);
nor U33057 (N_33057,N_27580,N_28112);
or U33058 (N_33058,N_26064,N_20419);
nor U33059 (N_33059,N_21554,N_23432);
xnor U33060 (N_33060,N_26442,N_26007);
nand U33061 (N_33061,N_29763,N_29119);
or U33062 (N_33062,N_20758,N_25497);
or U33063 (N_33063,N_20007,N_24439);
and U33064 (N_33064,N_26889,N_29377);
nor U33065 (N_33065,N_25630,N_20798);
xnor U33066 (N_33066,N_21123,N_28837);
nand U33067 (N_33067,N_22917,N_24676);
nand U33068 (N_33068,N_21065,N_23569);
nand U33069 (N_33069,N_26596,N_20378);
or U33070 (N_33070,N_24297,N_22253);
or U33071 (N_33071,N_23519,N_21003);
and U33072 (N_33072,N_20089,N_23539);
nand U33073 (N_33073,N_23931,N_20430);
xor U33074 (N_33074,N_20529,N_25749);
nor U33075 (N_33075,N_28203,N_28860);
nor U33076 (N_33076,N_26188,N_27867);
or U33077 (N_33077,N_25751,N_25638);
nor U33078 (N_33078,N_29212,N_29150);
xor U33079 (N_33079,N_20248,N_23337);
or U33080 (N_33080,N_29962,N_22305);
xnor U33081 (N_33081,N_22606,N_28804);
nor U33082 (N_33082,N_28338,N_20251);
or U33083 (N_33083,N_25077,N_20656);
and U33084 (N_33084,N_23146,N_29319);
nand U33085 (N_33085,N_26599,N_23227);
nand U33086 (N_33086,N_23530,N_26984);
and U33087 (N_33087,N_22689,N_23142);
nor U33088 (N_33088,N_22124,N_25225);
xnor U33089 (N_33089,N_29329,N_29134);
xor U33090 (N_33090,N_28643,N_24635);
nor U33091 (N_33091,N_22806,N_27332);
nand U33092 (N_33092,N_23940,N_21060);
and U33093 (N_33093,N_29148,N_27276);
nand U33094 (N_33094,N_25837,N_22212);
nand U33095 (N_33095,N_27169,N_20803);
nand U33096 (N_33096,N_26382,N_22936);
or U33097 (N_33097,N_28430,N_23645);
xnor U33098 (N_33098,N_29176,N_28396);
nand U33099 (N_33099,N_22576,N_23756);
xor U33100 (N_33100,N_27976,N_20606);
nand U33101 (N_33101,N_24806,N_23871);
xnor U33102 (N_33102,N_20231,N_29455);
and U33103 (N_33103,N_26611,N_21113);
nor U33104 (N_33104,N_23708,N_24503);
xor U33105 (N_33105,N_24212,N_25993);
and U33106 (N_33106,N_26815,N_27180);
and U33107 (N_33107,N_21219,N_26099);
and U33108 (N_33108,N_28154,N_28724);
nor U33109 (N_33109,N_22916,N_23244);
xnor U33110 (N_33110,N_26250,N_20727);
or U33111 (N_33111,N_21512,N_22528);
nand U33112 (N_33112,N_29247,N_23655);
nor U33113 (N_33113,N_26508,N_20245);
and U33114 (N_33114,N_27317,N_27348);
nand U33115 (N_33115,N_27946,N_23274);
nor U33116 (N_33116,N_25783,N_22410);
nor U33117 (N_33117,N_27309,N_24438);
and U33118 (N_33118,N_22550,N_28980);
nand U33119 (N_33119,N_24335,N_21329);
xnor U33120 (N_33120,N_25060,N_27298);
and U33121 (N_33121,N_22418,N_26784);
and U33122 (N_33122,N_27573,N_21209);
and U33123 (N_33123,N_29404,N_23442);
nor U33124 (N_33124,N_26324,N_24132);
nand U33125 (N_33125,N_27715,N_22096);
and U33126 (N_33126,N_24359,N_24655);
nor U33127 (N_33127,N_21598,N_29331);
or U33128 (N_33128,N_28379,N_24544);
xnor U33129 (N_33129,N_23611,N_20603);
nor U33130 (N_33130,N_22041,N_28326);
nand U33131 (N_33131,N_20959,N_29036);
or U33132 (N_33132,N_24442,N_27102);
nor U33133 (N_33133,N_25812,N_29479);
xor U33134 (N_33134,N_23350,N_21234);
and U33135 (N_33135,N_26084,N_27940);
nand U33136 (N_33136,N_25862,N_29637);
or U33137 (N_33137,N_21246,N_24533);
nand U33138 (N_33138,N_28475,N_26679);
or U33139 (N_33139,N_27054,N_29893);
or U33140 (N_33140,N_26153,N_21664);
nand U33141 (N_33141,N_26605,N_25803);
and U33142 (N_33142,N_22290,N_23022);
xnor U33143 (N_33143,N_29440,N_24521);
nand U33144 (N_33144,N_22082,N_24781);
nand U33145 (N_33145,N_26980,N_26540);
or U33146 (N_33146,N_22898,N_20607);
nor U33147 (N_33147,N_27644,N_23700);
or U33148 (N_33148,N_21332,N_21030);
and U33149 (N_33149,N_27452,N_25957);
nor U33150 (N_33150,N_24700,N_23294);
nor U33151 (N_33151,N_28977,N_20424);
nand U33152 (N_33152,N_27949,N_20579);
nand U33153 (N_33153,N_23922,N_25855);
nand U33154 (N_33154,N_28362,N_26803);
or U33155 (N_33155,N_27617,N_22812);
or U33156 (N_33156,N_28287,N_24332);
nand U33157 (N_33157,N_28464,N_25332);
and U33158 (N_33158,N_28762,N_28859);
or U33159 (N_33159,N_25275,N_28818);
xor U33160 (N_33160,N_20620,N_20292);
nand U33161 (N_33161,N_28375,N_25439);
xnor U33162 (N_33162,N_26659,N_25624);
and U33163 (N_33163,N_27677,N_20199);
xor U33164 (N_33164,N_22577,N_23293);
and U33165 (N_33165,N_22613,N_24839);
and U33166 (N_33166,N_22944,N_26947);
and U33167 (N_33167,N_25779,N_22639);
nor U33168 (N_33168,N_24250,N_26742);
or U33169 (N_33169,N_23465,N_26041);
xor U33170 (N_33170,N_26761,N_25910);
and U33171 (N_33171,N_26897,N_22312);
nand U33172 (N_33172,N_22229,N_29476);
nor U33173 (N_33173,N_20709,N_23506);
and U33174 (N_33174,N_26184,N_25835);
nor U33175 (N_33175,N_26124,N_27424);
xnor U33176 (N_33176,N_26576,N_28815);
nand U33177 (N_33177,N_20794,N_22906);
nand U33178 (N_33178,N_26629,N_26782);
nand U33179 (N_33179,N_21912,N_21229);
or U33180 (N_33180,N_22522,N_20195);
or U33181 (N_33181,N_26880,N_25308);
and U33182 (N_33182,N_23768,N_20190);
nand U33183 (N_33183,N_27751,N_28433);
or U33184 (N_33184,N_22913,N_20364);
xnor U33185 (N_33185,N_29473,N_29276);
nor U33186 (N_33186,N_26828,N_21356);
or U33187 (N_33187,N_27229,N_27408);
xnor U33188 (N_33188,N_22733,N_24155);
and U33189 (N_33189,N_29233,N_24986);
xor U33190 (N_33190,N_22357,N_26322);
xnor U33191 (N_33191,N_23624,N_24217);
xor U33192 (N_33192,N_20925,N_29363);
xor U33193 (N_33193,N_25883,N_25298);
or U33194 (N_33194,N_23387,N_24500);
nor U33195 (N_33195,N_20322,N_21756);
nand U33196 (N_33196,N_24028,N_28490);
or U33197 (N_33197,N_25027,N_21059);
nor U33198 (N_33198,N_22751,N_28884);
nor U33199 (N_33199,N_20716,N_25848);
nor U33200 (N_33200,N_23073,N_21369);
xor U33201 (N_33201,N_23822,N_29762);
xor U33202 (N_33202,N_25006,N_21924);
and U33203 (N_33203,N_28681,N_28080);
or U33204 (N_33204,N_24174,N_21276);
nand U33205 (N_33205,N_20492,N_21725);
xnor U33206 (N_33206,N_23584,N_22501);
nor U33207 (N_33207,N_26702,N_24111);
nor U33208 (N_33208,N_22995,N_21210);
nor U33209 (N_33209,N_29710,N_28786);
nand U33210 (N_33210,N_27869,N_28184);
nor U33211 (N_33211,N_24334,N_27206);
and U33212 (N_33212,N_20903,N_21110);
xnor U33213 (N_33213,N_24862,N_27395);
or U33214 (N_33214,N_21975,N_21399);
or U33215 (N_33215,N_22000,N_20970);
xnor U33216 (N_33216,N_26616,N_27592);
and U33217 (N_33217,N_24226,N_24836);
nor U33218 (N_33218,N_22183,N_20828);
or U33219 (N_33219,N_22095,N_29905);
and U33220 (N_33220,N_24280,N_23698);
nand U33221 (N_33221,N_22454,N_25360);
nand U33222 (N_33222,N_25405,N_24934);
nor U33223 (N_33223,N_24417,N_21205);
or U33224 (N_33224,N_25851,N_21998);
nor U33225 (N_33225,N_20940,N_26886);
nand U33226 (N_33226,N_23695,N_22117);
and U33227 (N_33227,N_27184,N_21389);
or U33228 (N_33228,N_23894,N_27563);
or U33229 (N_33229,N_23809,N_29271);
nor U33230 (N_33230,N_24465,N_28586);
nand U33231 (N_33231,N_20414,N_20218);
or U33232 (N_33232,N_28507,N_20019);
or U33233 (N_33233,N_29030,N_27966);
nor U33234 (N_33234,N_24845,N_23959);
nor U33235 (N_33235,N_24341,N_24116);
nor U33236 (N_33236,N_27864,N_29062);
or U33237 (N_33237,N_21159,N_29215);
xor U33238 (N_33238,N_26570,N_20109);
xor U33239 (N_33239,N_27703,N_22727);
xnor U33240 (N_33240,N_24966,N_26078);
or U33241 (N_33241,N_20265,N_28089);
xor U33242 (N_33242,N_28305,N_22774);
nand U33243 (N_33243,N_21727,N_26662);
xnor U33244 (N_33244,N_29604,N_28670);
nor U33245 (N_33245,N_28951,N_29796);
nor U33246 (N_33246,N_28495,N_20186);
or U33247 (N_33247,N_23631,N_24378);
or U33248 (N_33248,N_23627,N_22541);
and U33249 (N_33249,N_20816,N_26519);
nor U33250 (N_33250,N_29936,N_27972);
nor U33251 (N_33251,N_27361,N_29499);
or U33252 (N_33252,N_23176,N_22973);
and U33253 (N_33253,N_29322,N_21988);
nand U33254 (N_33254,N_24105,N_20886);
nor U33255 (N_33255,N_28374,N_20080);
nor U33256 (N_33256,N_22447,N_29197);
and U33257 (N_33257,N_25457,N_24829);
or U33258 (N_33258,N_29879,N_20117);
and U33259 (N_33259,N_21133,N_29005);
or U33260 (N_33260,N_21616,N_26530);
or U33261 (N_33261,N_25335,N_24668);
nand U33262 (N_33262,N_29775,N_20472);
nand U33263 (N_33263,N_27069,N_29052);
and U33264 (N_33264,N_28232,N_20678);
or U33265 (N_33265,N_28099,N_25260);
nor U33266 (N_33266,N_23371,N_29860);
nand U33267 (N_33267,N_25548,N_28558);
nor U33268 (N_33268,N_21023,N_21078);
nor U33269 (N_33269,N_26982,N_27003);
nor U33270 (N_33270,N_23716,N_21101);
nor U33271 (N_33271,N_22584,N_26025);
nor U33272 (N_33272,N_27654,N_27346);
or U33273 (N_33273,N_27607,N_24878);
xnor U33274 (N_33274,N_22743,N_21564);
xnor U33275 (N_33275,N_25948,N_23443);
nand U33276 (N_33276,N_25818,N_28864);
or U33277 (N_33277,N_22199,N_27280);
xnor U33278 (N_33278,N_26554,N_24610);
xor U33279 (N_33279,N_28369,N_26254);
xnor U33280 (N_33280,N_23254,N_20066);
xor U33281 (N_33281,N_24637,N_25515);
and U33282 (N_33282,N_24093,N_23399);
or U33283 (N_33283,N_28888,N_28029);
xor U33284 (N_33284,N_27848,N_26410);
and U33285 (N_33285,N_21089,N_27647);
nand U33286 (N_33286,N_25850,N_20115);
or U33287 (N_33287,N_24402,N_21692);
nand U33288 (N_33288,N_28794,N_21593);
xnor U33289 (N_33289,N_29253,N_26793);
nand U33290 (N_33290,N_29536,N_23522);
or U33291 (N_33291,N_24041,N_20343);
or U33292 (N_33292,N_29740,N_20463);
or U33293 (N_33293,N_29805,N_28699);
xnor U33294 (N_33294,N_27145,N_25535);
nor U33295 (N_33295,N_25709,N_21827);
nand U33296 (N_33296,N_25396,N_25408);
nor U33297 (N_33297,N_29658,N_20325);
or U33298 (N_33298,N_23000,N_27393);
and U33299 (N_33299,N_23837,N_23709);
and U33300 (N_33300,N_24065,N_20361);
and U33301 (N_33301,N_20467,N_28861);
nor U33302 (N_33302,N_22158,N_23221);
xnor U33303 (N_33303,N_20001,N_25687);
and U33304 (N_33304,N_25226,N_26904);
and U33305 (N_33305,N_26777,N_24581);
xnor U33306 (N_33306,N_22592,N_26938);
or U33307 (N_33307,N_27999,N_27638);
nand U33308 (N_33308,N_25316,N_25379);
nand U33309 (N_33309,N_23964,N_24802);
nor U33310 (N_33310,N_23881,N_29869);
nand U33311 (N_33311,N_26706,N_29556);
xnor U33312 (N_33312,N_22680,N_25280);
or U33313 (N_33313,N_27771,N_26336);
xor U33314 (N_33314,N_27441,N_26907);
xnor U33315 (N_33315,N_20641,N_20839);
and U33316 (N_33316,N_28187,N_25117);
nor U33317 (N_33317,N_24892,N_25959);
nor U33318 (N_33318,N_21795,N_22985);
or U33319 (N_33319,N_20917,N_28470);
or U33320 (N_33320,N_29105,N_27833);
xnor U33321 (N_33321,N_26238,N_27255);
and U33322 (N_33322,N_22921,N_28795);
nand U33323 (N_33323,N_22882,N_21353);
nand U33324 (N_33324,N_23347,N_25041);
and U33325 (N_33325,N_29038,N_26568);
nand U33326 (N_33326,N_25350,N_29021);
or U33327 (N_33327,N_21465,N_24669);
or U33328 (N_33328,N_29082,N_23024);
or U33329 (N_33329,N_26231,N_22504);
xor U33330 (N_33330,N_25358,N_23536);
or U33331 (N_33331,N_23331,N_22003);
or U33332 (N_33332,N_26840,N_21505);
nand U33333 (N_33333,N_22838,N_23783);
nand U33334 (N_33334,N_29028,N_22758);
and U33335 (N_33335,N_21165,N_24370);
or U33336 (N_33336,N_24790,N_22308);
nor U33337 (N_33337,N_24101,N_25777);
nand U33338 (N_33338,N_22267,N_29048);
and U33339 (N_33339,N_28224,N_25293);
and U33340 (N_33340,N_27007,N_28525);
nor U33341 (N_33341,N_29632,N_20236);
nand U33342 (N_33342,N_28469,N_26979);
or U33343 (N_33343,N_23817,N_26126);
xor U33344 (N_33344,N_24691,N_23517);
and U33345 (N_33345,N_27353,N_22489);
or U33346 (N_33346,N_20670,N_27335);
nor U33347 (N_33347,N_23893,N_23989);
nand U33348 (N_33348,N_24192,N_21152);
nor U33349 (N_33349,N_23058,N_28095);
nand U33350 (N_33350,N_24275,N_23540);
or U33351 (N_33351,N_28839,N_23189);
nor U33352 (N_33352,N_25409,N_28651);
or U33353 (N_33353,N_21252,N_25005);
and U33354 (N_33354,N_23340,N_27612);
nand U33355 (N_33355,N_25374,N_25951);
nor U33356 (N_33356,N_29509,N_28568);
or U33357 (N_33357,N_24273,N_26459);
nor U33358 (N_33358,N_24466,N_26376);
nand U33359 (N_33359,N_26709,N_22344);
nand U33360 (N_33360,N_21903,N_21286);
and U33361 (N_33361,N_20757,N_26933);
and U33362 (N_33362,N_28813,N_29463);
or U33363 (N_33363,N_23586,N_27297);
or U33364 (N_33364,N_29358,N_23490);
xor U33365 (N_33365,N_20146,N_28078);
xnor U33366 (N_33366,N_25013,N_23825);
nor U33367 (N_33367,N_26105,N_28295);
or U33368 (N_33368,N_22823,N_29738);
nand U33369 (N_33369,N_26526,N_20152);
nor U33370 (N_33370,N_26613,N_26368);
nor U33371 (N_33371,N_27172,N_25572);
nand U33372 (N_33372,N_24627,N_25897);
and U33373 (N_33373,N_26877,N_24063);
and U33374 (N_33374,N_29355,N_21095);
or U33375 (N_33375,N_23344,N_22180);
and U33376 (N_33376,N_23171,N_24369);
nand U33377 (N_33377,N_26887,N_29906);
xor U33378 (N_33378,N_23991,N_27702);
and U33379 (N_33379,N_21520,N_21925);
or U33380 (N_33380,N_25781,N_29672);
nand U33381 (N_33381,N_24406,N_27602);
nand U33382 (N_33382,N_28512,N_25091);
xnor U33383 (N_33383,N_27522,N_26441);
or U33384 (N_33384,N_21915,N_28351);
or U33385 (N_33385,N_21856,N_28905);
nor U33386 (N_33386,N_27981,N_27786);
nor U33387 (N_33387,N_24815,N_20846);
nand U33388 (N_33388,N_27698,N_28162);
xor U33389 (N_33389,N_29707,N_20613);
and U33390 (N_33390,N_28458,N_29330);
nor U33391 (N_33391,N_21553,N_24685);
xnor U33392 (N_33392,N_21873,N_21672);
nor U33393 (N_33393,N_28097,N_29114);
nand U33394 (N_33394,N_28373,N_27555);
and U33395 (N_33395,N_28976,N_20012);
nor U33396 (N_33396,N_29218,N_24074);
nand U33397 (N_33397,N_24022,N_23089);
nor U33398 (N_33398,N_28143,N_20316);
or U33399 (N_33399,N_24721,N_27103);
nor U33400 (N_33400,N_29564,N_21614);
and U33401 (N_33401,N_21559,N_26052);
nand U33402 (N_33402,N_27489,N_26972);
nand U33403 (N_33403,N_27561,N_28386);
nor U33404 (N_33404,N_28119,N_28552);
nor U33405 (N_33405,N_29865,N_21954);
or U33406 (N_33406,N_21754,N_22416);
nor U33407 (N_33407,N_28422,N_28767);
or U33408 (N_33408,N_24988,N_26245);
nor U33409 (N_33409,N_25333,N_28547);
or U33410 (N_33410,N_24958,N_22722);
and U33411 (N_33411,N_22950,N_29126);
or U33412 (N_33412,N_25895,N_21299);
xor U33413 (N_33413,N_29633,N_21893);
or U33414 (N_33414,N_22523,N_26117);
xor U33415 (N_33415,N_27925,N_29378);
nand U33416 (N_33416,N_22303,N_26546);
or U33417 (N_33417,N_27882,N_29087);
or U33418 (N_33418,N_29935,N_22941);
nor U33419 (N_33419,N_24104,N_28182);
xor U33420 (N_33420,N_20143,N_20335);
and U33421 (N_33421,N_21871,N_27415);
nand U33422 (N_33422,N_28933,N_21709);
or U33423 (N_33423,N_20078,N_28617);
nand U33424 (N_33424,N_21346,N_23356);
nor U33425 (N_33425,N_22757,N_25259);
nor U33426 (N_33426,N_24929,N_28996);
and U33427 (N_33427,N_20666,N_25098);
nand U33428 (N_33428,N_24476,N_23710);
or U33429 (N_33429,N_28949,N_25130);
and U33430 (N_33430,N_23602,N_22488);
nor U33431 (N_33431,N_29205,N_29008);
xnor U33432 (N_33432,N_23898,N_22019);
nand U33433 (N_33433,N_24603,N_27960);
xnor U33434 (N_33434,N_20669,N_26225);
and U33435 (N_33435,N_25575,N_27750);
nor U33436 (N_33436,N_21572,N_26983);
nand U33437 (N_33437,N_22220,N_29412);
xor U33438 (N_33438,N_22237,N_27970);
or U33439 (N_33439,N_29976,N_26038);
or U33440 (N_33440,N_22236,N_24876);
xor U33441 (N_33441,N_22795,N_20596);
or U33442 (N_33442,N_24918,N_25567);
xor U33443 (N_33443,N_29946,N_25625);
xnor U33444 (N_33444,N_29269,N_26913);
nand U33445 (N_33445,N_23312,N_23577);
or U33446 (N_33446,N_21775,N_25051);
or U33447 (N_33447,N_24358,N_29795);
or U33448 (N_33448,N_20836,N_20766);
nor U33449 (N_33449,N_21080,N_28755);
or U33450 (N_33450,N_21304,N_26481);
nand U33451 (N_33451,N_26043,N_22870);
nor U33452 (N_33452,N_28027,N_28009);
nand U33453 (N_33453,N_28105,N_23279);
and U33454 (N_33454,N_28335,N_29066);
nand U33455 (N_33455,N_28523,N_27400);
nor U33456 (N_33456,N_21696,N_28777);
nand U33457 (N_33457,N_21898,N_22072);
and U33458 (N_33458,N_22255,N_20614);
nand U33459 (N_33459,N_29582,N_28077);
nor U33460 (N_33460,N_23193,N_20887);
and U33461 (N_33461,N_24218,N_20483);
and U33462 (N_33462,N_20081,N_24771);
or U33463 (N_33463,N_28081,N_21841);
or U33464 (N_33464,N_28778,N_23963);
nor U33465 (N_33465,N_28429,N_26598);
or U33466 (N_33466,N_24258,N_26402);
and U33467 (N_33467,N_23373,N_21840);
xnor U33468 (N_33468,N_23565,N_24670);
nand U33469 (N_33469,N_28482,N_29683);
and U33470 (N_33470,N_21049,N_22785);
nor U33471 (N_33471,N_25394,N_24532);
nor U33472 (N_33472,N_25834,N_27039);
or U33473 (N_33473,N_24619,N_27275);
nor U33474 (N_33474,N_25043,N_26998);
or U33475 (N_33475,N_20815,N_25971);
and U33476 (N_33476,N_25900,N_20842);
xor U33477 (N_33477,N_24207,N_25703);
or U33478 (N_33478,N_26201,N_20500);
and U33479 (N_33479,N_28867,N_24943);
xnor U33480 (N_33480,N_28865,N_27620);
or U33481 (N_33481,N_26372,N_23101);
nand U33482 (N_33482,N_20617,N_29475);
and U33483 (N_33483,N_27731,N_21254);
xnor U33484 (N_33484,N_24726,N_26290);
nand U33485 (N_33485,N_23097,N_27942);
nor U33486 (N_33486,N_27876,N_20550);
and U33487 (N_33487,N_21137,N_22167);
xnor U33488 (N_33488,N_20031,N_20555);
nor U33489 (N_33489,N_23771,N_29470);
or U33490 (N_33490,N_23471,N_26359);
and U33491 (N_33491,N_26304,N_29348);
xor U33492 (N_33492,N_24542,N_25251);
nor U33493 (N_33493,N_25511,N_20215);
or U33494 (N_33494,N_28313,N_29989);
or U33495 (N_33495,N_22716,N_25351);
xor U33496 (N_33496,N_24185,N_20879);
nand U33497 (N_33497,N_22088,N_23204);
xnor U33498 (N_33498,N_28171,N_27014);
nand U33499 (N_33499,N_24546,N_27538);
or U33500 (N_33500,N_28026,N_25467);
and U33501 (N_33501,N_22764,N_25707);
xnor U33502 (N_33502,N_22905,N_22580);
xor U33503 (N_33503,N_22241,N_21847);
and U33504 (N_33504,N_21801,N_25868);
nor U33505 (N_33505,N_21722,N_21432);
nand U33506 (N_33506,N_24517,N_23127);
or U33507 (N_33507,N_23010,N_24117);
and U33508 (N_33508,N_26906,N_22444);
nor U33509 (N_33509,N_26626,N_28016);
and U33510 (N_33510,N_24650,N_25577);
xor U33511 (N_33511,N_28110,N_21523);
or U33512 (N_33512,N_20442,N_29995);
and U33513 (N_33513,N_25759,N_26766);
nor U33514 (N_33514,N_28432,N_27100);
nor U33515 (N_33515,N_24082,N_23676);
nor U33516 (N_33516,N_29060,N_26218);
and U33517 (N_33517,N_25532,N_25667);
xnor U33518 (N_33518,N_20914,N_27207);
or U33519 (N_33519,N_29513,N_24618);
nand U33520 (N_33520,N_27090,N_21260);
nand U33521 (N_33521,N_24498,N_20193);
xnor U33522 (N_33522,N_29668,N_29203);
or U33523 (N_33523,N_21241,N_25205);
or U33524 (N_33524,N_25208,N_26562);
and U33525 (N_33525,N_23632,N_21790);
xnor U33526 (N_33526,N_24677,N_29175);
or U33527 (N_33527,N_25465,N_27474);
xor U33528 (N_33528,N_26031,N_23084);
or U33529 (N_33529,N_28704,N_25029);
xnor U33530 (N_33530,N_22252,N_20761);
nand U33531 (N_33531,N_22546,N_20341);
nor U33532 (N_33532,N_27055,N_21396);
xnor U33533 (N_33533,N_20240,N_25038);
nand U33534 (N_33534,N_25124,N_24612);
xor U33535 (N_33535,N_21537,N_22002);
nand U33536 (N_33536,N_22261,N_22294);
nand U33537 (N_33537,N_24573,N_21400);
xnor U33538 (N_33538,N_21020,N_20895);
or U33539 (N_33539,N_29735,N_24278);
nor U33540 (N_33540,N_24911,N_24336);
nand U33541 (N_33541,N_23867,N_22808);
or U33542 (N_33542,N_25564,N_24286);
nor U33543 (N_33543,N_23601,N_29948);
xnor U33544 (N_33544,N_24772,N_22207);
and U33545 (N_33545,N_23612,N_24923);
nand U33546 (N_33546,N_25097,N_21693);
and U33547 (N_33547,N_21387,N_20026);
nand U33548 (N_33548,N_25056,N_22484);
or U33549 (N_33549,N_22329,N_22886);
xnor U33550 (N_33550,N_23915,N_29636);
or U33551 (N_33551,N_29894,N_20773);
and U33552 (N_33552,N_29777,N_29449);
and U33553 (N_33553,N_28510,N_28748);
or U33554 (N_33554,N_24638,N_23754);
xor U33555 (N_33555,N_27586,N_28652);
nand U33556 (N_33556,N_20863,N_25288);
nor U33557 (N_33557,N_27000,N_26801);
xnor U33558 (N_33558,N_23920,N_22455);
or U33559 (N_33559,N_28528,N_21724);
nor U33560 (N_33560,N_22643,N_26739);
nor U33561 (N_33561,N_24556,N_29725);
xnor U33562 (N_33562,N_26159,N_28066);
or U33563 (N_33563,N_22824,N_24950);
nor U33564 (N_33564,N_21532,N_27063);
xnor U33565 (N_33565,N_22790,N_25652);
or U33566 (N_33566,N_26206,N_27521);
and U33567 (N_33567,N_29299,N_27846);
or U33568 (N_33568,N_28161,N_28205);
or U33569 (N_33569,N_29057,N_26431);
xor U33570 (N_33570,N_28133,N_28042);
or U33571 (N_33571,N_23977,N_25810);
or U33572 (N_33572,N_29998,N_23026);
and U33573 (N_33573,N_22666,N_28248);
xnor U33574 (N_33574,N_23250,N_24812);
and U33575 (N_33575,N_26329,N_25927);
nand U33576 (N_33576,N_29840,N_27388);
nand U33577 (N_33577,N_23637,N_25522);
nor U33578 (N_33578,N_28743,N_27811);
nor U33579 (N_33579,N_28910,N_21331);
xnor U33580 (N_33580,N_25184,N_24821);
nor U33581 (N_33581,N_21778,N_22841);
and U33582 (N_33582,N_22140,N_22053);
or U33583 (N_33583,N_26847,N_26095);
and U33584 (N_33584,N_27674,N_28253);
nand U33585 (N_33585,N_26092,N_26830);
nand U33586 (N_33586,N_24684,N_24066);
or U33587 (N_33587,N_23280,N_28149);
xnor U33588 (N_33588,N_27221,N_27334);
xor U33589 (N_33589,N_29490,N_28049);
xnor U33590 (N_33590,N_20673,N_29024);
nor U33591 (N_33591,N_26357,N_21129);
xor U33592 (N_33592,N_27977,N_24909);
and U33593 (N_33593,N_22593,N_22789);
xnor U33594 (N_33594,N_24394,N_23427);
or U33595 (N_33595,N_24689,N_27666);
xor U33596 (N_33596,N_29665,N_25324);
nor U33597 (N_33597,N_28056,N_27508);
or U33598 (N_33598,N_20960,N_23315);
or U33599 (N_33599,N_27542,N_25477);
xor U33600 (N_33600,N_26707,N_22877);
xnor U33601 (N_33601,N_24930,N_22333);
or U33602 (N_33602,N_24783,N_27131);
xor U33603 (N_33603,N_24717,N_26331);
xnor U33604 (N_33604,N_22054,N_24632);
and U33605 (N_33605,N_26136,N_20189);
nor U33606 (N_33606,N_27075,N_20480);
or U33607 (N_33607,N_25539,N_25753);
nor U33608 (N_33608,N_25419,N_21618);
or U33609 (N_33609,N_26653,N_21634);
or U33610 (N_33610,N_27002,N_24495);
and U33611 (N_33611,N_28707,N_25470);
nor U33612 (N_33612,N_26986,N_29765);
or U33613 (N_33613,N_26622,N_26551);
nor U33614 (N_33614,N_24037,N_26230);
xor U33615 (N_33615,N_29964,N_25490);
nand U33616 (N_33616,N_21689,N_26749);
nor U33617 (N_33617,N_23564,N_22549);
nand U33618 (N_33618,N_27267,N_21497);
nand U33619 (N_33619,N_21204,N_28034);
xnor U33620 (N_33620,N_26158,N_27414);
and U33621 (N_33621,N_26624,N_23200);
xor U33622 (N_33622,N_20037,N_23362);
or U33623 (N_33623,N_23807,N_23242);
or U33624 (N_33624,N_27720,N_28984);
and U33625 (N_33625,N_28044,N_23697);
or U33626 (N_33626,N_28889,N_28862);
and U33627 (N_33627,N_20616,N_29904);
and U33628 (N_33628,N_24624,N_21605);
nor U33629 (N_33629,N_25050,N_23057);
xor U33630 (N_33630,N_29462,N_20170);
nor U33631 (N_33631,N_27512,N_28666);
nand U33632 (N_33632,N_21002,N_25362);
and U33633 (N_33633,N_21688,N_29282);
xor U33634 (N_33634,N_22040,N_21500);
xor U33635 (N_33635,N_29006,N_21509);
or U33636 (N_33636,N_26955,N_23613);
and U33637 (N_33637,N_28769,N_22087);
nor U33638 (N_33638,N_22776,N_29128);
xor U33639 (N_33639,N_24990,N_23734);
nand U33640 (N_33640,N_20820,N_21311);
or U33641 (N_33641,N_24338,N_29200);
nand U33642 (N_33642,N_28141,N_28472);
xnor U33643 (N_33643,N_22677,N_28461);
or U33644 (N_33644,N_29798,N_23410);
or U33645 (N_33645,N_23932,N_20972);
nand U33646 (N_33646,N_28215,N_21720);
nor U33647 (N_33647,N_23233,N_28921);
nand U33648 (N_33648,N_20552,N_26194);
nand U33649 (N_33649,N_22910,N_23489);
nand U33650 (N_33650,N_22583,N_23338);
nand U33651 (N_33651,N_29867,N_20721);
xnor U33652 (N_33652,N_21291,N_29389);
and U33653 (N_33653,N_29372,N_26969);
and U33654 (N_33654,N_25989,N_28689);
nand U33655 (N_33655,N_22370,N_24184);
or U33656 (N_33656,N_29851,N_23236);
nor U33657 (N_33657,N_27037,N_21989);
nand U33658 (N_33658,N_28088,N_20629);
or U33659 (N_33659,N_29934,N_21146);
nand U33660 (N_33660,N_25199,N_22736);
nor U33661 (N_33661,N_21151,N_20403);
nand U33662 (N_33662,N_20114,N_26299);
nor U33663 (N_33663,N_20788,N_28117);
or U33664 (N_33664,N_27585,N_22085);
nor U33665 (N_33665,N_28983,N_29533);
xnor U33666 (N_33666,N_25514,N_22107);
xnor U33667 (N_33667,N_25675,N_21117);
xor U33668 (N_33668,N_25137,N_29464);
and U33669 (N_33669,N_25857,N_28068);
xnor U33670 (N_33670,N_28275,N_21256);
or U33671 (N_33671,N_21300,N_29776);
nand U33672 (N_33672,N_21872,N_20829);
or U33673 (N_33673,N_24489,N_24384);
xor U33674 (N_33674,N_20127,N_24984);
and U33675 (N_33675,N_23199,N_23299);
xor U33676 (N_33676,N_27789,N_27423);
nor U33677 (N_33677,N_26090,N_23480);
and U33678 (N_33678,N_20943,N_23841);
nor U33679 (N_33679,N_27468,N_25454);
xnor U33680 (N_33680,N_22103,N_22493);
xor U33681 (N_33681,N_26026,N_27161);
and U33682 (N_33682,N_27281,N_23533);
nand U33683 (N_33683,N_24398,N_24843);
and U33684 (N_33684,N_24388,N_26781);
nand U33685 (N_33685,N_26346,N_25940);
nand U33686 (N_33686,N_27996,N_24951);
nand U33687 (N_33687,N_22943,N_21979);
nor U33688 (N_33688,N_22853,N_27366);
xor U33689 (N_33689,N_23534,N_23167);
or U33690 (N_33690,N_29981,N_27185);
nor U33691 (N_33691,N_22086,N_29524);
or U33692 (N_33692,N_20351,N_22153);
nand U33693 (N_33693,N_27449,N_23319);
nor U33694 (N_33694,N_25873,N_20439);
and U33695 (N_33695,N_21115,N_20284);
nor U33696 (N_33696,N_28421,N_25274);
xnor U33697 (N_33697,N_22388,N_20044);
and U33698 (N_33698,N_24566,N_22561);
nor U33699 (N_33699,N_25087,N_21679);
or U33700 (N_33700,N_21992,N_21424);
and U33701 (N_33701,N_24957,N_22740);
and U33702 (N_33702,N_23069,N_20288);
xor U33703 (N_33703,N_26283,N_27507);
xor U33704 (N_33704,N_26747,N_25584);
nand U33705 (N_33705,N_20126,N_21822);
nand U33706 (N_33706,N_26604,N_22897);
or U33707 (N_33707,N_27406,N_24644);
or U33708 (N_33708,N_27465,N_23450);
and U33709 (N_33709,N_22836,N_25762);
nor U33710 (N_33710,N_24099,N_20639);
and U33711 (N_33711,N_28800,N_23285);
nand U33712 (N_33712,N_23897,N_24162);
or U33713 (N_33713,N_23558,N_28358);
nand U33714 (N_33714,N_26617,N_21641);
nand U33715 (N_33715,N_25064,N_21243);
xor U33716 (N_33716,N_24816,N_21328);
nor U33717 (N_33717,N_26918,N_24697);
nand U33718 (N_33718,N_24289,N_20187);
nand U33719 (N_33719,N_25670,N_21968);
and U33720 (N_33720,N_28245,N_28956);
or U33721 (N_33721,N_20821,N_29297);
xor U33722 (N_33722,N_23493,N_27213);
nor U33723 (N_33723,N_24841,N_24764);
nand U33724 (N_33724,N_22895,N_24075);
xor U33725 (N_33725,N_26722,N_22645);
nor U33726 (N_33726,N_22010,N_24177);
xnor U33727 (N_33727,N_20523,N_21457);
nor U33728 (N_33728,N_22208,N_22835);
and U33729 (N_33729,N_23993,N_26339);
or U33730 (N_33730,N_23857,N_24695);
nand U33731 (N_33731,N_29961,N_21492);
nand U33732 (N_33732,N_20107,N_20531);
xnor U33733 (N_33733,N_25982,N_25113);
nand U33734 (N_33734,N_29878,N_20225);
and U33735 (N_33735,N_28711,N_29975);
or U33736 (N_33736,N_23252,N_27380);
xor U33737 (N_33737,N_27699,N_25828);
nand U33738 (N_33738,N_20789,N_21098);
or U33739 (N_33739,N_29067,N_22714);
and U33740 (N_33740,N_25219,N_24768);
or U33741 (N_33741,N_27958,N_25605);
nor U33742 (N_33742,N_24688,N_28920);
nor U33743 (N_33743,N_26759,N_20509);
nand U33744 (N_33744,N_27032,N_24435);
nor U33745 (N_33745,N_21788,N_25589);
or U33746 (N_33746,N_20088,N_26557);
nand U33747 (N_33747,N_22597,N_25192);
or U33748 (N_33748,N_28333,N_26522);
nor U33749 (N_33749,N_20400,N_20220);
nor U33750 (N_33750,N_22810,N_23358);
nand U33751 (N_33751,N_27557,N_26585);
xnor U33752 (N_33752,N_25966,N_21591);
and U33753 (N_33753,N_20106,N_27546);
and U33754 (N_33754,N_29681,N_28590);
xor U33755 (N_33755,N_24774,N_24767);
or U33756 (N_33756,N_29809,N_29328);
or U33757 (N_33757,N_21629,N_29671);
nor U33758 (N_33758,N_27500,N_27498);
nor U33759 (N_33759,N_28145,N_26929);
or U33760 (N_33760,N_25874,N_24920);
xor U33761 (N_33761,N_26365,N_26316);
nor U33762 (N_33762,N_25426,N_23566);
and U33763 (N_33763,N_28991,N_25480);
and U33764 (N_33764,N_28981,N_28010);
nand U33765 (N_33765,N_22629,N_23448);
and U33766 (N_33766,N_26247,N_23767);
and U33767 (N_33767,N_21610,N_22761);
nand U33768 (N_33768,N_23040,N_25822);
nand U33769 (N_33769,N_21464,N_27322);
and U33770 (N_33770,N_27325,N_29202);
or U33771 (N_33771,N_21921,N_23296);
xor U33772 (N_33772,N_28324,N_23126);
nand U33773 (N_33773,N_20014,N_22221);
and U33774 (N_33774,N_23003,N_29151);
and U33775 (N_33775,N_25181,N_22243);
or U33776 (N_33776,N_27814,N_28944);
or U33777 (N_33777,N_27018,N_27283);
xnor U33778 (N_33778,N_25144,N_21005);
xnor U33779 (N_33779,N_25318,N_23953);
and U33780 (N_33780,N_20874,N_27299);
nor U33781 (N_33781,N_28950,N_22374);
nor U33782 (N_33782,N_22129,N_29180);
xor U33783 (N_33783,N_26583,N_23433);
or U33784 (N_33784,N_25010,N_21714);
nand U33785 (N_33785,N_24647,N_29539);
and U33786 (N_33786,N_27989,N_28268);
or U33787 (N_33787,N_20601,N_21430);
or U33788 (N_33788,N_24811,N_26498);
and U33789 (N_33789,N_20033,N_26755);
nand U33790 (N_33790,N_21677,N_20967);
or U33791 (N_33791,N_27200,N_29059);
xor U33792 (N_33792,N_28148,N_20487);
or U33793 (N_33793,N_27842,N_20174);
and U33794 (N_33794,N_28201,N_28192);
nand U33795 (N_33795,N_21774,N_25663);
or U33796 (N_33796,N_28524,N_23647);
xor U33797 (N_33797,N_20401,N_29891);
nor U33798 (N_33798,N_28969,N_21530);
nor U33799 (N_33799,N_27154,N_23982);
or U33800 (N_33800,N_28827,N_27973);
or U33801 (N_33801,N_23711,N_23721);
nor U33802 (N_33802,N_23090,N_23153);
nor U33803 (N_33803,N_21105,N_23633);
or U33804 (N_33804,N_21571,N_23742);
or U33805 (N_33805,N_22126,N_25641);
or U33806 (N_33806,N_24972,N_26019);
or U33807 (N_33807,N_25157,N_24654);
or U33808 (N_33808,N_27170,N_27646);
nor U33809 (N_33809,N_26693,N_22198);
xor U33810 (N_33810,N_27634,N_20738);
or U33811 (N_33811,N_21965,N_27354);
xor U33812 (N_33812,N_29630,N_24804);
or U33813 (N_33813,N_22967,N_22125);
or U33814 (N_33814,N_22511,N_20219);
nor U33815 (N_33815,N_25268,N_27160);
or U33816 (N_33816,N_25807,N_24327);
nand U33817 (N_33817,N_22982,N_25221);
nand U33818 (N_33818,N_21058,N_23652);
nor U33819 (N_33819,N_22143,N_21076);
or U33820 (N_33820,N_22343,N_21628);
nor U33821 (N_33821,N_29978,N_27078);
nor U33822 (N_33822,N_27091,N_25899);
nor U33823 (N_33823,N_24813,N_26145);
and U33824 (N_33824,N_25561,N_21955);
xnor U33825 (N_33825,N_22793,N_22007);
nand U33826 (N_33826,N_26548,N_23663);
nand U33827 (N_33827,N_26104,N_29492);
nor U33828 (N_33828,N_25247,N_23482);
xor U33829 (N_33829,N_20647,N_27988);
and U33830 (N_33830,N_29830,N_23191);
or U33831 (N_33831,N_20547,N_21994);
nor U33832 (N_33832,N_27992,N_22293);
and U33833 (N_33833,N_27816,N_21437);
nor U33834 (N_33834,N_29930,N_20695);
xnor U33835 (N_33835,N_20869,N_20621);
nand U33836 (N_33836,N_29079,N_29207);
nand U33837 (N_33837,N_21093,N_24694);
xor U33838 (N_33838,N_21319,N_20806);
xnor U33839 (N_33839,N_24898,N_27471);
xor U33840 (N_33840,N_29387,N_29920);
nand U33841 (N_33841,N_21296,N_27809);
xnor U33842 (N_33842,N_21521,N_26743);
nor U33843 (N_33843,N_29152,N_22172);
or U33844 (N_33844,N_20331,N_28644);
xnor U33845 (N_33845,N_21676,N_28587);
or U33846 (N_33846,N_29001,N_21186);
and U33847 (N_33847,N_20840,N_21803);
or U33848 (N_33848,N_26394,N_22147);
or U33849 (N_33849,N_28792,N_26621);
nor U33850 (N_33850,N_20562,N_28058);
xor U33851 (N_33851,N_26354,N_24809);
nand U33852 (N_33852,N_26688,N_27403);
or U33853 (N_33853,N_22959,N_25122);
or U33854 (N_33854,N_27135,N_24309);
xnor U33855 (N_33855,N_20103,N_26638);
and U33856 (N_33856,N_27738,N_29310);
nor U33857 (N_33857,N_25833,N_26966);
xnor U33858 (N_33858,N_23001,N_26528);
nand U33859 (N_33859,N_24232,N_28812);
nand U33860 (N_33860,N_26485,N_28744);
or U33861 (N_33861,N_23019,N_23740);
and U33862 (N_33862,N_21584,N_21588);
or U33863 (N_33863,N_21484,N_26991);
nand U33864 (N_33864,N_23389,N_27540);
xor U33865 (N_33865,N_26447,N_27539);
nand U33866 (N_33866,N_22203,N_20544);
nand U33867 (N_33867,N_24328,N_23353);
or U33868 (N_33868,N_29927,N_28492);
nor U33869 (N_33869,N_20049,N_29580);
xnor U33870 (N_33870,N_23349,N_23949);
xor U33871 (N_33871,N_23346,N_24888);
or U33872 (N_33872,N_27800,N_20038);
xor U33873 (N_33873,N_22139,N_20353);
xnor U33874 (N_33874,N_23608,N_20457);
and U33875 (N_33875,N_25312,N_29771);
and U33876 (N_33876,N_21695,N_26377);
xnor U33877 (N_33877,N_21800,N_20443);
nand U33878 (N_33878,N_25826,N_29183);
nor U33879 (N_33879,N_27774,N_20832);
nor U33880 (N_33880,N_29501,N_28560);
nand U33881 (N_33881,N_26265,N_21447);
and U33882 (N_33882,N_20034,N_20889);
or U33883 (N_33883,N_23195,N_27359);
nand U33884 (N_33884,N_28629,N_21589);
or U33885 (N_33885,N_22092,N_23047);
nand U33886 (N_33886,N_25524,N_21312);
or U33887 (N_33887,N_26033,N_21318);
or U33888 (N_33888,N_26239,N_25277);
or U33889 (N_33889,N_28672,N_20743);
and U33890 (N_33890,N_23397,N_27951);
and U33891 (N_33891,N_24342,N_24223);
nor U33892 (N_33892,N_28334,N_24907);
nand U33893 (N_33893,N_21547,N_25666);
and U33894 (N_33894,N_28772,N_26569);
xnor U33895 (N_33895,N_25547,N_21874);
xnor U33896 (N_33896,N_20643,N_24137);
and U33897 (N_33897,N_26841,N_20163);
xor U33898 (N_33898,N_27006,N_23067);
xnor U33899 (N_33899,N_29634,N_26166);
xnor U33900 (N_33900,N_20899,N_27706);
nand U33901 (N_33901,N_29521,N_28372);
and U33902 (N_33902,N_24728,N_25972);
xor U33903 (N_33903,N_20518,N_23156);
and U33904 (N_33904,N_20164,N_26587);
nand U33905 (N_33905,N_23954,N_28822);
and U33906 (N_33906,N_20978,N_20672);
xnor U33907 (N_33907,N_26471,N_21066);
xnor U33908 (N_33908,N_20224,N_20488);
xnor U33909 (N_33909,N_28598,N_22186);
nor U33910 (N_33910,N_27064,N_27301);
and U33911 (N_33911,N_29789,N_26594);
nor U33912 (N_33912,N_20706,N_21858);
and U33913 (N_33913,N_22609,N_25261);
and U33914 (N_33914,N_29841,N_24158);
or U33915 (N_33915,N_23492,N_23345);
and U33916 (N_33916,N_22171,N_21007);
and U33917 (N_33917,N_28002,N_26242);
nor U33918 (N_33918,N_21556,N_28676);
and U33919 (N_33919,N_20354,N_29121);
nor U33920 (N_33920,N_22688,N_28828);
nand U33921 (N_33921,N_27511,N_26507);
nor U33922 (N_33922,N_28120,N_21429);
nor U33923 (N_33923,N_20173,N_27780);
or U33924 (N_33924,N_21488,N_25478);
and U33925 (N_33925,N_24189,N_22100);
and U33926 (N_33926,N_24152,N_26518);
or U33927 (N_33927,N_28247,N_21536);
nand U33928 (N_33928,N_28882,N_22839);
nand U33929 (N_33929,N_23382,N_26768);
nor U33930 (N_33930,N_29884,N_25551);
and U33931 (N_33931,N_28698,N_24100);
and U33932 (N_33932,N_27008,N_26307);
nor U33933 (N_33933,N_20422,N_26837);
or U33934 (N_33934,N_27012,N_25035);
nand U33935 (N_33935,N_26619,N_27819);
xnor U33936 (N_33936,N_29727,N_26209);
and U33937 (N_33937,N_21114,N_29284);
xnor U33938 (N_33938,N_29576,N_27475);
and U33939 (N_33939,N_25654,N_20545);
or U33940 (N_33940,N_21228,N_28990);
nor U33941 (N_33941,N_27320,N_26971);
nor U33942 (N_33942,N_27536,N_27695);
nand U33943 (N_33943,N_21266,N_26713);
or U33944 (N_33944,N_26057,N_26416);
nand U33945 (N_33945,N_24504,N_26405);
xor U33946 (N_33946,N_20272,N_22291);
and U33947 (N_33947,N_25384,N_22630);
nand U33948 (N_33948,N_22341,N_24446);
or U33949 (N_33949,N_26241,N_25588);
nand U33950 (N_33950,N_20530,N_25346);
nor U33951 (N_33951,N_22588,N_25676);
and U33952 (N_33952,N_24547,N_27316);
and U33953 (N_33953,N_25393,N_21685);
xor U33954 (N_33954,N_21261,N_23305);
nor U33955 (N_33955,N_29585,N_27149);
or U33956 (N_33956,N_29375,N_27983);
xnor U33957 (N_33957,N_22883,N_23230);
nor U33958 (N_33958,N_21880,N_21929);
xor U33959 (N_33959,N_22602,N_26831);
and U33960 (N_33960,N_20787,N_23138);
nor U33961 (N_33961,N_24925,N_28258);
or U33962 (N_33962,N_25656,N_25224);
or U33963 (N_33963,N_26682,N_23836);
xor U33964 (N_33964,N_27614,N_27416);
nand U33965 (N_33965,N_21702,N_21404);
nand U33966 (N_33966,N_25159,N_25804);
nand U33967 (N_33967,N_23495,N_24200);
xor U33968 (N_33968,N_26220,N_26850);
nand U33969 (N_33969,N_20876,N_22260);
or U33970 (N_33970,N_21932,N_20771);
or U33971 (N_33971,N_24853,N_24385);
and U33972 (N_33972,N_23958,N_26926);
xor U33973 (N_33973,N_28693,N_21411);
nor U33974 (N_33974,N_24933,N_29072);
nor U33975 (N_33975,N_28167,N_24520);
xnor U33976 (N_33976,N_29165,N_21455);
and U33977 (N_33977,N_28872,N_22256);
xnor U33978 (N_33978,N_24675,N_29592);
and U33979 (N_33979,N_28376,N_20611);
nor U33980 (N_33980,N_24873,N_21733);
or U33981 (N_33981,N_26686,N_20998);
nor U33982 (N_33982,N_25253,N_23278);
nand U33983 (N_33983,N_29145,N_22382);
xnor U33984 (N_33984,N_28488,N_28612);
or U33985 (N_33985,N_20810,N_23043);
or U33986 (N_33986,N_29794,N_21662);
or U33987 (N_33987,N_25796,N_22470);
or U33988 (N_33988,N_26727,N_21271);
nand U33989 (N_33989,N_23277,N_24720);
nor U33990 (N_33990,N_27944,N_21077);
nor U33991 (N_33991,N_25609,N_29915);
nand U33992 (N_33992,N_21468,N_22405);
nor U33993 (N_33993,N_22879,N_29713);
or U33994 (N_33994,N_25942,N_27336);
and U33995 (N_33995,N_24228,N_22544);
and U33996 (N_33996,N_21543,N_20992);
and U33997 (N_33997,N_24021,N_26993);
or U33998 (N_33998,N_24183,N_29264);
nand U33999 (N_33999,N_20229,N_26560);
and U34000 (N_34000,N_24895,N_23719);
and U34001 (N_34001,N_21585,N_29532);
xor U34002 (N_34002,N_29578,N_22240);
or U34003 (N_34003,N_21358,N_23797);
or U34004 (N_34004,N_20137,N_25328);
and U34005 (N_34005,N_20768,N_21638);
nand U34006 (N_34006,N_24238,N_26778);
nand U34007 (N_34007,N_23224,N_27183);
and U34008 (N_34008,N_24407,N_28107);
nor U34009 (N_34009,N_25103,N_20159);
xor U34010 (N_34010,N_20432,N_24064);
and U34011 (N_34011,N_20068,N_25430);
and U34012 (N_34012,N_24055,N_28845);
nor U34013 (N_34013,N_28346,N_21184);
and U34014 (N_34014,N_25193,N_21287);
and U34015 (N_34015,N_26412,N_29144);
xor U34016 (N_34016,N_26452,N_24565);
nor U34017 (N_34017,N_20969,N_22725);
and U34018 (N_34018,N_25623,N_20303);
nand U34019 (N_34019,N_21388,N_29211);
nand U34020 (N_34020,N_22384,N_26714);
and U34021 (N_34021,N_27384,N_25255);
nor U34022 (N_34022,N_28190,N_26974);
and U34023 (N_34023,N_29787,N_29399);
nand U34024 (N_34024,N_26082,N_28922);
nand U34025 (N_34025,N_28272,N_28898);
xnor U34026 (N_34026,N_26193,N_23701);
nor U34027 (N_34027,N_20214,N_20955);
or U34028 (N_34028,N_20433,N_24926);
nor U34029 (N_34029,N_29007,N_27044);
xor U34030 (N_34030,N_22141,N_26532);
nor U34031 (N_34031,N_20380,N_22176);
and U34032 (N_34032,N_27112,N_26216);
or U34033 (N_34033,N_23573,N_24824);
or U34034 (N_34034,N_23858,N_23434);
nor U34035 (N_34035,N_29571,N_26853);
xor U34036 (N_34036,N_22837,N_26102);
nor U34037 (N_34037,N_28442,N_20759);
nor U34038 (N_34038,N_27279,N_23106);
xor U34039 (N_34039,N_21281,N_28895);
nor U34040 (N_34040,N_23424,N_29461);
or U34041 (N_34041,N_25984,N_27822);
xor U34042 (N_34042,N_24611,N_24478);
nand U34043 (N_34043,N_23895,N_22623);
xnor U34044 (N_34044,N_27410,N_20389);
or U34045 (N_34045,N_22605,N_29845);
and U34046 (N_34046,N_28736,N_20983);
or U34047 (N_34047,N_25314,N_26647);
nor U34048 (N_34048,N_28866,N_21687);
nor U34049 (N_34049,N_25946,N_25481);
and U34050 (N_34050,N_29983,N_24414);
xnor U34051 (N_34051,N_26564,N_24970);
nand U34052 (N_34052,N_22414,N_29693);
nand U34053 (N_34053,N_28311,N_29065);
and U34054 (N_34054,N_24522,N_26077);
or U34055 (N_34055,N_29922,N_22336);
nand U34056 (N_34056,N_22801,N_25817);
and U34057 (N_34057,N_28233,N_26489);
nor U34058 (N_34058,N_20662,N_28686);
or U34059 (N_34059,N_25151,N_29799);
nand U34060 (N_34060,N_23576,N_20119);
and U34061 (N_34061,N_25083,N_23455);
xor U34062 (N_34062,N_28343,N_24103);
nor U34063 (N_34063,N_23753,N_26053);
nand U34064 (N_34064,N_21366,N_25816);
and U34065 (N_34065,N_20881,N_27094);
nand U34066 (N_34066,N_26816,N_29684);
xor U34067 (N_34067,N_24147,N_21522);
or U34068 (N_34068,N_24488,N_21107);
nand U34069 (N_34069,N_28588,N_23735);
and U34070 (N_34070,N_22902,N_27651);
and U34071 (N_34071,N_29257,N_24017);
xor U34072 (N_34072,N_27121,N_25747);
xor U34073 (N_34073,N_22923,N_21223);
xnor U34074 (N_34074,N_20650,N_20337);
xor U34075 (N_34075,N_26614,N_28240);
nand U34076 (N_34076,N_20348,N_21039);
nor U34077 (N_34077,N_25693,N_26975);
nor U34078 (N_34078,N_25256,N_20313);
and U34079 (N_34079,N_26656,N_22432);
and U34080 (N_34080,N_21177,N_21079);
xnor U34081 (N_34081,N_23914,N_27178);
nand U34082 (N_34082,N_23303,N_29535);
nor U34083 (N_34083,N_22996,N_21854);
nand U34084 (N_34084,N_25377,N_21083);
xor U34085 (N_34085,N_26343,N_24854);
nand U34086 (N_34086,N_22912,N_23056);
xor U34087 (N_34087,N_22473,N_20258);
nand U34088 (N_34088,N_29206,N_22825);
and U34089 (N_34089,N_27708,N_28366);
nand U34090 (N_34090,N_27672,N_26396);
xnor U34091 (N_34091,N_28825,N_24580);
or U34092 (N_34092,N_21490,N_29392);
nor U34093 (N_34093,N_25728,N_21728);
nor U34094 (N_34094,N_24552,N_20855);
xnor U34095 (N_34095,N_27532,N_22188);
or U34096 (N_34096,N_24292,N_21555);
nor U34097 (N_34097,N_28278,N_24072);
xnor U34098 (N_34098,N_24657,N_20104);
xor U34099 (N_34099,N_24393,N_25069);
xor U34100 (N_34100,N_28948,N_21034);
or U34101 (N_34101,N_21067,N_23328);
or U34102 (N_34102,N_29649,N_26854);
nand U34103 (N_34103,N_22254,N_26513);
nand U34104 (N_34104,N_27987,N_28784);
or U34105 (N_34105,N_24494,N_23720);
xor U34106 (N_34106,N_23635,N_27575);
or U34107 (N_34107,N_21240,N_21796);
nand U34108 (N_34108,N_20388,N_27880);
xnor U34109 (N_34109,N_25632,N_23411);
and U34110 (N_34110,N_21936,N_29194);
xor U34111 (N_34111,N_24087,N_26309);
nand U34112 (N_34112,N_21330,N_25085);
and U34113 (N_34113,N_25327,N_26192);
nor U34114 (N_34114,N_22642,N_21636);
nor U34115 (N_34115,N_24896,N_27622);
and U34116 (N_34116,N_20802,N_28371);
xor U34117 (N_34117,N_26717,N_28180);
or U34118 (N_34118,N_23377,N_27476);
xnor U34119 (N_34119,N_22338,N_25048);
and U34120 (N_34120,N_26636,N_25400);
xnor U34121 (N_34121,N_27982,N_20059);
and U34122 (N_34122,N_27534,N_25917);
or U34123 (N_34123,N_21935,N_20042);
or U34124 (N_34124,N_26701,N_26995);
and U34125 (N_34125,N_27256,N_23782);
nor U34126 (N_34126,N_28831,N_26473);
xnor U34127 (N_34127,N_23002,N_29661);
xnor U34128 (N_34128,N_20497,N_28690);
nor U34129 (N_34129,N_21916,N_23091);
and U34130 (N_34130,N_22459,N_28733);
nor U34131 (N_34131,N_26506,N_26580);
and U34132 (N_34132,N_27057,N_28817);
nand U34133 (N_34133,N_23456,N_23013);
nor U34134 (N_34134,N_29715,N_20609);
or U34135 (N_34135,N_22342,N_21908);
and U34136 (N_34136,N_22271,N_23732);
nand U34137 (N_34137,N_27123,N_24942);
nand U34138 (N_34138,N_26990,N_27803);
xnor U34139 (N_34139,N_20736,N_28039);
and U34140 (N_34140,N_26479,N_27525);
or U34141 (N_34141,N_21948,N_20664);
xnor U34142 (N_34142,N_20702,N_21127);
xnor U34143 (N_34143,N_28322,N_28797);
xor U34144 (N_34144,N_25070,N_24444);
nor U34145 (N_34145,N_20211,N_27554);
and U34146 (N_34146,N_24483,N_21780);
nand U34147 (N_34147,N_27902,N_25671);
xor U34148 (N_34148,N_25139,N_29019);
nand U34149 (N_34149,N_27232,N_25022);
and U34150 (N_34150,N_29174,N_23238);
xor U34151 (N_34151,N_22878,N_29096);
and U34152 (N_34152,N_20511,N_25686);
xnor U34153 (N_34153,N_27503,N_27589);
xor U34154 (N_34154,N_27001,N_27950);
and U34155 (N_34155,N_20418,N_29733);
and U34156 (N_34156,N_26353,N_29125);
nor U34157 (N_34157,N_26075,N_20036);
and U34158 (N_34158,N_22332,N_23812);
xor U34159 (N_34159,N_25464,N_24751);
nand U34160 (N_34160,N_23065,N_25120);
nor U34161 (N_34161,N_26155,N_28513);
and U34162 (N_34162,N_27565,N_22428);
nor U34163 (N_34163,N_21494,N_29520);
nand U34164 (N_34164,N_28750,N_25061);
or U34165 (N_34165,N_22500,N_26920);
nand U34166 (N_34166,N_23823,N_28633);
and U34167 (N_34167,N_24827,N_20281);
or U34168 (N_34168,N_21449,N_28011);
nand U34169 (N_34169,N_29305,N_25133);
and U34170 (N_34170,N_23414,N_28222);
nor U34171 (N_34171,N_28730,N_27596);
and U34172 (N_34172,N_25353,N_25530);
nor U34173 (N_34173,N_25082,N_29076);
or U34174 (N_34174,N_29142,N_27352);
or U34175 (N_34175,N_23775,N_25698);
nor U34176 (N_34176,N_21031,N_23656);
nor U34177 (N_34177,N_22109,N_28000);
xor U34178 (N_34178,N_23459,N_22509);
xnor U34179 (N_34179,N_20891,N_28297);
and U34180 (N_34180,N_28871,N_28070);
nor U34181 (N_34181,N_20006,N_23778);
xor U34182 (N_34182,N_29371,N_26468);
xor U34183 (N_34183,N_28986,N_22224);
or U34184 (N_34184,N_21474,N_21834);
xor U34185 (N_34185,N_20387,N_21557);
nand U34186 (N_34186,N_23690,N_27653);
nor U34187 (N_34187,N_25313,N_22744);
nor U34188 (N_34188,N_26202,N_21927);
and U34189 (N_34189,N_22295,N_25356);
and U34190 (N_34190,N_29338,N_21061);
xnor U34191 (N_34191,N_29870,N_28694);
xor U34192 (N_34192,N_20011,N_21595);
and U34193 (N_34193,N_29500,N_25691);
or U34194 (N_34194,N_28999,N_23976);
or U34195 (N_34195,N_26248,N_23575);
and U34196 (N_34196,N_29318,N_25744);
and U34197 (N_34197,N_26667,N_25127);
xnor U34198 (N_34198,N_24264,N_28597);
nand U34199 (N_34199,N_23234,N_26221);
xnor U34200 (N_34200,N_26932,N_21732);
nor U34201 (N_34201,N_23784,N_26649);
nor U34202 (N_34202,N_20319,N_21957);
and U34203 (N_34203,N_29730,N_26261);
xnor U34204 (N_34204,N_21451,N_22920);
nor U34205 (N_34205,N_25583,N_22892);
and U34206 (N_34206,N_28246,N_28835);
nand U34207 (N_34207,N_20627,N_27754);
nor U34208 (N_34208,N_23166,N_21395);
xnor U34209 (N_34209,N_22297,N_22872);
nor U34210 (N_34210,N_22015,N_24324);
nor U34211 (N_34211,N_29606,N_28109);
xor U34212 (N_34212,N_25504,N_21322);
or U34213 (N_34213,N_29303,N_22390);
and U34214 (N_34214,N_25052,N_20640);
nand U34215 (N_34215,N_29518,N_26039);
xor U34216 (N_34216,N_26697,N_22436);
or U34217 (N_34217,N_29911,N_23481);
nand U34218 (N_34218,N_24150,N_22223);
nand U34219 (N_34219,N_28580,N_29316);
nor U34220 (N_34220,N_23231,N_20052);
and U34221 (N_34221,N_27116,N_22231);
or U34222 (N_34222,N_23321,N_25452);
xnor U34223 (N_34223,N_24145,N_29752);
nand U34224 (N_34224,N_25299,N_27456);
and U34225 (N_34225,N_29110,N_26356);
and U34226 (N_34226,N_27081,N_24601);
and U34227 (N_34227,N_26884,N_25062);
nand U34228 (N_34228,N_29409,N_27870);
xnor U34229 (N_34229,N_23779,N_26609);
nor U34230 (N_34230,N_23736,N_21742);
or U34231 (N_34231,N_27047,N_25417);
nand U34232 (N_34232,N_22347,N_25287);
or U34233 (N_34233,N_27863,N_22396);
nand U34234 (N_34234,N_26421,N_22627);
or U34235 (N_34235,N_20499,N_28875);
and U34236 (N_34236,N_24948,N_27681);
nor U34237 (N_34237,N_24377,N_27487);
and U34238 (N_34238,N_20808,N_20566);
nor U34239 (N_34239,N_23600,N_29004);
nand U34240 (N_34240,N_28142,N_27917);
and U34241 (N_34241,N_21527,N_21428);
nand U34242 (N_34242,N_23031,N_24932);
nand U34243 (N_34243,N_20255,N_26379);
nor U34244 (N_34244,N_28172,N_24296);
xor U34245 (N_34245,N_22101,N_25770);
and U34246 (N_34246,N_25294,N_26798);
nor U34247 (N_34247,N_21335,N_29444);
and U34248 (N_34248,N_25739,N_27439);
and U34249 (N_34249,N_23508,N_20774);
nor U34250 (N_34250,N_26378,N_21514);
and U34251 (N_34251,N_20922,N_24051);
nand U34252 (N_34252,N_26822,N_26525);
nor U34253 (N_34253,N_28511,N_28139);
nand U34254 (N_34254,N_20635,N_29166);
nor U34255 (N_34255,N_26586,N_27841);
nor U34256 (N_34256,N_23269,N_24170);
nand U34257 (N_34257,N_26704,N_22829);
and U34258 (N_34258,N_23246,N_26808);
or U34259 (N_34259,N_22787,N_25936);
xor U34260 (N_34260,N_24979,N_22149);
or U34261 (N_34261,N_28771,N_20856);
xor U34262 (N_34262,N_20883,N_25746);
or U34263 (N_34263,N_20866,N_20349);
and U34264 (N_34264,N_25160,N_29091);
xor U34265 (N_34265,N_24219,N_27971);
xor U34266 (N_34266,N_23774,N_27448);
and U34267 (N_34267,N_22275,N_25977);
xnor U34268 (N_34268,N_20907,N_24486);
or U34269 (N_34269,N_29699,N_28685);
nand U34270 (N_34270,N_26590,N_29657);
nand U34271 (N_34271,N_25700,N_27953);
nand U34272 (N_34272,N_27597,N_23856);
and U34273 (N_34273,N_28018,N_24513);
xor U34274 (N_34274,N_24040,N_26572);
xor U34275 (N_34275,N_29311,N_21094);
and U34276 (N_34276,N_29285,N_26791);
nand U34277 (N_34277,N_24913,N_29938);
and U34278 (N_34278,N_24195,N_28989);
or U34279 (N_34279,N_25573,N_27828);
or U34280 (N_34280,N_23902,N_27223);
or U34281 (N_34281,N_21651,N_24723);
xor U34282 (N_34282,N_21220,N_21043);
or U34283 (N_34283,N_23470,N_29889);
xor U34284 (N_34284,N_25538,N_20102);
and U34285 (N_34285,N_26268,N_29545);
xnor U34286 (N_34286,N_27758,N_27564);
xor U34287 (N_34287,N_26438,N_29104);
xnor U34288 (N_34288,N_22017,N_23400);
and U34289 (N_34289,N_24807,N_20458);
or U34290 (N_34290,N_25101,N_22939);
and U34291 (N_34291,N_22873,N_26826);
nor U34292 (N_34292,N_20522,N_23352);
and U34293 (N_34293,N_29726,N_29414);
or U34294 (N_34294,N_29641,N_25386);
and U34295 (N_34295,N_24346,N_28819);
xnor U34296 (N_34296,N_27671,N_28302);
xor U34297 (N_34297,N_23119,N_25916);
xor U34298 (N_34298,N_21608,N_21905);
nor U34299 (N_34299,N_26285,N_29820);
nand U34300 (N_34300,N_24784,N_26281);
nand U34301 (N_34301,N_28725,N_26856);
and U34302 (N_34302,N_27092,N_25403);
xnor U34303 (N_34303,N_24863,N_28732);
nand U34304 (N_34304,N_29623,N_26453);
and U34305 (N_34305,N_27429,N_20230);
and U34306 (N_34306,N_20707,N_29700);
xnor U34307 (N_34307,N_26397,N_24560);
nor U34308 (N_34308,N_21018,N_23660);
nand U34309 (N_34309,N_22587,N_25979);
nand U34310 (N_34310,N_25307,N_29063);
or U34311 (N_34311,N_26664,N_23178);
and U34312 (N_34312,N_20217,N_28153);
xor U34313 (N_34313,N_21454,N_28393);
nor U34314 (N_34314,N_22659,N_22510);
and U34315 (N_34315,N_29945,N_28473);
nor U34316 (N_34316,N_24527,N_29204);
nor U34317 (N_34317,N_27641,N_22674);
or U34318 (N_34318,N_23838,N_26799);
and U34319 (N_34319,N_25385,N_21056);
and U34320 (N_34320,N_29088,N_25278);
and U34321 (N_34321,N_24993,N_26003);
nor U34322 (N_34322,N_28830,N_28663);
and U34323 (N_34323,N_23479,N_25962);
and U34324 (N_34324,N_24936,N_24403);
xor U34325 (N_34325,N_23828,N_28118);
or U34326 (N_34326,N_26020,N_23694);
xnor U34327 (N_34327,N_29778,N_23743);
nand U34328 (N_34328,N_28206,N_27293);
and U34329 (N_34329,N_25699,N_24320);
xnor U34330 (N_34330,N_29647,N_23223);
and U34331 (N_34331,N_24452,N_29393);
or U34332 (N_34332,N_20060,N_29139);
xnor U34333 (N_34333,N_29209,N_27723);
nor U34334 (N_34334,N_28569,N_26669);
nand U34335 (N_34335,N_28399,N_20915);
nand U34336 (N_34336,N_29434,N_22604);
xnor U34337 (N_34337,N_26868,N_24897);
or U34338 (N_34338,N_28606,N_24766);
and U34339 (N_34339,N_21063,N_26385);
nor U34340 (N_34340,N_24144,N_27625);
and U34341 (N_34341,N_26640,N_24303);
or U34342 (N_34342,N_22407,N_21181);
and U34343 (N_34343,N_24885,N_27068);
nand U34344 (N_34344,N_24859,N_27911);
nor U34345 (N_34345,N_28225,N_21887);
nor U34346 (N_34346,N_29819,N_23041);
and U34347 (N_34347,N_21122,N_21160);
nand U34348 (N_34348,N_28878,N_27688);
and U34349 (N_34349,N_25657,N_27661);
nand U34350 (N_34350,N_27168,N_25018);
nand U34351 (N_34351,N_22392,N_24124);
or U34352 (N_34352,N_29216,N_20685);
nor U34353 (N_34353,N_28390,N_21325);
xnor U34354 (N_34354,N_24716,N_28484);
or U34355 (N_34355,N_27871,N_23405);
nand U34356 (N_34356,N_20382,N_20593);
nor U34357 (N_34357,N_27025,N_28191);
xnor U34358 (N_34358,N_22189,N_27310);
nand U34359 (N_34359,N_25932,N_27426);
nand U34360 (N_34360,N_22929,N_22848);
nand U34361 (N_34361,N_23579,N_21409);
nand U34362 (N_34362,N_25918,N_24265);
nand U34363 (N_34363,N_20274,N_20333);
and U34364 (N_34364,N_29382,N_23752);
nor U34365 (N_34365,N_20595,N_22781);
and U34366 (N_34366,N_25968,N_26736);
nor U34367 (N_34367,N_21895,N_21971);
xnor U34368 (N_34368,N_29340,N_29443);
or U34369 (N_34369,N_28228,N_24415);
nand U34370 (N_34370,N_28436,N_21952);
and U34371 (N_34371,N_26190,N_24660);
or U34372 (N_34372,N_24139,N_22871);
and U34373 (N_34373,N_29214,N_24528);
or U34374 (N_34374,N_28057,N_24600);
xor U34375 (N_34375,N_23730,N_22773);
nor U34376 (N_34376,N_24375,N_28092);
xor U34377 (N_34377,N_22607,N_22521);
nor U34378 (N_34378,N_27046,N_24463);
or U34379 (N_34379,N_22073,N_20542);
nand U34380 (N_34380,N_24880,N_25146);
xor U34381 (N_34381,N_23786,N_24322);
nor U34382 (N_34382,N_21111,N_20885);
or U34383 (N_34383,N_22247,N_24215);
or U34384 (N_34384,N_22543,N_23672);
nor U34385 (N_34385,N_21746,N_27943);
nand U34386 (N_34386,N_29452,N_27853);
xor U34387 (N_34387,N_23416,N_29420);
xor U34388 (N_34388,N_28870,N_24775);
and U34389 (N_34389,N_20300,N_23163);
xor U34390 (N_34390,N_21875,N_25483);
and U34391 (N_34391,N_23748,N_24468);
and U34392 (N_34392,N_21583,N_26180);
nand U34393 (N_34393,N_26908,N_25161);
nor U34394 (N_34394,N_28427,N_21421);
xor U34395 (N_34395,N_22949,N_21044);
or U34396 (N_34396,N_20041,N_26865);
and U34397 (N_34397,N_27897,N_24982);
nand U34398 (N_34398,N_27261,N_24449);
or U34399 (N_34399,N_23164,N_24578);
or U34400 (N_34400,N_26810,N_27378);
or U34401 (N_34401,N_20747,N_25711);
xor U34402 (N_34402,N_20501,N_27743);
nand U34403 (N_34403,N_29376,N_23308);
xor U34404 (N_34404,N_28671,N_25466);
nand U34405 (N_34405,N_27248,N_27204);
nand U34406 (N_34406,N_22391,N_29397);
nand U34407 (N_34407,N_26076,N_20055);
or U34408 (N_34408,N_21533,N_23950);
nand U34409 (N_34409,N_21752,N_21945);
and U34410 (N_34410,N_29839,N_21507);
nor U34411 (N_34411,N_22353,N_21480);
xnor U34412 (N_34412,N_23726,N_24616);
nor U34413 (N_34413,N_22765,N_20304);
or U34414 (N_34414,N_27807,N_29772);
and U34415 (N_34415,N_28483,N_26048);
or U34416 (N_34416,N_25880,N_25915);
nor U34417 (N_34417,N_21761,N_24288);
nor U34418 (N_34418,N_26942,N_21582);
nand U34419 (N_34419,N_28479,N_21463);
nand U34420 (N_34420,N_22524,N_29230);
and U34421 (N_34421,N_28658,N_28697);
nand U34422 (N_34422,N_27379,N_25811);
and U34423 (N_34423,N_23380,N_20786);
nor U34424 (N_34424,N_22036,N_24994);
nand U34425 (N_34425,N_21997,N_27523);
nor U34426 (N_34426,N_21134,N_22051);
and U34427 (N_34427,N_25228,N_29141);
or U34428 (N_34428,N_22704,N_23248);
nor U34429 (N_34429,N_25964,N_26252);
xor U34430 (N_34430,N_20155,N_25109);
and U34431 (N_34431,N_20884,N_27859);
nand U34432 (N_34432,N_26957,N_26127);
xnor U34433 (N_34433,N_29538,N_27239);
and U34434 (N_34434,N_27872,N_25629);
xor U34435 (N_34435,N_28760,N_25484);
xor U34436 (N_34436,N_29951,N_25669);
or U34437 (N_34437,N_29107,N_27211);
xor U34438 (N_34438,N_23304,N_27203);
or U34439 (N_34439,N_25825,N_29857);
xnor U34440 (N_34440,N_22104,N_23654);
nor U34441 (N_34441,N_21118,N_25021);
or U34442 (N_34442,N_21010,N_21028);
nor U34443 (N_34443,N_28911,N_26310);
or U34444 (N_34444,N_26406,N_25644);
nand U34445 (N_34445,N_28398,N_26809);
xnor U34446 (N_34446,N_28709,N_21068);
or U34447 (N_34447,N_27331,N_25025);
nand U34448 (N_34448,N_26740,N_20826);
nor U34449 (N_34449,N_28807,N_26944);
and U34450 (N_34450,N_25591,N_29343);
nand U34451 (N_34451,N_29742,N_22962);
or U34452 (N_34452,N_25397,N_27164);
and U34453 (N_34453,N_22735,N_24490);
and U34454 (N_34454,N_29286,N_25784);
nand U34455 (N_34455,N_28551,N_21124);
xor U34456 (N_34456,N_20984,N_27212);
nor U34457 (N_34457,N_25920,N_24747);
or U34458 (N_34458,N_21906,N_20087);
or U34459 (N_34459,N_22696,N_20101);
and U34460 (N_34460,N_21195,N_27144);
nand U34461 (N_34461,N_28526,N_22745);
and U34462 (N_34462,N_25401,N_25585);
and U34463 (N_34463,N_22655,N_21937);
and U34464 (N_34464,N_25712,N_23995);
or U34465 (N_34465,N_26763,N_24586);
or U34466 (N_34466,N_26644,N_24234);
xnor U34467 (N_34467,N_26470,N_26046);
and U34468 (N_34468,N_23454,N_20604);
nor U34469 (N_34469,N_27404,N_25198);
nand U34470 (N_34470,N_24092,N_28189);
and U34471 (N_34471,N_25092,N_25076);
xor U34472 (N_34472,N_20453,N_26696);
and U34473 (N_34473,N_28349,N_29293);
xor U34474 (N_34474,N_21942,N_22508);
xnor U34475 (N_34475,N_25674,N_22463);
and U34476 (N_34476,N_23849,N_27307);
and U34477 (N_34477,N_21607,N_25766);
and U34478 (N_34478,N_25864,N_29786);
nand U34479 (N_34479,N_23847,N_20875);
and U34480 (N_34480,N_27618,N_20167);
nor U34481 (N_34481,N_24662,N_20147);
nand U34482 (N_34482,N_22031,N_20944);
and U34483 (N_34483,N_23076,N_28890);
or U34484 (N_34484,N_20357,N_21574);
nor U34485 (N_34485,N_21865,N_28832);
and U34486 (N_34486,N_27502,N_26773);
nor U34487 (N_34487,N_24931,N_21632);
xnor U34488 (N_34488,N_22960,N_22809);
nor U34489 (N_34489,N_28836,N_26458);
or U34490 (N_34490,N_20063,N_26870);
nand U34491 (N_34491,N_28869,N_23161);
nor U34492 (N_34492,N_22439,N_21149);
or U34493 (N_34493,N_22479,N_23483);
and U34494 (N_34494,N_28972,N_21141);
and U34495 (N_34495,N_24032,N_28614);
or U34496 (N_34496,N_20470,N_21599);
xor U34497 (N_34497,N_21493,N_24621);
or U34498 (N_34498,N_27108,N_21644);
nand U34499 (N_34499,N_21153,N_20942);
or U34500 (N_34500,N_26753,N_28004);
nor U34501 (N_34501,N_24634,N_20399);
and U34502 (N_34502,N_23831,N_26684);
xnor U34503 (N_34503,N_25248,N_29810);
nor U34504 (N_34504,N_20945,N_23634);
or U34505 (N_34505,N_27011,N_27305);
and U34506 (N_34506,N_21425,N_24910);
and U34507 (N_34507,N_26021,N_23485);
xor U34508 (N_34508,N_29788,N_28751);
or U34509 (N_34509,N_27024,N_28262);
and U34510 (N_34510,N_27428,N_27356);
nor U34511 (N_34511,N_24319,N_28023);
nand U34512 (N_34512,N_25876,N_25616);
xor U34513 (N_34513,N_24887,N_27722);
and U34514 (N_34514,N_28954,N_27721);
or U34515 (N_34515,N_22181,N_25925);
nor U34516 (N_34516,N_20772,N_20668);
or U34517 (N_34517,N_23606,N_21691);
xnor U34518 (N_34518,N_27692,N_28069);
nand U34519 (N_34519,N_21448,N_27517);
and U34520 (N_34520,N_24039,N_23228);
and U34521 (N_34521,N_28782,N_28494);
nand U34522 (N_34522,N_27886,N_28904);
xnor U34523 (N_34523,N_21845,N_20156);
and U34524 (N_34524,N_29365,N_28043);
nor U34525 (N_34525,N_23162,N_29235);
nand U34526 (N_34526,N_28821,N_25510);
xor U34527 (N_34527,N_29972,N_28674);
or U34528 (N_34528,N_24220,N_23412);
nand U34529 (N_34529,N_27640,N_25326);
nor U34530 (N_34530,N_23968,N_20352);
and U34531 (N_34531,N_25148,N_24568);
or U34532 (N_34532,N_25422,N_28250);
nand U34533 (N_34533,N_23286,N_27684);
or U34534 (N_34534,N_28995,N_22956);
xor U34535 (N_34535,N_29937,N_27690);
nand U34536 (N_34536,N_25410,N_22563);
nor U34537 (N_34537,N_28213,N_25172);
nor U34538 (N_34538,N_27321,N_23727);
or U34539 (N_34539,N_22251,N_20578);
and U34540 (N_34540,N_20696,N_24980);
and U34541 (N_34541,N_28100,N_23094);
or U34542 (N_34542,N_20365,N_26715);
and U34543 (N_34543,N_22937,N_23158);
xnor U34544 (N_34544,N_26658,N_23792);
nor U34545 (N_34545,N_23582,N_26122);
nand U34546 (N_34546,N_29602,N_27340);
or U34547 (N_34547,N_21397,N_25067);
and U34548 (N_34548,N_26516,N_22413);
nand U34549 (N_34549,N_22557,N_28582);
nand U34550 (N_34550,N_23447,N_23437);
nand U34551 (N_34551,N_22165,N_25482);
xor U34552 (N_34552,N_20256,N_27773);
or U34553 (N_34553,N_25592,N_26523);
or U34554 (N_34554,N_22925,N_25320);
nor U34555 (N_34555,N_27290,N_25516);
nand U34556 (N_34556,N_27177,N_29313);
xnor U34557 (N_34557,N_22490,N_23341);
xnor U34558 (N_34558,N_23555,N_21717);
nand U34559 (N_34559,N_22289,N_23886);
xnor U34560 (N_34560,N_26663,N_29124);
nor U34561 (N_34561,N_28785,N_27823);
xor U34562 (N_34562,N_25814,N_23994);
nand U34563 (N_34563,N_27009,N_28076);
nor U34564 (N_34564,N_22033,N_21528);
xnor U34565 (N_34565,N_25458,N_21973);
or U34566 (N_34566,N_24605,N_29039);
nor U34567 (N_34567,N_24939,N_28973);
nand U34568 (N_34568,N_27978,N_23808);
and U34569 (N_34569,N_23055,N_28197);
and U34570 (N_34570,N_26660,N_25690);
and U34571 (N_34571,N_28007,N_20605);
nor U34572 (N_34572,N_24791,N_26698);
and U34573 (N_34573,N_26273,N_20739);
and U34574 (N_34574,N_22011,N_23549);
nor U34575 (N_34575,N_26187,N_27918);
and U34576 (N_34576,N_27907,N_24405);
and U34577 (N_34577,N_26962,N_27166);
nor U34578 (N_34578,N_26451,N_29314);
nand U34579 (N_34579,N_27753,N_29011);
xnor U34580 (N_34580,N_24307,N_24424);
and U34581 (N_34581,N_25170,N_26284);
nor U34582 (N_34582,N_26301,N_24855);
nand U34583 (N_34583,N_25791,N_28434);
nor U34584 (N_34584,N_26257,N_28846);
nor U34585 (N_34585,N_25017,N_21171);
nor U34586 (N_34586,N_22854,N_29410);
and U34587 (N_34587,N_25244,N_28545);
nor U34588 (N_34588,N_20691,N_28319);
and U34589 (N_34589,N_23198,N_22190);
xor U34590 (N_34590,N_27425,N_28668);
xnor U34591 (N_34591,N_28576,N_29405);
nand U34592 (N_34592,N_24703,N_24516);
xor U34593 (N_34593,N_22686,N_26132);
nor U34594 (N_34594,N_23616,N_25164);
or U34595 (N_34595,N_28401,N_29943);
nor U34596 (N_34596,N_22089,N_28243);
and U34597 (N_34597,N_20965,N_28621);
or U34598 (N_34598,N_29489,N_23211);
and U34599 (N_34599,N_25361,N_21359);
xnor U34600 (N_34600,N_20200,N_25023);
nor U34601 (N_34601,N_20841,N_28677);
and U34602 (N_34602,N_25509,N_25545);
nor U34603 (N_34603,N_24945,N_26823);
nor U34604 (N_34604,N_27034,N_29094);
or U34605 (N_34605,N_26040,N_26999);
or U34606 (N_34606,N_29181,N_21623);
nor U34607 (N_34607,N_20513,N_29069);
nand U34608 (N_34608,N_29149,N_29351);
or U34609 (N_34609,N_28198,N_28497);
nor U34610 (N_34610,N_25727,N_24247);
xor U34611 (N_34611,N_29701,N_28802);
xnor U34612 (N_34612,N_24459,N_25365);
xor U34613 (N_34613,N_20308,N_28055);
nand U34614 (N_34614,N_22160,N_29268);
nand U34615 (N_34615,N_25614,N_29909);
or U34616 (N_34616,N_24757,N_26401);
or U34617 (N_34617,N_27921,N_27566);
nor U34618 (N_34618,N_25718,N_22918);
xor U34619 (N_34619,N_27802,N_27772);
xor U34620 (N_34620,N_27709,N_21999);
or U34621 (N_34621,N_23008,N_21213);
and U34622 (N_34622,N_27136,N_27077);
nand U34623 (N_34623,N_29140,N_21699);
nand U34624 (N_34624,N_29241,N_20847);
nand U34625 (N_34625,N_20375,N_26527);
nand U34626 (N_34626,N_22555,N_20021);
nor U34627 (N_34627,N_24692,N_20456);
xnor U34628 (N_34628,N_28385,N_26006);
nand U34629 (N_34629,N_28040,N_20138);
nor U34630 (N_34630,N_23082,N_25853);
and U34631 (N_34631,N_24357,N_26205);
or U34632 (N_34632,N_28964,N_22608);
xor U34633 (N_34633,N_23309,N_26011);
nand U34634 (N_34634,N_29494,N_24173);
nor U34635 (N_34635,N_27446,N_29635);
xor U34636 (N_34636,N_27501,N_24526);
nand U34637 (N_34637,N_20386,N_20581);
or U34638 (N_34638,N_23486,N_28462);
or U34639 (N_34639,N_23757,N_21747);
xnor U34640 (N_34640,N_23545,N_25169);
xnor U34641 (N_34641,N_25710,N_28356);
xor U34642 (N_34642,N_21755,N_25635);
nor U34643 (N_34643,N_20061,N_28209);
nor U34644 (N_34644,N_22653,N_27427);
xor U34645 (N_34645,N_25078,N_22658);
nand U34646 (N_34646,N_21798,N_20289);
nor U34647 (N_34647,N_22893,N_25028);
and U34648 (N_34648,N_21899,N_25960);
nand U34649 (N_34649,N_25518,N_22355);
or U34650 (N_34650,N_28966,N_21926);
xnor U34651 (N_34651,N_28688,N_28731);
or U34652 (N_34652,N_22094,N_27599);
xnor U34653 (N_34653,N_29747,N_29193);
nor U34654 (N_34654,N_21918,N_27804);
and U34655 (N_34655,N_22376,N_25449);
or U34656 (N_34656,N_25110,N_21890);
or U34657 (N_34657,N_27924,N_25965);
or U34658 (N_34658,N_28188,N_22926);
or U34659 (N_34659,N_24785,N_29932);
and U34660 (N_34660,N_23590,N_23585);
nand U34661 (N_34661,N_25185,N_20435);
nand U34662 (N_34662,N_26098,N_26244);
and U34663 (N_34663,N_21384,N_20405);
xnor U34664 (N_34664,N_23588,N_25634);
nor U34665 (N_34665,N_22536,N_25980);
nand U34666 (N_34666,N_27700,N_28806);
nand U34667 (N_34667,N_26848,N_23766);
nor U34668 (N_34668,N_28961,N_21920);
xor U34669 (N_34669,N_28714,N_21675);
and U34670 (N_34670,N_23578,N_22884);
and U34671 (N_34671,N_27070,N_23580);
nor U34672 (N_34672,N_20074,N_25722);
or U34673 (N_34673,N_21029,N_23524);
nor U34674 (N_34674,N_20918,N_27413);
nand U34675 (N_34675,N_22616,N_24707);
and U34676 (N_34676,N_27905,N_21784);
and U34677 (N_34677,N_24128,N_24604);
and U34678 (N_34678,N_24107,N_25741);
or U34679 (N_34679,N_20506,N_26802);
nor U34680 (N_34680,N_27747,N_26620);
nor U34681 (N_34681,N_25135,N_22784);
and U34682 (N_34682,N_25381,N_29583);
nand U34683 (N_34683,N_27337,N_27419);
xor U34684 (N_34684,N_22404,N_29137);
nor U34685 (N_34685,N_25664,N_29192);
nand U34686 (N_34686,N_27401,N_23075);
xnor U34687 (N_34687,N_28499,N_20342);
nand U34688 (N_34688,N_27845,N_26553);
or U34689 (N_34689,N_21370,N_21218);
xor U34690 (N_34690,N_29171,N_28060);
and U34691 (N_34691,N_24480,N_29967);
and U34692 (N_34692,N_21657,N_22840);
xnor U34693 (N_34693,N_28595,N_28739);
nor U34694 (N_34694,N_21562,N_23547);
nand U34695 (N_34695,N_22127,N_22474);
nor U34696 (N_34696,N_20657,N_29890);
and U34697 (N_34697,N_23712,N_29698);
and U34698 (N_34698,N_22118,N_22908);
nor U34699 (N_34699,N_21783,N_26422);
or U34700 (N_34700,N_28323,N_23972);
and U34701 (N_34701,N_23425,N_22752);
nor U34702 (N_34702,N_26347,N_26198);
xor U34703 (N_34703,N_22283,N_29505);
and U34704 (N_34704,N_21471,N_24749);
or U34705 (N_34705,N_28052,N_20795);
nor U34706 (N_34706,N_24817,N_22304);
and U34707 (N_34707,N_22318,N_25725);
nor U34708 (N_34708,N_23175,N_28241);
nand U34709 (N_34709,N_29367,N_23205);
or U34710 (N_34710,N_27370,N_24003);
nor U34711 (N_34711,N_20775,N_21024);
nand U34712 (N_34712,N_22395,N_21200);
nor U34713 (N_34713,N_23905,N_28940);
nor U34714 (N_34714,N_25118,N_25311);
nand U34715 (N_34715,N_27903,N_20129);
xnor U34716 (N_34716,N_29131,N_21475);
or U34717 (N_34717,N_24118,N_22768);
xnor U34718 (N_34718,N_21022,N_25032);
nor U34719 (N_34719,N_24502,N_27302);
xor U34720 (N_34720,N_29182,N_26296);
nand U34721 (N_34721,N_27493,N_23642);
and U34722 (N_34722,N_20197,N_26089);
and U34723 (N_34723,N_25571,N_26899);
nor U34724 (N_34724,N_21826,N_22703);
and U34725 (N_34725,N_23174,N_28439);
or U34726 (N_34726,N_28518,N_22734);
nor U34727 (N_34727,N_27381,N_28106);
nand U34728 (N_34728,N_27797,N_26927);
xnor U34729 (N_34729,N_21635,N_22350);
or U34730 (N_34730,N_23618,N_23587);
xnor U34731 (N_34731,N_24509,N_25881);
or U34732 (N_34732,N_22080,N_21166);
or U34733 (N_34733,N_29617,N_23050);
nand U34734 (N_34734,N_21383,N_28737);
or U34735 (N_34735,N_23614,N_27374);
nand U34736 (N_34736,N_29027,N_20428);
or U34737 (N_34737,N_24287,N_25080);
and U34738 (N_34738,N_20674,N_21976);
and U34739 (N_34739,N_20681,N_23561);
or U34740 (N_34740,N_23463,N_21273);
nand U34741 (N_34741,N_20330,N_23326);
and U34742 (N_34742,N_23667,N_21456);
nor U34743 (N_34743,N_26923,N_25904);
or U34744 (N_34744,N_21441,N_29843);
xor U34745 (N_34745,N_26829,N_23746);
nor U34746 (N_34746,N_24609,N_22972);
nor U34747 (N_34747,N_26503,N_26103);
nand U34748 (N_34748,N_20986,N_27878);
nor U34749 (N_34749,N_24081,N_22442);
or U34750 (N_34750,N_27218,N_26851);
or U34751 (N_34751,N_24056,N_24536);
nor U34752 (N_34752,N_21187,N_21072);
nor U34753 (N_34753,N_20340,N_28610);
or U34754 (N_34754,N_28467,N_20692);
nand U34755 (N_34755,N_23571,N_28923);
nor U34756 (N_34756,N_22668,N_21407);
xnor U34757 (N_34757,N_27778,N_22636);
nand U34758 (N_34758,N_28114,N_25523);
or U34759 (N_34759,N_23630,N_24364);
xor U34760 (N_34760,N_26852,N_20995);
or U34761 (N_34761,N_27947,N_24592);
xor U34762 (N_34762,N_28982,N_27300);
and U34763 (N_34763,N_26783,N_24304);
nor U34764 (N_34764,N_28210,N_25695);
or U34765 (N_34765,N_27360,N_20537);
nand U34766 (N_34766,N_25792,N_29031);
xor U34767 (N_34767,N_23677,N_24575);
and U34768 (N_34768,N_20067,N_25233);
and U34769 (N_34769,N_29089,N_25406);
and U34770 (N_34770,N_21907,N_20776);
xor U34771 (N_34771,N_23546,N_27581);
xor U34772 (N_34772,N_24629,N_27630);
nor U34773 (N_34773,N_29645,N_25754);
or U34774 (N_34774,N_26070,N_22928);
and U34775 (N_34775,N_28741,N_28716);
xnor U34776 (N_34776,N_23751,N_26943);
xnor U34777 (N_34777,N_23846,N_23803);
and U34778 (N_34778,N_24193,N_27285);
nor U34779 (N_34779,N_26237,N_27792);
and U34780 (N_34780,N_22431,N_29308);
or U34781 (N_34781,N_22049,N_22495);
or U34782 (N_34782,N_22534,N_27962);
nor U34783 (N_34783,N_24014,N_26915);
or U34784 (N_34784,N_22874,N_26300);
nor U34785 (N_34785,N_24029,N_27762);
nand U34786 (N_34786,N_20323,N_20783);
nand U34787 (N_34787,N_22946,N_21194);
nand U34788 (N_34788,N_21042,N_29113);
nand U34789 (N_34789,N_22496,N_21849);
or U34790 (N_34790,N_28085,N_28091);
and U34791 (N_34791,N_28682,N_24141);
or U34792 (N_34792,N_26066,N_27245);
or U34793 (N_34793,N_23216,N_24708);
xor U34794 (N_34794,N_22366,N_21236);
or U34795 (N_34795,N_26350,N_25794);
nor U34796 (N_34796,N_24870,N_21902);
xor U34797 (N_34797,N_22858,N_23264);
or U34798 (N_34798,N_25839,N_28312);
and U34799 (N_34799,N_26123,N_27694);
nand U34800 (N_34800,N_27058,N_22700);
nand U34801 (N_34801,N_29526,N_23440);
xnor U34802 (N_34802,N_20257,N_27478);
xnor U34803 (N_34803,N_25593,N_22311);
xnor U34804 (N_34804,N_20058,N_28273);
and U34805 (N_34805,N_29437,N_23257);
nand U34806 (N_34806,N_28005,N_21207);
and U34807 (N_34807,N_29291,N_28179);
nand U34808 (N_34808,N_27270,N_26427);
and U34809 (N_34809,N_26327,N_29925);
and U34810 (N_34810,N_28718,N_23827);
nor U34811 (N_34811,N_20486,N_28607);
nand U34812 (N_34812,N_27742,N_20132);
and U34813 (N_34813,N_25100,N_29153);
or U34814 (N_34814,N_29542,N_20688);
xnor U34815 (N_34815,N_20262,N_27761);
nand U34816 (N_34816,N_26464,N_29186);
nand U34817 (N_34817,N_23368,N_21173);
xor U34818 (N_34818,N_24724,N_29199);
and U34819 (N_34819,N_22050,N_21991);
xnor U34820 (N_34820,N_28868,N_26058);
nor U34821 (N_34821,N_23532,N_20988);
nor U34822 (N_34822,N_22520,N_21487);
nand U34823 (N_34823,N_29014,N_22539);
and U34824 (N_34824,N_25949,N_28847);
or U34825 (N_34825,N_28332,N_29254);
and U34826 (N_34826,N_29161,N_24457);
nand U34827 (N_34827,N_24413,N_28548);
nor U34828 (N_34828,N_20192,N_24059);
or U34829 (N_34829,N_23615,N_29590);
or U34830 (N_34830,N_21226,N_27885);
and U34831 (N_34831,N_26172,N_21157);
and U34832 (N_34832,N_22063,N_26341);
nand U34833 (N_34833,N_22994,N_27669);
nor U34834 (N_34834,N_29391,N_23168);
or U34835 (N_34835,N_29525,N_28636);
xnor U34836 (N_34836,N_29251,N_21392);
and U34837 (N_34837,N_27196,N_22560);
nor U34838 (N_34838,N_28656,N_25981);
nand U34839 (N_34839,N_25831,N_22915);
nor U34840 (N_34840,N_20301,N_26157);
xor U34841 (N_34841,N_25389,N_23921);
nor U34842 (N_34842,N_27941,N_27665);
nand U34843 (N_34843,N_25734,N_24891);
or U34844 (N_34844,N_26255,N_21212);
or U34845 (N_34845,N_21648,N_25586);
and U34846 (N_34846,N_27879,N_21349);
or U34847 (N_34847,N_28715,N_20394);
or U34848 (N_34848,N_27132,N_29852);
nand U34849 (N_34849,N_25872,N_24904);
xor U34850 (N_34850,N_20801,N_22983);
or U34851 (N_34851,N_22377,N_21100);
nand U34852 (N_34852,N_29054,N_25285);
nor U34853 (N_34853,N_20072,N_28226);
nand U34854 (N_34854,N_25411,N_26334);
xor U34855 (N_34855,N_26275,N_20134);
nor U34856 (N_34856,N_25367,N_26521);
nand U34857 (N_34857,N_24430,N_23496);
nor U34858 (N_34858,N_22866,N_23336);
or U34859 (N_34859,N_28274,N_20259);
xnor U34860 (N_34860,N_25543,N_22591);
or U34861 (N_34861,N_24115,N_26152);
xor U34862 (N_34862,N_22742,N_24538);
and U34863 (N_34863,N_20968,N_24941);
nand U34864 (N_34864,N_24360,N_21214);
or U34865 (N_34865,N_27326,N_24975);
xnor U34866 (N_34866,N_22860,N_20267);
and U34867 (N_34867,N_29746,N_23992);
or U34868 (N_34868,N_27916,N_24008);
and U34869 (N_34869,N_27569,N_25488);
xnor U34870 (N_34870,N_29980,N_25730);
and U34871 (N_34871,N_22206,N_25238);
or U34872 (N_34872,N_23901,N_23289);
nor U34873 (N_34873,N_23919,N_28357);
or U34874 (N_34874,N_22268,N_26606);
xor U34875 (N_34875,N_27051,N_20762);
nand U34876 (N_34876,N_29598,N_22945);
xor U34877 (N_34877,N_21704,N_29396);
and U34878 (N_34878,N_21303,N_20064);
xor U34879 (N_34879,N_21062,N_20232);
nor U34880 (N_34880,N_23306,N_28917);
and U34881 (N_34881,N_29928,N_28824);
nand U34882 (N_34882,N_21248,N_25334);
xor U34883 (N_34883,N_20381,N_21681);
or U34884 (N_34884,N_29828,N_29734);
xor U34885 (N_34885,N_22030,N_23874);
nand U34886 (N_34886,N_28678,N_25245);
or U34887 (N_34887,N_25336,N_20730);
xnor U34888 (N_34888,N_21144,N_27587);
nor U34889 (N_34889,N_26024,N_22475);
or U34890 (N_34890,N_20271,N_28425);
nor U34891 (N_34891,N_20612,N_26197);
and U34892 (N_34892,N_26500,N_28242);
xor U34893 (N_34893,N_28791,N_23798);
xnor U34894 (N_34894,N_28108,N_25542);
nand U34895 (N_34895,N_22146,N_22863);
nand U34896 (N_34896,N_27238,N_25642);
nor U34897 (N_34897,N_21825,N_27021);
nand U34898 (N_34898,N_22864,N_25407);
nand U34899 (N_34899,N_23907,N_20913);
or U34900 (N_34900,N_25125,N_27364);
xor U34901 (N_34901,N_26581,N_25111);
and U34902 (N_34902,N_22006,N_24753);
xnor U34903 (N_34903,N_23409,N_26195);
and U34904 (N_34904,N_23137,N_21538);
xnor U34905 (N_34905,N_22047,N_28906);
nand U34906 (N_34906,N_24696,N_24921);
nand U34907 (N_34907,N_21116,N_29885);
xnor U34908 (N_34908,N_21006,N_22077);
xnor U34909 (N_34909,N_27015,N_27174);
nand U34910 (N_34910,N_25913,N_25953);
nor U34911 (N_34911,N_28579,N_25338);
nand U34912 (N_34912,N_20477,N_24889);
nand U34913 (N_34913,N_24211,N_24543);
xor U34914 (N_34914,N_20278,N_25128);
nand U34915 (N_34915,N_26491,N_22280);
xnor U34916 (N_34916,N_26023,N_27740);
xnor U34917 (N_34917,N_27027,N_24440);
xor U34918 (N_34918,N_20648,N_27447);
nor U34919 (N_34919,N_23144,N_27714);
nor U34920 (N_34920,N_29835,N_21577);
nand U34921 (N_34921,N_27736,N_26332);
nor U34922 (N_34922,N_21135,N_20295);
xnor U34923 (N_34923,N_23814,N_27582);
and U34924 (N_34924,N_28608,N_20250);
and U34925 (N_34925,N_20926,N_29687);
nor U34926 (N_34926,N_27652,N_27133);
nand U34927 (N_34927,N_27056,N_24840);
xor U34928 (N_34928,N_24181,N_22142);
nand U34929 (N_34929,N_20466,N_28450);
nand U34930 (N_34930,N_22415,N_29259);
nor U34931 (N_34931,N_24018,N_23641);
or U34932 (N_34932,N_24474,N_28635);
xnor U34933 (N_34933,N_20016,N_23351);
xor U34934 (N_34934,N_27258,N_20676);
and U34935 (N_34935,N_20469,N_23525);
or U34936 (N_34936,N_27065,N_28384);
nand U34937 (N_34937,N_21496,N_22977);
and U34938 (N_34938,N_24738,N_25424);
or U34939 (N_34939,N_21371,N_28256);
or U34940 (N_34940,N_21604,N_22097);
nand U34941 (N_34941,N_26492,N_25677);
and U34942 (N_34942,N_27889,N_23644);
or U34943 (N_34943,N_25637,N_28615);
nor U34944 (N_34944,N_26060,N_25519);
or U34945 (N_34945,N_20697,N_22130);
nor U34946 (N_34946,N_26910,N_26593);
nor U34947 (N_34947,N_23081,N_27639);
xor U34948 (N_34948,N_25265,N_26085);
and U34949 (N_34949,N_27783,N_29663);
nor U34950 (N_34950,N_28059,N_24096);
nor U34951 (N_34951,N_20194,N_26045);
nor U34952 (N_34952,N_21436,N_27308);
and U34953 (N_34953,N_25487,N_26297);
nor U34954 (N_34954,N_28622,N_24471);
nor U34955 (N_34955,N_23802,N_21499);
and U34956 (N_34956,N_26796,N_23518);
nor U34957 (N_34957,N_20756,N_23276);
xor U34958 (N_34958,N_28971,N_29737);
xnor U34959 (N_34959,N_28914,N_24372);
and U34960 (N_34960,N_28735,N_21987);
nor U34961 (N_34961,N_24722,N_29353);
nand U34962 (N_34962,N_21282,N_29854);
nand U34963 (N_34963,N_28147,N_23510);
xor U34964 (N_34964,N_28104,N_20018);
and U34965 (N_34965,N_24310,N_21504);
xnor U34966 (N_34966,N_24256,N_24213);
and U34967 (N_34967,N_20427,N_28747);
xnor U34968 (N_34968,N_29722,N_26542);
xor U34969 (N_34969,N_24803,N_23478);
nand U34970 (N_34970,N_20931,N_20933);
and U34971 (N_34971,N_24432,N_27664);
nor U34972 (N_34972,N_21678,N_24908);
or U34973 (N_34973,N_22279,N_20658);
nor U34974 (N_34974,N_22685,N_29300);
xor U34975 (N_34975,N_20269,N_22288);
and U34976 (N_34976,N_22911,N_28025);
and U34977 (N_34977,N_24052,N_29581);
and U34978 (N_34978,N_22980,N_29090);
xnor U34979 (N_34979,N_27909,N_27510);
or U34980 (N_34980,N_24194,N_20176);
or U34981 (N_34981,N_24397,N_27053);
or U34982 (N_34982,N_24016,N_29400);
and U34983 (N_34983,N_29850,N_22121);
xor U34984 (N_34984,N_29195,N_24283);
nand U34985 (N_34985,N_23381,N_22325);
and U34986 (N_34986,N_27650,N_24156);
and U34987 (N_34987,N_28880,N_21884);
nor U34988 (N_34988,N_25943,N_20854);
and U34989 (N_34989,N_27243,N_21292);
and U34990 (N_34990,N_29729,N_22398);
nor U34991 (N_34991,N_22481,N_27873);
nor U34992 (N_34992,N_28924,N_20843);
or U34993 (N_34993,N_29669,N_27494);
xor U34994 (N_34994,N_25154,N_23986);
nand U34995 (N_34995,N_28410,N_21650);
and U34996 (N_34996,N_26967,N_24445);
and U34997 (N_34997,N_22448,N_25054);
or U34998 (N_34998,N_22861,N_29416);
and U34999 (N_34999,N_29252,N_28916);
xor U35000 (N_35000,N_29209,N_23273);
or U35001 (N_35001,N_20317,N_25005);
or U35002 (N_35002,N_26079,N_21256);
nor U35003 (N_35003,N_22292,N_24088);
nor U35004 (N_35004,N_20737,N_20817);
xor U35005 (N_35005,N_21830,N_29096);
xor U35006 (N_35006,N_28722,N_25074);
or U35007 (N_35007,N_24602,N_22103);
nor U35008 (N_35008,N_22739,N_21808);
nor U35009 (N_35009,N_24147,N_28047);
or U35010 (N_35010,N_27266,N_20356);
or U35011 (N_35011,N_28305,N_24623);
or U35012 (N_35012,N_23970,N_26879);
and U35013 (N_35013,N_25505,N_20063);
xnor U35014 (N_35014,N_27623,N_20097);
xnor U35015 (N_35015,N_23483,N_29067);
and U35016 (N_35016,N_22178,N_29409);
or U35017 (N_35017,N_29510,N_25675);
nor U35018 (N_35018,N_20194,N_23341);
nor U35019 (N_35019,N_20093,N_21287);
nand U35020 (N_35020,N_29340,N_23858);
or U35021 (N_35021,N_20054,N_27133);
nor U35022 (N_35022,N_23333,N_24955);
and U35023 (N_35023,N_26516,N_25704);
nand U35024 (N_35024,N_27422,N_22253);
xor U35025 (N_35025,N_23572,N_25300);
and U35026 (N_35026,N_24946,N_27901);
and U35027 (N_35027,N_24873,N_22781);
xor U35028 (N_35028,N_29444,N_25948);
nor U35029 (N_35029,N_21880,N_29668);
or U35030 (N_35030,N_22175,N_29586);
xor U35031 (N_35031,N_29934,N_29993);
or U35032 (N_35032,N_29208,N_20095);
xor U35033 (N_35033,N_29641,N_28806);
xnor U35034 (N_35034,N_26954,N_22755);
nor U35035 (N_35035,N_27864,N_29338);
or U35036 (N_35036,N_27295,N_23428);
nor U35037 (N_35037,N_24497,N_27618);
xnor U35038 (N_35038,N_24236,N_22770);
or U35039 (N_35039,N_23726,N_27426);
or U35040 (N_35040,N_20939,N_25239);
nor U35041 (N_35041,N_23269,N_21533);
nand U35042 (N_35042,N_26903,N_27937);
and U35043 (N_35043,N_25164,N_20388);
or U35044 (N_35044,N_22494,N_20645);
nor U35045 (N_35045,N_23448,N_23832);
and U35046 (N_35046,N_23780,N_29144);
or U35047 (N_35047,N_25220,N_22395);
or U35048 (N_35048,N_29009,N_25221);
and U35049 (N_35049,N_25966,N_21137);
and U35050 (N_35050,N_24158,N_20715);
nor U35051 (N_35051,N_23925,N_23694);
nor U35052 (N_35052,N_22034,N_23631);
nand U35053 (N_35053,N_21356,N_24397);
or U35054 (N_35054,N_25612,N_21486);
nor U35055 (N_35055,N_20246,N_28809);
and U35056 (N_35056,N_20539,N_26113);
or U35057 (N_35057,N_28539,N_26799);
xor U35058 (N_35058,N_20905,N_24169);
nor U35059 (N_35059,N_28748,N_27101);
xnor U35060 (N_35060,N_23457,N_27114);
and U35061 (N_35061,N_24900,N_25718);
nand U35062 (N_35062,N_28257,N_27691);
xnor U35063 (N_35063,N_20517,N_24903);
xor U35064 (N_35064,N_22236,N_22395);
xnor U35065 (N_35065,N_22778,N_21657);
xnor U35066 (N_35066,N_24491,N_22787);
and U35067 (N_35067,N_24896,N_26151);
and U35068 (N_35068,N_20024,N_29968);
and U35069 (N_35069,N_26900,N_27382);
xnor U35070 (N_35070,N_25214,N_26480);
nand U35071 (N_35071,N_28636,N_27378);
nand U35072 (N_35072,N_22905,N_22568);
nand U35073 (N_35073,N_24711,N_21693);
xnor U35074 (N_35074,N_28606,N_25514);
xor U35075 (N_35075,N_24693,N_22099);
and U35076 (N_35076,N_22001,N_27199);
xnor U35077 (N_35077,N_23017,N_26124);
nor U35078 (N_35078,N_29880,N_24531);
and U35079 (N_35079,N_23576,N_21411);
xnor U35080 (N_35080,N_21591,N_28044);
or U35081 (N_35081,N_25398,N_29705);
and U35082 (N_35082,N_26729,N_23511);
xnor U35083 (N_35083,N_23066,N_24234);
xnor U35084 (N_35084,N_21164,N_21930);
nor U35085 (N_35085,N_20538,N_28685);
xnor U35086 (N_35086,N_24072,N_27762);
nor U35087 (N_35087,N_27675,N_26246);
xor U35088 (N_35088,N_27549,N_21924);
or U35089 (N_35089,N_23484,N_20039);
nand U35090 (N_35090,N_23875,N_24789);
nor U35091 (N_35091,N_28296,N_21160);
nor U35092 (N_35092,N_22831,N_24212);
xnor U35093 (N_35093,N_25130,N_23678);
xnor U35094 (N_35094,N_21662,N_28081);
nor U35095 (N_35095,N_26582,N_23768);
or U35096 (N_35096,N_26180,N_24196);
and U35097 (N_35097,N_29677,N_23104);
nand U35098 (N_35098,N_24786,N_25741);
or U35099 (N_35099,N_21008,N_27111);
xor U35100 (N_35100,N_21572,N_23498);
xnor U35101 (N_35101,N_26112,N_24712);
nand U35102 (N_35102,N_28121,N_29262);
nand U35103 (N_35103,N_21225,N_28791);
and U35104 (N_35104,N_26453,N_20626);
nand U35105 (N_35105,N_20446,N_29410);
and U35106 (N_35106,N_22122,N_23494);
nor U35107 (N_35107,N_28038,N_21747);
or U35108 (N_35108,N_25798,N_22482);
or U35109 (N_35109,N_29322,N_27448);
and U35110 (N_35110,N_28970,N_21217);
xor U35111 (N_35111,N_21376,N_27851);
xor U35112 (N_35112,N_21553,N_28926);
xor U35113 (N_35113,N_20237,N_29994);
nor U35114 (N_35114,N_29225,N_22748);
nor U35115 (N_35115,N_22609,N_23455);
nand U35116 (N_35116,N_26042,N_21433);
and U35117 (N_35117,N_22638,N_27708);
and U35118 (N_35118,N_22678,N_29402);
or U35119 (N_35119,N_22875,N_26976);
and U35120 (N_35120,N_22335,N_26111);
xor U35121 (N_35121,N_21117,N_25185);
xnor U35122 (N_35122,N_27274,N_23565);
nor U35123 (N_35123,N_25392,N_21326);
or U35124 (N_35124,N_29775,N_23249);
nor U35125 (N_35125,N_23935,N_21702);
xor U35126 (N_35126,N_25036,N_29755);
xor U35127 (N_35127,N_20138,N_22096);
nand U35128 (N_35128,N_29526,N_27059);
or U35129 (N_35129,N_25983,N_22365);
or U35130 (N_35130,N_29893,N_28933);
nor U35131 (N_35131,N_20626,N_28548);
or U35132 (N_35132,N_20381,N_20008);
xnor U35133 (N_35133,N_21766,N_27969);
nor U35134 (N_35134,N_26129,N_28208);
nand U35135 (N_35135,N_22738,N_28791);
nand U35136 (N_35136,N_26816,N_23507);
xor U35137 (N_35137,N_28101,N_26743);
nor U35138 (N_35138,N_21091,N_29282);
nor U35139 (N_35139,N_20355,N_25491);
nand U35140 (N_35140,N_28125,N_21892);
nor U35141 (N_35141,N_27443,N_24555);
nor U35142 (N_35142,N_27039,N_25076);
nand U35143 (N_35143,N_21275,N_20390);
and U35144 (N_35144,N_21116,N_29034);
or U35145 (N_35145,N_21389,N_25876);
or U35146 (N_35146,N_21632,N_20811);
nor U35147 (N_35147,N_29879,N_29890);
nor U35148 (N_35148,N_20965,N_22255);
xor U35149 (N_35149,N_20452,N_28516);
and U35150 (N_35150,N_20131,N_21188);
nand U35151 (N_35151,N_23837,N_24757);
xor U35152 (N_35152,N_20581,N_26501);
nand U35153 (N_35153,N_24373,N_23002);
and U35154 (N_35154,N_24623,N_23082);
and U35155 (N_35155,N_27102,N_26567);
or U35156 (N_35156,N_21705,N_21452);
xnor U35157 (N_35157,N_29573,N_22114);
nor U35158 (N_35158,N_27028,N_26868);
xor U35159 (N_35159,N_25338,N_24832);
or U35160 (N_35160,N_29297,N_22825);
nor U35161 (N_35161,N_23727,N_26626);
or U35162 (N_35162,N_27887,N_23520);
or U35163 (N_35163,N_24081,N_28588);
nand U35164 (N_35164,N_27457,N_29070);
and U35165 (N_35165,N_25776,N_22284);
and U35166 (N_35166,N_27158,N_28719);
xor U35167 (N_35167,N_29695,N_28600);
and U35168 (N_35168,N_28634,N_23198);
nand U35169 (N_35169,N_22647,N_27981);
and U35170 (N_35170,N_23896,N_28149);
or U35171 (N_35171,N_22436,N_26017);
or U35172 (N_35172,N_20422,N_29113);
and U35173 (N_35173,N_23958,N_21033);
and U35174 (N_35174,N_21504,N_25525);
nor U35175 (N_35175,N_28910,N_21720);
and U35176 (N_35176,N_24892,N_23275);
xnor U35177 (N_35177,N_24997,N_23100);
xor U35178 (N_35178,N_29195,N_27966);
and U35179 (N_35179,N_20296,N_27062);
and U35180 (N_35180,N_21824,N_27953);
nor U35181 (N_35181,N_28387,N_25787);
nand U35182 (N_35182,N_24892,N_21732);
nand U35183 (N_35183,N_20225,N_24541);
and U35184 (N_35184,N_28621,N_29300);
nor U35185 (N_35185,N_29083,N_22632);
nand U35186 (N_35186,N_27598,N_26991);
xor U35187 (N_35187,N_27389,N_22857);
nand U35188 (N_35188,N_29775,N_29553);
nand U35189 (N_35189,N_21685,N_22072);
nor U35190 (N_35190,N_27447,N_25970);
and U35191 (N_35191,N_23356,N_25821);
and U35192 (N_35192,N_27107,N_22621);
nand U35193 (N_35193,N_23440,N_21805);
nand U35194 (N_35194,N_23337,N_29765);
nor U35195 (N_35195,N_22982,N_29639);
or U35196 (N_35196,N_29188,N_28448);
nand U35197 (N_35197,N_20103,N_24439);
xor U35198 (N_35198,N_27686,N_28827);
nand U35199 (N_35199,N_20553,N_24632);
xnor U35200 (N_35200,N_23008,N_22502);
nor U35201 (N_35201,N_28437,N_28069);
and U35202 (N_35202,N_20366,N_22926);
or U35203 (N_35203,N_25286,N_28049);
or U35204 (N_35204,N_21324,N_25188);
nor U35205 (N_35205,N_27592,N_23301);
and U35206 (N_35206,N_25018,N_29880);
xnor U35207 (N_35207,N_24378,N_25610);
nor U35208 (N_35208,N_27359,N_25839);
nor U35209 (N_35209,N_20203,N_22463);
nor U35210 (N_35210,N_23311,N_25426);
xnor U35211 (N_35211,N_28093,N_22299);
nand U35212 (N_35212,N_25932,N_21393);
nand U35213 (N_35213,N_28996,N_22990);
nand U35214 (N_35214,N_29336,N_25874);
or U35215 (N_35215,N_27230,N_23007);
and U35216 (N_35216,N_20512,N_21212);
nand U35217 (N_35217,N_26804,N_24413);
or U35218 (N_35218,N_22152,N_20186);
xnor U35219 (N_35219,N_21092,N_20743);
xor U35220 (N_35220,N_23620,N_23052);
and U35221 (N_35221,N_20144,N_25939);
and U35222 (N_35222,N_29664,N_28295);
or U35223 (N_35223,N_22222,N_28429);
nor U35224 (N_35224,N_21613,N_21542);
nand U35225 (N_35225,N_24138,N_27526);
or U35226 (N_35226,N_23710,N_23125);
xnor U35227 (N_35227,N_22336,N_24733);
or U35228 (N_35228,N_20425,N_28804);
nand U35229 (N_35229,N_29054,N_29871);
and U35230 (N_35230,N_21284,N_21311);
nand U35231 (N_35231,N_24913,N_23343);
nor U35232 (N_35232,N_25608,N_21454);
nand U35233 (N_35233,N_20041,N_22536);
xor U35234 (N_35234,N_22348,N_20844);
and U35235 (N_35235,N_20529,N_29708);
nor U35236 (N_35236,N_23312,N_28773);
xor U35237 (N_35237,N_20092,N_27283);
xor U35238 (N_35238,N_25248,N_25909);
and U35239 (N_35239,N_23408,N_22076);
or U35240 (N_35240,N_23115,N_28766);
and U35241 (N_35241,N_27076,N_23819);
and U35242 (N_35242,N_22574,N_22734);
or U35243 (N_35243,N_27978,N_26473);
or U35244 (N_35244,N_25582,N_21722);
or U35245 (N_35245,N_20705,N_28021);
and U35246 (N_35246,N_20387,N_21077);
and U35247 (N_35247,N_27658,N_23145);
and U35248 (N_35248,N_22548,N_23538);
and U35249 (N_35249,N_22239,N_22719);
xor U35250 (N_35250,N_24891,N_20658);
or U35251 (N_35251,N_25380,N_22888);
and U35252 (N_35252,N_25020,N_22264);
or U35253 (N_35253,N_25842,N_28211);
or U35254 (N_35254,N_26728,N_23062);
nor U35255 (N_35255,N_25075,N_28021);
and U35256 (N_35256,N_22404,N_26993);
and U35257 (N_35257,N_25450,N_22978);
and U35258 (N_35258,N_25992,N_26583);
nor U35259 (N_35259,N_23698,N_23123);
xnor U35260 (N_35260,N_22489,N_21027);
or U35261 (N_35261,N_29563,N_27078);
or U35262 (N_35262,N_24593,N_25339);
xor U35263 (N_35263,N_23641,N_20144);
and U35264 (N_35264,N_24851,N_22661);
nand U35265 (N_35265,N_29594,N_27709);
nor U35266 (N_35266,N_29150,N_29430);
xor U35267 (N_35267,N_29740,N_29609);
nand U35268 (N_35268,N_20707,N_22100);
and U35269 (N_35269,N_22442,N_29576);
and U35270 (N_35270,N_29759,N_27065);
nand U35271 (N_35271,N_25989,N_24240);
and U35272 (N_35272,N_24944,N_23880);
nand U35273 (N_35273,N_21804,N_24634);
nor U35274 (N_35274,N_22300,N_26501);
nand U35275 (N_35275,N_27121,N_23908);
nor U35276 (N_35276,N_23353,N_22318);
nor U35277 (N_35277,N_26142,N_23279);
or U35278 (N_35278,N_27388,N_25498);
nor U35279 (N_35279,N_27536,N_29633);
or U35280 (N_35280,N_29481,N_27887);
or U35281 (N_35281,N_23137,N_23131);
xnor U35282 (N_35282,N_25522,N_24353);
and U35283 (N_35283,N_28205,N_22598);
nand U35284 (N_35284,N_22082,N_22547);
nor U35285 (N_35285,N_26599,N_24047);
xor U35286 (N_35286,N_22836,N_28538);
and U35287 (N_35287,N_22568,N_22273);
or U35288 (N_35288,N_29169,N_20481);
nor U35289 (N_35289,N_22159,N_24764);
and U35290 (N_35290,N_24285,N_20378);
or U35291 (N_35291,N_21509,N_22805);
or U35292 (N_35292,N_28801,N_21725);
nor U35293 (N_35293,N_23388,N_28898);
and U35294 (N_35294,N_21076,N_26578);
nand U35295 (N_35295,N_23101,N_25731);
and U35296 (N_35296,N_25456,N_28889);
nand U35297 (N_35297,N_24475,N_27397);
and U35298 (N_35298,N_22762,N_24306);
xnor U35299 (N_35299,N_26903,N_26423);
and U35300 (N_35300,N_27520,N_25509);
xnor U35301 (N_35301,N_21672,N_21235);
or U35302 (N_35302,N_26870,N_21955);
xnor U35303 (N_35303,N_25131,N_24418);
xnor U35304 (N_35304,N_27393,N_23813);
and U35305 (N_35305,N_23323,N_23953);
and U35306 (N_35306,N_23836,N_24149);
and U35307 (N_35307,N_25487,N_29192);
nor U35308 (N_35308,N_26158,N_27472);
nand U35309 (N_35309,N_26042,N_24226);
nand U35310 (N_35310,N_24517,N_28843);
xnor U35311 (N_35311,N_22934,N_21148);
xnor U35312 (N_35312,N_25134,N_29042);
nand U35313 (N_35313,N_27566,N_29308);
nand U35314 (N_35314,N_24159,N_26873);
nand U35315 (N_35315,N_25145,N_25981);
and U35316 (N_35316,N_28096,N_20951);
and U35317 (N_35317,N_26302,N_27707);
xnor U35318 (N_35318,N_21222,N_24206);
nor U35319 (N_35319,N_27285,N_28266);
nand U35320 (N_35320,N_25843,N_22500);
nor U35321 (N_35321,N_20596,N_26112);
nor U35322 (N_35322,N_21040,N_22729);
or U35323 (N_35323,N_28572,N_21360);
and U35324 (N_35324,N_28932,N_29725);
xnor U35325 (N_35325,N_27008,N_22897);
or U35326 (N_35326,N_22686,N_27544);
xnor U35327 (N_35327,N_26886,N_23681);
nand U35328 (N_35328,N_21187,N_24312);
nand U35329 (N_35329,N_29699,N_27292);
xor U35330 (N_35330,N_28654,N_21071);
nand U35331 (N_35331,N_24935,N_28066);
xor U35332 (N_35332,N_25721,N_25270);
xnor U35333 (N_35333,N_23803,N_28809);
and U35334 (N_35334,N_29001,N_23296);
nor U35335 (N_35335,N_26293,N_23411);
nand U35336 (N_35336,N_28548,N_23972);
or U35337 (N_35337,N_23528,N_21255);
nor U35338 (N_35338,N_23791,N_29932);
xor U35339 (N_35339,N_21471,N_27266);
and U35340 (N_35340,N_27066,N_23534);
and U35341 (N_35341,N_25540,N_21717);
xnor U35342 (N_35342,N_28925,N_25697);
nand U35343 (N_35343,N_22208,N_22382);
nand U35344 (N_35344,N_21823,N_22283);
xnor U35345 (N_35345,N_28365,N_25256);
xnor U35346 (N_35346,N_25563,N_27590);
nand U35347 (N_35347,N_25301,N_29850);
nor U35348 (N_35348,N_28888,N_24901);
nor U35349 (N_35349,N_25353,N_27984);
nor U35350 (N_35350,N_24514,N_20325);
and U35351 (N_35351,N_20770,N_25057);
nand U35352 (N_35352,N_23815,N_20348);
xor U35353 (N_35353,N_20429,N_26528);
nand U35354 (N_35354,N_25739,N_26692);
xnor U35355 (N_35355,N_20103,N_23522);
nor U35356 (N_35356,N_28438,N_27213);
nor U35357 (N_35357,N_29679,N_28897);
or U35358 (N_35358,N_28357,N_28438);
xor U35359 (N_35359,N_20007,N_23345);
nor U35360 (N_35360,N_25029,N_20411);
nand U35361 (N_35361,N_27963,N_25029);
xor U35362 (N_35362,N_27730,N_22438);
and U35363 (N_35363,N_23747,N_21001);
xnor U35364 (N_35364,N_26247,N_22136);
and U35365 (N_35365,N_20696,N_22071);
nor U35366 (N_35366,N_22887,N_20953);
xor U35367 (N_35367,N_22204,N_22185);
xor U35368 (N_35368,N_27399,N_22910);
xnor U35369 (N_35369,N_28472,N_25311);
or U35370 (N_35370,N_20381,N_27185);
or U35371 (N_35371,N_21224,N_24092);
or U35372 (N_35372,N_26228,N_27361);
or U35373 (N_35373,N_20011,N_20044);
nor U35374 (N_35374,N_28629,N_25053);
and U35375 (N_35375,N_26673,N_21397);
nor U35376 (N_35376,N_28214,N_22849);
nand U35377 (N_35377,N_23416,N_25004);
and U35378 (N_35378,N_26682,N_26024);
or U35379 (N_35379,N_26293,N_20433);
nand U35380 (N_35380,N_22253,N_29210);
and U35381 (N_35381,N_29235,N_29699);
xor U35382 (N_35382,N_24138,N_23251);
and U35383 (N_35383,N_20848,N_20010);
or U35384 (N_35384,N_21032,N_29528);
or U35385 (N_35385,N_25489,N_23322);
or U35386 (N_35386,N_21862,N_22725);
or U35387 (N_35387,N_22925,N_24566);
nand U35388 (N_35388,N_21218,N_23723);
or U35389 (N_35389,N_26416,N_23394);
nand U35390 (N_35390,N_24820,N_23035);
or U35391 (N_35391,N_25860,N_23976);
and U35392 (N_35392,N_20236,N_21481);
nand U35393 (N_35393,N_20283,N_29275);
and U35394 (N_35394,N_26031,N_25717);
nand U35395 (N_35395,N_21560,N_20553);
xor U35396 (N_35396,N_20394,N_27784);
and U35397 (N_35397,N_25371,N_22774);
xor U35398 (N_35398,N_24326,N_29910);
and U35399 (N_35399,N_26675,N_27910);
or U35400 (N_35400,N_24831,N_25786);
and U35401 (N_35401,N_23131,N_23378);
nor U35402 (N_35402,N_28796,N_26805);
xnor U35403 (N_35403,N_23190,N_22485);
nor U35404 (N_35404,N_28450,N_20517);
nand U35405 (N_35405,N_26636,N_22680);
nor U35406 (N_35406,N_23019,N_23346);
or U35407 (N_35407,N_27631,N_25322);
nor U35408 (N_35408,N_21746,N_27793);
xor U35409 (N_35409,N_23279,N_28179);
nor U35410 (N_35410,N_20348,N_22419);
nor U35411 (N_35411,N_25083,N_27376);
xnor U35412 (N_35412,N_23092,N_21582);
and U35413 (N_35413,N_27882,N_22883);
xnor U35414 (N_35414,N_20831,N_22570);
and U35415 (N_35415,N_26009,N_26034);
xor U35416 (N_35416,N_22791,N_27031);
nand U35417 (N_35417,N_26156,N_28277);
nand U35418 (N_35418,N_20762,N_20967);
or U35419 (N_35419,N_24025,N_24079);
and U35420 (N_35420,N_25692,N_23677);
nand U35421 (N_35421,N_24254,N_28631);
and U35422 (N_35422,N_25286,N_24248);
nand U35423 (N_35423,N_23740,N_23977);
or U35424 (N_35424,N_21090,N_29232);
or U35425 (N_35425,N_26256,N_29994);
xor U35426 (N_35426,N_24539,N_24002);
nand U35427 (N_35427,N_22491,N_23685);
nand U35428 (N_35428,N_26821,N_28816);
or U35429 (N_35429,N_28241,N_25285);
xor U35430 (N_35430,N_26908,N_23396);
or U35431 (N_35431,N_25935,N_26218);
and U35432 (N_35432,N_27611,N_27193);
or U35433 (N_35433,N_25687,N_21581);
and U35434 (N_35434,N_29459,N_20461);
or U35435 (N_35435,N_26503,N_24720);
nand U35436 (N_35436,N_26744,N_26159);
xor U35437 (N_35437,N_28001,N_22322);
nand U35438 (N_35438,N_24913,N_26628);
xnor U35439 (N_35439,N_28759,N_26201);
and U35440 (N_35440,N_27189,N_29590);
nor U35441 (N_35441,N_20479,N_29058);
nor U35442 (N_35442,N_28130,N_20093);
xor U35443 (N_35443,N_21156,N_21080);
nand U35444 (N_35444,N_21176,N_27040);
or U35445 (N_35445,N_27414,N_25813);
and U35446 (N_35446,N_23174,N_27636);
nor U35447 (N_35447,N_24923,N_24559);
and U35448 (N_35448,N_25757,N_26384);
nand U35449 (N_35449,N_20001,N_24720);
nand U35450 (N_35450,N_20335,N_20825);
or U35451 (N_35451,N_24566,N_29009);
xnor U35452 (N_35452,N_20375,N_20754);
nand U35453 (N_35453,N_29376,N_22379);
nor U35454 (N_35454,N_22140,N_24686);
or U35455 (N_35455,N_22160,N_28736);
or U35456 (N_35456,N_24076,N_26643);
and U35457 (N_35457,N_27493,N_29901);
or U35458 (N_35458,N_21624,N_23871);
xor U35459 (N_35459,N_24338,N_22995);
and U35460 (N_35460,N_23471,N_27955);
or U35461 (N_35461,N_21096,N_22662);
and U35462 (N_35462,N_26770,N_23838);
nand U35463 (N_35463,N_29936,N_22360);
and U35464 (N_35464,N_28463,N_22087);
nor U35465 (N_35465,N_25464,N_26603);
and U35466 (N_35466,N_25615,N_21048);
nor U35467 (N_35467,N_21972,N_29156);
nor U35468 (N_35468,N_27466,N_27477);
or U35469 (N_35469,N_22346,N_27692);
xnor U35470 (N_35470,N_26634,N_22574);
nand U35471 (N_35471,N_28763,N_22140);
xor U35472 (N_35472,N_20936,N_27973);
nor U35473 (N_35473,N_27842,N_28710);
xnor U35474 (N_35474,N_21857,N_20426);
xnor U35475 (N_35475,N_20743,N_22796);
and U35476 (N_35476,N_20138,N_26012);
and U35477 (N_35477,N_29285,N_22376);
xnor U35478 (N_35478,N_26400,N_27765);
or U35479 (N_35479,N_26481,N_25629);
xnor U35480 (N_35480,N_29371,N_28795);
nand U35481 (N_35481,N_23683,N_29989);
and U35482 (N_35482,N_21339,N_28744);
or U35483 (N_35483,N_21729,N_20287);
xnor U35484 (N_35484,N_23719,N_23314);
and U35485 (N_35485,N_21887,N_26488);
or U35486 (N_35486,N_29139,N_25342);
xnor U35487 (N_35487,N_29819,N_27973);
nand U35488 (N_35488,N_24244,N_24864);
nor U35489 (N_35489,N_28384,N_29186);
nand U35490 (N_35490,N_24339,N_20824);
xnor U35491 (N_35491,N_25383,N_21240);
nor U35492 (N_35492,N_22067,N_27746);
nor U35493 (N_35493,N_20361,N_28755);
or U35494 (N_35494,N_24086,N_26169);
and U35495 (N_35495,N_22160,N_23192);
xnor U35496 (N_35496,N_26062,N_22578);
or U35497 (N_35497,N_22736,N_27417);
and U35498 (N_35498,N_25045,N_23805);
and U35499 (N_35499,N_22619,N_24909);
nand U35500 (N_35500,N_21652,N_27609);
or U35501 (N_35501,N_23944,N_29879);
or U35502 (N_35502,N_21659,N_24045);
xnor U35503 (N_35503,N_28321,N_20424);
nand U35504 (N_35504,N_22687,N_21615);
xor U35505 (N_35505,N_21231,N_28870);
nor U35506 (N_35506,N_29712,N_28795);
xor U35507 (N_35507,N_23671,N_24395);
nand U35508 (N_35508,N_21794,N_20838);
nor U35509 (N_35509,N_21891,N_22514);
nand U35510 (N_35510,N_22886,N_26919);
or U35511 (N_35511,N_24118,N_24174);
and U35512 (N_35512,N_27830,N_26454);
nand U35513 (N_35513,N_23905,N_28255);
or U35514 (N_35514,N_25695,N_21757);
or U35515 (N_35515,N_20417,N_28922);
nor U35516 (N_35516,N_28441,N_29916);
xor U35517 (N_35517,N_21840,N_22346);
or U35518 (N_35518,N_28452,N_26091);
and U35519 (N_35519,N_24861,N_27603);
xnor U35520 (N_35520,N_26013,N_29987);
nand U35521 (N_35521,N_24630,N_28345);
nand U35522 (N_35522,N_22880,N_24704);
or U35523 (N_35523,N_25558,N_22065);
xor U35524 (N_35524,N_24838,N_28402);
and U35525 (N_35525,N_28576,N_23835);
or U35526 (N_35526,N_23435,N_24740);
or U35527 (N_35527,N_26815,N_27695);
and U35528 (N_35528,N_27632,N_23609);
or U35529 (N_35529,N_23254,N_21053);
or U35530 (N_35530,N_27984,N_29149);
or U35531 (N_35531,N_21707,N_23690);
and U35532 (N_35532,N_22335,N_22169);
and U35533 (N_35533,N_29976,N_27657);
or U35534 (N_35534,N_22162,N_23090);
nand U35535 (N_35535,N_26825,N_21919);
xor U35536 (N_35536,N_21043,N_29144);
or U35537 (N_35537,N_29206,N_21217);
nor U35538 (N_35538,N_21635,N_20410);
or U35539 (N_35539,N_29007,N_28024);
xnor U35540 (N_35540,N_23098,N_23107);
nor U35541 (N_35541,N_21361,N_24206);
nand U35542 (N_35542,N_28957,N_27598);
or U35543 (N_35543,N_22010,N_26564);
nor U35544 (N_35544,N_27836,N_20887);
or U35545 (N_35545,N_25284,N_21518);
and U35546 (N_35546,N_28294,N_26011);
and U35547 (N_35547,N_27189,N_25733);
and U35548 (N_35548,N_23140,N_25746);
and U35549 (N_35549,N_22241,N_23378);
nand U35550 (N_35550,N_25931,N_21357);
nor U35551 (N_35551,N_23281,N_23396);
xnor U35552 (N_35552,N_25441,N_28489);
xor U35553 (N_35553,N_22077,N_22610);
nand U35554 (N_35554,N_24119,N_20048);
nor U35555 (N_35555,N_26198,N_23869);
nor U35556 (N_35556,N_26089,N_24163);
nand U35557 (N_35557,N_22888,N_29505);
or U35558 (N_35558,N_24003,N_25495);
or U35559 (N_35559,N_21861,N_27505);
and U35560 (N_35560,N_25451,N_26924);
nand U35561 (N_35561,N_21711,N_24215);
xnor U35562 (N_35562,N_24661,N_21989);
or U35563 (N_35563,N_22080,N_20434);
and U35564 (N_35564,N_25627,N_21933);
xnor U35565 (N_35565,N_26003,N_27592);
nand U35566 (N_35566,N_22443,N_28730);
nor U35567 (N_35567,N_24041,N_27566);
or U35568 (N_35568,N_20723,N_29000);
or U35569 (N_35569,N_24973,N_23093);
xor U35570 (N_35570,N_22921,N_23223);
nor U35571 (N_35571,N_28538,N_26317);
or U35572 (N_35572,N_28929,N_29510);
or U35573 (N_35573,N_22544,N_21192);
and U35574 (N_35574,N_22412,N_29577);
and U35575 (N_35575,N_22110,N_22045);
or U35576 (N_35576,N_21615,N_28861);
or U35577 (N_35577,N_21865,N_24782);
or U35578 (N_35578,N_20053,N_20069);
nor U35579 (N_35579,N_28554,N_20673);
or U35580 (N_35580,N_20081,N_26275);
or U35581 (N_35581,N_29154,N_21422);
nor U35582 (N_35582,N_21645,N_24184);
and U35583 (N_35583,N_21733,N_26025);
and U35584 (N_35584,N_21981,N_23164);
xor U35585 (N_35585,N_20819,N_20481);
or U35586 (N_35586,N_25321,N_27067);
or U35587 (N_35587,N_21750,N_21017);
and U35588 (N_35588,N_23266,N_29396);
or U35589 (N_35589,N_21591,N_27882);
or U35590 (N_35590,N_26191,N_23446);
nor U35591 (N_35591,N_22595,N_25468);
nand U35592 (N_35592,N_24721,N_28344);
nor U35593 (N_35593,N_28781,N_22404);
nand U35594 (N_35594,N_29238,N_25411);
nand U35595 (N_35595,N_22249,N_28720);
and U35596 (N_35596,N_29624,N_29936);
nor U35597 (N_35597,N_26185,N_29724);
and U35598 (N_35598,N_24351,N_25982);
nor U35599 (N_35599,N_25594,N_24327);
nand U35600 (N_35600,N_25769,N_23475);
xnor U35601 (N_35601,N_25627,N_28127);
xnor U35602 (N_35602,N_25105,N_27810);
or U35603 (N_35603,N_29383,N_23555);
nor U35604 (N_35604,N_29052,N_27971);
xor U35605 (N_35605,N_24101,N_27183);
and U35606 (N_35606,N_22165,N_27226);
or U35607 (N_35607,N_28703,N_20846);
nor U35608 (N_35608,N_24530,N_28137);
nor U35609 (N_35609,N_27356,N_28210);
and U35610 (N_35610,N_22228,N_27959);
and U35611 (N_35611,N_20851,N_25128);
or U35612 (N_35612,N_22971,N_27634);
xnor U35613 (N_35613,N_26722,N_23489);
nor U35614 (N_35614,N_28061,N_22910);
and U35615 (N_35615,N_20778,N_22427);
nor U35616 (N_35616,N_28726,N_22841);
nor U35617 (N_35617,N_26152,N_22974);
nor U35618 (N_35618,N_20528,N_25135);
nand U35619 (N_35619,N_22783,N_23981);
nand U35620 (N_35620,N_29574,N_27538);
nand U35621 (N_35621,N_21970,N_22526);
nor U35622 (N_35622,N_22415,N_28700);
nor U35623 (N_35623,N_29630,N_23865);
nand U35624 (N_35624,N_23920,N_28812);
xnor U35625 (N_35625,N_22253,N_26817);
xor U35626 (N_35626,N_27110,N_24618);
nor U35627 (N_35627,N_25179,N_25584);
xnor U35628 (N_35628,N_26397,N_25623);
or U35629 (N_35629,N_22724,N_26329);
xor U35630 (N_35630,N_26001,N_23427);
nor U35631 (N_35631,N_26235,N_23754);
xor U35632 (N_35632,N_22677,N_26711);
nor U35633 (N_35633,N_22289,N_28676);
nor U35634 (N_35634,N_24811,N_21403);
nor U35635 (N_35635,N_28467,N_27645);
or U35636 (N_35636,N_29735,N_22600);
or U35637 (N_35637,N_24322,N_20200);
xor U35638 (N_35638,N_20912,N_24727);
xnor U35639 (N_35639,N_27396,N_26282);
and U35640 (N_35640,N_26429,N_24626);
nor U35641 (N_35641,N_21002,N_21624);
or U35642 (N_35642,N_28914,N_26304);
xnor U35643 (N_35643,N_22210,N_23959);
and U35644 (N_35644,N_25113,N_27433);
nor U35645 (N_35645,N_20478,N_27614);
and U35646 (N_35646,N_26186,N_27652);
xor U35647 (N_35647,N_29473,N_20912);
nor U35648 (N_35648,N_29092,N_23921);
nor U35649 (N_35649,N_25833,N_21907);
xor U35650 (N_35650,N_23924,N_20068);
nand U35651 (N_35651,N_26586,N_20276);
or U35652 (N_35652,N_22407,N_27915);
nand U35653 (N_35653,N_24460,N_27812);
nand U35654 (N_35654,N_27321,N_22401);
nor U35655 (N_35655,N_21821,N_29918);
xor U35656 (N_35656,N_28717,N_24440);
and U35657 (N_35657,N_26094,N_23119);
nand U35658 (N_35658,N_26677,N_27211);
nor U35659 (N_35659,N_29302,N_26906);
and U35660 (N_35660,N_23483,N_25353);
nand U35661 (N_35661,N_25437,N_27576);
nand U35662 (N_35662,N_21332,N_29736);
xor U35663 (N_35663,N_24326,N_28378);
nand U35664 (N_35664,N_24315,N_24491);
and U35665 (N_35665,N_23210,N_20698);
xnor U35666 (N_35666,N_23741,N_28955);
xor U35667 (N_35667,N_21103,N_26874);
nand U35668 (N_35668,N_28366,N_23750);
nor U35669 (N_35669,N_25406,N_26159);
xnor U35670 (N_35670,N_21501,N_28300);
nand U35671 (N_35671,N_21045,N_25711);
nor U35672 (N_35672,N_21111,N_27748);
xor U35673 (N_35673,N_23090,N_22636);
or U35674 (N_35674,N_22093,N_25494);
or U35675 (N_35675,N_28876,N_24352);
xnor U35676 (N_35676,N_21764,N_26348);
or U35677 (N_35677,N_20789,N_25023);
and U35678 (N_35678,N_22992,N_25156);
nor U35679 (N_35679,N_21855,N_24300);
and U35680 (N_35680,N_29345,N_22025);
xnor U35681 (N_35681,N_27157,N_24706);
xor U35682 (N_35682,N_27272,N_22925);
and U35683 (N_35683,N_26716,N_29245);
nand U35684 (N_35684,N_28044,N_27075);
nand U35685 (N_35685,N_26322,N_20576);
and U35686 (N_35686,N_23914,N_23575);
and U35687 (N_35687,N_29232,N_24370);
xor U35688 (N_35688,N_29946,N_26262);
or U35689 (N_35689,N_26148,N_29263);
or U35690 (N_35690,N_27645,N_27706);
nor U35691 (N_35691,N_25959,N_25929);
or U35692 (N_35692,N_22955,N_21011);
or U35693 (N_35693,N_20976,N_23931);
or U35694 (N_35694,N_20250,N_21103);
xnor U35695 (N_35695,N_27515,N_22201);
nand U35696 (N_35696,N_20313,N_22562);
xnor U35697 (N_35697,N_24874,N_24760);
nand U35698 (N_35698,N_23744,N_25611);
nor U35699 (N_35699,N_28511,N_22053);
nand U35700 (N_35700,N_20265,N_22274);
xnor U35701 (N_35701,N_23191,N_22528);
nor U35702 (N_35702,N_26027,N_22005);
nand U35703 (N_35703,N_26047,N_27262);
and U35704 (N_35704,N_20203,N_24636);
nor U35705 (N_35705,N_24427,N_20463);
xnor U35706 (N_35706,N_28669,N_23470);
nor U35707 (N_35707,N_21652,N_29378);
nand U35708 (N_35708,N_24584,N_28800);
nor U35709 (N_35709,N_21560,N_27262);
nor U35710 (N_35710,N_20305,N_25882);
nand U35711 (N_35711,N_27308,N_27469);
or U35712 (N_35712,N_26346,N_28649);
xnor U35713 (N_35713,N_26464,N_27967);
nor U35714 (N_35714,N_23678,N_21017);
nand U35715 (N_35715,N_29875,N_24942);
nand U35716 (N_35716,N_24298,N_24250);
nor U35717 (N_35717,N_25013,N_25549);
or U35718 (N_35718,N_21682,N_26033);
nand U35719 (N_35719,N_20626,N_25519);
xor U35720 (N_35720,N_27763,N_21116);
or U35721 (N_35721,N_29406,N_20328);
and U35722 (N_35722,N_29551,N_22014);
nor U35723 (N_35723,N_23476,N_27891);
xor U35724 (N_35724,N_23795,N_29255);
xor U35725 (N_35725,N_25351,N_27401);
xor U35726 (N_35726,N_28176,N_21142);
nor U35727 (N_35727,N_29276,N_23591);
nand U35728 (N_35728,N_23394,N_24048);
nand U35729 (N_35729,N_23745,N_29333);
nand U35730 (N_35730,N_26964,N_24309);
nor U35731 (N_35731,N_27160,N_29302);
or U35732 (N_35732,N_24495,N_22345);
nand U35733 (N_35733,N_27492,N_21448);
xnor U35734 (N_35734,N_26462,N_23915);
nor U35735 (N_35735,N_21675,N_27216);
and U35736 (N_35736,N_26946,N_21168);
and U35737 (N_35737,N_21590,N_29778);
xor U35738 (N_35738,N_25453,N_23894);
or U35739 (N_35739,N_28260,N_22079);
xnor U35740 (N_35740,N_21925,N_21414);
nor U35741 (N_35741,N_24580,N_28454);
nor U35742 (N_35742,N_23174,N_22435);
nor U35743 (N_35743,N_22963,N_26167);
nor U35744 (N_35744,N_28479,N_21815);
or U35745 (N_35745,N_23268,N_29687);
xnor U35746 (N_35746,N_21796,N_22005);
and U35747 (N_35747,N_25514,N_29419);
or U35748 (N_35748,N_27578,N_26567);
nand U35749 (N_35749,N_21737,N_27193);
nand U35750 (N_35750,N_29731,N_26944);
nand U35751 (N_35751,N_28332,N_22043);
xnor U35752 (N_35752,N_25235,N_29851);
and U35753 (N_35753,N_23059,N_27379);
xnor U35754 (N_35754,N_25480,N_29107);
xor U35755 (N_35755,N_21422,N_27384);
nor U35756 (N_35756,N_28521,N_25028);
or U35757 (N_35757,N_22448,N_20915);
xor U35758 (N_35758,N_22463,N_26649);
nor U35759 (N_35759,N_24249,N_24129);
or U35760 (N_35760,N_23032,N_20285);
or U35761 (N_35761,N_27052,N_23901);
or U35762 (N_35762,N_20080,N_25471);
xor U35763 (N_35763,N_26141,N_22457);
xor U35764 (N_35764,N_27680,N_20023);
and U35765 (N_35765,N_27052,N_23475);
and U35766 (N_35766,N_29822,N_26574);
nand U35767 (N_35767,N_29801,N_25887);
and U35768 (N_35768,N_25988,N_20011);
xor U35769 (N_35769,N_21054,N_25777);
nand U35770 (N_35770,N_23999,N_29615);
or U35771 (N_35771,N_26505,N_22228);
xnor U35772 (N_35772,N_29720,N_20701);
xor U35773 (N_35773,N_28243,N_22640);
nand U35774 (N_35774,N_28209,N_26196);
nand U35775 (N_35775,N_27095,N_25686);
or U35776 (N_35776,N_28534,N_20468);
or U35777 (N_35777,N_22428,N_20550);
nand U35778 (N_35778,N_20800,N_26753);
xnor U35779 (N_35779,N_23410,N_27459);
nand U35780 (N_35780,N_26468,N_21004);
xnor U35781 (N_35781,N_26320,N_21399);
nor U35782 (N_35782,N_27353,N_25356);
and U35783 (N_35783,N_21009,N_27017);
nand U35784 (N_35784,N_27503,N_25232);
and U35785 (N_35785,N_28442,N_20577);
xor U35786 (N_35786,N_28444,N_21925);
nor U35787 (N_35787,N_27432,N_23595);
nand U35788 (N_35788,N_21312,N_25929);
or U35789 (N_35789,N_20331,N_25822);
xor U35790 (N_35790,N_24373,N_24862);
xnor U35791 (N_35791,N_21908,N_23964);
and U35792 (N_35792,N_27304,N_24231);
or U35793 (N_35793,N_25633,N_27161);
and U35794 (N_35794,N_26532,N_22604);
nand U35795 (N_35795,N_28316,N_22423);
or U35796 (N_35796,N_21642,N_24541);
or U35797 (N_35797,N_23064,N_26728);
xor U35798 (N_35798,N_24682,N_20178);
or U35799 (N_35799,N_23663,N_27938);
or U35800 (N_35800,N_24788,N_24444);
or U35801 (N_35801,N_29400,N_22168);
or U35802 (N_35802,N_20215,N_24656);
xor U35803 (N_35803,N_20334,N_25127);
nor U35804 (N_35804,N_27066,N_20016);
nor U35805 (N_35805,N_25784,N_23281);
and U35806 (N_35806,N_25528,N_27282);
and U35807 (N_35807,N_27875,N_29643);
or U35808 (N_35808,N_28774,N_23085);
or U35809 (N_35809,N_28354,N_27995);
nor U35810 (N_35810,N_28360,N_21282);
or U35811 (N_35811,N_26744,N_21923);
xnor U35812 (N_35812,N_21336,N_20874);
or U35813 (N_35813,N_22257,N_20033);
and U35814 (N_35814,N_20076,N_21734);
or U35815 (N_35815,N_23983,N_22553);
xnor U35816 (N_35816,N_29697,N_25143);
nand U35817 (N_35817,N_27706,N_22506);
and U35818 (N_35818,N_23272,N_25519);
or U35819 (N_35819,N_25067,N_25179);
and U35820 (N_35820,N_22469,N_24130);
nor U35821 (N_35821,N_29689,N_26133);
xnor U35822 (N_35822,N_23964,N_23249);
nand U35823 (N_35823,N_26544,N_27063);
nand U35824 (N_35824,N_25623,N_28318);
xnor U35825 (N_35825,N_29231,N_23249);
and U35826 (N_35826,N_26569,N_24264);
xor U35827 (N_35827,N_23899,N_26307);
or U35828 (N_35828,N_24814,N_24758);
and U35829 (N_35829,N_29380,N_26837);
xor U35830 (N_35830,N_20825,N_21814);
nor U35831 (N_35831,N_25359,N_21130);
nand U35832 (N_35832,N_23337,N_27277);
nor U35833 (N_35833,N_29107,N_22592);
nand U35834 (N_35834,N_25556,N_23631);
or U35835 (N_35835,N_22169,N_26626);
nor U35836 (N_35836,N_25260,N_29815);
nor U35837 (N_35837,N_25448,N_28361);
or U35838 (N_35838,N_28308,N_21168);
nand U35839 (N_35839,N_21367,N_20420);
and U35840 (N_35840,N_22236,N_29576);
or U35841 (N_35841,N_26961,N_24425);
nand U35842 (N_35842,N_21070,N_22134);
nand U35843 (N_35843,N_25017,N_22674);
nor U35844 (N_35844,N_29708,N_24802);
nor U35845 (N_35845,N_29491,N_20217);
nand U35846 (N_35846,N_24467,N_23481);
xor U35847 (N_35847,N_28247,N_28748);
nor U35848 (N_35848,N_26201,N_23064);
nand U35849 (N_35849,N_22721,N_23505);
nor U35850 (N_35850,N_28925,N_26645);
and U35851 (N_35851,N_24339,N_22086);
nor U35852 (N_35852,N_24549,N_29941);
nand U35853 (N_35853,N_22524,N_22610);
xor U35854 (N_35854,N_29737,N_25958);
nor U35855 (N_35855,N_26538,N_22997);
nand U35856 (N_35856,N_24581,N_21824);
nor U35857 (N_35857,N_27431,N_29295);
xor U35858 (N_35858,N_24921,N_25499);
nand U35859 (N_35859,N_28668,N_25742);
and U35860 (N_35860,N_22306,N_29443);
and U35861 (N_35861,N_25432,N_27844);
nand U35862 (N_35862,N_21155,N_28108);
xnor U35863 (N_35863,N_26413,N_26100);
nand U35864 (N_35864,N_28208,N_26374);
nand U35865 (N_35865,N_20432,N_21478);
and U35866 (N_35866,N_23000,N_29172);
xor U35867 (N_35867,N_28770,N_26608);
or U35868 (N_35868,N_24939,N_22435);
nand U35869 (N_35869,N_25321,N_28374);
and U35870 (N_35870,N_24742,N_24871);
and U35871 (N_35871,N_27341,N_29353);
nor U35872 (N_35872,N_29312,N_23135);
nand U35873 (N_35873,N_21560,N_22613);
and U35874 (N_35874,N_25745,N_22575);
xnor U35875 (N_35875,N_25786,N_23719);
or U35876 (N_35876,N_26492,N_27420);
xnor U35877 (N_35877,N_29407,N_27132);
nor U35878 (N_35878,N_28132,N_26403);
nor U35879 (N_35879,N_23441,N_27869);
nand U35880 (N_35880,N_22894,N_25331);
nand U35881 (N_35881,N_25263,N_29937);
or U35882 (N_35882,N_23921,N_26137);
and U35883 (N_35883,N_24982,N_22053);
xor U35884 (N_35884,N_21327,N_24852);
xnor U35885 (N_35885,N_24451,N_28855);
xor U35886 (N_35886,N_20220,N_22010);
nor U35887 (N_35887,N_22942,N_21206);
nand U35888 (N_35888,N_25975,N_23406);
nand U35889 (N_35889,N_26053,N_26712);
and U35890 (N_35890,N_29686,N_27566);
nor U35891 (N_35891,N_29611,N_22364);
nor U35892 (N_35892,N_26780,N_27551);
or U35893 (N_35893,N_21507,N_26097);
xnor U35894 (N_35894,N_25328,N_26045);
and U35895 (N_35895,N_26262,N_26872);
nor U35896 (N_35896,N_29959,N_24729);
and U35897 (N_35897,N_28751,N_20217);
xnor U35898 (N_35898,N_28815,N_28150);
nand U35899 (N_35899,N_28472,N_24260);
nor U35900 (N_35900,N_22563,N_27445);
and U35901 (N_35901,N_27291,N_27713);
and U35902 (N_35902,N_20359,N_25865);
and U35903 (N_35903,N_23586,N_24326);
and U35904 (N_35904,N_24925,N_26142);
and U35905 (N_35905,N_27129,N_29041);
or U35906 (N_35906,N_22052,N_20610);
xnor U35907 (N_35907,N_25051,N_28999);
nor U35908 (N_35908,N_25314,N_29630);
or U35909 (N_35909,N_20923,N_21205);
nand U35910 (N_35910,N_21210,N_25870);
or U35911 (N_35911,N_25842,N_29983);
xnor U35912 (N_35912,N_27190,N_23652);
and U35913 (N_35913,N_23671,N_23219);
xor U35914 (N_35914,N_29784,N_26237);
or U35915 (N_35915,N_22149,N_26690);
or U35916 (N_35916,N_26105,N_28775);
nand U35917 (N_35917,N_22251,N_29708);
nand U35918 (N_35918,N_20023,N_28620);
nand U35919 (N_35919,N_26795,N_28828);
or U35920 (N_35920,N_29195,N_20312);
and U35921 (N_35921,N_23839,N_24781);
nand U35922 (N_35922,N_25216,N_28663);
nor U35923 (N_35923,N_27811,N_21853);
or U35924 (N_35924,N_21704,N_22474);
xor U35925 (N_35925,N_26273,N_23063);
xor U35926 (N_35926,N_23930,N_26415);
xor U35927 (N_35927,N_26116,N_21613);
nor U35928 (N_35928,N_26907,N_21091);
and U35929 (N_35929,N_24621,N_27628);
or U35930 (N_35930,N_20846,N_29246);
xor U35931 (N_35931,N_23334,N_26206);
nor U35932 (N_35932,N_25809,N_20561);
nand U35933 (N_35933,N_24245,N_22248);
xnor U35934 (N_35934,N_27531,N_28020);
nor U35935 (N_35935,N_20656,N_23089);
xor U35936 (N_35936,N_28681,N_28560);
nand U35937 (N_35937,N_21963,N_29602);
and U35938 (N_35938,N_27051,N_29280);
and U35939 (N_35939,N_28871,N_28852);
nor U35940 (N_35940,N_26546,N_26371);
nor U35941 (N_35941,N_28123,N_25458);
nand U35942 (N_35942,N_27559,N_26644);
and U35943 (N_35943,N_22322,N_22116);
and U35944 (N_35944,N_28978,N_23373);
or U35945 (N_35945,N_28747,N_25516);
or U35946 (N_35946,N_23591,N_23343);
or U35947 (N_35947,N_24167,N_22473);
or U35948 (N_35948,N_21215,N_23086);
and U35949 (N_35949,N_25814,N_26319);
and U35950 (N_35950,N_28480,N_22795);
xnor U35951 (N_35951,N_27237,N_27553);
or U35952 (N_35952,N_28169,N_23017);
xnor U35953 (N_35953,N_28130,N_28541);
nor U35954 (N_35954,N_29990,N_20309);
nand U35955 (N_35955,N_26994,N_26714);
and U35956 (N_35956,N_20532,N_25348);
nand U35957 (N_35957,N_26193,N_20392);
xor U35958 (N_35958,N_28497,N_28996);
nand U35959 (N_35959,N_21081,N_23011);
nand U35960 (N_35960,N_20155,N_29086);
nand U35961 (N_35961,N_27021,N_23472);
and U35962 (N_35962,N_22346,N_28142);
or U35963 (N_35963,N_26987,N_29270);
and U35964 (N_35964,N_21015,N_24161);
and U35965 (N_35965,N_29969,N_22784);
nand U35966 (N_35966,N_23406,N_25558);
or U35967 (N_35967,N_27977,N_26675);
xor U35968 (N_35968,N_29389,N_22874);
and U35969 (N_35969,N_20336,N_21434);
xnor U35970 (N_35970,N_24991,N_25557);
or U35971 (N_35971,N_22704,N_20079);
nand U35972 (N_35972,N_22180,N_21956);
nor U35973 (N_35973,N_21624,N_22494);
nor U35974 (N_35974,N_24480,N_24870);
nand U35975 (N_35975,N_25012,N_27734);
nor U35976 (N_35976,N_21826,N_29918);
nor U35977 (N_35977,N_22189,N_27110);
xnor U35978 (N_35978,N_24999,N_21761);
or U35979 (N_35979,N_20321,N_29846);
and U35980 (N_35980,N_25877,N_28703);
and U35981 (N_35981,N_28241,N_21316);
nand U35982 (N_35982,N_29129,N_28760);
xor U35983 (N_35983,N_21111,N_26828);
and U35984 (N_35984,N_25817,N_26901);
and U35985 (N_35985,N_21577,N_21038);
xnor U35986 (N_35986,N_21629,N_20254);
and U35987 (N_35987,N_21532,N_21572);
or U35988 (N_35988,N_23853,N_24343);
or U35989 (N_35989,N_28505,N_21015);
and U35990 (N_35990,N_26848,N_28485);
xor U35991 (N_35991,N_27270,N_29590);
and U35992 (N_35992,N_21401,N_24383);
nand U35993 (N_35993,N_23091,N_21562);
or U35994 (N_35994,N_24739,N_26403);
and U35995 (N_35995,N_20379,N_22449);
nor U35996 (N_35996,N_28068,N_22129);
nor U35997 (N_35997,N_23963,N_26155);
and U35998 (N_35998,N_29213,N_26565);
or U35999 (N_35999,N_27715,N_21789);
and U36000 (N_36000,N_20685,N_28179);
xnor U36001 (N_36001,N_28484,N_22356);
xnor U36002 (N_36002,N_22766,N_20335);
or U36003 (N_36003,N_20109,N_28595);
nand U36004 (N_36004,N_29312,N_20506);
or U36005 (N_36005,N_29788,N_20836);
nor U36006 (N_36006,N_27738,N_23206);
or U36007 (N_36007,N_27132,N_21912);
and U36008 (N_36008,N_29112,N_22445);
and U36009 (N_36009,N_25583,N_28809);
nand U36010 (N_36010,N_23764,N_20796);
or U36011 (N_36011,N_26610,N_22362);
nand U36012 (N_36012,N_22271,N_21207);
or U36013 (N_36013,N_25687,N_24253);
nand U36014 (N_36014,N_20063,N_28285);
nor U36015 (N_36015,N_22368,N_25429);
and U36016 (N_36016,N_28237,N_20959);
nor U36017 (N_36017,N_27994,N_29953);
nor U36018 (N_36018,N_29129,N_26681);
nand U36019 (N_36019,N_27077,N_22920);
nand U36020 (N_36020,N_26813,N_20782);
nand U36021 (N_36021,N_20126,N_28376);
or U36022 (N_36022,N_20964,N_24511);
or U36023 (N_36023,N_20101,N_20385);
nand U36024 (N_36024,N_29547,N_26082);
or U36025 (N_36025,N_25005,N_20579);
xnor U36026 (N_36026,N_21878,N_27227);
xnor U36027 (N_36027,N_26899,N_28152);
or U36028 (N_36028,N_29837,N_20300);
nor U36029 (N_36029,N_23536,N_25566);
or U36030 (N_36030,N_25898,N_22065);
nor U36031 (N_36031,N_20750,N_28686);
or U36032 (N_36032,N_28614,N_25203);
and U36033 (N_36033,N_29154,N_27685);
and U36034 (N_36034,N_20240,N_28573);
or U36035 (N_36035,N_28855,N_20973);
and U36036 (N_36036,N_23780,N_25183);
xnor U36037 (N_36037,N_20935,N_28167);
and U36038 (N_36038,N_27326,N_20645);
nor U36039 (N_36039,N_25760,N_20909);
and U36040 (N_36040,N_22899,N_27928);
nand U36041 (N_36041,N_24255,N_25380);
or U36042 (N_36042,N_23490,N_20692);
nor U36043 (N_36043,N_22866,N_23796);
nor U36044 (N_36044,N_26882,N_21038);
xor U36045 (N_36045,N_26867,N_22691);
xnor U36046 (N_36046,N_22310,N_20226);
or U36047 (N_36047,N_28088,N_27433);
nor U36048 (N_36048,N_21142,N_25155);
or U36049 (N_36049,N_29514,N_26164);
nor U36050 (N_36050,N_27269,N_21271);
xor U36051 (N_36051,N_29232,N_23300);
nand U36052 (N_36052,N_24928,N_22382);
or U36053 (N_36053,N_28470,N_24087);
nand U36054 (N_36054,N_27245,N_29125);
nor U36055 (N_36055,N_26043,N_25168);
xor U36056 (N_36056,N_21564,N_26004);
or U36057 (N_36057,N_29971,N_23829);
nor U36058 (N_36058,N_26262,N_23562);
xnor U36059 (N_36059,N_22871,N_27505);
nand U36060 (N_36060,N_21548,N_23107);
nor U36061 (N_36061,N_26220,N_29918);
or U36062 (N_36062,N_20279,N_27107);
xnor U36063 (N_36063,N_20667,N_20196);
nand U36064 (N_36064,N_21062,N_24612);
nand U36065 (N_36065,N_22606,N_29625);
xnor U36066 (N_36066,N_26798,N_23236);
or U36067 (N_36067,N_28021,N_26148);
xnor U36068 (N_36068,N_22750,N_26663);
and U36069 (N_36069,N_21803,N_22119);
and U36070 (N_36070,N_25060,N_25423);
nand U36071 (N_36071,N_22608,N_20169);
or U36072 (N_36072,N_23389,N_28663);
xnor U36073 (N_36073,N_21419,N_27646);
xor U36074 (N_36074,N_23113,N_28378);
and U36075 (N_36075,N_22750,N_29354);
or U36076 (N_36076,N_27508,N_21444);
nand U36077 (N_36077,N_25754,N_21193);
nor U36078 (N_36078,N_20331,N_21541);
xnor U36079 (N_36079,N_27928,N_22994);
nand U36080 (N_36080,N_29894,N_28612);
or U36081 (N_36081,N_26207,N_22309);
xor U36082 (N_36082,N_24279,N_21331);
nor U36083 (N_36083,N_22425,N_20859);
xor U36084 (N_36084,N_25897,N_22088);
or U36085 (N_36085,N_24296,N_25111);
nand U36086 (N_36086,N_28231,N_25247);
nand U36087 (N_36087,N_28471,N_28712);
and U36088 (N_36088,N_21526,N_26621);
nor U36089 (N_36089,N_27162,N_23915);
xnor U36090 (N_36090,N_26013,N_24686);
and U36091 (N_36091,N_25179,N_20794);
or U36092 (N_36092,N_26349,N_28497);
nand U36093 (N_36093,N_22427,N_26470);
or U36094 (N_36094,N_22529,N_23989);
and U36095 (N_36095,N_26499,N_21374);
and U36096 (N_36096,N_28873,N_22870);
xor U36097 (N_36097,N_26307,N_24000);
nand U36098 (N_36098,N_27049,N_23113);
or U36099 (N_36099,N_28810,N_26201);
and U36100 (N_36100,N_28335,N_23964);
xnor U36101 (N_36101,N_22485,N_21144);
or U36102 (N_36102,N_23203,N_29908);
and U36103 (N_36103,N_25476,N_24490);
nor U36104 (N_36104,N_20296,N_20964);
and U36105 (N_36105,N_25048,N_24112);
xor U36106 (N_36106,N_21449,N_27345);
nor U36107 (N_36107,N_22493,N_27088);
nor U36108 (N_36108,N_23556,N_24231);
or U36109 (N_36109,N_24733,N_25708);
and U36110 (N_36110,N_23056,N_20832);
or U36111 (N_36111,N_20889,N_29908);
or U36112 (N_36112,N_28437,N_26409);
or U36113 (N_36113,N_28130,N_21703);
nor U36114 (N_36114,N_22422,N_27101);
xor U36115 (N_36115,N_24719,N_27370);
or U36116 (N_36116,N_24960,N_20644);
xnor U36117 (N_36117,N_20146,N_24322);
and U36118 (N_36118,N_24268,N_29616);
xnor U36119 (N_36119,N_28842,N_21032);
xor U36120 (N_36120,N_25460,N_21423);
or U36121 (N_36121,N_23994,N_29131);
nor U36122 (N_36122,N_26931,N_25217);
xor U36123 (N_36123,N_29736,N_25130);
xnor U36124 (N_36124,N_21053,N_22054);
and U36125 (N_36125,N_28252,N_29554);
nand U36126 (N_36126,N_24221,N_24096);
nor U36127 (N_36127,N_23511,N_20453);
nor U36128 (N_36128,N_29947,N_26189);
nor U36129 (N_36129,N_29629,N_28092);
and U36130 (N_36130,N_23668,N_21385);
nand U36131 (N_36131,N_21708,N_21536);
xor U36132 (N_36132,N_27534,N_25247);
nand U36133 (N_36133,N_23752,N_23474);
nand U36134 (N_36134,N_25351,N_25172);
and U36135 (N_36135,N_25928,N_22214);
xor U36136 (N_36136,N_28063,N_28136);
or U36137 (N_36137,N_28029,N_24150);
nor U36138 (N_36138,N_23367,N_26440);
nand U36139 (N_36139,N_21158,N_20614);
xnor U36140 (N_36140,N_29619,N_26248);
and U36141 (N_36141,N_28926,N_23518);
and U36142 (N_36142,N_24343,N_20391);
nor U36143 (N_36143,N_20143,N_23650);
and U36144 (N_36144,N_29386,N_28287);
nand U36145 (N_36145,N_24494,N_20063);
or U36146 (N_36146,N_21803,N_20567);
or U36147 (N_36147,N_20936,N_23917);
or U36148 (N_36148,N_27504,N_28058);
nor U36149 (N_36149,N_21468,N_27288);
xor U36150 (N_36150,N_26898,N_20428);
nor U36151 (N_36151,N_21866,N_28594);
nor U36152 (N_36152,N_24287,N_24395);
or U36153 (N_36153,N_28958,N_22705);
nor U36154 (N_36154,N_23142,N_23233);
xor U36155 (N_36155,N_22579,N_25822);
and U36156 (N_36156,N_27191,N_28984);
or U36157 (N_36157,N_24836,N_22415);
xor U36158 (N_36158,N_26208,N_20226);
or U36159 (N_36159,N_29640,N_25839);
or U36160 (N_36160,N_27058,N_26805);
and U36161 (N_36161,N_28584,N_25901);
nand U36162 (N_36162,N_26106,N_29901);
or U36163 (N_36163,N_20264,N_28061);
or U36164 (N_36164,N_29487,N_23913);
xnor U36165 (N_36165,N_27158,N_20585);
or U36166 (N_36166,N_26805,N_24403);
and U36167 (N_36167,N_21763,N_22851);
and U36168 (N_36168,N_24800,N_25310);
or U36169 (N_36169,N_23551,N_20566);
xor U36170 (N_36170,N_20671,N_23138);
nor U36171 (N_36171,N_28461,N_24776);
nand U36172 (N_36172,N_24680,N_28317);
and U36173 (N_36173,N_20166,N_26776);
xnor U36174 (N_36174,N_22741,N_23446);
and U36175 (N_36175,N_25893,N_27804);
and U36176 (N_36176,N_28166,N_21809);
and U36177 (N_36177,N_25086,N_25536);
or U36178 (N_36178,N_27473,N_20970);
xor U36179 (N_36179,N_28202,N_26738);
nor U36180 (N_36180,N_26988,N_22051);
xor U36181 (N_36181,N_24946,N_28736);
nor U36182 (N_36182,N_28009,N_25928);
nor U36183 (N_36183,N_29622,N_24416);
and U36184 (N_36184,N_25340,N_27043);
or U36185 (N_36185,N_24913,N_29430);
nand U36186 (N_36186,N_28406,N_22287);
xnor U36187 (N_36187,N_28880,N_23398);
nand U36188 (N_36188,N_26180,N_20852);
xnor U36189 (N_36189,N_24456,N_27409);
nand U36190 (N_36190,N_20002,N_26037);
nand U36191 (N_36191,N_28655,N_24256);
nand U36192 (N_36192,N_23784,N_27165);
and U36193 (N_36193,N_23898,N_21609);
and U36194 (N_36194,N_22396,N_24944);
nor U36195 (N_36195,N_23124,N_25108);
nand U36196 (N_36196,N_28470,N_26269);
and U36197 (N_36197,N_25032,N_21450);
and U36198 (N_36198,N_28277,N_24900);
nand U36199 (N_36199,N_25043,N_26661);
xnor U36200 (N_36200,N_22868,N_26949);
and U36201 (N_36201,N_25758,N_20300);
nor U36202 (N_36202,N_26415,N_28496);
xnor U36203 (N_36203,N_29760,N_20943);
nor U36204 (N_36204,N_23716,N_28155);
and U36205 (N_36205,N_25548,N_24591);
xor U36206 (N_36206,N_27040,N_27493);
or U36207 (N_36207,N_24775,N_29312);
or U36208 (N_36208,N_29994,N_28874);
nand U36209 (N_36209,N_22530,N_24229);
or U36210 (N_36210,N_27720,N_21933);
or U36211 (N_36211,N_26898,N_20760);
and U36212 (N_36212,N_20451,N_23702);
nand U36213 (N_36213,N_25483,N_27702);
xor U36214 (N_36214,N_28585,N_20719);
xor U36215 (N_36215,N_22293,N_23842);
or U36216 (N_36216,N_28551,N_23022);
nand U36217 (N_36217,N_25483,N_23243);
and U36218 (N_36218,N_25758,N_26759);
and U36219 (N_36219,N_24114,N_20627);
nor U36220 (N_36220,N_21069,N_23166);
nor U36221 (N_36221,N_23516,N_25343);
and U36222 (N_36222,N_22822,N_24272);
and U36223 (N_36223,N_22334,N_29831);
xnor U36224 (N_36224,N_28629,N_25732);
or U36225 (N_36225,N_25391,N_21800);
xnor U36226 (N_36226,N_20029,N_28793);
or U36227 (N_36227,N_29607,N_22995);
nor U36228 (N_36228,N_22828,N_28191);
xnor U36229 (N_36229,N_20716,N_26435);
nand U36230 (N_36230,N_28656,N_29900);
and U36231 (N_36231,N_28872,N_23263);
nand U36232 (N_36232,N_21962,N_26645);
xnor U36233 (N_36233,N_20554,N_26560);
xor U36234 (N_36234,N_22025,N_20972);
or U36235 (N_36235,N_27081,N_24004);
xnor U36236 (N_36236,N_24165,N_22918);
and U36237 (N_36237,N_28447,N_22738);
or U36238 (N_36238,N_21461,N_20714);
nand U36239 (N_36239,N_24684,N_29686);
nor U36240 (N_36240,N_29537,N_26004);
xnor U36241 (N_36241,N_21786,N_27451);
nand U36242 (N_36242,N_20311,N_25447);
nand U36243 (N_36243,N_21592,N_20498);
nor U36244 (N_36244,N_25818,N_22727);
nor U36245 (N_36245,N_21432,N_22778);
and U36246 (N_36246,N_23107,N_26143);
xnor U36247 (N_36247,N_20340,N_21663);
nand U36248 (N_36248,N_22210,N_21709);
or U36249 (N_36249,N_21472,N_20522);
nor U36250 (N_36250,N_28023,N_20461);
or U36251 (N_36251,N_29043,N_20506);
or U36252 (N_36252,N_20350,N_28449);
or U36253 (N_36253,N_27013,N_21325);
nor U36254 (N_36254,N_21076,N_20813);
or U36255 (N_36255,N_23354,N_23825);
or U36256 (N_36256,N_28129,N_24944);
or U36257 (N_36257,N_21653,N_29183);
xnor U36258 (N_36258,N_20999,N_24419);
nor U36259 (N_36259,N_26873,N_27486);
nand U36260 (N_36260,N_20165,N_21709);
xnor U36261 (N_36261,N_21992,N_26040);
xnor U36262 (N_36262,N_23153,N_22754);
nand U36263 (N_36263,N_28136,N_25333);
nor U36264 (N_36264,N_21935,N_21792);
nor U36265 (N_36265,N_22635,N_29755);
nor U36266 (N_36266,N_22531,N_24973);
and U36267 (N_36267,N_29151,N_27035);
and U36268 (N_36268,N_21223,N_20104);
and U36269 (N_36269,N_20446,N_20221);
nand U36270 (N_36270,N_24127,N_29224);
xnor U36271 (N_36271,N_23054,N_26386);
and U36272 (N_36272,N_28547,N_26473);
nor U36273 (N_36273,N_26245,N_25642);
nor U36274 (N_36274,N_24453,N_23771);
or U36275 (N_36275,N_24517,N_20797);
xnor U36276 (N_36276,N_22246,N_26985);
nand U36277 (N_36277,N_21026,N_20180);
or U36278 (N_36278,N_23010,N_21336);
xor U36279 (N_36279,N_21646,N_20262);
or U36280 (N_36280,N_26986,N_26419);
nor U36281 (N_36281,N_28941,N_23145);
xnor U36282 (N_36282,N_25434,N_25237);
or U36283 (N_36283,N_20830,N_27116);
nand U36284 (N_36284,N_27536,N_26577);
or U36285 (N_36285,N_20437,N_26924);
nand U36286 (N_36286,N_27929,N_27148);
xnor U36287 (N_36287,N_22483,N_24373);
xnor U36288 (N_36288,N_26832,N_27634);
nor U36289 (N_36289,N_26651,N_22616);
nand U36290 (N_36290,N_24290,N_28879);
and U36291 (N_36291,N_23702,N_22459);
nand U36292 (N_36292,N_23384,N_24021);
and U36293 (N_36293,N_28745,N_25416);
nor U36294 (N_36294,N_20916,N_23068);
xnor U36295 (N_36295,N_29547,N_24723);
or U36296 (N_36296,N_23928,N_22646);
xor U36297 (N_36297,N_26797,N_24830);
or U36298 (N_36298,N_23693,N_24120);
and U36299 (N_36299,N_29555,N_25002);
nand U36300 (N_36300,N_22775,N_27417);
nor U36301 (N_36301,N_27717,N_25552);
or U36302 (N_36302,N_22717,N_20603);
or U36303 (N_36303,N_21096,N_21498);
xor U36304 (N_36304,N_21400,N_21900);
xnor U36305 (N_36305,N_24462,N_27829);
and U36306 (N_36306,N_24622,N_20792);
nand U36307 (N_36307,N_22082,N_27878);
xnor U36308 (N_36308,N_27989,N_21410);
nand U36309 (N_36309,N_27893,N_20958);
nand U36310 (N_36310,N_28883,N_20962);
nand U36311 (N_36311,N_25950,N_25309);
xnor U36312 (N_36312,N_27314,N_29299);
or U36313 (N_36313,N_20143,N_27693);
nor U36314 (N_36314,N_29758,N_24843);
and U36315 (N_36315,N_24644,N_27041);
xnor U36316 (N_36316,N_23460,N_28649);
nor U36317 (N_36317,N_26941,N_27876);
and U36318 (N_36318,N_23616,N_22353);
nand U36319 (N_36319,N_25203,N_25456);
nor U36320 (N_36320,N_26327,N_27432);
xor U36321 (N_36321,N_27135,N_29722);
nor U36322 (N_36322,N_23323,N_25993);
and U36323 (N_36323,N_27864,N_26957);
nand U36324 (N_36324,N_28453,N_20033);
nor U36325 (N_36325,N_26894,N_29177);
nand U36326 (N_36326,N_23284,N_24993);
or U36327 (N_36327,N_24474,N_26725);
xnor U36328 (N_36328,N_23670,N_28305);
and U36329 (N_36329,N_22425,N_20512);
xnor U36330 (N_36330,N_20461,N_23957);
nand U36331 (N_36331,N_29135,N_25749);
xnor U36332 (N_36332,N_29230,N_21594);
nand U36333 (N_36333,N_26291,N_23399);
xor U36334 (N_36334,N_22936,N_27762);
xnor U36335 (N_36335,N_24036,N_22256);
xnor U36336 (N_36336,N_27198,N_28973);
nor U36337 (N_36337,N_28693,N_27525);
nand U36338 (N_36338,N_27029,N_25288);
and U36339 (N_36339,N_23810,N_23060);
nand U36340 (N_36340,N_28378,N_21603);
nor U36341 (N_36341,N_22422,N_20632);
nor U36342 (N_36342,N_20744,N_27548);
nor U36343 (N_36343,N_26682,N_23428);
and U36344 (N_36344,N_28703,N_23813);
nand U36345 (N_36345,N_27192,N_23293);
and U36346 (N_36346,N_26994,N_22317);
xnor U36347 (N_36347,N_27272,N_27531);
or U36348 (N_36348,N_27325,N_23117);
xnor U36349 (N_36349,N_28966,N_23688);
xor U36350 (N_36350,N_28854,N_21616);
nor U36351 (N_36351,N_27934,N_28869);
or U36352 (N_36352,N_29566,N_29351);
nand U36353 (N_36353,N_25329,N_27647);
and U36354 (N_36354,N_22987,N_23760);
xnor U36355 (N_36355,N_23385,N_28950);
nand U36356 (N_36356,N_24719,N_28636);
or U36357 (N_36357,N_26598,N_24424);
and U36358 (N_36358,N_27152,N_23913);
nor U36359 (N_36359,N_29723,N_24338);
xor U36360 (N_36360,N_24461,N_27601);
nand U36361 (N_36361,N_28286,N_26212);
nand U36362 (N_36362,N_23379,N_23422);
and U36363 (N_36363,N_25280,N_26465);
nor U36364 (N_36364,N_21227,N_27397);
and U36365 (N_36365,N_25439,N_26231);
and U36366 (N_36366,N_22489,N_20723);
nand U36367 (N_36367,N_29949,N_25561);
and U36368 (N_36368,N_26176,N_29836);
nor U36369 (N_36369,N_22476,N_26426);
and U36370 (N_36370,N_21684,N_23513);
nand U36371 (N_36371,N_27298,N_27548);
or U36372 (N_36372,N_23578,N_29385);
and U36373 (N_36373,N_20138,N_23092);
nand U36374 (N_36374,N_24070,N_28251);
or U36375 (N_36375,N_28343,N_20451);
or U36376 (N_36376,N_29795,N_22327);
xnor U36377 (N_36377,N_21825,N_27910);
or U36378 (N_36378,N_29563,N_29031);
nand U36379 (N_36379,N_21489,N_27702);
nor U36380 (N_36380,N_29312,N_23795);
nor U36381 (N_36381,N_26256,N_20802);
and U36382 (N_36382,N_23434,N_26103);
or U36383 (N_36383,N_24227,N_21253);
nor U36384 (N_36384,N_27355,N_25622);
xnor U36385 (N_36385,N_22289,N_25652);
nor U36386 (N_36386,N_24584,N_29002);
nand U36387 (N_36387,N_20270,N_27875);
nand U36388 (N_36388,N_25262,N_25743);
and U36389 (N_36389,N_26180,N_23449);
nand U36390 (N_36390,N_22646,N_25982);
nand U36391 (N_36391,N_21918,N_28967);
or U36392 (N_36392,N_28412,N_29622);
or U36393 (N_36393,N_22899,N_21441);
nand U36394 (N_36394,N_23587,N_23421);
nor U36395 (N_36395,N_29386,N_23132);
nand U36396 (N_36396,N_23693,N_26912);
nor U36397 (N_36397,N_27724,N_21276);
nor U36398 (N_36398,N_20469,N_20645);
and U36399 (N_36399,N_27023,N_27994);
xor U36400 (N_36400,N_20401,N_25036);
nor U36401 (N_36401,N_25775,N_24093);
and U36402 (N_36402,N_23530,N_22128);
or U36403 (N_36403,N_25144,N_28377);
nand U36404 (N_36404,N_25552,N_27168);
nor U36405 (N_36405,N_20371,N_25590);
and U36406 (N_36406,N_21914,N_21998);
nor U36407 (N_36407,N_25614,N_20590);
xnor U36408 (N_36408,N_21066,N_27211);
and U36409 (N_36409,N_20583,N_23332);
and U36410 (N_36410,N_28503,N_23637);
or U36411 (N_36411,N_29239,N_21511);
and U36412 (N_36412,N_29996,N_27263);
nand U36413 (N_36413,N_21574,N_20355);
nand U36414 (N_36414,N_26746,N_29152);
nor U36415 (N_36415,N_25383,N_28019);
nor U36416 (N_36416,N_28655,N_22799);
nor U36417 (N_36417,N_20141,N_23936);
nand U36418 (N_36418,N_24332,N_26880);
and U36419 (N_36419,N_28092,N_28561);
nor U36420 (N_36420,N_25911,N_23892);
nor U36421 (N_36421,N_29891,N_24860);
and U36422 (N_36422,N_25124,N_23327);
nor U36423 (N_36423,N_23823,N_23444);
xor U36424 (N_36424,N_26249,N_21028);
nor U36425 (N_36425,N_27761,N_27911);
and U36426 (N_36426,N_26171,N_25318);
nor U36427 (N_36427,N_21579,N_21765);
xnor U36428 (N_36428,N_27816,N_21800);
nand U36429 (N_36429,N_21852,N_29804);
or U36430 (N_36430,N_20070,N_20758);
xnor U36431 (N_36431,N_29851,N_21928);
xnor U36432 (N_36432,N_21301,N_22514);
nand U36433 (N_36433,N_24117,N_23369);
or U36434 (N_36434,N_22503,N_25891);
nor U36435 (N_36435,N_28531,N_22232);
or U36436 (N_36436,N_23888,N_22414);
or U36437 (N_36437,N_20468,N_27918);
nor U36438 (N_36438,N_29818,N_22873);
nand U36439 (N_36439,N_20218,N_27463);
xor U36440 (N_36440,N_27770,N_29642);
nand U36441 (N_36441,N_28090,N_29847);
or U36442 (N_36442,N_24455,N_26670);
or U36443 (N_36443,N_27208,N_26992);
xnor U36444 (N_36444,N_28067,N_29801);
nand U36445 (N_36445,N_25523,N_21535);
xnor U36446 (N_36446,N_26059,N_20983);
nor U36447 (N_36447,N_26696,N_28713);
and U36448 (N_36448,N_22748,N_22466);
or U36449 (N_36449,N_24600,N_28767);
nor U36450 (N_36450,N_21890,N_21587);
nor U36451 (N_36451,N_21644,N_23287);
or U36452 (N_36452,N_28844,N_27708);
nand U36453 (N_36453,N_26887,N_26142);
nor U36454 (N_36454,N_21409,N_22222);
nand U36455 (N_36455,N_20387,N_29927);
and U36456 (N_36456,N_26672,N_25410);
nor U36457 (N_36457,N_25796,N_20750);
or U36458 (N_36458,N_29235,N_29925);
and U36459 (N_36459,N_22939,N_29774);
nor U36460 (N_36460,N_26484,N_24818);
xor U36461 (N_36461,N_22208,N_24053);
nor U36462 (N_36462,N_21968,N_23688);
or U36463 (N_36463,N_24520,N_20764);
nor U36464 (N_36464,N_26252,N_28828);
or U36465 (N_36465,N_28927,N_22434);
nor U36466 (N_36466,N_24550,N_24151);
xnor U36467 (N_36467,N_25782,N_26592);
xnor U36468 (N_36468,N_23502,N_27817);
xor U36469 (N_36469,N_27673,N_24765);
xor U36470 (N_36470,N_23942,N_25275);
nor U36471 (N_36471,N_21440,N_22952);
nor U36472 (N_36472,N_21657,N_26246);
nor U36473 (N_36473,N_21128,N_20577);
or U36474 (N_36474,N_27506,N_29935);
or U36475 (N_36475,N_21061,N_27558);
nand U36476 (N_36476,N_23197,N_27790);
or U36477 (N_36477,N_27908,N_26033);
nand U36478 (N_36478,N_26113,N_23734);
nand U36479 (N_36479,N_22414,N_24599);
xnor U36480 (N_36480,N_26397,N_29319);
nand U36481 (N_36481,N_29188,N_21074);
nand U36482 (N_36482,N_24645,N_26336);
and U36483 (N_36483,N_20381,N_26546);
or U36484 (N_36484,N_27328,N_22163);
and U36485 (N_36485,N_20039,N_20549);
nor U36486 (N_36486,N_27011,N_22352);
nand U36487 (N_36487,N_21579,N_25728);
and U36488 (N_36488,N_24129,N_24011);
xor U36489 (N_36489,N_22950,N_28593);
or U36490 (N_36490,N_27657,N_29280);
or U36491 (N_36491,N_26858,N_26707);
nand U36492 (N_36492,N_26189,N_20213);
nand U36493 (N_36493,N_20163,N_25275);
or U36494 (N_36494,N_26906,N_27742);
nor U36495 (N_36495,N_25921,N_29014);
or U36496 (N_36496,N_22637,N_25926);
nor U36497 (N_36497,N_21519,N_24704);
xor U36498 (N_36498,N_26615,N_28683);
nand U36499 (N_36499,N_22223,N_21312);
or U36500 (N_36500,N_28904,N_29534);
nor U36501 (N_36501,N_22421,N_28502);
xnor U36502 (N_36502,N_20389,N_21858);
and U36503 (N_36503,N_24316,N_29278);
xor U36504 (N_36504,N_27196,N_23469);
nor U36505 (N_36505,N_20922,N_23252);
nand U36506 (N_36506,N_22750,N_24905);
and U36507 (N_36507,N_27114,N_25361);
nand U36508 (N_36508,N_25002,N_21930);
xor U36509 (N_36509,N_24877,N_20919);
and U36510 (N_36510,N_27449,N_20234);
and U36511 (N_36511,N_26483,N_23904);
or U36512 (N_36512,N_24613,N_21501);
or U36513 (N_36513,N_29801,N_25128);
or U36514 (N_36514,N_27547,N_23884);
xor U36515 (N_36515,N_26716,N_21647);
and U36516 (N_36516,N_23629,N_22442);
nand U36517 (N_36517,N_23332,N_29950);
xnor U36518 (N_36518,N_29722,N_29380);
or U36519 (N_36519,N_28826,N_20312);
nor U36520 (N_36520,N_20523,N_28974);
or U36521 (N_36521,N_29269,N_22843);
nor U36522 (N_36522,N_21412,N_26341);
nor U36523 (N_36523,N_23127,N_22803);
xnor U36524 (N_36524,N_22057,N_29697);
and U36525 (N_36525,N_26680,N_26060);
nand U36526 (N_36526,N_29162,N_27660);
xnor U36527 (N_36527,N_29579,N_25085);
or U36528 (N_36528,N_21286,N_25364);
xnor U36529 (N_36529,N_23924,N_25565);
and U36530 (N_36530,N_22678,N_21971);
nand U36531 (N_36531,N_24812,N_21110);
nor U36532 (N_36532,N_26238,N_29849);
or U36533 (N_36533,N_22108,N_21627);
nor U36534 (N_36534,N_29209,N_27575);
nor U36535 (N_36535,N_27549,N_23473);
nor U36536 (N_36536,N_21760,N_24601);
and U36537 (N_36537,N_22093,N_29044);
nand U36538 (N_36538,N_28463,N_23118);
xnor U36539 (N_36539,N_26564,N_26107);
nor U36540 (N_36540,N_29510,N_28955);
nand U36541 (N_36541,N_26054,N_29024);
xnor U36542 (N_36542,N_26774,N_21599);
nor U36543 (N_36543,N_25986,N_21845);
and U36544 (N_36544,N_26321,N_29785);
or U36545 (N_36545,N_26617,N_25753);
xor U36546 (N_36546,N_27721,N_24716);
nand U36547 (N_36547,N_25661,N_21673);
nand U36548 (N_36548,N_29719,N_23591);
xor U36549 (N_36549,N_20755,N_24868);
nand U36550 (N_36550,N_25608,N_26458);
xnor U36551 (N_36551,N_28752,N_23191);
nand U36552 (N_36552,N_28734,N_24624);
and U36553 (N_36553,N_25129,N_27042);
or U36554 (N_36554,N_20395,N_22235);
nor U36555 (N_36555,N_28126,N_23206);
xor U36556 (N_36556,N_25581,N_25269);
or U36557 (N_36557,N_23350,N_25402);
nor U36558 (N_36558,N_24709,N_22044);
nor U36559 (N_36559,N_22195,N_27413);
nor U36560 (N_36560,N_28601,N_26716);
and U36561 (N_36561,N_27487,N_27917);
nand U36562 (N_36562,N_27315,N_28648);
or U36563 (N_36563,N_27939,N_28805);
xnor U36564 (N_36564,N_24627,N_23430);
xnor U36565 (N_36565,N_20412,N_26805);
nand U36566 (N_36566,N_26321,N_26091);
or U36567 (N_36567,N_21710,N_20105);
nor U36568 (N_36568,N_26435,N_27376);
or U36569 (N_36569,N_21935,N_27161);
nand U36570 (N_36570,N_25122,N_29578);
and U36571 (N_36571,N_22090,N_20706);
or U36572 (N_36572,N_27737,N_27919);
nand U36573 (N_36573,N_28527,N_27312);
and U36574 (N_36574,N_20315,N_27324);
xnor U36575 (N_36575,N_28530,N_27384);
or U36576 (N_36576,N_23503,N_28586);
nor U36577 (N_36577,N_23071,N_27845);
xnor U36578 (N_36578,N_28027,N_23315);
or U36579 (N_36579,N_28797,N_20214);
and U36580 (N_36580,N_21986,N_26382);
nor U36581 (N_36581,N_26241,N_21591);
or U36582 (N_36582,N_26432,N_25276);
nand U36583 (N_36583,N_25382,N_26712);
nand U36584 (N_36584,N_29201,N_24696);
nor U36585 (N_36585,N_22929,N_28248);
nor U36586 (N_36586,N_25216,N_29359);
nand U36587 (N_36587,N_25435,N_24317);
nand U36588 (N_36588,N_29437,N_29036);
nor U36589 (N_36589,N_21198,N_24686);
and U36590 (N_36590,N_23956,N_24573);
nand U36591 (N_36591,N_25894,N_24797);
or U36592 (N_36592,N_29761,N_25506);
and U36593 (N_36593,N_23305,N_28428);
and U36594 (N_36594,N_27288,N_22460);
nand U36595 (N_36595,N_25715,N_27687);
nand U36596 (N_36596,N_29334,N_27993);
nand U36597 (N_36597,N_29494,N_26131);
nor U36598 (N_36598,N_20253,N_28062);
xnor U36599 (N_36599,N_21235,N_27297);
or U36600 (N_36600,N_28888,N_26989);
and U36601 (N_36601,N_21170,N_24318);
and U36602 (N_36602,N_29784,N_24156);
and U36603 (N_36603,N_23369,N_29262);
or U36604 (N_36604,N_27882,N_26629);
xnor U36605 (N_36605,N_29058,N_20350);
nand U36606 (N_36606,N_23735,N_28817);
nand U36607 (N_36607,N_28786,N_28686);
or U36608 (N_36608,N_25813,N_28859);
and U36609 (N_36609,N_28596,N_24365);
and U36610 (N_36610,N_26879,N_21792);
or U36611 (N_36611,N_21878,N_24430);
nand U36612 (N_36612,N_29798,N_20348);
nand U36613 (N_36613,N_26811,N_21813);
nand U36614 (N_36614,N_22428,N_22427);
or U36615 (N_36615,N_29828,N_24806);
and U36616 (N_36616,N_24736,N_28801);
xor U36617 (N_36617,N_20155,N_24128);
and U36618 (N_36618,N_21053,N_25605);
or U36619 (N_36619,N_28578,N_20900);
and U36620 (N_36620,N_24091,N_20574);
nor U36621 (N_36621,N_21963,N_23599);
and U36622 (N_36622,N_24826,N_24970);
and U36623 (N_36623,N_23390,N_20208);
nor U36624 (N_36624,N_20821,N_23565);
nand U36625 (N_36625,N_22629,N_23118);
nor U36626 (N_36626,N_23726,N_26881);
or U36627 (N_36627,N_27785,N_29618);
or U36628 (N_36628,N_23689,N_24576);
and U36629 (N_36629,N_25682,N_24665);
xor U36630 (N_36630,N_26667,N_22981);
or U36631 (N_36631,N_21344,N_26523);
or U36632 (N_36632,N_24598,N_29547);
xnor U36633 (N_36633,N_29548,N_27518);
or U36634 (N_36634,N_27580,N_21399);
and U36635 (N_36635,N_23932,N_29419);
and U36636 (N_36636,N_21647,N_29346);
and U36637 (N_36637,N_24534,N_28151);
nor U36638 (N_36638,N_21103,N_26392);
xnor U36639 (N_36639,N_24988,N_25618);
nor U36640 (N_36640,N_24462,N_26604);
xnor U36641 (N_36641,N_28515,N_25735);
nor U36642 (N_36642,N_28614,N_22061);
xnor U36643 (N_36643,N_25589,N_22341);
and U36644 (N_36644,N_25195,N_27891);
nand U36645 (N_36645,N_23139,N_20331);
or U36646 (N_36646,N_21734,N_27225);
and U36647 (N_36647,N_26874,N_24231);
nor U36648 (N_36648,N_23814,N_28041);
and U36649 (N_36649,N_20411,N_29516);
xnor U36650 (N_36650,N_24373,N_24354);
or U36651 (N_36651,N_24939,N_28934);
xor U36652 (N_36652,N_22514,N_20881);
nand U36653 (N_36653,N_24649,N_21245);
or U36654 (N_36654,N_25890,N_26749);
nor U36655 (N_36655,N_29572,N_27053);
nand U36656 (N_36656,N_28304,N_22608);
and U36657 (N_36657,N_23672,N_28259);
nand U36658 (N_36658,N_21304,N_22119);
or U36659 (N_36659,N_24562,N_23627);
nor U36660 (N_36660,N_26610,N_20781);
and U36661 (N_36661,N_25289,N_27416);
nand U36662 (N_36662,N_26256,N_22812);
nor U36663 (N_36663,N_22158,N_27907);
and U36664 (N_36664,N_23454,N_20736);
xnor U36665 (N_36665,N_26316,N_23864);
xor U36666 (N_36666,N_26301,N_24490);
or U36667 (N_36667,N_28152,N_24246);
nand U36668 (N_36668,N_24872,N_28566);
nor U36669 (N_36669,N_26713,N_24565);
nor U36670 (N_36670,N_28101,N_26222);
and U36671 (N_36671,N_26387,N_20753);
xor U36672 (N_36672,N_27368,N_27646);
xnor U36673 (N_36673,N_22442,N_20847);
or U36674 (N_36674,N_27622,N_27402);
and U36675 (N_36675,N_29763,N_29685);
xnor U36676 (N_36676,N_26519,N_22689);
and U36677 (N_36677,N_21299,N_28786);
or U36678 (N_36678,N_29047,N_26014);
and U36679 (N_36679,N_29522,N_28354);
nor U36680 (N_36680,N_20731,N_24015);
nand U36681 (N_36681,N_24778,N_23683);
and U36682 (N_36682,N_22067,N_29869);
and U36683 (N_36683,N_29529,N_24504);
and U36684 (N_36684,N_21295,N_24695);
nor U36685 (N_36685,N_27226,N_29513);
xnor U36686 (N_36686,N_22022,N_27096);
nor U36687 (N_36687,N_28651,N_25086);
nor U36688 (N_36688,N_28593,N_24686);
or U36689 (N_36689,N_28801,N_23954);
and U36690 (N_36690,N_24430,N_27207);
or U36691 (N_36691,N_26900,N_26732);
nand U36692 (N_36692,N_29221,N_21406);
xor U36693 (N_36693,N_25868,N_26884);
nand U36694 (N_36694,N_24291,N_24910);
xor U36695 (N_36695,N_27611,N_26618);
xnor U36696 (N_36696,N_21187,N_20798);
nor U36697 (N_36697,N_20467,N_22307);
and U36698 (N_36698,N_28206,N_25158);
and U36699 (N_36699,N_25295,N_24100);
xnor U36700 (N_36700,N_28892,N_25620);
nor U36701 (N_36701,N_27846,N_29584);
and U36702 (N_36702,N_27363,N_28670);
or U36703 (N_36703,N_23665,N_24157);
and U36704 (N_36704,N_21101,N_23440);
xor U36705 (N_36705,N_21291,N_25155);
and U36706 (N_36706,N_20449,N_28636);
and U36707 (N_36707,N_22312,N_27381);
or U36708 (N_36708,N_21773,N_21337);
and U36709 (N_36709,N_25539,N_29163);
xor U36710 (N_36710,N_23416,N_27881);
or U36711 (N_36711,N_25158,N_23575);
nor U36712 (N_36712,N_28638,N_23638);
nor U36713 (N_36713,N_24167,N_27803);
nor U36714 (N_36714,N_24806,N_21633);
nor U36715 (N_36715,N_29235,N_29059);
or U36716 (N_36716,N_21780,N_28266);
nand U36717 (N_36717,N_24029,N_24831);
and U36718 (N_36718,N_24514,N_29706);
xor U36719 (N_36719,N_23262,N_21532);
or U36720 (N_36720,N_23581,N_26430);
or U36721 (N_36721,N_26114,N_28928);
nor U36722 (N_36722,N_23476,N_27065);
or U36723 (N_36723,N_20926,N_26710);
nor U36724 (N_36724,N_26244,N_24400);
nor U36725 (N_36725,N_25661,N_29199);
and U36726 (N_36726,N_22800,N_27316);
nand U36727 (N_36727,N_21435,N_21109);
nand U36728 (N_36728,N_22557,N_28432);
nand U36729 (N_36729,N_23647,N_24517);
or U36730 (N_36730,N_21728,N_23623);
nor U36731 (N_36731,N_24432,N_21761);
xor U36732 (N_36732,N_24233,N_28186);
or U36733 (N_36733,N_22853,N_20920);
xnor U36734 (N_36734,N_28957,N_23963);
xor U36735 (N_36735,N_21149,N_26204);
and U36736 (N_36736,N_23361,N_28036);
nand U36737 (N_36737,N_26642,N_25985);
or U36738 (N_36738,N_27428,N_27734);
nor U36739 (N_36739,N_29524,N_24767);
xor U36740 (N_36740,N_21188,N_29066);
and U36741 (N_36741,N_24053,N_23780);
nand U36742 (N_36742,N_23960,N_20993);
or U36743 (N_36743,N_20026,N_20319);
or U36744 (N_36744,N_21501,N_23421);
nor U36745 (N_36745,N_27575,N_28431);
and U36746 (N_36746,N_24892,N_21855);
and U36747 (N_36747,N_29804,N_22922);
nand U36748 (N_36748,N_23729,N_25226);
xor U36749 (N_36749,N_20995,N_26544);
nand U36750 (N_36750,N_23376,N_21951);
nor U36751 (N_36751,N_21100,N_20124);
xnor U36752 (N_36752,N_24574,N_21310);
or U36753 (N_36753,N_23269,N_29949);
xor U36754 (N_36754,N_21374,N_23987);
or U36755 (N_36755,N_23218,N_26468);
nand U36756 (N_36756,N_20781,N_28292);
and U36757 (N_36757,N_21695,N_20321);
or U36758 (N_36758,N_24312,N_28447);
nor U36759 (N_36759,N_26712,N_29830);
xnor U36760 (N_36760,N_23206,N_27451);
nor U36761 (N_36761,N_26232,N_23318);
or U36762 (N_36762,N_24113,N_26576);
or U36763 (N_36763,N_22257,N_26016);
or U36764 (N_36764,N_27614,N_24510);
and U36765 (N_36765,N_29766,N_21732);
nand U36766 (N_36766,N_29006,N_27028);
nand U36767 (N_36767,N_25302,N_26056);
or U36768 (N_36768,N_24726,N_20128);
xor U36769 (N_36769,N_21096,N_22613);
nand U36770 (N_36770,N_24046,N_28982);
xor U36771 (N_36771,N_24082,N_26975);
and U36772 (N_36772,N_23182,N_26303);
and U36773 (N_36773,N_29548,N_23835);
xnor U36774 (N_36774,N_22564,N_28508);
nor U36775 (N_36775,N_23897,N_27147);
xnor U36776 (N_36776,N_26538,N_28362);
or U36777 (N_36777,N_29043,N_23137);
or U36778 (N_36778,N_22750,N_23793);
nor U36779 (N_36779,N_26517,N_23459);
xnor U36780 (N_36780,N_29113,N_29751);
or U36781 (N_36781,N_25174,N_22629);
and U36782 (N_36782,N_28992,N_26902);
xor U36783 (N_36783,N_24934,N_26559);
nor U36784 (N_36784,N_26360,N_23125);
nand U36785 (N_36785,N_25645,N_28698);
nor U36786 (N_36786,N_21759,N_29362);
nor U36787 (N_36787,N_23518,N_26446);
and U36788 (N_36788,N_27403,N_21063);
and U36789 (N_36789,N_28196,N_24450);
and U36790 (N_36790,N_29628,N_21518);
and U36791 (N_36791,N_20795,N_27724);
nand U36792 (N_36792,N_27763,N_28942);
nand U36793 (N_36793,N_26966,N_29944);
xor U36794 (N_36794,N_21826,N_22308);
nand U36795 (N_36795,N_29261,N_26651);
xor U36796 (N_36796,N_21668,N_24308);
xor U36797 (N_36797,N_23447,N_26459);
nor U36798 (N_36798,N_21467,N_24843);
nand U36799 (N_36799,N_29591,N_25568);
nand U36800 (N_36800,N_28407,N_21944);
or U36801 (N_36801,N_21946,N_29143);
xnor U36802 (N_36802,N_28966,N_22604);
nand U36803 (N_36803,N_29572,N_22633);
or U36804 (N_36804,N_28896,N_21281);
xnor U36805 (N_36805,N_22318,N_21522);
nand U36806 (N_36806,N_21982,N_26670);
nor U36807 (N_36807,N_20950,N_23384);
xor U36808 (N_36808,N_21225,N_23524);
xor U36809 (N_36809,N_24508,N_20941);
or U36810 (N_36810,N_28249,N_29084);
and U36811 (N_36811,N_27497,N_28503);
or U36812 (N_36812,N_24045,N_27905);
nor U36813 (N_36813,N_28637,N_23749);
xnor U36814 (N_36814,N_25934,N_23408);
xor U36815 (N_36815,N_28476,N_26324);
xor U36816 (N_36816,N_22514,N_27972);
or U36817 (N_36817,N_27880,N_26566);
nand U36818 (N_36818,N_24027,N_23558);
or U36819 (N_36819,N_22514,N_27789);
or U36820 (N_36820,N_24574,N_22117);
nand U36821 (N_36821,N_21426,N_24541);
or U36822 (N_36822,N_24774,N_28464);
nand U36823 (N_36823,N_24007,N_25579);
nor U36824 (N_36824,N_20849,N_29098);
nor U36825 (N_36825,N_24113,N_24607);
and U36826 (N_36826,N_28271,N_21307);
or U36827 (N_36827,N_24346,N_22209);
xor U36828 (N_36828,N_25229,N_24199);
xor U36829 (N_36829,N_26808,N_27398);
xnor U36830 (N_36830,N_26963,N_25218);
nor U36831 (N_36831,N_24964,N_22014);
xnor U36832 (N_36832,N_29717,N_26851);
and U36833 (N_36833,N_22373,N_21268);
and U36834 (N_36834,N_24481,N_20508);
or U36835 (N_36835,N_29355,N_27878);
nor U36836 (N_36836,N_27819,N_28986);
and U36837 (N_36837,N_22517,N_20606);
nand U36838 (N_36838,N_27017,N_28807);
and U36839 (N_36839,N_26592,N_24762);
and U36840 (N_36840,N_26448,N_24615);
xor U36841 (N_36841,N_20153,N_23148);
nor U36842 (N_36842,N_22472,N_27137);
nor U36843 (N_36843,N_29465,N_28238);
nor U36844 (N_36844,N_22484,N_29629);
and U36845 (N_36845,N_25460,N_22713);
or U36846 (N_36846,N_22655,N_24490);
xnor U36847 (N_36847,N_24098,N_24917);
and U36848 (N_36848,N_28404,N_23804);
or U36849 (N_36849,N_25273,N_29865);
nand U36850 (N_36850,N_22976,N_23937);
or U36851 (N_36851,N_22966,N_24272);
xor U36852 (N_36852,N_21021,N_27326);
or U36853 (N_36853,N_25909,N_20776);
nand U36854 (N_36854,N_29800,N_20864);
or U36855 (N_36855,N_22945,N_22635);
xnor U36856 (N_36856,N_24387,N_25643);
or U36857 (N_36857,N_28521,N_22942);
nor U36858 (N_36858,N_27381,N_22096);
xnor U36859 (N_36859,N_24562,N_22103);
or U36860 (N_36860,N_26189,N_21451);
nand U36861 (N_36861,N_28581,N_25280);
or U36862 (N_36862,N_22251,N_23246);
nand U36863 (N_36863,N_21780,N_21573);
or U36864 (N_36864,N_21926,N_21841);
and U36865 (N_36865,N_28367,N_22756);
nor U36866 (N_36866,N_28649,N_28046);
or U36867 (N_36867,N_29444,N_21040);
xnor U36868 (N_36868,N_21656,N_20757);
and U36869 (N_36869,N_22786,N_21653);
xnor U36870 (N_36870,N_21690,N_23451);
xor U36871 (N_36871,N_27912,N_25149);
or U36872 (N_36872,N_26582,N_20096);
xor U36873 (N_36873,N_24653,N_27524);
xnor U36874 (N_36874,N_20571,N_21749);
xor U36875 (N_36875,N_24653,N_24188);
nand U36876 (N_36876,N_23530,N_23056);
and U36877 (N_36877,N_25360,N_21105);
nor U36878 (N_36878,N_24293,N_24428);
nand U36879 (N_36879,N_25649,N_22055);
nor U36880 (N_36880,N_29397,N_24666);
nand U36881 (N_36881,N_24872,N_25533);
nand U36882 (N_36882,N_28885,N_22734);
or U36883 (N_36883,N_21289,N_21551);
nor U36884 (N_36884,N_23879,N_29036);
or U36885 (N_36885,N_29551,N_23043);
nor U36886 (N_36886,N_29886,N_21992);
nand U36887 (N_36887,N_21223,N_29040);
xor U36888 (N_36888,N_28979,N_23190);
nor U36889 (N_36889,N_24990,N_22094);
nand U36890 (N_36890,N_29063,N_28028);
nor U36891 (N_36891,N_23226,N_20882);
and U36892 (N_36892,N_25151,N_20596);
xor U36893 (N_36893,N_27380,N_25220);
nor U36894 (N_36894,N_20097,N_20381);
or U36895 (N_36895,N_27439,N_23424);
nand U36896 (N_36896,N_27225,N_27007);
xnor U36897 (N_36897,N_29279,N_23383);
nor U36898 (N_36898,N_24437,N_26930);
xor U36899 (N_36899,N_23795,N_20864);
nor U36900 (N_36900,N_23389,N_29649);
nand U36901 (N_36901,N_23731,N_23710);
or U36902 (N_36902,N_25852,N_20637);
xnor U36903 (N_36903,N_27917,N_29482);
nor U36904 (N_36904,N_23938,N_20897);
nor U36905 (N_36905,N_24789,N_20835);
or U36906 (N_36906,N_29360,N_23840);
and U36907 (N_36907,N_24339,N_28361);
nand U36908 (N_36908,N_27735,N_21222);
or U36909 (N_36909,N_22921,N_25234);
nand U36910 (N_36910,N_28639,N_23559);
or U36911 (N_36911,N_27681,N_26959);
nor U36912 (N_36912,N_26222,N_28474);
nor U36913 (N_36913,N_24418,N_23045);
nor U36914 (N_36914,N_23668,N_23718);
and U36915 (N_36915,N_28846,N_26688);
xor U36916 (N_36916,N_29303,N_29647);
and U36917 (N_36917,N_21466,N_26694);
nor U36918 (N_36918,N_26903,N_28111);
nand U36919 (N_36919,N_20829,N_25068);
or U36920 (N_36920,N_22929,N_28577);
nand U36921 (N_36921,N_26001,N_22753);
nor U36922 (N_36922,N_22198,N_21779);
nor U36923 (N_36923,N_22392,N_25311);
or U36924 (N_36924,N_23521,N_21940);
xor U36925 (N_36925,N_23536,N_28867);
nor U36926 (N_36926,N_20444,N_23427);
or U36927 (N_36927,N_20981,N_27916);
nand U36928 (N_36928,N_21725,N_20905);
xnor U36929 (N_36929,N_24418,N_22411);
nor U36930 (N_36930,N_28228,N_28877);
xor U36931 (N_36931,N_27155,N_23995);
or U36932 (N_36932,N_20675,N_24591);
and U36933 (N_36933,N_23839,N_20899);
nor U36934 (N_36934,N_21455,N_29444);
xnor U36935 (N_36935,N_25933,N_23489);
nor U36936 (N_36936,N_25929,N_21129);
or U36937 (N_36937,N_23976,N_23630);
nand U36938 (N_36938,N_26895,N_25287);
nor U36939 (N_36939,N_24028,N_29469);
or U36940 (N_36940,N_22613,N_27050);
nor U36941 (N_36941,N_22937,N_23572);
xnor U36942 (N_36942,N_22451,N_23656);
or U36943 (N_36943,N_24089,N_22832);
nand U36944 (N_36944,N_28874,N_24543);
and U36945 (N_36945,N_25769,N_20698);
or U36946 (N_36946,N_25984,N_21300);
xnor U36947 (N_36947,N_27687,N_22894);
xnor U36948 (N_36948,N_29206,N_24616);
nor U36949 (N_36949,N_22111,N_21380);
and U36950 (N_36950,N_29205,N_29429);
nand U36951 (N_36951,N_23634,N_26424);
nor U36952 (N_36952,N_28784,N_20441);
or U36953 (N_36953,N_25847,N_29055);
nor U36954 (N_36954,N_26016,N_21415);
nor U36955 (N_36955,N_21275,N_21110);
and U36956 (N_36956,N_23566,N_27115);
nor U36957 (N_36957,N_22821,N_24682);
or U36958 (N_36958,N_25018,N_21548);
nor U36959 (N_36959,N_27808,N_25556);
nand U36960 (N_36960,N_21706,N_21021);
nand U36961 (N_36961,N_29034,N_29190);
nor U36962 (N_36962,N_27537,N_24684);
or U36963 (N_36963,N_22993,N_23227);
or U36964 (N_36964,N_24775,N_24810);
nor U36965 (N_36965,N_22421,N_24181);
xor U36966 (N_36966,N_20429,N_28644);
nor U36967 (N_36967,N_20829,N_22077);
xor U36968 (N_36968,N_29769,N_22128);
nand U36969 (N_36969,N_29926,N_24404);
nand U36970 (N_36970,N_28146,N_25123);
nor U36971 (N_36971,N_22429,N_29433);
nand U36972 (N_36972,N_21863,N_25659);
xnor U36973 (N_36973,N_23403,N_25668);
xor U36974 (N_36974,N_29123,N_23353);
nand U36975 (N_36975,N_25645,N_29967);
and U36976 (N_36976,N_22881,N_20629);
and U36977 (N_36977,N_23829,N_23134);
or U36978 (N_36978,N_28248,N_25754);
xnor U36979 (N_36979,N_29261,N_25919);
nor U36980 (N_36980,N_23653,N_27562);
or U36981 (N_36981,N_29552,N_28324);
nand U36982 (N_36982,N_21116,N_23698);
and U36983 (N_36983,N_23539,N_26558);
nand U36984 (N_36984,N_22336,N_28399);
nor U36985 (N_36985,N_23386,N_24026);
nor U36986 (N_36986,N_26606,N_22338);
nor U36987 (N_36987,N_28264,N_29167);
or U36988 (N_36988,N_29618,N_29021);
and U36989 (N_36989,N_29563,N_24244);
nand U36990 (N_36990,N_23033,N_20239);
nor U36991 (N_36991,N_24443,N_28295);
nor U36992 (N_36992,N_26846,N_25968);
nand U36993 (N_36993,N_24581,N_20515);
or U36994 (N_36994,N_29425,N_25296);
nand U36995 (N_36995,N_29994,N_25526);
xor U36996 (N_36996,N_26972,N_27971);
or U36997 (N_36997,N_21630,N_25370);
xnor U36998 (N_36998,N_28942,N_25182);
nor U36999 (N_36999,N_20552,N_23573);
nor U37000 (N_37000,N_20267,N_23938);
xnor U37001 (N_37001,N_25983,N_25049);
or U37002 (N_37002,N_23919,N_25108);
and U37003 (N_37003,N_21941,N_26224);
or U37004 (N_37004,N_23065,N_20710);
and U37005 (N_37005,N_29478,N_22112);
or U37006 (N_37006,N_24954,N_28824);
xnor U37007 (N_37007,N_29106,N_22069);
xnor U37008 (N_37008,N_24215,N_24424);
and U37009 (N_37009,N_25968,N_27469);
and U37010 (N_37010,N_26733,N_29008);
nor U37011 (N_37011,N_24206,N_24696);
nor U37012 (N_37012,N_25787,N_26445);
nor U37013 (N_37013,N_24898,N_26574);
nor U37014 (N_37014,N_26004,N_20892);
xnor U37015 (N_37015,N_27055,N_22542);
or U37016 (N_37016,N_29962,N_23200);
nor U37017 (N_37017,N_26181,N_20474);
or U37018 (N_37018,N_24418,N_26197);
xnor U37019 (N_37019,N_20087,N_28506);
xnor U37020 (N_37020,N_21810,N_21417);
xnor U37021 (N_37021,N_23851,N_28050);
or U37022 (N_37022,N_26016,N_24022);
nor U37023 (N_37023,N_26435,N_26273);
nand U37024 (N_37024,N_27705,N_24466);
nand U37025 (N_37025,N_29906,N_25880);
or U37026 (N_37026,N_25810,N_26267);
or U37027 (N_37027,N_26376,N_21801);
and U37028 (N_37028,N_22188,N_27400);
or U37029 (N_37029,N_28134,N_25593);
or U37030 (N_37030,N_22160,N_26165);
nor U37031 (N_37031,N_28281,N_22433);
nand U37032 (N_37032,N_27406,N_21598);
xor U37033 (N_37033,N_21845,N_27580);
and U37034 (N_37034,N_26487,N_24087);
nand U37035 (N_37035,N_25576,N_26561);
and U37036 (N_37036,N_29586,N_28502);
and U37037 (N_37037,N_23180,N_28836);
nor U37038 (N_37038,N_21482,N_26213);
xor U37039 (N_37039,N_20541,N_22784);
and U37040 (N_37040,N_27503,N_22538);
xor U37041 (N_37041,N_22263,N_24823);
nand U37042 (N_37042,N_20316,N_26633);
xnor U37043 (N_37043,N_26709,N_25839);
and U37044 (N_37044,N_21098,N_26894);
nor U37045 (N_37045,N_22003,N_20367);
or U37046 (N_37046,N_25524,N_20661);
nor U37047 (N_37047,N_23169,N_22272);
and U37048 (N_37048,N_27234,N_24516);
xor U37049 (N_37049,N_28823,N_28968);
or U37050 (N_37050,N_22905,N_22684);
xor U37051 (N_37051,N_28550,N_28656);
nand U37052 (N_37052,N_27440,N_20085);
nor U37053 (N_37053,N_21738,N_27260);
nor U37054 (N_37054,N_20765,N_29706);
nor U37055 (N_37055,N_25452,N_25505);
xnor U37056 (N_37056,N_27648,N_27488);
nor U37057 (N_37057,N_26705,N_20047);
and U37058 (N_37058,N_28724,N_24604);
xnor U37059 (N_37059,N_21759,N_24660);
nor U37060 (N_37060,N_29877,N_25448);
xor U37061 (N_37061,N_20238,N_29716);
xnor U37062 (N_37062,N_24655,N_21748);
xnor U37063 (N_37063,N_27397,N_27361);
nor U37064 (N_37064,N_20281,N_24098);
or U37065 (N_37065,N_25609,N_26879);
nor U37066 (N_37066,N_29270,N_26282);
xor U37067 (N_37067,N_26480,N_29165);
xor U37068 (N_37068,N_29732,N_27466);
nor U37069 (N_37069,N_20898,N_28670);
xor U37070 (N_37070,N_28705,N_26903);
nand U37071 (N_37071,N_25993,N_28642);
and U37072 (N_37072,N_28532,N_29921);
xnor U37073 (N_37073,N_24429,N_25269);
nand U37074 (N_37074,N_26251,N_24670);
or U37075 (N_37075,N_27237,N_20219);
or U37076 (N_37076,N_29249,N_25394);
nor U37077 (N_37077,N_22382,N_28647);
nand U37078 (N_37078,N_22017,N_27224);
and U37079 (N_37079,N_22863,N_20173);
and U37080 (N_37080,N_22118,N_23329);
or U37081 (N_37081,N_26482,N_21716);
nand U37082 (N_37082,N_24792,N_27449);
nand U37083 (N_37083,N_20529,N_25831);
xnor U37084 (N_37084,N_22407,N_22442);
or U37085 (N_37085,N_25364,N_27414);
and U37086 (N_37086,N_28389,N_21588);
xor U37087 (N_37087,N_24468,N_20223);
and U37088 (N_37088,N_28762,N_20711);
and U37089 (N_37089,N_26198,N_20756);
xor U37090 (N_37090,N_23413,N_25368);
xnor U37091 (N_37091,N_27863,N_24258);
and U37092 (N_37092,N_20166,N_26972);
nor U37093 (N_37093,N_29936,N_22274);
nand U37094 (N_37094,N_21181,N_24933);
or U37095 (N_37095,N_27657,N_23876);
xnor U37096 (N_37096,N_23685,N_26500);
nand U37097 (N_37097,N_22972,N_26982);
nand U37098 (N_37098,N_29269,N_21231);
nand U37099 (N_37099,N_20298,N_20204);
xor U37100 (N_37100,N_22475,N_27257);
and U37101 (N_37101,N_26001,N_29487);
or U37102 (N_37102,N_21722,N_22162);
xnor U37103 (N_37103,N_21386,N_28811);
nand U37104 (N_37104,N_22997,N_20433);
nor U37105 (N_37105,N_27551,N_29624);
nor U37106 (N_37106,N_20349,N_26385);
or U37107 (N_37107,N_21696,N_27242);
or U37108 (N_37108,N_25354,N_24965);
or U37109 (N_37109,N_23767,N_24329);
xor U37110 (N_37110,N_27609,N_28798);
or U37111 (N_37111,N_21367,N_26539);
xnor U37112 (N_37112,N_27207,N_20073);
xnor U37113 (N_37113,N_22975,N_28515);
and U37114 (N_37114,N_28027,N_27977);
xnor U37115 (N_37115,N_27415,N_26771);
xor U37116 (N_37116,N_20799,N_26265);
or U37117 (N_37117,N_24408,N_29417);
nor U37118 (N_37118,N_23743,N_20719);
nor U37119 (N_37119,N_25891,N_23622);
nor U37120 (N_37120,N_25147,N_26515);
nor U37121 (N_37121,N_23013,N_22053);
xnor U37122 (N_37122,N_24068,N_29085);
nor U37123 (N_37123,N_23375,N_22635);
and U37124 (N_37124,N_23123,N_28470);
xnor U37125 (N_37125,N_22190,N_29192);
nand U37126 (N_37126,N_29606,N_28938);
xor U37127 (N_37127,N_28891,N_27414);
and U37128 (N_37128,N_24398,N_22228);
nand U37129 (N_37129,N_22952,N_21324);
or U37130 (N_37130,N_24179,N_25007);
nand U37131 (N_37131,N_27674,N_20011);
and U37132 (N_37132,N_24624,N_26442);
or U37133 (N_37133,N_25875,N_29431);
nand U37134 (N_37134,N_21179,N_25881);
nor U37135 (N_37135,N_27101,N_20362);
nor U37136 (N_37136,N_29339,N_24107);
or U37137 (N_37137,N_27056,N_23015);
and U37138 (N_37138,N_21610,N_27330);
or U37139 (N_37139,N_26769,N_21720);
nand U37140 (N_37140,N_29527,N_29606);
and U37141 (N_37141,N_25207,N_25980);
nor U37142 (N_37142,N_27850,N_25536);
nor U37143 (N_37143,N_26381,N_21690);
nand U37144 (N_37144,N_28876,N_21012);
xnor U37145 (N_37145,N_22293,N_21355);
and U37146 (N_37146,N_20592,N_23509);
nor U37147 (N_37147,N_22534,N_23732);
or U37148 (N_37148,N_28002,N_24649);
nor U37149 (N_37149,N_27123,N_26463);
xnor U37150 (N_37150,N_23748,N_29195);
and U37151 (N_37151,N_28160,N_28789);
or U37152 (N_37152,N_22462,N_29325);
or U37153 (N_37153,N_20235,N_22505);
nor U37154 (N_37154,N_22258,N_20587);
nand U37155 (N_37155,N_27720,N_23590);
nand U37156 (N_37156,N_28234,N_23052);
and U37157 (N_37157,N_27438,N_24610);
or U37158 (N_37158,N_27437,N_23481);
nor U37159 (N_37159,N_22032,N_21464);
xor U37160 (N_37160,N_23807,N_25811);
xnor U37161 (N_37161,N_29775,N_21174);
xnor U37162 (N_37162,N_20201,N_24565);
nand U37163 (N_37163,N_23198,N_21492);
nand U37164 (N_37164,N_21417,N_22567);
and U37165 (N_37165,N_21456,N_24849);
or U37166 (N_37166,N_27431,N_26162);
and U37167 (N_37167,N_29302,N_22017);
or U37168 (N_37168,N_21535,N_26736);
or U37169 (N_37169,N_24449,N_28776);
nand U37170 (N_37170,N_21700,N_21654);
nor U37171 (N_37171,N_22499,N_24053);
nand U37172 (N_37172,N_22034,N_26846);
xor U37173 (N_37173,N_28170,N_24387);
or U37174 (N_37174,N_29153,N_20059);
nor U37175 (N_37175,N_28158,N_23660);
and U37176 (N_37176,N_23160,N_23925);
nand U37177 (N_37177,N_23455,N_23210);
nor U37178 (N_37178,N_23167,N_27281);
and U37179 (N_37179,N_27519,N_27486);
nor U37180 (N_37180,N_28732,N_23750);
or U37181 (N_37181,N_25118,N_24368);
nand U37182 (N_37182,N_25804,N_23416);
xor U37183 (N_37183,N_20088,N_25696);
or U37184 (N_37184,N_21773,N_21898);
nor U37185 (N_37185,N_29200,N_24356);
or U37186 (N_37186,N_26277,N_24703);
xor U37187 (N_37187,N_28332,N_27860);
xnor U37188 (N_37188,N_29156,N_25376);
nor U37189 (N_37189,N_23137,N_25718);
nor U37190 (N_37190,N_23830,N_20926);
nor U37191 (N_37191,N_20569,N_22777);
xor U37192 (N_37192,N_24884,N_20623);
or U37193 (N_37193,N_28352,N_26910);
and U37194 (N_37194,N_27742,N_28214);
nand U37195 (N_37195,N_24780,N_27834);
and U37196 (N_37196,N_24113,N_24360);
nand U37197 (N_37197,N_27515,N_27273);
or U37198 (N_37198,N_29575,N_26091);
nor U37199 (N_37199,N_25008,N_28545);
xnor U37200 (N_37200,N_22462,N_29767);
or U37201 (N_37201,N_28839,N_25966);
nor U37202 (N_37202,N_28629,N_20856);
and U37203 (N_37203,N_28305,N_27215);
nand U37204 (N_37204,N_27822,N_28277);
nor U37205 (N_37205,N_26860,N_28404);
xor U37206 (N_37206,N_23276,N_27055);
xor U37207 (N_37207,N_22716,N_27810);
nor U37208 (N_37208,N_21334,N_26016);
nand U37209 (N_37209,N_25332,N_27945);
nand U37210 (N_37210,N_29126,N_29985);
nand U37211 (N_37211,N_22087,N_24303);
nand U37212 (N_37212,N_29858,N_26106);
nand U37213 (N_37213,N_24160,N_26958);
and U37214 (N_37214,N_23871,N_22092);
xor U37215 (N_37215,N_27703,N_21631);
nand U37216 (N_37216,N_25780,N_20574);
nor U37217 (N_37217,N_22098,N_24362);
or U37218 (N_37218,N_22792,N_20302);
or U37219 (N_37219,N_28991,N_23830);
nor U37220 (N_37220,N_22625,N_22969);
or U37221 (N_37221,N_27451,N_26555);
nor U37222 (N_37222,N_26176,N_20281);
nand U37223 (N_37223,N_20652,N_26979);
or U37224 (N_37224,N_26660,N_28740);
nand U37225 (N_37225,N_22402,N_23852);
nor U37226 (N_37226,N_25851,N_20283);
and U37227 (N_37227,N_26822,N_22488);
nand U37228 (N_37228,N_28746,N_29850);
xor U37229 (N_37229,N_29501,N_20603);
nand U37230 (N_37230,N_26853,N_27669);
nor U37231 (N_37231,N_28367,N_28118);
nor U37232 (N_37232,N_26228,N_28737);
and U37233 (N_37233,N_23119,N_21626);
nor U37234 (N_37234,N_20155,N_26858);
nor U37235 (N_37235,N_24470,N_27980);
or U37236 (N_37236,N_27851,N_28582);
xor U37237 (N_37237,N_23386,N_21717);
nor U37238 (N_37238,N_20595,N_29513);
or U37239 (N_37239,N_25259,N_20465);
or U37240 (N_37240,N_22911,N_24917);
and U37241 (N_37241,N_23517,N_29967);
or U37242 (N_37242,N_26595,N_22767);
nand U37243 (N_37243,N_22480,N_27680);
xnor U37244 (N_37244,N_25863,N_23429);
and U37245 (N_37245,N_27711,N_26478);
xnor U37246 (N_37246,N_28396,N_22294);
nor U37247 (N_37247,N_27743,N_21166);
or U37248 (N_37248,N_29004,N_29016);
or U37249 (N_37249,N_21680,N_20544);
nor U37250 (N_37250,N_21115,N_21360);
or U37251 (N_37251,N_21174,N_27435);
and U37252 (N_37252,N_21476,N_29752);
nand U37253 (N_37253,N_20721,N_25607);
xnor U37254 (N_37254,N_22730,N_25030);
xor U37255 (N_37255,N_22856,N_25390);
and U37256 (N_37256,N_23609,N_29617);
nand U37257 (N_37257,N_26045,N_23633);
and U37258 (N_37258,N_27312,N_28149);
nand U37259 (N_37259,N_26468,N_22501);
or U37260 (N_37260,N_26550,N_29073);
nand U37261 (N_37261,N_21811,N_25400);
and U37262 (N_37262,N_22246,N_25829);
nor U37263 (N_37263,N_21649,N_22568);
nand U37264 (N_37264,N_25954,N_24275);
xor U37265 (N_37265,N_29121,N_24481);
nor U37266 (N_37266,N_26657,N_24898);
or U37267 (N_37267,N_27444,N_24183);
nor U37268 (N_37268,N_26092,N_22981);
nor U37269 (N_37269,N_24964,N_21355);
or U37270 (N_37270,N_21974,N_26733);
and U37271 (N_37271,N_25360,N_28257);
nor U37272 (N_37272,N_20522,N_23846);
xnor U37273 (N_37273,N_21534,N_22592);
or U37274 (N_37274,N_26666,N_29738);
nor U37275 (N_37275,N_28674,N_24398);
nand U37276 (N_37276,N_27829,N_24890);
or U37277 (N_37277,N_29658,N_24440);
nand U37278 (N_37278,N_26133,N_25624);
or U37279 (N_37279,N_24730,N_21672);
or U37280 (N_37280,N_23582,N_27789);
and U37281 (N_37281,N_27181,N_20855);
nor U37282 (N_37282,N_28050,N_24529);
nand U37283 (N_37283,N_24552,N_27236);
xnor U37284 (N_37284,N_26737,N_25449);
or U37285 (N_37285,N_22530,N_22100);
xor U37286 (N_37286,N_23061,N_23321);
and U37287 (N_37287,N_27323,N_22780);
and U37288 (N_37288,N_23447,N_22249);
or U37289 (N_37289,N_24556,N_23617);
and U37290 (N_37290,N_28959,N_25426);
xnor U37291 (N_37291,N_27438,N_29092);
or U37292 (N_37292,N_22475,N_27337);
nor U37293 (N_37293,N_28687,N_25833);
nor U37294 (N_37294,N_23833,N_27622);
nand U37295 (N_37295,N_29680,N_26265);
nor U37296 (N_37296,N_29931,N_24231);
nor U37297 (N_37297,N_29144,N_27603);
nor U37298 (N_37298,N_23665,N_28933);
and U37299 (N_37299,N_24134,N_28713);
and U37300 (N_37300,N_27754,N_20821);
xor U37301 (N_37301,N_29821,N_23802);
nand U37302 (N_37302,N_27507,N_26328);
nand U37303 (N_37303,N_27652,N_25861);
or U37304 (N_37304,N_25222,N_22448);
nand U37305 (N_37305,N_29609,N_22255);
and U37306 (N_37306,N_21604,N_24246);
xnor U37307 (N_37307,N_28021,N_23454);
nor U37308 (N_37308,N_20270,N_23236);
nor U37309 (N_37309,N_25864,N_27484);
xor U37310 (N_37310,N_25378,N_27875);
nor U37311 (N_37311,N_24359,N_28563);
and U37312 (N_37312,N_27533,N_22748);
and U37313 (N_37313,N_22780,N_24919);
xor U37314 (N_37314,N_24155,N_24694);
nor U37315 (N_37315,N_21275,N_22044);
xnor U37316 (N_37316,N_24826,N_26654);
xor U37317 (N_37317,N_25368,N_22725);
nand U37318 (N_37318,N_26371,N_20064);
xnor U37319 (N_37319,N_23945,N_29748);
xor U37320 (N_37320,N_23223,N_23583);
nand U37321 (N_37321,N_26251,N_25931);
and U37322 (N_37322,N_27884,N_28791);
nor U37323 (N_37323,N_21150,N_29293);
xor U37324 (N_37324,N_27244,N_24532);
or U37325 (N_37325,N_25560,N_20448);
xor U37326 (N_37326,N_26166,N_21244);
xor U37327 (N_37327,N_28813,N_20773);
nand U37328 (N_37328,N_20431,N_20397);
and U37329 (N_37329,N_23202,N_27604);
and U37330 (N_37330,N_25021,N_21374);
and U37331 (N_37331,N_21085,N_27986);
nor U37332 (N_37332,N_24812,N_22118);
nand U37333 (N_37333,N_21339,N_23904);
nor U37334 (N_37334,N_25521,N_29144);
xnor U37335 (N_37335,N_26977,N_25478);
nor U37336 (N_37336,N_29793,N_20699);
or U37337 (N_37337,N_25772,N_21569);
or U37338 (N_37338,N_25049,N_22389);
or U37339 (N_37339,N_29770,N_26545);
or U37340 (N_37340,N_28028,N_26297);
nor U37341 (N_37341,N_20444,N_24862);
or U37342 (N_37342,N_27641,N_25725);
xnor U37343 (N_37343,N_25912,N_21273);
or U37344 (N_37344,N_28193,N_27313);
or U37345 (N_37345,N_26702,N_29746);
or U37346 (N_37346,N_27367,N_23601);
and U37347 (N_37347,N_20388,N_27216);
xnor U37348 (N_37348,N_21396,N_26318);
nor U37349 (N_37349,N_20030,N_22169);
and U37350 (N_37350,N_23892,N_25195);
nor U37351 (N_37351,N_29983,N_24177);
and U37352 (N_37352,N_20626,N_25111);
and U37353 (N_37353,N_21372,N_28648);
nor U37354 (N_37354,N_22459,N_21789);
nand U37355 (N_37355,N_28260,N_20040);
nor U37356 (N_37356,N_23952,N_25661);
or U37357 (N_37357,N_26519,N_26907);
or U37358 (N_37358,N_24885,N_20009);
or U37359 (N_37359,N_29115,N_24783);
or U37360 (N_37360,N_22557,N_20157);
nand U37361 (N_37361,N_21947,N_20534);
nand U37362 (N_37362,N_26410,N_21657);
and U37363 (N_37363,N_23796,N_28322);
nand U37364 (N_37364,N_20548,N_20060);
nor U37365 (N_37365,N_29680,N_21250);
xor U37366 (N_37366,N_27352,N_28181);
nor U37367 (N_37367,N_22717,N_27570);
xor U37368 (N_37368,N_27414,N_25852);
or U37369 (N_37369,N_24195,N_23334);
and U37370 (N_37370,N_23123,N_21393);
xor U37371 (N_37371,N_28611,N_25682);
nand U37372 (N_37372,N_29902,N_21700);
and U37373 (N_37373,N_28254,N_28040);
xnor U37374 (N_37374,N_23486,N_26311);
or U37375 (N_37375,N_24969,N_28741);
nand U37376 (N_37376,N_20240,N_27347);
nor U37377 (N_37377,N_26924,N_22343);
and U37378 (N_37378,N_26911,N_23627);
nor U37379 (N_37379,N_27041,N_28823);
xor U37380 (N_37380,N_28965,N_27559);
or U37381 (N_37381,N_29635,N_20669);
or U37382 (N_37382,N_20935,N_23266);
nand U37383 (N_37383,N_23526,N_21853);
or U37384 (N_37384,N_20650,N_23299);
xnor U37385 (N_37385,N_26461,N_28719);
or U37386 (N_37386,N_23277,N_22806);
nand U37387 (N_37387,N_23624,N_24148);
and U37388 (N_37388,N_24731,N_29116);
nor U37389 (N_37389,N_21108,N_29233);
and U37390 (N_37390,N_27559,N_29760);
or U37391 (N_37391,N_23480,N_28960);
nor U37392 (N_37392,N_26791,N_29433);
nor U37393 (N_37393,N_28613,N_23241);
or U37394 (N_37394,N_24982,N_22974);
nor U37395 (N_37395,N_25680,N_26464);
and U37396 (N_37396,N_28892,N_25393);
nand U37397 (N_37397,N_26583,N_29305);
or U37398 (N_37398,N_20068,N_22636);
and U37399 (N_37399,N_22309,N_24604);
or U37400 (N_37400,N_27790,N_21372);
or U37401 (N_37401,N_28011,N_28126);
xnor U37402 (N_37402,N_21677,N_29589);
nor U37403 (N_37403,N_23716,N_29657);
and U37404 (N_37404,N_20981,N_23789);
or U37405 (N_37405,N_26057,N_20327);
or U37406 (N_37406,N_29204,N_25576);
nor U37407 (N_37407,N_25669,N_29227);
nand U37408 (N_37408,N_24707,N_22985);
or U37409 (N_37409,N_25512,N_22338);
nor U37410 (N_37410,N_26697,N_26233);
xnor U37411 (N_37411,N_20791,N_26537);
xor U37412 (N_37412,N_26505,N_26519);
xor U37413 (N_37413,N_26242,N_27644);
nor U37414 (N_37414,N_29416,N_24076);
and U37415 (N_37415,N_23060,N_22693);
nand U37416 (N_37416,N_26732,N_24653);
nor U37417 (N_37417,N_21313,N_28496);
or U37418 (N_37418,N_21786,N_23868);
nor U37419 (N_37419,N_26913,N_24828);
xnor U37420 (N_37420,N_28447,N_26331);
or U37421 (N_37421,N_22374,N_23533);
nand U37422 (N_37422,N_25831,N_21193);
or U37423 (N_37423,N_24171,N_24036);
and U37424 (N_37424,N_21063,N_29406);
nor U37425 (N_37425,N_25680,N_23618);
nor U37426 (N_37426,N_29068,N_27224);
xnor U37427 (N_37427,N_23493,N_21550);
nand U37428 (N_37428,N_23976,N_20136);
nand U37429 (N_37429,N_24793,N_21517);
or U37430 (N_37430,N_24020,N_28166);
xor U37431 (N_37431,N_22977,N_28211);
xor U37432 (N_37432,N_28067,N_28747);
or U37433 (N_37433,N_28548,N_27482);
and U37434 (N_37434,N_28328,N_21406);
xor U37435 (N_37435,N_27533,N_28864);
nand U37436 (N_37436,N_27116,N_23865);
and U37437 (N_37437,N_26252,N_28431);
and U37438 (N_37438,N_29101,N_20814);
and U37439 (N_37439,N_22177,N_28369);
and U37440 (N_37440,N_23904,N_28094);
and U37441 (N_37441,N_24040,N_27531);
xor U37442 (N_37442,N_21926,N_24534);
xor U37443 (N_37443,N_23572,N_20854);
or U37444 (N_37444,N_27648,N_27979);
or U37445 (N_37445,N_23501,N_27219);
or U37446 (N_37446,N_27597,N_20601);
nand U37447 (N_37447,N_28740,N_26389);
nand U37448 (N_37448,N_23028,N_29364);
xor U37449 (N_37449,N_21328,N_21433);
or U37450 (N_37450,N_23677,N_24593);
or U37451 (N_37451,N_22937,N_25682);
nor U37452 (N_37452,N_25355,N_21280);
nor U37453 (N_37453,N_29089,N_21912);
nor U37454 (N_37454,N_29273,N_25586);
or U37455 (N_37455,N_26951,N_29286);
or U37456 (N_37456,N_24603,N_20457);
or U37457 (N_37457,N_20452,N_29909);
xor U37458 (N_37458,N_22273,N_20535);
xnor U37459 (N_37459,N_23197,N_28331);
nor U37460 (N_37460,N_27471,N_20134);
or U37461 (N_37461,N_29233,N_20192);
or U37462 (N_37462,N_25614,N_23990);
and U37463 (N_37463,N_22771,N_27475);
nor U37464 (N_37464,N_20547,N_22283);
nor U37465 (N_37465,N_26669,N_25524);
nand U37466 (N_37466,N_26071,N_24870);
or U37467 (N_37467,N_25648,N_23751);
nand U37468 (N_37468,N_23125,N_23751);
or U37469 (N_37469,N_26675,N_22394);
or U37470 (N_37470,N_21077,N_25915);
xor U37471 (N_37471,N_21250,N_26468);
xor U37472 (N_37472,N_24169,N_22073);
xnor U37473 (N_37473,N_22096,N_26826);
and U37474 (N_37474,N_26831,N_26941);
xor U37475 (N_37475,N_20145,N_23781);
or U37476 (N_37476,N_21332,N_22321);
xor U37477 (N_37477,N_23846,N_21954);
nand U37478 (N_37478,N_22769,N_23901);
xor U37479 (N_37479,N_27109,N_29878);
nor U37480 (N_37480,N_26210,N_28854);
and U37481 (N_37481,N_27614,N_23219);
xnor U37482 (N_37482,N_27870,N_25326);
xnor U37483 (N_37483,N_20787,N_20342);
or U37484 (N_37484,N_24287,N_21960);
nand U37485 (N_37485,N_27240,N_25848);
nor U37486 (N_37486,N_29001,N_23987);
nand U37487 (N_37487,N_20680,N_29173);
or U37488 (N_37488,N_29679,N_29911);
or U37489 (N_37489,N_28407,N_21229);
nor U37490 (N_37490,N_20156,N_26170);
or U37491 (N_37491,N_20391,N_20920);
nor U37492 (N_37492,N_21887,N_29793);
nand U37493 (N_37493,N_21772,N_26248);
xnor U37494 (N_37494,N_25787,N_20246);
and U37495 (N_37495,N_21708,N_28256);
or U37496 (N_37496,N_26400,N_20545);
nor U37497 (N_37497,N_29017,N_20967);
nor U37498 (N_37498,N_20240,N_23011);
and U37499 (N_37499,N_21978,N_29137);
nor U37500 (N_37500,N_27778,N_24377);
and U37501 (N_37501,N_24050,N_21945);
xor U37502 (N_37502,N_29357,N_27472);
xor U37503 (N_37503,N_22173,N_28202);
xnor U37504 (N_37504,N_26761,N_24020);
and U37505 (N_37505,N_28240,N_21829);
nand U37506 (N_37506,N_25534,N_22017);
nor U37507 (N_37507,N_27606,N_20574);
xnor U37508 (N_37508,N_27178,N_25871);
nand U37509 (N_37509,N_21984,N_28034);
nor U37510 (N_37510,N_20136,N_27866);
nor U37511 (N_37511,N_25593,N_22899);
nor U37512 (N_37512,N_26416,N_24574);
xor U37513 (N_37513,N_29729,N_27391);
nor U37514 (N_37514,N_22426,N_25192);
nor U37515 (N_37515,N_27586,N_22387);
or U37516 (N_37516,N_21815,N_25451);
and U37517 (N_37517,N_29490,N_23862);
and U37518 (N_37518,N_25853,N_26064);
nand U37519 (N_37519,N_26085,N_25497);
nor U37520 (N_37520,N_25145,N_26323);
or U37521 (N_37521,N_25259,N_26712);
or U37522 (N_37522,N_23907,N_20947);
nor U37523 (N_37523,N_22048,N_21846);
and U37524 (N_37524,N_20871,N_20134);
or U37525 (N_37525,N_20598,N_22403);
nand U37526 (N_37526,N_27188,N_29845);
and U37527 (N_37527,N_24517,N_24961);
or U37528 (N_37528,N_28341,N_27271);
nor U37529 (N_37529,N_26844,N_21742);
and U37530 (N_37530,N_20344,N_29286);
nand U37531 (N_37531,N_20807,N_23316);
nor U37532 (N_37532,N_26674,N_25493);
nor U37533 (N_37533,N_23425,N_21084);
and U37534 (N_37534,N_25271,N_21536);
nor U37535 (N_37535,N_20842,N_29563);
nand U37536 (N_37536,N_23238,N_22410);
or U37537 (N_37537,N_25914,N_24945);
xor U37538 (N_37538,N_25776,N_28397);
nor U37539 (N_37539,N_25604,N_28958);
xor U37540 (N_37540,N_22079,N_22821);
nand U37541 (N_37541,N_25634,N_20124);
nand U37542 (N_37542,N_23527,N_24251);
xor U37543 (N_37543,N_21740,N_27883);
xor U37544 (N_37544,N_26069,N_25275);
nor U37545 (N_37545,N_28355,N_29051);
nand U37546 (N_37546,N_29890,N_28512);
and U37547 (N_37547,N_20136,N_20857);
or U37548 (N_37548,N_24009,N_20834);
or U37549 (N_37549,N_25027,N_25207);
nand U37550 (N_37550,N_21859,N_28946);
xor U37551 (N_37551,N_26877,N_28173);
xnor U37552 (N_37552,N_27764,N_27261);
or U37553 (N_37553,N_26422,N_27200);
nand U37554 (N_37554,N_25685,N_22219);
or U37555 (N_37555,N_22302,N_25692);
or U37556 (N_37556,N_23730,N_28980);
or U37557 (N_37557,N_27997,N_28690);
nand U37558 (N_37558,N_20854,N_28822);
nor U37559 (N_37559,N_20370,N_29980);
xnor U37560 (N_37560,N_26111,N_23050);
or U37561 (N_37561,N_27847,N_27133);
nor U37562 (N_37562,N_24897,N_20283);
nand U37563 (N_37563,N_22352,N_27933);
and U37564 (N_37564,N_22808,N_29423);
nand U37565 (N_37565,N_25547,N_20846);
and U37566 (N_37566,N_24833,N_23254);
xnor U37567 (N_37567,N_29816,N_23933);
or U37568 (N_37568,N_21024,N_20976);
or U37569 (N_37569,N_28771,N_25713);
or U37570 (N_37570,N_22303,N_20213);
and U37571 (N_37571,N_29720,N_21384);
nor U37572 (N_37572,N_23358,N_28626);
nand U37573 (N_37573,N_26201,N_28912);
nor U37574 (N_37574,N_26715,N_20477);
xnor U37575 (N_37575,N_22499,N_27869);
nand U37576 (N_37576,N_21405,N_27287);
xor U37577 (N_37577,N_25840,N_26276);
xor U37578 (N_37578,N_21128,N_28806);
nor U37579 (N_37579,N_24551,N_27316);
xor U37580 (N_37580,N_29547,N_22844);
nand U37581 (N_37581,N_29403,N_21523);
nor U37582 (N_37582,N_26272,N_29340);
and U37583 (N_37583,N_25561,N_28984);
and U37584 (N_37584,N_29024,N_25307);
or U37585 (N_37585,N_21035,N_28166);
nor U37586 (N_37586,N_25550,N_23145);
nor U37587 (N_37587,N_27028,N_24821);
or U37588 (N_37588,N_25117,N_27352);
xor U37589 (N_37589,N_22974,N_20451);
xor U37590 (N_37590,N_26663,N_27820);
nand U37591 (N_37591,N_22824,N_28021);
or U37592 (N_37592,N_28490,N_21047);
nand U37593 (N_37593,N_23722,N_26567);
xnor U37594 (N_37594,N_22490,N_28195);
or U37595 (N_37595,N_23551,N_20217);
and U37596 (N_37596,N_28674,N_24660);
nand U37597 (N_37597,N_28907,N_20007);
and U37598 (N_37598,N_26432,N_28532);
xnor U37599 (N_37599,N_22019,N_26045);
or U37600 (N_37600,N_25270,N_21592);
and U37601 (N_37601,N_28389,N_25007);
nor U37602 (N_37602,N_26121,N_22386);
nor U37603 (N_37603,N_25401,N_20575);
nand U37604 (N_37604,N_29411,N_25891);
and U37605 (N_37605,N_28295,N_20119);
or U37606 (N_37606,N_29497,N_23495);
or U37607 (N_37607,N_25780,N_27702);
and U37608 (N_37608,N_28396,N_23275);
or U37609 (N_37609,N_27105,N_24797);
nor U37610 (N_37610,N_21636,N_26088);
or U37611 (N_37611,N_25061,N_20322);
nor U37612 (N_37612,N_20604,N_27375);
nor U37613 (N_37613,N_28695,N_21691);
and U37614 (N_37614,N_25341,N_25613);
xnor U37615 (N_37615,N_24385,N_25174);
and U37616 (N_37616,N_26835,N_29157);
nand U37617 (N_37617,N_25929,N_28722);
nor U37618 (N_37618,N_25067,N_25397);
or U37619 (N_37619,N_29487,N_23129);
or U37620 (N_37620,N_21239,N_27287);
xnor U37621 (N_37621,N_24854,N_28085);
xor U37622 (N_37622,N_20975,N_25405);
nor U37623 (N_37623,N_27364,N_28215);
nand U37624 (N_37624,N_26317,N_26392);
xor U37625 (N_37625,N_24672,N_21907);
nor U37626 (N_37626,N_29138,N_28392);
and U37627 (N_37627,N_27659,N_22718);
nand U37628 (N_37628,N_28624,N_22185);
or U37629 (N_37629,N_27541,N_29200);
nor U37630 (N_37630,N_25211,N_26383);
and U37631 (N_37631,N_28576,N_24347);
xor U37632 (N_37632,N_23839,N_25039);
or U37633 (N_37633,N_28084,N_25557);
nand U37634 (N_37634,N_29893,N_23766);
nand U37635 (N_37635,N_20401,N_24606);
nand U37636 (N_37636,N_21035,N_28004);
or U37637 (N_37637,N_26594,N_26280);
xnor U37638 (N_37638,N_28924,N_20440);
nor U37639 (N_37639,N_22414,N_28298);
or U37640 (N_37640,N_27089,N_20040);
nor U37641 (N_37641,N_24971,N_27510);
nor U37642 (N_37642,N_22426,N_28961);
nor U37643 (N_37643,N_24080,N_21312);
nor U37644 (N_37644,N_29642,N_24501);
nor U37645 (N_37645,N_27629,N_28630);
xnor U37646 (N_37646,N_27325,N_25884);
nand U37647 (N_37647,N_29641,N_21038);
xor U37648 (N_37648,N_21169,N_21147);
and U37649 (N_37649,N_20084,N_21019);
nand U37650 (N_37650,N_28584,N_23595);
nor U37651 (N_37651,N_26569,N_28844);
and U37652 (N_37652,N_26539,N_20211);
xnor U37653 (N_37653,N_24345,N_23811);
or U37654 (N_37654,N_26210,N_23964);
nor U37655 (N_37655,N_29236,N_24257);
and U37656 (N_37656,N_23421,N_25453);
and U37657 (N_37657,N_25828,N_28686);
nor U37658 (N_37658,N_23209,N_21335);
nor U37659 (N_37659,N_26043,N_24384);
nor U37660 (N_37660,N_22195,N_23803);
or U37661 (N_37661,N_21457,N_23595);
and U37662 (N_37662,N_28919,N_26118);
and U37663 (N_37663,N_21381,N_28557);
xnor U37664 (N_37664,N_23995,N_24183);
xor U37665 (N_37665,N_27167,N_24221);
or U37666 (N_37666,N_24034,N_26218);
nand U37667 (N_37667,N_21373,N_20943);
or U37668 (N_37668,N_22642,N_25617);
nor U37669 (N_37669,N_29291,N_27204);
xor U37670 (N_37670,N_21279,N_21482);
xnor U37671 (N_37671,N_27577,N_24557);
and U37672 (N_37672,N_25296,N_28022);
xnor U37673 (N_37673,N_22317,N_26901);
xnor U37674 (N_37674,N_24573,N_28268);
xor U37675 (N_37675,N_28963,N_26085);
and U37676 (N_37676,N_20574,N_20981);
and U37677 (N_37677,N_26385,N_29986);
nor U37678 (N_37678,N_22544,N_21546);
nor U37679 (N_37679,N_27283,N_26167);
or U37680 (N_37680,N_20256,N_26849);
nor U37681 (N_37681,N_22679,N_27211);
nand U37682 (N_37682,N_23549,N_24164);
or U37683 (N_37683,N_29916,N_20628);
xnor U37684 (N_37684,N_22996,N_22488);
nor U37685 (N_37685,N_23493,N_20346);
nor U37686 (N_37686,N_22837,N_29064);
and U37687 (N_37687,N_29143,N_22792);
and U37688 (N_37688,N_24558,N_24909);
xor U37689 (N_37689,N_27306,N_28409);
xnor U37690 (N_37690,N_25443,N_26447);
and U37691 (N_37691,N_21656,N_23044);
and U37692 (N_37692,N_20144,N_20090);
nor U37693 (N_37693,N_24913,N_21286);
xnor U37694 (N_37694,N_22992,N_26950);
xor U37695 (N_37695,N_26662,N_22757);
or U37696 (N_37696,N_26037,N_23190);
nor U37697 (N_37697,N_27568,N_26274);
or U37698 (N_37698,N_26230,N_25266);
xor U37699 (N_37699,N_27032,N_21301);
nand U37700 (N_37700,N_27054,N_21210);
xnor U37701 (N_37701,N_28757,N_29773);
and U37702 (N_37702,N_29131,N_28614);
nor U37703 (N_37703,N_20167,N_25406);
xor U37704 (N_37704,N_27349,N_26464);
xor U37705 (N_37705,N_26682,N_25616);
xnor U37706 (N_37706,N_26465,N_24333);
nor U37707 (N_37707,N_23787,N_28932);
nor U37708 (N_37708,N_27028,N_26869);
xor U37709 (N_37709,N_28160,N_24010);
and U37710 (N_37710,N_29339,N_22162);
or U37711 (N_37711,N_20107,N_26858);
nand U37712 (N_37712,N_29232,N_20436);
and U37713 (N_37713,N_23161,N_21647);
nand U37714 (N_37714,N_21859,N_23529);
xnor U37715 (N_37715,N_26256,N_28400);
xnor U37716 (N_37716,N_29398,N_23652);
or U37717 (N_37717,N_20817,N_29115);
xnor U37718 (N_37718,N_23550,N_28121);
xor U37719 (N_37719,N_26841,N_29147);
and U37720 (N_37720,N_20723,N_21357);
or U37721 (N_37721,N_25501,N_20767);
or U37722 (N_37722,N_25809,N_25604);
and U37723 (N_37723,N_28395,N_23532);
or U37724 (N_37724,N_27334,N_24687);
nor U37725 (N_37725,N_24124,N_23697);
nor U37726 (N_37726,N_23287,N_24455);
nand U37727 (N_37727,N_26011,N_24914);
nor U37728 (N_37728,N_23314,N_20214);
and U37729 (N_37729,N_22199,N_24918);
or U37730 (N_37730,N_28224,N_28013);
or U37731 (N_37731,N_27895,N_22761);
xor U37732 (N_37732,N_24930,N_28894);
xnor U37733 (N_37733,N_28226,N_22815);
xor U37734 (N_37734,N_29544,N_22756);
xnor U37735 (N_37735,N_20957,N_20005);
nor U37736 (N_37736,N_25812,N_25795);
or U37737 (N_37737,N_22997,N_26489);
and U37738 (N_37738,N_25028,N_21085);
nor U37739 (N_37739,N_24673,N_24127);
and U37740 (N_37740,N_24142,N_21131);
or U37741 (N_37741,N_26238,N_22372);
xnor U37742 (N_37742,N_29722,N_27714);
xor U37743 (N_37743,N_20401,N_26083);
xnor U37744 (N_37744,N_27633,N_27486);
xor U37745 (N_37745,N_24440,N_26706);
xnor U37746 (N_37746,N_22669,N_28785);
nor U37747 (N_37747,N_22726,N_22922);
nor U37748 (N_37748,N_20236,N_21427);
xnor U37749 (N_37749,N_28256,N_28572);
and U37750 (N_37750,N_21806,N_23572);
and U37751 (N_37751,N_28661,N_25724);
and U37752 (N_37752,N_20252,N_24005);
or U37753 (N_37753,N_29346,N_23960);
nand U37754 (N_37754,N_25195,N_22175);
nor U37755 (N_37755,N_23784,N_28559);
nand U37756 (N_37756,N_27260,N_24659);
nor U37757 (N_37757,N_22463,N_20022);
and U37758 (N_37758,N_22432,N_29558);
and U37759 (N_37759,N_28842,N_21726);
nor U37760 (N_37760,N_29303,N_23445);
nor U37761 (N_37761,N_20552,N_27463);
or U37762 (N_37762,N_20884,N_27793);
nor U37763 (N_37763,N_22760,N_27198);
xnor U37764 (N_37764,N_27366,N_29571);
or U37765 (N_37765,N_23977,N_25746);
or U37766 (N_37766,N_25545,N_20774);
and U37767 (N_37767,N_25535,N_28128);
xor U37768 (N_37768,N_21975,N_28156);
nor U37769 (N_37769,N_25821,N_20847);
nor U37770 (N_37770,N_28001,N_27620);
or U37771 (N_37771,N_24802,N_25596);
or U37772 (N_37772,N_24426,N_23241);
and U37773 (N_37773,N_25421,N_26461);
xnor U37774 (N_37774,N_23050,N_27106);
nand U37775 (N_37775,N_26433,N_21812);
and U37776 (N_37776,N_22727,N_28955);
xor U37777 (N_37777,N_21062,N_28557);
nand U37778 (N_37778,N_23885,N_25962);
and U37779 (N_37779,N_24824,N_20207);
nor U37780 (N_37780,N_29820,N_25524);
xnor U37781 (N_37781,N_24123,N_25500);
nor U37782 (N_37782,N_22901,N_21937);
xnor U37783 (N_37783,N_20204,N_26385);
nand U37784 (N_37784,N_21534,N_22037);
nor U37785 (N_37785,N_25509,N_27983);
nor U37786 (N_37786,N_28351,N_22643);
or U37787 (N_37787,N_20718,N_26135);
nor U37788 (N_37788,N_23914,N_26373);
nand U37789 (N_37789,N_29265,N_25088);
nand U37790 (N_37790,N_22288,N_20394);
or U37791 (N_37791,N_21063,N_25195);
or U37792 (N_37792,N_23828,N_29915);
and U37793 (N_37793,N_27161,N_26672);
nand U37794 (N_37794,N_27789,N_23116);
nor U37795 (N_37795,N_26895,N_24540);
xnor U37796 (N_37796,N_23276,N_26236);
nand U37797 (N_37797,N_20795,N_21611);
xnor U37798 (N_37798,N_28574,N_23808);
and U37799 (N_37799,N_22983,N_27710);
or U37800 (N_37800,N_20527,N_22244);
xnor U37801 (N_37801,N_23890,N_28058);
nor U37802 (N_37802,N_23129,N_29370);
nor U37803 (N_37803,N_25458,N_20788);
or U37804 (N_37804,N_28090,N_20491);
nor U37805 (N_37805,N_24684,N_22482);
and U37806 (N_37806,N_20527,N_22794);
xor U37807 (N_37807,N_27590,N_22267);
nand U37808 (N_37808,N_28865,N_29599);
xor U37809 (N_37809,N_25600,N_26931);
or U37810 (N_37810,N_24990,N_20232);
nor U37811 (N_37811,N_25136,N_20901);
nor U37812 (N_37812,N_28306,N_20091);
xor U37813 (N_37813,N_28699,N_22829);
xor U37814 (N_37814,N_29820,N_20726);
xor U37815 (N_37815,N_25934,N_21340);
and U37816 (N_37816,N_27192,N_23505);
and U37817 (N_37817,N_27331,N_25987);
nand U37818 (N_37818,N_28214,N_25108);
or U37819 (N_37819,N_28707,N_21486);
xnor U37820 (N_37820,N_27291,N_28960);
xor U37821 (N_37821,N_27499,N_29788);
nor U37822 (N_37822,N_22861,N_22608);
nor U37823 (N_37823,N_29634,N_27112);
xor U37824 (N_37824,N_28719,N_23159);
or U37825 (N_37825,N_28028,N_26587);
nand U37826 (N_37826,N_25552,N_25943);
nor U37827 (N_37827,N_28819,N_25586);
xnor U37828 (N_37828,N_20879,N_21956);
xnor U37829 (N_37829,N_23712,N_23918);
and U37830 (N_37830,N_28120,N_25384);
or U37831 (N_37831,N_28450,N_24579);
nor U37832 (N_37832,N_26169,N_28697);
or U37833 (N_37833,N_28878,N_26557);
nor U37834 (N_37834,N_26188,N_21158);
and U37835 (N_37835,N_25097,N_29780);
or U37836 (N_37836,N_20190,N_29221);
or U37837 (N_37837,N_24698,N_28456);
or U37838 (N_37838,N_24749,N_27636);
xor U37839 (N_37839,N_23465,N_20753);
or U37840 (N_37840,N_29074,N_26451);
nand U37841 (N_37841,N_28785,N_26685);
xor U37842 (N_37842,N_20979,N_21154);
nand U37843 (N_37843,N_26246,N_27427);
nand U37844 (N_37844,N_29402,N_25522);
xor U37845 (N_37845,N_29259,N_27953);
nand U37846 (N_37846,N_22116,N_29652);
and U37847 (N_37847,N_21198,N_21564);
or U37848 (N_37848,N_21477,N_24495);
and U37849 (N_37849,N_27523,N_29048);
nand U37850 (N_37850,N_24519,N_25074);
and U37851 (N_37851,N_20111,N_25283);
xnor U37852 (N_37852,N_24079,N_25998);
nand U37853 (N_37853,N_28968,N_28825);
nor U37854 (N_37854,N_29472,N_28348);
nand U37855 (N_37855,N_28951,N_25642);
and U37856 (N_37856,N_27022,N_23303);
or U37857 (N_37857,N_25378,N_24525);
or U37858 (N_37858,N_27571,N_28568);
nand U37859 (N_37859,N_20280,N_28857);
nor U37860 (N_37860,N_21814,N_21284);
and U37861 (N_37861,N_22416,N_25999);
nor U37862 (N_37862,N_22349,N_24320);
nand U37863 (N_37863,N_27067,N_26403);
and U37864 (N_37864,N_21670,N_25897);
nor U37865 (N_37865,N_22334,N_29718);
or U37866 (N_37866,N_23407,N_25654);
xnor U37867 (N_37867,N_26824,N_20213);
or U37868 (N_37868,N_22715,N_27736);
nand U37869 (N_37869,N_22978,N_27671);
nor U37870 (N_37870,N_26588,N_23301);
nand U37871 (N_37871,N_25680,N_27956);
and U37872 (N_37872,N_28178,N_23318);
and U37873 (N_37873,N_26652,N_21529);
nor U37874 (N_37874,N_29381,N_25491);
or U37875 (N_37875,N_28191,N_21359);
nand U37876 (N_37876,N_22877,N_26125);
and U37877 (N_37877,N_28056,N_29174);
nor U37878 (N_37878,N_26899,N_28748);
nand U37879 (N_37879,N_24347,N_29618);
nor U37880 (N_37880,N_24685,N_28247);
nor U37881 (N_37881,N_22206,N_20616);
or U37882 (N_37882,N_28958,N_29120);
or U37883 (N_37883,N_28256,N_20594);
or U37884 (N_37884,N_24994,N_27833);
or U37885 (N_37885,N_23968,N_26639);
or U37886 (N_37886,N_23543,N_29317);
xnor U37887 (N_37887,N_25823,N_28006);
nor U37888 (N_37888,N_23862,N_28798);
and U37889 (N_37889,N_23187,N_23492);
or U37890 (N_37890,N_26494,N_27190);
or U37891 (N_37891,N_28885,N_29287);
nand U37892 (N_37892,N_25543,N_26239);
or U37893 (N_37893,N_28252,N_29049);
nand U37894 (N_37894,N_20427,N_24518);
or U37895 (N_37895,N_21040,N_20053);
nand U37896 (N_37896,N_22906,N_27406);
and U37897 (N_37897,N_26643,N_23360);
or U37898 (N_37898,N_28551,N_27018);
and U37899 (N_37899,N_27795,N_23694);
and U37900 (N_37900,N_20080,N_26923);
and U37901 (N_37901,N_22421,N_24848);
nand U37902 (N_37902,N_27725,N_28854);
xor U37903 (N_37903,N_21993,N_28670);
nor U37904 (N_37904,N_23754,N_28230);
and U37905 (N_37905,N_28050,N_27015);
or U37906 (N_37906,N_23008,N_22661);
and U37907 (N_37907,N_28306,N_25217);
nor U37908 (N_37908,N_21719,N_27854);
nor U37909 (N_37909,N_22368,N_22140);
xnor U37910 (N_37910,N_24131,N_28372);
and U37911 (N_37911,N_26155,N_25835);
or U37912 (N_37912,N_21914,N_20388);
xor U37913 (N_37913,N_22399,N_29465);
nand U37914 (N_37914,N_22507,N_29974);
nand U37915 (N_37915,N_22072,N_28344);
xor U37916 (N_37916,N_20572,N_20848);
or U37917 (N_37917,N_24024,N_29789);
nand U37918 (N_37918,N_24815,N_28691);
or U37919 (N_37919,N_22249,N_22567);
and U37920 (N_37920,N_20918,N_23040);
and U37921 (N_37921,N_20643,N_29922);
or U37922 (N_37922,N_28083,N_29518);
or U37923 (N_37923,N_24867,N_28152);
nor U37924 (N_37924,N_25635,N_22282);
or U37925 (N_37925,N_23793,N_23436);
nand U37926 (N_37926,N_28171,N_29773);
or U37927 (N_37927,N_26791,N_27671);
nand U37928 (N_37928,N_23785,N_28795);
and U37929 (N_37929,N_20782,N_22192);
nand U37930 (N_37930,N_23378,N_28863);
and U37931 (N_37931,N_25581,N_21849);
nor U37932 (N_37932,N_26521,N_22507);
nand U37933 (N_37933,N_28126,N_23634);
xor U37934 (N_37934,N_26028,N_20983);
xnor U37935 (N_37935,N_21163,N_23506);
nor U37936 (N_37936,N_26640,N_22427);
xnor U37937 (N_37937,N_29140,N_25217);
nor U37938 (N_37938,N_22823,N_27447);
and U37939 (N_37939,N_20605,N_23848);
nand U37940 (N_37940,N_23301,N_28761);
nand U37941 (N_37941,N_28820,N_23187);
nand U37942 (N_37942,N_24149,N_27570);
nor U37943 (N_37943,N_29885,N_23237);
or U37944 (N_37944,N_27182,N_24707);
xnor U37945 (N_37945,N_23735,N_24306);
nor U37946 (N_37946,N_29374,N_21897);
and U37947 (N_37947,N_28773,N_25535);
xnor U37948 (N_37948,N_24891,N_28147);
nor U37949 (N_37949,N_24726,N_22946);
xor U37950 (N_37950,N_23671,N_22858);
nand U37951 (N_37951,N_26253,N_28864);
nand U37952 (N_37952,N_29794,N_23528);
nor U37953 (N_37953,N_21907,N_23343);
nand U37954 (N_37954,N_20734,N_29162);
nor U37955 (N_37955,N_21451,N_21025);
nor U37956 (N_37956,N_21917,N_28539);
nand U37957 (N_37957,N_20772,N_26479);
and U37958 (N_37958,N_21358,N_23794);
xor U37959 (N_37959,N_21395,N_23701);
nand U37960 (N_37960,N_27931,N_27107);
and U37961 (N_37961,N_23453,N_22220);
or U37962 (N_37962,N_21415,N_24895);
and U37963 (N_37963,N_26716,N_28981);
nor U37964 (N_37964,N_27213,N_24865);
xor U37965 (N_37965,N_25769,N_28578);
nand U37966 (N_37966,N_26620,N_29328);
and U37967 (N_37967,N_25881,N_27258);
nor U37968 (N_37968,N_28048,N_27324);
or U37969 (N_37969,N_28259,N_25543);
and U37970 (N_37970,N_20365,N_20613);
xor U37971 (N_37971,N_28865,N_24382);
or U37972 (N_37972,N_21964,N_27818);
nor U37973 (N_37973,N_25782,N_25019);
nand U37974 (N_37974,N_22878,N_26195);
nand U37975 (N_37975,N_27247,N_26912);
nor U37976 (N_37976,N_28770,N_23981);
or U37977 (N_37977,N_29751,N_21286);
or U37978 (N_37978,N_23120,N_25426);
nor U37979 (N_37979,N_26062,N_26307);
nand U37980 (N_37980,N_27991,N_25037);
nand U37981 (N_37981,N_25612,N_21137);
and U37982 (N_37982,N_23177,N_29007);
nor U37983 (N_37983,N_24270,N_23712);
nor U37984 (N_37984,N_24959,N_26750);
nand U37985 (N_37985,N_21738,N_22945);
nor U37986 (N_37986,N_29920,N_27519);
or U37987 (N_37987,N_20374,N_22705);
and U37988 (N_37988,N_23472,N_23530);
nor U37989 (N_37989,N_27383,N_28666);
xor U37990 (N_37990,N_24357,N_24354);
and U37991 (N_37991,N_28323,N_23361);
nor U37992 (N_37992,N_24496,N_27847);
nand U37993 (N_37993,N_20719,N_21083);
and U37994 (N_37994,N_25393,N_25512);
and U37995 (N_37995,N_25148,N_20509);
xnor U37996 (N_37996,N_20895,N_29012);
nand U37997 (N_37997,N_28372,N_28787);
xor U37998 (N_37998,N_27626,N_25197);
nor U37999 (N_37999,N_21365,N_24889);
nand U38000 (N_38000,N_25464,N_20813);
xor U38001 (N_38001,N_21540,N_28718);
nor U38002 (N_38002,N_24946,N_27286);
xnor U38003 (N_38003,N_28779,N_29498);
nor U38004 (N_38004,N_20208,N_23472);
or U38005 (N_38005,N_22516,N_27062);
and U38006 (N_38006,N_20285,N_20074);
nand U38007 (N_38007,N_28321,N_22295);
and U38008 (N_38008,N_22388,N_28300);
nor U38009 (N_38009,N_26236,N_20913);
or U38010 (N_38010,N_27485,N_28471);
and U38011 (N_38011,N_25201,N_22914);
nor U38012 (N_38012,N_24791,N_27671);
or U38013 (N_38013,N_29499,N_22623);
nand U38014 (N_38014,N_22323,N_22674);
nor U38015 (N_38015,N_27409,N_23063);
or U38016 (N_38016,N_27395,N_20518);
and U38017 (N_38017,N_22773,N_28966);
nor U38018 (N_38018,N_27815,N_22310);
or U38019 (N_38019,N_25714,N_25814);
nand U38020 (N_38020,N_27576,N_20485);
and U38021 (N_38021,N_22283,N_28987);
xnor U38022 (N_38022,N_21513,N_26032);
and U38023 (N_38023,N_23303,N_20755);
nand U38024 (N_38024,N_20158,N_25917);
nor U38025 (N_38025,N_25097,N_28073);
nand U38026 (N_38026,N_28174,N_25919);
nand U38027 (N_38027,N_29928,N_28943);
and U38028 (N_38028,N_25465,N_29972);
or U38029 (N_38029,N_23375,N_23277);
xnor U38030 (N_38030,N_22235,N_26411);
xnor U38031 (N_38031,N_27503,N_28407);
nor U38032 (N_38032,N_28923,N_24595);
or U38033 (N_38033,N_25420,N_29774);
nand U38034 (N_38034,N_22643,N_24836);
or U38035 (N_38035,N_21387,N_20293);
and U38036 (N_38036,N_22356,N_23770);
nor U38037 (N_38037,N_25640,N_21506);
nand U38038 (N_38038,N_25387,N_29289);
and U38039 (N_38039,N_29776,N_24848);
and U38040 (N_38040,N_22634,N_26476);
nor U38041 (N_38041,N_21706,N_25685);
nand U38042 (N_38042,N_28872,N_26386);
xor U38043 (N_38043,N_25545,N_23334);
and U38044 (N_38044,N_21445,N_25221);
or U38045 (N_38045,N_25899,N_27304);
nor U38046 (N_38046,N_20058,N_23669);
or U38047 (N_38047,N_28039,N_22366);
xor U38048 (N_38048,N_28423,N_25415);
nor U38049 (N_38049,N_26138,N_21312);
or U38050 (N_38050,N_24935,N_22038);
nor U38051 (N_38051,N_25116,N_24736);
or U38052 (N_38052,N_26693,N_28062);
xor U38053 (N_38053,N_26614,N_26525);
nand U38054 (N_38054,N_20278,N_22284);
or U38055 (N_38055,N_26062,N_25356);
or U38056 (N_38056,N_24106,N_20157);
nor U38057 (N_38057,N_27872,N_22551);
nor U38058 (N_38058,N_24775,N_21514);
and U38059 (N_38059,N_22128,N_20255);
or U38060 (N_38060,N_29816,N_24813);
nand U38061 (N_38061,N_27055,N_20758);
nand U38062 (N_38062,N_27626,N_21610);
nand U38063 (N_38063,N_28039,N_25893);
or U38064 (N_38064,N_24270,N_20925);
nor U38065 (N_38065,N_24969,N_27467);
nand U38066 (N_38066,N_26486,N_29974);
or U38067 (N_38067,N_24842,N_22906);
nor U38068 (N_38068,N_22772,N_25750);
or U38069 (N_38069,N_25599,N_22429);
nand U38070 (N_38070,N_27365,N_23928);
and U38071 (N_38071,N_20152,N_28547);
or U38072 (N_38072,N_24393,N_22664);
or U38073 (N_38073,N_22890,N_20938);
or U38074 (N_38074,N_21604,N_22942);
and U38075 (N_38075,N_22546,N_24857);
nor U38076 (N_38076,N_23291,N_23748);
and U38077 (N_38077,N_28655,N_21240);
nor U38078 (N_38078,N_23909,N_25556);
and U38079 (N_38079,N_29386,N_27794);
xor U38080 (N_38080,N_24869,N_25948);
nor U38081 (N_38081,N_25738,N_24959);
nand U38082 (N_38082,N_24373,N_22752);
nor U38083 (N_38083,N_26472,N_24754);
xor U38084 (N_38084,N_24781,N_25583);
nand U38085 (N_38085,N_26610,N_24957);
nor U38086 (N_38086,N_24846,N_26484);
xor U38087 (N_38087,N_24945,N_21969);
or U38088 (N_38088,N_28252,N_20670);
nand U38089 (N_38089,N_26991,N_26912);
xnor U38090 (N_38090,N_26407,N_27682);
or U38091 (N_38091,N_23490,N_22735);
or U38092 (N_38092,N_21583,N_28499);
nor U38093 (N_38093,N_20764,N_25427);
nand U38094 (N_38094,N_22888,N_21662);
or U38095 (N_38095,N_20581,N_25717);
or U38096 (N_38096,N_23788,N_29252);
nand U38097 (N_38097,N_24238,N_24059);
xor U38098 (N_38098,N_29015,N_22705);
and U38099 (N_38099,N_28388,N_28491);
and U38100 (N_38100,N_23601,N_23435);
nand U38101 (N_38101,N_28844,N_20323);
xnor U38102 (N_38102,N_26750,N_27568);
xor U38103 (N_38103,N_23173,N_28946);
nor U38104 (N_38104,N_22689,N_23342);
nand U38105 (N_38105,N_27712,N_22455);
xor U38106 (N_38106,N_20590,N_20094);
xnor U38107 (N_38107,N_25025,N_27190);
or U38108 (N_38108,N_24470,N_27520);
and U38109 (N_38109,N_25669,N_24252);
nand U38110 (N_38110,N_26517,N_21676);
or U38111 (N_38111,N_29369,N_27687);
or U38112 (N_38112,N_27124,N_28115);
nor U38113 (N_38113,N_25025,N_22747);
xor U38114 (N_38114,N_27054,N_21020);
xor U38115 (N_38115,N_25642,N_28927);
or U38116 (N_38116,N_25971,N_28595);
nor U38117 (N_38117,N_21509,N_29520);
nand U38118 (N_38118,N_24566,N_23152);
nor U38119 (N_38119,N_24902,N_22138);
nor U38120 (N_38120,N_28502,N_20897);
or U38121 (N_38121,N_25563,N_20478);
or U38122 (N_38122,N_24880,N_29569);
xor U38123 (N_38123,N_20699,N_27320);
nand U38124 (N_38124,N_22964,N_23649);
xnor U38125 (N_38125,N_23006,N_28841);
nor U38126 (N_38126,N_26551,N_22646);
or U38127 (N_38127,N_28733,N_29795);
nand U38128 (N_38128,N_26459,N_23978);
nand U38129 (N_38129,N_29717,N_23456);
xnor U38130 (N_38130,N_20625,N_23379);
nand U38131 (N_38131,N_25396,N_26406);
nand U38132 (N_38132,N_24581,N_22319);
xor U38133 (N_38133,N_28352,N_22779);
or U38134 (N_38134,N_22395,N_24716);
or U38135 (N_38135,N_20514,N_28586);
xor U38136 (N_38136,N_23367,N_26476);
nand U38137 (N_38137,N_21817,N_20134);
nor U38138 (N_38138,N_22561,N_21049);
nand U38139 (N_38139,N_25618,N_23355);
xnor U38140 (N_38140,N_28217,N_20115);
nand U38141 (N_38141,N_22117,N_23197);
xor U38142 (N_38142,N_27017,N_26127);
and U38143 (N_38143,N_28916,N_20479);
xnor U38144 (N_38144,N_23236,N_29795);
and U38145 (N_38145,N_22704,N_22858);
xor U38146 (N_38146,N_23698,N_27658);
xor U38147 (N_38147,N_22463,N_22029);
and U38148 (N_38148,N_29227,N_29499);
and U38149 (N_38149,N_23713,N_21354);
xnor U38150 (N_38150,N_26887,N_27039);
xnor U38151 (N_38151,N_20238,N_21905);
nand U38152 (N_38152,N_29585,N_20456);
xor U38153 (N_38153,N_25446,N_24889);
xor U38154 (N_38154,N_28062,N_27181);
and U38155 (N_38155,N_28208,N_21404);
or U38156 (N_38156,N_21861,N_21789);
xnor U38157 (N_38157,N_27045,N_22583);
xnor U38158 (N_38158,N_22208,N_25421);
and U38159 (N_38159,N_23156,N_20944);
nor U38160 (N_38160,N_29631,N_22774);
and U38161 (N_38161,N_24526,N_23002);
xnor U38162 (N_38162,N_25686,N_21499);
and U38163 (N_38163,N_27222,N_28895);
or U38164 (N_38164,N_26970,N_23843);
xor U38165 (N_38165,N_28278,N_29083);
and U38166 (N_38166,N_24357,N_23313);
xnor U38167 (N_38167,N_22516,N_28055);
xor U38168 (N_38168,N_28043,N_27293);
and U38169 (N_38169,N_20972,N_29723);
nand U38170 (N_38170,N_25658,N_26093);
xor U38171 (N_38171,N_20950,N_24964);
or U38172 (N_38172,N_25304,N_20429);
and U38173 (N_38173,N_20266,N_28064);
nor U38174 (N_38174,N_21933,N_27615);
xnor U38175 (N_38175,N_26353,N_21964);
nor U38176 (N_38176,N_29156,N_29007);
and U38177 (N_38177,N_20852,N_26841);
nor U38178 (N_38178,N_22092,N_22652);
nor U38179 (N_38179,N_28304,N_29619);
nand U38180 (N_38180,N_27327,N_22993);
xor U38181 (N_38181,N_23280,N_28082);
nand U38182 (N_38182,N_28938,N_22724);
xnor U38183 (N_38183,N_26756,N_20069);
xnor U38184 (N_38184,N_29782,N_25809);
nor U38185 (N_38185,N_20054,N_28226);
nand U38186 (N_38186,N_24871,N_27716);
nand U38187 (N_38187,N_28593,N_25380);
or U38188 (N_38188,N_26510,N_23954);
xor U38189 (N_38189,N_28652,N_25987);
xor U38190 (N_38190,N_28669,N_29008);
or U38191 (N_38191,N_23573,N_22346);
nor U38192 (N_38192,N_25092,N_27946);
and U38193 (N_38193,N_20728,N_28466);
and U38194 (N_38194,N_28819,N_23281);
xor U38195 (N_38195,N_29202,N_24264);
xnor U38196 (N_38196,N_25573,N_21228);
xnor U38197 (N_38197,N_25756,N_22475);
nand U38198 (N_38198,N_26697,N_29910);
nand U38199 (N_38199,N_26865,N_21030);
and U38200 (N_38200,N_26201,N_22962);
nand U38201 (N_38201,N_21437,N_24791);
and U38202 (N_38202,N_29206,N_21015);
xor U38203 (N_38203,N_28351,N_26654);
or U38204 (N_38204,N_25084,N_23625);
or U38205 (N_38205,N_26690,N_22438);
nor U38206 (N_38206,N_21861,N_23581);
nand U38207 (N_38207,N_23105,N_26450);
nand U38208 (N_38208,N_24713,N_25138);
nor U38209 (N_38209,N_28024,N_22321);
xnor U38210 (N_38210,N_20692,N_26355);
xor U38211 (N_38211,N_25370,N_21306);
xor U38212 (N_38212,N_22877,N_26458);
and U38213 (N_38213,N_27450,N_20299);
nor U38214 (N_38214,N_20960,N_22067);
nand U38215 (N_38215,N_25122,N_25640);
nor U38216 (N_38216,N_27666,N_29588);
or U38217 (N_38217,N_27151,N_20213);
nor U38218 (N_38218,N_25022,N_23780);
or U38219 (N_38219,N_29950,N_24457);
nand U38220 (N_38220,N_23242,N_25286);
and U38221 (N_38221,N_29627,N_29833);
nor U38222 (N_38222,N_23316,N_23475);
nor U38223 (N_38223,N_28854,N_20520);
and U38224 (N_38224,N_20947,N_24539);
and U38225 (N_38225,N_24446,N_25035);
xnor U38226 (N_38226,N_20546,N_21631);
and U38227 (N_38227,N_27827,N_26139);
or U38228 (N_38228,N_28918,N_20458);
nand U38229 (N_38229,N_29790,N_22146);
or U38230 (N_38230,N_20253,N_23954);
nand U38231 (N_38231,N_24548,N_29668);
and U38232 (N_38232,N_26484,N_26704);
nand U38233 (N_38233,N_24137,N_21645);
xnor U38234 (N_38234,N_20535,N_21643);
xnor U38235 (N_38235,N_28457,N_25509);
nand U38236 (N_38236,N_20102,N_26002);
or U38237 (N_38237,N_22557,N_21926);
nand U38238 (N_38238,N_25904,N_26207);
nand U38239 (N_38239,N_26789,N_23636);
or U38240 (N_38240,N_21516,N_23016);
and U38241 (N_38241,N_29695,N_28963);
or U38242 (N_38242,N_24443,N_21706);
nand U38243 (N_38243,N_28736,N_28406);
nand U38244 (N_38244,N_26476,N_22137);
or U38245 (N_38245,N_28783,N_26224);
or U38246 (N_38246,N_20466,N_28086);
nor U38247 (N_38247,N_27544,N_25465);
or U38248 (N_38248,N_28802,N_20980);
nor U38249 (N_38249,N_29399,N_22728);
xnor U38250 (N_38250,N_25252,N_27930);
or U38251 (N_38251,N_24390,N_22674);
nor U38252 (N_38252,N_22838,N_28638);
nor U38253 (N_38253,N_23039,N_21819);
nor U38254 (N_38254,N_21569,N_28287);
and U38255 (N_38255,N_20003,N_24312);
nand U38256 (N_38256,N_27513,N_28720);
nand U38257 (N_38257,N_21427,N_25161);
nor U38258 (N_38258,N_21334,N_21794);
nor U38259 (N_38259,N_24519,N_29863);
nand U38260 (N_38260,N_22103,N_27011);
or U38261 (N_38261,N_28924,N_24363);
nor U38262 (N_38262,N_25373,N_23884);
or U38263 (N_38263,N_24628,N_20199);
or U38264 (N_38264,N_21178,N_22047);
or U38265 (N_38265,N_24325,N_23131);
and U38266 (N_38266,N_28539,N_27580);
and U38267 (N_38267,N_21511,N_21290);
and U38268 (N_38268,N_23928,N_24029);
or U38269 (N_38269,N_22314,N_24330);
or U38270 (N_38270,N_25946,N_25371);
nand U38271 (N_38271,N_29870,N_29128);
xnor U38272 (N_38272,N_22474,N_28906);
and U38273 (N_38273,N_24029,N_21510);
or U38274 (N_38274,N_28899,N_23644);
nor U38275 (N_38275,N_21246,N_28630);
nand U38276 (N_38276,N_26262,N_20697);
nand U38277 (N_38277,N_26841,N_20776);
or U38278 (N_38278,N_22211,N_29199);
and U38279 (N_38279,N_25255,N_27847);
and U38280 (N_38280,N_27613,N_28200);
nor U38281 (N_38281,N_29759,N_22834);
nand U38282 (N_38282,N_22352,N_25974);
nor U38283 (N_38283,N_22331,N_27598);
xor U38284 (N_38284,N_23229,N_27494);
nor U38285 (N_38285,N_28403,N_22834);
and U38286 (N_38286,N_24314,N_26553);
nor U38287 (N_38287,N_27107,N_20389);
nor U38288 (N_38288,N_20777,N_20922);
nand U38289 (N_38289,N_23963,N_23764);
nor U38290 (N_38290,N_25774,N_27703);
nor U38291 (N_38291,N_24788,N_27300);
xnor U38292 (N_38292,N_29192,N_23959);
nand U38293 (N_38293,N_28190,N_27449);
and U38294 (N_38294,N_29925,N_27647);
and U38295 (N_38295,N_25652,N_26392);
and U38296 (N_38296,N_22504,N_27753);
or U38297 (N_38297,N_25075,N_26720);
or U38298 (N_38298,N_28416,N_23724);
xnor U38299 (N_38299,N_23255,N_25014);
or U38300 (N_38300,N_24857,N_28774);
nor U38301 (N_38301,N_23404,N_28830);
or U38302 (N_38302,N_24339,N_27729);
xor U38303 (N_38303,N_22969,N_28182);
nor U38304 (N_38304,N_29762,N_24309);
xnor U38305 (N_38305,N_26266,N_28593);
and U38306 (N_38306,N_21833,N_27830);
or U38307 (N_38307,N_20801,N_22594);
nand U38308 (N_38308,N_27213,N_21257);
nor U38309 (N_38309,N_26024,N_21366);
nor U38310 (N_38310,N_22958,N_28218);
nor U38311 (N_38311,N_22037,N_22914);
nand U38312 (N_38312,N_26490,N_29664);
or U38313 (N_38313,N_25586,N_23645);
or U38314 (N_38314,N_24742,N_21311);
or U38315 (N_38315,N_25539,N_21267);
or U38316 (N_38316,N_22894,N_25151);
nor U38317 (N_38317,N_25967,N_21304);
and U38318 (N_38318,N_29940,N_25139);
or U38319 (N_38319,N_26672,N_21997);
or U38320 (N_38320,N_26737,N_27114);
xnor U38321 (N_38321,N_20447,N_24291);
and U38322 (N_38322,N_22131,N_23857);
nand U38323 (N_38323,N_27871,N_22593);
nor U38324 (N_38324,N_27408,N_27295);
or U38325 (N_38325,N_21776,N_26634);
xnor U38326 (N_38326,N_23673,N_23807);
nand U38327 (N_38327,N_21779,N_24767);
or U38328 (N_38328,N_21011,N_29697);
nor U38329 (N_38329,N_28546,N_24856);
or U38330 (N_38330,N_28882,N_24402);
nand U38331 (N_38331,N_26206,N_24982);
and U38332 (N_38332,N_25295,N_25628);
nor U38333 (N_38333,N_26004,N_26632);
xnor U38334 (N_38334,N_27462,N_23343);
or U38335 (N_38335,N_27826,N_23534);
and U38336 (N_38336,N_26010,N_22235);
nand U38337 (N_38337,N_20330,N_24321);
nor U38338 (N_38338,N_20271,N_25427);
or U38339 (N_38339,N_29752,N_27440);
nand U38340 (N_38340,N_24439,N_27108);
nand U38341 (N_38341,N_29787,N_23190);
and U38342 (N_38342,N_25963,N_24219);
and U38343 (N_38343,N_27447,N_24595);
nand U38344 (N_38344,N_20999,N_20606);
or U38345 (N_38345,N_25547,N_20863);
xnor U38346 (N_38346,N_20768,N_24705);
and U38347 (N_38347,N_23313,N_23777);
and U38348 (N_38348,N_22296,N_29636);
or U38349 (N_38349,N_29690,N_24039);
or U38350 (N_38350,N_22348,N_24819);
and U38351 (N_38351,N_24483,N_27850);
nor U38352 (N_38352,N_20231,N_22898);
nand U38353 (N_38353,N_20230,N_22883);
nand U38354 (N_38354,N_28939,N_20674);
and U38355 (N_38355,N_21690,N_26183);
or U38356 (N_38356,N_24176,N_24698);
and U38357 (N_38357,N_21604,N_23684);
nand U38358 (N_38358,N_25154,N_21739);
and U38359 (N_38359,N_21884,N_23474);
or U38360 (N_38360,N_25651,N_20476);
nand U38361 (N_38361,N_22840,N_24086);
xor U38362 (N_38362,N_26561,N_23782);
or U38363 (N_38363,N_28641,N_21256);
xnor U38364 (N_38364,N_27132,N_24214);
and U38365 (N_38365,N_23238,N_25925);
nor U38366 (N_38366,N_26876,N_22497);
nand U38367 (N_38367,N_29792,N_20894);
and U38368 (N_38368,N_27138,N_27118);
or U38369 (N_38369,N_21317,N_28611);
and U38370 (N_38370,N_20160,N_23575);
nor U38371 (N_38371,N_29044,N_25783);
and U38372 (N_38372,N_20430,N_27052);
nand U38373 (N_38373,N_29191,N_29239);
nand U38374 (N_38374,N_28618,N_21507);
or U38375 (N_38375,N_22367,N_28258);
nand U38376 (N_38376,N_23221,N_29537);
and U38377 (N_38377,N_27817,N_22628);
and U38378 (N_38378,N_22001,N_22403);
nand U38379 (N_38379,N_26925,N_22632);
or U38380 (N_38380,N_26200,N_27994);
nand U38381 (N_38381,N_25932,N_27410);
nand U38382 (N_38382,N_23264,N_28179);
and U38383 (N_38383,N_29363,N_21551);
nand U38384 (N_38384,N_25343,N_25546);
and U38385 (N_38385,N_22746,N_25602);
or U38386 (N_38386,N_27303,N_26286);
or U38387 (N_38387,N_22971,N_20972);
xnor U38388 (N_38388,N_22818,N_27537);
xnor U38389 (N_38389,N_27154,N_29609);
nor U38390 (N_38390,N_21159,N_29783);
or U38391 (N_38391,N_20078,N_21609);
nand U38392 (N_38392,N_21967,N_24910);
or U38393 (N_38393,N_20961,N_22921);
nor U38394 (N_38394,N_23740,N_25808);
or U38395 (N_38395,N_26840,N_25736);
and U38396 (N_38396,N_20980,N_22900);
or U38397 (N_38397,N_22635,N_28879);
nor U38398 (N_38398,N_24189,N_28781);
or U38399 (N_38399,N_24776,N_29871);
nor U38400 (N_38400,N_27274,N_24650);
nand U38401 (N_38401,N_23459,N_25160);
and U38402 (N_38402,N_23283,N_29888);
nand U38403 (N_38403,N_29254,N_21843);
xnor U38404 (N_38404,N_22983,N_21649);
and U38405 (N_38405,N_24382,N_27343);
or U38406 (N_38406,N_23922,N_28085);
nand U38407 (N_38407,N_20099,N_20343);
xnor U38408 (N_38408,N_25566,N_21471);
nor U38409 (N_38409,N_23354,N_29716);
nand U38410 (N_38410,N_23473,N_28887);
nand U38411 (N_38411,N_25707,N_23067);
or U38412 (N_38412,N_21731,N_26645);
nor U38413 (N_38413,N_27929,N_21241);
xor U38414 (N_38414,N_27310,N_21452);
and U38415 (N_38415,N_20531,N_21103);
nand U38416 (N_38416,N_20725,N_26060);
nor U38417 (N_38417,N_22062,N_20543);
nor U38418 (N_38418,N_26746,N_29033);
and U38419 (N_38419,N_28105,N_25626);
xnor U38420 (N_38420,N_28694,N_20583);
or U38421 (N_38421,N_26292,N_29626);
and U38422 (N_38422,N_24147,N_27266);
nand U38423 (N_38423,N_20986,N_21273);
nand U38424 (N_38424,N_24605,N_27735);
and U38425 (N_38425,N_29235,N_23876);
nand U38426 (N_38426,N_21816,N_21715);
nor U38427 (N_38427,N_26113,N_29003);
and U38428 (N_38428,N_24214,N_25305);
nand U38429 (N_38429,N_28790,N_23407);
nand U38430 (N_38430,N_26362,N_25006);
nor U38431 (N_38431,N_26040,N_29615);
and U38432 (N_38432,N_29476,N_26160);
nand U38433 (N_38433,N_29838,N_24495);
or U38434 (N_38434,N_25338,N_27810);
nor U38435 (N_38435,N_20014,N_25492);
or U38436 (N_38436,N_23615,N_29753);
nor U38437 (N_38437,N_25333,N_29953);
nand U38438 (N_38438,N_22523,N_20393);
nand U38439 (N_38439,N_26718,N_22525);
and U38440 (N_38440,N_21009,N_20978);
nand U38441 (N_38441,N_24809,N_21704);
xor U38442 (N_38442,N_27819,N_21593);
and U38443 (N_38443,N_21879,N_20066);
xor U38444 (N_38444,N_26876,N_21870);
xnor U38445 (N_38445,N_23920,N_24976);
or U38446 (N_38446,N_27520,N_27488);
and U38447 (N_38447,N_27166,N_24816);
nand U38448 (N_38448,N_21279,N_27141);
and U38449 (N_38449,N_25517,N_20206);
and U38450 (N_38450,N_23188,N_20983);
and U38451 (N_38451,N_28812,N_29126);
xor U38452 (N_38452,N_26294,N_23690);
or U38453 (N_38453,N_26384,N_28164);
xor U38454 (N_38454,N_21443,N_26723);
xor U38455 (N_38455,N_24265,N_24617);
nor U38456 (N_38456,N_22439,N_20678);
nand U38457 (N_38457,N_23461,N_27798);
nor U38458 (N_38458,N_22058,N_22424);
nand U38459 (N_38459,N_23986,N_25721);
nor U38460 (N_38460,N_27648,N_20952);
or U38461 (N_38461,N_29040,N_24246);
and U38462 (N_38462,N_26456,N_27473);
or U38463 (N_38463,N_24407,N_28319);
and U38464 (N_38464,N_23514,N_21549);
or U38465 (N_38465,N_23486,N_23016);
and U38466 (N_38466,N_27132,N_23300);
nand U38467 (N_38467,N_29944,N_21353);
xor U38468 (N_38468,N_25484,N_26018);
nor U38469 (N_38469,N_20592,N_28056);
nor U38470 (N_38470,N_21936,N_24453);
and U38471 (N_38471,N_22991,N_20719);
and U38472 (N_38472,N_24111,N_24575);
and U38473 (N_38473,N_26235,N_29180);
nor U38474 (N_38474,N_21492,N_20169);
and U38475 (N_38475,N_22043,N_24252);
and U38476 (N_38476,N_29033,N_20240);
and U38477 (N_38477,N_29525,N_28795);
nand U38478 (N_38478,N_24976,N_22794);
or U38479 (N_38479,N_22665,N_20693);
xor U38480 (N_38480,N_22522,N_29497);
xor U38481 (N_38481,N_22673,N_24208);
nand U38482 (N_38482,N_21670,N_24107);
nor U38483 (N_38483,N_21313,N_25367);
or U38484 (N_38484,N_20774,N_22656);
xnor U38485 (N_38485,N_20199,N_22067);
or U38486 (N_38486,N_27184,N_29893);
and U38487 (N_38487,N_24251,N_21794);
or U38488 (N_38488,N_28161,N_20457);
nor U38489 (N_38489,N_27369,N_26171);
nor U38490 (N_38490,N_29704,N_25492);
nand U38491 (N_38491,N_21818,N_21905);
or U38492 (N_38492,N_21537,N_24531);
xor U38493 (N_38493,N_26279,N_21597);
or U38494 (N_38494,N_20892,N_22751);
or U38495 (N_38495,N_29945,N_26781);
and U38496 (N_38496,N_28341,N_26274);
xor U38497 (N_38497,N_24002,N_26194);
nor U38498 (N_38498,N_22468,N_22393);
xor U38499 (N_38499,N_29534,N_20028);
nand U38500 (N_38500,N_21773,N_25504);
xor U38501 (N_38501,N_27818,N_28769);
xnor U38502 (N_38502,N_27420,N_25005);
xnor U38503 (N_38503,N_20297,N_21933);
or U38504 (N_38504,N_22245,N_25914);
or U38505 (N_38505,N_29340,N_23927);
xor U38506 (N_38506,N_24011,N_23241);
nor U38507 (N_38507,N_23232,N_28937);
nand U38508 (N_38508,N_25996,N_28194);
nor U38509 (N_38509,N_21565,N_26326);
nand U38510 (N_38510,N_27555,N_28760);
and U38511 (N_38511,N_20721,N_22339);
and U38512 (N_38512,N_29013,N_24739);
or U38513 (N_38513,N_25007,N_26134);
nand U38514 (N_38514,N_23340,N_23266);
xor U38515 (N_38515,N_26873,N_20528);
xor U38516 (N_38516,N_21035,N_28007);
xnor U38517 (N_38517,N_28802,N_24970);
nor U38518 (N_38518,N_21935,N_22043);
or U38519 (N_38519,N_22925,N_20817);
or U38520 (N_38520,N_26179,N_27396);
nand U38521 (N_38521,N_25875,N_27054);
nor U38522 (N_38522,N_24883,N_25857);
xnor U38523 (N_38523,N_26777,N_27891);
or U38524 (N_38524,N_24544,N_28375);
or U38525 (N_38525,N_24878,N_23689);
and U38526 (N_38526,N_28727,N_26983);
or U38527 (N_38527,N_27625,N_26986);
xnor U38528 (N_38528,N_24525,N_24078);
nor U38529 (N_38529,N_21028,N_25400);
nand U38530 (N_38530,N_28125,N_24800);
xnor U38531 (N_38531,N_27511,N_28374);
xor U38532 (N_38532,N_24616,N_28291);
nor U38533 (N_38533,N_20538,N_20975);
xor U38534 (N_38534,N_23361,N_25550);
or U38535 (N_38535,N_20626,N_28762);
xnor U38536 (N_38536,N_28824,N_22017);
xor U38537 (N_38537,N_27843,N_27293);
nor U38538 (N_38538,N_28754,N_25249);
nand U38539 (N_38539,N_23333,N_24341);
nor U38540 (N_38540,N_25818,N_28020);
or U38541 (N_38541,N_26039,N_20897);
and U38542 (N_38542,N_27337,N_28086);
and U38543 (N_38543,N_26388,N_26572);
nand U38544 (N_38544,N_25910,N_24404);
and U38545 (N_38545,N_28368,N_23260);
or U38546 (N_38546,N_22242,N_22435);
nand U38547 (N_38547,N_26245,N_29511);
nor U38548 (N_38548,N_23034,N_24345);
xor U38549 (N_38549,N_29708,N_22616);
or U38550 (N_38550,N_28502,N_22734);
xor U38551 (N_38551,N_26930,N_28244);
and U38552 (N_38552,N_22760,N_20015);
nor U38553 (N_38553,N_27592,N_20282);
xnor U38554 (N_38554,N_20908,N_24661);
or U38555 (N_38555,N_23063,N_26824);
xor U38556 (N_38556,N_26313,N_24311);
nand U38557 (N_38557,N_21313,N_26791);
or U38558 (N_38558,N_27650,N_27561);
nor U38559 (N_38559,N_25997,N_28143);
nand U38560 (N_38560,N_28757,N_20670);
nor U38561 (N_38561,N_25871,N_28587);
xnor U38562 (N_38562,N_28697,N_28310);
and U38563 (N_38563,N_26294,N_26819);
nor U38564 (N_38564,N_26145,N_29534);
or U38565 (N_38565,N_27707,N_22222);
and U38566 (N_38566,N_23510,N_28935);
or U38567 (N_38567,N_21136,N_24092);
nand U38568 (N_38568,N_20904,N_24223);
nor U38569 (N_38569,N_27107,N_27920);
or U38570 (N_38570,N_26974,N_20649);
or U38571 (N_38571,N_21526,N_26325);
nor U38572 (N_38572,N_28091,N_24087);
nor U38573 (N_38573,N_25884,N_21646);
and U38574 (N_38574,N_24415,N_28439);
xor U38575 (N_38575,N_25974,N_21441);
xnor U38576 (N_38576,N_21434,N_28064);
and U38577 (N_38577,N_23116,N_28547);
nor U38578 (N_38578,N_22540,N_20211);
and U38579 (N_38579,N_22646,N_21348);
nor U38580 (N_38580,N_21975,N_21655);
nand U38581 (N_38581,N_27878,N_24228);
xnor U38582 (N_38582,N_22391,N_25791);
xor U38583 (N_38583,N_24603,N_26992);
nand U38584 (N_38584,N_23880,N_21262);
nor U38585 (N_38585,N_26621,N_24552);
and U38586 (N_38586,N_21237,N_28862);
and U38587 (N_38587,N_25706,N_21243);
or U38588 (N_38588,N_20314,N_26999);
or U38589 (N_38589,N_20064,N_20280);
nor U38590 (N_38590,N_20735,N_29472);
nor U38591 (N_38591,N_22431,N_26055);
nand U38592 (N_38592,N_20205,N_25309);
or U38593 (N_38593,N_28364,N_23955);
or U38594 (N_38594,N_24877,N_20623);
or U38595 (N_38595,N_21559,N_22345);
nor U38596 (N_38596,N_21166,N_28112);
or U38597 (N_38597,N_25906,N_20989);
nor U38598 (N_38598,N_24946,N_22943);
xor U38599 (N_38599,N_24705,N_26318);
nor U38600 (N_38600,N_20612,N_23003);
nand U38601 (N_38601,N_21360,N_24794);
xnor U38602 (N_38602,N_27690,N_20078);
xnor U38603 (N_38603,N_23767,N_20155);
nor U38604 (N_38604,N_21335,N_25352);
and U38605 (N_38605,N_20820,N_24499);
or U38606 (N_38606,N_26247,N_20631);
xnor U38607 (N_38607,N_23621,N_27592);
or U38608 (N_38608,N_20168,N_24373);
nor U38609 (N_38609,N_28047,N_28130);
and U38610 (N_38610,N_27380,N_20577);
nand U38611 (N_38611,N_28710,N_23625);
or U38612 (N_38612,N_23966,N_27213);
and U38613 (N_38613,N_25856,N_23429);
and U38614 (N_38614,N_21316,N_27547);
nand U38615 (N_38615,N_29352,N_29333);
or U38616 (N_38616,N_25115,N_20186);
nand U38617 (N_38617,N_21258,N_28910);
and U38618 (N_38618,N_22348,N_25588);
or U38619 (N_38619,N_22711,N_25096);
nand U38620 (N_38620,N_25035,N_20733);
nand U38621 (N_38621,N_21246,N_21186);
nor U38622 (N_38622,N_24866,N_28186);
xor U38623 (N_38623,N_28657,N_28559);
or U38624 (N_38624,N_29495,N_25937);
xnor U38625 (N_38625,N_24727,N_25316);
nor U38626 (N_38626,N_22463,N_23599);
or U38627 (N_38627,N_25026,N_20876);
nor U38628 (N_38628,N_23128,N_22541);
nor U38629 (N_38629,N_24055,N_28675);
or U38630 (N_38630,N_23394,N_25234);
nand U38631 (N_38631,N_21903,N_20513);
nor U38632 (N_38632,N_23093,N_25696);
nand U38633 (N_38633,N_24444,N_26367);
xnor U38634 (N_38634,N_25643,N_29993);
and U38635 (N_38635,N_20798,N_23145);
and U38636 (N_38636,N_26243,N_26610);
and U38637 (N_38637,N_22696,N_26660);
nor U38638 (N_38638,N_24234,N_25929);
nand U38639 (N_38639,N_22383,N_29593);
and U38640 (N_38640,N_21410,N_20455);
and U38641 (N_38641,N_24375,N_28887);
or U38642 (N_38642,N_20895,N_26810);
xnor U38643 (N_38643,N_23852,N_28887);
nor U38644 (N_38644,N_28531,N_28970);
or U38645 (N_38645,N_29698,N_28632);
nor U38646 (N_38646,N_21791,N_23517);
and U38647 (N_38647,N_26116,N_24944);
nand U38648 (N_38648,N_22587,N_25743);
nand U38649 (N_38649,N_21294,N_24301);
nor U38650 (N_38650,N_25551,N_26431);
or U38651 (N_38651,N_28137,N_27115);
and U38652 (N_38652,N_23368,N_23990);
or U38653 (N_38653,N_25644,N_24186);
or U38654 (N_38654,N_23721,N_28842);
or U38655 (N_38655,N_23676,N_26334);
nor U38656 (N_38656,N_28467,N_23340);
xor U38657 (N_38657,N_26928,N_22651);
nor U38658 (N_38658,N_29666,N_28362);
or U38659 (N_38659,N_29749,N_25250);
nand U38660 (N_38660,N_20837,N_26639);
nand U38661 (N_38661,N_24983,N_22030);
nor U38662 (N_38662,N_20995,N_24463);
or U38663 (N_38663,N_29888,N_21917);
nand U38664 (N_38664,N_24445,N_28054);
nor U38665 (N_38665,N_25659,N_25082);
or U38666 (N_38666,N_29066,N_25108);
and U38667 (N_38667,N_23368,N_23063);
or U38668 (N_38668,N_23573,N_26461);
nand U38669 (N_38669,N_28150,N_29678);
nand U38670 (N_38670,N_27621,N_23441);
xor U38671 (N_38671,N_24959,N_20306);
nor U38672 (N_38672,N_27921,N_29433);
or U38673 (N_38673,N_23184,N_25563);
and U38674 (N_38674,N_26782,N_21947);
nor U38675 (N_38675,N_20277,N_21835);
nor U38676 (N_38676,N_29890,N_25201);
nor U38677 (N_38677,N_23422,N_27786);
and U38678 (N_38678,N_24463,N_27471);
and U38679 (N_38679,N_27733,N_20552);
or U38680 (N_38680,N_22097,N_20573);
and U38681 (N_38681,N_20692,N_20351);
nand U38682 (N_38682,N_24303,N_22745);
nor U38683 (N_38683,N_22858,N_20664);
or U38684 (N_38684,N_26276,N_24673);
nand U38685 (N_38685,N_27762,N_22768);
or U38686 (N_38686,N_20055,N_27398);
xor U38687 (N_38687,N_24452,N_20579);
or U38688 (N_38688,N_24348,N_22264);
nand U38689 (N_38689,N_27962,N_29344);
xnor U38690 (N_38690,N_24800,N_28175);
nand U38691 (N_38691,N_24522,N_21610);
nor U38692 (N_38692,N_29565,N_24377);
and U38693 (N_38693,N_24597,N_20125);
xor U38694 (N_38694,N_28314,N_29295);
xnor U38695 (N_38695,N_20234,N_29552);
and U38696 (N_38696,N_26663,N_22408);
nand U38697 (N_38697,N_28045,N_27613);
and U38698 (N_38698,N_26155,N_26899);
and U38699 (N_38699,N_25866,N_22455);
nand U38700 (N_38700,N_27375,N_22570);
nand U38701 (N_38701,N_22122,N_22029);
nor U38702 (N_38702,N_22561,N_21634);
nor U38703 (N_38703,N_26775,N_28369);
nand U38704 (N_38704,N_29168,N_22629);
nor U38705 (N_38705,N_26201,N_21339);
nand U38706 (N_38706,N_23596,N_27409);
nor U38707 (N_38707,N_29654,N_20959);
nand U38708 (N_38708,N_26103,N_27298);
nor U38709 (N_38709,N_28459,N_28782);
and U38710 (N_38710,N_26044,N_21145);
and U38711 (N_38711,N_21202,N_26213);
nor U38712 (N_38712,N_24338,N_24189);
or U38713 (N_38713,N_27124,N_25682);
and U38714 (N_38714,N_27706,N_23996);
or U38715 (N_38715,N_26817,N_20832);
nand U38716 (N_38716,N_24835,N_29827);
and U38717 (N_38717,N_21624,N_27628);
nor U38718 (N_38718,N_25247,N_27088);
nand U38719 (N_38719,N_27018,N_27293);
xnor U38720 (N_38720,N_25435,N_25875);
nor U38721 (N_38721,N_20118,N_27594);
xor U38722 (N_38722,N_20400,N_25256);
nand U38723 (N_38723,N_25226,N_29825);
nand U38724 (N_38724,N_24945,N_20325);
nand U38725 (N_38725,N_23629,N_28968);
xnor U38726 (N_38726,N_27550,N_26575);
xor U38727 (N_38727,N_26810,N_24839);
and U38728 (N_38728,N_27099,N_22628);
nand U38729 (N_38729,N_23560,N_26829);
or U38730 (N_38730,N_20935,N_22138);
nor U38731 (N_38731,N_26598,N_27725);
xnor U38732 (N_38732,N_25684,N_28477);
or U38733 (N_38733,N_29955,N_29126);
nor U38734 (N_38734,N_29751,N_26578);
and U38735 (N_38735,N_22592,N_24633);
or U38736 (N_38736,N_28913,N_22710);
nor U38737 (N_38737,N_23340,N_26130);
nor U38738 (N_38738,N_27264,N_21866);
or U38739 (N_38739,N_26380,N_20437);
nor U38740 (N_38740,N_25219,N_21448);
nor U38741 (N_38741,N_22154,N_22506);
or U38742 (N_38742,N_28164,N_20074);
and U38743 (N_38743,N_22601,N_25765);
xnor U38744 (N_38744,N_21929,N_26615);
and U38745 (N_38745,N_24091,N_29634);
nand U38746 (N_38746,N_23698,N_26156);
nand U38747 (N_38747,N_20017,N_21240);
and U38748 (N_38748,N_28294,N_20504);
nand U38749 (N_38749,N_22119,N_22720);
nor U38750 (N_38750,N_28732,N_29461);
xor U38751 (N_38751,N_29972,N_28913);
nand U38752 (N_38752,N_28388,N_21456);
nor U38753 (N_38753,N_25861,N_27112);
xor U38754 (N_38754,N_24172,N_21662);
nor U38755 (N_38755,N_26614,N_22931);
nand U38756 (N_38756,N_29509,N_21622);
nand U38757 (N_38757,N_28024,N_22399);
or U38758 (N_38758,N_21951,N_23770);
and U38759 (N_38759,N_24216,N_26163);
xnor U38760 (N_38760,N_29867,N_22226);
and U38761 (N_38761,N_27756,N_25052);
nand U38762 (N_38762,N_20457,N_27199);
xor U38763 (N_38763,N_29388,N_22166);
and U38764 (N_38764,N_21712,N_23475);
xor U38765 (N_38765,N_29435,N_29123);
nand U38766 (N_38766,N_22128,N_22657);
and U38767 (N_38767,N_22995,N_21796);
or U38768 (N_38768,N_25217,N_20714);
or U38769 (N_38769,N_27526,N_29735);
nand U38770 (N_38770,N_23295,N_28088);
nor U38771 (N_38771,N_21522,N_24672);
and U38772 (N_38772,N_27639,N_23530);
xor U38773 (N_38773,N_24336,N_24338);
or U38774 (N_38774,N_29738,N_21236);
nor U38775 (N_38775,N_29991,N_25729);
nand U38776 (N_38776,N_24417,N_28197);
or U38777 (N_38777,N_28425,N_23929);
or U38778 (N_38778,N_26639,N_22911);
or U38779 (N_38779,N_20554,N_27677);
nor U38780 (N_38780,N_28254,N_20682);
nor U38781 (N_38781,N_23186,N_29437);
or U38782 (N_38782,N_27143,N_25002);
nand U38783 (N_38783,N_28376,N_23125);
xor U38784 (N_38784,N_26660,N_21746);
or U38785 (N_38785,N_21289,N_20979);
xnor U38786 (N_38786,N_22049,N_28759);
nand U38787 (N_38787,N_29536,N_24430);
xor U38788 (N_38788,N_29326,N_29435);
and U38789 (N_38789,N_29948,N_23412);
xor U38790 (N_38790,N_21180,N_28302);
nor U38791 (N_38791,N_28466,N_21043);
nand U38792 (N_38792,N_20999,N_27763);
nand U38793 (N_38793,N_26073,N_25162);
xor U38794 (N_38794,N_29065,N_24233);
nand U38795 (N_38795,N_21174,N_26325);
and U38796 (N_38796,N_28326,N_20539);
and U38797 (N_38797,N_29041,N_22020);
or U38798 (N_38798,N_26440,N_27052);
nand U38799 (N_38799,N_20315,N_20549);
and U38800 (N_38800,N_27404,N_25083);
or U38801 (N_38801,N_23259,N_26197);
and U38802 (N_38802,N_29650,N_21560);
or U38803 (N_38803,N_22902,N_28750);
nand U38804 (N_38804,N_28274,N_21424);
xnor U38805 (N_38805,N_24781,N_26092);
nor U38806 (N_38806,N_23968,N_20919);
nor U38807 (N_38807,N_23995,N_20287);
xor U38808 (N_38808,N_21474,N_28101);
nand U38809 (N_38809,N_26840,N_25978);
or U38810 (N_38810,N_20336,N_22920);
and U38811 (N_38811,N_20128,N_28822);
nor U38812 (N_38812,N_27128,N_20307);
and U38813 (N_38813,N_29476,N_20730);
nand U38814 (N_38814,N_25800,N_23905);
nand U38815 (N_38815,N_27169,N_23021);
or U38816 (N_38816,N_28714,N_21021);
and U38817 (N_38817,N_22025,N_23315);
and U38818 (N_38818,N_24980,N_23357);
or U38819 (N_38819,N_28745,N_27588);
nand U38820 (N_38820,N_25553,N_20155);
and U38821 (N_38821,N_29772,N_29566);
or U38822 (N_38822,N_29985,N_22133);
xnor U38823 (N_38823,N_26901,N_22073);
nand U38824 (N_38824,N_27929,N_24296);
xnor U38825 (N_38825,N_22638,N_20455);
or U38826 (N_38826,N_20026,N_29077);
or U38827 (N_38827,N_22417,N_23031);
nor U38828 (N_38828,N_25060,N_24650);
xnor U38829 (N_38829,N_28071,N_26503);
nor U38830 (N_38830,N_22626,N_24241);
and U38831 (N_38831,N_24091,N_24972);
xor U38832 (N_38832,N_29606,N_20788);
or U38833 (N_38833,N_29225,N_27914);
nor U38834 (N_38834,N_23916,N_28972);
and U38835 (N_38835,N_22712,N_23986);
nand U38836 (N_38836,N_26308,N_21882);
nor U38837 (N_38837,N_23527,N_21180);
and U38838 (N_38838,N_24811,N_26681);
nand U38839 (N_38839,N_24911,N_28314);
or U38840 (N_38840,N_23584,N_25424);
nand U38841 (N_38841,N_26527,N_25983);
nor U38842 (N_38842,N_24352,N_26070);
or U38843 (N_38843,N_25831,N_22692);
nand U38844 (N_38844,N_26428,N_29670);
xnor U38845 (N_38845,N_20700,N_28790);
and U38846 (N_38846,N_28482,N_24300);
xor U38847 (N_38847,N_28804,N_29706);
nor U38848 (N_38848,N_29433,N_25295);
xor U38849 (N_38849,N_24174,N_24768);
or U38850 (N_38850,N_22511,N_24430);
or U38851 (N_38851,N_28275,N_21746);
xnor U38852 (N_38852,N_20602,N_26908);
xor U38853 (N_38853,N_25065,N_21209);
or U38854 (N_38854,N_21533,N_28457);
xor U38855 (N_38855,N_22630,N_21544);
nand U38856 (N_38856,N_23148,N_22729);
and U38857 (N_38857,N_23768,N_25804);
nand U38858 (N_38858,N_22975,N_24882);
nor U38859 (N_38859,N_20637,N_23013);
or U38860 (N_38860,N_22412,N_26048);
or U38861 (N_38861,N_23294,N_21011);
xnor U38862 (N_38862,N_22531,N_21091);
or U38863 (N_38863,N_21944,N_21142);
xor U38864 (N_38864,N_29209,N_28993);
nor U38865 (N_38865,N_20731,N_28307);
nand U38866 (N_38866,N_26040,N_20836);
nand U38867 (N_38867,N_22283,N_25843);
xor U38868 (N_38868,N_22293,N_26986);
and U38869 (N_38869,N_23151,N_29397);
nand U38870 (N_38870,N_21787,N_20396);
and U38871 (N_38871,N_24845,N_29673);
and U38872 (N_38872,N_20462,N_26462);
or U38873 (N_38873,N_24588,N_26825);
and U38874 (N_38874,N_20665,N_23908);
xnor U38875 (N_38875,N_21402,N_22914);
nor U38876 (N_38876,N_26567,N_21103);
or U38877 (N_38877,N_28828,N_26960);
nor U38878 (N_38878,N_23487,N_22846);
and U38879 (N_38879,N_23595,N_25224);
and U38880 (N_38880,N_20997,N_22171);
or U38881 (N_38881,N_29025,N_26239);
or U38882 (N_38882,N_20617,N_24559);
xor U38883 (N_38883,N_21468,N_23029);
or U38884 (N_38884,N_26743,N_29201);
nand U38885 (N_38885,N_24644,N_23655);
xnor U38886 (N_38886,N_21996,N_20272);
xor U38887 (N_38887,N_24175,N_22953);
and U38888 (N_38888,N_25007,N_25150);
nand U38889 (N_38889,N_25908,N_22355);
nor U38890 (N_38890,N_20056,N_25886);
and U38891 (N_38891,N_25269,N_28792);
nor U38892 (N_38892,N_27012,N_21906);
and U38893 (N_38893,N_28550,N_22998);
nand U38894 (N_38894,N_27650,N_27850);
nand U38895 (N_38895,N_26118,N_22387);
and U38896 (N_38896,N_24980,N_26448);
and U38897 (N_38897,N_25023,N_20916);
xor U38898 (N_38898,N_27542,N_24536);
nor U38899 (N_38899,N_23750,N_21350);
and U38900 (N_38900,N_26032,N_23597);
nand U38901 (N_38901,N_29788,N_26593);
and U38902 (N_38902,N_27509,N_27506);
nand U38903 (N_38903,N_25252,N_22425);
nor U38904 (N_38904,N_29099,N_26010);
and U38905 (N_38905,N_24036,N_24191);
or U38906 (N_38906,N_26591,N_22161);
and U38907 (N_38907,N_27853,N_25132);
or U38908 (N_38908,N_26810,N_26185);
or U38909 (N_38909,N_21971,N_27807);
and U38910 (N_38910,N_27810,N_26160);
nand U38911 (N_38911,N_26506,N_26836);
and U38912 (N_38912,N_20865,N_25805);
and U38913 (N_38913,N_22970,N_20388);
nor U38914 (N_38914,N_20854,N_25858);
and U38915 (N_38915,N_21148,N_27384);
nor U38916 (N_38916,N_27891,N_22719);
nor U38917 (N_38917,N_27611,N_23860);
nand U38918 (N_38918,N_28880,N_21655);
and U38919 (N_38919,N_21032,N_21483);
xor U38920 (N_38920,N_22615,N_28991);
or U38921 (N_38921,N_28397,N_23084);
or U38922 (N_38922,N_29171,N_20049);
or U38923 (N_38923,N_23614,N_24873);
xor U38924 (N_38924,N_29014,N_23380);
and U38925 (N_38925,N_28176,N_24838);
nand U38926 (N_38926,N_28090,N_26864);
xor U38927 (N_38927,N_26452,N_27766);
or U38928 (N_38928,N_23962,N_27128);
or U38929 (N_38929,N_22020,N_26154);
xor U38930 (N_38930,N_24417,N_25813);
and U38931 (N_38931,N_24860,N_28459);
and U38932 (N_38932,N_25027,N_28870);
or U38933 (N_38933,N_27211,N_25865);
nand U38934 (N_38934,N_25775,N_27204);
nand U38935 (N_38935,N_22043,N_20626);
and U38936 (N_38936,N_23248,N_23682);
nor U38937 (N_38937,N_25587,N_25408);
nand U38938 (N_38938,N_20317,N_28891);
xor U38939 (N_38939,N_25268,N_20933);
nand U38940 (N_38940,N_22751,N_24621);
nand U38941 (N_38941,N_23005,N_25777);
or U38942 (N_38942,N_28035,N_25767);
or U38943 (N_38943,N_26067,N_27646);
nor U38944 (N_38944,N_23090,N_23802);
nand U38945 (N_38945,N_29390,N_24562);
and U38946 (N_38946,N_29941,N_29617);
xor U38947 (N_38947,N_24745,N_20497);
nand U38948 (N_38948,N_26238,N_20825);
or U38949 (N_38949,N_28992,N_21401);
or U38950 (N_38950,N_20470,N_25370);
or U38951 (N_38951,N_29442,N_20618);
or U38952 (N_38952,N_22242,N_23503);
nand U38953 (N_38953,N_21771,N_28142);
nor U38954 (N_38954,N_20342,N_23098);
or U38955 (N_38955,N_23719,N_29859);
and U38956 (N_38956,N_29754,N_24382);
xnor U38957 (N_38957,N_29208,N_27779);
nor U38958 (N_38958,N_22566,N_20625);
xnor U38959 (N_38959,N_27058,N_25828);
or U38960 (N_38960,N_21023,N_24467);
nand U38961 (N_38961,N_28254,N_27656);
xor U38962 (N_38962,N_21967,N_21249);
and U38963 (N_38963,N_27107,N_25890);
or U38964 (N_38964,N_25942,N_28506);
xor U38965 (N_38965,N_24666,N_24047);
and U38966 (N_38966,N_22687,N_23863);
nor U38967 (N_38967,N_25117,N_29685);
nand U38968 (N_38968,N_24336,N_24774);
xnor U38969 (N_38969,N_23976,N_28543);
and U38970 (N_38970,N_21404,N_21708);
nor U38971 (N_38971,N_28323,N_24209);
or U38972 (N_38972,N_28783,N_25650);
xnor U38973 (N_38973,N_21112,N_20057);
and U38974 (N_38974,N_23181,N_20035);
and U38975 (N_38975,N_28064,N_21634);
or U38976 (N_38976,N_23714,N_21000);
or U38977 (N_38977,N_20502,N_24334);
nand U38978 (N_38978,N_27683,N_21647);
and U38979 (N_38979,N_20757,N_25622);
or U38980 (N_38980,N_25616,N_23165);
or U38981 (N_38981,N_28228,N_21499);
or U38982 (N_38982,N_27876,N_26222);
xor U38983 (N_38983,N_21176,N_23037);
nand U38984 (N_38984,N_21350,N_26597);
nor U38985 (N_38985,N_23606,N_21455);
nor U38986 (N_38986,N_28431,N_23077);
or U38987 (N_38987,N_23240,N_24514);
nand U38988 (N_38988,N_28158,N_24455);
xnor U38989 (N_38989,N_28616,N_25441);
and U38990 (N_38990,N_24433,N_27736);
and U38991 (N_38991,N_28132,N_24464);
or U38992 (N_38992,N_25574,N_20247);
or U38993 (N_38993,N_26061,N_25522);
xnor U38994 (N_38994,N_29210,N_23031);
nor U38995 (N_38995,N_24460,N_29060);
and U38996 (N_38996,N_26553,N_21516);
xnor U38997 (N_38997,N_22305,N_21552);
nor U38998 (N_38998,N_27849,N_29012);
nand U38999 (N_38999,N_25433,N_28161);
or U39000 (N_39000,N_28361,N_27853);
xor U39001 (N_39001,N_21040,N_23847);
nor U39002 (N_39002,N_20106,N_25717);
and U39003 (N_39003,N_24270,N_26209);
xnor U39004 (N_39004,N_23724,N_21729);
nor U39005 (N_39005,N_29127,N_22206);
or U39006 (N_39006,N_27517,N_29990);
xnor U39007 (N_39007,N_28804,N_28932);
and U39008 (N_39008,N_23623,N_28781);
nor U39009 (N_39009,N_21717,N_26912);
nand U39010 (N_39010,N_26038,N_25754);
nand U39011 (N_39011,N_25665,N_26566);
or U39012 (N_39012,N_29324,N_22619);
nand U39013 (N_39013,N_29231,N_24465);
xnor U39014 (N_39014,N_21113,N_26433);
nor U39015 (N_39015,N_20003,N_24487);
or U39016 (N_39016,N_29135,N_22301);
xnor U39017 (N_39017,N_29402,N_21422);
and U39018 (N_39018,N_24572,N_24173);
xnor U39019 (N_39019,N_20090,N_21361);
nor U39020 (N_39020,N_20836,N_24160);
or U39021 (N_39021,N_25936,N_22023);
or U39022 (N_39022,N_22057,N_28807);
and U39023 (N_39023,N_20558,N_22487);
and U39024 (N_39024,N_20935,N_26541);
or U39025 (N_39025,N_25026,N_26300);
nand U39026 (N_39026,N_21693,N_21097);
nor U39027 (N_39027,N_22892,N_22783);
nor U39028 (N_39028,N_25413,N_27821);
or U39029 (N_39029,N_25420,N_29258);
nor U39030 (N_39030,N_29241,N_24902);
and U39031 (N_39031,N_22220,N_23885);
nor U39032 (N_39032,N_21740,N_23479);
nand U39033 (N_39033,N_22526,N_28261);
or U39034 (N_39034,N_28204,N_23933);
xnor U39035 (N_39035,N_26240,N_26456);
xnor U39036 (N_39036,N_26965,N_22442);
and U39037 (N_39037,N_25806,N_23389);
nand U39038 (N_39038,N_28416,N_25689);
nor U39039 (N_39039,N_24718,N_28063);
and U39040 (N_39040,N_25364,N_22825);
xnor U39041 (N_39041,N_28825,N_28740);
nor U39042 (N_39042,N_23233,N_25675);
and U39043 (N_39043,N_28850,N_20973);
nor U39044 (N_39044,N_21518,N_20733);
xnor U39045 (N_39045,N_23992,N_29353);
nand U39046 (N_39046,N_29212,N_26072);
or U39047 (N_39047,N_28482,N_22744);
and U39048 (N_39048,N_22487,N_21000);
and U39049 (N_39049,N_28433,N_29927);
nor U39050 (N_39050,N_27412,N_20000);
or U39051 (N_39051,N_21393,N_22660);
nand U39052 (N_39052,N_20328,N_20722);
xor U39053 (N_39053,N_23056,N_26197);
or U39054 (N_39054,N_28154,N_29135);
and U39055 (N_39055,N_29807,N_22582);
nor U39056 (N_39056,N_23115,N_21381);
nand U39057 (N_39057,N_28296,N_23161);
or U39058 (N_39058,N_23992,N_24183);
and U39059 (N_39059,N_22764,N_26797);
nand U39060 (N_39060,N_23329,N_23914);
xnor U39061 (N_39061,N_20659,N_22913);
xor U39062 (N_39062,N_25533,N_26820);
and U39063 (N_39063,N_24736,N_25852);
xor U39064 (N_39064,N_26748,N_21778);
nor U39065 (N_39065,N_22486,N_28078);
xnor U39066 (N_39066,N_27134,N_21630);
nand U39067 (N_39067,N_24732,N_27932);
and U39068 (N_39068,N_22417,N_26054);
or U39069 (N_39069,N_29582,N_29467);
and U39070 (N_39070,N_20259,N_22796);
or U39071 (N_39071,N_22372,N_29721);
xor U39072 (N_39072,N_24553,N_29624);
and U39073 (N_39073,N_27610,N_20674);
and U39074 (N_39074,N_27100,N_26003);
nor U39075 (N_39075,N_21472,N_20483);
or U39076 (N_39076,N_21369,N_23085);
and U39077 (N_39077,N_25170,N_22850);
nand U39078 (N_39078,N_22292,N_20615);
nor U39079 (N_39079,N_29372,N_20344);
or U39080 (N_39080,N_22420,N_24846);
or U39081 (N_39081,N_27179,N_22194);
xor U39082 (N_39082,N_20733,N_20764);
nand U39083 (N_39083,N_21691,N_22181);
nand U39084 (N_39084,N_21844,N_28854);
nor U39085 (N_39085,N_27254,N_21843);
and U39086 (N_39086,N_28766,N_28459);
xor U39087 (N_39087,N_25343,N_28220);
and U39088 (N_39088,N_20525,N_23104);
and U39089 (N_39089,N_20663,N_23068);
and U39090 (N_39090,N_28354,N_23297);
xor U39091 (N_39091,N_21736,N_23992);
or U39092 (N_39092,N_22248,N_20167);
nand U39093 (N_39093,N_23070,N_28065);
and U39094 (N_39094,N_29905,N_29238);
nor U39095 (N_39095,N_27952,N_24067);
and U39096 (N_39096,N_26470,N_28751);
xor U39097 (N_39097,N_26236,N_27103);
or U39098 (N_39098,N_27672,N_29060);
and U39099 (N_39099,N_27191,N_22130);
nand U39100 (N_39100,N_21053,N_24506);
nand U39101 (N_39101,N_26041,N_20953);
and U39102 (N_39102,N_20177,N_28390);
nand U39103 (N_39103,N_23029,N_21115);
or U39104 (N_39104,N_26295,N_23760);
xnor U39105 (N_39105,N_25748,N_25745);
xnor U39106 (N_39106,N_25918,N_24821);
nor U39107 (N_39107,N_24742,N_24141);
or U39108 (N_39108,N_21600,N_23436);
and U39109 (N_39109,N_21039,N_24274);
or U39110 (N_39110,N_27560,N_26641);
nor U39111 (N_39111,N_28149,N_23957);
or U39112 (N_39112,N_28339,N_26038);
nor U39113 (N_39113,N_22779,N_28821);
and U39114 (N_39114,N_20549,N_22399);
or U39115 (N_39115,N_27732,N_29097);
and U39116 (N_39116,N_25205,N_28018);
nor U39117 (N_39117,N_23006,N_26556);
nand U39118 (N_39118,N_24741,N_27115);
or U39119 (N_39119,N_28099,N_25526);
or U39120 (N_39120,N_21221,N_20048);
xnor U39121 (N_39121,N_28025,N_24196);
nand U39122 (N_39122,N_24716,N_25690);
nor U39123 (N_39123,N_23991,N_22752);
or U39124 (N_39124,N_27509,N_24460);
nand U39125 (N_39125,N_29507,N_20630);
and U39126 (N_39126,N_20463,N_26975);
nor U39127 (N_39127,N_23925,N_21550);
xnor U39128 (N_39128,N_21452,N_20599);
nor U39129 (N_39129,N_25718,N_23435);
xor U39130 (N_39130,N_20318,N_27132);
nand U39131 (N_39131,N_27234,N_21776);
xnor U39132 (N_39132,N_26339,N_23921);
xor U39133 (N_39133,N_23381,N_27028);
xnor U39134 (N_39134,N_20021,N_21250);
and U39135 (N_39135,N_20939,N_24280);
and U39136 (N_39136,N_20351,N_23547);
and U39137 (N_39137,N_21737,N_25096);
and U39138 (N_39138,N_25059,N_29797);
nor U39139 (N_39139,N_25974,N_20176);
nor U39140 (N_39140,N_25538,N_20867);
or U39141 (N_39141,N_29321,N_20575);
or U39142 (N_39142,N_26831,N_29314);
nor U39143 (N_39143,N_25230,N_27390);
or U39144 (N_39144,N_24503,N_28511);
or U39145 (N_39145,N_21331,N_25210);
nand U39146 (N_39146,N_28579,N_26787);
nor U39147 (N_39147,N_20039,N_20634);
or U39148 (N_39148,N_26755,N_21507);
and U39149 (N_39149,N_24555,N_21535);
and U39150 (N_39150,N_22289,N_26902);
or U39151 (N_39151,N_28326,N_25032);
and U39152 (N_39152,N_20999,N_20875);
nor U39153 (N_39153,N_23416,N_21700);
nor U39154 (N_39154,N_20375,N_24520);
xor U39155 (N_39155,N_23294,N_24962);
nand U39156 (N_39156,N_25333,N_23083);
nor U39157 (N_39157,N_20841,N_24023);
nand U39158 (N_39158,N_21542,N_26934);
nor U39159 (N_39159,N_29809,N_21040);
and U39160 (N_39160,N_20854,N_25157);
xnor U39161 (N_39161,N_23796,N_27443);
and U39162 (N_39162,N_26946,N_23647);
and U39163 (N_39163,N_24430,N_25956);
nand U39164 (N_39164,N_25323,N_28699);
nand U39165 (N_39165,N_25857,N_28136);
xnor U39166 (N_39166,N_26214,N_23229);
and U39167 (N_39167,N_27795,N_27096);
and U39168 (N_39168,N_22441,N_21817);
and U39169 (N_39169,N_28502,N_26385);
nand U39170 (N_39170,N_21078,N_28994);
nor U39171 (N_39171,N_23060,N_20439);
and U39172 (N_39172,N_21697,N_29028);
nor U39173 (N_39173,N_27772,N_20208);
and U39174 (N_39174,N_20338,N_28677);
nor U39175 (N_39175,N_26039,N_26461);
and U39176 (N_39176,N_27402,N_22902);
xnor U39177 (N_39177,N_24716,N_26759);
or U39178 (N_39178,N_21351,N_26601);
or U39179 (N_39179,N_22488,N_20823);
nor U39180 (N_39180,N_25408,N_27035);
nand U39181 (N_39181,N_29223,N_23298);
nand U39182 (N_39182,N_25580,N_27846);
and U39183 (N_39183,N_26266,N_23310);
and U39184 (N_39184,N_21156,N_23579);
xnor U39185 (N_39185,N_20135,N_22227);
xor U39186 (N_39186,N_26590,N_28539);
nand U39187 (N_39187,N_21850,N_25067);
or U39188 (N_39188,N_23360,N_27289);
or U39189 (N_39189,N_23387,N_26096);
nor U39190 (N_39190,N_26967,N_26550);
xor U39191 (N_39191,N_23484,N_23432);
and U39192 (N_39192,N_26658,N_28467);
nand U39193 (N_39193,N_29701,N_25749);
nor U39194 (N_39194,N_20187,N_24377);
nor U39195 (N_39195,N_21531,N_27180);
and U39196 (N_39196,N_27061,N_29374);
nor U39197 (N_39197,N_27373,N_24909);
nand U39198 (N_39198,N_25904,N_20091);
nand U39199 (N_39199,N_26867,N_23636);
and U39200 (N_39200,N_29123,N_29971);
nand U39201 (N_39201,N_24298,N_21204);
nor U39202 (N_39202,N_25869,N_25219);
or U39203 (N_39203,N_29177,N_23062);
nand U39204 (N_39204,N_22167,N_27356);
and U39205 (N_39205,N_27714,N_29342);
xnor U39206 (N_39206,N_22839,N_24954);
nor U39207 (N_39207,N_29398,N_27935);
xnor U39208 (N_39208,N_28899,N_22483);
and U39209 (N_39209,N_20467,N_20899);
nor U39210 (N_39210,N_28644,N_22676);
nor U39211 (N_39211,N_28408,N_28335);
xnor U39212 (N_39212,N_25092,N_28638);
nor U39213 (N_39213,N_24347,N_27453);
nand U39214 (N_39214,N_25345,N_20943);
or U39215 (N_39215,N_20244,N_29670);
nand U39216 (N_39216,N_20650,N_25434);
nand U39217 (N_39217,N_22334,N_24506);
or U39218 (N_39218,N_28255,N_27465);
nand U39219 (N_39219,N_20673,N_25012);
nor U39220 (N_39220,N_27655,N_25665);
nand U39221 (N_39221,N_25473,N_28747);
nor U39222 (N_39222,N_20557,N_23798);
xor U39223 (N_39223,N_20623,N_21427);
xor U39224 (N_39224,N_23187,N_20667);
and U39225 (N_39225,N_29457,N_26991);
nand U39226 (N_39226,N_22410,N_28563);
and U39227 (N_39227,N_22893,N_23996);
nand U39228 (N_39228,N_28482,N_22702);
xnor U39229 (N_39229,N_20965,N_28183);
nand U39230 (N_39230,N_22095,N_23369);
or U39231 (N_39231,N_20360,N_22251);
and U39232 (N_39232,N_29633,N_28455);
or U39233 (N_39233,N_28278,N_26379);
nor U39234 (N_39234,N_21666,N_22414);
xor U39235 (N_39235,N_21643,N_23236);
xnor U39236 (N_39236,N_20254,N_20325);
xnor U39237 (N_39237,N_27963,N_28081);
nand U39238 (N_39238,N_22662,N_20622);
nor U39239 (N_39239,N_24349,N_20592);
or U39240 (N_39240,N_22800,N_20140);
nor U39241 (N_39241,N_25756,N_23897);
xor U39242 (N_39242,N_29300,N_23230);
xor U39243 (N_39243,N_21154,N_20190);
xor U39244 (N_39244,N_25909,N_23082);
and U39245 (N_39245,N_25554,N_25379);
nor U39246 (N_39246,N_22038,N_29883);
or U39247 (N_39247,N_25082,N_25182);
or U39248 (N_39248,N_23432,N_28736);
nand U39249 (N_39249,N_25590,N_24262);
nand U39250 (N_39250,N_22506,N_26618);
or U39251 (N_39251,N_24269,N_28829);
nor U39252 (N_39252,N_23771,N_29139);
or U39253 (N_39253,N_22013,N_22795);
and U39254 (N_39254,N_27486,N_23139);
xnor U39255 (N_39255,N_22395,N_20160);
nand U39256 (N_39256,N_26059,N_27523);
xnor U39257 (N_39257,N_28002,N_27532);
nor U39258 (N_39258,N_24739,N_24084);
or U39259 (N_39259,N_26047,N_26345);
nand U39260 (N_39260,N_26405,N_20953);
xnor U39261 (N_39261,N_27539,N_21293);
nand U39262 (N_39262,N_26867,N_23938);
nor U39263 (N_39263,N_28584,N_24063);
or U39264 (N_39264,N_27747,N_25174);
and U39265 (N_39265,N_24874,N_26970);
xnor U39266 (N_39266,N_24705,N_23633);
and U39267 (N_39267,N_28370,N_23076);
nand U39268 (N_39268,N_20355,N_22603);
xnor U39269 (N_39269,N_29225,N_20818);
or U39270 (N_39270,N_23067,N_23940);
xor U39271 (N_39271,N_26188,N_27834);
xnor U39272 (N_39272,N_27261,N_25363);
or U39273 (N_39273,N_24306,N_24495);
and U39274 (N_39274,N_24635,N_21033);
nand U39275 (N_39275,N_27866,N_29976);
or U39276 (N_39276,N_28528,N_27866);
nor U39277 (N_39277,N_21617,N_25052);
nand U39278 (N_39278,N_21517,N_20135);
or U39279 (N_39279,N_29103,N_21516);
xnor U39280 (N_39280,N_23604,N_21582);
or U39281 (N_39281,N_28410,N_24874);
nor U39282 (N_39282,N_21450,N_26851);
nor U39283 (N_39283,N_23819,N_29550);
nor U39284 (N_39284,N_22893,N_26638);
and U39285 (N_39285,N_24237,N_25520);
xor U39286 (N_39286,N_26456,N_28860);
xor U39287 (N_39287,N_24941,N_22016);
nor U39288 (N_39288,N_29087,N_28105);
and U39289 (N_39289,N_25987,N_28590);
and U39290 (N_39290,N_21025,N_25867);
or U39291 (N_39291,N_20296,N_21870);
nand U39292 (N_39292,N_23089,N_22968);
nor U39293 (N_39293,N_21818,N_24420);
and U39294 (N_39294,N_29553,N_23952);
nand U39295 (N_39295,N_23719,N_23832);
nand U39296 (N_39296,N_27465,N_26140);
nand U39297 (N_39297,N_21231,N_23292);
and U39298 (N_39298,N_23811,N_25504);
nor U39299 (N_39299,N_20255,N_22578);
xor U39300 (N_39300,N_20653,N_29527);
or U39301 (N_39301,N_23721,N_20286);
nand U39302 (N_39302,N_28710,N_27954);
nand U39303 (N_39303,N_20057,N_22154);
nand U39304 (N_39304,N_27935,N_21446);
nand U39305 (N_39305,N_28852,N_26783);
nand U39306 (N_39306,N_22590,N_27930);
or U39307 (N_39307,N_29209,N_24106);
and U39308 (N_39308,N_25900,N_20624);
nand U39309 (N_39309,N_23016,N_20840);
nor U39310 (N_39310,N_25317,N_23901);
or U39311 (N_39311,N_25637,N_27588);
nor U39312 (N_39312,N_27787,N_23995);
xnor U39313 (N_39313,N_29775,N_29840);
xor U39314 (N_39314,N_23261,N_27445);
xnor U39315 (N_39315,N_21121,N_29434);
or U39316 (N_39316,N_20995,N_25751);
or U39317 (N_39317,N_21401,N_29951);
and U39318 (N_39318,N_23644,N_23671);
or U39319 (N_39319,N_22450,N_20466);
nand U39320 (N_39320,N_21950,N_29538);
or U39321 (N_39321,N_27231,N_27980);
nor U39322 (N_39322,N_22834,N_29330);
or U39323 (N_39323,N_28806,N_26891);
nand U39324 (N_39324,N_20923,N_20939);
nor U39325 (N_39325,N_24089,N_20815);
nor U39326 (N_39326,N_28970,N_20253);
xnor U39327 (N_39327,N_28605,N_25542);
or U39328 (N_39328,N_22230,N_29708);
and U39329 (N_39329,N_27380,N_29612);
nor U39330 (N_39330,N_27811,N_28891);
nand U39331 (N_39331,N_27579,N_21888);
nand U39332 (N_39332,N_24792,N_26547);
xor U39333 (N_39333,N_27526,N_28612);
or U39334 (N_39334,N_25921,N_24559);
and U39335 (N_39335,N_28757,N_23368);
nand U39336 (N_39336,N_21838,N_27516);
nor U39337 (N_39337,N_23696,N_24808);
xor U39338 (N_39338,N_26273,N_28574);
and U39339 (N_39339,N_24922,N_21436);
xnor U39340 (N_39340,N_21359,N_21874);
nor U39341 (N_39341,N_28332,N_25471);
or U39342 (N_39342,N_27424,N_21405);
and U39343 (N_39343,N_21669,N_27068);
nand U39344 (N_39344,N_21658,N_28991);
or U39345 (N_39345,N_25533,N_21124);
and U39346 (N_39346,N_23192,N_22430);
xnor U39347 (N_39347,N_24790,N_20215);
nand U39348 (N_39348,N_23659,N_29842);
xnor U39349 (N_39349,N_26706,N_25797);
and U39350 (N_39350,N_28331,N_24190);
nor U39351 (N_39351,N_22863,N_26467);
xnor U39352 (N_39352,N_22944,N_27442);
or U39353 (N_39353,N_28806,N_23002);
and U39354 (N_39354,N_28861,N_21771);
nand U39355 (N_39355,N_25331,N_25148);
nor U39356 (N_39356,N_28467,N_20136);
or U39357 (N_39357,N_20510,N_23988);
or U39358 (N_39358,N_28014,N_27785);
nor U39359 (N_39359,N_21584,N_22619);
nand U39360 (N_39360,N_25110,N_27339);
or U39361 (N_39361,N_23772,N_24830);
or U39362 (N_39362,N_28594,N_28619);
or U39363 (N_39363,N_20133,N_20695);
nand U39364 (N_39364,N_24014,N_28910);
xnor U39365 (N_39365,N_25855,N_23652);
xor U39366 (N_39366,N_25415,N_23101);
nor U39367 (N_39367,N_29452,N_27305);
nor U39368 (N_39368,N_25468,N_26645);
xor U39369 (N_39369,N_29612,N_21874);
nor U39370 (N_39370,N_20569,N_27646);
nor U39371 (N_39371,N_26320,N_24406);
xor U39372 (N_39372,N_20124,N_23015);
nor U39373 (N_39373,N_21656,N_23382);
nor U39374 (N_39374,N_28422,N_20180);
nor U39375 (N_39375,N_29827,N_27346);
or U39376 (N_39376,N_22105,N_27094);
and U39377 (N_39377,N_29181,N_22912);
xnor U39378 (N_39378,N_28922,N_29804);
nand U39379 (N_39379,N_20959,N_28664);
nor U39380 (N_39380,N_21632,N_27087);
nor U39381 (N_39381,N_29469,N_24319);
nor U39382 (N_39382,N_26243,N_26407);
or U39383 (N_39383,N_28552,N_21781);
xnor U39384 (N_39384,N_21558,N_25337);
nor U39385 (N_39385,N_29021,N_21968);
nor U39386 (N_39386,N_21730,N_22972);
nand U39387 (N_39387,N_21046,N_24356);
or U39388 (N_39388,N_22211,N_21350);
nand U39389 (N_39389,N_28958,N_29350);
nand U39390 (N_39390,N_23574,N_27163);
and U39391 (N_39391,N_23061,N_21849);
nand U39392 (N_39392,N_27875,N_29582);
and U39393 (N_39393,N_24154,N_26149);
or U39394 (N_39394,N_27624,N_22487);
nor U39395 (N_39395,N_26406,N_20658);
or U39396 (N_39396,N_20270,N_21841);
nor U39397 (N_39397,N_28519,N_23411);
or U39398 (N_39398,N_25240,N_20710);
or U39399 (N_39399,N_27952,N_27651);
and U39400 (N_39400,N_21115,N_28765);
or U39401 (N_39401,N_23787,N_27802);
nand U39402 (N_39402,N_21102,N_23454);
and U39403 (N_39403,N_20025,N_22343);
xor U39404 (N_39404,N_23105,N_24103);
or U39405 (N_39405,N_22940,N_29108);
nor U39406 (N_39406,N_22290,N_23450);
or U39407 (N_39407,N_21355,N_20015);
nor U39408 (N_39408,N_23136,N_20385);
and U39409 (N_39409,N_23046,N_22191);
xnor U39410 (N_39410,N_22980,N_22599);
nor U39411 (N_39411,N_25926,N_28398);
or U39412 (N_39412,N_26200,N_21873);
nor U39413 (N_39413,N_21281,N_22615);
or U39414 (N_39414,N_25289,N_20668);
nor U39415 (N_39415,N_22978,N_22413);
nand U39416 (N_39416,N_28903,N_28464);
xor U39417 (N_39417,N_27996,N_27802);
xor U39418 (N_39418,N_28270,N_21756);
nor U39419 (N_39419,N_21882,N_20236);
or U39420 (N_39420,N_26884,N_20139);
or U39421 (N_39421,N_26135,N_21718);
xor U39422 (N_39422,N_25238,N_24838);
nand U39423 (N_39423,N_23173,N_29408);
nand U39424 (N_39424,N_27597,N_28546);
nand U39425 (N_39425,N_21287,N_22025);
nand U39426 (N_39426,N_25479,N_23250);
nor U39427 (N_39427,N_29668,N_21995);
or U39428 (N_39428,N_25143,N_29262);
and U39429 (N_39429,N_20622,N_27659);
xnor U39430 (N_39430,N_24885,N_23326);
xor U39431 (N_39431,N_23649,N_27083);
nand U39432 (N_39432,N_28238,N_25385);
nor U39433 (N_39433,N_29727,N_24359);
or U39434 (N_39434,N_20161,N_28348);
or U39435 (N_39435,N_20125,N_26359);
nor U39436 (N_39436,N_28052,N_28989);
or U39437 (N_39437,N_27516,N_26600);
and U39438 (N_39438,N_24560,N_25999);
and U39439 (N_39439,N_22579,N_22935);
nor U39440 (N_39440,N_29372,N_27640);
or U39441 (N_39441,N_21395,N_27671);
and U39442 (N_39442,N_20481,N_23167);
nand U39443 (N_39443,N_20186,N_21886);
xnor U39444 (N_39444,N_22431,N_25910);
nand U39445 (N_39445,N_29670,N_29767);
and U39446 (N_39446,N_24999,N_20685);
nor U39447 (N_39447,N_29617,N_25430);
nor U39448 (N_39448,N_25313,N_25636);
and U39449 (N_39449,N_24388,N_25075);
or U39450 (N_39450,N_27587,N_24677);
xor U39451 (N_39451,N_22643,N_26148);
xnor U39452 (N_39452,N_28310,N_28360);
and U39453 (N_39453,N_29226,N_20092);
xnor U39454 (N_39454,N_27414,N_23447);
or U39455 (N_39455,N_20629,N_23516);
nand U39456 (N_39456,N_28122,N_22817);
xnor U39457 (N_39457,N_29962,N_25904);
nor U39458 (N_39458,N_25798,N_29486);
or U39459 (N_39459,N_27558,N_26088);
xor U39460 (N_39460,N_27123,N_23297);
nor U39461 (N_39461,N_24146,N_29163);
nand U39462 (N_39462,N_22238,N_29662);
or U39463 (N_39463,N_26736,N_25143);
or U39464 (N_39464,N_26245,N_27688);
or U39465 (N_39465,N_21010,N_23579);
nor U39466 (N_39466,N_26450,N_26696);
nand U39467 (N_39467,N_20051,N_20647);
or U39468 (N_39468,N_26004,N_26558);
or U39469 (N_39469,N_24571,N_20073);
and U39470 (N_39470,N_24972,N_28101);
or U39471 (N_39471,N_24666,N_29506);
nand U39472 (N_39472,N_29228,N_20517);
nor U39473 (N_39473,N_23497,N_28145);
or U39474 (N_39474,N_29362,N_23300);
or U39475 (N_39475,N_22157,N_20484);
and U39476 (N_39476,N_22187,N_27637);
nand U39477 (N_39477,N_24105,N_27498);
and U39478 (N_39478,N_21002,N_20990);
and U39479 (N_39479,N_20807,N_23000);
xor U39480 (N_39480,N_26756,N_28111);
xnor U39481 (N_39481,N_25705,N_27969);
nor U39482 (N_39482,N_23290,N_29756);
and U39483 (N_39483,N_24522,N_27596);
or U39484 (N_39484,N_20725,N_29537);
nor U39485 (N_39485,N_23141,N_24501);
xor U39486 (N_39486,N_28233,N_22428);
and U39487 (N_39487,N_24202,N_22930);
and U39488 (N_39488,N_22146,N_29894);
nand U39489 (N_39489,N_27065,N_24554);
nand U39490 (N_39490,N_20736,N_28750);
or U39491 (N_39491,N_22962,N_20462);
nor U39492 (N_39492,N_29132,N_28997);
xnor U39493 (N_39493,N_20392,N_20266);
and U39494 (N_39494,N_24703,N_21531);
nand U39495 (N_39495,N_20502,N_20259);
and U39496 (N_39496,N_25051,N_23839);
nor U39497 (N_39497,N_29087,N_25151);
and U39498 (N_39498,N_25018,N_23833);
and U39499 (N_39499,N_20360,N_21076);
nand U39500 (N_39500,N_20910,N_29030);
nor U39501 (N_39501,N_21061,N_20134);
or U39502 (N_39502,N_21776,N_28444);
nor U39503 (N_39503,N_29378,N_28180);
nand U39504 (N_39504,N_21303,N_23563);
or U39505 (N_39505,N_25574,N_26189);
xnor U39506 (N_39506,N_25485,N_23841);
xnor U39507 (N_39507,N_28710,N_26461);
nand U39508 (N_39508,N_29206,N_21331);
xor U39509 (N_39509,N_24526,N_24866);
nor U39510 (N_39510,N_29671,N_25621);
nand U39511 (N_39511,N_20883,N_22077);
nand U39512 (N_39512,N_29563,N_28107);
nand U39513 (N_39513,N_29246,N_20385);
and U39514 (N_39514,N_23833,N_26269);
xnor U39515 (N_39515,N_26222,N_24360);
or U39516 (N_39516,N_27073,N_23696);
and U39517 (N_39517,N_22859,N_21847);
and U39518 (N_39518,N_20438,N_25889);
nand U39519 (N_39519,N_20843,N_24714);
and U39520 (N_39520,N_26813,N_24210);
or U39521 (N_39521,N_25928,N_25317);
xor U39522 (N_39522,N_24009,N_20236);
nor U39523 (N_39523,N_20830,N_26862);
nand U39524 (N_39524,N_25869,N_29745);
nor U39525 (N_39525,N_24202,N_23593);
or U39526 (N_39526,N_21553,N_22798);
nor U39527 (N_39527,N_28252,N_26795);
xnor U39528 (N_39528,N_22172,N_21653);
nand U39529 (N_39529,N_26078,N_28872);
and U39530 (N_39530,N_20674,N_25641);
and U39531 (N_39531,N_28520,N_21632);
xnor U39532 (N_39532,N_26432,N_26392);
and U39533 (N_39533,N_26534,N_20271);
nor U39534 (N_39534,N_25369,N_23912);
xnor U39535 (N_39535,N_28294,N_26084);
nor U39536 (N_39536,N_22043,N_27495);
nand U39537 (N_39537,N_27479,N_22724);
nand U39538 (N_39538,N_27828,N_21306);
xor U39539 (N_39539,N_27598,N_21837);
and U39540 (N_39540,N_24001,N_23854);
xor U39541 (N_39541,N_26618,N_23782);
nor U39542 (N_39542,N_21664,N_22646);
nand U39543 (N_39543,N_20908,N_24904);
or U39544 (N_39544,N_27759,N_28512);
nor U39545 (N_39545,N_27746,N_29752);
and U39546 (N_39546,N_27099,N_25137);
or U39547 (N_39547,N_24445,N_27691);
nand U39548 (N_39548,N_28727,N_28520);
xnor U39549 (N_39549,N_28361,N_28279);
nor U39550 (N_39550,N_23897,N_28137);
and U39551 (N_39551,N_23045,N_20570);
nand U39552 (N_39552,N_29755,N_25437);
and U39553 (N_39553,N_20379,N_29363);
and U39554 (N_39554,N_20677,N_28934);
or U39555 (N_39555,N_24494,N_26195);
and U39556 (N_39556,N_23763,N_22661);
nand U39557 (N_39557,N_21615,N_21686);
or U39558 (N_39558,N_22640,N_23617);
xnor U39559 (N_39559,N_23798,N_25453);
and U39560 (N_39560,N_21266,N_23973);
nor U39561 (N_39561,N_25530,N_21492);
or U39562 (N_39562,N_22954,N_29984);
and U39563 (N_39563,N_24156,N_21673);
nand U39564 (N_39564,N_21998,N_24392);
or U39565 (N_39565,N_20849,N_23021);
or U39566 (N_39566,N_21992,N_25581);
nand U39567 (N_39567,N_29297,N_23757);
or U39568 (N_39568,N_23644,N_25887);
nand U39569 (N_39569,N_23260,N_22028);
nand U39570 (N_39570,N_24886,N_25232);
nor U39571 (N_39571,N_22587,N_24787);
xnor U39572 (N_39572,N_28393,N_23310);
xor U39573 (N_39573,N_20450,N_26299);
and U39574 (N_39574,N_25329,N_29918);
and U39575 (N_39575,N_23008,N_27147);
or U39576 (N_39576,N_29056,N_29249);
xor U39577 (N_39577,N_24947,N_27672);
nand U39578 (N_39578,N_21207,N_20726);
xnor U39579 (N_39579,N_23178,N_23002);
nor U39580 (N_39580,N_24555,N_27919);
xnor U39581 (N_39581,N_24108,N_23950);
nand U39582 (N_39582,N_22970,N_29182);
nor U39583 (N_39583,N_22869,N_29817);
nand U39584 (N_39584,N_23039,N_29023);
and U39585 (N_39585,N_27062,N_28144);
xnor U39586 (N_39586,N_26158,N_29356);
or U39587 (N_39587,N_24235,N_28507);
nand U39588 (N_39588,N_27158,N_27539);
nor U39589 (N_39589,N_26220,N_23818);
nor U39590 (N_39590,N_25554,N_23067);
nor U39591 (N_39591,N_20156,N_25922);
nor U39592 (N_39592,N_26783,N_21107);
or U39593 (N_39593,N_21932,N_27644);
or U39594 (N_39594,N_28060,N_20342);
nor U39595 (N_39595,N_27125,N_23003);
or U39596 (N_39596,N_24744,N_28313);
and U39597 (N_39597,N_23628,N_20167);
nand U39598 (N_39598,N_20893,N_26272);
nand U39599 (N_39599,N_26579,N_27409);
and U39600 (N_39600,N_25101,N_22637);
xnor U39601 (N_39601,N_27117,N_25878);
xnor U39602 (N_39602,N_25878,N_21788);
nand U39603 (N_39603,N_23610,N_22712);
or U39604 (N_39604,N_24360,N_23762);
and U39605 (N_39605,N_27805,N_21275);
or U39606 (N_39606,N_29624,N_25267);
and U39607 (N_39607,N_24852,N_29691);
nor U39608 (N_39608,N_26980,N_28913);
and U39609 (N_39609,N_22076,N_25130);
or U39610 (N_39610,N_20999,N_29603);
or U39611 (N_39611,N_21051,N_26291);
nor U39612 (N_39612,N_23600,N_29158);
nor U39613 (N_39613,N_23378,N_28792);
nor U39614 (N_39614,N_22345,N_27030);
and U39615 (N_39615,N_28710,N_25674);
or U39616 (N_39616,N_25970,N_24787);
nand U39617 (N_39617,N_24467,N_26314);
xor U39618 (N_39618,N_29271,N_21313);
and U39619 (N_39619,N_22035,N_25810);
nand U39620 (N_39620,N_20597,N_27163);
nor U39621 (N_39621,N_26698,N_26988);
nor U39622 (N_39622,N_22017,N_25255);
nor U39623 (N_39623,N_23380,N_29824);
xor U39624 (N_39624,N_20723,N_25432);
or U39625 (N_39625,N_20650,N_28541);
nor U39626 (N_39626,N_23276,N_21401);
nor U39627 (N_39627,N_23104,N_23780);
and U39628 (N_39628,N_21707,N_24438);
nand U39629 (N_39629,N_27749,N_21956);
xor U39630 (N_39630,N_24391,N_21113);
xor U39631 (N_39631,N_29238,N_28879);
or U39632 (N_39632,N_29825,N_20070);
or U39633 (N_39633,N_28291,N_20982);
xnor U39634 (N_39634,N_25899,N_24727);
or U39635 (N_39635,N_28250,N_26426);
or U39636 (N_39636,N_23676,N_28039);
nor U39637 (N_39637,N_22630,N_24131);
and U39638 (N_39638,N_26352,N_27304);
nand U39639 (N_39639,N_24135,N_25426);
or U39640 (N_39640,N_25637,N_29514);
xnor U39641 (N_39641,N_26951,N_25662);
nand U39642 (N_39642,N_26936,N_29130);
and U39643 (N_39643,N_24578,N_25017);
xor U39644 (N_39644,N_20082,N_21852);
nor U39645 (N_39645,N_24971,N_27795);
nor U39646 (N_39646,N_24273,N_23014);
and U39647 (N_39647,N_28352,N_23048);
nor U39648 (N_39648,N_21915,N_27940);
xnor U39649 (N_39649,N_28901,N_26143);
or U39650 (N_39650,N_26643,N_29714);
nand U39651 (N_39651,N_26579,N_29740);
nor U39652 (N_39652,N_20384,N_26891);
xor U39653 (N_39653,N_27437,N_21210);
and U39654 (N_39654,N_22727,N_22191);
nand U39655 (N_39655,N_22745,N_26542);
and U39656 (N_39656,N_27274,N_28389);
and U39657 (N_39657,N_21115,N_28666);
and U39658 (N_39658,N_20630,N_26832);
xnor U39659 (N_39659,N_26597,N_27287);
nand U39660 (N_39660,N_21622,N_20561);
nor U39661 (N_39661,N_25728,N_20450);
nor U39662 (N_39662,N_29159,N_22531);
xnor U39663 (N_39663,N_24843,N_22634);
xor U39664 (N_39664,N_22846,N_20962);
and U39665 (N_39665,N_23359,N_29970);
nand U39666 (N_39666,N_29366,N_24944);
nand U39667 (N_39667,N_27928,N_24357);
nand U39668 (N_39668,N_20673,N_22336);
nor U39669 (N_39669,N_24397,N_27359);
nor U39670 (N_39670,N_22594,N_23531);
nor U39671 (N_39671,N_21142,N_25644);
or U39672 (N_39672,N_26172,N_21539);
and U39673 (N_39673,N_29342,N_25477);
or U39674 (N_39674,N_21855,N_20346);
xor U39675 (N_39675,N_24225,N_24289);
nand U39676 (N_39676,N_24064,N_21064);
nand U39677 (N_39677,N_29187,N_25762);
nand U39678 (N_39678,N_23860,N_29634);
xnor U39679 (N_39679,N_23438,N_28031);
xor U39680 (N_39680,N_20941,N_26998);
or U39681 (N_39681,N_23248,N_28013);
xnor U39682 (N_39682,N_25976,N_20399);
or U39683 (N_39683,N_25247,N_20307);
nor U39684 (N_39684,N_27743,N_29571);
nand U39685 (N_39685,N_24837,N_20702);
nor U39686 (N_39686,N_25150,N_28828);
xnor U39687 (N_39687,N_27285,N_22510);
or U39688 (N_39688,N_22614,N_20665);
nand U39689 (N_39689,N_22497,N_23893);
or U39690 (N_39690,N_22899,N_26040);
nor U39691 (N_39691,N_20388,N_24680);
and U39692 (N_39692,N_21886,N_28371);
xnor U39693 (N_39693,N_29578,N_21095);
nand U39694 (N_39694,N_26960,N_24693);
or U39695 (N_39695,N_26527,N_22377);
or U39696 (N_39696,N_23784,N_29519);
nor U39697 (N_39697,N_23362,N_20104);
nor U39698 (N_39698,N_29339,N_29455);
and U39699 (N_39699,N_26819,N_25255);
nor U39700 (N_39700,N_29236,N_22125);
or U39701 (N_39701,N_24743,N_25331);
nand U39702 (N_39702,N_28768,N_27050);
nand U39703 (N_39703,N_28299,N_24629);
nand U39704 (N_39704,N_29950,N_29280);
and U39705 (N_39705,N_29282,N_29379);
or U39706 (N_39706,N_26768,N_22788);
nand U39707 (N_39707,N_26317,N_23898);
nand U39708 (N_39708,N_23680,N_26916);
or U39709 (N_39709,N_20672,N_20608);
xor U39710 (N_39710,N_22542,N_25296);
nand U39711 (N_39711,N_24868,N_28111);
xor U39712 (N_39712,N_22415,N_20736);
nand U39713 (N_39713,N_23352,N_22163);
and U39714 (N_39714,N_24993,N_22592);
nand U39715 (N_39715,N_26101,N_26907);
and U39716 (N_39716,N_20226,N_26601);
nor U39717 (N_39717,N_21333,N_29496);
or U39718 (N_39718,N_20258,N_27646);
nand U39719 (N_39719,N_26654,N_22134);
xor U39720 (N_39720,N_23884,N_28651);
xor U39721 (N_39721,N_28792,N_23511);
nor U39722 (N_39722,N_29944,N_20138);
or U39723 (N_39723,N_28683,N_23059);
nor U39724 (N_39724,N_22400,N_25210);
nor U39725 (N_39725,N_23667,N_24543);
xnor U39726 (N_39726,N_27140,N_21449);
nand U39727 (N_39727,N_20850,N_27632);
or U39728 (N_39728,N_20711,N_27784);
and U39729 (N_39729,N_20945,N_20850);
nor U39730 (N_39730,N_20987,N_26535);
nor U39731 (N_39731,N_27302,N_29843);
nor U39732 (N_39732,N_20346,N_20062);
nor U39733 (N_39733,N_23780,N_23003);
and U39734 (N_39734,N_22965,N_22450);
nand U39735 (N_39735,N_25661,N_20904);
and U39736 (N_39736,N_26496,N_22241);
or U39737 (N_39737,N_28039,N_27114);
or U39738 (N_39738,N_27824,N_29854);
or U39739 (N_39739,N_24817,N_21264);
and U39740 (N_39740,N_24501,N_27879);
nand U39741 (N_39741,N_24882,N_21632);
and U39742 (N_39742,N_22890,N_26605);
or U39743 (N_39743,N_21020,N_27793);
xor U39744 (N_39744,N_26241,N_25903);
xor U39745 (N_39745,N_20294,N_21138);
xnor U39746 (N_39746,N_20624,N_22184);
and U39747 (N_39747,N_28464,N_21441);
and U39748 (N_39748,N_22880,N_20140);
nand U39749 (N_39749,N_24932,N_21787);
nand U39750 (N_39750,N_20746,N_29032);
or U39751 (N_39751,N_29249,N_20682);
and U39752 (N_39752,N_29364,N_26850);
xnor U39753 (N_39753,N_28782,N_27217);
xor U39754 (N_39754,N_27049,N_27533);
or U39755 (N_39755,N_27060,N_29730);
xor U39756 (N_39756,N_21644,N_23818);
and U39757 (N_39757,N_20924,N_23119);
xor U39758 (N_39758,N_22295,N_22424);
xor U39759 (N_39759,N_25554,N_26521);
nor U39760 (N_39760,N_23841,N_20946);
xnor U39761 (N_39761,N_23279,N_27100);
and U39762 (N_39762,N_25515,N_28071);
nor U39763 (N_39763,N_24152,N_25309);
and U39764 (N_39764,N_25803,N_21500);
or U39765 (N_39765,N_23903,N_24520);
or U39766 (N_39766,N_26824,N_24991);
and U39767 (N_39767,N_26446,N_26676);
or U39768 (N_39768,N_27555,N_20435);
nand U39769 (N_39769,N_26704,N_27051);
xor U39770 (N_39770,N_21701,N_26056);
nand U39771 (N_39771,N_22434,N_24342);
nor U39772 (N_39772,N_22829,N_25747);
xnor U39773 (N_39773,N_26644,N_27530);
and U39774 (N_39774,N_23840,N_27873);
nor U39775 (N_39775,N_20358,N_26199);
xor U39776 (N_39776,N_28350,N_21276);
xor U39777 (N_39777,N_20580,N_21469);
and U39778 (N_39778,N_28922,N_27634);
nor U39779 (N_39779,N_28579,N_26898);
and U39780 (N_39780,N_28559,N_29772);
nor U39781 (N_39781,N_25287,N_21387);
xor U39782 (N_39782,N_20133,N_23985);
nor U39783 (N_39783,N_20403,N_27577);
or U39784 (N_39784,N_24636,N_22925);
nand U39785 (N_39785,N_23265,N_26381);
or U39786 (N_39786,N_22169,N_25704);
and U39787 (N_39787,N_27139,N_27785);
nand U39788 (N_39788,N_22033,N_26251);
or U39789 (N_39789,N_22481,N_23072);
and U39790 (N_39790,N_20091,N_22755);
nor U39791 (N_39791,N_25876,N_20339);
and U39792 (N_39792,N_29000,N_28202);
nand U39793 (N_39793,N_22211,N_25609);
and U39794 (N_39794,N_23426,N_27861);
nor U39795 (N_39795,N_25043,N_27658);
xor U39796 (N_39796,N_21085,N_29662);
nor U39797 (N_39797,N_29617,N_23871);
and U39798 (N_39798,N_24389,N_24656);
and U39799 (N_39799,N_28309,N_27579);
nor U39800 (N_39800,N_27998,N_21692);
xor U39801 (N_39801,N_25204,N_28704);
nand U39802 (N_39802,N_28163,N_22528);
and U39803 (N_39803,N_22018,N_29175);
or U39804 (N_39804,N_27391,N_23790);
and U39805 (N_39805,N_24057,N_28958);
xnor U39806 (N_39806,N_20032,N_24317);
nor U39807 (N_39807,N_26105,N_24431);
or U39808 (N_39808,N_25336,N_29158);
and U39809 (N_39809,N_24409,N_21250);
nand U39810 (N_39810,N_25049,N_22934);
nand U39811 (N_39811,N_27836,N_21255);
xnor U39812 (N_39812,N_20121,N_27341);
xor U39813 (N_39813,N_29391,N_23983);
or U39814 (N_39814,N_22081,N_23132);
xnor U39815 (N_39815,N_24634,N_20355);
and U39816 (N_39816,N_28467,N_26332);
nor U39817 (N_39817,N_26252,N_21023);
nor U39818 (N_39818,N_28033,N_26337);
nor U39819 (N_39819,N_29261,N_24345);
nand U39820 (N_39820,N_29172,N_29277);
or U39821 (N_39821,N_22723,N_29313);
nor U39822 (N_39822,N_28568,N_20628);
xor U39823 (N_39823,N_22612,N_29813);
xnor U39824 (N_39824,N_29907,N_20917);
nand U39825 (N_39825,N_22615,N_28546);
nor U39826 (N_39826,N_20078,N_20027);
or U39827 (N_39827,N_20564,N_22533);
nor U39828 (N_39828,N_21686,N_20502);
or U39829 (N_39829,N_26340,N_20161);
and U39830 (N_39830,N_20107,N_23200);
and U39831 (N_39831,N_22095,N_24523);
xnor U39832 (N_39832,N_27912,N_29561);
xnor U39833 (N_39833,N_22874,N_25108);
or U39834 (N_39834,N_29940,N_25100);
or U39835 (N_39835,N_21230,N_24773);
and U39836 (N_39836,N_26264,N_23491);
xnor U39837 (N_39837,N_28616,N_21472);
and U39838 (N_39838,N_27356,N_23968);
xnor U39839 (N_39839,N_20088,N_27409);
and U39840 (N_39840,N_26339,N_22501);
or U39841 (N_39841,N_28914,N_29559);
xnor U39842 (N_39842,N_20909,N_24749);
xnor U39843 (N_39843,N_24321,N_24355);
or U39844 (N_39844,N_27985,N_24299);
or U39845 (N_39845,N_25063,N_24666);
nand U39846 (N_39846,N_29014,N_23637);
or U39847 (N_39847,N_20915,N_21328);
nor U39848 (N_39848,N_26622,N_21885);
nand U39849 (N_39849,N_28398,N_28232);
nand U39850 (N_39850,N_26533,N_27623);
or U39851 (N_39851,N_25032,N_27591);
nor U39852 (N_39852,N_26559,N_21193);
xor U39853 (N_39853,N_23486,N_22085);
xor U39854 (N_39854,N_25139,N_20315);
or U39855 (N_39855,N_23729,N_28322);
xor U39856 (N_39856,N_26471,N_25044);
nor U39857 (N_39857,N_27557,N_26423);
xor U39858 (N_39858,N_27371,N_27422);
nor U39859 (N_39859,N_27925,N_25394);
nor U39860 (N_39860,N_23051,N_20114);
and U39861 (N_39861,N_22154,N_27442);
nor U39862 (N_39862,N_25323,N_27945);
and U39863 (N_39863,N_25843,N_25044);
or U39864 (N_39864,N_29839,N_20804);
nand U39865 (N_39865,N_24004,N_24124);
and U39866 (N_39866,N_20801,N_25758);
nand U39867 (N_39867,N_24056,N_26736);
nor U39868 (N_39868,N_20101,N_22961);
xnor U39869 (N_39869,N_21501,N_28311);
and U39870 (N_39870,N_20649,N_22901);
or U39871 (N_39871,N_25782,N_27342);
xor U39872 (N_39872,N_20814,N_22260);
and U39873 (N_39873,N_28375,N_22107);
and U39874 (N_39874,N_26560,N_21077);
or U39875 (N_39875,N_25963,N_20803);
nor U39876 (N_39876,N_29409,N_22384);
and U39877 (N_39877,N_26624,N_22554);
and U39878 (N_39878,N_22927,N_24772);
xor U39879 (N_39879,N_25880,N_25585);
nand U39880 (N_39880,N_25396,N_29164);
or U39881 (N_39881,N_27957,N_20882);
and U39882 (N_39882,N_25692,N_29277);
or U39883 (N_39883,N_28778,N_25281);
xnor U39884 (N_39884,N_27592,N_22274);
nor U39885 (N_39885,N_25623,N_23964);
or U39886 (N_39886,N_21941,N_22637);
and U39887 (N_39887,N_22675,N_25771);
and U39888 (N_39888,N_22516,N_25221);
and U39889 (N_39889,N_29516,N_26422);
nor U39890 (N_39890,N_20374,N_27850);
or U39891 (N_39891,N_29699,N_22916);
nand U39892 (N_39892,N_22667,N_28229);
nand U39893 (N_39893,N_22529,N_26906);
xnor U39894 (N_39894,N_27337,N_20494);
xor U39895 (N_39895,N_20702,N_26260);
nand U39896 (N_39896,N_25931,N_27616);
or U39897 (N_39897,N_21183,N_23172);
and U39898 (N_39898,N_29885,N_23828);
nand U39899 (N_39899,N_23776,N_24554);
xnor U39900 (N_39900,N_24271,N_23336);
nor U39901 (N_39901,N_25262,N_24154);
nand U39902 (N_39902,N_24838,N_23896);
nand U39903 (N_39903,N_26612,N_27816);
nand U39904 (N_39904,N_26030,N_28707);
and U39905 (N_39905,N_20604,N_25103);
nor U39906 (N_39906,N_26322,N_24450);
nand U39907 (N_39907,N_20625,N_20747);
nand U39908 (N_39908,N_26075,N_28133);
xor U39909 (N_39909,N_24263,N_20420);
nor U39910 (N_39910,N_23770,N_20214);
nand U39911 (N_39911,N_23017,N_26081);
nor U39912 (N_39912,N_20347,N_25168);
or U39913 (N_39913,N_27668,N_29215);
and U39914 (N_39914,N_25217,N_20543);
xnor U39915 (N_39915,N_25487,N_25146);
or U39916 (N_39916,N_24045,N_20777);
and U39917 (N_39917,N_21175,N_29529);
xor U39918 (N_39918,N_21339,N_26327);
nand U39919 (N_39919,N_29385,N_25405);
and U39920 (N_39920,N_28184,N_24799);
nor U39921 (N_39921,N_22084,N_23935);
or U39922 (N_39922,N_23018,N_24281);
nor U39923 (N_39923,N_25735,N_24730);
and U39924 (N_39924,N_29386,N_27032);
and U39925 (N_39925,N_29316,N_27879);
xnor U39926 (N_39926,N_28525,N_23243);
nand U39927 (N_39927,N_21617,N_28312);
xnor U39928 (N_39928,N_23612,N_25598);
nand U39929 (N_39929,N_23973,N_29901);
nand U39930 (N_39930,N_23509,N_25159);
and U39931 (N_39931,N_27579,N_21173);
and U39932 (N_39932,N_23670,N_24500);
xnor U39933 (N_39933,N_21831,N_25024);
nor U39934 (N_39934,N_23419,N_21913);
or U39935 (N_39935,N_24201,N_28330);
nor U39936 (N_39936,N_27995,N_28522);
nor U39937 (N_39937,N_28674,N_22654);
or U39938 (N_39938,N_26874,N_25092);
nor U39939 (N_39939,N_22510,N_20983);
or U39940 (N_39940,N_21930,N_28906);
nor U39941 (N_39941,N_22087,N_22987);
or U39942 (N_39942,N_24695,N_22660);
and U39943 (N_39943,N_20061,N_22344);
or U39944 (N_39944,N_26864,N_27155);
or U39945 (N_39945,N_29494,N_28244);
nand U39946 (N_39946,N_25271,N_26684);
nand U39947 (N_39947,N_29064,N_26877);
xnor U39948 (N_39948,N_26410,N_24493);
or U39949 (N_39949,N_21303,N_21804);
or U39950 (N_39950,N_28231,N_22970);
xor U39951 (N_39951,N_20627,N_26761);
and U39952 (N_39952,N_21299,N_25737);
nor U39953 (N_39953,N_20547,N_26927);
nor U39954 (N_39954,N_28943,N_23288);
or U39955 (N_39955,N_23742,N_23893);
or U39956 (N_39956,N_29657,N_22381);
nand U39957 (N_39957,N_23755,N_26480);
or U39958 (N_39958,N_28875,N_20662);
nor U39959 (N_39959,N_24698,N_22375);
nor U39960 (N_39960,N_27765,N_22158);
and U39961 (N_39961,N_23696,N_29105);
or U39962 (N_39962,N_26336,N_20770);
nor U39963 (N_39963,N_22688,N_23701);
and U39964 (N_39964,N_20637,N_24038);
and U39965 (N_39965,N_23482,N_23456);
or U39966 (N_39966,N_28582,N_28304);
nor U39967 (N_39967,N_29495,N_28048);
xor U39968 (N_39968,N_26247,N_28336);
nand U39969 (N_39969,N_25409,N_29281);
nor U39970 (N_39970,N_20356,N_26440);
xnor U39971 (N_39971,N_24937,N_20002);
nor U39972 (N_39972,N_23468,N_23022);
xnor U39973 (N_39973,N_29626,N_26928);
or U39974 (N_39974,N_28344,N_21065);
nand U39975 (N_39975,N_29093,N_20988);
nand U39976 (N_39976,N_29288,N_29646);
nor U39977 (N_39977,N_23082,N_28671);
and U39978 (N_39978,N_22216,N_28015);
or U39979 (N_39979,N_23216,N_26164);
nor U39980 (N_39980,N_23028,N_28198);
or U39981 (N_39981,N_29016,N_24118);
nor U39982 (N_39982,N_23623,N_22338);
and U39983 (N_39983,N_23950,N_25593);
and U39984 (N_39984,N_20472,N_23444);
xnor U39985 (N_39985,N_21692,N_28699);
and U39986 (N_39986,N_26418,N_20834);
or U39987 (N_39987,N_25350,N_24065);
xor U39988 (N_39988,N_29139,N_20569);
or U39989 (N_39989,N_22365,N_28465);
nor U39990 (N_39990,N_21032,N_22288);
nand U39991 (N_39991,N_25806,N_20834);
xor U39992 (N_39992,N_26920,N_23479);
xor U39993 (N_39993,N_28989,N_25986);
or U39994 (N_39994,N_23346,N_22440);
and U39995 (N_39995,N_28506,N_21892);
xnor U39996 (N_39996,N_27977,N_21959);
nor U39997 (N_39997,N_28918,N_29313);
nor U39998 (N_39998,N_20450,N_26429);
nor U39999 (N_39999,N_21188,N_24383);
or U40000 (N_40000,N_39170,N_36592);
and U40001 (N_40001,N_32596,N_38366);
xor U40002 (N_40002,N_30996,N_33355);
nand U40003 (N_40003,N_33193,N_38726);
nor U40004 (N_40004,N_37517,N_37618);
or U40005 (N_40005,N_34997,N_31821);
and U40006 (N_40006,N_31766,N_30735);
xor U40007 (N_40007,N_31746,N_35195);
and U40008 (N_40008,N_35666,N_38397);
xor U40009 (N_40009,N_37152,N_34507);
nor U40010 (N_40010,N_35765,N_35657);
or U40011 (N_40011,N_31603,N_30997);
xnor U40012 (N_40012,N_39007,N_36812);
and U40013 (N_40013,N_31896,N_31576);
xnor U40014 (N_40014,N_36604,N_32117);
nor U40015 (N_40015,N_39915,N_36331);
nand U40016 (N_40016,N_34889,N_33917);
nand U40017 (N_40017,N_39069,N_32160);
nor U40018 (N_40018,N_30740,N_39533);
xnor U40019 (N_40019,N_38701,N_39630);
or U40020 (N_40020,N_35351,N_33559);
nor U40021 (N_40021,N_34002,N_30844);
or U40022 (N_40022,N_38999,N_38911);
and U40023 (N_40023,N_35529,N_35031);
or U40024 (N_40024,N_32539,N_38024);
and U40025 (N_40025,N_33424,N_30354);
and U40026 (N_40026,N_30777,N_33745);
or U40027 (N_40027,N_32244,N_30050);
xnor U40028 (N_40028,N_37626,N_38359);
or U40029 (N_40029,N_38810,N_39948);
or U40030 (N_40030,N_38161,N_37584);
nor U40031 (N_40031,N_37923,N_36386);
or U40032 (N_40032,N_39378,N_30455);
nand U40033 (N_40033,N_30813,N_35285);
nor U40034 (N_40034,N_36351,N_32191);
nor U40035 (N_40035,N_34829,N_36783);
nor U40036 (N_40036,N_39256,N_30310);
and U40037 (N_40037,N_33812,N_31569);
and U40038 (N_40038,N_31742,N_30960);
or U40039 (N_40039,N_34781,N_39566);
nor U40040 (N_40040,N_34280,N_33976);
or U40041 (N_40041,N_33581,N_36194);
nand U40042 (N_40042,N_37253,N_34783);
nor U40043 (N_40043,N_33501,N_33012);
nand U40044 (N_40044,N_34995,N_34826);
and U40045 (N_40045,N_37762,N_33208);
or U40046 (N_40046,N_38164,N_38058);
xor U40047 (N_40047,N_35770,N_32826);
or U40048 (N_40048,N_34100,N_35672);
or U40049 (N_40049,N_30421,N_39552);
and U40050 (N_40050,N_38186,N_39964);
and U40051 (N_40051,N_34805,N_34957);
or U40052 (N_40052,N_32934,N_34285);
or U40053 (N_40053,N_39708,N_33342);
xor U40054 (N_40054,N_37644,N_33196);
or U40055 (N_40055,N_31253,N_30600);
and U40056 (N_40056,N_36537,N_31056);
and U40057 (N_40057,N_39923,N_37023);
xnor U40058 (N_40058,N_33945,N_34969);
nand U40059 (N_40059,N_34110,N_34648);
xor U40060 (N_40060,N_34261,N_39308);
and U40061 (N_40061,N_36020,N_37222);
nor U40062 (N_40062,N_35947,N_36023);
or U40063 (N_40063,N_37579,N_31709);
nand U40064 (N_40064,N_35861,N_38669);
and U40065 (N_40065,N_35948,N_36927);
and U40066 (N_40066,N_34204,N_34160);
or U40067 (N_40067,N_30937,N_31340);
nand U40068 (N_40068,N_36790,N_39640);
nor U40069 (N_40069,N_38070,N_34707);
or U40070 (N_40070,N_36650,N_39084);
and U40071 (N_40071,N_37126,N_32995);
nor U40072 (N_40072,N_36244,N_39614);
or U40073 (N_40073,N_35725,N_30432);
nor U40074 (N_40074,N_35302,N_36958);
xnor U40075 (N_40075,N_37702,N_34152);
or U40076 (N_40076,N_35906,N_39786);
nand U40077 (N_40077,N_31157,N_33431);
or U40078 (N_40078,N_36833,N_34134);
xor U40079 (N_40079,N_36229,N_36251);
nor U40080 (N_40080,N_31502,N_35495);
or U40081 (N_40081,N_36926,N_39156);
and U40082 (N_40082,N_38025,N_30678);
xor U40083 (N_40083,N_33029,N_38878);
nor U40084 (N_40084,N_37337,N_30144);
nand U40085 (N_40085,N_36085,N_30139);
or U40086 (N_40086,N_36853,N_35581);
and U40087 (N_40087,N_37563,N_31016);
or U40088 (N_40088,N_35373,N_39992);
nand U40089 (N_40089,N_32711,N_31680);
nand U40090 (N_40090,N_34510,N_38901);
or U40091 (N_40091,N_30918,N_31130);
and U40092 (N_40092,N_31833,N_34586);
nor U40093 (N_40093,N_36755,N_38430);
or U40094 (N_40094,N_38286,N_31822);
xnor U40095 (N_40095,N_38087,N_34190);
and U40096 (N_40096,N_32757,N_31879);
nand U40097 (N_40097,N_36613,N_35273);
or U40098 (N_40098,N_31198,N_39743);
xnor U40099 (N_40099,N_34474,N_38806);
and U40100 (N_40100,N_35157,N_37919);
xnor U40101 (N_40101,N_37353,N_36193);
and U40102 (N_40102,N_35460,N_30296);
or U40103 (N_40103,N_31917,N_35257);
nand U40104 (N_40104,N_32975,N_32053);
xor U40105 (N_40105,N_35989,N_39840);
xnor U40106 (N_40106,N_30917,N_34464);
xor U40107 (N_40107,N_31074,N_33489);
or U40108 (N_40108,N_38884,N_32509);
or U40109 (N_40109,N_32305,N_39876);
nor U40110 (N_40110,N_34535,N_35835);
xnor U40111 (N_40111,N_37578,N_34643);
or U40112 (N_40112,N_37371,N_38222);
or U40113 (N_40113,N_33503,N_32601);
or U40114 (N_40114,N_32806,N_32518);
nor U40115 (N_40115,N_37121,N_32953);
xor U40116 (N_40116,N_33135,N_30157);
xor U40117 (N_40117,N_36630,N_35106);
nand U40118 (N_40118,N_32331,N_31700);
xor U40119 (N_40119,N_34135,N_38332);
nor U40120 (N_40120,N_33477,N_39206);
and U40121 (N_40121,N_37080,N_33632);
nor U40122 (N_40122,N_33218,N_36629);
or U40123 (N_40123,N_39961,N_39150);
and U40124 (N_40124,N_34545,N_33353);
and U40125 (N_40125,N_32389,N_37120);
xnor U40126 (N_40126,N_35970,N_34999);
or U40127 (N_40127,N_33289,N_39398);
nor U40128 (N_40128,N_30214,N_31175);
xnor U40129 (N_40129,N_36907,N_33443);
or U40130 (N_40130,N_39292,N_36533);
or U40131 (N_40131,N_33893,N_37770);
or U40132 (N_40132,N_37603,N_38303);
nand U40133 (N_40133,N_33921,N_37409);
nor U40134 (N_40134,N_33275,N_34131);
xnor U40135 (N_40135,N_34562,N_38352);
and U40136 (N_40136,N_34668,N_36401);
nand U40137 (N_40137,N_38188,N_38441);
or U40138 (N_40138,N_30905,N_34048);
or U40139 (N_40139,N_37532,N_33832);
or U40140 (N_40140,N_39208,N_32944);
and U40141 (N_40141,N_32778,N_37986);
nand U40142 (N_40142,N_30908,N_31254);
and U40143 (N_40143,N_39360,N_37103);
nand U40144 (N_40144,N_39502,N_31421);
xnor U40145 (N_40145,N_33024,N_38549);
nand U40146 (N_40146,N_32795,N_33091);
nand U40147 (N_40147,N_33594,N_37464);
and U40148 (N_40148,N_37412,N_38892);
or U40149 (N_40149,N_32215,N_36339);
xnor U40150 (N_40150,N_38723,N_33237);
nor U40151 (N_40151,N_36036,N_39189);
or U40152 (N_40152,N_34466,N_30229);
and U40153 (N_40153,N_32484,N_30130);
nor U40154 (N_40154,N_34671,N_39483);
nand U40155 (N_40155,N_38107,N_39355);
nand U40156 (N_40156,N_34614,N_36614);
nand U40157 (N_40157,N_39938,N_32118);
nand U40158 (N_40158,N_30665,N_38801);
nor U40159 (N_40159,N_32306,N_30829);
or U40160 (N_40160,N_39392,N_33294);
nor U40161 (N_40161,N_32132,N_34169);
xor U40162 (N_40162,N_34684,N_32572);
and U40163 (N_40163,N_30867,N_36204);
xor U40164 (N_40164,N_31278,N_35613);
and U40165 (N_40165,N_36273,N_34666);
and U40166 (N_40166,N_35566,N_39551);
xnor U40167 (N_40167,N_39489,N_35342);
xnor U40168 (N_40168,N_35082,N_34813);
and U40169 (N_40169,N_33049,N_30344);
nor U40170 (N_40170,N_36071,N_33607);
and U40171 (N_40171,N_39463,N_31462);
nand U40172 (N_40172,N_36113,N_35689);
or U40173 (N_40173,N_30962,N_32649);
or U40174 (N_40174,N_33017,N_32514);
or U40175 (N_40175,N_33671,N_35251);
or U40176 (N_40176,N_31834,N_36561);
nor U40177 (N_40177,N_32024,N_36149);
nand U40178 (N_40178,N_30709,N_32497);
nand U40179 (N_40179,N_32230,N_39271);
nor U40180 (N_40180,N_38460,N_36298);
xor U40181 (N_40181,N_35510,N_37311);
and U40182 (N_40182,N_37073,N_38822);
and U40183 (N_40183,N_32663,N_33171);
and U40184 (N_40184,N_36024,N_30430);
nor U40185 (N_40185,N_37436,N_38106);
xnor U40186 (N_40186,N_34469,N_35958);
or U40187 (N_40187,N_39092,N_34955);
nand U40188 (N_40188,N_33247,N_33401);
and U40189 (N_40189,N_32499,N_30210);
nor U40190 (N_40190,N_36782,N_34254);
xor U40191 (N_40191,N_31868,N_36901);
xor U40192 (N_40192,N_35057,N_35079);
nor U40193 (N_40193,N_36482,N_33537);
and U40194 (N_40194,N_33777,N_32202);
nand U40195 (N_40195,N_30264,N_34639);
nor U40196 (N_40196,N_33156,N_33755);
nand U40197 (N_40197,N_35467,N_33357);
xnor U40198 (N_40198,N_38381,N_38653);
nand U40199 (N_40199,N_33839,N_38264);
and U40200 (N_40200,N_38679,N_32654);
and U40201 (N_40201,N_33323,N_34594);
or U40202 (N_40202,N_37239,N_30878);
or U40203 (N_40203,N_39372,N_38076);
nor U40204 (N_40204,N_39823,N_32843);
nand U40205 (N_40205,N_31855,N_32164);
xnor U40206 (N_40206,N_38829,N_31374);
and U40207 (N_40207,N_31574,N_35368);
nor U40208 (N_40208,N_31108,N_35269);
and U40209 (N_40209,N_38900,N_35232);
nand U40210 (N_40210,N_31059,N_34393);
nand U40211 (N_40211,N_33441,N_34461);
nand U40212 (N_40212,N_36662,N_37641);
and U40213 (N_40213,N_31748,N_35642);
and U40214 (N_40214,N_36679,N_38190);
nand U40215 (N_40215,N_37444,N_36064);
nor U40216 (N_40216,N_37031,N_36004);
and U40217 (N_40217,N_37289,N_34034);
and U40218 (N_40218,N_31804,N_39249);
xor U40219 (N_40219,N_30909,N_34253);
nor U40220 (N_40220,N_37056,N_35254);
or U40221 (N_40221,N_36364,N_38592);
nor U40222 (N_40222,N_30401,N_33784);
nand U40223 (N_40223,N_37482,N_33059);
nand U40224 (N_40224,N_30358,N_32688);
or U40225 (N_40225,N_37585,N_39088);
and U40226 (N_40226,N_32114,N_35454);
xnor U40227 (N_40227,N_34916,N_39982);
xor U40228 (N_40228,N_36252,N_30550);
or U40229 (N_40229,N_35793,N_32436);
xnor U40230 (N_40230,N_39612,N_35651);
xor U40231 (N_40231,N_32796,N_35029);
nand U40232 (N_40232,N_38557,N_32977);
xnor U40233 (N_40233,N_30887,N_36306);
nand U40234 (N_40234,N_32985,N_37571);
and U40235 (N_40235,N_38895,N_34654);
nor U40236 (N_40236,N_36959,N_31900);
xor U40237 (N_40237,N_30817,N_39265);
nor U40238 (N_40238,N_39373,N_36779);
and U40239 (N_40239,N_35927,N_38992);
nor U40240 (N_40240,N_33541,N_35653);
or U40241 (N_40241,N_30062,N_33269);
nand U40242 (N_40242,N_33308,N_37297);
xnor U40243 (N_40243,N_31832,N_30171);
and U40244 (N_40244,N_36921,N_39247);
xnor U40245 (N_40245,N_37556,N_34624);
nor U40246 (N_40246,N_31427,N_38432);
or U40247 (N_40247,N_30435,N_30220);
and U40248 (N_40248,N_38338,N_37065);
and U40249 (N_40249,N_34619,N_36269);
nand U40250 (N_40250,N_30679,N_36741);
nand U40251 (N_40251,N_39456,N_39830);
and U40252 (N_40252,N_36432,N_35261);
nor U40253 (N_40253,N_39179,N_30675);
and U40254 (N_40254,N_37396,N_39268);
nor U40255 (N_40255,N_38135,N_33154);
xnor U40256 (N_40256,N_35239,N_35663);
xnor U40257 (N_40257,N_36624,N_32968);
nor U40258 (N_40258,N_33788,N_39324);
nand U40259 (N_40259,N_39998,N_38849);
and U40260 (N_40260,N_30570,N_34233);
nor U40261 (N_40261,N_31031,N_38554);
xor U40262 (N_40262,N_39736,N_39541);
and U40263 (N_40263,N_35518,N_38240);
and U40264 (N_40264,N_36731,N_35789);
xor U40265 (N_40265,N_35625,N_36439);
nand U40266 (N_40266,N_36483,N_30630);
or U40267 (N_40267,N_33924,N_39760);
nand U40268 (N_40268,N_36235,N_33414);
or U40269 (N_40269,N_39592,N_31135);
nor U40270 (N_40270,N_39861,N_36658);
nand U40271 (N_40271,N_33348,N_31506);
xnor U40272 (N_40272,N_30333,N_36261);
xor U40273 (N_40273,N_34968,N_37540);
xnor U40274 (N_40274,N_37053,N_39590);
or U40275 (N_40275,N_34747,N_33300);
nand U40276 (N_40276,N_30206,N_34455);
or U40277 (N_40277,N_37098,N_31755);
xnor U40278 (N_40278,N_38238,N_36325);
and U40279 (N_40279,N_36574,N_35867);
and U40280 (N_40280,N_31629,N_30102);
nor U40281 (N_40281,N_37359,N_38559);
nand U40282 (N_40282,N_35309,N_35218);
and U40283 (N_40283,N_37700,N_34788);
and U40284 (N_40284,N_33530,N_37953);
and U40285 (N_40285,N_31751,N_30190);
xnor U40286 (N_40286,N_38828,N_36348);
nand U40287 (N_40287,N_37821,N_36725);
nor U40288 (N_40288,N_37831,N_35217);
and U40289 (N_40289,N_33699,N_36195);
and U40290 (N_40290,N_33078,N_33066);
and U40291 (N_40291,N_34574,N_31286);
nand U40292 (N_40292,N_34255,N_30546);
and U40293 (N_40293,N_38093,N_39101);
or U40294 (N_40294,N_30127,N_34141);
nand U40295 (N_40295,N_38062,N_39564);
nand U40296 (N_40296,N_36358,N_38817);
nor U40297 (N_40297,N_39433,N_37000);
xor U40298 (N_40298,N_32676,N_31850);
nor U40299 (N_40299,N_35104,N_31568);
nor U40300 (N_40300,N_30477,N_34956);
xor U40301 (N_40301,N_33292,N_30521);
and U40302 (N_40302,N_33800,N_39675);
xnor U40303 (N_40303,N_32410,N_37048);
and U40304 (N_40304,N_36890,N_33318);
and U40305 (N_40305,N_36014,N_33822);
and U40306 (N_40306,N_34154,N_31885);
xnor U40307 (N_40307,N_33250,N_36322);
or U40308 (N_40308,N_33402,N_33056);
or U40309 (N_40309,N_36724,N_32814);
or U40310 (N_40310,N_39581,N_37471);
xnor U40311 (N_40311,N_33031,N_30170);
and U40312 (N_40312,N_34918,N_36259);
nor U40313 (N_40313,N_39722,N_34682);
nand U40314 (N_40314,N_37734,N_35441);
nor U40315 (N_40315,N_37835,N_37713);
nand U40316 (N_40316,N_39495,N_39266);
nand U40317 (N_40317,N_32480,N_30099);
xnor U40318 (N_40318,N_32470,N_31282);
or U40319 (N_40319,N_37674,N_37234);
nor U40320 (N_40320,N_39738,N_38871);
and U40321 (N_40321,N_30987,N_38585);
nor U40322 (N_40322,N_30213,N_38143);
nor U40323 (N_40323,N_32319,N_33975);
and U40324 (N_40324,N_32235,N_35627);
nand U40325 (N_40325,N_30769,N_32072);
nor U40326 (N_40326,N_36478,N_33715);
nor U40327 (N_40327,N_32219,N_37845);
xnor U40328 (N_40328,N_38044,N_31317);
nor U40329 (N_40329,N_35860,N_33930);
nand U40330 (N_40330,N_39157,N_38328);
or U40331 (N_40331,N_36743,N_34570);
nor U40332 (N_40332,N_32693,N_32987);
or U40333 (N_40333,N_31396,N_38162);
nand U40334 (N_40334,N_35509,N_31276);
xor U40335 (N_40335,N_30388,N_31444);
and U40336 (N_40336,N_37271,N_34333);
or U40337 (N_40337,N_34281,N_35694);
nor U40338 (N_40338,N_34884,N_37173);
nand U40339 (N_40339,N_33490,N_39971);
nor U40340 (N_40340,N_33377,N_31600);
or U40341 (N_40341,N_35857,N_30682);
nor U40342 (N_40342,N_34667,N_31435);
nand U40343 (N_40343,N_36840,N_33844);
xor U40344 (N_40344,N_30199,N_34827);
xor U40345 (N_40345,N_37564,N_37561);
nor U40346 (N_40346,N_39250,N_36615);
and U40347 (N_40347,N_33825,N_38533);
xor U40348 (N_40348,N_35372,N_33046);
nor U40349 (N_40349,N_30319,N_38204);
and U40350 (N_40350,N_37841,N_35396);
xor U40351 (N_40351,N_37320,N_34547);
nand U40352 (N_40352,N_35626,N_32091);
xor U40353 (N_40353,N_33714,N_33560);
nand U40354 (N_40354,N_32699,N_30003);
or U40355 (N_40355,N_35681,N_36153);
xor U40356 (N_40356,N_37625,N_38803);
or U40357 (N_40357,N_39568,N_33068);
nor U40358 (N_40358,N_34998,N_37962);
and U40359 (N_40359,N_32150,N_35300);
or U40360 (N_40360,N_36808,N_30552);
xnor U40361 (N_40361,N_35856,N_36506);
or U40362 (N_40362,N_31187,N_38777);
or U40363 (N_40363,N_33586,N_37972);
and U40364 (N_40364,N_32682,N_34677);
xnor U40365 (N_40365,N_34198,N_30470);
xnor U40366 (N_40366,N_36437,N_36215);
or U40367 (N_40367,N_30362,N_35698);
xnor U40368 (N_40368,N_30737,N_31669);
nor U40369 (N_40369,N_37358,N_38142);
or U40370 (N_40370,N_33635,N_31474);
or U40371 (N_40371,N_37782,N_37410);
nand U40372 (N_40372,N_33067,N_38289);
xnor U40373 (N_40373,N_34246,N_33325);
nand U40374 (N_40374,N_36616,N_39070);
xnor U40375 (N_40375,N_33992,N_37435);
xor U40376 (N_40376,N_39727,N_33876);
nand U40377 (N_40377,N_34114,N_34436);
xnor U40378 (N_40378,N_30954,N_32505);
xnor U40379 (N_40379,N_37500,N_34818);
nor U40380 (N_40380,N_34681,N_31251);
xnor U40381 (N_40381,N_30481,N_38261);
and U40382 (N_40382,N_33077,N_31214);
nor U40383 (N_40383,N_39406,N_31429);
or U40384 (N_40384,N_32149,N_35552);
nand U40385 (N_40385,N_30591,N_39718);
nor U40386 (N_40386,N_34387,N_37523);
and U40387 (N_40387,N_32898,N_37495);
xnor U40388 (N_40388,N_33816,N_30669);
nor U40389 (N_40389,N_31649,N_31263);
xnor U40390 (N_40390,N_35167,N_33799);
or U40391 (N_40391,N_38475,N_39775);
and U40392 (N_40392,N_30270,N_37880);
and U40393 (N_40393,N_31118,N_39939);
nand U40394 (N_40394,N_36067,N_31332);
nor U40395 (N_40395,N_37350,N_33284);
nor U40396 (N_40396,N_37913,N_34795);
nor U40397 (N_40397,N_30991,N_31392);
xnor U40398 (N_40398,N_39023,N_37966);
or U40399 (N_40399,N_39458,N_30431);
xor U40400 (N_40400,N_30778,N_37441);
nand U40401 (N_40401,N_33551,N_31871);
xor U40402 (N_40402,N_34375,N_34180);
or U40403 (N_40403,N_35829,N_31371);
and U40404 (N_40404,N_33287,N_37251);
nor U40405 (N_40405,N_31580,N_33644);
nor U40406 (N_40406,N_33556,N_39677);
and U40407 (N_40407,N_30309,N_38156);
or U40408 (N_40408,N_37695,N_33257);
and U40409 (N_40409,N_39571,N_35719);
xnor U40410 (N_40410,N_39237,N_32580);
nand U40411 (N_40411,N_36718,N_33449);
and U40412 (N_40412,N_33994,N_33487);
nand U40413 (N_40413,N_30766,N_34457);
and U40414 (N_40414,N_34628,N_32366);
or U40415 (N_40415,N_34480,N_31012);
xnor U40416 (N_40416,N_38239,N_39908);
nand U40417 (N_40417,N_34277,N_32055);
and U40418 (N_40418,N_35574,N_36497);
xor U40419 (N_40419,N_31109,N_34028);
nor U40420 (N_40420,N_33923,N_37930);
nor U40421 (N_40421,N_36970,N_34496);
nor U40422 (N_40422,N_32128,N_30352);
or U40423 (N_40423,N_39450,N_37007);
nor U40424 (N_40424,N_31705,N_30248);
nor U40425 (N_40425,N_31092,N_31139);
nor U40426 (N_40426,N_37951,N_31794);
nor U40427 (N_40427,N_38619,N_36530);
xnor U40428 (N_40428,N_33422,N_39046);
or U40429 (N_40429,N_33080,N_35158);
xnor U40430 (N_40430,N_33895,N_34903);
or U40431 (N_40431,N_36197,N_35497);
xor U40432 (N_40432,N_38127,N_31323);
or U40433 (N_40433,N_32489,N_34075);
and U40434 (N_40434,N_37983,N_32491);
and U40435 (N_40435,N_34740,N_34683);
and U40436 (N_40436,N_30635,N_30230);
or U40437 (N_40437,N_38456,N_36266);
nand U40438 (N_40438,N_30594,N_35123);
nand U40439 (N_40439,N_36220,N_31769);
nor U40440 (N_40440,N_38514,N_34650);
and U40441 (N_40441,N_36988,N_37077);
nor U40442 (N_40442,N_30695,N_31131);
nor U40443 (N_40443,N_38981,N_33460);
and U40444 (N_40444,N_33691,N_35920);
xnor U40445 (N_40445,N_39492,N_37419);
xnor U40446 (N_40446,N_34404,N_39141);
nor U40447 (N_40447,N_39213,N_34822);
nor U40448 (N_40448,N_33969,N_35228);
nor U40449 (N_40449,N_30166,N_32359);
xor U40450 (N_40450,N_36019,N_32506);
xor U40451 (N_40451,N_37748,N_33925);
xor U40452 (N_40452,N_34336,N_36335);
xnor U40453 (N_40453,N_36795,N_38390);
nor U40454 (N_40454,N_31385,N_37487);
or U40455 (N_40455,N_39093,N_32827);
nor U40456 (N_40456,N_38593,N_30577);
nand U40457 (N_40457,N_30450,N_35744);
or U40458 (N_40458,N_32408,N_39269);
and U40459 (N_40459,N_34528,N_34537);
xor U40460 (N_40460,N_37623,N_36507);
nand U40461 (N_40461,N_38171,N_34565);
and U40462 (N_40462,N_31901,N_33946);
xnor U40463 (N_40463,N_37383,N_32268);
or U40464 (N_40464,N_30859,N_35570);
xor U40465 (N_40465,N_35282,N_32208);
and U40466 (N_40466,N_36665,N_30267);
or U40467 (N_40467,N_37530,N_30400);
or U40468 (N_40468,N_31265,N_30820);
or U40469 (N_40469,N_31053,N_34943);
nand U40470 (N_40470,N_38422,N_36281);
or U40471 (N_40471,N_38485,N_30952);
nor U40472 (N_40472,N_31888,N_33748);
or U40473 (N_40473,N_38975,N_30676);
and U40474 (N_40474,N_33179,N_36874);
or U40475 (N_40475,N_36379,N_35586);
nor U40476 (N_40476,N_38713,N_34658);
and U40477 (N_40477,N_36203,N_31102);
xnor U40478 (N_40478,N_30294,N_37881);
and U40479 (N_40479,N_32146,N_36385);
and U40480 (N_40480,N_34766,N_38212);
xnor U40481 (N_40481,N_35221,N_37418);
xor U40482 (N_40482,N_37887,N_37593);
nand U40483 (N_40483,N_35832,N_38956);
and U40484 (N_40484,N_39205,N_37308);
xor U40485 (N_40485,N_36960,N_39231);
or U40486 (N_40486,N_38082,N_36257);
nor U40487 (N_40487,N_39798,N_37064);
and U40488 (N_40488,N_35364,N_37392);
and U40489 (N_40489,N_39678,N_39076);
nor U40490 (N_40490,N_37589,N_39874);
xnor U40491 (N_40491,N_34768,N_34569);
or U40492 (N_40492,N_33576,N_39476);
nor U40493 (N_40493,N_31757,N_35640);
and U40494 (N_40494,N_30473,N_31233);
nand U40495 (N_40495,N_38147,N_38545);
nor U40496 (N_40496,N_35577,N_39839);
nor U40497 (N_40497,N_39868,N_39696);
xor U40498 (N_40498,N_39331,N_30637);
nand U40499 (N_40499,N_37453,N_33086);
nand U40500 (N_40500,N_31986,N_39638);
or U40501 (N_40501,N_33915,N_32612);
and U40502 (N_40502,N_37654,N_35448);
and U40503 (N_40503,N_30771,N_37160);
nor U40504 (N_40504,N_38636,N_31466);
and U40505 (N_40505,N_36643,N_32714);
xor U40506 (N_40506,N_34580,N_35420);
nand U40507 (N_40507,N_32272,N_32095);
nor U40508 (N_40508,N_35402,N_37638);
nor U40509 (N_40509,N_31687,N_36253);
or U40510 (N_40510,N_39517,N_30005);
nor U40511 (N_40511,N_38918,N_39739);
nor U40512 (N_40512,N_33598,N_33986);
or U40513 (N_40513,N_35466,N_34129);
nand U40514 (N_40514,N_30943,N_38098);
xor U40515 (N_40515,N_38666,N_34244);
xor U40516 (N_40516,N_31594,N_35965);
xnor U40517 (N_40517,N_36106,N_35598);
xnor U40518 (N_40518,N_34990,N_32104);
nand U40519 (N_40519,N_33148,N_36223);
or U40520 (N_40520,N_37724,N_39668);
nand U40521 (N_40521,N_30612,N_39479);
xnor U40522 (N_40522,N_36999,N_32168);
nor U40523 (N_40523,N_32116,N_32392);
nor U40524 (N_40524,N_33139,N_36882);
nand U40525 (N_40525,N_38620,N_30956);
xor U40526 (N_40526,N_34806,N_38189);
nor U40527 (N_40527,N_39885,N_33214);
nor U40528 (N_40528,N_36017,N_30701);
nand U40529 (N_40529,N_35652,N_39952);
and U40530 (N_40530,N_34659,N_30459);
nand U40531 (N_40531,N_35916,N_38350);
and U40532 (N_40532,N_36154,N_36706);
and U40533 (N_40533,N_37391,N_34062);
or U40534 (N_40534,N_35365,N_34268);
xor U40535 (N_40535,N_39768,N_31839);
or U40536 (N_40536,N_36357,N_31204);
and U40537 (N_40537,N_39949,N_34530);
and U40538 (N_40538,N_31291,N_38906);
nor U40539 (N_40539,N_35236,N_35099);
nand U40540 (N_40540,N_36097,N_30080);
xnor U40541 (N_40541,N_34548,N_38897);
and U40542 (N_40542,N_30014,N_30095);
xor U40543 (N_40543,N_35997,N_33680);
nand U40544 (N_40544,N_31230,N_38103);
nand U40545 (N_40545,N_33213,N_35243);
and U40546 (N_40546,N_31514,N_32720);
and U40547 (N_40547,N_32618,N_30071);
xnor U40548 (N_40548,N_35699,N_38199);
and U40549 (N_40549,N_38919,N_39192);
nand U40550 (N_40550,N_34676,N_32726);
or U40551 (N_40551,N_33122,N_35140);
nand U40552 (N_40552,N_34159,N_33571);
xor U40553 (N_40553,N_37955,N_36247);
and U40554 (N_40554,N_32617,N_30364);
nand U40555 (N_40555,N_34984,N_34311);
or U40556 (N_40556,N_35609,N_35683);
and U40557 (N_40557,N_32967,N_30822);
xor U40558 (N_40558,N_36954,N_31178);
or U40559 (N_40559,N_33793,N_33311);
or U40560 (N_40560,N_36906,N_38023);
xnor U40561 (N_40561,N_34330,N_34313);
and U40562 (N_40562,N_36005,N_32309);
or U40563 (N_40563,N_33941,N_31487);
or U40564 (N_40564,N_33260,N_34481);
xnor U40565 (N_40565,N_32195,N_39124);
nand U40566 (N_40566,N_36425,N_30356);
or U40567 (N_40567,N_33456,N_30645);
nor U40568 (N_40568,N_31965,N_33900);
nand U40569 (N_40569,N_39881,N_37148);
nand U40570 (N_40570,N_33483,N_32263);
or U40571 (N_40571,N_30348,N_31202);
or U40572 (N_40572,N_31524,N_36034);
or U40573 (N_40573,N_38949,N_37302);
nor U40574 (N_40574,N_31566,N_34043);
and U40575 (N_40575,N_34019,N_37617);
nor U40576 (N_40576,N_39538,N_35612);
or U40577 (N_40577,N_31107,N_39212);
xor U40578 (N_40578,N_35423,N_37321);
xor U40579 (N_40579,N_31872,N_35736);
nor U40580 (N_40580,N_36199,N_39434);
and U40581 (N_40581,N_36167,N_32681);
and U40582 (N_40582,N_33362,N_35664);
and U40583 (N_40583,N_34724,N_30619);
nor U40584 (N_40584,N_32517,N_30054);
nand U40585 (N_40585,N_34801,N_34420);
or U40586 (N_40586,N_39981,N_38749);
nor U40587 (N_40587,N_39799,N_38128);
or U40588 (N_40588,N_32932,N_33102);
nand U40589 (N_40589,N_33302,N_39086);
xnor U40590 (N_40590,N_33178,N_32100);
nand U40591 (N_40591,N_31761,N_36456);
xnor U40592 (N_40592,N_35704,N_34780);
or U40593 (N_40593,N_37811,N_34315);
nor U40594 (N_40594,N_33539,N_32362);
xnor U40595 (N_40595,N_38440,N_33221);
nor U40596 (N_40596,N_32052,N_38271);
nor U40597 (N_40597,N_33519,N_35980);
nand U40598 (N_40598,N_30195,N_35130);
or U40599 (N_40599,N_31841,N_38925);
xor U40600 (N_40600,N_30088,N_30075);
nand U40601 (N_40601,N_31115,N_33873);
nor U40602 (N_40602,N_36488,N_37975);
nor U40603 (N_40603,N_36081,N_34241);
nand U40604 (N_40604,N_30493,N_39548);
xor U40605 (N_40605,N_39290,N_32836);
or U40606 (N_40606,N_33564,N_36326);
or U40607 (N_40607,N_32749,N_32194);
xnor U40608 (N_40608,N_38519,N_30098);
xnor U40609 (N_40609,N_39731,N_39123);
or U40610 (N_40610,N_30208,N_39145);
and U40611 (N_40611,N_31765,N_36594);
and U40612 (N_40612,N_34199,N_37504);
nand U40613 (N_40613,N_32181,N_38754);
nand U40614 (N_40614,N_35579,N_39100);
nor U40615 (N_40615,N_35884,N_30583);
and U40616 (N_40616,N_31382,N_36118);
nor U40617 (N_40617,N_30387,N_30781);
and U40618 (N_40618,N_30707,N_35485);
xor U40619 (N_40619,N_36242,N_30205);
nor U40620 (N_40620,N_36291,N_30060);
nand U40621 (N_40621,N_37833,N_36139);
nor U40622 (N_40622,N_34820,N_32815);
xnor U40623 (N_40623,N_30703,N_34056);
xnor U40624 (N_40624,N_35516,N_39703);
and U40625 (N_40625,N_30442,N_33709);
nand U40626 (N_40626,N_32466,N_33481);
and U40627 (N_40627,N_32363,N_33430);
nand U40628 (N_40628,N_33716,N_33765);
nand U40629 (N_40629,N_35935,N_37197);
nor U40630 (N_40630,N_32603,N_37689);
xor U40631 (N_40631,N_33200,N_32798);
nor U40632 (N_40632,N_37733,N_37791);
nor U40633 (N_40633,N_33124,N_38132);
nand U40634 (N_40634,N_30239,N_37079);
xor U40635 (N_40635,N_32808,N_31163);
and U40636 (N_40636,N_32587,N_38640);
nor U40637 (N_40637,N_37040,N_34531);
nor U40638 (N_40638,N_33701,N_35558);
xnor U40639 (N_40639,N_34446,N_39350);
or U40640 (N_40640,N_39730,N_36295);
nand U40641 (N_40641,N_30168,N_35520);
nand U40642 (N_40642,N_30113,N_36621);
nand U40643 (N_40643,N_39922,N_31912);
and U40644 (N_40644,N_34516,N_36605);
or U40645 (N_40645,N_39515,N_37965);
xnor U40646 (N_40646,N_39781,N_33399);
and U40647 (N_40647,N_34511,N_36249);
or U40648 (N_40648,N_39304,N_30288);
and U40649 (N_40649,N_33911,N_34153);
xnor U40650 (N_40650,N_39669,N_39357);
and U40651 (N_40651,N_34275,N_38997);
and U40652 (N_40652,N_38146,N_30469);
nor U40653 (N_40653,N_33630,N_35033);
nor U40654 (N_40654,N_35353,N_31030);
nand U40655 (N_40655,N_30728,N_36565);
and U40656 (N_40656,N_37496,N_30924);
xnor U40657 (N_40657,N_36278,N_31905);
xnor U40658 (N_40658,N_38774,N_35910);
nor U40659 (N_40659,N_35840,N_32350);
or U40660 (N_40660,N_32754,N_37931);
or U40661 (N_40661,N_39310,N_33256);
and U40662 (N_40662,N_32087,N_35177);
nand U40663 (N_40663,N_34409,N_33712);
nand U40664 (N_40664,N_37813,N_37278);
nor U40665 (N_40665,N_36728,N_38616);
xor U40666 (N_40666,N_32443,N_31754);
xnor U40667 (N_40667,N_32210,N_33398);
nand U40668 (N_40668,N_38770,N_34926);
xnor U40669 (N_40669,N_39282,N_30048);
or U40670 (N_40670,N_30532,N_37003);
nor U40671 (N_40671,N_37807,N_36500);
nor U40672 (N_40672,N_39136,N_34693);
or U40673 (N_40673,N_31819,N_30237);
xnor U40674 (N_40674,N_35943,N_31377);
or U40675 (N_40675,N_36968,N_39772);
or U40676 (N_40676,N_39241,N_37765);
nand U40677 (N_40677,N_33982,N_32615);
nand U40678 (N_40678,N_31980,N_37870);
xor U40679 (N_40679,N_31732,N_34981);
and U40680 (N_40680,N_39283,N_31560);
and U40681 (N_40681,N_34151,N_31076);
nand U40682 (N_40682,N_39199,N_37280);
xor U40683 (N_40683,N_36851,N_31063);
or U40684 (N_40684,N_37046,N_32412);
nand U40685 (N_40685,N_37764,N_34611);
xnor U40686 (N_40686,N_32273,N_30361);
and U40687 (N_40687,N_33910,N_34010);
nand U40688 (N_40688,N_34573,N_39340);
or U40689 (N_40689,N_30936,N_32899);
xor U40690 (N_40690,N_30920,N_35024);
xor U40691 (N_40691,N_36844,N_32765);
nor U40692 (N_40692,N_36541,N_37135);
and U40693 (N_40693,N_30762,N_39294);
nand U40694 (N_40694,N_30337,N_38618);
xor U40695 (N_40695,N_37070,N_37978);
or U40696 (N_40696,N_35159,N_34854);
nor U40697 (N_40697,N_36975,N_32919);
nand U40698 (N_40698,N_30965,N_36567);
xor U40699 (N_40699,N_34687,N_33637);
nand U40700 (N_40700,N_36221,N_31161);
and U40701 (N_40701,N_34546,N_33723);
or U40702 (N_40702,N_35173,N_34513);
or U40703 (N_40703,N_33574,N_34533);
and U40704 (N_40704,N_37442,N_32015);
xnor U40705 (N_40705,N_30716,N_36653);
nor U40706 (N_40706,N_31450,N_35695);
xor U40707 (N_40707,N_31084,N_36239);
nand U40708 (N_40708,N_37566,N_33686);
or U40709 (N_40709,N_39171,N_35245);
xnor U40710 (N_40710,N_37027,N_34590);
and U40711 (N_40711,N_39491,N_33657);
nor U40712 (N_40712,N_35645,N_39219);
nand U40713 (N_40713,N_35045,N_39653);
nor U40714 (N_40714,N_39754,N_39724);
xor U40715 (N_40715,N_37551,N_31174);
or U40716 (N_40716,N_34458,N_39774);
or U40717 (N_40717,N_30330,N_33126);
nor U40718 (N_40718,N_36686,N_39792);
nor U40719 (N_40719,N_37544,N_37036);
xor U40720 (N_40720,N_33484,N_34072);
nor U40721 (N_40721,N_33869,N_31715);
xnor U40722 (N_40722,N_32488,N_38648);
nand U40723 (N_40723,N_32739,N_31518);
or U40724 (N_40724,N_31788,N_33198);
and U40725 (N_40725,N_37633,N_32544);
nand U40726 (N_40726,N_33051,N_38170);
or U40727 (N_40727,N_35755,N_35688);
and U40728 (N_40728,N_34213,N_34857);
xnor U40729 (N_40729,N_38879,N_38002);
nor U40730 (N_40730,N_39748,N_32056);
nand U40731 (N_40731,N_36454,N_36109);
nand U40732 (N_40732,N_31026,N_35258);
nor U40733 (N_40733,N_39063,N_36576);
or U40734 (N_40734,N_30788,N_36920);
nor U40735 (N_40735,N_32427,N_31020);
or U40736 (N_40736,N_39198,N_31784);
nand U40737 (N_40737,N_34980,N_32939);
xnor U40738 (N_40738,N_37491,N_32344);
nand U40739 (N_40739,N_30461,N_35149);
and U40740 (N_40740,N_33585,N_32355);
xor U40741 (N_40741,N_37393,N_33116);
xnor U40742 (N_40742,N_33902,N_31380);
nor U40743 (N_40743,N_35411,N_31646);
or U40744 (N_40744,N_37249,N_30539);
and U40745 (N_40745,N_35040,N_38457);
nor U40746 (N_40746,N_31455,N_37117);
and U40747 (N_40747,N_35279,N_37067);
and U40748 (N_40748,N_35067,N_30444);
nand U40749 (N_40749,N_30422,N_35504);
nand U40750 (N_40750,N_39174,N_33343);
xnor U40751 (N_40751,N_35549,N_36848);
or U40752 (N_40752,N_36771,N_32418);
and U40753 (N_40753,N_30302,N_36582);
xor U40754 (N_40754,N_36633,N_31098);
nor U40755 (N_40755,N_33664,N_39787);
nor U40756 (N_40756,N_38325,N_39666);
or U40757 (N_40757,N_38542,N_38614);
nor U40758 (N_40758,N_31388,N_32692);
and U40759 (N_40759,N_37287,N_37763);
or U40760 (N_40760,N_34568,N_33550);
xor U40761 (N_40761,N_34424,N_38021);
xnor U40762 (N_40762,N_37140,N_31671);
nor U40763 (N_40763,N_34495,N_33886);
nand U40764 (N_40764,N_32454,N_34081);
or U40765 (N_40765,N_30866,N_39029);
xnor U40766 (N_40766,N_37451,N_38279);
or U40767 (N_40767,N_34307,N_35298);
nand U40768 (N_40768,N_31285,N_33276);
or U40769 (N_40769,N_34411,N_38940);
and U40770 (N_40770,N_39776,N_38506);
nand U40771 (N_40771,N_38202,N_34251);
or U40772 (N_40772,N_33336,N_34050);
and U40773 (N_40773,N_36864,N_33958);
xor U40774 (N_40774,N_38693,N_38138);
nor U40775 (N_40775,N_30879,N_30201);
xnor U40776 (N_40776,N_30313,N_30957);
nor U40777 (N_40777,N_34479,N_39587);
or U40778 (N_40778,N_33429,N_32879);
xnor U40779 (N_40779,N_33497,N_36595);
and U40780 (N_40780,N_35112,N_39239);
and U40781 (N_40781,N_37475,N_31232);
xnor U40782 (N_40782,N_32270,N_37182);
or U40783 (N_40783,N_33648,N_37501);
xnor U40784 (N_40784,N_39374,N_38526);
nand U40785 (N_40785,N_38287,N_31540);
nand U40786 (N_40786,N_38373,N_34064);
xnor U40787 (N_40787,N_34575,N_38599);
nor U40788 (N_40788,N_33439,N_31773);
nor U40789 (N_40789,N_34076,N_39033);
and U40790 (N_40790,N_38462,N_35841);
or U40791 (N_40791,N_39807,N_37397);
and U40792 (N_40792,N_35341,N_37741);
nor U40793 (N_40793,N_32213,N_33264);
nor U40794 (N_40794,N_33511,N_36992);
nor U40795 (N_40795,N_36581,N_31195);
and U40796 (N_40796,N_35489,N_34680);
or U40797 (N_40797,N_38617,N_31228);
and U40798 (N_40798,N_35735,N_31508);
or U40799 (N_40799,N_38230,N_37347);
nand U40800 (N_40800,N_38675,N_39665);
nand U40801 (N_40801,N_38140,N_37658);
nand U40802 (N_40802,N_38466,N_39055);
and U40803 (N_40803,N_38178,N_38400);
and U40804 (N_40804,N_35531,N_33662);
and U40805 (N_40805,N_35169,N_33633);
and U40806 (N_40806,N_33595,N_35933);
nor U40807 (N_40807,N_38905,N_36387);
or U40808 (N_40808,N_36035,N_38972);
xor U40809 (N_40809,N_31425,N_30634);
and U40810 (N_40810,N_32724,N_35409);
nor U40811 (N_40811,N_37708,N_37991);
and U40812 (N_40812,N_33689,N_32256);
nand U40813 (N_40813,N_32734,N_37349);
or U40814 (N_40814,N_37430,N_38129);
nand U40815 (N_40815,N_39615,N_35187);
or U40816 (N_40816,N_31951,N_37974);
nand U40817 (N_40817,N_34491,N_30410);
nor U40818 (N_40818,N_31712,N_39077);
and U40819 (N_40819,N_39813,N_35790);
nand U40820 (N_40820,N_36111,N_39227);
xnor U40821 (N_40821,N_33615,N_38576);
and U40822 (N_40822,N_35419,N_30833);
or U40823 (N_40823,N_39129,N_35492);
or U40824 (N_40824,N_38125,N_37233);
nand U40825 (N_40825,N_39633,N_30207);
or U40826 (N_40826,N_30966,N_34178);
and U40827 (N_40827,N_34422,N_32167);
xor U40828 (N_40828,N_38085,N_34176);
xor U40829 (N_40829,N_39493,N_32007);
or U40830 (N_40830,N_39108,N_30058);
xor U40831 (N_40831,N_37727,N_36829);
or U40832 (N_40832,N_39257,N_35815);
nor U40833 (N_40833,N_36781,N_36699);
nor U40834 (N_40834,N_38739,N_34116);
xnor U40835 (N_40835,N_30417,N_34206);
xnor U40836 (N_40836,N_31859,N_31181);
nor U40837 (N_40837,N_30652,N_34201);
xor U40838 (N_40838,N_33096,N_36880);
or U40839 (N_40839,N_31268,N_39589);
or U40840 (N_40840,N_30743,N_34911);
nor U40841 (N_40841,N_38857,N_39215);
and U40842 (N_40842,N_39041,N_35008);
and U40843 (N_40843,N_33374,N_39296);
or U40844 (N_40844,N_33944,N_34390);
nor U40845 (N_40845,N_34262,N_36179);
or U40846 (N_40846,N_32969,N_38214);
and U40847 (N_40847,N_35784,N_39002);
or U40848 (N_40848,N_37245,N_31823);
nor U40849 (N_40849,N_37587,N_38715);
and U40850 (N_40850,N_34622,N_39715);
nand U40851 (N_40851,N_32990,N_34278);
xor U40852 (N_40852,N_34005,N_37291);
and U40853 (N_40853,N_39769,N_32286);
nor U40854 (N_40854,N_37902,N_30486);
and U40855 (N_40855,N_38802,N_36121);
nor U40856 (N_40856,N_34381,N_31176);
nor U40857 (N_40857,N_31378,N_36177);
nand U40858 (N_40858,N_39609,N_30038);
xor U40859 (N_40859,N_35862,N_32710);
or U40860 (N_40860,N_39149,N_30837);
nor U40861 (N_40861,N_35847,N_30850);
and U40862 (N_40862,N_38012,N_33746);
or U40863 (N_40863,N_33692,N_38579);
nor U40864 (N_40864,N_38116,N_36155);
and U40865 (N_40865,N_31598,N_38964);
or U40866 (N_40866,N_31534,N_34193);
and U40867 (N_40867,N_37545,N_37690);
nor U40868 (N_40868,N_35710,N_32570);
nor U40869 (N_40869,N_35054,N_35163);
xor U40870 (N_40870,N_30082,N_31005);
xnor U40871 (N_40871,N_31820,N_31458);
or U40872 (N_40872,N_31362,N_36947);
xor U40873 (N_40873,N_30608,N_35237);
xnor U40874 (N_40874,N_35556,N_30801);
or U40875 (N_40875,N_34625,N_39652);
nand U40876 (N_40876,N_33344,N_35788);
xor U40877 (N_40877,N_32828,N_32546);
and U40878 (N_40878,N_38097,N_32906);
nand U40879 (N_40879,N_30968,N_38458);
or U40880 (N_40880,N_32391,N_36051);
xor U40881 (N_40881,N_31364,N_35413);
nor U40882 (N_40882,N_32159,N_36933);
and U40883 (N_40883,N_33569,N_33734);
nor U40884 (N_40884,N_30882,N_38417);
xor U40885 (N_40885,N_30639,N_33770);
xor U40886 (N_40886,N_31281,N_37100);
and U40887 (N_40887,N_30475,N_33631);
nor U40888 (N_40888,N_30377,N_39601);
nor U40889 (N_40889,N_36219,N_38258);
or U40890 (N_40890,N_35046,N_30946);
nand U40891 (N_40891,N_34164,N_38193);
or U40892 (N_40892,N_33589,N_33565);
nand U40893 (N_40893,N_36224,N_30511);
nor U40894 (N_40894,N_32881,N_36485);
or U40895 (N_40895,N_32310,N_31931);
nor U40896 (N_40896,N_38018,N_33025);
and U40897 (N_40897,N_30584,N_31783);
and U40898 (N_40898,N_32069,N_36591);
or U40899 (N_40899,N_35209,N_37645);
xnor U40900 (N_40900,N_39036,N_38040);
or U40901 (N_40901,N_35678,N_32907);
or U40902 (N_40902,N_39561,N_38039);
xnor U40903 (N_40903,N_38769,N_33695);
nand U40904 (N_40904,N_36072,N_38952);
or U40905 (N_40905,N_39235,N_34074);
or U40906 (N_40906,N_37463,N_33673);
or U40907 (N_40907,N_31060,N_39090);
xnor U40908 (N_40908,N_35382,N_31149);
xor U40909 (N_40909,N_39918,N_39679);
or U40910 (N_40910,N_33099,N_37680);
nand U40911 (N_40911,N_39820,N_35447);
or U40912 (N_40912,N_32751,N_37543);
and U40913 (N_40913,N_31763,N_34431);
xor U40914 (N_40914,N_39339,N_31357);
or U40915 (N_40915,N_33803,N_35412);
xor U40916 (N_40916,N_38498,N_36008);
nor U40917 (N_40917,N_34636,N_33114);
nor U40918 (N_40918,N_34366,N_34354);
or U40919 (N_40919,N_31510,N_30569);
or U40920 (N_40920,N_35009,N_39983);
nand U40921 (N_40921,N_34452,N_34819);
or U40922 (N_40922,N_31664,N_37301);
xnor U40923 (N_40923,N_39997,N_32851);
or U40924 (N_40924,N_37257,N_32481);
nor U40925 (N_40925,N_35713,N_35165);
and U40926 (N_40926,N_33338,N_33954);
or U40927 (N_40927,N_33596,N_32036);
nand U40928 (N_40928,N_33005,N_31704);
nor U40929 (N_40929,N_39713,N_32325);
nand U40930 (N_40930,N_36584,N_34257);
nor U40931 (N_40931,N_38365,N_35141);
nor U40932 (N_40932,N_33403,N_33085);
nand U40933 (N_40933,N_34966,N_37403);
nand U40934 (N_40934,N_36375,N_39190);
or U40935 (N_40935,N_32605,N_34758);
xor U40936 (N_40936,N_35205,N_32988);
nor U40937 (N_40937,N_38160,N_36602);
and U40938 (N_40938,N_34416,N_30365);
nor U40939 (N_40939,N_36598,N_32368);
xnor U40940 (N_40940,N_39278,N_30854);
nand U40941 (N_40941,N_32018,N_31802);
nor U40942 (N_40942,N_30154,N_34032);
or U40943 (N_40943,N_35985,N_36997);
nor U40944 (N_40944,N_31950,N_31509);
or U40945 (N_40945,N_30689,N_38612);
xor U40946 (N_40946,N_39197,N_37772);
xor U40947 (N_40947,N_36393,N_30699);
or U40948 (N_40948,N_39642,N_39267);
and U40949 (N_40949,N_37017,N_31352);
nor U40950 (N_40950,N_32314,N_35576);
nand U40951 (N_40951,N_34274,N_38783);
or U40952 (N_40952,N_39058,N_39109);
xnor U40953 (N_40953,N_30277,N_36191);
xnor U40954 (N_40954,N_39853,N_39726);
nand U40955 (N_40955,N_30687,N_32948);
xor U40956 (N_40956,N_31595,N_35191);
nor U40957 (N_40957,N_31869,N_33390);
nand U40958 (N_40958,N_35071,N_34814);
xor U40959 (N_40959,N_30858,N_34156);
or U40960 (N_40960,N_36037,N_39003);
and U40961 (N_40961,N_30298,N_30826);
or U40962 (N_40962,N_32209,N_36619);
nand U40963 (N_40963,N_33903,N_30106);
nor U40964 (N_40964,N_38883,N_32728);
and U40965 (N_40965,N_35204,N_37273);
nor U40966 (N_40966,N_34448,N_33623);
nor U40967 (N_40967,N_37926,N_31919);
and U40968 (N_40968,N_32648,N_38382);
nand U40969 (N_40969,N_38250,N_35611);
xnor U40970 (N_40970,N_30384,N_30597);
nand U40971 (N_40971,N_35624,N_38104);
and U40972 (N_40972,N_31528,N_30233);
nand U40973 (N_40973,N_36389,N_34329);
and U40974 (N_40974,N_38959,N_30963);
and U40975 (N_40975,N_35820,N_32413);
or U40976 (N_40976,N_30913,N_30508);
nand U40977 (N_40977,N_36166,N_35296);
or U40978 (N_40978,N_30981,N_30811);
nand U40979 (N_40979,N_33007,N_32846);
and U40980 (N_40980,N_32671,N_34498);
xnor U40981 (N_40981,N_32105,N_31185);
nand U40982 (N_40982,N_30992,N_38402);
nor U40983 (N_40983,N_38237,N_33045);
nor U40984 (N_40984,N_33211,N_33044);
or U40985 (N_40985,N_33132,N_35921);
or U40986 (N_40986,N_33433,N_33769);
nor U40987 (N_40987,N_34289,N_39958);
and U40988 (N_40988,N_39485,N_35750);
nor U40989 (N_40989,N_32250,N_36657);
nand U40990 (N_40990,N_36666,N_39512);
and U40991 (N_40991,N_31328,N_33894);
or U40992 (N_40992,N_37605,N_31008);
and U40993 (N_40993,N_31947,N_31719);
nor U40994 (N_40994,N_32294,N_30610);
or U40995 (N_40995,N_31134,N_39795);
nand U40996 (N_40996,N_30370,N_33580);
or U40997 (N_40997,N_37388,N_30134);
and U40998 (N_40998,N_39121,N_36467);
xnor U40999 (N_40999,N_37269,N_32642);
xor U41000 (N_41000,N_30501,N_31476);
and U41001 (N_41001,N_39275,N_31258);
xnor U41002 (N_41002,N_32046,N_36416);
nor U41003 (N_41003,N_31736,N_35733);
nand U41004 (N_41004,N_35186,N_37520);
nor U41005 (N_41005,N_38522,N_39051);
nor U41006 (N_41006,N_35042,N_35836);
nand U41007 (N_41007,N_31847,N_35208);
or U41008 (N_41008,N_33420,N_37113);
and U41009 (N_41009,N_35950,N_38583);
xor U41010 (N_41010,N_36381,N_32872);
nand U41011 (N_41011,N_32030,N_33389);
or U41012 (N_41012,N_31500,N_37922);
and U41013 (N_41013,N_31080,N_38932);
or U41014 (N_41014,N_31169,N_30232);
xnor U41015 (N_41015,N_37848,N_36867);
nand U41016 (N_41016,N_30057,N_36490);
or U41017 (N_41017,N_38020,N_32970);
or U41018 (N_41018,N_33345,N_33069);
xor U41019 (N_41019,N_34472,N_35103);
and U41020 (N_41020,N_32535,N_30085);
and U41021 (N_41021,N_32262,N_38733);
nand U41022 (N_41022,N_30899,N_33908);
or U41023 (N_41023,N_33540,N_32238);
xnor U41024 (N_41024,N_31609,N_36477);
or U41025 (N_41025,N_38035,N_31222);
and U41026 (N_41026,N_38889,N_35528);
xnor U41027 (N_41027,N_31619,N_37950);
or U41028 (N_41028,N_34909,N_35823);
xor U41029 (N_41029,N_39490,N_31471);
nor U41030 (N_41030,N_32060,N_35174);
or U41031 (N_41031,N_33948,N_37707);
nor U41032 (N_41032,N_30581,N_38476);
nand U41033 (N_41033,N_39691,N_35667);
nor U41034 (N_41034,N_34004,N_31963);
or U41035 (N_41035,N_37051,N_33531);
nand U41036 (N_41036,N_36018,N_37455);
xor U41037 (N_41037,N_33707,N_37376);
nand U41038 (N_41038,N_30662,N_35281);
xnor U41039 (N_41039,N_36793,N_35843);
and U41040 (N_41040,N_30681,N_36363);
and U41041 (N_41041,N_37976,N_30873);
xor U41042 (N_41042,N_39976,N_33231);
and U41043 (N_41043,N_35432,N_32955);
nand U41044 (N_41044,N_34784,N_34267);
or U41045 (N_41045,N_36283,N_31111);
and U41046 (N_41046,N_36524,N_34951);
or U41047 (N_41047,N_31284,N_34174);
nand U41048 (N_41048,N_37738,N_32696);
nand U41049 (N_41049,N_31696,N_32914);
xnor U41050 (N_41050,N_35839,N_31191);
or U41051 (N_41051,N_33259,N_36701);
xor U41052 (N_41052,N_31132,N_35670);
nand U41053 (N_41053,N_37599,N_36305);
or U41054 (N_41054,N_37852,N_39854);
nor U41055 (N_41055,N_37216,N_32915);
nor U41056 (N_41056,N_39154,N_32121);
nand U41057 (N_41057,N_32643,N_30719);
or U41058 (N_41058,N_37527,N_38823);
and U41059 (N_41059,N_38141,N_38378);
nand U41060 (N_41060,N_39187,N_39320);
or U41061 (N_41061,N_33036,N_36881);
xnor U41062 (N_41062,N_30734,N_37304);
xnor U41063 (N_41063,N_32360,N_30588);
nor U41064 (N_41064,N_37760,N_39681);
xnor U41065 (N_41065,N_37071,N_31325);
nand U41066 (N_41066,N_38661,N_38067);
or U41067 (N_41067,N_33710,N_33647);
nand U41068 (N_41068,N_32375,N_38707);
or U41069 (N_41069,N_36030,N_34853);
xnor U41070 (N_41070,N_35569,N_34442);
and U41071 (N_41071,N_32865,N_34047);
nand U41072 (N_41072,N_34564,N_35010);
nand U41073 (N_41073,N_38716,N_33458);
and U41074 (N_41074,N_37427,N_37712);
or U41075 (N_41075,N_39391,N_35679);
and U41076 (N_41076,N_34954,N_34309);
nand U41077 (N_41077,N_30698,N_36211);
nand U41078 (N_41078,N_31636,N_36168);
and U41079 (N_41079,N_33775,N_34595);
and U41080 (N_41080,N_30143,N_37607);
nor U41081 (N_41081,N_39523,N_34727);
or U41082 (N_41082,N_32725,N_38353);
or U41083 (N_41083,N_35949,N_38235);
and U41084 (N_41084,N_34579,N_31953);
xor U41085 (N_41085,N_38943,N_30240);
and U41086 (N_41086,N_32746,N_38562);
nand U41087 (N_41087,N_38649,N_31442);
or U41088 (N_41088,N_35709,N_34022);
xor U41089 (N_41089,N_31194,N_39302);
xnor U41090 (N_41090,N_31607,N_34484);
and U41091 (N_41091,N_34095,N_38113);
nor U41092 (N_41092,N_37370,N_34733);
xnor U41093 (N_41093,N_34230,N_30121);
and U41094 (N_41094,N_32165,N_35608);
nor U41095 (N_41095,N_34776,N_31575);
nor U41096 (N_41096,N_37559,N_39175);
or U41097 (N_41097,N_32526,N_31189);
xor U41098 (N_41098,N_34702,N_36207);
nand U41099 (N_41099,N_32674,N_34816);
and U41100 (N_41100,N_32293,N_37088);
xor U41101 (N_41101,N_33753,N_35658);
xor U41102 (N_41102,N_30636,N_37081);
and U41103 (N_41103,N_36366,N_35774);
or U41104 (N_41104,N_30066,N_30861);
and U41105 (N_41105,N_39383,N_38786);
and U41106 (N_41106,N_37784,N_35247);
and U41107 (N_41107,N_33255,N_37715);
and U41108 (N_41108,N_36466,N_31675);
or U41109 (N_41109,N_33376,N_36668);
xor U41110 (N_41110,N_34463,N_34556);
or U41111 (N_41111,N_31154,N_35766);
xnor U41112 (N_41112,N_36400,N_34369);
nor U41113 (N_41113,N_37382,N_33450);
or U41114 (N_41114,N_38063,N_37854);
or U41115 (N_41115,N_32631,N_30579);
xor U41116 (N_41116,N_30790,N_32278);
nand U41117 (N_41117,N_31968,N_35349);
and U41118 (N_41118,N_37228,N_39550);
nor U41119 (N_41119,N_38071,N_35120);
nor U41120 (N_41120,N_32797,N_34536);
and U41121 (N_41121,N_33363,N_38183);
or U41122 (N_41122,N_30935,N_30116);
nor U41123 (N_41123,N_38608,N_31790);
xnor U41124 (N_41124,N_38862,N_34147);
nor U41125 (N_41125,N_36041,N_31625);
nand U41126 (N_41126,N_37299,N_36498);
xnor U41127 (N_41127,N_35798,N_31612);
nor U41128 (N_41128,N_31808,N_38929);
xor U41129 (N_41129,N_36761,N_31256);
and U41130 (N_41130,N_39883,N_33407);
nand U41131 (N_41131,N_31199,N_31882);
and U41132 (N_41132,N_38765,N_35126);
and U41133 (N_41133,N_36641,N_33870);
nor U41134 (N_41134,N_37990,N_35879);
nand U41135 (N_41135,N_32709,N_39252);
or U41136 (N_41136,N_32741,N_35377);
nor U41137 (N_41137,N_35166,N_31177);
or U41138 (N_41138,N_33665,N_31881);
and U41139 (N_41139,N_35589,N_31812);
or U41140 (N_41140,N_31720,N_30037);
and U41141 (N_41141,N_32088,N_37616);
or U41142 (N_41142,N_33104,N_30628);
and U41143 (N_41143,N_30729,N_34991);
xor U41144 (N_41144,N_38568,N_37057);
and U41145 (N_41145,N_39132,N_32722);
or U41146 (N_41146,N_38662,N_37942);
and U41147 (N_41147,N_33129,N_30761);
and U41148 (N_41148,N_34090,N_31811);
and U41149 (N_41149,N_39815,N_33601);
nor U41150 (N_41150,N_34292,N_35384);
and U41151 (N_41151,N_32838,N_34874);
xnor U41152 (N_41152,N_36294,N_30183);
and U41153 (N_41153,N_36789,N_36282);
xor U41154 (N_41154,N_35020,N_36025);
or U41155 (N_41155,N_38451,N_30509);
and U41156 (N_41156,N_36780,N_35853);
or U41157 (N_41157,N_39686,N_36209);
nand U41158 (N_41158,N_39196,N_32982);
nand U41159 (N_41159,N_37622,N_33379);
nand U41160 (N_41160,N_34143,N_37981);
nand U41161 (N_41161,N_35015,N_38697);
xnor U41162 (N_41162,N_35438,N_35392);
or U41163 (N_41163,N_38831,N_35942);
or U41164 (N_41164,N_31590,N_30347);
or U41165 (N_41165,N_34649,N_35998);
or U41166 (N_41166,N_32379,N_36847);
or U41167 (N_41167,N_31123,N_38567);
nand U41168 (N_41168,N_38584,N_33023);
nand U41169 (N_41169,N_36794,N_30339);
and U41170 (N_41170,N_33891,N_30504);
nand U41171 (N_41171,N_35869,N_30732);
or U41172 (N_41172,N_38004,N_30725);
nor U41173 (N_41173,N_30541,N_37711);
or U41174 (N_41174,N_32567,N_34232);
nand U41175 (N_41175,N_36832,N_39432);
or U41176 (N_41176,N_34197,N_30623);
xor U41177 (N_41177,N_35211,N_39955);
or U41178 (N_41178,N_34402,N_37834);
nand U41179 (N_41179,N_34713,N_32264);
nand U41180 (N_41180,N_30671,N_34119);
and U41181 (N_41181,N_38577,N_38848);
nand U41182 (N_41182,N_38725,N_34017);
xnor U41183 (N_41183,N_33050,N_38312);
nor U41184 (N_41184,N_30454,N_38336);
xor U41185 (N_41185,N_37142,N_33155);
xor U41186 (N_41186,N_34195,N_39091);
xor U41187 (N_41187,N_32070,N_34848);
and U41188 (N_41188,N_32027,N_31585);
nand U41189 (N_41189,N_33679,N_32033);
and U41190 (N_41190,N_39079,N_37001);
nand U41191 (N_41191,N_32613,N_32924);
nor U41192 (N_41192,N_34367,N_34634);
nor U41193 (N_41193,N_37016,N_38863);
nand U41194 (N_41194,N_31605,N_37925);
or U41195 (N_41195,N_39851,N_34982);
nand U41196 (N_41196,N_36969,N_36869);
xnor U41197 (N_41197,N_30856,N_36813);
xor U41198 (N_41198,N_33113,N_35922);
or U41199 (N_41199,N_35502,N_30731);
nand U41200 (N_41200,N_32330,N_34322);
nand U41201 (N_41201,N_32818,N_33584);
nand U41202 (N_41202,N_34497,N_30587);
nand U41203 (N_41203,N_34526,N_32867);
nor U41204 (N_41204,N_34815,N_39365);
and U41205 (N_41205,N_34602,N_32916);
nor U41206 (N_41206,N_35868,N_38658);
or U41207 (N_41207,N_33750,N_31103);
and U41208 (N_41208,N_33317,N_39221);
and U41209 (N_41209,N_38866,N_39333);
nand U41210 (N_41210,N_39356,N_35825);
and U41211 (N_41211,N_37361,N_38727);
or U41212 (N_41212,N_34245,N_31353);
or U41213 (N_41213,N_36090,N_33165);
and U41214 (N_41214,N_35483,N_34939);
or U41215 (N_41215,N_30985,N_38885);
and U41216 (N_41216,N_35909,N_35132);
or U41217 (N_41217,N_39440,N_30835);
nand U41218 (N_41218,N_38105,N_38314);
or U41219 (N_41219,N_35185,N_36169);
and U41220 (N_41220,N_38667,N_35964);
and U41221 (N_41221,N_31106,N_31724);
xor U41222 (N_41222,N_31961,N_37037);
nor U41223 (N_41223,N_32579,N_35982);
nand U41224 (N_41224,N_37255,N_36288);
and U41225 (N_41225,N_36418,N_32656);
nor U41226 (N_41226,N_36099,N_35972);
nor U41227 (N_41227,N_37904,N_39937);
nand U41228 (N_41228,N_35181,N_38163);
nand U41229 (N_41229,N_35595,N_34852);
nand U41230 (N_41230,N_36320,N_37008);
nor U41231 (N_41231,N_32801,N_38712);
nor U41232 (N_41232,N_34929,N_32832);
or U41233 (N_41233,N_34557,N_38784);
nor U41234 (N_41234,N_35025,N_37649);
nand U41235 (N_41235,N_30251,N_38159);
nand U41236 (N_41236,N_34352,N_30792);
or U41237 (N_41237,N_38061,N_35358);
or U41238 (N_41238,N_34485,N_35712);
xor U41239 (N_41239,N_34534,N_32162);
and U41240 (N_41240,N_34865,N_33011);
or U41241 (N_41241,N_37481,N_37567);
or U41242 (N_41242,N_37390,N_37426);
nor U41243 (N_41243,N_31395,N_38263);
or U41244 (N_41244,N_35979,N_30089);
nor U41245 (N_41245,N_37192,N_32819);
xnor U41246 (N_41246,N_36528,N_30180);
and U41247 (N_41247,N_36688,N_39351);
or U41248 (N_41248,N_31800,N_39107);
nor U41249 (N_41249,N_32207,N_36929);
nor U41250 (N_41250,N_38277,N_36419);
and U41251 (N_41251,N_35352,N_39804);
or U41252 (N_41252,N_32322,N_38273);
xor U41253 (N_41253,N_39470,N_31555);
or U41254 (N_41254,N_30783,N_31801);
nor U41255 (N_41255,N_32035,N_37610);
nand U41256 (N_41256,N_34070,N_36730);
xor U41257 (N_41257,N_32809,N_32864);
nand U41258 (N_41258,N_34380,N_31731);
and U41259 (N_41259,N_38322,N_35523);
or U41260 (N_41260,N_32425,N_39242);
or U41261 (N_41261,N_39635,N_32635);
and U41262 (N_41262,N_30360,N_30006);
and U41263 (N_41263,N_30368,N_35677);
nor U41264 (N_41264,N_38502,N_36977);
nand U41265 (N_41265,N_39138,N_31055);
xnor U41266 (N_41266,N_30883,N_33008);
nor U41267 (N_41267,N_31863,N_32483);
or U41268 (N_41268,N_31681,N_31403);
nor U41269 (N_41269,N_39455,N_32371);
and U41270 (N_41270,N_33552,N_33434);
xor U41271 (N_41271,N_37739,N_32667);
nand U41272 (N_41272,N_35818,N_33143);
and U41273 (N_41273,N_34096,N_36459);
nor U41274 (N_41274,N_37993,N_34025);
or U41275 (N_41275,N_33731,N_34900);
nor U41276 (N_41276,N_35224,N_37819);
nor U41277 (N_41277,N_32420,N_35914);
or U41278 (N_41278,N_30970,N_32373);
or U41279 (N_41279,N_30808,N_36311);
xnor U41280 (N_41280,N_33493,N_32673);
xnor U41281 (N_41281,N_37341,N_38100);
xnor U41282 (N_41282,N_31140,N_30265);
xnor U41283 (N_41283,N_30979,N_36769);
nand U41284 (N_41284,N_33549,N_33767);
and U41285 (N_41285,N_38064,N_36693);
xor U41286 (N_41286,N_36695,N_33057);
nor U41287 (N_41287,N_36564,N_39599);
xor U41288 (N_41288,N_30159,N_34800);
and U41289 (N_41289,N_38993,N_39957);
or U41290 (N_41290,N_32775,N_37406);
nand U41291 (N_41291,N_33566,N_36819);
and U41292 (N_41292,N_30211,N_33807);
and U41293 (N_41293,N_37217,N_32856);
nand U41294 (N_41294,N_33232,N_37890);
xor U41295 (N_41295,N_33238,N_35153);
and U41296 (N_41296,N_38575,N_34286);
nand U41297 (N_41297,N_38194,N_37354);
or U41298 (N_41298,N_37206,N_36413);
nand U41299 (N_41299,N_39661,N_32093);
and U41300 (N_41300,N_37818,N_34224);
xor U41301 (N_41301,N_32581,N_39771);
or U41302 (N_41302,N_35094,N_36909);
xor U41303 (N_41303,N_38604,N_38446);
or U41304 (N_41304,N_34856,N_35771);
xnor U41305 (N_41305,N_38793,N_39075);
xor U41306 (N_41306,N_34235,N_34049);
and U41307 (N_41307,N_32632,N_36684);
nand U41308 (N_41308,N_36893,N_34031);
nand U41309 (N_41309,N_30070,N_31062);
and U41310 (N_41310,N_34438,N_34127);
and U41311 (N_41311,N_30407,N_35139);
nand U41312 (N_41312,N_31128,N_37264);
and U41313 (N_41313,N_34287,N_37314);
or U41314 (N_41314,N_30386,N_34872);
nor U41315 (N_41315,N_34148,N_35193);
nor U41316 (N_41316,N_33779,N_36750);
nor U41317 (N_41317,N_31606,N_39114);
and U41318 (N_41318,N_37212,N_34000);
nand U41319 (N_41319,N_30606,N_30857);
xnor U41320 (N_41320,N_39127,N_36313);
and U41321 (N_41321,N_34211,N_35452);
nor U41322 (N_41322,N_35035,N_37108);
nor U41323 (N_41323,N_35714,N_34890);
and U41324 (N_41324,N_35988,N_31401);
xor U41325 (N_41325,N_31021,N_31365);
nand U41326 (N_41326,N_38371,N_36031);
nand U41327 (N_41327,N_37398,N_30403);
nor U41328 (N_41328,N_33391,N_38761);
nand U41329 (N_41329,N_35685,N_37157);
xnor U41330 (N_41330,N_36013,N_33713);
or U41331 (N_41331,N_35363,N_34749);
and U41332 (N_41332,N_35408,N_31851);
nor U41333 (N_41333,N_32557,N_32460);
or U41334 (N_41334,N_32348,N_32320);
nor U41335 (N_41335,N_37793,N_35501);
or U41336 (N_41336,N_36898,N_37078);
nand U41337 (N_41337,N_38771,N_36770);
nor U41338 (N_41338,N_30614,N_34248);
or U41339 (N_41339,N_31190,N_33646);
xnor U41340 (N_41340,N_37166,N_35830);
nor U41341 (N_41341,N_39466,N_32861);
nand U41342 (N_41342,N_34519,N_35622);
or U41343 (N_41343,N_35479,N_39048);
xnor U41344 (N_41344,N_38320,N_36719);
nor U41345 (N_41345,N_31155,N_37395);
nor U41346 (N_41346,N_32857,N_30998);
xor U41347 (N_41347,N_33199,N_34714);
and U41348 (N_41348,N_31662,N_32630);
and U41349 (N_41349,N_39210,N_36858);
and U41350 (N_41350,N_37263,N_34196);
or U41351 (N_41351,N_34443,N_37889);
nand U41352 (N_41352,N_32478,N_36631);
nor U41353 (N_41353,N_32930,N_36087);
or U41354 (N_41354,N_35366,N_36544);
and U41355 (N_41355,N_36952,N_32102);
nand U41356 (N_41356,N_33016,N_39245);
xor U41357 (N_41357,N_31764,N_30663);
nand U41358 (N_41358,N_34417,N_34983);
and U41359 (N_41359,N_33229,N_38300);
nor U41360 (N_41360,N_34708,N_33110);
and U41361 (N_41361,N_31217,N_32542);
nor U41362 (N_41362,N_31663,N_34217);
xnor U41363 (N_41363,N_31399,N_39693);
xor U41364 (N_41364,N_38681,N_38090);
nor U41365 (N_41365,N_38056,N_38075);
xnor U41366 (N_41366,N_39902,N_37237);
xnor U41367 (N_41367,N_31780,N_37535);
or U41368 (N_41368,N_33191,N_33805);
and U41369 (N_41369,N_38225,N_35050);
nor U41370 (N_41370,N_33253,N_31749);
xnor U41371 (N_41371,N_35344,N_37367);
and U41372 (N_41372,N_32153,N_39146);
xnor U41373 (N_41373,N_31730,N_32884);
and U41374 (N_41374,N_37591,N_34179);
nor U41375 (N_41375,N_39700,N_33771);
and U41376 (N_41376,N_30897,N_39732);
xor U41377 (N_41377,N_31104,N_37909);
nand U41378 (N_41378,N_38556,N_30012);
nand U41379 (N_41379,N_38078,N_36378);
and U41380 (N_41380,N_33841,N_35246);
and U41381 (N_41381,N_37209,N_33157);
nor U41382 (N_41382,N_35568,N_30609);
or U41383 (N_41383,N_33058,N_32192);
or U41384 (N_41384,N_34522,N_38486);
nor U41385 (N_41385,N_32713,N_38504);
and U41386 (N_41386,N_38411,N_34428);
nor U41387 (N_41387,N_35990,N_36337);
xnor U41388 (N_41388,N_35812,N_34578);
or U41389 (N_41389,N_39152,N_38102);
and U41390 (N_41390,N_30632,N_35999);
xor U41391 (N_41391,N_32830,N_33545);
and U41392 (N_41392,N_38994,N_34811);
and U41393 (N_41393,N_36593,N_31706);
and U41394 (N_41394,N_38724,N_35325);
or U41395 (N_41395,N_32231,N_35135);
and U41396 (N_41396,N_33756,N_34834);
nand U41397 (N_41397,N_38494,N_34488);
nand U41398 (N_41398,N_39761,N_34385);
nor U41399 (N_41399,N_38887,N_36713);
nand U41400 (N_41400,N_35541,N_33423);
xnor U41401 (N_41401,N_35044,N_37223);
nand U41402 (N_41402,N_32558,N_31913);
or U41403 (N_41403,N_36979,N_32530);
nand U41404 (N_41404,N_36632,N_39300);
nor U41405 (N_41405,N_32821,N_32817);
or U41406 (N_41406,N_34231,N_34603);
and U41407 (N_41407,N_30537,N_38031);
or U41408 (N_41408,N_35439,N_30869);
xnor U41409 (N_41409,N_36186,N_31537);
and U41410 (N_41410,N_31734,N_37794);
xor U41411 (N_41411,N_32575,N_34105);
nor U41412 (N_41412,N_31315,N_39327);
nor U41413 (N_41413,N_32935,N_31018);
xor U41414 (N_41414,N_37198,N_31305);
xnor U41415 (N_41415,N_36384,N_38427);
nand U41416 (N_41416,N_37825,N_31525);
nand U41417 (N_41417,N_36554,N_38588);
nor U41418 (N_41418,N_38958,N_36923);
or U41419 (N_41419,N_35817,N_39286);
xor U41420 (N_41420,N_36644,N_39901);
xnor U41421 (N_41421,N_37022,N_39067);
or U41422 (N_41422,N_32844,N_36353);
nand U41423 (N_41423,N_38781,N_39097);
and U41424 (N_41424,N_34504,N_35007);
and U41425 (N_41425,N_30398,N_32863);
or U41426 (N_41426,N_32388,N_33093);
and U41427 (N_41427,N_38449,N_34210);
nand U41428 (N_41428,N_30518,N_39848);
xor U41429 (N_41429,N_32212,N_38006);
or U41430 (N_41430,N_39382,N_31361);
nor U41431 (N_41431,N_36917,N_35219);
xnor U41432 (N_41432,N_32111,N_36279);
or U41433 (N_41433,N_35616,N_39595);
nor U41434 (N_41434,N_31946,N_38896);
and U41435 (N_41435,N_30929,N_36671);
or U41436 (N_41436,N_39780,N_30124);
xor U41437 (N_41437,N_39120,N_35406);
or U41438 (N_41438,N_32664,N_33307);
or U41439 (N_41439,N_36346,N_39346);
or U41440 (N_41440,N_30657,N_31349);
or U41441 (N_41441,N_39168,N_39859);
nor U41442 (N_41442,N_37162,N_32356);
nand U41443 (N_41443,N_37322,N_35212);
xnor U41444 (N_41444,N_35319,N_37411);
xnor U41445 (N_41445,N_39648,N_39478);
and U41446 (N_41446,N_38254,N_33425);
nand U41447 (N_41447,N_37373,N_36690);
nor U41448 (N_41448,N_34607,N_37038);
or U41449 (N_41449,N_33055,N_37174);
nor U41450 (N_41450,N_39427,N_36255);
and U41451 (N_41451,N_35499,N_31698);
xnor U41452 (N_41452,N_37723,N_33792);
nor U41453 (N_41453,N_37085,N_37988);
xnor U41454 (N_41454,N_36334,N_35544);
or U41455 (N_41455,N_38624,N_31295);
nand U41456 (N_41456,N_31889,N_37864);
nor U41457 (N_41457,N_37872,N_31368);
nand U41458 (N_41458,N_37528,N_32536);
xnor U41459 (N_41459,N_39006,N_37631);
and U41460 (N_41460,N_31344,N_35226);
nor U41461 (N_41461,N_36826,N_31554);
or U41462 (N_41462,N_35493,N_34843);
or U41463 (N_41463,N_32825,N_35833);
nor U41464 (N_41464,N_38463,N_38654);
nand U41465 (N_41465,N_30188,N_37019);
nor U41466 (N_41466,N_36577,N_38974);
or U41467 (N_41467,N_39999,N_39261);
and U41468 (N_41468,N_33706,N_31086);
or U41469 (N_41469,N_30246,N_31778);
xor U41470 (N_41470,N_31999,N_39697);
nand U41471 (N_41471,N_38933,N_38242);
or U41472 (N_41472,N_38850,N_37509);
and U41473 (N_41473,N_36866,N_31383);
or U41474 (N_41474,N_35779,N_31703);
nor U41475 (N_41475,N_35846,N_33451);
nand U41476 (N_41476,N_39892,N_30626);
or U41477 (N_41477,N_39153,N_32485);
and U41478 (N_41478,N_30834,N_39388);
and U41479 (N_41479,N_33774,N_33000);
xor U41480 (N_41480,N_38833,N_30338);
or U41481 (N_41481,N_32963,N_32061);
nand U41482 (N_41482,N_35593,N_34426);
xnor U41483 (N_41483,N_32299,N_37804);
nor U41484 (N_41484,N_35290,N_30898);
nand U41485 (N_41485,N_34372,N_33967);
nor U41486 (N_41486,N_39318,N_33997);
or U41487 (N_41487,N_35571,N_39203);
and U41488 (N_41488,N_36356,N_37254);
xor U41489 (N_41489,N_37885,N_34588);
or U41490 (N_41490,N_38790,N_39867);
nor U41491 (N_41491,N_33020,N_38945);
xor U41492 (N_41492,N_36971,N_38088);
nor U41493 (N_41493,N_36012,N_35255);
nand U41494 (N_41494,N_39043,N_36849);
or U41495 (N_41495,N_32415,N_38503);
nor U41496 (N_41496,N_37323,N_37281);
and U41497 (N_41497,N_30044,N_34945);
nor U41498 (N_41498,N_35680,N_31110);
and U41499 (N_41499,N_34960,N_31923);
or U41500 (N_41500,N_34468,N_31994);
nor U41501 (N_41501,N_36763,N_32122);
xor U41502 (N_41502,N_39690,N_30375);
and U41503 (N_41503,N_33314,N_30491);
and U41504 (N_41504,N_32358,N_36580);
or U41505 (N_41505,N_38094,N_37677);
or U41506 (N_41506,N_35484,N_35831);
nor U41507 (N_41507,N_32107,N_36513);
xor U41508 (N_41508,N_35721,N_30056);
xnor U41509 (N_41509,N_30958,N_36827);
and U41510 (N_41510,N_35090,N_32511);
xnor U41511 (N_41511,N_31439,N_37840);
and U41512 (N_41512,N_31069,N_36088);
or U41513 (N_41513,N_38842,N_37394);
nor U41514 (N_41514,N_30527,N_36340);
and U41515 (N_41515,N_39234,N_34460);
and U41516 (N_41516,N_30487,N_35761);
nand U41517 (N_41517,N_31302,N_32155);
or U41518 (N_41518,N_39366,N_35944);
and U41519 (N_41519,N_32662,N_37959);
and U41520 (N_41520,N_31623,N_32258);
nand U41521 (N_41521,N_35500,N_34739);
nor U41522 (N_41522,N_32777,N_36714);
or U41523 (N_41523,N_33937,N_33966);
and U41524 (N_41524,N_37005,N_38423);
xnor U41525 (N_41525,N_33272,N_38292);
nand U41526 (N_41526,N_39507,N_36068);
and U41527 (N_41527,N_31866,N_36372);
nand U41528 (N_41528,N_31587,N_32079);
nor U41529 (N_41529,N_35014,N_31926);
xor U41530 (N_41530,N_37348,N_39934);
nand U41531 (N_41531,N_32685,N_34226);
xor U41532 (N_41532,N_34012,N_30007);
or U41533 (N_41533,N_35742,N_38167);
or U41534 (N_41534,N_35307,N_36905);
nor U41535 (N_41535,N_31956,N_33654);
nor U41536 (N_41536,N_39352,N_31976);
xnor U41537 (N_41537,N_30726,N_35124);
or U41538 (N_41538,N_30816,N_33995);
or U41539 (N_41539,N_38077,N_36987);
or U41540 (N_41540,N_39454,N_37756);
and U41541 (N_41541,N_33542,N_32960);
nand U41542 (N_41542,N_37333,N_34343);
or U41543 (N_41543,N_33983,N_33097);
xnor U41544 (N_41544,N_37717,N_32326);
or U41545 (N_41545,N_34873,N_33328);
or U41546 (N_41546,N_33105,N_35286);
xnor U41547 (N_41547,N_30463,N_37785);
and U41548 (N_41548,N_32556,N_36314);
nand U41549 (N_41549,N_39487,N_36130);
and U41550 (N_41550,N_30314,N_38965);
and U41551 (N_41551,N_35095,N_35545);
and U41552 (N_41552,N_34831,N_38477);
nand U41553 (N_41553,N_38886,N_39528);
nor U41554 (N_41554,N_32892,N_38680);
nor U41555 (N_41555,N_38484,N_35478);
or U41556 (N_41556,N_30202,N_30683);
xor U41557 (N_41557,N_33411,N_35329);
nor U41558 (N_41558,N_37284,N_32139);
nor U41559 (N_41559,N_39628,N_35314);
nor U41560 (N_41560,N_35749,N_37687);
xnor U41561 (N_41561,N_31856,N_39348);
nand U41562 (N_41562,N_30629,N_36768);
and U41563 (N_41563,N_32697,N_30544);
nor U41564 (N_41564,N_34200,N_34501);
nand U41565 (N_41565,N_35878,N_34069);
nor U41566 (N_41566,N_38920,N_36055);
xnor U41567 (N_41567,N_30573,N_34986);
xnor U41568 (N_41568,N_37729,N_32211);
and U41569 (N_41569,N_30437,N_38229);
nand U41570 (N_41570,N_36074,N_38215);
or U41571 (N_41571,N_32226,N_32729);
xor U41572 (N_41572,N_35350,N_31512);
nand U41573 (N_41573,N_31989,N_35096);
and U41574 (N_41574,N_30172,N_32568);
or U41575 (N_41575,N_34809,N_30994);
or U41576 (N_41576,N_36293,N_38068);
and U41577 (N_41577,N_39577,N_39394);
or U41578 (N_41578,N_34301,N_35294);
xor U41579 (N_41579,N_39384,N_33852);
or U41580 (N_41580,N_31998,N_39894);
or U41581 (N_41581,N_34778,N_37836);
or U41582 (N_41582,N_34688,N_32386);
and U41583 (N_41583,N_35644,N_33393);
xnor U41584 (N_41584,N_34921,N_34613);
nand U41585 (N_41585,N_35888,N_33936);
and U41586 (N_41586,N_30002,N_39306);
xor U41587 (N_41587,N_36412,N_36972);
or U41588 (N_41588,N_37460,N_31775);
nand U41589 (N_41589,N_36966,N_30483);
nand U41590 (N_41590,N_30039,N_32295);
xnor U41591 (N_41591,N_33728,N_33324);
and U41592 (N_41592,N_31902,N_32744);
or U41593 (N_41593,N_38369,N_38388);
and U41594 (N_41594,N_37282,N_30884);
and U41595 (N_41595,N_30000,N_38358);
nand U41596 (N_41596,N_34168,N_39746);
and U41597 (N_41597,N_31840,N_31050);
xnor U41598 (N_41598,N_38750,N_34863);
and U41599 (N_41599,N_38605,N_31259);
and U41600 (N_41600,N_30704,N_33061);
and U41601 (N_41601,N_32971,N_34558);
nor U41602 (N_41602,N_30590,N_35235);
nand U41603 (N_41603,N_32241,N_35244);
xnor U41604 (N_41604,N_31038,N_39554);
xor U41605 (N_41605,N_33197,N_34757);
and U41606 (N_41606,N_33120,N_35939);
or U41607 (N_41607,N_38873,N_37596);
or U41608 (N_41608,N_32938,N_35114);
xor U41609 (N_41609,N_33837,N_39887);
or U41610 (N_41610,N_30163,N_34512);
or U41611 (N_41611,N_33742,N_37577);
or U41612 (N_41612,N_30948,N_35442);
nand U41613 (N_41613,N_34249,N_34212);
and U41614 (N_41614,N_32203,N_32147);
nand U41615 (N_41615,N_38709,N_39113);
nor U41616 (N_41616,N_35051,N_33963);
nand U41617 (N_41617,N_30389,N_34054);
or U41618 (N_41618,N_35081,N_35496);
xor U41619 (N_41619,N_36806,N_30574);
nor U41620 (N_41620,N_35304,N_37386);
xnor U41621 (N_41621,N_33628,N_30827);
or U41622 (N_41622,N_36648,N_36039);
and U41623 (N_41623,N_33996,N_39767);
xnor U41624 (N_41624,N_32400,N_32220);
nor U41625 (N_41625,N_38412,N_38054);
or U41626 (N_41626,N_39410,N_31519);
or U41627 (N_41627,N_35780,N_31027);
nand U41628 (N_41628,N_37363,N_31932);
nor U41629 (N_41629,N_34797,N_38227);
or U41630 (N_41630,N_36327,N_31039);
xnor U41631 (N_41631,N_36804,N_35227);
nand U41632 (N_41632,N_35800,N_37858);
and U41633 (N_41633,N_32951,N_30367);
xor U41634 (N_41634,N_32129,N_30851);
xnor U41635 (N_41635,N_35056,N_31618);
xor U41636 (N_41636,N_37498,N_31722);
xor U41637 (N_41637,N_35331,N_32450);
and U41638 (N_41638,N_31375,N_36586);
nand U41639 (N_41639,N_31423,N_34108);
and U41640 (N_41640,N_34101,N_34616);
nand U41641 (N_41641,N_31133,N_34895);
nand U41642 (N_41642,N_35706,N_38072);
nand U41643 (N_41643,N_30563,N_32154);
or U41644 (N_41644,N_34358,N_38590);
nand U41645 (N_41645,N_32467,N_39941);
nand U41646 (N_41646,N_33169,N_30902);
xnor U41647 (N_41647,N_32887,N_36523);
and U41648 (N_41648,N_32718,N_32228);
or U41649 (N_41649,N_39273,N_30269);
nor U41650 (N_41650,N_30872,N_37549);
nand U41651 (N_41651,N_39900,N_37447);
nand U41652 (N_41652,N_31298,N_30667);
nor U41653 (N_41653,N_30567,N_35073);
and U41654 (N_41654,N_37522,N_39670);
or U41655 (N_41655,N_36089,N_32496);
nor U41656 (N_41656,N_36319,N_38305);
and U41657 (N_41657,N_39529,N_36757);
nand U41658 (N_41658,N_38923,N_32520);
xor U41659 (N_41659,N_38482,N_31082);
nand U41660 (N_41660,N_37293,N_39499);
nor U41661 (N_41661,N_34338,N_37639);
or U41662 (N_41662,N_39064,N_31497);
xnor U41663 (N_41663,N_31200,N_30382);
xor U41664 (N_41664,N_36995,N_36764);
xor U41665 (N_41665,N_35397,N_33505);
and U41666 (N_41666,N_34828,N_36098);
nand U41667 (N_41667,N_36172,N_37146);
nor U41668 (N_41668,N_38148,N_30015);
nor U41669 (N_41669,N_30196,N_30641);
nand U41670 (N_41670,N_37875,N_38398);
and U41671 (N_41671,N_34647,N_36627);
xnor U41672 (N_41672,N_30616,N_34444);
xnor U41673 (N_41673,N_33472,N_32507);
nand U41674 (N_41674,N_30433,N_35724);
nor U41675 (N_41675,N_39119,N_37477);
and U41676 (N_41676,N_38898,N_31070);
nor U41677 (N_41677,N_31006,N_34662);
nor U41678 (N_41678,N_38114,N_33006);
xor U41679 (N_41679,N_39974,N_34415);
nor U41680 (N_41680,N_32182,N_36377);
nand U41681 (N_41681,N_37944,N_37260);
nor U41682 (N_41682,N_38019,N_34880);
xor U41683 (N_41683,N_35429,N_32390);
xor U41684 (N_41684,N_33502,N_35198);
xnor U41685 (N_41685,N_32456,N_30809);
nor U41686 (N_41686,N_33039,N_34525);
or U41687 (N_41687,N_30757,N_38218);
nand U41688 (N_41688,N_34345,N_35111);
nand U41689 (N_41689,N_32559,N_31151);
or U41690 (N_41690,N_38665,N_37842);
and U41691 (N_41691,N_37446,N_32885);
nor U41692 (N_41692,N_34055,N_37769);
nand U41693 (N_41693,N_30831,N_34059);
and U41694 (N_41694,N_38043,N_32513);
or U41695 (N_41695,N_30141,N_31791);
nand U41696 (N_41696,N_36246,N_38854);
nor U41697 (N_41697,N_32453,N_35564);
and U41698 (N_41698,N_35076,N_33905);
nand U41699 (N_41699,N_36002,N_37116);
nand U41700 (N_41700,N_38748,N_35472);
nor U41701 (N_41701,N_37945,N_30280);
or U41702 (N_41702,N_37985,N_35615);
or U41703 (N_41703,N_31122,N_38615);
or U41704 (N_41704,N_37010,N_39330);
nor U41705 (N_41705,N_36188,N_34018);
and U41706 (N_41706,N_39817,N_32577);
xnor U41707 (N_41707,N_32039,N_30322);
xor U41708 (N_41708,N_30331,N_35711);
xnor U41709 (N_41709,N_30714,N_30142);
and U41710 (N_41710,N_31630,N_31927);
and U41711 (N_41711,N_37768,N_39297);
nor U41712 (N_41712,N_36190,N_37746);
xor U41713 (N_41713,N_37570,N_37179);
nor U41714 (N_41714,N_37346,N_35400);
xor U41715 (N_41715,N_32384,N_37164);
and U41716 (N_41716,N_33720,N_36368);
or U41717 (N_41717,N_39737,N_35320);
nor U41718 (N_41718,N_33846,N_34256);
or U41719 (N_41719,N_31409,N_34934);
xnor U41720 (N_41720,N_36046,N_31126);
xor U41721 (N_41721,N_32823,N_34370);
and U41722 (N_41722,N_31241,N_33696);
and U41723 (N_41723,N_34273,N_36531);
and U41724 (N_41724,N_37275,N_36672);
nor U41725 (N_41725,N_34218,N_37161);
nand U41726 (N_41726,N_33404,N_37837);
xor U41727 (N_41727,N_38221,N_31260);
xor U41728 (N_41728,N_38450,N_31213);
nand U41729 (N_41729,N_35822,N_32773);
nand U41730 (N_41730,N_35418,N_30534);
or U41731 (N_41731,N_38010,N_39759);
or U41732 (N_41732,N_31843,N_31577);
nand U41733 (N_41733,N_36173,N_33857);
xor U41734 (N_41734,N_38938,N_39160);
and U41735 (N_41735,N_36669,N_37989);
and U41736 (N_41736,N_30480,N_36877);
and U41737 (N_41737,N_38182,N_34920);
and U41738 (N_41738,N_34785,N_33798);
nand U41739 (N_41739,N_30059,N_37914);
or U41740 (N_41740,N_30169,N_39845);
nor U41741 (N_41741,N_32589,N_37068);
or U41742 (N_41742,N_37177,N_34542);
xor U41743 (N_41743,N_39184,N_34341);
and U41744 (N_41744,N_38826,N_36433);
nor U41745 (N_41745,N_34540,N_35074);
nor U41746 (N_41746,N_39354,N_35393);
nand U41747 (N_41747,N_35975,N_35176);
and U41748 (N_41748,N_35747,N_35323);
nor U41749 (N_41749,N_34896,N_36553);
nor U41750 (N_41750,N_32501,N_36452);
xnor U41751 (N_41751,N_34851,N_34701);
or U41752 (N_41752,N_35292,N_32620);
or U41753 (N_41753,N_35085,N_33757);
or U41754 (N_41754,N_30949,N_38553);
and U41755 (N_41755,N_38455,N_31145);
xor U41756 (N_41756,N_39707,N_30064);
xnor U41757 (N_41757,N_38756,N_37315);
xor U41758 (N_41758,N_34187,N_32633);
or U41759 (N_41759,N_34094,N_34621);
and U41760 (N_41760,N_37759,N_35785);
nand U41761 (N_41761,N_33235,N_35312);
xor U41762 (N_41762,N_32998,N_30090);
xnor U41763 (N_41763,N_30343,N_36735);
nor U41764 (N_41764,N_39475,N_37327);
xor U41765 (N_41765,N_36296,N_32316);
and U41766 (N_41766,N_33621,N_30892);
nor U41767 (N_41767,N_36268,N_37324);
or U41768 (N_41768,N_37757,N_34606);
nor U41769 (N_41769,N_38429,N_34875);
nor U41770 (N_41770,N_32110,N_37292);
or U41771 (N_41771,N_39508,N_31304);
xor U41772 (N_41772,N_38939,N_35385);
or U41773 (N_41773,N_33108,N_30692);
nand U41774 (N_41774,N_34111,N_37524);
nand U41775 (N_41775,N_37801,N_31227);
nand U41776 (N_41776,N_36711,N_39408);
xnor U41777 (N_41777,N_31061,N_30193);
nor U41778 (N_41778,N_33215,N_37600);
nor U41779 (N_41779,N_39802,N_32419);
nor U41780 (N_41780,N_31984,N_39040);
nand U41781 (N_41781,N_38513,N_31556);
or U41782 (N_41782,N_32666,N_32054);
and U41783 (N_41783,N_39814,N_35355);
and U41784 (N_41784,N_32839,N_37006);
nand U41785 (N_41785,N_39588,N_32651);
nor U41786 (N_41786,N_39647,N_37365);
nand U41787 (N_41787,N_31632,N_37921);
and U41788 (N_41788,N_39403,N_31660);
and U41789 (N_41789,N_31970,N_35260);
nor U41790 (N_41790,N_36647,N_38180);
or U41791 (N_41791,N_30794,N_34098);
nand U41792 (N_41792,N_39337,N_33727);
xnor U41793 (N_41793,N_34403,N_39909);
nand U41794 (N_41794,N_30497,N_35850);
nand U41795 (N_41795,N_39699,N_31234);
and U41796 (N_41796,N_32156,N_39694);
nand U41797 (N_41797,N_30250,N_35630);
or U41798 (N_41798,N_39449,N_33918);
nor U41799 (N_41799,N_30441,N_37492);
nand U41800 (N_41800,N_38970,N_39389);
nor U41801 (N_41801,N_33739,N_36010);
or U41802 (N_41802,N_33334,N_34166);
nor U41803 (N_41803,N_36563,N_36994);
xor U41804 (N_41804,N_32198,N_33901);
and U41805 (N_41805,N_34172,N_35945);
nor U41806 (N_41806,N_32037,N_32637);
nor U41807 (N_41807,N_33159,N_38080);
nor U41808 (N_41808,N_30372,N_38490);
nand U41809 (N_41809,N_31209,N_36110);
or U41810 (N_41810,N_30286,N_30263);
and U41811 (N_41811,N_34601,N_38946);
or U41812 (N_41812,N_35827,N_39045);
xor U41813 (N_41813,N_31015,N_33137);
nor U41814 (N_41814,N_32135,N_36079);
xnor U41815 (N_41815,N_35974,N_37279);
nand U41816 (N_41816,N_37691,N_32313);
nand U41817 (N_41817,N_36402,N_34471);
nor U41818 (N_41818,N_30311,N_36955);
nand U41819 (N_41819,N_30889,N_38582);
nand U41820 (N_41820,N_31322,N_33252);
nand U41821 (N_41821,N_34935,N_34894);
or U41822 (N_41822,N_36450,N_33687);
nand U41823 (N_41823,N_30845,N_36572);
nand U41824 (N_41824,N_36562,N_35834);
nand U41825 (N_41825,N_34459,N_31659);
or U41826 (N_41826,N_39756,N_39765);
and U41827 (N_41827,N_35940,N_31224);
and U41828 (N_41828,N_36133,N_37063);
xnor U41829 (N_41829,N_36332,N_35743);
nand U41830 (N_41830,N_30830,N_30321);
and U41831 (N_41831,N_36534,N_32566);
xnor U41832 (N_41832,N_36468,N_37650);
or U41833 (N_41833,N_36953,N_36164);
nand U41834 (N_41834,N_36558,N_36527);
nand U41835 (N_41835,N_38903,N_37136);
or U41836 (N_41836,N_35903,N_31539);
xor U41837 (N_41837,N_37732,N_33083);
nand U41838 (N_41838,N_33659,N_34128);
and U41839 (N_41839,N_38934,N_38065);
xnor U41840 (N_41840,N_36300,N_39078);
xor U41841 (N_41841,N_39689,N_31048);
and U41842 (N_41842,N_39947,N_36070);
nand U41843 (N_41843,N_32221,N_32307);
and U41844 (N_41844,N_32380,N_38788);
nand U41845 (N_41845,N_30796,N_32193);
nor U41846 (N_41846,N_33759,N_30526);
nor U41847 (N_41847,N_31597,N_32917);
nand U41848 (N_41848,N_30598,N_37941);
and U41849 (N_41849,N_31236,N_38594);
and U41850 (N_41850,N_34158,N_38089);
nand U41851 (N_41851,N_38243,N_33991);
xnor U41852 (N_41852,N_36075,N_37294);
nor U41853 (N_41853,N_34373,N_35038);
nand U41854 (N_41854,N_34397,N_34432);
xnor U41855 (N_41855,N_35776,N_35804);
xnor U41856 (N_41856,N_31745,N_38220);
nor U41857 (N_41857,N_38165,N_34449);
xnor U41858 (N_41858,N_35004,N_36744);
xnor U41859 (N_41859,N_36336,N_36555);
nand U41860 (N_41860,N_31333,N_33089);
nor U41861 (N_41861,N_36058,N_36237);
or U41862 (N_41862,N_31088,N_33369);
nor U41863 (N_41863,N_39978,N_35875);
nor U41864 (N_41864,N_38034,N_31225);
and U41865 (N_41865,N_32014,N_39779);
and U41866 (N_41866,N_37167,N_34024);
xor U41867 (N_41867,N_38537,N_34228);
and U41868 (N_41868,N_38629,N_30710);
nand U41869 (N_41869,N_34136,N_36822);
xor U41870 (N_41870,N_34290,N_35525);
nand U41871 (N_41871,N_35127,N_30815);
xor U41872 (N_41872,N_33101,N_34789);
xor U41873 (N_41873,N_33871,N_36112);
or U41874 (N_41874,N_30601,N_32871);
nor U41875 (N_41875,N_33382,N_31948);
nand U41876 (N_41876,N_39562,N_35180);
and U41877 (N_41877,N_34346,N_37087);
or U41878 (N_41878,N_32767,N_30194);
and U41879 (N_41879,N_34717,N_35006);
nand U41880 (N_41880,N_34125,N_39844);
nand U41881 (N_41881,N_32065,N_31058);
nand U41882 (N_41882,N_31469,N_39065);
nand U41883 (N_41883,N_31546,N_32837);
and U41884 (N_41884,N_39530,N_39089);
xor U41885 (N_41885,N_32829,N_34794);
or U41886 (N_41886,N_35431,N_32327);
or U41887 (N_41887,N_36270,N_34500);
and U41888 (N_41888,N_32690,N_35745);
xnor U41889 (N_41889,N_38036,N_38570);
xor U41890 (N_41890,N_30785,N_36618);
nor U41891 (N_41891,N_30126,N_32974);
xor U41892 (N_41892,N_34400,N_35797);
nor U41893 (N_41893,N_38283,N_39094);
nand U41894 (N_41894,N_33142,N_35264);
or U41895 (N_41895,N_35864,N_36996);
xnor U41896 (N_41896,N_36998,N_36308);
nor U41897 (N_41897,N_34989,N_38836);
nor U41898 (N_41898,N_33013,N_36061);
and U41899 (N_41899,N_39553,N_38092);
and U41900 (N_41900,N_33508,N_33181);
or U41901 (N_41901,N_33217,N_30499);
or U41902 (N_41902,N_36717,N_36144);
xnor U41903 (N_41903,N_31393,N_37042);
or U41904 (N_41904,N_32999,N_34071);
and U41905 (N_41905,N_31536,N_36925);
and U41906 (N_41906,N_33889,N_30543);
and U41907 (N_41907,N_30261,N_33634);
and U41908 (N_41908,N_38780,N_36944);
or U41909 (N_41909,N_35934,N_34036);
or U41910 (N_41910,N_32913,N_31465);
nor U41911 (N_41911,N_38702,N_32976);
xor U41912 (N_41912,N_38915,N_33141);
nor U41913 (N_41913,N_32173,N_30888);
nor U41914 (N_41914,N_33248,N_35242);
and U41915 (N_41915,N_33087,N_32922);
nor U41916 (N_41916,N_38700,N_37286);
nor U41917 (N_41917,N_33136,N_35345);
xor U41918 (N_41918,N_31743,N_34793);
or U41919 (N_41919,N_33140,N_30720);
nor U41920 (N_41920,N_38281,N_39316);
and U41921 (N_41921,N_33381,N_32791);
nand U41922 (N_41922,N_33312,N_34840);
nand U41923 (N_41923,N_36622,N_37565);
nor U41924 (N_41924,N_38927,N_37634);
nor U41925 (N_41925,N_34716,N_33970);
and U41926 (N_41926,N_35356,N_36404);
or U41927 (N_41927,N_33121,N_36948);
xnor U41928 (N_41928,N_35468,N_39602);
and U41929 (N_41929,N_31445,N_39371);
and U41930 (N_41930,N_36123,N_34678);
xor U41931 (N_41931,N_39134,N_36066);
and U41932 (N_41932,N_33461,N_31289);
nand U41933 (N_41933,N_34571,N_35928);
or U41934 (N_41934,N_30040,N_35540);
nor U41935 (N_41935,N_37244,N_39506);
nor U41936 (N_41936,N_39608,N_36884);
xor U41937 (N_41937,N_31261,N_30073);
or U41938 (N_41938,N_34149,N_37456);
and U41939 (N_41939,N_34439,N_35893);
or U41940 (N_41940,N_38708,N_37452);
and U41941 (N_41941,N_39597,N_36608);
and U41942 (N_41942,N_39344,N_33053);
or U41943 (N_41943,N_35553,N_39311);
or U41944 (N_41944,N_38776,N_33613);
nor U41945 (N_41945,N_32860,N_34553);
nor U41946 (N_41946,N_37478,N_38195);
nor U41947 (N_41947,N_31987,N_35692);
nor U41948 (N_41948,N_38406,N_39395);
nand U41949 (N_41949,N_35803,N_38119);
nand U41950 (N_41950,N_33412,N_34799);
xnor U41951 (N_41951,N_33616,N_39663);
or U41952 (N_41952,N_38051,N_37469);
nand U41953 (N_41953,N_34008,N_34374);
and U41954 (N_41954,N_32369,N_31141);
and U41955 (N_41955,N_30812,N_35386);
and U41956 (N_41956,N_37673,N_38841);
xor U41957 (N_41957,N_32184,N_31017);
nand U41958 (N_41958,N_32016,N_39822);
nand U41959 (N_41959,N_39843,N_36198);
or U41960 (N_41960,N_34490,N_35701);
nor U41961 (N_41961,N_32225,N_31116);
and U41962 (N_41962,N_37494,N_31143);
or U41963 (N_41963,N_34462,N_32680);
or U41964 (N_41964,N_33610,N_36365);
or U41965 (N_41965,N_36902,N_39341);
xor U41966 (N_41966,N_30950,N_38995);
nand U41967 (N_41967,N_33109,N_31004);
xor U41968 (N_41968,N_31033,N_35597);
nor U41969 (N_41969,N_31441,N_39917);
xor U41970 (N_41970,N_30103,N_39618);
nor U41971 (N_41971,N_36936,N_32965);
xor U41972 (N_41972,N_31809,N_31887);
xnor U41973 (N_41973,N_30702,N_31089);
or U41974 (N_41974,N_33395,N_37947);
nor U41975 (N_41975,N_34299,N_32598);
and U41976 (N_41976,N_34651,N_34208);
or U41977 (N_41977,N_31824,N_37588);
and U41978 (N_41978,N_32768,N_38346);
and U41979 (N_41979,N_30841,N_31785);
or U41980 (N_41980,N_35061,N_38516);
xnor U41981 (N_41981,N_35102,N_39710);
and U41982 (N_41982,N_32291,N_32800);
nand U41983 (N_41983,N_38508,N_30198);
nor U41984 (N_41984,N_31369,N_39404);
and U41985 (N_41985,N_36202,N_34958);
xor U41986 (N_41986,N_31964,N_31848);
xor U41987 (N_41987,N_38950,N_38634);
xor U41988 (N_41988,N_39565,N_31582);
xnor U41989 (N_41989,N_32177,N_31239);
and U41990 (N_41990,N_39946,N_38672);
nand U41991 (N_41991,N_30696,N_38492);
and U41992 (N_41992,N_34084,N_38038);
or U41993 (N_41993,N_34294,N_39202);
or U41994 (N_41994,N_37062,N_39442);
nand U41995 (N_41995,N_31316,N_35960);
nand U41996 (N_41996,N_30793,N_35633);
or U41997 (N_41997,N_35340,N_32151);
nor U41998 (N_41998,N_30545,N_39430);
and U41999 (N_41999,N_38638,N_35952);
and U42000 (N_42000,N_37518,N_33683);
nor U42001 (N_42001,N_35088,N_38630);
and U42002 (N_42002,N_30148,N_31342);
nand U42003 (N_42003,N_31634,N_38607);
nand U42004 (N_42004,N_32334,N_39721);
nand U42005 (N_42005,N_39082,N_32691);
nor U42006 (N_42006,N_35786,N_30391);
xor U42007 (N_42007,N_33725,N_31411);
nor U42008 (N_42008,N_32954,N_35444);
xor U42009 (N_42009,N_31495,N_35333);
xnor U42010 (N_42010,N_39810,N_37531);
and U42011 (N_42011,N_35026,N_33321);
and U42012 (N_42012,N_32783,N_32136);
nor U42013 (N_42013,N_39701,N_39531);
nor U42014 (N_42014,N_31701,N_32140);
and U42015 (N_42015,N_37111,N_34335);
or U42016 (N_42016,N_33776,N_39654);
or U42017 (N_42017,N_33303,N_38251);
nand U42018 (N_42018,N_35563,N_31522);
xor U42019 (N_42019,N_31688,N_35805);
nor U42020 (N_42020,N_36522,N_38091);
and U42021 (N_42021,N_31616,N_31306);
nand U42022 (N_42022,N_38845,N_34391);
and U42023 (N_42023,N_34202,N_31591);
nand U42024 (N_42024,N_32911,N_38882);
nand U42025 (N_42025,N_36451,N_37490);
or U42026 (N_42026,N_34554,N_37191);
and U42027 (N_42027,N_35582,N_31159);
or U42028 (N_42028,N_36016,N_32233);
nand U42029 (N_42029,N_33752,N_39147);
xnor U42030 (N_42030,N_39906,N_34209);
nor U42031 (N_42031,N_32357,N_38835);
or U42032 (N_42032,N_31034,N_36876);
or U42033 (N_42033,N_33134,N_34657);
xor U42034 (N_42034,N_35572,N_35781);
xor U42035 (N_42035,N_36391,N_31876);
nand U42036 (N_42036,N_34021,N_39916);
xor U42037 (N_42037,N_31100,N_31643);
and U42038 (N_42038,N_36991,N_36854);
and U42039 (N_42039,N_31370,N_31277);
and U42040 (N_42040,N_37886,N_36265);
nand U42041 (N_42041,N_38699,N_35769);
nor U42042 (N_42042,N_39397,N_33570);
nor U42043 (N_42043,N_38507,N_34883);
or U42044 (N_42044,N_36924,N_33579);
or U42045 (N_42045,N_37325,N_30036);
or U42046 (N_42046,N_30489,N_36861);
xnor U42047 (N_42047,N_36078,N_34053);
and U42048 (N_42048,N_39828,N_35782);
and U42049 (N_42049,N_36899,N_36342);
and U42050 (N_42050,N_37706,N_32144);
nand U42051 (N_42051,N_39910,N_32929);
or U42052 (N_42052,N_35369,N_30803);
or U42053 (N_42053,N_33366,N_38573);
and U42054 (N_42054,N_33617,N_34596);
nand U42055 (N_42055,N_32979,N_35638);
and U42056 (N_42056,N_33557,N_35043);
or U42057 (N_42057,N_35543,N_34288);
xor U42058 (N_42058,N_33724,N_39329);
xnor U42059 (N_42059,N_32548,N_31460);
nor U42060 (N_42060,N_34664,N_30593);
or U42061 (N_42061,N_37093,N_30292);
nand U42062 (N_42062,N_36040,N_37984);
xnor U42063 (N_42063,N_38963,N_39627);
nor U42064 (N_42064,N_33073,N_34761);
nor U42065 (N_42065,N_31066,N_36453);
and U42066 (N_42066,N_34207,N_31515);
nor U42067 (N_42067,N_37401,N_33536);
and U42068 (N_42068,N_38834,N_34271);
or U42069 (N_42069,N_37817,N_32271);
nor U42070 (N_42070,N_37431,N_36178);
nor U42071 (N_42071,N_36521,N_32890);
nor U42072 (N_42072,N_34642,N_37404);
nor U42073 (N_42073,N_35810,N_33939);
nor U42074 (N_42074,N_31386,N_39896);
nand U42075 (N_42075,N_38729,N_31105);
nand U42076 (N_42076,N_37742,N_34016);
nor U42077 (N_42077,N_34597,N_38744);
xnor U42078 (N_42078,N_30520,N_36551);
nand U42079 (N_42079,N_33572,N_35379);
nor U42080 (N_42080,N_38368,N_33778);
and U42081 (N_42081,N_36777,N_34312);
and U42082 (N_42082,N_39752,N_37877);
or U42083 (N_42083,N_33418,N_37020);
or U42084 (N_42084,N_35003,N_39284);
nor U42085 (N_42085,N_35764,N_32942);
nor U42086 (N_42086,N_31336,N_31721);
or U42087 (N_42087,N_35849,N_38688);
nor U42088 (N_42088,N_34317,N_38348);
nand U42089 (N_42089,N_37266,N_34823);
or U42090 (N_42090,N_36903,N_30087);
nand U42091 (N_42091,N_36263,N_30353);
or U42092 (N_42092,N_34767,N_38158);
and U42093 (N_42093,N_30001,N_33440);
or U42094 (N_42094,N_39262,N_30290);
or U42095 (N_42095,N_31010,N_37648);
or U42096 (N_42096,N_31338,N_33349);
or U42097 (N_42097,N_38659,N_30930);
nand U42098 (N_42098,N_33787,N_39543);
nand U42099 (N_42099,N_37423,N_31908);
and U42100 (N_42100,N_34418,N_37312);
and U42101 (N_42101,N_31960,N_35306);
and U42102 (N_42102,N_36838,N_35705);
or U42103 (N_42103,N_35421,N_33957);
xnor U42104 (N_42104,N_37754,N_39393);
nand U42105 (N_42105,N_39183,N_39362);
and U42106 (N_42106,N_37241,N_37915);
and U42107 (N_42107,N_32494,N_31301);
nor U42108 (N_42108,N_38228,N_37957);
and U42109 (N_42109,N_37466,N_33498);
xnor U42110 (N_42110,N_35092,N_36405);
nor U42111 (N_42111,N_38852,N_39126);
and U42112 (N_42112,N_37054,N_37199);
xnor U42113 (N_42113,N_34163,N_36569);
nor U42114 (N_42114,N_36285,N_36938);
nor U42115 (N_42115,N_31180,N_35215);
or U42116 (N_42116,N_35192,N_33955);
xor U42117 (N_42117,N_38136,N_34871);
nor U42118 (N_42118,N_34992,N_31679);
and U42119 (N_42119,N_39674,N_37969);
or U42120 (N_42120,N_37416,N_35089);
and U42121 (N_42121,N_30097,N_34962);
nor U42122 (N_42122,N_38404,N_39233);
and U42123 (N_42123,N_36707,N_34615);
nor U42124 (N_42124,N_35188,N_35870);
xor U42125 (N_42125,N_32125,N_31567);
and U42126 (N_42126,N_38428,N_36436);
and U42127 (N_42127,N_34295,N_38489);
nor U42128 (N_42128,N_38499,N_30999);
nor U42129 (N_42129,N_36916,N_30846);
nand U42130 (N_42130,N_35741,N_37897);
nand U42131 (N_42131,N_33868,N_39178);
nor U42132 (N_42132,N_32223,N_32247);
nor U42133 (N_42133,N_38501,N_31813);
xnor U42134 (N_42134,N_31559,N_33684);
or U42135 (N_42135,N_30307,N_36274);
nor U42136 (N_42136,N_30395,N_38384);
nand U42137 (N_42137,N_31627,N_32896);
xor U42138 (N_42138,N_38379,N_36739);
nor U42139 (N_42139,N_38217,N_34137);
or U42140 (N_42140,N_31857,N_39586);
xor U42141 (N_42141,N_32076,N_39172);
xnor U42142 (N_42142,N_32217,N_38921);
nand U42143 (N_42143,N_36175,N_31635);
or U42144 (N_42144,N_38875,N_30045);
nor U42145 (N_42145,N_35814,N_32586);
and U42146 (N_42146,N_33346,N_37480);
nor U42147 (N_42147,N_38937,N_37882);
and U42148 (N_42148,N_35953,N_31150);
nand U42149 (N_42149,N_31667,N_39683);
nor U42150 (N_42150,N_39435,N_35021);
nor U42151 (N_42151,N_33785,N_31229);
nor U42152 (N_42152,N_39864,N_31699);
xor U42153 (N_42153,N_30693,N_35795);
or U42154 (N_42154,N_35567,N_36805);
xnor U42155 (N_42155,N_32719,N_39000);
nor U42156 (N_42156,N_36607,N_31207);
or U42157 (N_42157,N_30259,N_35986);
and U42158 (N_42158,N_32641,N_36458);
xnor U42159 (N_42159,N_38650,N_33014);
nand U42160 (N_42160,N_32747,N_33859);
nand U42161 (N_42161,N_32206,N_37725);
xor U42162 (N_42162,N_32188,N_33828);
nor U42163 (N_42163,N_34723,N_39104);
xor U42164 (N_42164,N_33794,N_30592);
nor U42165 (N_42165,N_32788,N_39545);
nor U42166 (N_42166,N_30538,N_33660);
nor U42167 (N_42167,N_30119,N_31831);
nor U42168 (N_42168,N_37686,N_34541);
nand U42169 (N_42169,N_37407,N_38014);
nand U42170 (N_42170,N_35116,N_32031);
nor U42171 (N_42171,N_30711,N_36504);
and U42172 (N_42172,N_34214,N_30804);
xnor U42173 (N_42173,N_31513,N_36983);
xor U42174 (N_42174,N_33090,N_32966);
or U42175 (N_42175,N_35631,N_39682);
xnor U42176 (N_42176,N_38187,N_38473);
xor U42177 (N_42177,N_34965,N_31420);
and U42178 (N_42178,N_32927,N_38676);
xor U42179 (N_42179,N_33383,N_35538);
and U42180 (N_42180,N_37894,N_31842);
xor U42181 (N_42181,N_39358,N_33322);
and U42182 (N_42182,N_36476,N_33203);
or U42183 (N_42183,N_39494,N_33754);
and U42184 (N_42184,N_33951,N_39717);
or U42185 (N_42185,N_37342,N_32743);
nor U42186 (N_42186,N_34477,N_30376);
xor U42187 (N_42187,N_39521,N_37832);
or U42188 (N_42188,N_39913,N_35791);
xnor U42189 (N_42189,N_36824,N_39558);
nor U42190 (N_42190,N_32365,N_36116);
nand U42191 (N_42191,N_38437,N_39481);
or U42192 (N_42192,N_30032,N_31308);
or U42193 (N_42193,N_32745,N_39204);
and U42194 (N_42194,N_34910,N_37660);
or U42195 (N_42195,N_36338,N_38968);
xnor U42196 (N_42196,N_33790,N_38561);
nor U42197 (N_42197,N_32989,N_32874);
or U42198 (N_42198,N_31242,N_35461);
nor U42199 (N_42199,N_30764,N_35539);
or U42200 (N_42200,N_32888,N_31959);
xor U42201 (N_42201,N_30580,N_38772);
nor U42202 (N_42202,N_36785,N_30955);
nand U42203 (N_42203,N_37857,N_38226);
or U42204 (N_42204,N_37461,N_34769);
xnor U42205 (N_42205,N_36547,N_38042);
nand U42206 (N_42206,N_38856,N_37851);
xnor U42207 (N_42207,N_33313,N_31212);
nand U42208 (N_42208,N_39880,N_35913);
nor U42209 (N_42209,N_33166,N_38157);
nor U42210 (N_42210,N_39522,N_38028);
nand U42211 (N_42211,N_33088,N_36429);
nor U42212 (N_42212,N_39424,N_39467);
and U42213 (N_42213,N_33397,N_31124);
nand U42214 (N_42214,N_31216,N_37935);
or U42215 (N_42215,N_30549,N_38267);
nand U42216 (N_42216,N_35498,N_37595);
nor U42217 (N_42217,N_31491,N_31578);
nand U42218 (N_42218,N_33719,N_36481);
or U42219 (N_42219,N_31891,N_33688);
nand U42220 (N_42220,N_31744,N_31543);
nor U42221 (N_42221,N_36799,N_37936);
xnor U42222 (N_42222,N_39445,N_33854);
or U42223 (N_42223,N_30115,N_33241);
xor U42224 (N_42224,N_34821,N_33111);
xor U42225 (N_42225,N_33872,N_35018);
and U42226 (N_42226,N_35748,N_32457);
xor U42227 (N_42227,N_32787,N_32900);
nand U42228 (N_42228,N_39826,N_32434);
or U42229 (N_42229,N_37118,N_39015);
nand U42230 (N_42230,N_32081,N_35375);
and U42231 (N_42231,N_39871,N_38596);
or U42232 (N_42232,N_36102,N_39945);
nand U42233 (N_42233,N_38710,N_30404);
nor U42234 (N_42234,N_33047,N_36980);
xor U42235 (N_42235,N_35767,N_35842);
nand U42236 (N_42236,N_30225,N_30911);
nand U42237 (N_42237,N_33452,N_33619);
and U42238 (N_42238,N_31320,N_35405);
nand U42239 (N_42239,N_39605,N_35272);
nor U42240 (N_42240,N_30916,N_37030);
nand U42241 (N_42241,N_30959,N_31563);
and U42242 (N_42242,N_33956,N_37621);
and U42243 (N_42243,N_39486,N_36542);
nand U42244 (N_42244,N_34710,N_32339);
xnor U42245 (N_42245,N_32451,N_35016);
nand U42246 (N_42246,N_39539,N_32113);
and U42247 (N_42247,N_33406,N_31127);
or U42248 (N_42248,N_34107,N_30434);
nand U42249 (N_42249,N_38673,N_37331);
and U42250 (N_42250,N_36919,N_38331);
xor U42251 (N_42251,N_30009,N_37076);
xnor U42252 (N_42252,N_30284,N_31538);
and U42253 (N_42253,N_31152,N_33437);
xor U42254 (N_42254,N_36536,N_34753);
and U42255 (N_42255,N_37149,N_36258);
nand U42256 (N_42256,N_31468,N_32868);
xnor U42257 (N_42257,N_33494,N_37916);
xor U42258 (N_42258,N_31415,N_32218);
and U42259 (N_42259,N_33764,N_31078);
and U42260 (N_42260,N_37855,N_32563);
and U42261 (N_42261,N_38360,N_31639);
and U42262 (N_42262,N_37352,N_38926);
nor U42263 (N_42263,N_38280,N_39970);
or U42264 (N_42264,N_36709,N_35503);
xnor U42265 (N_42265,N_30212,N_39893);
nor U42266 (N_42266,N_35536,N_30471);
nand U42267 (N_42267,N_30525,N_31433);
nor U42268 (N_42268,N_31511,N_35072);
or U42269 (N_42269,N_39763,N_32381);
xor U42270 (N_42270,N_36791,N_37973);
nor U42271 (N_42271,N_31921,N_30378);
and U42272 (N_42272,N_30490,N_33998);
or U42273 (N_42273,N_36845,N_32524);
xor U42274 (N_42274,N_39956,N_36248);
and U42275 (N_42275,N_30149,N_38558);
or U42276 (N_42276,N_38595,N_37229);
nand U42277 (N_42277,N_33408,N_37137);
and U42278 (N_42278,N_37998,N_32190);
xor U42279 (N_42279,N_37066,N_39169);
xor U42280 (N_42280,N_39925,N_34502);
nand U42281 (N_42281,N_30767,N_36520);
nand U42282 (N_42282,N_37555,N_36417);
xnor U42283 (N_42283,N_37839,N_30448);
nand U42284 (N_42284,N_36474,N_32854);
nand U42285 (N_42285,N_36302,N_39872);
and U42286 (N_42286,N_39569,N_39053);
nand U42287 (N_42287,N_36284,N_36912);
xnor U42288 (N_42288,N_37795,N_36986);
and U42289 (N_42289,N_38807,N_37405);
or U42290 (N_42290,N_38017,N_37236);
and U42291 (N_42291,N_33669,N_32399);
nand U42292 (N_42292,N_30806,N_39447);
nand U42293 (N_42293,N_37356,N_39277);
nor U42294 (N_42294,N_36931,N_31818);
or U42295 (N_42295,N_38442,N_37710);
nor U42296 (N_42296,N_37326,N_39944);
and U42297 (N_42297,N_37097,N_31443);
and U42298 (N_42298,N_30986,N_32686);
nand U42299 (N_42299,N_38572,N_33797);
or U42300 (N_42300,N_32429,N_38310);
nand U42301 (N_42301,N_37433,N_37158);
nand U42302 (N_42302,N_37614,N_39071);
and U42303 (N_42303,N_36609,N_35981);
xnor U42304 (N_42304,N_31807,N_37170);
or U42305 (N_42305,N_32493,N_31542);
nor U42306 (N_42306,N_34796,N_30072);
or U42307 (N_42307,N_37277,N_36192);
or U42308 (N_42308,N_38767,N_39066);
or U42309 (N_42309,N_34454,N_35717);
nor U42310 (N_42310,N_34503,N_35656);
nor U42311 (N_42311,N_30466,N_33340);
xor U42312 (N_42312,N_36697,N_32205);
or U42313 (N_42313,N_30231,N_34838);
nor U42314 (N_42314,N_37766,N_39649);
nor U42315 (N_42315,N_31799,N_36617);
xnor U42316 (N_42316,N_37796,N_32983);
and U42317 (N_42317,N_37378,N_33117);
nor U42318 (N_42318,N_33405,N_36264);
nand U42319 (N_42319,N_34291,N_31193);
nor U42320 (N_42320,N_36559,N_35992);
or U42321 (N_42321,N_31551,N_39620);
xnor U42322 (N_42322,N_39837,N_35757);
nand U42323 (N_42323,N_35201,N_38196);
or U42324 (N_42324,N_39130,N_36232);
and U42325 (N_42325,N_38511,N_33076);
nand U42326 (N_42326,N_38627,N_37893);
xor U42327 (N_42327,N_39472,N_30738);
and U42328 (N_42328,N_32452,N_32180);
nor U42329 (N_42329,N_31504,N_33360);
nand U42330 (N_42330,N_36749,N_35437);
or U42331 (N_42331,N_36625,N_33476);
nand U42332 (N_42332,N_31798,N_35590);
xor U42333 (N_42333,N_32435,N_38323);
nor U42334 (N_42334,N_32342,N_33528);
xor U42335 (N_42335,N_35534,N_30341);
nand U42336 (N_42336,N_38488,N_37306);
xnor U42337 (N_42337,N_31324,N_31310);
nor U42338 (N_42338,N_33234,N_31521);
nand U42339 (N_42339,N_32003,N_34626);
or U42340 (N_42340,N_30415,N_36028);
or U42341 (N_42341,N_37208,N_34353);
or U42342 (N_42342,N_32658,N_32043);
or U42343 (N_42343,N_37636,N_32553);
nand U42344 (N_42344,N_31608,N_33251);
or U42345 (N_42345,N_35107,N_30484);
or U42346 (N_42346,N_37932,N_37878);
or U42347 (N_42347,N_38977,N_32576);
or U42348 (N_42348,N_35618,N_31280);
nor U42349 (N_42349,N_31995,N_38813);
or U42350 (N_42350,N_35891,N_35852);
or U42351 (N_42351,N_34447,N_32038);
nor U42352 (N_42352,N_35052,N_36620);
nor U42353 (N_42353,N_37859,N_38922);
nand U42354 (N_42354,N_33791,N_32712);
and U42355 (N_42355,N_35395,N_30406);
xnor U42356 (N_42356,N_31803,N_39988);
xnor U42357 (N_42357,N_35802,N_34551);
or U42358 (N_42358,N_32010,N_33749);
or U42359 (N_42359,N_32878,N_30519);
or U42360 (N_42360,N_30439,N_36185);
xor U42361 (N_42361,N_34932,N_34205);
nand U42362 (N_42362,N_38248,N_33054);
nor U42363 (N_42363,N_32423,N_30445);
and U42364 (N_42364,N_36316,N_32126);
nand U42365 (N_42365,N_39098,N_35900);
and U42366 (N_42366,N_35819,N_38307);
nand U42367 (N_42367,N_31924,N_38867);
xnor U42368 (N_42368,N_31482,N_38394);
or U42369 (N_42369,N_34899,N_32004);
xor U42370 (N_42370,N_30371,N_36753);
xnor U42371 (N_42371,N_32516,N_32172);
and U42372 (N_42372,N_34327,N_35955);
and U42373 (N_42373,N_39307,N_35378);
or U42374 (N_42374,N_37122,N_35259);
nor U42375 (N_42375,N_37178,N_32265);
nor U42376 (N_42376,N_30604,N_34223);
and U42377 (N_42377,N_35202,N_30236);
xnor U42378 (N_42378,N_38481,N_36000);
nor U42379 (N_42379,N_39211,N_35561);
nand U42380 (N_42380,N_38245,N_32931);
nand U42381 (N_42381,N_34539,N_36540);
xor U42382 (N_42382,N_31893,N_36222);
nand U42383 (N_42383,N_38798,N_36494);
nor U42384 (N_42384,N_39778,N_32405);
xor U42385 (N_42385,N_38340,N_39714);
nor U42386 (N_42386,N_35708,N_37049);
nand U42387 (N_42387,N_37534,N_32569);
xor U42388 (N_42388,N_31240,N_39415);
xor U42389 (N_42389,N_33125,N_31440);
nor U42390 (N_42390,N_31596,N_31862);
nand U42391 (N_42391,N_32292,N_32703);
or U42392 (N_42392,N_35669,N_34567);
nor U42393 (N_42393,N_35512,N_34919);
xnor U42394 (N_42394,N_37159,N_35376);
nand U42395 (N_42395,N_35763,N_38364);
and U42396 (N_42396,N_34282,N_34771);
or U42397 (N_42397,N_34066,N_36801);
nand U42398 (N_42398,N_39072,N_32296);
xor U42399 (N_42399,N_33856,N_30823);
or U42400 (N_42400,N_34037,N_30472);
or U42401 (N_42401,N_36132,N_30548);
and U42402 (N_42402,N_38396,N_38291);
nand U42403 (N_42403,N_31617,N_35490);
or U42404 (N_42404,N_31250,N_32261);
nand U42405 (N_42405,N_34082,N_33295);
nor U42406 (N_42406,N_33212,N_36380);
nand U42407 (N_42407,N_37798,N_34188);
or U42408 (N_42408,N_30786,N_31269);
xor U42409 (N_42409,N_33845,N_36738);
nand U42410 (N_42410,N_33516,N_31044);
nor U42411 (N_42411,N_38877,N_35473);
nor U42412 (N_42412,N_38996,N_34798);
and U42413 (N_42413,N_32469,N_34936);
or U42414 (N_42414,N_36599,N_35951);
nor U42415 (N_42415,N_32269,N_39448);
and U42416 (N_42416,N_39994,N_32996);
xnor U42417 (N_42417,N_31827,N_30901);
xnor U42418 (N_42418,N_30247,N_32275);
nor U42419 (N_42419,N_32952,N_34238);
xnor U42420 (N_42420,N_37115,N_36982);
nor U42421 (N_42421,N_38785,N_37823);
or U42422 (N_42422,N_37696,N_39860);
nand U42423 (N_42423,N_32058,N_37896);
nor U42424 (N_42424,N_30385,N_38953);
nor U42425 (N_42425,N_35866,N_39073);
nor U42426 (N_42426,N_33562,N_33285);
or U42427 (N_42427,N_36094,N_37705);
xnor U42428 (N_42428,N_30482,N_33453);
or U42429 (N_42429,N_33624,N_31201);
or U42430 (N_42430,N_38600,N_36092);
or U42431 (N_42431,N_35643,N_31446);
and U42432 (N_42432,N_32109,N_30257);
nand U42433 (N_42433,N_37474,N_30449);
nor U42434 (N_42434,N_39319,N_37637);
and U42435 (N_42435,N_37369,N_38718);
or U42436 (N_42436,N_30517,N_31975);
nand U42437 (N_42437,N_37138,N_38491);
nand U42438 (N_42438,N_37597,N_36276);
and U42439 (N_42439,N_35519,N_32115);
nand U42440 (N_42440,N_34520,N_35389);
nand U42441 (N_42441,N_33929,N_32500);
nand U42442 (N_42442,N_37664,N_33953);
and U42443 (N_42443,N_33877,N_36511);
nand U42444 (N_42444,N_30938,N_39325);
xor U42445 (N_42445,N_33512,N_30279);
or U42446 (N_42446,N_31428,N_37659);
nor U42447 (N_42447,N_33736,N_30326);
xor U42448 (N_42448,N_34065,N_35937);
nor U42449 (N_42449,N_34382,N_37127);
and U42450 (N_42450,N_39480,N_32335);
nand U42451 (N_42451,N_30020,N_31095);
or U42452 (N_42452,N_36855,N_31081);
or U42453 (N_42453,N_37592,N_35401);
nand U42454 (N_42454,N_39862,N_37871);
nor U42455 (N_42455,N_37283,N_38698);
nand U42456 (N_42456,N_31179,N_39274);
or U42457 (N_42457,N_37758,N_35610);
xnor U42458 (N_42458,N_36289,N_33534);
nor U42459 (N_42459,N_36287,N_31697);
nand U42460 (N_42460,N_30203,N_31014);
xnor U42461 (N_42461,N_36119,N_30478);
nand U42462 (N_42462,N_37472,N_35559);
nor U42463 (N_42463,N_32822,N_37797);
nand U42464 (N_42464,N_30651,N_37124);
nor U42465 (N_42465,N_35083,N_38433);
nor U42466 (N_42466,N_31573,N_30625);
xor U42467 (N_42467,N_38962,N_34103);
nor U42468 (N_42468,N_33820,N_33587);
or U42469 (N_42469,N_30451,N_32945);
nand U42470 (N_42470,N_38824,N_35374);
nor U42471 (N_42471,N_37072,N_33228);
xor U42472 (N_42472,N_36441,N_31505);
nor U42473 (N_42473,N_34585,N_35305);
nand U42474 (N_42474,N_31211,N_30680);
xnor U42475 (N_42475,N_36141,N_37662);
nor U42476 (N_42476,N_38540,N_36398);
xnor U42477 (N_42477,N_36649,N_39164);
nor U42478 (N_42478,N_39429,N_37340);
xnor U42479 (N_42479,N_35328,N_39741);
nand U42480 (N_42480,N_35183,N_36645);
nor U42481 (N_42481,N_38565,N_34652);
or U42482 (N_42482,N_32440,N_36756);
or U42483 (N_42483,N_34434,N_32142);
nor U42484 (N_42484,N_35199,N_39645);
and U42485 (N_42485,N_35154,N_30585);
and U42486 (N_42486,N_38029,N_31830);
and U42487 (N_42487,N_36721,N_36448);
nor U42488 (N_42488,N_31693,N_32920);
or U42489 (N_42489,N_30017,N_32646);
xor U42490 (N_42490,N_30802,N_32477);
nor U42491 (N_42491,N_30456,N_32019);
nor U42492 (N_42492,N_38016,N_37924);
or U42493 (N_42493,N_37139,N_39022);
and U42494 (N_42494,N_35826,N_31729);
nor U42495 (N_42495,N_34623,N_34365);
or U42496 (N_42496,N_38663,N_32657);
and U42497 (N_42497,N_32257,N_34885);
xor U42498 (N_42498,N_37145,N_39293);
nand U42499 (N_42499,N_31529,N_30770);
and U42500 (N_42500,N_37226,N_39593);
xnor U42501 (N_42501,N_35380,N_31309);
and U42502 (N_42502,N_39060,N_31464);
nand U42503 (N_42503,N_39122,N_35521);
nor U42504 (N_42504,N_31579,N_32738);
nor U42505 (N_42505,N_35621,N_32179);
nand U42506 (N_42506,N_33291,N_38234);
and U42507 (N_42507,N_30136,N_33814);
nand U42508 (N_42508,N_37319,N_33261);
xor U42509 (N_42509,N_36715,N_30427);
nand U42510 (N_42510,N_39989,N_39716);
xor U42511 (N_42511,N_37681,N_38452);
nor U42512 (N_42512,N_33347,N_33112);
xnor U42513 (N_42513,N_31708,N_32891);
nor U42514 (N_42514,N_36823,N_33567);
or U42515 (N_42515,N_30412,N_39194);
and U42516 (N_42516,N_35179,N_34847);
nor U42517 (N_42517,N_39985,N_38979);
nand U42518 (N_42518,N_38357,N_36245);
xor U42519 (N_42519,N_37908,N_34583);
xnor U42520 (N_42520,N_30528,N_38139);
nand U42521 (N_42521,N_36573,N_30468);
and U42522 (N_42522,N_35318,N_31047);
and U42523 (N_42523,N_38434,N_36206);
nand U42524 (N_42524,N_34825,N_38668);
and U42525 (N_42525,N_33388,N_33826);
or U42526 (N_42526,N_30522,N_34978);
or U42527 (N_42527,N_32345,N_33801);
nor U42528 (N_42528,N_32222,N_34979);
xnor U42529 (N_42529,N_36407,N_36091);
or U42530 (N_42530,N_39381,N_33042);
and U42531 (N_42531,N_36637,N_39137);
and U42532 (N_42532,N_34730,N_33522);
and U42533 (N_42533,N_38472,N_38980);
nand U42534 (N_42534,N_35162,N_30721);
nand U42535 (N_42535,N_39827,N_36101);
nand U42536 (N_42536,N_39244,N_37868);
and U42537 (N_42537,N_33070,N_33019);
nand U42538 (N_42538,N_33984,N_32312);
nor U42539 (N_42539,N_31756,N_35731);
xor U42540 (N_42540,N_31311,N_37128);
xnor U42541 (N_42541,N_37248,N_37503);
and U42542 (N_42542,N_36798,N_38714);
and U42543 (N_42543,N_35426,N_34808);
or U42544 (N_42544,N_39399,N_39634);
nand U42545 (N_42545,N_38574,N_34221);
nor U42546 (N_42546,N_34270,N_33717);
nor U42547 (N_42547,N_37777,N_39125);
xor U42548 (N_42548,N_34858,N_36740);
nand U42549 (N_42549,N_30332,N_35760);
nor U42550 (N_42550,N_34804,N_37133);
and U42551 (N_42551,N_30414,N_35585);
and U42552 (N_42552,N_32026,N_37901);
and U42553 (N_42553,N_30476,N_32593);
nor U42554 (N_42554,N_38426,N_38847);
nand U42555 (N_42555,N_38757,N_38252);
nor U42556 (N_42556,N_39253,N_33062);
and U42557 (N_42557,N_35601,N_39195);
nand U42558 (N_42558,N_38603,N_32152);
xnor U42559 (N_42559,N_38376,N_32742);
nor U42560 (N_42560,N_35641,N_36800);
or U42561 (N_42561,N_32464,N_39042);
nand U42562 (N_42562,N_32736,N_36773);
nor U42563 (N_42563,N_34117,N_39426);
xor U42564 (N_42564,N_39921,N_37683);
and U42565 (N_42565,N_36445,N_31077);
and U42566 (N_42566,N_32707,N_35524);
nor U42567 (N_42567,N_35471,N_34704);
nand U42568 (N_42568,N_34123,N_39272);
xor U42569 (N_42569,N_32329,N_38580);
nor U42570 (N_42570,N_31836,N_39140);
or U42571 (N_42571,N_37402,N_38055);
xor U42572 (N_42572,N_37670,N_30494);
xnor U42573 (N_42573,N_33107,N_30759);
and U42574 (N_42574,N_30947,N_31437);
xor U42575 (N_42575,N_34177,N_33293);
or U42576 (N_42576,N_32858,N_34429);
and U42577 (N_42577,N_36937,N_39425);
or U42578 (N_42578,N_38942,N_36115);
nand U42579 (N_42579,N_33964,N_33729);
and U42580 (N_42580,N_37151,N_36514);
or U42581 (N_42581,N_33525,N_36444);
nand U42582 (N_42582,N_31878,N_38660);
or U42583 (N_42583,N_32727,N_36307);
nor U42584 (N_42584,N_39687,N_32991);
xnor U42585 (N_42585,N_39757,N_38260);
and U42586 (N_42586,N_34532,N_30690);
or U42587 (N_42587,N_35060,N_39191);
or U42588 (N_42588,N_35175,N_33931);
nor U42589 (N_42589,N_35535,N_35172);
and U42590 (N_42590,N_33740,N_30542);
and U42591 (N_42591,N_37613,N_37256);
nor U42592 (N_42592,N_38179,N_31678);
xor U42593 (N_42593,N_31279,N_30191);
and U42594 (N_42594,N_33943,N_39969);
nor U42595 (N_42595,N_36403,N_30492);
nor U42596 (N_42596,N_32227,N_32106);
or U42597 (N_42597,N_37163,N_35654);
nor U42598 (N_42598,N_39096,N_32098);
xor U42599 (N_42599,N_32659,N_38181);
nand U42600 (N_42600,N_39214,N_35845);
or U42601 (N_42601,N_31290,N_35729);
and U42602 (N_42602,N_35283,N_30065);
or U42603 (N_42603,N_37900,N_37075);
and U42604 (N_42604,N_35070,N_34297);
xnor U42605 (N_42605,N_30555,N_34033);
xor U42606 (N_42606,N_31928,N_35078);
nand U42607 (N_42607,N_32704,N_39762);
nor U42608 (N_42608,N_35354,N_31895);
and U42609 (N_42609,N_32537,N_38859);
xnor U42610 (N_42610,N_33672,N_37039);
and U42611 (N_42611,N_36473,N_31345);
and U42612 (N_42612,N_32730,N_38894);
or U42613 (N_42613,N_36048,N_39563);
and U42614 (N_42614,N_32044,N_30460);
and U42615 (N_42615,N_31347,N_37671);
xor U42616 (N_42616,N_39524,N_34132);
xnor U42617 (N_42617,N_33592,N_39979);
nand U42618 (N_42618,N_36420,N_36426);
xnor U42619 (N_42619,N_35012,N_33435);
xnor U42620 (N_42620,N_30717,N_32705);
and U42621 (N_42621,N_30227,N_30672);
nor U42622 (N_42622,N_36182,N_32848);
or U42623 (N_42623,N_38419,N_32008);
and U42624 (N_42624,N_31348,N_38671);
or U42625 (N_42625,N_36006,N_35594);
and U42626 (N_42626,N_31865,N_31376);
xnor U42627 (N_42627,N_34220,N_35455);
xnor U42628 (N_42628,N_34901,N_37615);
or U42629 (N_42629,N_38602,N_31727);
nand U42630 (N_42630,N_34326,N_37259);
nor U42631 (N_42631,N_39139,N_30565);
or U42632 (N_42632,N_32781,N_36710);
and U42633 (N_42633,N_35904,N_33245);
and U42634 (N_42634,N_33041,N_31707);
nor U42635 (N_42635,N_38048,N_33840);
nor U42636 (N_42636,N_36162,N_30252);
nand U42637 (N_42637,N_39520,N_37861);
or U42638 (N_42638,N_39583,N_38819);
or U42639 (N_42639,N_31113,N_34907);
and U42640 (N_42640,N_39904,N_37632);
xnor U42641 (N_42641,N_38909,N_36512);
xnor U42642 (N_42642,N_32785,N_35371);
nor U42643 (N_42643,N_37262,N_36949);
or U42644 (N_42644,N_39805,N_38535);
or U42645 (N_42645,N_30752,N_38705);
nand U42646 (N_42646,N_32928,N_30424);
and U42647 (N_42647,N_35346,N_37586);
xnor U42648 (N_42648,N_34001,N_30748);
xnor U42649 (N_42649,N_39672,N_32120);
or U42650 (N_42650,N_38762,N_37788);
nor U42651 (N_42651,N_37728,N_35753);
nor U42652 (N_42652,N_38393,N_38496);
and U42653 (N_42653,N_39509,N_37389);
nand U42654 (N_42654,N_30122,N_38333);
nor U42655 (N_42655,N_38695,N_30226);
nor U42656 (N_42656,N_35275,N_36716);
nand U42657 (N_42657,N_35322,N_33708);
and U42658 (N_42658,N_39705,N_35926);
or U42659 (N_42659,N_38041,N_34627);
and U42660 (N_42660,N_31255,N_31192);
nor U42661 (N_42661,N_33935,N_34527);
nand U42662 (N_42662,N_38764,N_35223);
nand U42663 (N_42663,N_33380,N_37153);
or U42664 (N_42664,N_32602,N_33513);
nor U42665 (N_42665,N_30013,N_38960);
nor U42666 (N_42666,N_35293,N_34364);
or U42667 (N_42667,N_35303,N_39972);
nand U42668 (N_42668,N_38335,N_31672);
or U42669 (N_42669,N_33267,N_35348);
nand U42670 (N_42670,N_32561,N_37826);
or U42671 (N_42671,N_34320,N_34862);
xor U42672 (N_42672,N_31035,N_32407);
or U42673 (N_42673,N_32252,N_36137);
xnor U42674 (N_42674,N_35115,N_39255);
nor U42675 (N_42675,N_34711,N_31120);
and U42676 (N_42676,N_37368,N_38413);
or U42677 (N_42677,N_38818,N_38957);
nor U42678 (N_42678,N_31075,N_30513);
nor U42679 (N_42679,N_30896,N_33981);
or U42680 (N_42680,N_38375,N_35425);
or U42681 (N_42681,N_38529,N_32583);
and U42682 (N_42682,N_33486,N_34089);
xor U42683 (N_42683,N_38741,N_33650);
or U42684 (N_42684,N_35977,N_39664);
nand U42685 (N_42685,N_38079,N_31164);
or U42686 (N_42686,N_39057,N_39836);
and U42687 (N_42687,N_35330,N_36060);
nand U42688 (N_42688,N_39646,N_34810);
xor U42689 (N_42689,N_38206,N_37803);
xnor U42690 (N_42690,N_39017,N_36496);
nor U42691 (N_42691,N_33339,N_38329);
or U42692 (N_42692,N_37720,N_39637);
xor U42693 (N_42693,N_30069,N_36214);
nor U42694 (N_42694,N_36732,N_31381);
nand U42695 (N_42695,N_33833,N_33436);
xnor U42696 (N_42696,N_33732,N_34905);
or U42697 (N_42697,N_31363,N_30174);
xor U42698 (N_42698,N_34351,N_33372);
nand U42699 (N_42699,N_33145,N_38414);
nand U42700 (N_42700,N_33663,N_37290);
nor U42701 (N_42701,N_39527,N_38354);
nor U42702 (N_42702,N_30557,N_38742);
nand U42703 (N_42703,N_30011,N_36816);
and U42704 (N_42704,N_32196,N_30034);
nand U42705 (N_42705,N_30964,N_37355);
or U42706 (N_42706,N_34167,N_39062);
or U42707 (N_42707,N_30512,N_36610);
nor U42708 (N_42708,N_35161,N_38541);
or U42709 (N_42709,N_30041,N_33103);
xnor U42710 (N_42710,N_30336,N_39842);
and U42711 (N_42711,N_30895,N_30200);
nor U42712 (N_42712,N_35410,N_36272);
xnor U42713 (N_42713,N_37948,N_39280);
nor U42714 (N_42714,N_33032,N_38967);
and U42715 (N_42715,N_38387,N_34631);
nand U42716 (N_42716,N_31545,N_36868);
nor U42717 (N_42717,N_34656,N_32080);
nand U42718 (N_42718,N_39099,N_36472);
nor U42719 (N_42719,N_35189,N_30366);
nand U42720 (N_42720,N_39367,N_31943);
and U42721 (N_42721,N_36549,N_38099);
xor U42722 (N_42722,N_33319,N_30222);
nor U42723 (N_42723,N_35573,N_33184);
xor U42724 (N_42724,N_34802,N_37698);
and U42725 (N_42725,N_39744,N_35930);
nand U42726 (N_42726,N_37961,N_34165);
nor U42727 (N_42727,N_36689,N_31853);
nor U42728 (N_42728,N_38613,N_30457);
xnor U42729 (N_42729,N_38444,N_30758);
xnor U42730 (N_42730,N_37744,N_36886);
xnor U42731 (N_42731,N_38326,N_38986);
xnor U42732 (N_42732,N_38528,N_37052);
or U42733 (N_42733,N_32936,N_37843);
and U42734 (N_42734,N_39230,N_34079);
and U42735 (N_42735,N_38597,N_30599);
and U42736 (N_42736,N_35122,N_33677);
or U42737 (N_42737,N_34412,N_31894);
nand U42738 (N_42738,N_38611,N_31782);
xor U42739 (N_42739,N_31676,N_37417);
nand U42740 (N_42740,N_36587,N_38198);
or U42741 (N_42741,N_34040,N_36552);
or U42742 (N_42742,N_36694,N_31838);
nand U42743 (N_42743,N_38385,N_36939);
xnor U42744 (N_42744,N_39821,N_38469);
nand U42745 (N_42745,N_35533,N_38745);
and U42746 (N_42746,N_33003,N_36461);
nor U42747 (N_42747,N_34376,N_38902);
and U42748 (N_42748,N_36484,N_33188);
nand U42749 (N_42749,N_37235,N_36708);
xnor U42750 (N_42750,N_34876,N_35138);
nor U42751 (N_42751,N_36321,N_37787);
nor U42752 (N_42752,N_34632,N_37862);
nand U42753 (N_42753,N_31099,N_39954);
and U42754 (N_42754,N_38030,N_31267);
nor U42755 (N_42755,N_35726,N_34423);
and U42756 (N_42756,N_30100,N_36842);
and U42757 (N_42757,N_32274,N_35554);
and U42758 (N_42758,N_38746,N_30578);
nand U42759 (N_42759,N_31398,N_34020);
nand U42760 (N_42760,N_32786,N_37215);
and U42761 (N_42761,N_37580,N_35047);
nand U42762 (N_42762,N_30624,N_33666);
nand U42763 (N_42763,N_31631,N_35308);
nand U42764 (N_42764,N_38846,N_31958);
and U42765 (N_42765,N_30245,N_38154);
nor U42766 (N_42766,N_39685,N_33147);
nor U42767 (N_42767,N_35752,N_37033);
and U42768 (N_42768,N_33880,N_35634);
nand U42769 (N_42769,N_39047,N_39975);
or U42770 (N_42770,N_38203,N_35084);
or U42771 (N_42771,N_30910,N_36516);
nor U42772 (N_42772,N_31645,N_37838);
or U42773 (N_42773,N_35808,N_36946);
nor U42774 (N_42774,N_31692,N_35210);
and U42775 (N_42775,N_30932,N_31029);
or U42776 (N_42776,N_34772,N_37958);
nand U42777 (N_42777,N_38256,N_39929);
nand U42778 (N_42778,N_38948,N_30819);
xor U42779 (N_42779,N_31860,N_36788);
nor U42780 (N_42780,N_38647,N_38224);
xor U42781 (N_42781,N_37525,N_33830);
or U42782 (N_42782,N_30773,N_36093);
xnor U42783 (N_42783,N_30474,N_38145);
nand U42784 (N_42784,N_37242,N_30192);
nand U42785 (N_42785,N_30035,N_35526);
xnor U42786 (N_42786,N_37675,N_38682);
and U42787 (N_42787,N_34561,N_31117);
or U42788 (N_42788,N_34927,N_39303);
nand U42789 (N_42789,N_33167,N_30016);
nand U42790 (N_42790,N_33465,N_31983);
xor U42791 (N_42791,N_36122,N_39240);
or U42792 (N_42792,N_37101,N_32735);
nor U42793 (N_42793,N_38971,N_39264);
nand U42794 (N_42794,N_31343,N_31270);
xor U42795 (N_42795,N_33890,N_39285);
nor U42796 (N_42796,N_39870,N_35458);
nand U42797 (N_42797,N_38308,N_34371);
and U42798 (N_42798,N_34264,N_35890);
or U42799 (N_42799,N_33162,N_39068);
or U42800 (N_42800,N_33365,N_36722);
nand U42801 (N_42801,N_34762,N_31602);
nor U42802 (N_42802,N_33043,N_35728);
nor U42803 (N_42803,N_31844,N_35200);
and U42804 (N_42804,N_35316,N_36052);
and U42805 (N_42805,N_33396,N_34155);
and U42806 (N_42806,N_32687,N_31654);
or U42807 (N_42807,N_39118,N_35404);
nor U42808 (N_42808,N_30077,N_36945);
or U42809 (N_42809,N_32057,N_31904);
or U42810 (N_42810,N_35619,N_38209);
nand U42811 (N_42811,N_34598,N_31028);
and U42812 (N_42812,N_35816,N_37413);
and U42813 (N_42813,N_37620,N_34741);
nand U42814 (N_42814,N_37186,N_32013);
and U42815 (N_42815,N_32259,N_35796);
or U42816 (N_42816,N_35794,N_38244);
nor U42817 (N_42817,N_31475,N_32799);
nand U42818 (N_42818,N_38453,N_33783);
xnor U42819 (N_42819,N_38421,N_36396);
nand U42820 (N_42820,N_34706,N_32528);
and U42821 (N_42821,N_33474,N_33968);
and U42822 (N_42822,N_33207,N_31779);
xor U42823 (N_42823,N_36628,N_37415);
nand U42824 (N_42824,N_35080,N_35637);
or U42825 (N_42825,N_31817,N_33417);
nand U42826 (N_42826,N_31318,N_36810);
or U42827 (N_42827,N_35911,N_33667);
or U42828 (N_42828,N_30243,N_39376);
nor U42829 (N_42829,N_30658,N_39556);
xnor U42830 (N_42830,N_36411,N_38912);
nor U42831 (N_42831,N_37876,N_31910);
xnor U42832 (N_42832,N_39501,N_38622);
xor U42833 (N_42833,N_32761,N_30244);
or U42834 (N_42834,N_32943,N_37344);
nor U42835 (N_42835,N_34679,N_30084);
or U42836 (N_42836,N_32364,N_39185);
nand U42837 (N_42837,N_37004,N_31648);
nor U42838 (N_42838,N_39639,N_39263);
nand U42839 (N_42839,N_31837,N_30768);
or U42840 (N_42840,N_35925,N_30691);
and U42841 (N_42841,N_35844,N_32811);
nor U42842 (N_42842,N_31218,N_30033);
nand U42843 (N_42843,N_38917,N_33195);
nand U42844 (N_42844,N_37099,N_33428);
nor U42845 (N_42845,N_32550,N_33004);
and U42846 (N_42846,N_32883,N_32197);
nand U42847 (N_42847,N_30055,N_38543);
xnor U42848 (N_42848,N_30941,N_30510);
and U42849 (N_42849,N_31933,N_36495);
and U42850 (N_42850,N_35550,N_36125);
nor U42851 (N_42851,N_38306,N_37364);
nor U42852 (N_42852,N_31404,N_37934);
xnor U42853 (N_42853,N_31165,N_37790);
or U42854 (N_42854,N_35617,N_39270);
nor U42855 (N_42855,N_32277,N_31436);
xor U42856 (N_42856,N_36535,N_30893);
xnor U42857 (N_42857,N_37483,N_31735);
or U42858 (N_42858,N_37533,N_39361);
nand U42859 (N_42859,N_32805,N_34044);
or U42860 (N_42860,N_39542,N_31523);
xor U42861 (N_42861,N_36850,N_34971);
nand U42862 (N_42862,N_32243,N_37867);
or U42863 (N_42863,N_30425,N_38908);
or U42864 (N_42864,N_35222,N_38779);
xnor U42865 (N_42865,N_32402,N_39422);
nor U42866 (N_42866,N_32547,N_30426);
and U42867 (N_42867,N_34378,N_32343);
and U42868 (N_42868,N_33933,N_39514);
or U42869 (N_42869,N_33446,N_33988);
nand U42870 (N_42870,N_35148,N_32614);
xnor U42871 (N_42871,N_33563,N_38598);
nand U42872 (N_42872,N_39162,N_36117);
nand U42873 (N_42873,N_37806,N_30807);
nor U42874 (N_42874,N_33220,N_30505);
nand U42875 (N_42875,N_39831,N_38152);
and U42876 (N_42876,N_31890,N_37493);
nand U42877 (N_42877,N_35991,N_30755);
or U42878 (N_42878,N_39176,N_34121);
nor U42879 (N_42879,N_32455,N_34913);
and U42880 (N_42880,N_32439,N_39709);
nor U42881 (N_42881,N_36388,N_38853);
and U42882 (N_42882,N_30763,N_39012);
nand U42883 (N_42883,N_33855,N_34961);
nand U42884 (N_42884,N_38536,N_34237);
or U42885 (N_42885,N_30776,N_38383);
or U42886 (N_42886,N_34234,N_30797);
nor U42887 (N_42887,N_38008,N_36626);
nand U42888 (N_42888,N_38988,N_37513);
and U42889 (N_42889,N_31592,N_37102);
or U42890 (N_42890,N_30107,N_37484);
or U42891 (N_42891,N_36675,N_30516);
xnor U42892 (N_42892,N_31011,N_35602);
and U42893 (N_42893,N_31072,N_31389);
nand U42894 (N_42894,N_31480,N_30355);
nand U42895 (N_42895,N_33509,N_34140);
xnor U42896 (N_42896,N_35407,N_36883);
nor U42897 (N_42897,N_32474,N_33942);
nand U42898 (N_42898,N_30568,N_34293);
nand U42899 (N_42899,N_37999,N_38532);
xnor U42900 (N_42900,N_34061,N_32698);
or U42901 (N_42901,N_30140,N_37181);
xnor U42902 (N_42902,N_37653,N_30800);
or U42903 (N_42903,N_36309,N_37134);
xor U42904 (N_42904,N_35315,N_38539);
or U42905 (N_42905,N_37628,N_36096);
xor U42906 (N_42906,N_32283,N_38330);
nand U42907 (N_42907,N_30109,N_36373);
or U42908 (N_42908,N_38232,N_34725);
nand U42909 (N_42909,N_37874,N_34543);
or U42910 (N_42910,N_32459,N_38468);
xor U42911 (N_42911,N_30524,N_33885);
xnor U42912 (N_42912,N_31674,N_34735);
nand U42913 (N_42913,N_39336,N_34406);
nor U42914 (N_42914,N_35182,N_34728);
and U42915 (N_42915,N_31533,N_36003);
and U42916 (N_42916,N_36491,N_35915);
and U42917 (N_42917,N_32594,N_33618);
or U42918 (N_42918,N_31032,N_38355);
nand U42919 (N_42919,N_33473,N_36566);
and U42920 (N_42920,N_32607,N_33413);
xnor U42921 (N_42921,N_36208,N_36742);
or U42922 (N_42922,N_36150,N_36974);
and U42923 (N_42923,N_31346,N_38110);
xnor U42924 (N_42924,N_31922,N_37499);
or U42925 (N_42925,N_37247,N_37849);
or U42926 (N_42926,N_37722,N_33590);
nand U42927 (N_42927,N_32432,N_31354);
nand U42928 (N_42928,N_38951,N_35108);
and U42929 (N_42929,N_33682,N_39549);
and U42930 (N_42930,N_35427,N_32471);
or U42931 (N_42931,N_31883,N_38789);
nand U42932 (N_42932,N_38443,N_31914);
nand U42933 (N_42933,N_31771,N_36471);
nor U42934 (N_42934,N_32185,N_30784);
or U42935 (N_42935,N_38207,N_35734);
nor U42936 (N_42936,N_37652,N_32395);
and U42937 (N_42937,N_36083,N_38047);
nor U42938 (N_42938,N_32463,N_36465);
and U42939 (N_42939,N_39580,N_30603);
and U42940 (N_42940,N_39728,N_39027);
and U42941 (N_42941,N_34836,N_37963);
nor U42942 (N_42942,N_31967,N_32071);
nand U42943 (N_42943,N_32063,N_31666);
nor U42944 (N_42944,N_35477,N_38947);
xnor U42945 (N_42945,N_32397,N_34867);
xor U42946 (N_42946,N_34591,N_35758);
or U42947 (N_42947,N_37091,N_38755);
xnor U42948 (N_42948,N_30125,N_35877);
or U42949 (N_42949,N_35414,N_39052);
xnor U42950 (N_42950,N_37143,N_30291);
xnor U42951 (N_42951,N_33591,N_31009);
and U42952 (N_42952,N_34038,N_32174);
xor U42953 (N_42953,N_34760,N_39544);
nor U42954 (N_42954,N_31941,N_36590);
nor U42955 (N_42955,N_30615,N_31432);
xnor U42956 (N_42956,N_39818,N_34773);
xor U42957 (N_42957,N_33337,N_35555);
nor U42958 (N_42958,N_34709,N_33829);
and U42959 (N_42959,N_39291,N_34011);
xnor U42960 (N_42960,N_31503,N_33938);
or U42961 (N_42961,N_33588,N_39513);
nor U42962 (N_42962,N_30746,N_37661);
nand U42963 (N_42963,N_38192,N_31188);
and U42964 (N_42964,N_36406,N_39416);
or U42965 (N_42965,N_36830,N_38983);
or U42966 (N_42966,N_33034,N_37799);
or U42967 (N_42967,N_35144,N_30744);
nor U42968 (N_42968,N_36651,N_30705);
and U42969 (N_42969,N_33216,N_30318);
or U42970 (N_42970,N_31670,N_34112);
xnor U42971 (N_42971,N_31424,N_35959);
and U42972 (N_42972,N_38343,N_33808);
and U42973 (N_42973,N_34308,N_30915);
nor U42974 (N_42974,N_34952,N_39785);
nor U42975 (N_42975,N_37424,N_36138);
nand U42976 (N_42976,N_39030,N_38201);
nor U42977 (N_42977,N_38425,N_37511);
xor U42978 (N_42978,N_37154,N_37918);
nand U42979 (N_42979,N_32341,N_33813);
xnor U42980 (N_42980,N_30409,N_39166);
xnor U42981 (N_42981,N_32543,N_31738);
or U42982 (N_42982,N_35265,N_36942);
nor U42983 (N_42983,N_30919,N_39832);
xor U42984 (N_42984,N_38796,N_32012);
or U42985 (N_42985,N_32492,N_30649);
and U42986 (N_42986,N_34674,N_31001);
nor U42987 (N_42987,N_33645,N_30496);
nor U42988 (N_42988,N_39613,N_38646);
and U42989 (N_42989,N_35068,N_34633);
and U42990 (N_42990,N_37193,N_32078);
xor U42991 (N_42991,N_32048,N_31210);
nand U42992 (N_42992,N_33288,N_35022);
xor U42993 (N_42993,N_37379,N_35604);
or U42994 (N_42994,N_32187,N_32926);
xor U42995 (N_42995,N_37443,N_35266);
and U42996 (N_42996,N_33327,N_39816);
and U42997 (N_42997,N_33789,N_35486);
xnor U42998 (N_42998,N_34524,N_30030);
xor U42999 (N_42999,N_37879,N_38493);
nand U43000 (N_43000,N_36815,N_35956);
nor U43001 (N_43001,N_37865,N_33824);
and U43002 (N_43002,N_39334,N_31153);
and U43003 (N_43003,N_39177,N_33273);
xor U43004 (N_43004,N_35463,N_36601);
nand U43005 (N_43005,N_39155,N_31915);
and U43006 (N_43006,N_38037,N_32893);
nand U43007 (N_43007,N_31360,N_35607);
or U43008 (N_43008,N_34720,N_32833);
xor U43009 (N_43009,N_36124,N_39085);
xnor U43010 (N_43010,N_35690,N_36349);
nor U43011 (N_43011,N_30572,N_30535);
and U43012 (N_43012,N_39570,N_39106);
and U43013 (N_43013,N_34589,N_34937);
xnor U43014 (N_43014,N_34368,N_35584);
or U43015 (N_43015,N_35880,N_39951);
nand U43016 (N_43016,N_33978,N_35768);
nand U43017 (N_43017,N_34835,N_38111);
and U43018 (N_43018,N_32835,N_38587);
nand U43019 (N_43019,N_32009,N_36449);
nor U43020 (N_43020,N_37329,N_34608);
nand U43021 (N_43021,N_39990,N_30605);
nor U43022 (N_43022,N_38550,N_38735);
nand U43023 (N_43023,N_34988,N_39400);
xor U43024 (N_43024,N_34130,N_39471);
and U43025 (N_43025,N_39222,N_30123);
or U43026 (N_43026,N_36571,N_31683);
xor U43027 (N_43027,N_30047,N_31849);
nor U43028 (N_43028,N_37608,N_31997);
or U43029 (N_43029,N_34355,N_38101);
nand U43030 (N_43030,N_39151,N_36431);
nand U43031 (N_43031,N_37771,N_39806);
nor U43032 (N_43032,N_36736,N_33927);
nand U43033 (N_43033,N_39671,N_30747);
or U43034 (N_43034,N_35324,N_36611);
nor U43035 (N_43035,N_39390,N_36347);
nand U43036 (N_43036,N_34846,N_39031);
or U43037 (N_43037,N_33001,N_32763);
and U43038 (N_43038,N_37906,N_39850);
nand U43039 (N_43039,N_38635,N_36226);
xor U43040 (N_43040,N_30824,N_35287);
or U43041 (N_43041,N_31418,N_39186);
or U43042 (N_43042,N_38880,N_34035);
nor U43043 (N_43043,N_32700,N_34560);
xnor U43044 (N_43044,N_31372,N_33818);
nor U43045 (N_43045,N_34779,N_33438);
nand U43046 (N_43046,N_30674,N_37884);
xnor U43047 (N_43047,N_31861,N_35063);
or U43048 (N_43048,N_33283,N_36639);
xnor U43049 (N_43049,N_35660,N_32022);
nand U43050 (N_43050,N_37188,N_37165);
nand U43051 (N_43051,N_39847,N_38339);
xnor U43052 (N_43052,N_34518,N_31041);
nor U43053 (N_43053,N_35969,N_37360);
nand U43054 (N_43054,N_30507,N_32034);
nor U43055 (N_43055,N_30131,N_34085);
and U43056 (N_43056,N_36872,N_38827);
or U43057 (N_43057,N_33499,N_30880);
xnor U43058 (N_43058,N_35457,N_30942);
nand U43059 (N_43059,N_34750,N_32308);
xor U43060 (N_43060,N_33568,N_31644);
nor U43061 (N_43061,N_34377,N_39457);
xor U43062 (N_43062,N_31407,N_32766);
or U43063 (N_43063,N_30028,N_30736);
nand U43064 (N_43064,N_38517,N_32609);
xnor U43065 (N_43065,N_30818,N_35848);
nand U43066 (N_43066,N_39305,N_38686);
and U43067 (N_43067,N_39702,N_37508);
xnor U43068 (N_43068,N_33674,N_30043);
nand U43069 (N_43069,N_34770,N_36369);
and U43070 (N_43070,N_32964,N_36505);
xnor U43071 (N_43071,N_33106,N_31993);
or U43072 (N_43072,N_34912,N_35252);
or U43073 (N_43073,N_38814,N_31787);
nor U43074 (N_43074,N_32802,N_32255);
nor U43075 (N_43075,N_31087,N_38454);
nor U43076 (N_43076,N_39793,N_37850);
or U43077 (N_43077,N_32248,N_33457);
xor U43078 (N_43078,N_36915,N_35732);
nand U43079 (N_43079,N_38888,N_31828);
or U43080 (N_43080,N_36103,N_34635);
xnor U43081 (N_43081,N_30282,N_37204);
xor U43082 (N_43082,N_30068,N_38799);
xor U43083 (N_43083,N_30753,N_35311);
xnor U43084 (N_43084,N_36127,N_37200);
nand U43085 (N_43085,N_39451,N_39246);
and U43086 (N_43086,N_32716,N_32957);
nor U43087 (N_43087,N_39676,N_38515);
xnor U43088 (N_43088,N_32538,N_35032);
nor U43089 (N_43089,N_32171,N_30969);
nor U43090 (N_43090,N_33258,N_37473);
nor U43091 (N_43091,N_38112,N_33172);
or U43092 (N_43092,N_33309,N_32502);
or U43093 (N_43093,N_32629,N_32849);
xor U43094 (N_43094,N_32229,N_30156);
nor U43095 (N_43095,N_36355,N_32804);
or U43096 (N_43096,N_36606,N_31942);
nor U43097 (N_43097,N_38524,N_31002);
or U43098 (N_43098,N_37964,N_36667);
or U43099 (N_43099,N_30633,N_39631);
xnor U43100 (N_43100,N_35160,N_32050);
nor U43101 (N_43101,N_34729,N_38495);
nand U43102 (N_43102,N_34581,N_32771);
xnor U43103 (N_43103,N_38210,N_37643);
xor U43104 (N_43104,N_32555,N_32624);
nand U43105 (N_43105,N_38832,N_39511);
nor U43106 (N_43106,N_30178,N_38205);
or U43107 (N_43107,N_32921,N_35537);
nor U43108 (N_43108,N_38563,N_33762);
or U43109 (N_43109,N_32702,N_38296);
nor U43110 (N_43110,N_35398,N_38166);
nor U43111 (N_43111,N_36784,N_37651);
nand U43112 (N_43112,N_38766,N_37059);
nand U43113 (N_43113,N_35449,N_32374);
nand U43114 (N_43114,N_39758,N_32297);
nand U43115 (N_43115,N_35194,N_34941);
and U43116 (N_43116,N_38174,N_37432);
and U43117 (N_43117,N_32112,N_36344);
nand U43118 (N_43118,N_35203,N_36434);
nor U43119 (N_43119,N_32701,N_38200);
and U43120 (N_43120,N_33546,N_30925);
and U43121 (N_43121,N_36807,N_31658);
nor U43122 (N_43122,N_34240,N_30285);
nor U43123 (N_43123,N_32169,N_39891);
nand U43124 (N_43124,N_33600,N_32525);
and U43125 (N_43125,N_30135,N_38720);
xor U43126 (N_43126,N_36510,N_39555);
nand U43127 (N_43127,N_31944,N_39777);
and U43128 (N_43128,N_30301,N_39926);
nand U43129 (N_43129,N_34243,N_37873);
nor U43130 (N_43130,N_31351,N_34482);
nor U43131 (N_43131,N_31852,N_39667);
or U43132 (N_43132,N_30262,N_36673);
or U43133 (N_43133,N_39600,N_38363);
nand U43134 (N_43134,N_30503,N_36486);
nor U43135 (N_43135,N_35887,N_36082);
and U43136 (N_43136,N_32608,N_35993);
and U43137 (N_43137,N_36303,N_30004);
and U43138 (N_43138,N_39764,N_32508);
and U43139 (N_43139,N_34499,N_38415);
xor U43140 (N_43140,N_32317,N_31992);
nor U43141 (N_43141,N_34304,N_32442);
and U43142 (N_43142,N_37912,N_36077);
and U43143 (N_43143,N_36654,N_31768);
xor U43144 (N_43144,N_34051,N_30750);
xnor U43145 (N_43145,N_36128,N_31991);
nand U43146 (N_43146,N_36825,N_31571);
xor U43147 (N_43147,N_32647,N_38820);
and U43148 (N_43148,N_30138,N_33971);
nand U43149 (N_43149,N_37400,N_37467);
and U43150 (N_43150,N_35898,N_37572);
and U43151 (N_43151,N_32910,N_38133);
xnor U43152 (N_43152,N_39610,N_37185);
nor U43153 (N_43153,N_36820,N_30145);
or U43154 (N_43154,N_34686,N_33676);
xor U43155 (N_43155,N_30128,N_38173);
nor U43156 (N_43156,N_30254,N_37552);
or U43157 (N_43157,N_30317,N_31614);
xnor U43158 (N_43158,N_37977,N_32847);
or U43159 (N_43159,N_33506,N_37183);
nor U43160 (N_43160,N_39698,N_34410);
xnor U43161 (N_43161,N_35109,N_37753);
nand U43162 (N_43162,N_34470,N_34839);
xnor U43163 (N_43163,N_39359,N_34296);
xnor U43164 (N_43164,N_33907,N_39008);
xnor U43165 (N_43165,N_38095,N_31753);
nand U43166 (N_43166,N_39617,N_33627);
and U43167 (N_43167,N_31854,N_32925);
xor U43168 (N_43168,N_36292,N_36135);
and U43169 (N_43169,N_30688,N_30742);
nand U43170 (N_43170,N_36047,N_35954);
nor U43171 (N_43171,N_39462,N_38479);
nand U43172 (N_43172,N_36212,N_32214);
nand U43173 (N_43173,N_34515,N_38409);
nand U43174 (N_43174,N_36290,N_32905);
xnor U43175 (N_43175,N_33341,N_33281);
nor U43176 (N_43176,N_33851,N_37786);
nand U43177 (N_43177,N_36360,N_39321);
or U43178 (N_43178,N_37703,N_33651);
xor U43179 (N_43179,N_38670,N_33625);
xnor U43180 (N_43180,N_37021,N_39474);
nor U43181 (N_43181,N_35055,N_32138);
or U43182 (N_43182,N_31496,N_31858);
and U43183 (N_43183,N_37929,N_30181);
or U43184 (N_43184,N_31593,N_33751);
or U43185 (N_43185,N_36568,N_30197);
nand U43186 (N_43186,N_38169,N_31589);
xnor U43187 (N_43187,N_34973,N_39751);
nor U43188 (N_43188,N_35837,N_34388);
nor U43189 (N_43189,N_33127,N_36596);
xor U43190 (N_43190,N_32253,N_36700);
or U43191 (N_43191,N_38445,N_30383);
nor U43192 (N_43192,N_33848,N_32756);
nand U43193 (N_43193,N_32866,N_36733);
xnor U43194 (N_43194,N_35034,N_35262);
or U43195 (N_43195,N_38812,N_30185);
or U43196 (N_43196,N_37895,N_32853);
xor U43197 (N_43197,N_39734,N_37313);
or U43198 (N_43198,N_37575,N_37582);
and U43199 (N_43199,N_30092,N_31023);
and U43200 (N_43200,N_33675,N_33678);
nor U43201 (N_43201,N_30078,N_33711);
and U43202 (N_43202,N_32889,N_32794);
xor U43203 (N_43203,N_37816,N_35066);
or U43204 (N_43204,N_38395,N_31221);
xnor U43205 (N_43205,N_37201,N_33761);
nor U43206 (N_43206,N_36509,N_33064);
and U43207 (N_43207,N_39019,N_33194);
nand U43208 (N_43208,N_34803,N_39973);
xor U43209 (N_43209,N_32610,N_38759);
and U43210 (N_43210,N_31770,N_39498);
nor U43211 (N_43211,N_37276,N_33582);
xnor U43212 (N_43212,N_32877,N_38464);
or U43213 (N_43213,N_38272,N_34191);
nand U43214 (N_43214,N_38732,N_37092);
xor U43215 (N_43215,N_33298,N_37489);
nor U43216 (N_43216,N_38066,N_30464);
and U43217 (N_43217,N_38623,N_31313);
and U43218 (N_43218,N_39436,N_33095);
and U43219 (N_43219,N_36585,N_34670);
and U43220 (N_43220,N_33864,N_36703);
and U43221 (N_43221,N_34475,N_35230);
xnor U43222 (N_43222,N_33470,N_39625);
nand U43223 (N_43223,N_32495,N_38274);
nor U43224 (N_43224,N_33721,N_38083);
nor U43225 (N_43225,N_31615,N_34303);
and U43226 (N_43226,N_36205,N_36603);
xnor U43227 (N_43227,N_36734,N_30653);
or U43228 (N_43228,N_32997,N_33492);
xnor U43229 (N_43229,N_33469,N_31626);
or U43230 (N_43230,N_34473,N_30613);
and U43231 (N_43231,N_36275,N_39866);
xnor U43232 (N_43232,N_33040,N_34763);
nor U43233 (N_43233,N_37938,N_36932);
and U43234 (N_43234,N_36670,N_30779);
nand U43235 (N_43235,N_30051,N_34908);
or U43236 (N_43236,N_37510,N_38049);
or U43237 (N_43237,N_34183,N_39193);
and U43238 (N_43238,N_38721,N_31459);
or U43239 (N_43239,N_37997,N_34630);
nor U43240 (N_43240,N_34122,N_36323);
xnor U43241 (N_43241,N_37105,N_30756);
and U43242 (N_43242,N_31438,N_35023);
or U43243 (N_43243,N_35233,N_34699);
nand U43244 (N_43244,N_32124,N_36519);
and U43245 (N_43245,N_39980,N_38751);
or U43246 (N_43246,N_38304,N_33932);
or U43247 (N_43247,N_30079,N_30787);
nor U43248 (N_43248,N_36361,N_33934);
and U43249 (N_43249,N_36989,N_37045);
or U43250 (N_43250,N_34866,N_37547);
or U43251 (N_43251,N_31650,N_31620);
nand U43252 (N_43252,N_36256,N_38301);
and U43253 (N_43253,N_36797,N_31979);
xor U43254 (N_43254,N_34328,N_33849);
xor U43255 (N_43255,N_34552,N_34881);
and U43256 (N_43256,N_39238,N_31419);
xnor U43257 (N_43257,N_31647,N_31473);
nor U43258 (N_43258,N_32157,N_38566);
or U43259 (N_43259,N_35445,N_39026);
and U43260 (N_43260,N_30074,N_32023);
nor U43261 (N_43261,N_38175,N_39438);
nand U43262 (N_43262,N_38717,N_33500);
nor U43263 (N_43263,N_36333,N_35762);
nor U43264 (N_43264,N_37640,N_37642);
xnor U43265 (N_43265,N_32565,N_38284);
or U43266 (N_43266,N_34138,N_30971);
and U43267 (N_43267,N_39005,N_32372);
nor U43268 (N_43268,N_31952,N_33578);
and U43269 (N_43269,N_35583,N_39409);
or U43270 (N_43270,N_33658,N_37996);
xor U43271 (N_43271,N_34109,N_37150);
xor U43272 (N_43272,N_32677,N_31815);
xnor U43273 (N_43273,N_35775,N_33092);
nand U43274 (N_43274,N_36588,N_37737);
nor U43275 (N_43275,N_37553,N_32678);
and U43276 (N_43276,N_39338,N_39180);
nor U43277 (N_43277,N_31341,N_34398);
or U43278 (N_43278,N_36397,N_31203);
and U43279 (N_43279,N_37328,N_33315);
nor U43280 (N_43280,N_33649,N_39829);
and U43281 (N_43281,N_36745,N_36941);
or U43282 (N_43282,N_30067,N_35450);
nor U43283 (N_43283,N_31206,N_38525);
nor U43284 (N_43284,N_33392,N_30224);
nor U43285 (N_43285,N_35152,N_39173);
xnor U43286 (N_43286,N_33219,N_34599);
nor U43287 (N_43287,N_34045,N_33333);
or U43288 (N_43288,N_32042,N_33028);
nor U43289 (N_43289,N_38074,N_33225);
nor U43290 (N_43290,N_33693,N_36646);
nor U43291 (N_43291,N_37601,N_36059);
nor U43292 (N_43292,N_36897,N_37420);
nor U43293 (N_43293,N_36159,N_38969);
nand U43294 (N_43294,N_30523,N_37827);
xnor U43295 (N_43295,N_38869,N_32406);
nor U43296 (N_43296,N_38743,N_34013);
nand U43297 (N_43297,N_39660,N_31477);
and U43298 (N_43298,N_31877,N_33641);
nor U43299 (N_43299,N_33118,N_32634);
and U43300 (N_43300,N_36501,N_38032);
nand U43301 (N_43301,N_35881,N_38124);
xor U43302 (N_43302,N_37044,N_32020);
xnor U43303 (N_43303,N_38606,N_32582);
xnor U43304 (N_43304,N_37657,N_33685);
or U43305 (N_43305,N_38677,N_32237);
xor U43306 (N_43306,N_33897,N_32239);
nand U43307 (N_43307,N_33535,N_34830);
xnor U43308 (N_43308,N_31461,N_31327);
nand U43309 (N_43309,N_39148,N_36811);
and U43310 (N_43310,N_30155,N_35515);
or U43311 (N_43311,N_39882,N_32695);
or U43312 (N_43312,N_33306,N_37002);
and U43313 (N_43313,N_34672,N_38150);
xnor U43314 (N_43314,N_37221,N_34476);
nand U43315 (N_43315,N_33639,N_35098);
xnor U43316 (N_43316,N_36796,N_31520);
or U43317 (N_43317,N_34563,N_33874);
nand U43318 (N_43318,N_30255,N_36228);
nor U43319 (N_43319,N_33074,N_38438);
xnor U43320 (N_43320,N_38626,N_39216);
nand U43321 (N_43321,N_37519,N_33246);
xor U43322 (N_43322,N_34252,N_38448);
nand U43323 (N_43323,N_31911,N_36918);
nand U43324 (N_43324,N_38899,N_34660);
or U43325 (N_43325,N_33843,N_38052);
nor U43326 (N_43326,N_36663,N_38924);
xor U43327 (N_43327,N_39182,N_38208);
or U43328 (N_43328,N_32869,N_34203);
nor U43329 (N_43329,N_30399,N_35077);
or U43330 (N_43330,N_37506,N_38151);
nor U43331 (N_43331,N_39260,N_38177);
nor U43332 (N_43332,N_36776,N_38792);
nand U43333 (N_43333,N_33538,N_36271);
nor U43334 (N_43334,N_36042,N_33875);
nand U43335 (N_43335,N_36727,N_30993);
nand U43336 (N_43336,N_36887,N_38259);
nand U43337 (N_43337,N_32912,N_39965);
nor U43338 (N_43338,N_33082,N_32346);
and U43339 (N_43339,N_35403,N_30561);
and U43340 (N_43340,N_35151,N_31223);
or U43341 (N_43341,N_37529,N_33426);
nand U43342 (N_43342,N_37375,N_31713);
nor U43343 (N_43343,N_35838,N_35513);
and U43344 (N_43344,N_34362,N_39181);
and U43345 (N_43345,N_37971,N_33514);
nor U43346 (N_43346,N_36729,N_38815);
nand U43347 (N_43347,N_30419,N_31846);
and U43348 (N_43348,N_39903,N_38531);
nor U43349 (N_43349,N_30547,N_35924);
xnor U43350 (N_43350,N_33326,N_32041);
nand U43351 (N_43351,N_35005,N_38257);
or U43352 (N_43352,N_32625,N_35435);
and U43353 (N_43353,N_32946,N_35313);
nor U43354 (N_43354,N_38275,N_37812);
xor U43355 (N_43355,N_34430,N_36857);
and U43356 (N_43356,N_33804,N_32541);
nor U43357 (N_43357,N_38609,N_37335);
or U43358 (N_43358,N_36659,N_33529);
xnor U43359 (N_43359,N_37685,N_33009);
and U43360 (N_43360,N_36737,N_37820);
nor U43361 (N_43361,N_34389,N_38213);
or U43362 (N_43362,N_39729,N_30241);
or U43363 (N_43363,N_32103,N_35299);
nor U43364 (N_43364,N_39258,N_32638);
xnor U43365 (N_43365,N_39335,N_31899);
nand U43366 (N_43366,N_34042,N_34126);
and U43367 (N_43367,N_34576,N_35754);
nand U43368 (N_43368,N_38470,N_32875);
xor U43369 (N_43369,N_31955,N_30272);
and U43370 (N_43370,N_33959,N_30093);
nand U43371 (N_43371,N_35703,N_34555);
and U43372 (N_43372,N_33861,N_31527);
xor U43373 (N_43373,N_30187,N_39332);
or U43374 (N_43374,N_39889,N_33467);
xor U43375 (N_43375,N_31093,N_35359);
nor U43376 (N_43376,N_37465,N_34332);
or U43377 (N_43377,N_31814,N_33527);
or U43378 (N_43378,N_38510,N_39229);
xor U43379 (N_43379,N_38876,N_37176);
xnor U43380 (N_43380,N_32937,N_35897);
nand U43381 (N_43381,N_34925,N_38655);
or U43382 (N_43382,N_30700,N_36234);
nor U43383 (N_43383,N_39879,N_32178);
or U43384 (N_43384,N_30673,N_39037);
or U43385 (N_43385,N_39380,N_32515);
nand U43386 (N_43386,N_39504,N_33916);
and U43387 (N_43387,N_30621,N_34950);
nor U43388 (N_43388,N_37604,N_33468);
and U43389 (N_43389,N_39773,N_31065);
or U43390 (N_43390,N_34655,N_33835);
nand U43391 (N_43391,N_34087,N_38966);
or U43392 (N_43392,N_30114,N_39295);
or U43393 (N_43393,N_32981,N_39326);
nor U43394 (N_43394,N_38874,N_39128);
or U43395 (N_43395,N_37084,N_38825);
or U43396 (N_43396,N_38294,N_36696);
and U43397 (N_43397,N_39510,N_33254);
and U43398 (N_43398,N_36376,N_33370);
nor U43399 (N_43399,N_35145,N_38349);
and U43400 (N_43400,N_32855,N_30863);
xor U43401 (N_43401,N_30877,N_37558);
xnor U43402 (N_43402,N_30428,N_39740);
and U43403 (N_43403,N_30274,N_30162);
and U43404 (N_43404,N_33375,N_33940);
nand U43405 (N_43405,N_35002,N_37339);
or U43406 (N_43406,N_30418,N_35121);
xor U43407 (N_43407,N_39987,N_35291);
xor U43408 (N_43408,N_31499,N_32770);
and U43409 (N_43409,N_31796,N_36940);
and U43410 (N_43410,N_32552,N_31293);
or U43411 (N_43411,N_37232,N_37119);
nor U43412 (N_43412,N_37357,N_38081);
nor U43413 (N_43413,N_34864,N_30334);
and U43414 (N_43414,N_34697,N_37667);
nand U43415 (N_43415,N_33236,N_35603);
or U43416 (N_43416,N_31806,N_32772);
xnor U43417 (N_43417,N_32604,N_39080);
nand U43418 (N_43418,N_35019,N_31463);
nor U43419 (N_43419,N_34994,N_30175);
nand U43420 (N_43420,N_35746,N_31422);
nand U43421 (N_43421,N_38000,N_36043);
and U43422 (N_43422,N_32224,N_32282);
nor U43423 (N_43423,N_32527,N_34091);
or U43424 (N_43424,N_39414,N_32644);
xnor U43425 (N_43425,N_32201,N_36469);
and U43426 (N_43426,N_37267,N_35876);
and U43427 (N_43427,N_37050,N_36957);
nand U43428 (N_43428,N_34339,N_34637);
xor U43429 (N_43429,N_35737,N_32523);
nor U43430 (N_43430,N_31068,N_31307);
xor U43431 (N_43431,N_37144,N_39226);
and U43432 (N_43432,N_33263,N_39516);
or U43433 (N_43433,N_38505,N_33265);
and U43434 (N_43434,N_36754,N_33462);
nand U43435 (N_43435,N_35337,N_36802);
and U43436 (N_43436,N_38722,N_38954);
xnor U43437 (N_43437,N_31248,N_34170);
xor U43438 (N_43438,N_37476,N_30467);
nor U43439 (N_43439,N_37550,N_31430);
nand U43440 (N_43440,N_36487,N_39933);
or U43441 (N_43441,N_34685,N_32841);
and U43442 (N_43442,N_32378,N_36655);
nor U43443 (N_43443,N_31314,N_38276);
or U43444 (N_43444,N_36142,N_31638);
and U43445 (N_43445,N_33653,N_33781);
nand U43446 (N_43446,N_36241,N_38808);
xor U43447 (N_43447,N_39518,N_35963);
and U43448 (N_43448,N_36831,N_39049);
xnor U43449 (N_43449,N_33243,N_35707);
xnor U43450 (N_43450,N_34306,N_35039);
nor U43451 (N_43451,N_33882,N_35229);
and U43452 (N_43452,N_34698,N_39418);
xnor U43453 (N_43453,N_33979,N_39603);
nand U43454 (N_43454,N_31182,N_39812);
or U43455 (N_43455,N_30260,N_31170);
xor U43456 (N_43456,N_31962,N_30914);
or U43457 (N_43457,N_33496,N_39632);
xnor U43458 (N_43458,N_35451,N_32351);
nand U43459 (N_43459,N_38973,N_33661);
nand U43460 (N_43460,N_33700,N_37343);
or U43461 (N_43461,N_32652,N_36973);
and U43462 (N_43462,N_37899,N_32189);
nor U43463 (N_43463,N_31940,N_37960);
nor U43464 (N_43464,N_37032,N_32813);
xnor U43465 (N_43465,N_33297,N_32183);
or U43466 (N_43466,N_35919,N_39855);
nand U43467 (N_43467,N_36747,N_36860);
xnor U43468 (N_43468,N_36879,N_34765);
and U43469 (N_43469,N_38374,N_38134);
nand U43470 (N_43470,N_36225,N_36935);
nor U43471 (N_43471,N_31337,N_38011);
and U43472 (N_43472,N_38351,N_37853);
nor U43473 (N_43473,N_39800,N_35491);
nor U43474 (N_43474,N_30223,N_37982);
and U43475 (N_43475,N_39825,N_34250);
nand U43476 (N_43476,N_39745,N_32068);
or U43477 (N_43477,N_31025,N_36174);
nor U43478 (N_43478,N_31321,N_38868);
xor U43479 (N_43479,N_30453,N_30083);
and U43480 (N_43480,N_35297,N_37627);
nor U43481 (N_43481,N_33608,N_39797);
and U43482 (N_43482,N_39967,N_38436);
xor U43483 (N_43483,N_33183,N_34347);
or U43484 (N_43484,N_34887,N_33772);
or U43485 (N_43485,N_37169,N_32281);
nand U43486 (N_43486,N_33410,N_37187);
and U43487 (N_43487,N_39742,N_35361);
or U43488 (N_43488,N_38989,N_36140);
nand U43489 (N_43489,N_38704,N_31303);
and U43490 (N_43490,N_38991,N_32234);
or U43491 (N_43491,N_39526,N_34521);
nor U43492 (N_43492,N_32468,N_32655);
nand U43493 (N_43493,N_32170,N_38155);
or U43494 (N_43494,N_39841,N_36213);
or U43495 (N_43495,N_33583,N_30324);
and U43496 (N_43496,N_39452,N_35284);
nand U43497 (N_43497,N_34673,N_36383);
and U43498 (N_43498,N_33296,N_30328);
xnor U43499 (N_43499,N_31186,N_30870);
nand U43500 (N_43500,N_35360,N_36993);
nor U43501 (N_43501,N_34265,N_33620);
nand U43502 (N_43502,N_34544,N_31805);
and U43503 (N_43503,N_37678,N_37345);
nand U43504 (N_43504,N_35062,N_39413);
xnor U43505 (N_43505,N_33454,N_31447);
xor U43506 (N_43506,N_37749,N_31414);
and U43507 (N_43507,N_30722,N_30268);
and U43508 (N_43508,N_31774,N_30602);
nor U43509 (N_43509,N_35289,N_37940);
xnor U43510 (N_43510,N_31394,N_30042);
nand U43511 (N_43511,N_36435,N_30133);
nand U43512 (N_43512,N_39243,N_39688);
or U43513 (N_43513,N_35168,N_38003);
nor U43514 (N_43514,N_39616,N_37655);
and U43515 (N_43515,N_35339,N_31051);
nor U43516 (N_43516,N_35087,N_37422);
xor U43517 (N_43517,N_36532,N_32090);
xnor U43518 (N_43518,N_31112,N_37515);
nand U43519 (N_43519,N_38474,N_31584);
xnor U43520 (N_43520,N_36767,N_35696);
xor U43521 (N_43521,N_30446,N_39953);
nand U43522 (N_43522,N_37258,N_36896);
xor U43523 (N_43523,N_36165,N_34587);
nor U43524 (N_43524,N_37954,N_31686);
and U43525 (N_43525,N_38317,N_30650);
or U43526 (N_43526,N_33906,N_36069);
xor U43527 (N_43527,N_30234,N_34775);
and U43528 (N_43528,N_34083,N_35301);
xor U43529 (N_43529,N_35270,N_32780);
nor U43530 (N_43530,N_31173,N_33960);
and U43531 (N_43531,N_39248,N_30423);
or U43532 (N_43532,N_31892,N_34298);
or U43533 (N_43533,N_31795,N_31283);
nor U43534 (N_43534,N_35310,N_31400);
or U43535 (N_43535,N_34734,N_39188);
xnor U43536 (N_43536,N_30640,N_30644);
or U43537 (N_43537,N_39930,N_36297);
nand U43538 (N_43538,N_34726,N_32383);
nor U43539 (N_43539,N_35196,N_34759);
xor U43540 (N_43540,N_38976,N_30891);
nor U43541 (N_43541,N_34970,N_31726);
nor U43542 (N_43542,N_33504,N_36843);
or U43543 (N_43543,N_38057,N_37041);
nor U43544 (N_43544,N_38571,N_30923);
nor U43545 (N_43545,N_30094,N_33821);
nor U43546 (N_43546,N_37261,N_31091);
or U43547 (N_43547,N_30749,N_39963);
and U43548 (N_43548,N_39704,N_34467);
and U43549 (N_43549,N_34902,N_39942);
and U43550 (N_43550,N_35546,N_39453);
nand U43551 (N_43551,N_35142,N_34027);
nor U43552 (N_43552,N_31402,N_33495);
xor U43553 (N_43553,N_33599,N_34026);
nor U43554 (N_43554,N_30405,N_33652);
nand U43555 (N_43555,N_38405,N_31682);
or U43556 (N_43556,N_30146,N_30556);
nand U43557 (N_43557,N_32127,N_36766);
nor U43558 (N_43558,N_37219,N_30216);
xnor U43559 (N_43559,N_32562,N_32880);
and U43560 (N_43560,N_31929,N_33523);
nand U43561 (N_43561,N_34924,N_34751);
or U43562 (N_43562,N_31183,N_38478);
and U43563 (N_43563,N_34600,N_32077);
and U43564 (N_43564,N_35474,N_31243);
and U43565 (N_43565,N_35962,N_35317);
and U43566 (N_43566,N_30010,N_32564);
nand U43567 (N_43567,N_36146,N_30739);
nor U43568 (N_43568,N_38191,N_38930);
nand U43569 (N_43569,N_33488,N_33350);
and U43570 (N_43570,N_34731,N_39464);
nand U43571 (N_43571,N_38523,N_32532);
nand U43572 (N_43572,N_30150,N_38928);
and U43573 (N_43573,N_37548,N_39852);
and U43574 (N_43574,N_32141,N_39834);
nand U43575 (N_43575,N_31758,N_38461);
nor U43576 (N_43576,N_37285,N_34106);
nand U43577 (N_43577,N_33993,N_32522);
nand U43578 (N_43578,N_34104,N_37863);
or U43579 (N_43579,N_31762,N_32626);
xor U43580 (N_43580,N_34419,N_33131);
nor U43581 (N_43581,N_37202,N_34509);
xor U43582 (N_43582,N_30564,N_31453);
and U43583 (N_43583,N_32803,N_33282);
nor U43584 (N_43584,N_31835,N_31604);
nor U43585 (N_43585,N_35792,N_32683);
xor U43586 (N_43586,N_31457,N_33299);
and U43587 (N_43587,N_30049,N_38512);
nand U43588 (N_43588,N_38342,N_36315);
xnor U43589 (N_43589,N_38022,N_35646);
or U43590 (N_43590,N_30558,N_39469);
nand U43591 (N_43591,N_38560,N_35773);
nand U43592 (N_43592,N_35917,N_39606);
xnor U43593 (N_43593,N_30571,N_35973);
nor U43594 (N_43594,N_33510,N_30369);
nand U43595 (N_43595,N_32465,N_36280);
xor U43596 (N_43596,N_39897,N_34383);
or U43597 (N_43597,N_33515,N_32733);
nand U43598 (N_43598,N_31257,N_32498);
and U43599 (N_43599,N_32670,N_34786);
xor U43600 (N_43600,N_38652,N_38262);
and U43601 (N_43601,N_34914,N_32694);
and U43602 (N_43602,N_35430,N_30108);
and U43603 (N_43603,N_38775,N_39477);
nand U43604 (N_43604,N_35605,N_31655);
and U43605 (N_43605,N_33973,N_32287);
nor U43606 (N_43606,N_36922,N_30973);
nand U43607 (N_43607,N_31387,N_37635);
nor U43608 (N_43608,N_32737,N_35882);
xnor U43609 (N_43609,N_36217,N_31252);
and U43610 (N_43610,N_33763,N_39407);
nand U43611 (N_43611,N_34897,N_38538);
and U43612 (N_43612,N_35675,N_37692);
and U43613 (N_43613,N_35100,N_34629);
nor U43614 (N_43614,N_32280,N_36525);
xnor U43615 (N_43615,N_36371,N_35101);
and U43616 (N_43616,N_39112,N_38643);
nand U43617 (N_43617,N_31816,N_32675);
nand U43618 (N_43618,N_31541,N_38115);
nor U43619 (N_43619,N_30153,N_31391);
nor U43620 (N_43620,N_34745,N_33815);
nor U43621 (N_43621,N_38907,N_30775);
xor U43622 (N_43622,N_32289,N_34976);
xnor U43623 (N_43623,N_31096,N_33553);
nand U43624 (N_43624,N_34689,N_35929);
xor U43625 (N_43625,N_38399,N_32175);
nand U43626 (N_43626,N_37454,N_36216);
or U43627 (N_43627,N_31501,N_32108);
xor U43628 (N_43628,N_34192,N_33354);
xor U43629 (N_43629,N_31057,N_39962);
nand U43630 (N_43630,N_33819,N_32137);
nor U43631 (N_43631,N_37338,N_38690);
xor U43632 (N_43632,N_35899,N_32134);
or U43633 (N_43633,N_37939,N_30554);
or U43634 (N_43634,N_30934,N_30860);
and U43635 (N_43635,N_33543,N_36934);
and U43636 (N_43636,N_31184,N_36557);
or U43637 (N_43637,N_32304,N_30315);
and U43638 (N_43638,N_36136,N_34088);
xnor U43639 (N_43639,N_30868,N_36702);
xnor U43640 (N_43640,N_31052,N_30278);
nand U43641 (N_43641,N_36640,N_33175);
xor U43642 (N_43642,N_39503,N_36892);
xnor U43643 (N_43643,N_38591,N_30686);
xor U43644 (N_43644,N_32393,N_37933);
xor U43645 (N_43645,N_38246,N_31936);
nor U43646 (N_43646,N_34236,N_35146);
xor U43647 (N_43647,N_36184,N_38851);
or U43648 (N_43648,N_34609,N_31489);
nor U43649 (N_43649,N_33018,N_34514);
or U43650 (N_43650,N_32482,N_30989);
or U43651 (N_43651,N_30306,N_33079);
or U43652 (N_43652,N_38219,N_31565);
nor U43653 (N_43653,N_35013,N_34483);
or U43654 (N_43654,N_36171,N_35118);
or U43655 (N_43655,N_39940,N_32472);
xor U43656 (N_43656,N_34691,N_38278);
nand U43657 (N_43657,N_32774,N_34644);
and U43658 (N_43658,N_38778,N_38408);
xor U43659 (N_43659,N_36157,N_33836);
nor U43660 (N_43660,N_30283,N_31094);
nand U43661 (N_43661,N_32302,N_37428);
nand U43662 (N_43662,N_38447,N_37035);
or U43663 (N_43663,N_37449,N_35655);
xor U43664 (N_43664,N_34738,N_36200);
or U43665 (N_43665,N_30540,N_36240);
nand U43666 (N_43666,N_33860,N_37112);
nand U43667 (N_43667,N_32186,N_39584);
nor U43668 (N_43668,N_39747,N_33867);
xor U43669 (N_43669,N_32606,N_37830);
nor U43670 (N_43670,N_35030,N_39695);
nor U43671 (N_43671,N_32812,N_34215);
nor U43672 (N_43672,N_36076,N_31090);
xnor U43673 (N_43673,N_37905,N_31710);
nand U43674 (N_43674,N_33030,N_33071);
xnor U43675 (N_43675,N_38864,N_33780);
and U43676 (N_43676,N_30485,N_30654);
xnor U43677 (N_43677,N_32398,N_30052);
nand U43678 (N_43678,N_39931,N_37704);
and U43679 (N_43679,N_36978,N_36600);
xnor U43680 (N_43680,N_31208,N_30760);
nor U43681 (N_43681,N_39692,N_39912);
or U43682 (N_43682,N_34774,N_33985);
nand U43683 (N_43683,N_30727,N_32782);
and U43684 (N_43684,N_39163,N_35436);
or U43685 (N_43685,N_39650,N_39133);
nor U43686 (N_43686,N_39784,N_36457);
nand U43687 (N_43687,N_37736,N_34898);
nor U43688 (N_43688,N_32021,N_34663);
nand U43689 (N_43689,N_35957,N_32200);
nor U43690 (N_43690,N_36746,N_32972);
nand U43691 (N_43691,N_33888,N_34113);
or U43692 (N_43692,N_32519,N_39347);
or U43693 (N_43693,N_32684,N_37231);
and U43694 (N_43694,N_32445,N_36930);
nor U43695 (N_43695,N_31296,N_34923);
xor U43696 (N_43696,N_33478,N_37666);
or U43697 (N_43697,N_37270,N_34029);
and U43698 (N_43698,N_35394,N_39536);
xnor U43699 (N_43699,N_37184,N_35966);
and U43700 (N_43700,N_31413,N_37104);
nand U43701 (N_43701,N_30875,N_35976);
and U43702 (N_43702,N_32161,N_31685);
xor U43703 (N_43703,N_33239,N_37274);
nor U43704 (N_43704,N_37903,N_33002);
xor U43705 (N_43705,N_30795,N_30101);
or U43706 (N_43706,N_32740,N_31517);
nand U43707 (N_43707,N_33847,N_34356);
xnor U43708 (N_43708,N_30907,N_37468);
or U43709 (N_43709,N_39789,N_31410);
xnor U43710 (N_43710,N_33459,N_30754);
or U43711 (N_43711,N_33316,N_31552);
or U43712 (N_43712,N_39288,N_37055);
or U43713 (N_43713,N_30906,N_31776);
or U43714 (N_43714,N_36508,N_33703);
nand U43715 (N_43715,N_36129,N_35274);
or U43716 (N_43716,N_37699,N_30327);
or U43717 (N_43717,N_37907,N_33150);
and U43718 (N_43718,N_33697,N_31129);
and U43719 (N_43719,N_36660,N_36908);
or U43720 (N_43720,N_30685,N_35137);
or U43721 (N_43721,N_35885,N_30995);
and U43722 (N_43722,N_31481,N_39856);
and U43723 (N_43723,N_38266,N_32204);
nand U43724 (N_43724,N_31266,N_38015);
nand U43725 (N_43725,N_35855,N_37408);
xor U43726 (N_43726,N_37647,N_35821);
or U43727 (N_43727,N_35216,N_36885);
xnor U43728 (N_43728,N_35907,N_30876);
xnor U43729 (N_43729,N_34931,N_32404);
and U43730 (N_43730,N_34433,N_34421);
nand U43731 (N_43731,N_34344,N_37609);
nand U43732 (N_43732,N_32840,N_36545);
or U43733 (N_43733,N_36480,N_31750);
and U43734 (N_43734,N_31733,N_38753);
and U43735 (N_43735,N_33912,N_36518);
xor U43736 (N_43736,N_33980,N_38657);
and U43737 (N_43737,N_35011,N_34791);
or U43738 (N_43738,N_31611,N_35334);
or U43739 (N_43739,N_35720,N_32933);
or U43740 (N_43740,N_35635,N_30670);
nand U43741 (N_43741,N_37303,N_39056);
nor U43742 (N_43742,N_31661,N_34700);
xor U43743 (N_43743,N_31581,N_31390);
nand U43744 (N_43744,N_37719,N_31610);
nor U43745 (N_43745,N_35548,N_34175);
nand U43746 (N_43746,N_30462,N_30983);
nor U43747 (N_43747,N_36345,N_34302);
and U43748 (N_43748,N_37438,N_35522);
nand U43749 (N_43749,N_32886,N_35288);
xnor U43750 (N_43750,N_35596,N_32403);
or U43751 (N_43751,N_35575,N_32619);
nor U43752 (N_43752,N_35125,N_33262);
nand U43753 (N_43753,N_34517,N_37507);
nor U43754 (N_43754,N_30865,N_32441);
and U43755 (N_43755,N_39441,N_32994);
xor U43756 (N_43756,N_36493,N_37316);
and U43757 (N_43757,N_39790,N_35662);
nand U43758 (N_43758,N_38601,N_30111);
and U43759 (N_43759,N_33485,N_37829);
xor U43760 (N_43760,N_38288,N_30712);
nor U43761 (N_43761,N_34904,N_36084);
nor U43762 (N_43762,N_31003,N_30664);
and U43763 (N_43763,N_32752,N_38073);
and U43764 (N_43764,N_37676,N_34258);
nand U43765 (N_43765,N_31695,N_36026);
or U43766 (N_43766,N_35801,N_32732);
or U43767 (N_43767,N_38253,N_35041);
or U43768 (N_43768,N_35155,N_38046);
or U43769 (N_43769,N_39115,N_32895);
or U43770 (N_43770,N_33899,N_32382);
or U43771 (N_43771,N_37701,N_35505);
xnor U43772 (N_43772,N_32850,N_35684);
and U43773 (N_43773,N_34506,N_38144);
nand U43774 (N_43774,N_34959,N_33335);
nor U43775 (N_43775,N_39873,N_39899);
xor U43776 (N_43776,N_35476,N_36045);
nor U43777 (N_43777,N_38131,N_33419);
and U43778 (N_43778,N_39309,N_34039);
or U43779 (N_43779,N_39788,N_38060);
nor U43780 (N_43780,N_34743,N_30118);
nor U43781 (N_43781,N_30931,N_30677);
and U43782 (N_43782,N_34715,N_39546);
nor U43783 (N_43783,N_37318,N_35787);
and U43784 (N_43784,N_33972,N_31526);
nor U43785 (N_43785,N_38380,N_31601);
xor U43786 (N_43786,N_38736,N_36163);
xnor U43787 (N_43787,N_31406,N_31245);
and U43788 (N_43788,N_34092,N_39103);
nand U43789 (N_43789,N_36664,N_30029);
xnor U43790 (N_43790,N_34987,N_30105);
xnor U43791 (N_43791,N_31985,N_36515);
or U43792 (N_43792,N_37920,N_38632);
nand U43793 (N_43793,N_33884,N_34777);
and U43794 (N_43794,N_33331,N_39411);
nand U43795 (N_43795,N_34408,N_39018);
and U43796 (N_43796,N_30300,N_31789);
or U43797 (N_43797,N_35415,N_30304);
and U43798 (N_43798,N_32461,N_33385);
nand U43799 (N_43799,N_35036,N_33865);
nand U43800 (N_43800,N_33133,N_39314);
or U43801 (N_43801,N_34604,N_31797);
nand U43802 (N_43802,N_31479,N_30287);
xnor U43803 (N_43803,N_35851,N_39228);
nand U43804 (N_43804,N_34318,N_38367);
xnor U43805 (N_43805,N_31146,N_36455);
and U43806 (N_43806,N_32679,N_35399);
xnor U43807 (N_43807,N_32585,N_34173);
or U43808 (N_43808,N_32199,N_30668);
xnor U43809 (N_43809,N_35517,N_36636);
xor U43810 (N_43810,N_30741,N_36772);
or U43811 (N_43811,N_36774,N_35723);
nand U43812 (N_43812,N_35462,N_38231);
and U43813 (N_43813,N_39712,N_31725);
or U43814 (N_43814,N_31197,N_36007);
nor U43815 (N_43815,N_30551,N_38315);
nor U43816 (N_43816,N_38122,N_38108);
nor U43817 (N_43817,N_34171,N_37992);
and U43818 (N_43818,N_30502,N_31570);
nor U43819 (N_43819,N_30514,N_34963);
nand U43820 (N_43820,N_38401,N_36705);
nor U43821 (N_43821,N_35606,N_37083);
nor U43822 (N_43822,N_30303,N_37190);
nand U43823 (N_43823,N_35883,N_33947);
nand U43824 (N_43824,N_37970,N_31652);
and U43825 (N_43825,N_34996,N_35665);
or U43826 (N_43826,N_38547,N_36350);
nor U43827 (N_43827,N_31019,N_33475);
nand U43828 (N_43828,N_33161,N_38059);
and U43829 (N_43829,N_37822,N_36105);
xor U43830 (N_43830,N_38581,N_37074);
nor U43831 (N_43831,N_33173,N_30218);
or U43832 (N_43832,N_30498,N_31397);
nor U43833 (N_43833,N_36928,N_38509);
and U43834 (N_43834,N_32236,N_30061);
or U43835 (N_43835,N_37995,N_35994);
xor U43836 (N_43836,N_37735,N_37028);
nand U43837 (N_43837,N_36676,N_30396);
or U43838 (N_43838,N_37125,N_32475);
nor U43839 (N_43839,N_37672,N_30990);
or U43840 (N_43840,N_35530,N_31996);
nand U43841 (N_43841,N_33271,N_34566);
nand U43842 (N_43842,N_32760,N_33806);
or U43843 (N_43843,N_37130,N_36464);
nand U43844 (N_43844,N_32073,N_36230);
nand U43845 (N_43845,N_37429,N_33400);
nand U43846 (N_43846,N_39201,N_35967);
nor U43847 (N_43847,N_37731,N_32894);
or U43848 (N_43848,N_37385,N_37718);
nand U43849 (N_43849,N_30275,N_31792);
or U43850 (N_43850,N_38149,N_39986);
xor U43851 (N_43851,N_31690,N_33611);
nor U43852 (N_43852,N_33735,N_33597);
nand U43853 (N_43853,N_31886,N_36834);
nor U43854 (N_43854,N_35676,N_38548);
xnor U43855 (N_43855,N_33442,N_39835);
nand U43856 (N_43856,N_34849,N_39484);
nor U43857 (N_43857,N_39117,N_33733);
nand U43858 (N_43858,N_37752,N_36317);
nand U43859 (N_43859,N_32980,N_30642);
or U43860 (N_43860,N_39343,N_34888);
nor U43861 (N_43861,N_39323,N_31326);
nand U43862 (N_43862,N_36395,N_37709);
nor U43863 (N_43863,N_39888,N_33532);
xnor U43864 (N_43864,N_35777,N_34219);
nor U43865 (N_43865,N_39276,N_35901);
and U43866 (N_43866,N_38001,N_35470);
xor U43867 (N_43867,N_39420,N_38914);
nand U43868 (N_43868,N_36428,N_36086);
nor U43869 (N_43869,N_35129,N_33384);
and U43870 (N_43870,N_32590,N_35995);
nor U43871 (N_43871,N_38870,N_31897);
and U43872 (N_43872,N_30847,N_32668);
and U43873 (N_43873,N_38656,N_39315);
or U43874 (N_43874,N_39995,N_30864);
xor U43875 (N_43875,N_37180,N_35514);
xnor U43876 (N_43876,N_36415,N_38763);
or U43877 (N_43877,N_39312,N_30182);
and U43878 (N_43878,N_38126,N_39385);
xor U43879 (N_43879,N_33668,N_37132);
nor U43880 (N_43880,N_36180,N_37374);
nand U43881 (N_43881,N_30132,N_39858);
nand U43882 (N_43882,N_31272,N_36726);
nand U43883 (N_43883,N_31558,N_36685);
nor U43884 (N_43884,N_32446,N_30506);
nand U43885 (N_43885,N_38804,N_34077);
xnor U43886 (N_43886,N_34067,N_37828);
and U43887 (N_43887,N_31494,N_32986);
nand U43888 (N_43888,N_30394,N_38407);
xnor U43889 (N_43889,N_39087,N_32089);
nor U43890 (N_43890,N_38910,N_31741);
xor U43891 (N_43891,N_31677,N_36529);
or U43892 (N_43892,N_34349,N_30008);
and U43893 (N_43893,N_37334,N_37943);
and U43894 (N_43894,N_37694,N_39035);
and U43895 (N_43895,N_33544,N_39386);
or U43896 (N_43896,N_37230,N_38773);
nor U43897 (N_43897,N_38285,N_36462);
nor U43898 (N_43898,N_37486,N_31334);
and U43899 (N_43899,N_35674,N_36143);
nor U43900 (N_43900,N_35931,N_33738);
nand U43901 (N_43901,N_35971,N_35416);
nor U43902 (N_43902,N_35481,N_32085);
nor U43903 (N_43903,N_36967,N_32148);
nor U43904 (N_43904,N_35075,N_36589);
nor U43905 (N_43905,N_37612,N_37194);
xnor U43906 (N_43906,N_33367,N_39808);
or U43907 (N_43907,N_31488,N_32628);
nor U43908 (N_43908,N_32958,N_38797);
and U43909 (N_43909,N_31867,N_33786);
or U43910 (N_43910,N_36950,N_33226);
nor U43911 (N_43911,N_31148,N_34041);
nand U43912 (N_43912,N_39281,N_39750);
and U43913 (N_43913,N_38197,N_32903);
xor U43914 (N_43914,N_39534,N_34868);
nand U43915 (N_43915,N_35912,N_31147);
xor U43916 (N_43916,N_37778,N_34582);
or U43917 (N_43917,N_37539,N_38069);
and U43918 (N_43918,N_30026,N_32627);
nand U43919 (N_43919,N_33802,N_37502);
and U43920 (N_43920,N_33914,N_30349);
xor U43921 (N_43921,N_31226,N_32909);
xor U43922 (N_43922,N_39622,N_31486);
and U43923 (N_43923,N_35620,N_36550);
nor U43924 (N_43924,N_34523,N_31158);
xor U43925 (N_43925,N_37026,N_39907);
nor U43926 (N_43926,N_33464,N_33361);
nor U43927 (N_43927,N_34440,N_35278);
or U43928 (N_43928,N_32396,N_37096);
nor U43929 (N_43929,N_31760,N_33990);
nor U43930 (N_43930,N_39596,N_36201);
or U43931 (N_43931,N_36114,N_39142);
or U43932 (N_43932,N_36539,N_39014);
and U43933 (N_43933,N_37665,N_37238);
or U43934 (N_43934,N_33656,N_35053);
or U43935 (N_43935,N_35213,N_39299);
xor U43936 (N_43936,N_39927,N_33704);
nand U43937 (N_43937,N_38651,N_32599);
nor U43938 (N_43938,N_36134,N_36463);
xnor U43939 (N_43939,N_37521,N_34260);
and U43940 (N_43940,N_34675,N_37069);
or U43941 (N_43941,N_33329,N_36856);
xnor U43942 (N_43942,N_34142,N_38313);
nand U43943 (N_43943,N_34605,N_39465);
nand U43944 (N_43944,N_37937,N_33351);
nand U43945 (N_43945,N_34845,N_30238);
xnor U43946 (N_43946,N_35434,N_39582);
xor U43947 (N_43947,N_38860,N_36236);
nand U43948 (N_43948,N_31747,N_30825);
nor U43949 (N_43949,N_36871,N_34493);
or U43950 (N_43950,N_37745,N_37265);
and U43951 (N_43951,N_37761,N_37606);
nand U43952 (N_43952,N_39039,N_39110);
nor U43953 (N_43953,N_33809,N_38327);
and U43954 (N_43954,N_34859,N_39009);
nand U43955 (N_43955,N_39598,N_35156);
or U43956 (N_43956,N_30164,N_31451);
nand U43957 (N_43957,N_36312,N_35806);
nand U43958 (N_43958,N_35873,N_32904);
and U43959 (N_43959,N_32430,N_37781);
or U43960 (N_43960,N_33614,N_30832);
xnor U43961 (N_43961,N_33471,N_39377);
nor U43962 (N_43962,N_31085,N_39540);
nor U43963 (N_43963,N_30086,N_38109);
and U43964 (N_43964,N_34833,N_39289);
xor U43965 (N_43965,N_34917,N_38347);
or U43966 (N_43966,N_31319,N_33705);
or U43967 (N_43967,N_32428,N_31384);
or U43968 (N_43968,N_31547,N_35693);
and U43969 (N_43969,N_32301,N_37573);
and U43970 (N_43970,N_32285,N_35321);
or U43971 (N_43971,N_31137,N_33548);
or U43972 (N_43972,N_32715,N_31668);
nor U43973 (N_43973,N_32842,N_35065);
and U43974 (N_43974,N_31244,N_30533);
nand U43975 (N_43975,N_33858,N_39105);
and U43976 (N_43976,N_30890,N_36678);
nor U43977 (N_43977,N_35069,N_36859);
and U43978 (N_43978,N_38731,N_33842);
nand U43979 (N_43979,N_35440,N_39783);
nand U43980 (N_43980,N_33626,N_35908);
nor U43981 (N_43981,N_38639,N_37910);
nand U43982 (N_43982,N_38837,N_35614);
xor U43983 (N_43983,N_37095,N_37211);
nor U43984 (N_43984,N_35424,N_33158);
xnor U43985 (N_43985,N_31024,N_39074);
nand U43986 (N_43986,N_32424,N_36623);
xor U43987 (N_43987,N_36517,N_37497);
nor U43988 (N_43988,N_33278,N_33163);
nor U43989 (N_43989,N_38678,N_34877);
nor U43990 (N_43990,N_38564,N_37268);
or U43991 (N_43991,N_38527,N_31156);
nand U43992 (N_43992,N_38096,N_39505);
and U43993 (N_43993,N_35892,N_34242);
nor U43994 (N_43994,N_33305,N_31431);
nand U43995 (N_43995,N_35256,N_39443);
or U43996 (N_43996,N_30617,N_31637);
nand U43997 (N_43997,N_35702,N_34985);
nand U43998 (N_43998,N_35428,N_39559);
xnor U43999 (N_43999,N_33766,N_31561);
or U44000 (N_44000,N_37994,N_30853);
nand U44001 (N_44001,N_36803,N_39573);
nand U44002 (N_44002,N_35813,N_36022);
or U44003 (N_44003,N_37668,N_39431);
xnor U44004 (N_44004,N_38641,N_32431);
and U44005 (N_44005,N_30465,N_35238);
and U44006 (N_44006,N_39809,N_38730);
and U44007 (N_44007,N_36862,N_37310);
and U44008 (N_44008,N_33416,N_30926);
and U44009 (N_44009,N_32049,N_31172);
nor U44010 (N_44010,N_34360,N_32852);
and U44011 (N_44011,N_31572,N_38683);
and U44012 (N_44012,N_35456,N_33747);
nor U44013 (N_44013,N_32000,N_30221);
or U44014 (N_44014,N_30242,N_39021);
nor U44015 (N_44015,N_37189,N_36027);
and U44016 (N_44016,N_38990,N_32433);
and U44017 (N_44017,N_38987,N_35049);
and U44018 (N_44018,N_35347,N_32426);
xor U44019 (N_44019,N_33128,N_36056);
xor U44020 (N_44020,N_35506,N_39733);
nor U44021 (N_44021,N_32753,N_35058);
and U44022 (N_44022,N_31864,N_32665);
and U44023 (N_44023,N_37421,N_39658);
and U44024 (N_44024,N_30308,N_36063);
or U44025 (N_44025,N_30904,N_32862);
nand U44026 (N_44026,N_39824,N_31826);
and U44027 (N_44027,N_30529,N_37783);
xor U44028 (N_44028,N_33950,N_32961);
or U44029 (N_44029,N_32414,N_39643);
nand U44030 (N_44030,N_33352,N_34712);
or U44031 (N_44031,N_30204,N_36870);
nor U44032 (N_44032,N_32242,N_39437);
nand U44033 (N_44033,N_37106,N_33520);
or U44034 (N_44034,N_32600,N_37574);
nor U44035 (N_44035,N_34435,N_33604);
or U44036 (N_44036,N_35231,N_31171);
or U44037 (N_44037,N_32645,N_32333);
or U44038 (N_44038,N_39936,N_30373);
or U44039 (N_44039,N_36990,N_38471);
or U44040 (N_44040,N_34284,N_39532);
xnor U44041 (N_44041,N_35370,N_33330);
or U44042 (N_44042,N_36218,N_36029);
nand U44043 (N_44043,N_31934,N_35772);
nor U44044 (N_44044,N_34538,N_34324);
xnor U44045 (N_44045,N_32708,N_39928);
xnor U44046 (N_44046,N_36878,N_33831);
xnor U44047 (N_44047,N_33304,N_33773);
nand U44048 (N_44048,N_39924,N_35446);
xnor U44049 (N_44049,N_32347,N_35086);
or U44050 (N_44050,N_32017,N_39024);
nor U44051 (N_44051,N_33146,N_37775);
nor U44052 (N_44052,N_32086,N_31138);
and U44053 (N_44053,N_31628,N_35028);
xor U44054 (N_44054,N_39579,N_39317);
nor U44055 (N_44055,N_32092,N_31231);
xor U44056 (N_44056,N_37094,N_30814);
nand U44057 (N_44057,N_32597,N_33021);
nand U44058 (N_44058,N_30586,N_30117);
xor U44059 (N_44059,N_39591,N_35557);
or U44060 (N_44060,N_34229,N_30715);
nor U44061 (N_44061,N_31470,N_34386);
or U44062 (N_44062,N_36579,N_37656);
or U44063 (N_44063,N_35131,N_32447);
or U44064 (N_44064,N_36479,N_34841);
nor U44065 (N_44065,N_30656,N_37155);
nor U44066 (N_44066,N_30411,N_32549);
nand U44067 (N_44067,N_31759,N_39059);
xor U44068 (N_44068,N_36324,N_37669);
and U44069 (N_44069,N_38674,N_36985);
and U44070 (N_44070,N_37141,N_38084);
or U44071 (N_44071,N_32166,N_35858);
or U44072 (N_44072,N_33223,N_38176);
and U44073 (N_44073,N_36187,N_35686);
and U44074 (N_44074,N_34003,N_36120);
or U44075 (N_44075,N_39723,N_31977);
and U44076 (N_44076,N_30027,N_35722);
or U44077 (N_44077,N_35600,N_33904);
and U44078 (N_44078,N_32882,N_39232);
xnor U44079 (N_44079,N_32011,N_37968);
and U44080 (N_44080,N_37952,N_34949);
nand U44081 (N_44081,N_31367,N_35422);
nand U44082 (N_44082,N_35874,N_39766);
and U44083 (N_44083,N_37824,N_33896);
xnor U44084 (N_44084,N_39167,N_36421);
or U44085 (N_44085,N_33726,N_38625);
nand U44086 (N_44086,N_30885,N_34276);
or U44087 (N_44087,N_39996,N_39594);
xnor U44088 (N_44088,N_39547,N_34146);
xnor U44089 (N_44089,N_36692,N_31054);
nor U44090 (N_44090,N_32764,N_37485);
xnor U44091 (N_44091,N_39419,N_30215);
nand U44092 (N_44092,N_30984,N_38791);
nor U44093 (N_44093,N_37866,N_35326);
and U44094 (N_44094,N_31366,N_35171);
nor U44095 (N_44095,N_39849,N_38431);
nand U44096 (N_44096,N_32276,N_35113);
nand U44097 (N_44097,N_34300,N_37917);
nand U44098 (N_44098,N_34549,N_30531);
and U44099 (N_44099,N_31653,N_32284);
xor U44100 (N_44100,N_39865,N_34331);
or U44101 (N_44101,N_30980,N_39863);
and U44102 (N_44102,N_39869,N_38026);
and U44103 (N_44103,N_37381,N_38318);
or U44104 (N_44104,N_36408,N_33427);
or U44105 (N_44105,N_38589,N_34405);
and U44106 (N_44106,N_30438,N_39001);
nor U44107 (N_44107,N_39342,N_33153);
nor U44108 (N_44108,N_36751,N_33081);
or U44109 (N_44109,N_32001,N_34073);
xor U44110 (N_44110,N_31588,N_36852);
xnor U44111 (N_44111,N_31125,N_33015);
nor U44112 (N_44112,N_38480,N_34752);
or U44113 (N_44113,N_31870,N_31829);
and U44114 (N_44114,N_37210,N_35487);
nand U44115 (N_44115,N_31408,N_34161);
nor U44116 (N_44116,N_35465,N_35671);
xnor U44117 (N_44117,N_31168,N_32349);
or U44118 (N_44118,N_37131,N_38809);
xnor U44119 (N_44119,N_31484,N_30562);
and U44120 (N_44120,N_34869,N_38403);
and U44121 (N_44121,N_33098,N_34316);
and U44122 (N_44122,N_32790,N_36422);
xnor U44123 (N_44123,N_35494,N_37425);
xor U44124 (N_44124,N_33744,N_31238);
nand U44125 (N_44125,N_34194,N_31925);
nand U44126 (N_44126,N_36095,N_37663);
xor U44127 (N_44127,N_39279,N_32323);
nand U44128 (N_44128,N_34052,N_31205);
and U44129 (N_44129,N_30323,N_34394);
nor U44130 (N_44130,N_38050,N_37967);
nand U44131 (N_44131,N_33743,N_35946);
and U44132 (N_44132,N_33123,N_33037);
and U44133 (N_44133,N_39496,N_39604);
nor U44134 (N_44134,N_38916,N_39353);
nor U44135 (N_44135,N_36723,N_36546);
nor U44136 (N_44136,N_38297,N_37987);
or U44137 (N_44137,N_37714,N_38268);
nor U44138 (N_44138,N_38893,N_35783);
nor U44139 (N_44139,N_33524,N_31472);
xnor U44140 (N_44140,N_35443,N_39680);
xnor U44141 (N_44141,N_32759,N_34015);
and U44142 (N_44142,N_38255,N_32377);
or U44143 (N_44143,N_30944,N_34186);
xnor U44144 (N_44144,N_35097,N_38009);
or U44145 (N_44145,N_39379,N_38941);
xnor U44146 (N_44146,N_32621,N_34030);
and U44147 (N_44147,N_35134,N_30357);
nor U44148 (N_44148,N_38416,N_30293);
nand U44149 (N_44149,N_36147,N_37459);
nand U44150 (N_44150,N_34755,N_31793);
and U44151 (N_44151,N_32028,N_35143);
xnor U44152 (N_44152,N_34653,N_35150);
nor U44153 (N_44153,N_30184,N_31564);
or U44154 (N_44154,N_33373,N_31036);
nand U44155 (N_44155,N_30977,N_33189);
and U44156 (N_44156,N_31454,N_39459);
nand U44157 (N_44157,N_31772,N_33602);
or U44158 (N_44158,N_30553,N_35932);
nand U44159 (N_44159,N_38293,N_35250);
and U44160 (N_44160,N_31049,N_39950);
nand U44161 (N_44161,N_30666,N_35978);
or U44162 (N_44162,N_38692,N_38270);
nand U44163 (N_44163,N_36661,N_34068);
and U44164 (N_44164,N_31557,N_32158);
xor U44165 (N_44165,N_34145,N_35718);
or U44166 (N_44166,N_31114,N_39218);
or U44167 (N_44167,N_35588,N_36254);
xnor U44168 (N_44168,N_30848,N_37846);
and U44169 (N_44169,N_31624,N_36704);
xnor U44170 (N_44170,N_33974,N_30894);
nor U44171 (N_44171,N_32476,N_30927);
nand U44172 (N_44172,N_31219,N_39884);
nand U44173 (N_44173,N_32006,N_36846);
and U44174 (N_44174,N_33517,N_34944);
nand U44175 (N_44175,N_32367,N_34363);
xnor U44176 (N_44176,N_37109,N_37684);
nor U44177 (N_44177,N_31516,N_31299);
or U44178 (N_44178,N_39287,N_37168);
nand U44179 (N_44179,N_30258,N_32260);
nand U44180 (N_44180,N_37317,N_32290);
and U44181 (N_44181,N_37089,N_30151);
and U44182 (N_44182,N_33387,N_33827);
or U44183 (N_44183,N_36911,N_35547);
xor U44184 (N_44184,N_36888,N_38316);
nor U44185 (N_44185,N_37554,N_31777);
or U44186 (N_44186,N_37009,N_36243);
xor U44187 (N_44187,N_38392,N_35824);
xor U44188 (N_44188,N_34893,N_39655);
xor U44189 (N_44189,N_38935,N_39396);
and U44190 (N_44190,N_30852,N_32479);
xor U44191 (N_44191,N_36438,N_32978);
nand U44192 (N_44192,N_38424,N_31673);
nor U44193 (N_44193,N_34577,N_36267);
nor U44194 (N_44194,N_35336,N_35562);
or U44195 (N_44195,N_30912,N_33048);
nand U44196 (N_44196,N_31037,N_32328);
nand U44197 (N_44197,N_34120,N_34529);
and U44198 (N_44198,N_39838,N_38555);
nand U44199 (N_44199,N_37114,N_31973);
nor U44200 (N_44200,N_30160,N_34882);
nand U44201 (N_44201,N_33368,N_39662);
or U44202 (N_44202,N_34144,N_39328);
nand U44203 (N_44203,N_35987,N_37214);
nor U44204 (N_44204,N_34099,N_35357);
nand U44205 (N_44205,N_30495,N_38760);
and U44206 (N_44206,N_33655,N_33926);
nand U44207 (N_44207,N_33466,N_38309);
xnor U44208 (N_44208,N_38696,N_32923);
and U44209 (N_44209,N_33206,N_37207);
xor U44210 (N_44210,N_34696,N_32101);
nand U44211 (N_44211,N_38420,N_30147);
nor U44212 (N_44212,N_38740,N_38269);
or U44213 (N_44213,N_38631,N_35578);
and U44214 (N_44214,N_38033,N_35647);
nand U44215 (N_44215,N_37296,N_31898);
nand U44216 (N_44216,N_37450,N_33240);
xor U44217 (N_44217,N_31101,N_35649);
xor U44218 (N_44218,N_36775,N_32962);
nor U44219 (N_44219,N_34227,N_31903);
nand U44220 (N_44220,N_37646,N_33987);
nand U44221 (N_44221,N_38955,N_30219);
nor U44222 (N_44222,N_31356,N_33482);
xor U44223 (N_44223,N_31166,N_36841);
or U44224 (N_44224,N_35206,N_36390);
nor U44225 (N_44225,N_39225,N_35691);
nor U44226 (N_44226,N_33192,N_37336);
xnor U44227 (N_44227,N_34946,N_38086);
nor U44228 (N_44228,N_39659,N_37726);
nor U44229 (N_44229,N_30340,N_32689);
and U44230 (N_44230,N_38321,N_39159);
or U44231 (N_44231,N_31000,N_33758);
nand U44232 (N_44232,N_39991,N_37856);
and U44233 (N_44233,N_30799,N_38544);
nand U44234 (N_44234,N_35240,N_32321);
or U44235 (N_44235,N_33977,N_31728);
and U44236 (N_44236,N_39143,N_37888);
and U44237 (N_44237,N_36873,N_31972);
or U44238 (N_44238,N_39791,N_38719);
and U44239 (N_44239,N_33160,N_36828);
xnor U44240 (N_44240,N_33301,N_34401);
nand U44241 (N_44241,N_38685,N_32267);
nor U44242 (N_44242,N_37300,N_30390);
nand U44243 (N_44243,N_37693,N_37802);
nand U44244 (N_44244,N_32779,N_32588);
nand U44245 (N_44245,N_30393,N_31957);
and U44246 (N_44246,N_35648,N_36758);
and U44247 (N_44247,N_39801,N_38628);
or U44248 (N_44248,N_31274,N_37018);
or U44249 (N_44249,N_39560,N_31694);
xnor U44250 (N_44250,N_33060,N_34407);
or U44251 (N_44251,N_33702,N_37243);
nand U44252 (N_44252,N_35968,N_32338);
nand U44253 (N_44253,N_38299,N_35271);
xnor U44254 (N_44254,N_35433,N_34933);
nor U44255 (N_44255,N_32462,N_39144);
xnor U44256 (N_44256,N_30447,N_38130);
xnor U44257 (N_44257,N_32387,N_38337);
nor U44258 (N_44258,N_39298,N_39846);
or U44259 (N_44259,N_32807,N_38013);
nand U44260 (N_44260,N_34938,N_33277);
or U44261 (N_44261,N_33027,N_36352);
nor U44262 (N_44262,N_33084,N_30559);
nand U44263 (N_44263,N_35482,N_32540);
xnor U44264 (N_44264,N_36104,N_37380);
and U44265 (N_44265,N_35128,N_32504);
or U44266 (N_44266,N_37175,N_39626);
xnor U44267 (N_44267,N_37815,N_37809);
nand U44268 (N_44268,N_36682,N_38839);
or U44269 (N_44269,N_38361,N_39460);
and U44270 (N_44270,N_35391,N_33920);
nand U44271 (N_44271,N_38978,N_35715);
and U44272 (N_44272,N_36126,N_34269);
xor U44273 (N_44273,N_35700,N_39977);
and U44274 (N_44274,N_33152,N_30335);
or U44275 (N_44275,N_38694,N_35048);
nand U44276 (N_44276,N_37015,N_36913);
and U44277 (N_44277,N_32653,N_36652);
or U44278 (N_44278,N_39439,N_35220);
and U44279 (N_44279,N_34184,N_31880);
nand U44280 (N_44280,N_37060,N_39102);
nand U44281 (N_44281,N_34225,N_35225);
or U44282 (N_44282,N_32531,N_33421);
xor U44283 (N_44283,N_33547,N_31549);
or U44284 (N_44284,N_30413,N_34489);
nor U44285 (N_44285,N_32584,N_37012);
nand U44286 (N_44286,N_37956,N_39575);
and U44287 (N_44287,N_31966,N_34115);
or U44288 (N_44288,N_31550,N_33185);
or U44289 (N_44289,N_34824,N_34337);
or U44290 (N_44290,N_32834,N_38711);
nor U44291 (N_44291,N_31978,N_39083);
nor U44292 (N_44292,N_33094,N_36009);
or U44293 (N_44293,N_37107,N_38530);
nand U44294 (N_44294,N_39032,N_37488);
xor U44295 (N_44295,N_36183,N_36080);
xor U44296 (N_44296,N_34661,N_37767);
nand U44297 (N_44297,N_36889,N_38117);
and U44298 (N_44298,N_33760,N_39050);
nand U44299 (N_44299,N_39651,N_36430);
and U44300 (N_44300,N_32075,N_34764);
and U44301 (N_44301,N_36100,N_37332);
xnor U44302 (N_44302,N_38569,N_31162);
and U44303 (N_44303,N_30871,N_35253);
nor U44304 (N_44304,N_34009,N_35807);
xnor U44305 (N_44305,N_35591,N_38045);
nand U44306 (N_44306,N_34453,N_34892);
and U44307 (N_44307,N_33270,N_35587);
nor U44308 (N_44308,N_38241,N_30643);
or U44309 (N_44309,N_31339,N_39607);
xor U44310 (N_44310,N_32300,N_33491);
or U44311 (N_44311,N_37630,N_34456);
xnor U44312 (N_44312,N_34737,N_30299);
nand U44313 (N_44313,N_32336,N_32449);
and U44314 (N_44314,N_33690,N_30408);
or U44315 (N_44315,N_36065,N_37682);
nor U44316 (N_44316,N_31702,N_33151);
or U44317 (N_44317,N_37814,N_37110);
nor U44318 (N_44318,N_39644,N_31097);
xnor U44319 (N_44319,N_38389,N_31043);
or U44320 (N_44320,N_39811,N_32438);
nor U44321 (N_44321,N_36964,N_37309);
nor U44322 (N_44322,N_33913,N_32959);
nor U44323 (N_44323,N_39004,N_34906);
nor U44324 (N_44324,N_36642,N_38236);
xor U44325 (N_44325,N_34792,N_30595);
xnor U44326 (N_44326,N_37025,N_37086);
or U44327 (N_44327,N_36865,N_36612);
and U44328 (N_44328,N_38913,N_30978);
or U44329 (N_44329,N_30765,N_31119);
nand U44330 (N_44330,N_36894,N_30179);
or U44331 (N_44331,N_31548,N_30019);
nand U44332 (N_44332,N_38795,N_33823);
nor U44333 (N_44333,N_33892,N_36156);
nand U44334 (N_44334,N_39641,N_31930);
and U44335 (N_44335,N_37594,N_33182);
nor U44336 (N_44336,N_36839,N_30024);
nand U44337 (N_44337,N_32640,N_35580);
or U44338 (N_44338,N_31235,N_31656);
and U44339 (N_44339,N_39135,N_34703);
and U44340 (N_44340,N_38633,N_37730);
nor U44341 (N_44341,N_37196,N_31498);
nor U44342 (N_44342,N_30046,N_39572);
xnor U44343 (N_44343,N_35133,N_31246);
nor U44344 (N_44344,N_34185,N_30945);
or U44345 (N_44345,N_34790,N_38520);
or U44346 (N_44346,N_31287,N_31981);
and U44347 (N_44347,N_34093,N_35091);
xor U44348 (N_44348,N_35263,N_38728);
xor U44349 (N_44349,N_30312,N_34878);
nand U44350 (N_44350,N_35234,N_36414);
nand U44351 (N_44351,N_39446,N_37470);
and U44352 (N_44352,N_37024,N_33838);
and U44353 (N_44353,N_32529,N_38645);
and U44354 (N_44354,N_30724,N_30772);
or U44355 (N_44355,N_32810,N_37440);
nand U44356 (N_44356,N_36656,N_33177);
or U44357 (N_44357,N_32458,N_31417);
xor U44358 (N_44358,N_33642,N_35759);
nand U44359 (N_44359,N_35918,N_31456);
xnor U44360 (N_44360,N_34063,N_30953);
nor U44361 (N_44361,N_32824,N_37568);
xor U44362 (N_44362,N_36233,N_36765);
and U44363 (N_44363,N_39236,N_32660);
or U44364 (N_44364,N_34486,N_35863);
nand U44365 (N_44365,N_31767,N_32592);
xnor U44366 (N_44366,N_38610,N_39158);
nand U44367 (N_44367,N_37457,N_39217);
or U44368 (N_44368,N_39919,N_36424);
nor U44369 (N_44369,N_33358,N_34692);
nor U44370 (N_44370,N_35488,N_31691);
or U44371 (N_44371,N_30076,N_30798);
xor U44372 (N_44372,N_32758,N_37462);
and U44373 (N_44373,N_32533,N_36570);
or U44374 (N_44374,N_36891,N_36492);
nand U44375 (N_44375,N_34465,N_32130);
and U44376 (N_44376,N_35628,N_39984);
nand U44377 (N_44377,N_34046,N_33409);
or U44378 (N_44378,N_35716,N_32385);
xnor U44379 (N_44379,N_32831,N_34861);
nor U44380 (N_44380,N_32820,N_32908);
and U44381 (N_44381,N_35859,N_37560);
or U44382 (N_44382,N_39749,N_39932);
nor U44383 (N_44383,N_34837,N_30176);
or U44384 (N_44384,N_31426,N_33606);
and U44385 (N_44385,N_31355,N_37750);
nor U44386 (N_44386,N_33518,N_37298);
nor U44387 (N_44387,N_31553,N_32411);
nand U44388 (N_44388,N_35388,N_30627);
nand U44389 (N_44389,N_38311,N_30325);
xnor U44390 (N_44390,N_31640,N_30922);
or U44391 (N_44391,N_33201,N_34007);
and U44392 (N_44392,N_36836,N_30158);
nand U44393 (N_44393,N_33850,N_34342);
nand U44394 (N_44394,N_35136,N_34150);
and U44395 (N_44395,N_39567,N_31988);
nand U44396 (N_44396,N_34593,N_30129);
nand U44397 (N_44397,N_30289,N_39993);
and U44398 (N_44398,N_36835,N_32409);
nor U44399 (N_44399,N_33887,N_39819);
xnor U44400 (N_44400,N_30631,N_30392);
or U44401 (N_44401,N_32340,N_38738);
xor U44402 (N_44402,N_33210,N_36151);
or U44403 (N_44403,N_30025,N_36015);
or U44404 (N_44404,N_37362,N_37780);
nor U44405 (N_44405,N_37171,N_33909);
nand U44406 (N_44406,N_35508,N_36762);
or U44407 (N_44407,N_34006,N_36330);
or U44408 (N_44408,N_32571,N_35027);
nor U44409 (N_44409,N_34323,N_33063);
and U44410 (N_44410,N_34832,N_36382);
or U44411 (N_44411,N_39619,N_30452);
and U44412 (N_44412,N_31405,N_38982);
or U44413 (N_44413,N_33371,N_30694);
nor U44414 (N_44414,N_39755,N_33230);
or U44415 (N_44415,N_38344,N_30708);
nor U44416 (N_44416,N_32784,N_33432);
and U44417 (N_44417,N_39857,N_38290);
nor U44418 (N_44418,N_31874,N_38621);
or U44419 (N_44419,N_35469,N_39624);
xor U44420 (N_44420,N_31937,N_39482);
xnor U44421 (N_44421,N_38865,N_36196);
and U44422 (N_44422,N_38534,N_31684);
and U44423 (N_44423,N_32354,N_38843);
nor U44424 (N_44424,N_35197,N_35894);
xnor U44425 (N_44425,N_38185,N_33507);
xor U44426 (N_44426,N_30659,N_37949);
nand U44427 (N_44427,N_30622,N_30091);
nor U44428 (N_44428,N_33072,N_39578);
or U44429 (N_44429,N_37272,N_31067);
xor U44430 (N_44430,N_31622,N_39875);
or U44431 (N_44431,N_38644,N_30596);
and U44432 (N_44432,N_33603,N_39968);
or U44433 (N_44433,N_33768,N_35267);
nand U44434 (N_44434,N_36410,N_33922);
nor U44435 (N_44435,N_32051,N_30402);
nor U44436 (N_44436,N_32083,N_36299);
xor U44437 (N_44437,N_39161,N_34427);
and U44438 (N_44438,N_31292,N_38687);
or U44439 (N_44439,N_36681,N_35001);
xnor U44440 (N_44440,N_38805,N_39473);
xnor U44441 (N_44441,N_33455,N_36329);
nor U44442 (N_44442,N_34057,N_33928);
and U44443 (N_44443,N_37792,N_34842);
and U44444 (N_44444,N_36189,N_37014);
nand U44445 (N_44445,N_33898,N_32545);
or U44446 (N_44446,N_30458,N_30840);
nand U44447 (N_44447,N_34384,N_35507);
nand U44448 (N_44448,N_33149,N_33332);
nand U44449 (N_44449,N_30096,N_32361);
xor U44450 (N_44450,N_38800,N_36720);
xnor U44451 (N_44451,N_30320,N_31262);
nand U44452 (N_44452,N_33279,N_37512);
nand U44453 (N_44453,N_37082,N_38861);
and U44454 (N_44454,N_37458,N_39796);
and U44455 (N_44455,N_35895,N_39345);
and U44456 (N_44456,N_37716,N_30967);
nor U44457 (N_44457,N_36310,N_35697);
nor U44458 (N_44458,N_30137,N_35532);
or U44459 (N_44459,N_30420,N_33879);
xnor U44460 (N_44460,N_36914,N_33965);
xnor U44461 (N_44461,N_35740,N_35905);
xnor U44462 (N_44462,N_37437,N_33310);
and U44463 (N_44463,N_39401,N_33176);
or U44464 (N_44464,N_33205,N_36354);
nand U44465 (N_44465,N_32859,N_33266);
xor U44466 (N_44466,N_33698,N_36053);
nand U44467 (N_44467,N_37330,N_37011);
nor U44468 (N_44468,N_30350,N_34157);
xnor U44469 (N_44469,N_37351,N_36691);
nor U44470 (N_44470,N_39753,N_36304);
and U44471 (N_44471,N_33180,N_32623);
and U44472 (N_44472,N_32487,N_36158);
and U44473 (N_44473,N_39525,N_36399);
xnor U44474 (N_44474,N_34665,N_34414);
and U44475 (N_44475,N_35248,N_31215);
nor U44476 (N_44476,N_38551,N_30018);
nor U44477 (N_44477,N_35064,N_32401);
or U44478 (N_44478,N_39914,N_32669);
nand U44479 (N_44479,N_30611,N_34392);
or U44480 (N_44480,N_38787,N_30780);
or U44481 (N_44481,N_31249,N_37377);
nand U44482 (N_44482,N_37773,N_36778);
xor U44483 (N_44483,N_36033,N_38985);
nor U44484 (N_44484,N_34748,N_39259);
nand U44485 (N_44485,N_32251,N_34450);
xor U44486 (N_44486,N_32066,N_36038);
and U44487 (N_44487,N_33168,N_32245);
or U44488 (N_44488,N_30828,N_33593);
or U44489 (N_44489,N_38418,N_31716);
xnor U44490 (N_44490,N_39428,N_32486);
nor U44491 (N_44491,N_36910,N_36875);
nor U44492 (N_44492,N_31136,N_31982);
nor U44493 (N_44493,N_30620,N_32512);
or U44494 (N_44494,N_33130,N_37305);
xnor U44495 (N_44495,N_30982,N_33378);
or U44496 (N_44496,N_38840,N_34870);
and U44497 (N_44497,N_37240,N_30443);
xor U44498 (N_44498,N_36362,N_30436);
nor U44499 (N_44499,N_34646,N_31873);
and U44500 (N_44500,N_35367,N_38782);
xor U44501 (N_44501,N_35961,N_34612);
and U44502 (N_44502,N_33033,N_39421);
xnor U44503 (N_44503,N_38118,N_31740);
xnor U44504 (N_44504,N_34844,N_35280);
nand U44505 (N_44505,N_32002,N_39111);
and U44506 (N_44506,N_37946,N_35332);
nand U44507 (N_44507,N_34645,N_37047);
and U44508 (N_44508,N_38123,N_39574);
and U44509 (N_44509,N_39363,N_36683);
nand U44510 (N_44510,N_35459,N_39657);
xnor U44511 (N_44511,N_31532,N_38931);
nor U44512 (N_44512,N_31264,N_33035);
xnor U44513 (N_44513,N_33629,N_39044);
or U44514 (N_44514,N_32094,N_33834);
nand U44515 (N_44515,N_33561,N_34756);
xnor U44516 (N_44516,N_31064,N_34967);
and U44517 (N_44517,N_37061,N_38341);
xor U44518 (N_44518,N_38439,N_32816);
or U44519 (N_44519,N_36442,N_30607);
or U44520 (N_44520,N_31641,N_31825);
nor U44521 (N_44521,N_37740,N_31642);
and U44522 (N_44522,N_30961,N_32025);
and U44523 (N_44523,N_31718,N_38546);
xnor U44524 (N_44524,N_39254,N_34940);
nor U44525 (N_44525,N_31492,N_31535);
xnor U44526 (N_44526,N_32731,N_39402);
nand U44527 (N_44527,N_32984,N_31621);
or U44528 (N_44528,N_31449,N_34572);
nor U44529 (N_44529,N_31714,N_37399);
or U44530 (N_44530,N_37227,N_39368);
xnor U44531 (N_44531,N_38377,N_33853);
nand U44532 (N_44532,N_34617,N_30618);
xor U44533 (N_44533,N_34396,N_32901);
xor U44534 (N_44534,N_34348,N_30235);
nor U44535 (N_44535,N_39905,N_37679);
nor U44536 (N_44536,N_35362,N_34610);
nor U44537 (N_44537,N_38521,N_34855);
xor U44538 (N_44538,N_31271,N_39013);
or U44539 (N_44539,N_37123,N_33320);
nor U44540 (N_44540,N_30782,N_36341);
nor U44541 (N_44541,N_31071,N_35093);
or U44542 (N_44542,N_35560,N_37218);
xor U44543 (N_44543,N_35938,N_34283);
and U44544 (N_44544,N_32059,N_35453);
nor U44545 (N_44545,N_32266,N_35017);
nor U44546 (N_44546,N_34263,N_37810);
nor U44547 (N_44547,N_36062,N_39611);
nand U44548 (N_44548,N_35809,N_36181);
or U44549 (N_44549,N_34086,N_34736);
nor U44550 (N_44550,N_30855,N_31531);
xor U44551 (N_44551,N_31288,N_32560);
nor U44552 (N_44552,N_33164,N_32503);
or U44553 (N_44553,N_37980,N_34690);
or U44554 (N_44554,N_30975,N_31329);
or U44555 (N_44555,N_37147,N_30397);
nor U44556 (N_44556,N_31275,N_35110);
xnor U44557 (N_44557,N_39468,N_39423);
xor U44558 (N_44558,N_37583,N_35599);
nor U44559 (N_44559,N_33138,N_39375);
nand U44560 (N_44560,N_35673,N_35661);
and U44561 (N_44561,N_30566,N_35327);
or U44562 (N_44562,N_32721,N_33878);
xnor U44563 (N_44563,N_37526,N_37445);
xnor U44564 (N_44564,N_36548,N_36427);
and U44565 (N_44565,N_34620,N_31467);
nand U44566 (N_44566,N_39735,N_36409);
nand U44567 (N_44567,N_36054,N_35343);
and U44568 (N_44568,N_37755,N_39387);
nor U44569 (N_44569,N_32591,N_33866);
nand U44570 (N_44570,N_34695,N_38936);
xnor U44571 (N_44571,N_34023,N_36981);
nor U44572 (N_44572,N_35147,N_38007);
xor U44573 (N_44573,N_36583,N_31781);
nand U44574 (N_44574,N_36073,N_31845);
nor U44575 (N_44575,N_39803,N_32650);
xor U44576 (N_44576,N_34669,N_37688);
nand U44577 (N_44577,N_32993,N_38282);
nand U44578 (N_44578,N_30380,N_34487);
nor U44579 (N_44579,N_35475,N_36965);
or U44580 (N_44580,N_36809,N_39833);
nor U44581 (N_44581,N_35996,N_31416);
xnor U44582 (N_44582,N_34948,N_37516);
and U44583 (N_44583,N_38467,N_31013);
and U44584 (N_44584,N_30021,N_37697);
nor U44585 (N_44585,N_38998,N_36638);
nand U44586 (N_44586,N_35390,N_36575);
xor U44587 (N_44587,N_37562,N_32163);
nor U44588 (N_44588,N_35865,N_31954);
and U44589 (N_44589,N_34550,N_30440);
or U44590 (N_44590,N_38844,N_32376);
nand U44591 (N_44591,N_34266,N_37891);
xnor U44592 (N_44592,N_37220,N_33575);
nor U44593 (N_44593,N_39220,N_39770);
nand U44594 (N_44594,N_35623,N_30266);
nor U44595 (N_44595,N_30345,N_37808);
nor U44596 (N_44596,N_36107,N_32064);
nand U44597 (N_44597,N_30862,N_34721);
or U44598 (N_44598,N_30791,N_38172);
xnor U44599 (N_44599,N_35105,N_37624);
xor U44600 (N_44600,N_34445,N_39878);
or U44601 (N_44601,N_36635,N_39165);
and U44602 (N_44602,N_35756,N_33119);
nor U44603 (N_44603,N_32616,N_36900);
nand U44604 (N_44604,N_32776,N_35936);
xor U44605 (N_44605,N_31300,N_32748);
nand U44606 (N_44606,N_39488,N_38794);
or U44607 (N_44607,N_31312,N_31562);
and U44608 (N_44608,N_31412,N_30789);
xnor U44609 (N_44609,N_33386,N_39673);
xnor U44610 (N_44610,N_38891,N_34640);
xnor U44611 (N_44611,N_37569,N_32370);
or U44612 (N_44612,N_30297,N_30416);
or U44613 (N_44613,N_34746,N_30081);
or U44614 (N_44614,N_31237,N_33949);
and U44615 (N_44615,N_37911,N_37779);
nand U44616 (N_44616,N_30988,N_30560);
xnor U44617 (N_44617,N_32337,N_38768);
or U44618 (N_44618,N_39656,N_33881);
nor U44619 (N_44619,N_32947,N_33065);
or U44620 (N_44620,N_33187,N_34379);
nor U44621 (N_44621,N_32554,N_36976);
xnor U44622 (N_44622,N_32315,N_38459);
xnor U44623 (N_44623,N_31483,N_30342);
xnor U44624 (N_44624,N_32417,N_36984);
xor U44625 (N_44625,N_35811,N_38247);
xor U44626 (N_44626,N_36392,N_31160);
and U44627 (N_44627,N_31613,N_30031);
xnor U44628 (N_44628,N_32353,N_30167);
xor U44629 (N_44629,N_31358,N_30177);
or U44630 (N_44630,N_35778,N_30751);
xor U44631 (N_44631,N_30839,N_31144);
and U44632 (N_44632,N_36634,N_34807);
or U44633 (N_44633,N_34359,N_37224);
nand U44634 (N_44634,N_37898,N_33274);
xnor U44635 (N_44635,N_37611,N_34879);
nand U44636 (N_44636,N_38370,N_30933);
nand U44637 (N_44637,N_33242,N_30305);
nand U44638 (N_44638,N_37774,N_39725);
nand U44639 (N_44639,N_37034,N_32084);
nand U44640 (N_44640,N_35923,N_31651);
nor U44641 (N_44641,N_31935,N_37366);
nand U44642 (N_44642,N_34930,N_36131);
nor U44643 (N_44643,N_34977,N_35650);
xor U44644 (N_44644,N_33463,N_37195);
xor U44645 (N_44645,N_36475,N_32769);
and U44646 (N_44646,N_31335,N_31220);
and U44647 (N_44647,N_30940,N_31938);
nand U44648 (N_44648,N_39877,N_30638);
and U44649 (N_44649,N_38435,N_37928);
nand U44650 (N_44650,N_30253,N_32950);
or U44651 (N_44651,N_32551,N_32032);
nand U44652 (N_44652,N_38838,N_38345);
xnor U44653 (N_44653,N_33521,N_39322);
nor U44654 (N_44654,N_34162,N_31737);
and U44655 (N_44655,N_34492,N_32249);
and U44656 (N_44656,N_36001,N_31452);
xor U44657 (N_44657,N_37205,N_35592);
nor U44658 (N_44658,N_39629,N_34395);
and U44659 (N_44659,N_35387,N_32792);
nand U44660 (N_44660,N_39497,N_30655);
xor U44661 (N_44661,N_37747,N_32949);
nand U44662 (N_44662,N_38053,N_33394);
xnor U44663 (N_44663,N_33190,N_33356);
nor U44664 (N_44664,N_37883,N_33989);
nand U44665 (N_44665,N_33447,N_39911);
nor U44666 (N_44666,N_38356,N_30381);
nor U44667 (N_44667,N_30359,N_30273);
or U44668 (N_44668,N_34357,N_31478);
nor U44669 (N_44669,N_32119,N_35117);
nor U44670 (N_44670,N_36895,N_37434);
xor U44671 (N_44671,N_36821,N_31042);
and U44672 (N_44672,N_38881,N_30706);
nand U44673 (N_44673,N_33782,N_38211);
nand U44674 (N_44674,N_33526,N_36176);
and U44675 (N_44675,N_33010,N_31294);
nand U44676 (N_44676,N_36057,N_31196);
nor U44677 (N_44677,N_33817,N_35277);
and U44678 (N_44678,N_36597,N_38137);
xnor U44679 (N_44679,N_33170,N_32762);
nand U44680 (N_44680,N_38586,N_36108);
or U44681 (N_44681,N_34584,N_32897);
xnor U44682 (N_44682,N_36814,N_35984);
and U44683 (N_44683,N_32324,N_33811);
or U44684 (N_44684,N_39209,N_30022);
nor U44685 (N_44685,N_37479,N_34189);
xor U44686 (N_44686,N_30228,N_32789);
and U44687 (N_44687,N_32005,N_38637);
nor U44688 (N_44688,N_36963,N_35636);
nor U44689 (N_44689,N_35276,N_39364);
xnor U44690 (N_44690,N_30346,N_30316);
or U44691 (N_44691,N_33286,N_33638);
and U44692 (N_44692,N_38487,N_34947);
or U44693 (N_44693,N_36556,N_30842);
and U44694 (N_44694,N_32473,N_32672);
nor U44695 (N_44695,N_34886,N_33222);
nor U44696 (N_44696,N_34559,N_36543);
nand U44697 (N_44697,N_30730,N_38302);
and U44698 (N_44698,N_35565,N_36698);
xor U44699 (N_44699,N_39706,N_34860);
and U44700 (N_44700,N_33022,N_34974);
xnor U44701 (N_44701,N_31448,N_32992);
and U44702 (N_44702,N_31022,N_39782);
or U44703 (N_44703,N_30104,N_35178);
xor U44704 (N_44704,N_37252,N_36011);
xor U44705 (N_44705,N_34891,N_34964);
or U44706 (N_44706,N_30582,N_36367);
and U44707 (N_44707,N_34451,N_38216);
nor U44708 (N_44708,N_35739,N_38706);
nand U44709 (N_44709,N_30488,N_38821);
and U44710 (N_44710,N_39223,N_36526);
nand U44711 (N_44711,N_38391,N_34118);
and U44712 (N_44712,N_36152,N_34058);
and U44713 (N_44713,N_33480,N_38855);
xor U44714 (N_44714,N_39920,N_33359);
and U44715 (N_44715,N_36748,N_30972);
and U44716 (N_44716,N_32941,N_37538);
or U44717 (N_44717,N_36161,N_32303);
nand U44718 (N_44718,N_32279,N_34787);
nand U44719 (N_44719,N_36260,N_32062);
or U44720 (N_44720,N_34259,N_33233);
and U44721 (N_44721,N_30249,N_32661);
or U44722 (N_44722,N_37372,N_33730);
nand U44723 (N_44723,N_39444,N_36145);
nor U44724 (N_44724,N_39207,N_37043);
nor U44725 (N_44725,N_31359,N_35668);
xnor U44726 (N_44726,N_30697,N_35659);
nor U44727 (N_44727,N_34508,N_33174);
and U44728 (N_44728,N_37927,N_37542);
and U44729 (N_44729,N_34505,N_39557);
xnor U44730 (N_44730,N_36277,N_34618);
and U44731 (N_44731,N_36560,N_34782);
and U44732 (N_44732,N_30429,N_30374);
xnor U44733 (N_44733,N_38027,N_32437);
nor U44734 (N_44734,N_32097,N_36227);
or U44735 (N_44735,N_30281,N_38265);
nor U44736 (N_44736,N_32521,N_30329);
or U44737 (N_44737,N_33038,N_34638);
and U44738 (N_44738,N_31909,N_36286);
nand U44739 (N_44739,N_34694,N_31073);
nor U44740 (N_44740,N_30881,N_30152);
nor U44741 (N_44741,N_35854,N_34993);
and U44742 (N_44742,N_33605,N_32131);
xor U44743 (N_44743,N_37058,N_35730);
and U44744 (N_44744,N_34239,N_32723);
nand U44745 (N_44745,N_30849,N_30276);
xor U44746 (N_44746,N_39095,N_30921);
nor U44747 (N_44747,N_38465,N_34361);
or U44748 (N_44748,N_38984,N_35417);
nor U44749 (N_44749,N_38324,N_32254);
nand U44750 (N_44750,N_35941,N_31083);
and U44751 (N_44751,N_34314,N_30874);
xnor U44752 (N_44752,N_35381,N_35511);
xnor U44753 (N_44753,N_30900,N_37557);
nand U44754 (N_44754,N_36394,N_35551);
and U44755 (N_44755,N_39054,N_39412);
nor U44756 (N_44756,N_33670,N_33555);
or U44757 (N_44757,N_39935,N_38858);
xor U44758 (N_44758,N_32133,N_30576);
xor U44759 (N_44759,N_38689,N_36489);
and U44760 (N_44760,N_37129,N_35872);
or U44761 (N_44761,N_39369,N_33718);
and U44762 (N_44762,N_37090,N_31434);
or U44763 (N_44763,N_35727,N_38830);
and U44764 (N_44764,N_33640,N_33622);
or U44765 (N_44765,N_32956,N_34182);
nand U44766 (N_44766,N_37013,N_38961);
nand U44767 (N_44767,N_30976,N_31045);
nor U44768 (N_44768,N_32216,N_38153);
nand U44769 (N_44769,N_32422,N_33694);
nor U44770 (N_44770,N_39405,N_30363);
or U44771 (N_44771,N_35184,N_37213);
nor U44772 (N_44772,N_33052,N_33280);
xor U44773 (N_44773,N_39898,N_32717);
nor U44774 (N_44774,N_31711,N_36170);
or U44775 (N_44775,N_39038,N_30271);
xnor U44776 (N_44776,N_32755,N_33115);
nor U44777 (N_44777,N_36951,N_36818);
and U44778 (N_44778,N_35338,N_35383);
nand U44779 (N_44779,N_36499,N_34139);
xnor U44780 (N_44780,N_34334,N_36578);
nand U44781 (N_44781,N_38168,N_30479);
nand U44782 (N_44782,N_33883,N_36961);
nand U44783 (N_44783,N_36787,N_37225);
xnor U44784 (N_44784,N_39890,N_34247);
xor U44785 (N_44785,N_30217,N_39011);
nand U44786 (N_44786,N_34850,N_30646);
xor U44787 (N_44787,N_35335,N_34705);
xnor U44788 (N_44788,N_35164,N_39417);
nor U44789 (N_44789,N_31916,N_39061);
xnor U44790 (N_44790,N_38811,N_34216);
or U44791 (N_44791,N_32074,N_37414);
or U44792 (N_44792,N_36370,N_33577);
nor U44793 (N_44793,N_31485,N_30774);
xor U44794 (N_44794,N_38816,N_31167);
and U44795 (N_44795,N_33227,N_34097);
nand U44796 (N_44796,N_36792,N_33554);
xor U44797 (N_44797,N_39200,N_34272);
nand U44798 (N_44798,N_31689,N_33862);
nand U44799 (N_44799,N_30805,N_30063);
or U44800 (N_44800,N_30647,N_36538);
nand U44801 (N_44801,N_31907,N_33100);
nor U44802 (N_44802,N_36343,N_39519);
or U44803 (N_44803,N_31297,N_37869);
nand U44804 (N_44804,N_37288,N_32029);
and U44805 (N_44805,N_32595,N_31544);
xor U44806 (N_44806,N_32870,N_35682);
and U44807 (N_44807,N_35542,N_32973);
nor U44808 (N_44808,N_33249,N_34817);
or U44809 (N_44809,N_39116,N_36374);
nand U44810 (N_44810,N_36503,N_31875);
or U44811 (N_44811,N_30684,N_30733);
xnor U44812 (N_44812,N_35000,N_37514);
nor U44813 (N_44813,N_36050,N_38642);
or U44814 (N_44814,N_32246,N_37805);
and U44815 (N_44815,N_31810,N_30209);
nand U44816 (N_44816,N_30379,N_38223);
xnor U44817 (N_44817,N_31007,N_33810);
or U44818 (N_44818,N_35249,N_33722);
or U44819 (N_44819,N_32318,N_33448);
nand U44820 (N_44820,N_32123,N_39623);
xor U44821 (N_44821,N_30536,N_38334);
nor U44822 (N_44822,N_31350,N_31945);
nand U44823 (N_44823,N_38005,N_39576);
xnor U44824 (N_44824,N_30648,N_36863);
nand U44825 (N_44825,N_36443,N_32574);
or U44826 (N_44826,N_34718,N_37979);
xor U44827 (N_44827,N_36502,N_36359);
and U44828 (N_44828,N_38319,N_30256);
nand U44829 (N_44829,N_37439,N_35738);
or U44830 (N_44830,N_36318,N_36687);
nor U44831 (N_44831,N_36238,N_39224);
nor U44832 (N_44832,N_34124,N_39370);
or U44833 (N_44833,N_32573,N_37546);
nor U44834 (N_44834,N_30023,N_33796);
and U44835 (N_44835,N_39895,N_39794);
xnor U44836 (N_44836,N_32232,N_31990);
nor U44837 (N_44837,N_34437,N_34305);
or U44838 (N_44838,N_36447,N_30165);
nand U44839 (N_44839,N_34413,N_32611);
xor U44840 (N_44840,N_39034,N_37844);
nand U44841 (N_44841,N_36328,N_33636);
and U44842 (N_44842,N_33204,N_34181);
and U44843 (N_44843,N_35037,N_35896);
or U44844 (N_44844,N_33681,N_33209);
and U44845 (N_44845,N_39081,N_39461);
and U44846 (N_44846,N_33268,N_31507);
and U44847 (N_44847,N_37892,N_34494);
or U44848 (N_44848,N_31331,N_33533);
nand U44849 (N_44849,N_39966,N_34719);
or U44850 (N_44850,N_38372,N_31717);
xnor U44851 (N_44851,N_30745,N_34641);
nand U44852 (N_44852,N_39301,N_31969);
nor U44853 (N_44853,N_33741,N_37743);
nand U44854 (N_44854,N_33186,N_33961);
xor U44855 (N_44855,N_34102,N_32352);
xnor U44856 (N_44856,N_39535,N_36262);
xnor U44857 (N_44857,N_37789,N_33573);
or U44858 (N_44858,N_30186,N_31752);
nor U44859 (N_44859,N_33737,N_30886);
nand U44860 (N_44860,N_35629,N_39636);
nand U44861 (N_44861,N_34812,N_31530);
xnor U44862 (N_44862,N_31939,N_37250);
nand U44863 (N_44863,N_39684,N_37602);
or U44864 (N_44864,N_30713,N_36032);
nor U44865 (N_44865,N_39020,N_31599);
nand U44866 (N_44866,N_30810,N_37751);
xor U44867 (N_44867,N_32176,N_33026);
or U44868 (N_44868,N_34060,N_36760);
or U44869 (N_44869,N_32096,N_32750);
and U44870 (N_44870,N_34592,N_38386);
or U44871 (N_44871,N_34744,N_30951);
nor U44872 (N_44872,N_38518,N_36423);
and U44873 (N_44873,N_35889,N_36160);
xor U44874 (N_44874,N_31490,N_32311);
nand U44875 (N_44875,N_35268,N_31079);
or U44876 (N_44876,N_33445,N_38295);
and U44877 (N_44877,N_31723,N_30660);
nand U44878 (N_44878,N_34928,N_32902);
and U44879 (N_44879,N_36440,N_39131);
nor U44880 (N_44880,N_31920,N_34922);
or U44881 (N_44881,N_30718,N_39943);
nand U44882 (N_44882,N_33999,N_32145);
xnor U44883 (N_44883,N_33479,N_39537);
xnor U44884 (N_44884,N_36148,N_31974);
and U44885 (N_44885,N_34732,N_30530);
xnor U44886 (N_44886,N_37536,N_37156);
nor U44887 (N_44887,N_37800,N_30575);
and U44888 (N_44888,N_36049,N_38904);
and U44889 (N_44889,N_38249,N_39016);
and U44890 (N_44890,N_36680,N_32578);
or U44891 (N_44891,N_30351,N_30836);
nand U44892 (N_44892,N_38298,N_30661);
and U44893 (N_44893,N_31657,N_38120);
or U44894 (N_44894,N_36677,N_33144);
nand U44895 (N_44895,N_39010,N_38703);
xnor U44896 (N_44896,N_38410,N_36817);
or U44897 (N_44897,N_39960,N_30120);
nor U44898 (N_44898,N_32288,N_30500);
nor U44899 (N_44899,N_30515,N_32298);
or U44900 (N_44900,N_34279,N_34080);
nor U44901 (N_44901,N_31586,N_36446);
or U44902 (N_44902,N_37576,N_30843);
nand U44903 (N_44903,N_39719,N_32639);
or U44904 (N_44904,N_33075,N_35241);
and U44905 (N_44905,N_37860,N_38684);
or U44906 (N_44906,N_33643,N_34014);
and U44907 (N_44907,N_35527,N_32918);
nor U44908 (N_44908,N_39251,N_32394);
and U44909 (N_44909,N_37203,N_37387);
or U44910 (N_44910,N_30821,N_38578);
or U44911 (N_44911,N_32448,N_30928);
xnor U44912 (N_44912,N_30173,N_36956);
xnor U44913 (N_44913,N_30589,N_33202);
nand U44914 (N_44914,N_35687,N_38752);
xor U44915 (N_44915,N_39585,N_36044);
xnor U44916 (N_44916,N_38552,N_35119);
xnor U44917 (N_44917,N_32067,N_33863);
xor U44918 (N_44918,N_33795,N_38664);
or U44919 (N_44919,N_38734,N_36250);
and U44920 (N_44920,N_37590,N_39313);
nor U44921 (N_44921,N_37448,N_31247);
nand U44922 (N_44922,N_30053,N_37307);
and U44923 (N_44923,N_38184,N_37847);
or U44924 (N_44924,N_30974,N_30110);
or U44925 (N_44925,N_38691,N_37541);
and U44926 (N_44926,N_34478,N_32876);
or U44927 (N_44927,N_34441,N_35480);
or U44928 (N_44928,N_35828,N_39959);
nor U44929 (N_44929,N_35902,N_31040);
or U44930 (N_44930,N_34975,N_32332);
xor U44931 (N_44931,N_38500,N_31949);
nor U44932 (N_44932,N_31046,N_34325);
and U44933 (N_44933,N_36752,N_31330);
xnor U44934 (N_44934,N_36962,N_30723);
nor U44935 (N_44935,N_37384,N_35190);
and U44936 (N_44936,N_36904,N_35871);
and U44937 (N_44937,N_33558,N_32099);
xnor U44938 (N_44938,N_37598,N_37721);
and U44939 (N_44939,N_31583,N_31273);
nand U44940 (N_44940,N_37537,N_31633);
or U44941 (N_44941,N_32421,N_36674);
nor U44942 (N_44942,N_31142,N_34972);
nor U44943 (N_44943,N_39720,N_33919);
xnor U44944 (N_44944,N_33415,N_32047);
nor U44945 (N_44945,N_38233,N_31918);
nand U44946 (N_44946,N_36837,N_31884);
nor U44947 (N_44947,N_37029,N_39711);
xor U44948 (N_44948,N_39025,N_35464);
nand U44949 (N_44949,N_31906,N_35639);
nand U44950 (N_44950,N_31373,N_34222);
nor U44951 (N_44951,N_34321,N_32636);
or U44952 (N_44952,N_37172,N_31379);
nand U44953 (N_44953,N_32622,N_30295);
or U44954 (N_44954,N_38497,N_39349);
nand U44955 (N_44955,N_34722,N_30161);
and U44956 (N_44956,N_34399,N_34953);
nor U44957 (N_44957,N_34319,N_31665);
or U44958 (N_44958,N_38944,N_36460);
or U44959 (N_44959,N_35295,N_38747);
xnor U44960 (N_44960,N_34340,N_35886);
nor U44961 (N_44961,N_37505,N_33244);
nand U44962 (N_44962,N_37581,N_32940);
xnor U44963 (N_44963,N_39886,N_30838);
nor U44964 (N_44964,N_31786,N_33952);
or U44965 (N_44965,N_35632,N_39028);
and U44966 (N_44966,N_32444,N_33612);
and U44967 (N_44967,N_32534,N_33962);
or U44968 (N_44968,N_36759,N_38737);
or U44969 (N_44969,N_38121,N_34310);
nand U44970 (N_44970,N_36712,N_36301);
xnor U44971 (N_44971,N_34133,N_33290);
or U44972 (N_44972,N_32706,N_37246);
nor U44973 (N_44973,N_36786,N_38890);
nand U44974 (N_44974,N_35799,N_30189);
xor U44975 (N_44975,N_32845,N_30112);
and U44976 (N_44976,N_32416,N_37629);
nand U44977 (N_44977,N_33609,N_38872);
xor U44978 (N_44978,N_30939,N_32082);
or U44979 (N_44979,N_36470,N_31493);
and U44980 (N_44980,N_36231,N_34078);
nand U44981 (N_44981,N_32240,N_32045);
or U44982 (N_44982,N_35170,N_33224);
nor U44983 (N_44983,N_34425,N_38362);
nor U44984 (N_44984,N_39500,N_31739);
and U44985 (N_44985,N_31121,N_32510);
and U44986 (N_44986,N_38758,N_36210);
or U44987 (N_44987,N_31971,N_30903);
nor U44988 (N_44988,N_35214,N_32793);
xor U44989 (N_44989,N_37776,N_35207);
xor U44990 (N_44990,N_33364,N_37619);
nand U44991 (N_44991,N_38483,N_34754);
or U44992 (N_44992,N_34350,N_32490);
and U44993 (N_44993,N_32873,N_35983);
nand U44994 (N_44994,N_33444,N_34942);
and U44995 (N_44995,N_37295,N_34915);
nand U44996 (N_44996,N_32040,N_35059);
nor U44997 (N_44997,N_35751,N_34742);
or U44998 (N_44998,N_32143,N_39621);
or U44999 (N_44999,N_36021,N_36943);
and U45000 (N_45000,N_34009,N_36516);
nor U45001 (N_45001,N_32578,N_37852);
xor U45002 (N_45002,N_33408,N_35076);
nor U45003 (N_45003,N_37576,N_34816);
and U45004 (N_45004,N_36045,N_37674);
or U45005 (N_45005,N_35250,N_32045);
nor U45006 (N_45006,N_35639,N_33968);
or U45007 (N_45007,N_32834,N_34240);
nand U45008 (N_45008,N_37931,N_32529);
nand U45009 (N_45009,N_36545,N_30869);
nand U45010 (N_45010,N_34305,N_37566);
xor U45011 (N_45011,N_36572,N_36199);
or U45012 (N_45012,N_37492,N_34164);
and U45013 (N_45013,N_37474,N_30833);
nand U45014 (N_45014,N_34393,N_36625);
nand U45015 (N_45015,N_38428,N_37514);
and U45016 (N_45016,N_39531,N_35829);
xor U45017 (N_45017,N_31145,N_36960);
nand U45018 (N_45018,N_32090,N_34543);
or U45019 (N_45019,N_38556,N_38426);
nand U45020 (N_45020,N_37408,N_34155);
nor U45021 (N_45021,N_32199,N_36384);
nor U45022 (N_45022,N_30874,N_31414);
nor U45023 (N_45023,N_36884,N_30943);
or U45024 (N_45024,N_33624,N_39648);
nand U45025 (N_45025,N_37562,N_37898);
or U45026 (N_45026,N_39787,N_36271);
nor U45027 (N_45027,N_38121,N_34763);
nor U45028 (N_45028,N_33980,N_33820);
and U45029 (N_45029,N_31745,N_37490);
and U45030 (N_45030,N_38710,N_30934);
and U45031 (N_45031,N_39203,N_34836);
xor U45032 (N_45032,N_32983,N_37252);
or U45033 (N_45033,N_37594,N_32716);
xor U45034 (N_45034,N_39427,N_34544);
nand U45035 (N_45035,N_37228,N_39837);
and U45036 (N_45036,N_31973,N_33011);
nand U45037 (N_45037,N_35253,N_39836);
or U45038 (N_45038,N_38831,N_30736);
or U45039 (N_45039,N_32445,N_32922);
or U45040 (N_45040,N_38679,N_30289);
xor U45041 (N_45041,N_39278,N_37635);
and U45042 (N_45042,N_33757,N_36139);
and U45043 (N_45043,N_32583,N_35928);
xnor U45044 (N_45044,N_35316,N_32198);
nor U45045 (N_45045,N_38708,N_36115);
and U45046 (N_45046,N_32419,N_31634);
or U45047 (N_45047,N_32791,N_36666);
nor U45048 (N_45048,N_37210,N_31798);
nor U45049 (N_45049,N_36963,N_36936);
and U45050 (N_45050,N_33692,N_37332);
nor U45051 (N_45051,N_30691,N_36035);
and U45052 (N_45052,N_35943,N_35803);
and U45053 (N_45053,N_32461,N_34882);
and U45054 (N_45054,N_36130,N_34469);
xor U45055 (N_45055,N_31077,N_38098);
xnor U45056 (N_45056,N_35824,N_38375);
or U45057 (N_45057,N_37303,N_31886);
nor U45058 (N_45058,N_33035,N_36561);
xnor U45059 (N_45059,N_33182,N_34880);
or U45060 (N_45060,N_38239,N_36418);
or U45061 (N_45061,N_39611,N_38882);
or U45062 (N_45062,N_36223,N_32612);
xnor U45063 (N_45063,N_39176,N_39533);
and U45064 (N_45064,N_30122,N_30110);
nand U45065 (N_45065,N_37656,N_38470);
or U45066 (N_45066,N_35640,N_39690);
or U45067 (N_45067,N_38355,N_37356);
nand U45068 (N_45068,N_37744,N_32275);
or U45069 (N_45069,N_35599,N_34450);
or U45070 (N_45070,N_32016,N_35847);
and U45071 (N_45071,N_30194,N_32092);
and U45072 (N_45072,N_35766,N_39572);
nor U45073 (N_45073,N_38263,N_31222);
xor U45074 (N_45074,N_33258,N_38004);
or U45075 (N_45075,N_35409,N_31159);
nand U45076 (N_45076,N_33202,N_30606);
nand U45077 (N_45077,N_39835,N_34717);
and U45078 (N_45078,N_39423,N_32523);
nand U45079 (N_45079,N_34663,N_33146);
and U45080 (N_45080,N_30298,N_37239);
nand U45081 (N_45081,N_39669,N_37496);
or U45082 (N_45082,N_34422,N_33074);
or U45083 (N_45083,N_30130,N_36816);
nor U45084 (N_45084,N_37546,N_32062);
xnor U45085 (N_45085,N_38707,N_38531);
nor U45086 (N_45086,N_35780,N_34998);
xor U45087 (N_45087,N_30498,N_32683);
xnor U45088 (N_45088,N_37735,N_33999);
or U45089 (N_45089,N_30731,N_32905);
and U45090 (N_45090,N_31188,N_31817);
and U45091 (N_45091,N_30157,N_34605);
xnor U45092 (N_45092,N_39152,N_30695);
nor U45093 (N_45093,N_37116,N_35571);
nor U45094 (N_45094,N_36571,N_39883);
nor U45095 (N_45095,N_30631,N_31917);
nand U45096 (N_45096,N_32851,N_35261);
or U45097 (N_45097,N_38486,N_38225);
xor U45098 (N_45098,N_31197,N_38573);
xnor U45099 (N_45099,N_34544,N_38510);
and U45100 (N_45100,N_31986,N_31951);
nand U45101 (N_45101,N_38541,N_34539);
or U45102 (N_45102,N_35325,N_39988);
and U45103 (N_45103,N_32941,N_31598);
or U45104 (N_45104,N_38016,N_36332);
or U45105 (N_45105,N_36740,N_30600);
or U45106 (N_45106,N_32041,N_39181);
nand U45107 (N_45107,N_33864,N_39303);
nor U45108 (N_45108,N_38709,N_38743);
nor U45109 (N_45109,N_33685,N_30450);
and U45110 (N_45110,N_39800,N_39441);
nor U45111 (N_45111,N_31843,N_38383);
nand U45112 (N_45112,N_33556,N_33655);
and U45113 (N_45113,N_34873,N_38873);
or U45114 (N_45114,N_38190,N_35610);
xnor U45115 (N_45115,N_36902,N_32038);
nand U45116 (N_45116,N_36903,N_30741);
nand U45117 (N_45117,N_38909,N_32987);
nor U45118 (N_45118,N_30234,N_36546);
nor U45119 (N_45119,N_33906,N_39920);
xor U45120 (N_45120,N_37455,N_33812);
nor U45121 (N_45121,N_32100,N_32646);
nor U45122 (N_45122,N_32361,N_39307);
xor U45123 (N_45123,N_32117,N_36009);
nor U45124 (N_45124,N_38830,N_31110);
xnor U45125 (N_45125,N_37418,N_37279);
or U45126 (N_45126,N_37621,N_33690);
or U45127 (N_45127,N_34432,N_34997);
and U45128 (N_45128,N_30397,N_37337);
and U45129 (N_45129,N_34848,N_37857);
or U45130 (N_45130,N_37952,N_32158);
or U45131 (N_45131,N_39973,N_34525);
nand U45132 (N_45132,N_33113,N_35610);
nor U45133 (N_45133,N_34866,N_38256);
nand U45134 (N_45134,N_34328,N_32542);
and U45135 (N_45135,N_36388,N_37030);
or U45136 (N_45136,N_36336,N_34807);
xnor U45137 (N_45137,N_36662,N_31764);
or U45138 (N_45138,N_34826,N_34808);
nand U45139 (N_45139,N_32266,N_38782);
or U45140 (N_45140,N_31110,N_34039);
and U45141 (N_45141,N_34049,N_34208);
and U45142 (N_45142,N_32500,N_37224);
xnor U45143 (N_45143,N_33993,N_38083);
or U45144 (N_45144,N_39996,N_38727);
and U45145 (N_45145,N_34747,N_32080);
xor U45146 (N_45146,N_37007,N_35876);
xor U45147 (N_45147,N_32619,N_30097);
or U45148 (N_45148,N_36195,N_38831);
nand U45149 (N_45149,N_30747,N_30029);
xnor U45150 (N_45150,N_30423,N_39148);
nor U45151 (N_45151,N_30052,N_35723);
nand U45152 (N_45152,N_37547,N_32519);
nand U45153 (N_45153,N_37231,N_32353);
xnor U45154 (N_45154,N_31608,N_35089);
nand U45155 (N_45155,N_35413,N_32031);
xor U45156 (N_45156,N_37753,N_39710);
or U45157 (N_45157,N_33745,N_35412);
nor U45158 (N_45158,N_37814,N_36584);
nor U45159 (N_45159,N_32148,N_37242);
or U45160 (N_45160,N_35541,N_32561);
and U45161 (N_45161,N_39131,N_38561);
or U45162 (N_45162,N_31428,N_33926);
or U45163 (N_45163,N_37309,N_36421);
and U45164 (N_45164,N_32213,N_37847);
xnor U45165 (N_45165,N_39814,N_36412);
nand U45166 (N_45166,N_32547,N_37985);
nand U45167 (N_45167,N_30715,N_36327);
nand U45168 (N_45168,N_36434,N_39453);
nand U45169 (N_45169,N_30099,N_31016);
or U45170 (N_45170,N_36998,N_33112);
nor U45171 (N_45171,N_31638,N_35082);
xor U45172 (N_45172,N_38781,N_37696);
xnor U45173 (N_45173,N_37497,N_38545);
xnor U45174 (N_45174,N_37685,N_39116);
nand U45175 (N_45175,N_36823,N_31550);
xnor U45176 (N_45176,N_34099,N_31778);
and U45177 (N_45177,N_32184,N_33295);
xor U45178 (N_45178,N_38873,N_37771);
nor U45179 (N_45179,N_37832,N_36343);
nor U45180 (N_45180,N_32441,N_38274);
xnor U45181 (N_45181,N_39991,N_39425);
or U45182 (N_45182,N_37198,N_35017);
xnor U45183 (N_45183,N_39089,N_32591);
or U45184 (N_45184,N_32050,N_32943);
xnor U45185 (N_45185,N_38739,N_35837);
xor U45186 (N_45186,N_38779,N_30472);
nor U45187 (N_45187,N_39580,N_30841);
xor U45188 (N_45188,N_39459,N_38580);
or U45189 (N_45189,N_35814,N_37451);
and U45190 (N_45190,N_31113,N_35715);
nand U45191 (N_45191,N_38504,N_30449);
or U45192 (N_45192,N_35419,N_32790);
nand U45193 (N_45193,N_32237,N_30356);
xor U45194 (N_45194,N_39668,N_33336);
nor U45195 (N_45195,N_33034,N_37664);
xor U45196 (N_45196,N_39262,N_34542);
nand U45197 (N_45197,N_36589,N_35108);
xnor U45198 (N_45198,N_37843,N_33154);
and U45199 (N_45199,N_35082,N_38036);
and U45200 (N_45200,N_39208,N_34539);
nor U45201 (N_45201,N_37132,N_33335);
or U45202 (N_45202,N_34851,N_37305);
nor U45203 (N_45203,N_38857,N_39665);
or U45204 (N_45204,N_38230,N_33148);
and U45205 (N_45205,N_31005,N_33119);
or U45206 (N_45206,N_34934,N_33081);
and U45207 (N_45207,N_36138,N_38574);
nand U45208 (N_45208,N_30917,N_31769);
nand U45209 (N_45209,N_38224,N_39311);
or U45210 (N_45210,N_37711,N_32218);
nand U45211 (N_45211,N_36330,N_37390);
nand U45212 (N_45212,N_37980,N_31761);
or U45213 (N_45213,N_39042,N_31291);
or U45214 (N_45214,N_30793,N_38639);
or U45215 (N_45215,N_37022,N_37010);
and U45216 (N_45216,N_37982,N_35713);
xor U45217 (N_45217,N_37209,N_33139);
nor U45218 (N_45218,N_34151,N_36022);
nor U45219 (N_45219,N_35514,N_38985);
nand U45220 (N_45220,N_36538,N_31475);
or U45221 (N_45221,N_38500,N_37635);
nand U45222 (N_45222,N_34374,N_30382);
nand U45223 (N_45223,N_37852,N_30507);
and U45224 (N_45224,N_32730,N_31117);
nand U45225 (N_45225,N_39921,N_38115);
and U45226 (N_45226,N_37859,N_37596);
nand U45227 (N_45227,N_36807,N_38435);
xor U45228 (N_45228,N_33546,N_31449);
nor U45229 (N_45229,N_38167,N_38632);
and U45230 (N_45230,N_36548,N_30524);
and U45231 (N_45231,N_33813,N_39390);
nand U45232 (N_45232,N_31441,N_38168);
or U45233 (N_45233,N_35545,N_38708);
and U45234 (N_45234,N_35367,N_31144);
xor U45235 (N_45235,N_32147,N_38471);
nand U45236 (N_45236,N_37504,N_30849);
xnor U45237 (N_45237,N_35044,N_37063);
xor U45238 (N_45238,N_37141,N_39156);
xnor U45239 (N_45239,N_37186,N_33687);
or U45240 (N_45240,N_31754,N_33554);
xor U45241 (N_45241,N_34024,N_37905);
xnor U45242 (N_45242,N_35544,N_32011);
and U45243 (N_45243,N_30373,N_39559);
or U45244 (N_45244,N_33896,N_34915);
and U45245 (N_45245,N_35292,N_31259);
nor U45246 (N_45246,N_34889,N_39126);
and U45247 (N_45247,N_38639,N_33273);
and U45248 (N_45248,N_30924,N_35146);
nor U45249 (N_45249,N_36270,N_34349);
nor U45250 (N_45250,N_33184,N_39258);
and U45251 (N_45251,N_37740,N_33834);
nand U45252 (N_45252,N_38317,N_39532);
nand U45253 (N_45253,N_38524,N_38544);
nor U45254 (N_45254,N_34955,N_34229);
xnor U45255 (N_45255,N_36264,N_36680);
or U45256 (N_45256,N_39640,N_34751);
xnor U45257 (N_45257,N_38464,N_37039);
and U45258 (N_45258,N_30390,N_39607);
and U45259 (N_45259,N_30911,N_32032);
and U45260 (N_45260,N_39866,N_34767);
xor U45261 (N_45261,N_31411,N_32628);
nand U45262 (N_45262,N_37604,N_32881);
nor U45263 (N_45263,N_34971,N_37023);
and U45264 (N_45264,N_33709,N_34959);
or U45265 (N_45265,N_33520,N_32201);
nand U45266 (N_45266,N_30198,N_34554);
nor U45267 (N_45267,N_36164,N_32873);
or U45268 (N_45268,N_37616,N_39980);
or U45269 (N_45269,N_31346,N_32748);
and U45270 (N_45270,N_36037,N_38678);
xor U45271 (N_45271,N_39133,N_36210);
and U45272 (N_45272,N_31110,N_34111);
or U45273 (N_45273,N_38471,N_39425);
xnor U45274 (N_45274,N_32045,N_31107);
nor U45275 (N_45275,N_32907,N_35444);
xor U45276 (N_45276,N_33355,N_31272);
or U45277 (N_45277,N_37880,N_35788);
or U45278 (N_45278,N_32936,N_30411);
or U45279 (N_45279,N_30262,N_33341);
or U45280 (N_45280,N_39627,N_34077);
nand U45281 (N_45281,N_32394,N_36898);
nand U45282 (N_45282,N_32476,N_31796);
or U45283 (N_45283,N_36008,N_36141);
nor U45284 (N_45284,N_36393,N_39321);
and U45285 (N_45285,N_39805,N_36806);
nor U45286 (N_45286,N_37438,N_36534);
xnor U45287 (N_45287,N_36687,N_34861);
nand U45288 (N_45288,N_35988,N_34705);
or U45289 (N_45289,N_38310,N_33077);
or U45290 (N_45290,N_30356,N_34636);
or U45291 (N_45291,N_37813,N_37853);
xor U45292 (N_45292,N_30045,N_32674);
and U45293 (N_45293,N_34630,N_38203);
or U45294 (N_45294,N_39523,N_36360);
xnor U45295 (N_45295,N_31198,N_34734);
nor U45296 (N_45296,N_31819,N_31498);
or U45297 (N_45297,N_34167,N_36584);
xor U45298 (N_45298,N_30071,N_37300);
and U45299 (N_45299,N_36084,N_32447);
nand U45300 (N_45300,N_39946,N_38289);
or U45301 (N_45301,N_33754,N_39412);
xor U45302 (N_45302,N_36597,N_33212);
nand U45303 (N_45303,N_33019,N_32993);
nand U45304 (N_45304,N_33161,N_37379);
nand U45305 (N_45305,N_34783,N_38812);
and U45306 (N_45306,N_35621,N_37867);
or U45307 (N_45307,N_39739,N_34963);
and U45308 (N_45308,N_34224,N_39320);
and U45309 (N_45309,N_38778,N_33840);
and U45310 (N_45310,N_39082,N_33465);
nor U45311 (N_45311,N_33830,N_35844);
nand U45312 (N_45312,N_31395,N_36842);
or U45313 (N_45313,N_31703,N_30661);
nand U45314 (N_45314,N_38782,N_36577);
nand U45315 (N_45315,N_30052,N_38818);
xnor U45316 (N_45316,N_37233,N_37653);
and U45317 (N_45317,N_30660,N_31748);
nor U45318 (N_45318,N_37484,N_34910);
xor U45319 (N_45319,N_35115,N_35383);
nor U45320 (N_45320,N_38802,N_32245);
or U45321 (N_45321,N_33498,N_38921);
and U45322 (N_45322,N_37582,N_33708);
and U45323 (N_45323,N_36238,N_33649);
xor U45324 (N_45324,N_39516,N_34001);
nor U45325 (N_45325,N_31530,N_37479);
or U45326 (N_45326,N_36833,N_31336);
nor U45327 (N_45327,N_32646,N_35355);
nand U45328 (N_45328,N_33584,N_30090);
nor U45329 (N_45329,N_39114,N_37306);
nor U45330 (N_45330,N_39161,N_39422);
nand U45331 (N_45331,N_35879,N_36814);
xnor U45332 (N_45332,N_37864,N_32240);
nand U45333 (N_45333,N_34975,N_38123);
and U45334 (N_45334,N_30901,N_30473);
nand U45335 (N_45335,N_33235,N_30659);
and U45336 (N_45336,N_34881,N_38358);
xnor U45337 (N_45337,N_37675,N_36211);
and U45338 (N_45338,N_32181,N_36746);
and U45339 (N_45339,N_35012,N_36784);
or U45340 (N_45340,N_39704,N_30773);
or U45341 (N_45341,N_32238,N_32843);
xor U45342 (N_45342,N_36995,N_31368);
nand U45343 (N_45343,N_35701,N_38232);
nand U45344 (N_45344,N_38640,N_36228);
nor U45345 (N_45345,N_38433,N_39230);
and U45346 (N_45346,N_34522,N_31330);
nor U45347 (N_45347,N_37749,N_32007);
nand U45348 (N_45348,N_30024,N_30915);
or U45349 (N_45349,N_36600,N_33204);
or U45350 (N_45350,N_35385,N_34302);
xnor U45351 (N_45351,N_33435,N_35184);
and U45352 (N_45352,N_32375,N_38394);
and U45353 (N_45353,N_31468,N_36614);
nor U45354 (N_45354,N_37859,N_37443);
xnor U45355 (N_45355,N_35557,N_39366);
or U45356 (N_45356,N_39061,N_38563);
nor U45357 (N_45357,N_36809,N_35202);
or U45358 (N_45358,N_34938,N_37246);
and U45359 (N_45359,N_31787,N_31840);
and U45360 (N_45360,N_35960,N_33193);
nor U45361 (N_45361,N_38919,N_36432);
xor U45362 (N_45362,N_33609,N_32410);
and U45363 (N_45363,N_34139,N_39857);
and U45364 (N_45364,N_38662,N_34234);
or U45365 (N_45365,N_37109,N_39490);
or U45366 (N_45366,N_34709,N_39690);
and U45367 (N_45367,N_33873,N_31814);
xnor U45368 (N_45368,N_31696,N_37903);
nor U45369 (N_45369,N_35472,N_33326);
nor U45370 (N_45370,N_30763,N_30076);
nand U45371 (N_45371,N_38553,N_38917);
nor U45372 (N_45372,N_34464,N_36087);
nand U45373 (N_45373,N_30122,N_39914);
and U45374 (N_45374,N_38386,N_33010);
xor U45375 (N_45375,N_30076,N_36534);
nor U45376 (N_45376,N_39746,N_39736);
nor U45377 (N_45377,N_33118,N_32497);
nand U45378 (N_45378,N_38289,N_38444);
nand U45379 (N_45379,N_33915,N_37929);
or U45380 (N_45380,N_32795,N_33686);
nor U45381 (N_45381,N_38954,N_30694);
nand U45382 (N_45382,N_39092,N_31026);
nand U45383 (N_45383,N_39503,N_34134);
and U45384 (N_45384,N_34281,N_35500);
and U45385 (N_45385,N_38027,N_38619);
or U45386 (N_45386,N_31752,N_30860);
and U45387 (N_45387,N_31140,N_36784);
nor U45388 (N_45388,N_38146,N_32472);
or U45389 (N_45389,N_37200,N_31047);
nor U45390 (N_45390,N_36855,N_34841);
and U45391 (N_45391,N_30950,N_33008);
nor U45392 (N_45392,N_33486,N_38671);
nor U45393 (N_45393,N_32737,N_30458);
and U45394 (N_45394,N_31132,N_38905);
nor U45395 (N_45395,N_39980,N_36307);
xor U45396 (N_45396,N_34620,N_38930);
or U45397 (N_45397,N_36378,N_39329);
and U45398 (N_45398,N_38354,N_37408);
xnor U45399 (N_45399,N_38735,N_34520);
nor U45400 (N_45400,N_30352,N_32287);
nand U45401 (N_45401,N_32933,N_34890);
nand U45402 (N_45402,N_35877,N_31078);
and U45403 (N_45403,N_39833,N_33409);
nand U45404 (N_45404,N_37956,N_34984);
xor U45405 (N_45405,N_30065,N_34097);
nand U45406 (N_45406,N_32130,N_37056);
xor U45407 (N_45407,N_35677,N_34193);
and U45408 (N_45408,N_34357,N_33552);
xor U45409 (N_45409,N_38696,N_32769);
nor U45410 (N_45410,N_31462,N_38190);
nand U45411 (N_45411,N_34494,N_39453);
nor U45412 (N_45412,N_34691,N_35815);
nand U45413 (N_45413,N_37241,N_35859);
or U45414 (N_45414,N_38743,N_37310);
xnor U45415 (N_45415,N_31649,N_34687);
or U45416 (N_45416,N_38442,N_38588);
and U45417 (N_45417,N_38201,N_34894);
xor U45418 (N_45418,N_39369,N_38038);
nand U45419 (N_45419,N_30526,N_36296);
xor U45420 (N_45420,N_31611,N_34700);
nand U45421 (N_45421,N_38435,N_32284);
nand U45422 (N_45422,N_31705,N_31368);
or U45423 (N_45423,N_38123,N_34002);
or U45424 (N_45424,N_39276,N_38264);
nand U45425 (N_45425,N_35174,N_36216);
or U45426 (N_45426,N_39421,N_30896);
nand U45427 (N_45427,N_39540,N_38258);
and U45428 (N_45428,N_35441,N_32570);
nand U45429 (N_45429,N_34709,N_32822);
xnor U45430 (N_45430,N_38280,N_34268);
xnor U45431 (N_45431,N_37120,N_31535);
nor U45432 (N_45432,N_35358,N_30341);
or U45433 (N_45433,N_39580,N_36828);
nor U45434 (N_45434,N_31918,N_37493);
nor U45435 (N_45435,N_38484,N_35035);
nor U45436 (N_45436,N_30412,N_37393);
nor U45437 (N_45437,N_31323,N_31343);
and U45438 (N_45438,N_31705,N_39311);
nand U45439 (N_45439,N_32886,N_33992);
nand U45440 (N_45440,N_36505,N_35679);
nand U45441 (N_45441,N_34731,N_30247);
and U45442 (N_45442,N_31302,N_37892);
nand U45443 (N_45443,N_31876,N_37486);
nand U45444 (N_45444,N_35175,N_38023);
or U45445 (N_45445,N_31175,N_39341);
nor U45446 (N_45446,N_37215,N_35084);
nor U45447 (N_45447,N_39472,N_33051);
or U45448 (N_45448,N_39430,N_33103);
nor U45449 (N_45449,N_39563,N_32614);
nand U45450 (N_45450,N_36234,N_33253);
and U45451 (N_45451,N_32609,N_39795);
xor U45452 (N_45452,N_32093,N_31379);
nor U45453 (N_45453,N_31238,N_32002);
or U45454 (N_45454,N_39037,N_31855);
and U45455 (N_45455,N_39879,N_32875);
nand U45456 (N_45456,N_35895,N_30929);
nand U45457 (N_45457,N_37227,N_37561);
xor U45458 (N_45458,N_30988,N_38089);
and U45459 (N_45459,N_33536,N_35364);
xor U45460 (N_45460,N_39227,N_30871);
and U45461 (N_45461,N_37439,N_38372);
or U45462 (N_45462,N_34364,N_31324);
nor U45463 (N_45463,N_36496,N_37046);
nand U45464 (N_45464,N_34292,N_35264);
nand U45465 (N_45465,N_38171,N_35225);
and U45466 (N_45466,N_37415,N_36966);
or U45467 (N_45467,N_35358,N_34658);
nand U45468 (N_45468,N_30023,N_38235);
nand U45469 (N_45469,N_32920,N_35648);
xor U45470 (N_45470,N_33574,N_37003);
or U45471 (N_45471,N_35593,N_33502);
nor U45472 (N_45472,N_38919,N_33863);
xnor U45473 (N_45473,N_33612,N_38610);
and U45474 (N_45474,N_34136,N_32455);
and U45475 (N_45475,N_33102,N_36235);
nand U45476 (N_45476,N_32997,N_35577);
and U45477 (N_45477,N_38052,N_33831);
nor U45478 (N_45478,N_36527,N_36011);
nor U45479 (N_45479,N_35851,N_39281);
nand U45480 (N_45480,N_39539,N_37575);
nor U45481 (N_45481,N_30133,N_31447);
nor U45482 (N_45482,N_39685,N_33027);
nand U45483 (N_45483,N_34314,N_36982);
nor U45484 (N_45484,N_35445,N_30605);
or U45485 (N_45485,N_31286,N_34434);
or U45486 (N_45486,N_37989,N_39861);
nand U45487 (N_45487,N_39844,N_31125);
or U45488 (N_45488,N_37317,N_39550);
xor U45489 (N_45489,N_37175,N_38361);
xor U45490 (N_45490,N_32806,N_39969);
or U45491 (N_45491,N_39074,N_34660);
xnor U45492 (N_45492,N_37872,N_32283);
and U45493 (N_45493,N_35918,N_30568);
nor U45494 (N_45494,N_33833,N_35670);
nand U45495 (N_45495,N_38533,N_38446);
xor U45496 (N_45496,N_32969,N_32322);
nor U45497 (N_45497,N_38771,N_34332);
nor U45498 (N_45498,N_32200,N_36220);
nand U45499 (N_45499,N_38062,N_30386);
or U45500 (N_45500,N_38264,N_38484);
and U45501 (N_45501,N_39552,N_37387);
and U45502 (N_45502,N_37447,N_35240);
and U45503 (N_45503,N_30862,N_37223);
xor U45504 (N_45504,N_32891,N_37472);
xnor U45505 (N_45505,N_38071,N_30911);
nand U45506 (N_45506,N_31029,N_30987);
xnor U45507 (N_45507,N_34179,N_34723);
and U45508 (N_45508,N_33065,N_31955);
or U45509 (N_45509,N_34579,N_32067);
nor U45510 (N_45510,N_34437,N_33681);
or U45511 (N_45511,N_39261,N_37509);
and U45512 (N_45512,N_36693,N_36613);
and U45513 (N_45513,N_35261,N_33026);
xor U45514 (N_45514,N_39855,N_35091);
nand U45515 (N_45515,N_39366,N_38348);
nor U45516 (N_45516,N_32268,N_36736);
and U45517 (N_45517,N_37845,N_39431);
and U45518 (N_45518,N_32293,N_39417);
nor U45519 (N_45519,N_31236,N_31237);
nand U45520 (N_45520,N_33200,N_34427);
nand U45521 (N_45521,N_34563,N_39928);
or U45522 (N_45522,N_34399,N_36808);
nand U45523 (N_45523,N_36562,N_37811);
and U45524 (N_45524,N_31699,N_37949);
xor U45525 (N_45525,N_33062,N_38543);
nand U45526 (N_45526,N_30730,N_37582);
and U45527 (N_45527,N_39518,N_38079);
nor U45528 (N_45528,N_38158,N_36454);
nand U45529 (N_45529,N_34617,N_31350);
xnor U45530 (N_45530,N_33872,N_36550);
and U45531 (N_45531,N_39375,N_32360);
and U45532 (N_45532,N_38833,N_30258);
and U45533 (N_45533,N_33633,N_34279);
or U45534 (N_45534,N_39282,N_34054);
and U45535 (N_45535,N_37976,N_38885);
or U45536 (N_45536,N_35177,N_31680);
or U45537 (N_45537,N_38407,N_34503);
nor U45538 (N_45538,N_30508,N_31452);
nor U45539 (N_45539,N_36573,N_38683);
nand U45540 (N_45540,N_33258,N_38373);
or U45541 (N_45541,N_37851,N_33695);
nor U45542 (N_45542,N_35308,N_39963);
and U45543 (N_45543,N_36736,N_33374);
and U45544 (N_45544,N_39748,N_39296);
nor U45545 (N_45545,N_38378,N_36017);
or U45546 (N_45546,N_31165,N_32926);
nor U45547 (N_45547,N_37501,N_31124);
nand U45548 (N_45548,N_36794,N_37307);
xor U45549 (N_45549,N_30076,N_32179);
nand U45550 (N_45550,N_37397,N_32950);
and U45551 (N_45551,N_39218,N_34684);
nand U45552 (N_45552,N_31567,N_37224);
and U45553 (N_45553,N_37223,N_39482);
or U45554 (N_45554,N_30397,N_33956);
and U45555 (N_45555,N_36580,N_32627);
nor U45556 (N_45556,N_32473,N_35428);
nand U45557 (N_45557,N_35214,N_30383);
and U45558 (N_45558,N_35840,N_35613);
nor U45559 (N_45559,N_39908,N_30904);
nor U45560 (N_45560,N_32125,N_39080);
nand U45561 (N_45561,N_39656,N_32149);
xnor U45562 (N_45562,N_36091,N_32669);
xnor U45563 (N_45563,N_37002,N_38480);
nand U45564 (N_45564,N_32978,N_32141);
nor U45565 (N_45565,N_38639,N_38543);
nand U45566 (N_45566,N_34540,N_30332);
nand U45567 (N_45567,N_36870,N_31757);
nand U45568 (N_45568,N_37358,N_35634);
xor U45569 (N_45569,N_36296,N_30432);
or U45570 (N_45570,N_36341,N_32432);
nand U45571 (N_45571,N_36838,N_30391);
or U45572 (N_45572,N_38096,N_34887);
and U45573 (N_45573,N_38376,N_35065);
nand U45574 (N_45574,N_39375,N_38901);
and U45575 (N_45575,N_32908,N_31389);
or U45576 (N_45576,N_34787,N_39173);
xor U45577 (N_45577,N_37182,N_32227);
and U45578 (N_45578,N_39047,N_34770);
xor U45579 (N_45579,N_35669,N_33176);
nor U45580 (N_45580,N_31025,N_32099);
nor U45581 (N_45581,N_31848,N_31031);
and U45582 (N_45582,N_36415,N_32745);
nand U45583 (N_45583,N_32757,N_30464);
xnor U45584 (N_45584,N_35135,N_37343);
nand U45585 (N_45585,N_38243,N_30375);
nor U45586 (N_45586,N_33877,N_34720);
or U45587 (N_45587,N_34904,N_38211);
and U45588 (N_45588,N_35519,N_35091);
nor U45589 (N_45589,N_30589,N_34808);
nor U45590 (N_45590,N_34302,N_35115);
xnor U45591 (N_45591,N_35073,N_36234);
nor U45592 (N_45592,N_34765,N_31308);
nand U45593 (N_45593,N_31765,N_36609);
xor U45594 (N_45594,N_30953,N_35336);
or U45595 (N_45595,N_33079,N_33324);
nand U45596 (N_45596,N_32741,N_33300);
or U45597 (N_45597,N_30836,N_31581);
nor U45598 (N_45598,N_33588,N_39942);
nor U45599 (N_45599,N_31119,N_36774);
nor U45600 (N_45600,N_30893,N_36306);
or U45601 (N_45601,N_33069,N_32096);
and U45602 (N_45602,N_32542,N_39993);
or U45603 (N_45603,N_39498,N_37886);
nand U45604 (N_45604,N_34009,N_31008);
or U45605 (N_45605,N_38418,N_31455);
xor U45606 (N_45606,N_33115,N_33656);
and U45607 (N_45607,N_37434,N_30795);
nand U45608 (N_45608,N_35114,N_39370);
xnor U45609 (N_45609,N_34031,N_34820);
xnor U45610 (N_45610,N_38604,N_39059);
nor U45611 (N_45611,N_36538,N_32068);
xor U45612 (N_45612,N_32114,N_31494);
or U45613 (N_45613,N_38336,N_31268);
xor U45614 (N_45614,N_31819,N_36983);
nor U45615 (N_45615,N_32361,N_37567);
or U45616 (N_45616,N_39957,N_33155);
or U45617 (N_45617,N_32705,N_34723);
and U45618 (N_45618,N_37188,N_37356);
and U45619 (N_45619,N_37701,N_33772);
nor U45620 (N_45620,N_37380,N_38991);
xnor U45621 (N_45621,N_37414,N_38430);
xnor U45622 (N_45622,N_37348,N_32119);
or U45623 (N_45623,N_30889,N_37760);
and U45624 (N_45624,N_35707,N_35271);
and U45625 (N_45625,N_35232,N_39136);
and U45626 (N_45626,N_38343,N_34303);
and U45627 (N_45627,N_32344,N_37297);
nor U45628 (N_45628,N_31507,N_33061);
and U45629 (N_45629,N_32174,N_36036);
or U45630 (N_45630,N_35529,N_31752);
nand U45631 (N_45631,N_30599,N_33096);
nor U45632 (N_45632,N_32927,N_33746);
nand U45633 (N_45633,N_39922,N_34318);
nand U45634 (N_45634,N_39662,N_36001);
nor U45635 (N_45635,N_39756,N_37062);
xnor U45636 (N_45636,N_36156,N_36413);
or U45637 (N_45637,N_31859,N_32323);
or U45638 (N_45638,N_37493,N_36375);
or U45639 (N_45639,N_33849,N_30881);
or U45640 (N_45640,N_38496,N_32334);
nand U45641 (N_45641,N_32082,N_39566);
or U45642 (N_45642,N_30614,N_32781);
nor U45643 (N_45643,N_33537,N_30235);
and U45644 (N_45644,N_34315,N_38397);
or U45645 (N_45645,N_39801,N_36553);
or U45646 (N_45646,N_32012,N_34495);
xor U45647 (N_45647,N_39517,N_33706);
nor U45648 (N_45648,N_37638,N_36543);
or U45649 (N_45649,N_33362,N_31512);
nand U45650 (N_45650,N_33932,N_34697);
nand U45651 (N_45651,N_31036,N_35690);
xnor U45652 (N_45652,N_39000,N_38301);
nor U45653 (N_45653,N_31302,N_35047);
and U45654 (N_45654,N_34391,N_34812);
and U45655 (N_45655,N_36433,N_38031);
and U45656 (N_45656,N_37025,N_31315);
xnor U45657 (N_45657,N_32571,N_33824);
nor U45658 (N_45658,N_37126,N_36143);
xnor U45659 (N_45659,N_39620,N_39581);
nor U45660 (N_45660,N_36841,N_35361);
and U45661 (N_45661,N_36197,N_35206);
xor U45662 (N_45662,N_37940,N_34072);
and U45663 (N_45663,N_37580,N_32147);
nand U45664 (N_45664,N_34186,N_37655);
and U45665 (N_45665,N_32354,N_34379);
or U45666 (N_45666,N_31551,N_35571);
or U45667 (N_45667,N_31911,N_31605);
nand U45668 (N_45668,N_30579,N_36956);
nor U45669 (N_45669,N_35195,N_30954);
nand U45670 (N_45670,N_34545,N_30795);
xor U45671 (N_45671,N_36380,N_32633);
nand U45672 (N_45672,N_39009,N_31640);
nor U45673 (N_45673,N_39578,N_39386);
and U45674 (N_45674,N_36970,N_38104);
and U45675 (N_45675,N_35662,N_37074);
or U45676 (N_45676,N_32692,N_36646);
and U45677 (N_45677,N_38855,N_31667);
and U45678 (N_45678,N_33068,N_37739);
xor U45679 (N_45679,N_39869,N_37380);
and U45680 (N_45680,N_37084,N_33255);
nor U45681 (N_45681,N_32617,N_33525);
and U45682 (N_45682,N_36036,N_34322);
nand U45683 (N_45683,N_36562,N_31289);
or U45684 (N_45684,N_33605,N_31218);
xnor U45685 (N_45685,N_39979,N_37182);
and U45686 (N_45686,N_38537,N_36403);
or U45687 (N_45687,N_32231,N_31273);
nand U45688 (N_45688,N_34604,N_32575);
nand U45689 (N_45689,N_30760,N_33092);
xnor U45690 (N_45690,N_36098,N_36372);
nor U45691 (N_45691,N_37949,N_30053);
nand U45692 (N_45692,N_32834,N_34657);
nor U45693 (N_45693,N_39705,N_36878);
or U45694 (N_45694,N_36875,N_34235);
nand U45695 (N_45695,N_37560,N_34363);
nor U45696 (N_45696,N_34396,N_32016);
xnor U45697 (N_45697,N_35367,N_35869);
nand U45698 (N_45698,N_38743,N_32691);
or U45699 (N_45699,N_32407,N_39226);
nor U45700 (N_45700,N_38861,N_34872);
or U45701 (N_45701,N_39815,N_30959);
xnor U45702 (N_45702,N_34314,N_38676);
xnor U45703 (N_45703,N_31964,N_37902);
xor U45704 (N_45704,N_36724,N_38143);
nor U45705 (N_45705,N_36979,N_37474);
or U45706 (N_45706,N_35246,N_31935);
nor U45707 (N_45707,N_39738,N_32201);
nor U45708 (N_45708,N_36193,N_34301);
or U45709 (N_45709,N_39763,N_30148);
xnor U45710 (N_45710,N_32270,N_34784);
nand U45711 (N_45711,N_34762,N_35940);
or U45712 (N_45712,N_32382,N_35371);
or U45713 (N_45713,N_34838,N_36021);
xor U45714 (N_45714,N_30524,N_33143);
nand U45715 (N_45715,N_39968,N_39135);
nor U45716 (N_45716,N_31516,N_35385);
or U45717 (N_45717,N_34198,N_31574);
xor U45718 (N_45718,N_31404,N_34896);
and U45719 (N_45719,N_33672,N_37280);
or U45720 (N_45720,N_30588,N_34458);
or U45721 (N_45721,N_35342,N_36271);
and U45722 (N_45722,N_34170,N_34951);
nor U45723 (N_45723,N_33224,N_32770);
nand U45724 (N_45724,N_38136,N_35135);
nand U45725 (N_45725,N_31803,N_31258);
and U45726 (N_45726,N_38925,N_37447);
nor U45727 (N_45727,N_38887,N_35748);
nand U45728 (N_45728,N_35723,N_34684);
nand U45729 (N_45729,N_31013,N_31071);
nor U45730 (N_45730,N_38729,N_39444);
and U45731 (N_45731,N_35990,N_31234);
nor U45732 (N_45732,N_32316,N_36407);
nor U45733 (N_45733,N_39311,N_34636);
xnor U45734 (N_45734,N_38809,N_38897);
xor U45735 (N_45735,N_30604,N_36584);
xnor U45736 (N_45736,N_30889,N_36658);
xor U45737 (N_45737,N_37022,N_38843);
xnor U45738 (N_45738,N_38978,N_31805);
nor U45739 (N_45739,N_36540,N_31836);
nor U45740 (N_45740,N_32703,N_33558);
or U45741 (N_45741,N_31904,N_38752);
xor U45742 (N_45742,N_39044,N_36206);
nor U45743 (N_45743,N_34988,N_33935);
and U45744 (N_45744,N_36038,N_38163);
nand U45745 (N_45745,N_36747,N_33899);
nand U45746 (N_45746,N_37343,N_37975);
xor U45747 (N_45747,N_33767,N_34299);
nor U45748 (N_45748,N_38602,N_34168);
or U45749 (N_45749,N_39370,N_35352);
and U45750 (N_45750,N_37213,N_34566);
nand U45751 (N_45751,N_30391,N_34012);
or U45752 (N_45752,N_30068,N_35125);
and U45753 (N_45753,N_35691,N_37129);
nor U45754 (N_45754,N_33235,N_39764);
nor U45755 (N_45755,N_37189,N_37670);
xor U45756 (N_45756,N_33182,N_36019);
xor U45757 (N_45757,N_39714,N_33227);
nor U45758 (N_45758,N_31832,N_35226);
or U45759 (N_45759,N_32710,N_37194);
nor U45760 (N_45760,N_33954,N_35499);
xnor U45761 (N_45761,N_34117,N_36894);
or U45762 (N_45762,N_30245,N_30363);
or U45763 (N_45763,N_31524,N_38722);
nor U45764 (N_45764,N_34149,N_32509);
nor U45765 (N_45765,N_31288,N_37911);
nand U45766 (N_45766,N_34982,N_31180);
nor U45767 (N_45767,N_36926,N_33335);
and U45768 (N_45768,N_39345,N_36696);
nor U45769 (N_45769,N_38823,N_31846);
nor U45770 (N_45770,N_34925,N_37746);
xnor U45771 (N_45771,N_35695,N_35802);
xor U45772 (N_45772,N_36060,N_32635);
or U45773 (N_45773,N_33572,N_39701);
nor U45774 (N_45774,N_30802,N_31465);
and U45775 (N_45775,N_34903,N_37366);
or U45776 (N_45776,N_36272,N_38748);
or U45777 (N_45777,N_33662,N_35645);
xnor U45778 (N_45778,N_31718,N_30721);
xor U45779 (N_45779,N_35417,N_38934);
xnor U45780 (N_45780,N_39651,N_36857);
or U45781 (N_45781,N_32672,N_39896);
nand U45782 (N_45782,N_33316,N_35502);
or U45783 (N_45783,N_34169,N_38089);
or U45784 (N_45784,N_37574,N_37522);
and U45785 (N_45785,N_37426,N_37805);
nand U45786 (N_45786,N_36420,N_34017);
and U45787 (N_45787,N_34906,N_39976);
nand U45788 (N_45788,N_39658,N_32954);
or U45789 (N_45789,N_36800,N_32079);
xnor U45790 (N_45790,N_32375,N_36556);
or U45791 (N_45791,N_33747,N_34567);
or U45792 (N_45792,N_39218,N_34481);
nand U45793 (N_45793,N_35888,N_30020);
or U45794 (N_45794,N_32724,N_35605);
nor U45795 (N_45795,N_38067,N_31235);
and U45796 (N_45796,N_31449,N_36900);
nand U45797 (N_45797,N_37513,N_33586);
and U45798 (N_45798,N_33667,N_39800);
nor U45799 (N_45799,N_33013,N_37316);
nor U45800 (N_45800,N_38178,N_39420);
xnor U45801 (N_45801,N_30358,N_37751);
nand U45802 (N_45802,N_32296,N_30240);
nor U45803 (N_45803,N_34818,N_37579);
nand U45804 (N_45804,N_31700,N_32785);
xor U45805 (N_45805,N_36482,N_39171);
nor U45806 (N_45806,N_33589,N_32855);
nand U45807 (N_45807,N_38977,N_32372);
nand U45808 (N_45808,N_39216,N_37655);
nand U45809 (N_45809,N_39771,N_38023);
and U45810 (N_45810,N_35666,N_38599);
nor U45811 (N_45811,N_37651,N_38327);
nor U45812 (N_45812,N_37973,N_31170);
or U45813 (N_45813,N_39632,N_38804);
nor U45814 (N_45814,N_34639,N_38154);
or U45815 (N_45815,N_33269,N_34034);
and U45816 (N_45816,N_30028,N_37530);
nand U45817 (N_45817,N_37822,N_34568);
or U45818 (N_45818,N_34597,N_35426);
nand U45819 (N_45819,N_39456,N_32086);
or U45820 (N_45820,N_34938,N_34295);
nand U45821 (N_45821,N_30145,N_33239);
xor U45822 (N_45822,N_39181,N_34657);
and U45823 (N_45823,N_36210,N_37897);
nand U45824 (N_45824,N_36263,N_30406);
and U45825 (N_45825,N_31939,N_32252);
and U45826 (N_45826,N_37217,N_36709);
nor U45827 (N_45827,N_33881,N_32095);
or U45828 (N_45828,N_31920,N_35694);
and U45829 (N_45829,N_31550,N_35259);
and U45830 (N_45830,N_33401,N_34789);
and U45831 (N_45831,N_32512,N_37974);
and U45832 (N_45832,N_36990,N_32651);
and U45833 (N_45833,N_33764,N_32819);
nand U45834 (N_45834,N_38082,N_38873);
nand U45835 (N_45835,N_32985,N_36964);
nand U45836 (N_45836,N_38862,N_39395);
xor U45837 (N_45837,N_38596,N_30289);
or U45838 (N_45838,N_37004,N_34231);
xor U45839 (N_45839,N_35947,N_39108);
nand U45840 (N_45840,N_36782,N_35489);
xnor U45841 (N_45841,N_38541,N_39987);
nand U45842 (N_45842,N_32438,N_39447);
nand U45843 (N_45843,N_35697,N_31888);
nor U45844 (N_45844,N_31314,N_33494);
nor U45845 (N_45845,N_38816,N_30039);
xor U45846 (N_45846,N_36577,N_33292);
nand U45847 (N_45847,N_31723,N_38592);
and U45848 (N_45848,N_37369,N_31247);
xor U45849 (N_45849,N_34060,N_32739);
nand U45850 (N_45850,N_31777,N_32186);
nor U45851 (N_45851,N_35491,N_33801);
nor U45852 (N_45852,N_33523,N_33959);
nand U45853 (N_45853,N_39201,N_39870);
or U45854 (N_45854,N_31561,N_38782);
nor U45855 (N_45855,N_36512,N_38664);
nor U45856 (N_45856,N_31393,N_34881);
or U45857 (N_45857,N_39481,N_39066);
or U45858 (N_45858,N_39017,N_31819);
and U45859 (N_45859,N_35663,N_31506);
xnor U45860 (N_45860,N_36194,N_36734);
xor U45861 (N_45861,N_35175,N_30717);
xnor U45862 (N_45862,N_31320,N_37342);
nand U45863 (N_45863,N_33887,N_34260);
or U45864 (N_45864,N_39141,N_37903);
nor U45865 (N_45865,N_31634,N_39525);
xnor U45866 (N_45866,N_34010,N_36781);
and U45867 (N_45867,N_35162,N_34159);
nor U45868 (N_45868,N_39008,N_39327);
nor U45869 (N_45869,N_35521,N_31445);
nor U45870 (N_45870,N_36919,N_34678);
or U45871 (N_45871,N_38024,N_35644);
xnor U45872 (N_45872,N_30004,N_31115);
or U45873 (N_45873,N_33562,N_35499);
xor U45874 (N_45874,N_34072,N_35019);
nand U45875 (N_45875,N_39271,N_33873);
xnor U45876 (N_45876,N_36688,N_35404);
or U45877 (N_45877,N_36458,N_30224);
nor U45878 (N_45878,N_39723,N_38922);
or U45879 (N_45879,N_30060,N_32367);
xnor U45880 (N_45880,N_36413,N_30738);
xnor U45881 (N_45881,N_35569,N_34220);
nand U45882 (N_45882,N_37710,N_39161);
or U45883 (N_45883,N_37030,N_34247);
nor U45884 (N_45884,N_30644,N_33829);
or U45885 (N_45885,N_33456,N_30539);
nand U45886 (N_45886,N_31638,N_31919);
or U45887 (N_45887,N_37528,N_30803);
or U45888 (N_45888,N_38707,N_31795);
xnor U45889 (N_45889,N_32910,N_34560);
xor U45890 (N_45890,N_37969,N_32330);
nor U45891 (N_45891,N_38325,N_31737);
and U45892 (N_45892,N_31333,N_33187);
nor U45893 (N_45893,N_35328,N_33714);
or U45894 (N_45894,N_32858,N_34184);
nor U45895 (N_45895,N_31374,N_38824);
or U45896 (N_45896,N_39392,N_34741);
nand U45897 (N_45897,N_35909,N_33269);
xor U45898 (N_45898,N_31023,N_30868);
nand U45899 (N_45899,N_34282,N_36714);
xor U45900 (N_45900,N_39932,N_38635);
nor U45901 (N_45901,N_38154,N_32566);
nor U45902 (N_45902,N_36513,N_36506);
and U45903 (N_45903,N_37757,N_39148);
and U45904 (N_45904,N_38972,N_36213);
xor U45905 (N_45905,N_35232,N_36558);
nor U45906 (N_45906,N_35656,N_30382);
xor U45907 (N_45907,N_34596,N_35687);
nor U45908 (N_45908,N_37329,N_39277);
or U45909 (N_45909,N_35650,N_37073);
or U45910 (N_45910,N_36645,N_39882);
nor U45911 (N_45911,N_39611,N_34860);
or U45912 (N_45912,N_39489,N_35882);
xor U45913 (N_45913,N_38015,N_39398);
and U45914 (N_45914,N_35071,N_31775);
or U45915 (N_45915,N_31229,N_36039);
nand U45916 (N_45916,N_35400,N_38515);
nor U45917 (N_45917,N_38017,N_39045);
xor U45918 (N_45918,N_37137,N_39551);
nand U45919 (N_45919,N_38967,N_37132);
xor U45920 (N_45920,N_37470,N_38175);
nor U45921 (N_45921,N_31758,N_33752);
nand U45922 (N_45922,N_35433,N_37111);
nand U45923 (N_45923,N_37623,N_35654);
nand U45924 (N_45924,N_32864,N_30762);
xor U45925 (N_45925,N_39693,N_36827);
nand U45926 (N_45926,N_32355,N_31260);
nand U45927 (N_45927,N_34678,N_32552);
or U45928 (N_45928,N_39283,N_35081);
nand U45929 (N_45929,N_39407,N_35889);
or U45930 (N_45930,N_33073,N_34088);
nand U45931 (N_45931,N_33498,N_33853);
nand U45932 (N_45932,N_38676,N_39954);
or U45933 (N_45933,N_39799,N_34891);
nand U45934 (N_45934,N_39904,N_31115);
xnor U45935 (N_45935,N_31145,N_39392);
nand U45936 (N_45936,N_38745,N_38085);
and U45937 (N_45937,N_33859,N_36676);
or U45938 (N_45938,N_33400,N_30062);
xnor U45939 (N_45939,N_36682,N_34237);
nor U45940 (N_45940,N_31894,N_37106);
or U45941 (N_45941,N_30225,N_35424);
or U45942 (N_45942,N_36396,N_35259);
nor U45943 (N_45943,N_38394,N_37518);
and U45944 (N_45944,N_30743,N_34740);
nor U45945 (N_45945,N_36805,N_32962);
and U45946 (N_45946,N_32514,N_32618);
or U45947 (N_45947,N_34009,N_33977);
or U45948 (N_45948,N_33964,N_36074);
nor U45949 (N_45949,N_39268,N_36272);
xnor U45950 (N_45950,N_33033,N_33884);
xor U45951 (N_45951,N_32597,N_37601);
nor U45952 (N_45952,N_35129,N_30049);
xnor U45953 (N_45953,N_36328,N_33969);
and U45954 (N_45954,N_34121,N_35834);
or U45955 (N_45955,N_31162,N_37765);
or U45956 (N_45956,N_38822,N_39001);
and U45957 (N_45957,N_36550,N_33405);
xor U45958 (N_45958,N_30217,N_33045);
xor U45959 (N_45959,N_38378,N_38111);
and U45960 (N_45960,N_38585,N_38952);
xnor U45961 (N_45961,N_38967,N_36726);
nor U45962 (N_45962,N_36380,N_35258);
nor U45963 (N_45963,N_30649,N_35960);
xor U45964 (N_45964,N_31230,N_39379);
xor U45965 (N_45965,N_32871,N_33139);
xnor U45966 (N_45966,N_33224,N_37493);
or U45967 (N_45967,N_35785,N_39416);
and U45968 (N_45968,N_37283,N_39579);
nor U45969 (N_45969,N_35074,N_34229);
nor U45970 (N_45970,N_34826,N_33942);
xnor U45971 (N_45971,N_35592,N_32425);
and U45972 (N_45972,N_39449,N_36356);
xor U45973 (N_45973,N_32748,N_37169);
and U45974 (N_45974,N_33336,N_31038);
nor U45975 (N_45975,N_30747,N_37615);
xor U45976 (N_45976,N_30990,N_37606);
or U45977 (N_45977,N_32737,N_30970);
and U45978 (N_45978,N_36687,N_37024);
and U45979 (N_45979,N_31266,N_34950);
and U45980 (N_45980,N_34884,N_35010);
nor U45981 (N_45981,N_35064,N_30048);
nor U45982 (N_45982,N_38163,N_32533);
nand U45983 (N_45983,N_33153,N_38354);
xnor U45984 (N_45984,N_34113,N_34174);
xnor U45985 (N_45985,N_35601,N_38700);
or U45986 (N_45986,N_34141,N_32144);
or U45987 (N_45987,N_33424,N_34737);
nand U45988 (N_45988,N_30090,N_38314);
or U45989 (N_45989,N_31258,N_30608);
and U45990 (N_45990,N_34159,N_32516);
xor U45991 (N_45991,N_38446,N_31567);
nor U45992 (N_45992,N_31298,N_35845);
nand U45993 (N_45993,N_33592,N_39448);
or U45994 (N_45994,N_35324,N_37684);
nor U45995 (N_45995,N_32808,N_37799);
or U45996 (N_45996,N_37412,N_39571);
and U45997 (N_45997,N_32639,N_31664);
nand U45998 (N_45998,N_31892,N_32915);
and U45999 (N_45999,N_39917,N_34337);
or U46000 (N_46000,N_31195,N_38517);
nor U46001 (N_46001,N_33128,N_34466);
or U46002 (N_46002,N_39830,N_38667);
nand U46003 (N_46003,N_34566,N_34967);
and U46004 (N_46004,N_34445,N_30935);
nor U46005 (N_46005,N_35648,N_35253);
nand U46006 (N_46006,N_36314,N_34501);
or U46007 (N_46007,N_33604,N_37026);
xor U46008 (N_46008,N_37988,N_34386);
or U46009 (N_46009,N_30762,N_37848);
nand U46010 (N_46010,N_37349,N_39702);
nand U46011 (N_46011,N_30375,N_39933);
nor U46012 (N_46012,N_31126,N_35349);
nand U46013 (N_46013,N_38590,N_38418);
nand U46014 (N_46014,N_31210,N_32707);
or U46015 (N_46015,N_38753,N_32778);
nor U46016 (N_46016,N_33185,N_35497);
or U46017 (N_46017,N_35385,N_31708);
xor U46018 (N_46018,N_33555,N_39237);
or U46019 (N_46019,N_37482,N_35915);
and U46020 (N_46020,N_34028,N_37669);
nand U46021 (N_46021,N_34023,N_39375);
nand U46022 (N_46022,N_37821,N_32197);
nand U46023 (N_46023,N_37084,N_39099);
and U46024 (N_46024,N_36222,N_39089);
nor U46025 (N_46025,N_39017,N_35029);
or U46026 (N_46026,N_39370,N_37832);
nand U46027 (N_46027,N_30880,N_36873);
xnor U46028 (N_46028,N_39206,N_38481);
or U46029 (N_46029,N_32546,N_38507);
xnor U46030 (N_46030,N_38406,N_30426);
xnor U46031 (N_46031,N_37809,N_33477);
nand U46032 (N_46032,N_31724,N_31069);
nor U46033 (N_46033,N_38006,N_39551);
and U46034 (N_46034,N_37325,N_30561);
nand U46035 (N_46035,N_35742,N_38219);
nor U46036 (N_46036,N_37719,N_37471);
and U46037 (N_46037,N_36923,N_35019);
xor U46038 (N_46038,N_31526,N_33006);
nand U46039 (N_46039,N_35720,N_36365);
or U46040 (N_46040,N_36006,N_37535);
xor U46041 (N_46041,N_38584,N_37299);
or U46042 (N_46042,N_33012,N_36222);
nor U46043 (N_46043,N_39901,N_30569);
xnor U46044 (N_46044,N_38898,N_33537);
or U46045 (N_46045,N_32576,N_33153);
xor U46046 (N_46046,N_34651,N_36239);
nor U46047 (N_46047,N_36734,N_39367);
xnor U46048 (N_46048,N_33243,N_34698);
xor U46049 (N_46049,N_31770,N_31948);
or U46050 (N_46050,N_35629,N_31410);
and U46051 (N_46051,N_32971,N_34979);
nor U46052 (N_46052,N_35500,N_30657);
xor U46053 (N_46053,N_31444,N_38965);
and U46054 (N_46054,N_35214,N_37911);
nor U46055 (N_46055,N_32281,N_34347);
nand U46056 (N_46056,N_39295,N_33590);
nor U46057 (N_46057,N_33901,N_39675);
and U46058 (N_46058,N_34276,N_32792);
xor U46059 (N_46059,N_33545,N_31591);
or U46060 (N_46060,N_35328,N_39181);
xor U46061 (N_46061,N_38269,N_38858);
xnor U46062 (N_46062,N_34299,N_31502);
or U46063 (N_46063,N_30395,N_32610);
or U46064 (N_46064,N_35013,N_39057);
and U46065 (N_46065,N_32710,N_31066);
nand U46066 (N_46066,N_32806,N_38483);
xnor U46067 (N_46067,N_39075,N_32452);
or U46068 (N_46068,N_39023,N_34325);
and U46069 (N_46069,N_31727,N_35026);
and U46070 (N_46070,N_30865,N_31746);
nand U46071 (N_46071,N_38390,N_35240);
nand U46072 (N_46072,N_30527,N_36207);
or U46073 (N_46073,N_30279,N_34092);
nor U46074 (N_46074,N_32899,N_31741);
nor U46075 (N_46075,N_34424,N_34755);
or U46076 (N_46076,N_30175,N_39050);
or U46077 (N_46077,N_33630,N_37134);
nand U46078 (N_46078,N_39062,N_38632);
nand U46079 (N_46079,N_30559,N_36942);
xnor U46080 (N_46080,N_38890,N_34950);
xnor U46081 (N_46081,N_36541,N_31404);
xnor U46082 (N_46082,N_39776,N_36033);
nand U46083 (N_46083,N_39771,N_30985);
nor U46084 (N_46084,N_34609,N_34393);
nor U46085 (N_46085,N_37941,N_35298);
and U46086 (N_46086,N_35505,N_30705);
nor U46087 (N_46087,N_32217,N_36772);
and U46088 (N_46088,N_32929,N_32672);
nor U46089 (N_46089,N_36856,N_31743);
nand U46090 (N_46090,N_37477,N_37951);
or U46091 (N_46091,N_35722,N_35111);
or U46092 (N_46092,N_34354,N_31224);
and U46093 (N_46093,N_32990,N_31551);
and U46094 (N_46094,N_37032,N_33061);
nor U46095 (N_46095,N_34131,N_32901);
xor U46096 (N_46096,N_32251,N_36623);
nor U46097 (N_46097,N_35586,N_33883);
and U46098 (N_46098,N_33284,N_35230);
or U46099 (N_46099,N_37620,N_32594);
nor U46100 (N_46100,N_37715,N_39150);
xor U46101 (N_46101,N_39793,N_39958);
or U46102 (N_46102,N_32695,N_32209);
nor U46103 (N_46103,N_32907,N_30149);
nand U46104 (N_46104,N_38402,N_32509);
xnor U46105 (N_46105,N_32644,N_33193);
nand U46106 (N_46106,N_33068,N_36387);
and U46107 (N_46107,N_32859,N_38292);
or U46108 (N_46108,N_35969,N_39228);
xor U46109 (N_46109,N_30148,N_34933);
nor U46110 (N_46110,N_32752,N_37389);
or U46111 (N_46111,N_33628,N_33550);
nand U46112 (N_46112,N_37036,N_31860);
xor U46113 (N_46113,N_31187,N_39389);
nand U46114 (N_46114,N_35356,N_30710);
or U46115 (N_46115,N_34341,N_30290);
nor U46116 (N_46116,N_35663,N_34249);
or U46117 (N_46117,N_36565,N_37666);
nor U46118 (N_46118,N_32689,N_36599);
and U46119 (N_46119,N_39256,N_39360);
xor U46120 (N_46120,N_33357,N_39547);
or U46121 (N_46121,N_35191,N_31537);
or U46122 (N_46122,N_39284,N_31843);
or U46123 (N_46123,N_38865,N_33216);
xor U46124 (N_46124,N_39392,N_39829);
or U46125 (N_46125,N_31538,N_39677);
or U46126 (N_46126,N_35383,N_35878);
xor U46127 (N_46127,N_30092,N_38109);
or U46128 (N_46128,N_34268,N_33012);
nor U46129 (N_46129,N_36546,N_37457);
nand U46130 (N_46130,N_39177,N_33219);
and U46131 (N_46131,N_39623,N_31959);
nand U46132 (N_46132,N_34161,N_32335);
and U46133 (N_46133,N_33517,N_36574);
xnor U46134 (N_46134,N_31106,N_36015);
xor U46135 (N_46135,N_30186,N_37664);
nor U46136 (N_46136,N_33580,N_33124);
nor U46137 (N_46137,N_31677,N_39696);
xor U46138 (N_46138,N_30466,N_37230);
or U46139 (N_46139,N_37136,N_31034);
and U46140 (N_46140,N_31110,N_33201);
nor U46141 (N_46141,N_35009,N_32111);
xor U46142 (N_46142,N_33233,N_35338);
and U46143 (N_46143,N_30101,N_35924);
nor U46144 (N_46144,N_30067,N_30551);
and U46145 (N_46145,N_34577,N_37834);
or U46146 (N_46146,N_33508,N_38493);
nor U46147 (N_46147,N_33127,N_35545);
or U46148 (N_46148,N_38573,N_31600);
xnor U46149 (N_46149,N_39154,N_33736);
xnor U46150 (N_46150,N_37465,N_37543);
nor U46151 (N_46151,N_36882,N_39557);
or U46152 (N_46152,N_37322,N_37651);
xnor U46153 (N_46153,N_31018,N_36460);
and U46154 (N_46154,N_38392,N_30978);
nor U46155 (N_46155,N_37859,N_39841);
or U46156 (N_46156,N_31872,N_32223);
nor U46157 (N_46157,N_36810,N_36794);
nor U46158 (N_46158,N_30119,N_33818);
or U46159 (N_46159,N_33516,N_37169);
or U46160 (N_46160,N_35609,N_32238);
nor U46161 (N_46161,N_33556,N_33452);
nand U46162 (N_46162,N_37312,N_30147);
xor U46163 (N_46163,N_37480,N_35149);
nor U46164 (N_46164,N_38312,N_31454);
nand U46165 (N_46165,N_34244,N_34783);
nand U46166 (N_46166,N_30124,N_36416);
and U46167 (N_46167,N_36594,N_39244);
nand U46168 (N_46168,N_38500,N_38145);
and U46169 (N_46169,N_34768,N_30271);
and U46170 (N_46170,N_36019,N_32091);
or U46171 (N_46171,N_34014,N_31712);
or U46172 (N_46172,N_39275,N_33576);
xor U46173 (N_46173,N_33055,N_37488);
xor U46174 (N_46174,N_36935,N_36244);
or U46175 (N_46175,N_30401,N_33610);
and U46176 (N_46176,N_34607,N_36104);
nor U46177 (N_46177,N_33001,N_33204);
xnor U46178 (N_46178,N_35247,N_36949);
and U46179 (N_46179,N_38000,N_30530);
or U46180 (N_46180,N_34025,N_39734);
or U46181 (N_46181,N_30379,N_37809);
xnor U46182 (N_46182,N_36521,N_38080);
and U46183 (N_46183,N_31586,N_35471);
and U46184 (N_46184,N_34178,N_36590);
or U46185 (N_46185,N_34799,N_32128);
xnor U46186 (N_46186,N_30323,N_31254);
and U46187 (N_46187,N_39649,N_35431);
nor U46188 (N_46188,N_36968,N_36021);
and U46189 (N_46189,N_38519,N_32249);
xor U46190 (N_46190,N_32125,N_34488);
and U46191 (N_46191,N_32214,N_32313);
xor U46192 (N_46192,N_30108,N_37518);
or U46193 (N_46193,N_34339,N_34351);
or U46194 (N_46194,N_31045,N_39454);
xnor U46195 (N_46195,N_32071,N_34219);
nor U46196 (N_46196,N_38782,N_34839);
nand U46197 (N_46197,N_31072,N_35305);
nor U46198 (N_46198,N_32148,N_35948);
xnor U46199 (N_46199,N_39906,N_38030);
xor U46200 (N_46200,N_35468,N_31512);
nor U46201 (N_46201,N_38926,N_38083);
nand U46202 (N_46202,N_32509,N_35086);
or U46203 (N_46203,N_34916,N_34516);
or U46204 (N_46204,N_34627,N_31733);
and U46205 (N_46205,N_35372,N_32966);
xor U46206 (N_46206,N_36681,N_38481);
or U46207 (N_46207,N_39128,N_39408);
xnor U46208 (N_46208,N_33966,N_32805);
and U46209 (N_46209,N_38787,N_34844);
xnor U46210 (N_46210,N_33553,N_37416);
xor U46211 (N_46211,N_38353,N_38335);
nand U46212 (N_46212,N_39124,N_30770);
xor U46213 (N_46213,N_39670,N_38904);
and U46214 (N_46214,N_33002,N_31835);
nand U46215 (N_46215,N_37846,N_30155);
and U46216 (N_46216,N_37994,N_31938);
and U46217 (N_46217,N_35559,N_35087);
nor U46218 (N_46218,N_35326,N_37629);
xnor U46219 (N_46219,N_35729,N_30406);
xnor U46220 (N_46220,N_35139,N_34286);
nor U46221 (N_46221,N_30740,N_32513);
or U46222 (N_46222,N_38506,N_35730);
nor U46223 (N_46223,N_34989,N_30645);
and U46224 (N_46224,N_37536,N_32025);
nand U46225 (N_46225,N_32502,N_32816);
xnor U46226 (N_46226,N_32839,N_38458);
nand U46227 (N_46227,N_38846,N_35120);
nand U46228 (N_46228,N_37574,N_30282);
nor U46229 (N_46229,N_35833,N_34319);
xor U46230 (N_46230,N_34189,N_32954);
nand U46231 (N_46231,N_30490,N_31432);
nor U46232 (N_46232,N_38921,N_39062);
and U46233 (N_46233,N_34016,N_37390);
nand U46234 (N_46234,N_37562,N_35639);
xnor U46235 (N_46235,N_36832,N_30570);
nand U46236 (N_46236,N_37879,N_32420);
and U46237 (N_46237,N_33577,N_37347);
nor U46238 (N_46238,N_36974,N_37359);
xor U46239 (N_46239,N_32035,N_34854);
or U46240 (N_46240,N_33156,N_34716);
and U46241 (N_46241,N_34157,N_37394);
nor U46242 (N_46242,N_33059,N_32460);
nor U46243 (N_46243,N_32206,N_37840);
nand U46244 (N_46244,N_34103,N_34580);
or U46245 (N_46245,N_35721,N_30079);
or U46246 (N_46246,N_32650,N_34612);
or U46247 (N_46247,N_37337,N_39648);
nand U46248 (N_46248,N_34854,N_36128);
nand U46249 (N_46249,N_30651,N_34927);
nor U46250 (N_46250,N_32863,N_39673);
nand U46251 (N_46251,N_36542,N_31632);
nand U46252 (N_46252,N_33706,N_38856);
and U46253 (N_46253,N_37273,N_34710);
nand U46254 (N_46254,N_35198,N_33016);
nand U46255 (N_46255,N_30984,N_35951);
and U46256 (N_46256,N_37584,N_36289);
or U46257 (N_46257,N_32627,N_39253);
and U46258 (N_46258,N_34219,N_30530);
and U46259 (N_46259,N_38262,N_35642);
nand U46260 (N_46260,N_39113,N_35171);
and U46261 (N_46261,N_37640,N_32080);
xnor U46262 (N_46262,N_31957,N_30275);
nand U46263 (N_46263,N_39952,N_39250);
nand U46264 (N_46264,N_34258,N_37015);
nand U46265 (N_46265,N_32379,N_33575);
or U46266 (N_46266,N_35114,N_33084);
nor U46267 (N_46267,N_36590,N_34375);
and U46268 (N_46268,N_32101,N_31313);
or U46269 (N_46269,N_38740,N_38871);
xnor U46270 (N_46270,N_33222,N_39596);
nand U46271 (N_46271,N_34899,N_34433);
or U46272 (N_46272,N_30671,N_32816);
or U46273 (N_46273,N_31679,N_38078);
xor U46274 (N_46274,N_32972,N_30800);
and U46275 (N_46275,N_34927,N_39595);
nand U46276 (N_46276,N_32536,N_39608);
nand U46277 (N_46277,N_34061,N_30380);
nor U46278 (N_46278,N_39242,N_38235);
and U46279 (N_46279,N_39756,N_36546);
nor U46280 (N_46280,N_35587,N_31475);
nand U46281 (N_46281,N_38714,N_37582);
and U46282 (N_46282,N_34897,N_38544);
nand U46283 (N_46283,N_38100,N_39651);
or U46284 (N_46284,N_33072,N_37943);
and U46285 (N_46285,N_38546,N_30461);
nand U46286 (N_46286,N_35081,N_32875);
xor U46287 (N_46287,N_30234,N_34673);
nor U46288 (N_46288,N_36799,N_30857);
and U46289 (N_46289,N_33876,N_33364);
and U46290 (N_46290,N_34499,N_31593);
and U46291 (N_46291,N_34637,N_36658);
nor U46292 (N_46292,N_39096,N_39645);
or U46293 (N_46293,N_34164,N_38175);
xor U46294 (N_46294,N_37220,N_32061);
xor U46295 (N_46295,N_32549,N_36796);
nand U46296 (N_46296,N_39141,N_30370);
nor U46297 (N_46297,N_34710,N_39582);
or U46298 (N_46298,N_38560,N_33995);
nor U46299 (N_46299,N_35690,N_30445);
nor U46300 (N_46300,N_36030,N_34313);
xor U46301 (N_46301,N_33323,N_33870);
xnor U46302 (N_46302,N_36583,N_37409);
and U46303 (N_46303,N_39487,N_31758);
xor U46304 (N_46304,N_38528,N_34604);
and U46305 (N_46305,N_36749,N_30946);
xnor U46306 (N_46306,N_35276,N_31052);
nor U46307 (N_46307,N_36583,N_32386);
nand U46308 (N_46308,N_33574,N_36416);
and U46309 (N_46309,N_37619,N_31014);
xor U46310 (N_46310,N_38158,N_35542);
and U46311 (N_46311,N_35084,N_35989);
nor U46312 (N_46312,N_35307,N_33970);
or U46313 (N_46313,N_38377,N_39025);
xnor U46314 (N_46314,N_38232,N_31579);
and U46315 (N_46315,N_37532,N_34256);
nor U46316 (N_46316,N_32334,N_35491);
xor U46317 (N_46317,N_31721,N_30555);
and U46318 (N_46318,N_36175,N_32233);
nand U46319 (N_46319,N_36972,N_31246);
or U46320 (N_46320,N_30800,N_32322);
xnor U46321 (N_46321,N_34848,N_38798);
nor U46322 (N_46322,N_35536,N_38570);
nor U46323 (N_46323,N_39744,N_33724);
xnor U46324 (N_46324,N_38829,N_39451);
xnor U46325 (N_46325,N_36673,N_31249);
and U46326 (N_46326,N_32158,N_35282);
or U46327 (N_46327,N_37771,N_33573);
nor U46328 (N_46328,N_36514,N_30056);
xnor U46329 (N_46329,N_32279,N_33560);
nand U46330 (N_46330,N_30786,N_31351);
and U46331 (N_46331,N_37621,N_33472);
or U46332 (N_46332,N_32413,N_31666);
and U46333 (N_46333,N_38277,N_34328);
or U46334 (N_46334,N_38904,N_35231);
nor U46335 (N_46335,N_35684,N_39702);
nor U46336 (N_46336,N_30989,N_38963);
nor U46337 (N_46337,N_37560,N_30234);
nand U46338 (N_46338,N_35897,N_35521);
nor U46339 (N_46339,N_33977,N_38265);
or U46340 (N_46340,N_30662,N_37753);
or U46341 (N_46341,N_37572,N_39814);
and U46342 (N_46342,N_32089,N_32767);
xnor U46343 (N_46343,N_38913,N_33876);
or U46344 (N_46344,N_37670,N_31826);
nor U46345 (N_46345,N_30736,N_32571);
nand U46346 (N_46346,N_36583,N_39493);
nor U46347 (N_46347,N_30823,N_31276);
nor U46348 (N_46348,N_32562,N_33858);
nand U46349 (N_46349,N_33371,N_37703);
nand U46350 (N_46350,N_31905,N_35699);
nor U46351 (N_46351,N_39365,N_37071);
and U46352 (N_46352,N_31823,N_33682);
nor U46353 (N_46353,N_33694,N_33363);
nand U46354 (N_46354,N_31652,N_38334);
nand U46355 (N_46355,N_33977,N_38716);
xnor U46356 (N_46356,N_34821,N_30364);
nand U46357 (N_46357,N_39394,N_31486);
nor U46358 (N_46358,N_31549,N_33971);
and U46359 (N_46359,N_35292,N_33279);
xor U46360 (N_46360,N_34904,N_31267);
nor U46361 (N_46361,N_38042,N_30867);
nand U46362 (N_46362,N_33227,N_35985);
nor U46363 (N_46363,N_30000,N_33095);
xor U46364 (N_46364,N_30309,N_30994);
nor U46365 (N_46365,N_30265,N_35993);
and U46366 (N_46366,N_30805,N_38246);
or U46367 (N_46367,N_31320,N_38325);
or U46368 (N_46368,N_38064,N_33648);
and U46369 (N_46369,N_32577,N_37094);
nand U46370 (N_46370,N_33873,N_39599);
nand U46371 (N_46371,N_37244,N_35969);
nor U46372 (N_46372,N_34782,N_31069);
nand U46373 (N_46373,N_37962,N_38982);
nor U46374 (N_46374,N_38254,N_33634);
xnor U46375 (N_46375,N_31486,N_32733);
or U46376 (N_46376,N_38535,N_34495);
xor U46377 (N_46377,N_38955,N_38039);
xor U46378 (N_46378,N_31551,N_30496);
and U46379 (N_46379,N_32061,N_32302);
xnor U46380 (N_46380,N_38978,N_30803);
xor U46381 (N_46381,N_34174,N_35842);
xnor U46382 (N_46382,N_39867,N_39501);
nand U46383 (N_46383,N_36327,N_30459);
and U46384 (N_46384,N_30786,N_30799);
xnor U46385 (N_46385,N_31064,N_39388);
nor U46386 (N_46386,N_31901,N_30226);
or U46387 (N_46387,N_33656,N_39299);
and U46388 (N_46388,N_35182,N_33679);
xnor U46389 (N_46389,N_33910,N_31940);
or U46390 (N_46390,N_38038,N_31778);
and U46391 (N_46391,N_31878,N_36893);
nand U46392 (N_46392,N_30040,N_37692);
and U46393 (N_46393,N_39330,N_34556);
or U46394 (N_46394,N_35975,N_31287);
or U46395 (N_46395,N_30377,N_37051);
nand U46396 (N_46396,N_36109,N_31131);
xnor U46397 (N_46397,N_35178,N_37024);
or U46398 (N_46398,N_32111,N_34797);
xnor U46399 (N_46399,N_35824,N_38482);
nor U46400 (N_46400,N_31164,N_31836);
nor U46401 (N_46401,N_36826,N_37611);
xnor U46402 (N_46402,N_38871,N_37340);
and U46403 (N_46403,N_37795,N_37228);
and U46404 (N_46404,N_37828,N_37626);
nor U46405 (N_46405,N_35756,N_35440);
nor U46406 (N_46406,N_34193,N_38211);
and U46407 (N_46407,N_31490,N_32836);
nand U46408 (N_46408,N_36473,N_37734);
nor U46409 (N_46409,N_37600,N_33300);
or U46410 (N_46410,N_32506,N_32250);
nor U46411 (N_46411,N_35963,N_38014);
nor U46412 (N_46412,N_37739,N_33066);
nand U46413 (N_46413,N_37244,N_37148);
and U46414 (N_46414,N_35822,N_36967);
xor U46415 (N_46415,N_33865,N_39712);
xor U46416 (N_46416,N_33485,N_33241);
or U46417 (N_46417,N_34772,N_37700);
xnor U46418 (N_46418,N_33669,N_36916);
nor U46419 (N_46419,N_36117,N_35498);
nand U46420 (N_46420,N_31991,N_31202);
or U46421 (N_46421,N_36415,N_39141);
and U46422 (N_46422,N_31463,N_33369);
or U46423 (N_46423,N_36628,N_36243);
and U46424 (N_46424,N_33066,N_36240);
nand U46425 (N_46425,N_31157,N_33362);
and U46426 (N_46426,N_30491,N_30929);
and U46427 (N_46427,N_35364,N_38788);
xor U46428 (N_46428,N_31265,N_39857);
or U46429 (N_46429,N_36471,N_31153);
or U46430 (N_46430,N_31075,N_30825);
nand U46431 (N_46431,N_30632,N_35762);
nor U46432 (N_46432,N_33505,N_34889);
nor U46433 (N_46433,N_37444,N_35075);
xnor U46434 (N_46434,N_38293,N_35369);
nand U46435 (N_46435,N_33000,N_31666);
nor U46436 (N_46436,N_38863,N_30252);
xnor U46437 (N_46437,N_39723,N_30556);
nor U46438 (N_46438,N_38579,N_35540);
and U46439 (N_46439,N_32836,N_30399);
nor U46440 (N_46440,N_37285,N_31747);
xnor U46441 (N_46441,N_36547,N_33865);
nand U46442 (N_46442,N_35183,N_38298);
xnor U46443 (N_46443,N_38684,N_33953);
nand U46444 (N_46444,N_30457,N_31850);
xor U46445 (N_46445,N_38232,N_32113);
nand U46446 (N_46446,N_36147,N_30309);
nor U46447 (N_46447,N_30620,N_32961);
or U46448 (N_46448,N_35360,N_37548);
xnor U46449 (N_46449,N_35201,N_36554);
and U46450 (N_46450,N_35618,N_39912);
xor U46451 (N_46451,N_34270,N_35319);
xor U46452 (N_46452,N_32464,N_36089);
xnor U46453 (N_46453,N_32096,N_35998);
nand U46454 (N_46454,N_39785,N_39511);
xnor U46455 (N_46455,N_32017,N_37403);
or U46456 (N_46456,N_37000,N_33488);
xnor U46457 (N_46457,N_39278,N_37034);
nand U46458 (N_46458,N_30731,N_38286);
and U46459 (N_46459,N_37127,N_34662);
or U46460 (N_46460,N_33842,N_38494);
or U46461 (N_46461,N_37848,N_37081);
xnor U46462 (N_46462,N_33815,N_33473);
or U46463 (N_46463,N_31586,N_30726);
nand U46464 (N_46464,N_35856,N_31676);
nor U46465 (N_46465,N_30607,N_34223);
nor U46466 (N_46466,N_33152,N_37036);
nand U46467 (N_46467,N_34187,N_31822);
nand U46468 (N_46468,N_30389,N_37337);
xor U46469 (N_46469,N_33306,N_31075);
nand U46470 (N_46470,N_34407,N_35025);
nand U46471 (N_46471,N_32094,N_32638);
and U46472 (N_46472,N_37722,N_33653);
and U46473 (N_46473,N_34923,N_36246);
xor U46474 (N_46474,N_36149,N_37759);
or U46475 (N_46475,N_32309,N_33557);
xnor U46476 (N_46476,N_34003,N_38009);
xor U46477 (N_46477,N_33348,N_30879);
xor U46478 (N_46478,N_37281,N_34288);
nor U46479 (N_46479,N_35541,N_31385);
or U46480 (N_46480,N_31454,N_31736);
and U46481 (N_46481,N_30739,N_30068);
xnor U46482 (N_46482,N_35380,N_34375);
nor U46483 (N_46483,N_37298,N_31207);
and U46484 (N_46484,N_32981,N_35899);
and U46485 (N_46485,N_32785,N_38510);
xor U46486 (N_46486,N_38903,N_31141);
and U46487 (N_46487,N_34671,N_39576);
or U46488 (N_46488,N_32496,N_38485);
and U46489 (N_46489,N_38757,N_33087);
or U46490 (N_46490,N_37458,N_35195);
and U46491 (N_46491,N_38992,N_38145);
or U46492 (N_46492,N_33797,N_34690);
and U46493 (N_46493,N_33080,N_30453);
and U46494 (N_46494,N_32050,N_39378);
nand U46495 (N_46495,N_37923,N_38391);
and U46496 (N_46496,N_36039,N_38291);
or U46497 (N_46497,N_39546,N_31249);
and U46498 (N_46498,N_39572,N_31556);
or U46499 (N_46499,N_31923,N_38809);
xnor U46500 (N_46500,N_34202,N_38858);
or U46501 (N_46501,N_35091,N_35504);
nor U46502 (N_46502,N_32175,N_34700);
and U46503 (N_46503,N_30048,N_39199);
and U46504 (N_46504,N_32462,N_30094);
nand U46505 (N_46505,N_36358,N_30114);
xnor U46506 (N_46506,N_37155,N_38933);
and U46507 (N_46507,N_34336,N_34230);
nor U46508 (N_46508,N_32725,N_38308);
and U46509 (N_46509,N_30112,N_39295);
nor U46510 (N_46510,N_35569,N_32140);
and U46511 (N_46511,N_34951,N_32488);
nand U46512 (N_46512,N_39074,N_35117);
xor U46513 (N_46513,N_31907,N_35584);
nor U46514 (N_46514,N_35253,N_38647);
nor U46515 (N_46515,N_31306,N_32443);
and U46516 (N_46516,N_31150,N_32326);
nand U46517 (N_46517,N_34166,N_33720);
nor U46518 (N_46518,N_33482,N_38742);
nor U46519 (N_46519,N_34339,N_30042);
nand U46520 (N_46520,N_30323,N_38759);
nor U46521 (N_46521,N_36490,N_38459);
nand U46522 (N_46522,N_37572,N_32387);
nand U46523 (N_46523,N_31183,N_35591);
or U46524 (N_46524,N_38709,N_39668);
xor U46525 (N_46525,N_38400,N_31046);
xnor U46526 (N_46526,N_31920,N_30871);
nand U46527 (N_46527,N_37218,N_33169);
or U46528 (N_46528,N_32372,N_31783);
nand U46529 (N_46529,N_33481,N_32614);
and U46530 (N_46530,N_30513,N_35101);
or U46531 (N_46531,N_32769,N_30280);
xor U46532 (N_46532,N_33089,N_34321);
or U46533 (N_46533,N_37349,N_34056);
nand U46534 (N_46534,N_35996,N_35747);
and U46535 (N_46535,N_31017,N_37363);
nor U46536 (N_46536,N_39584,N_35255);
nand U46537 (N_46537,N_32773,N_33616);
and U46538 (N_46538,N_31260,N_30351);
nand U46539 (N_46539,N_38366,N_33026);
and U46540 (N_46540,N_38287,N_39339);
or U46541 (N_46541,N_32380,N_30886);
nor U46542 (N_46542,N_39851,N_39773);
nor U46543 (N_46543,N_32454,N_39105);
nor U46544 (N_46544,N_32081,N_31189);
or U46545 (N_46545,N_30405,N_34949);
nand U46546 (N_46546,N_38212,N_33133);
and U46547 (N_46547,N_39193,N_39355);
xor U46548 (N_46548,N_37014,N_32674);
xor U46549 (N_46549,N_30580,N_35286);
or U46550 (N_46550,N_33124,N_31826);
nand U46551 (N_46551,N_39811,N_39219);
and U46552 (N_46552,N_39332,N_39133);
xor U46553 (N_46553,N_38954,N_33081);
and U46554 (N_46554,N_34956,N_36770);
xor U46555 (N_46555,N_30958,N_38642);
or U46556 (N_46556,N_35468,N_31625);
and U46557 (N_46557,N_34175,N_39949);
or U46558 (N_46558,N_31805,N_38727);
nor U46559 (N_46559,N_30918,N_34354);
nand U46560 (N_46560,N_30651,N_34772);
nor U46561 (N_46561,N_31354,N_32895);
or U46562 (N_46562,N_38661,N_31547);
and U46563 (N_46563,N_33599,N_33534);
or U46564 (N_46564,N_34764,N_30959);
xor U46565 (N_46565,N_36958,N_32749);
xor U46566 (N_46566,N_35391,N_38405);
nand U46567 (N_46567,N_33147,N_39209);
nor U46568 (N_46568,N_37284,N_38359);
xor U46569 (N_46569,N_38021,N_38214);
nor U46570 (N_46570,N_39321,N_39742);
and U46571 (N_46571,N_33969,N_37129);
or U46572 (N_46572,N_38983,N_30888);
xor U46573 (N_46573,N_34989,N_34400);
nor U46574 (N_46574,N_38094,N_37844);
or U46575 (N_46575,N_32243,N_39941);
or U46576 (N_46576,N_34882,N_32412);
or U46577 (N_46577,N_31861,N_32116);
xor U46578 (N_46578,N_36346,N_37255);
or U46579 (N_46579,N_33646,N_37690);
nor U46580 (N_46580,N_34333,N_36083);
nand U46581 (N_46581,N_37430,N_30345);
nand U46582 (N_46582,N_32045,N_30387);
or U46583 (N_46583,N_30098,N_31016);
and U46584 (N_46584,N_31959,N_36535);
xnor U46585 (N_46585,N_34629,N_34370);
and U46586 (N_46586,N_36462,N_33853);
and U46587 (N_46587,N_37499,N_33559);
nor U46588 (N_46588,N_32634,N_39571);
or U46589 (N_46589,N_31250,N_33088);
and U46590 (N_46590,N_38364,N_37459);
nand U46591 (N_46591,N_31027,N_36142);
xnor U46592 (N_46592,N_33410,N_36496);
xnor U46593 (N_46593,N_35257,N_38867);
or U46594 (N_46594,N_36708,N_33751);
xor U46595 (N_46595,N_34393,N_35255);
nor U46596 (N_46596,N_39645,N_34877);
nand U46597 (N_46597,N_38217,N_30946);
xnor U46598 (N_46598,N_31687,N_38887);
nor U46599 (N_46599,N_38019,N_35363);
nor U46600 (N_46600,N_32947,N_31244);
nor U46601 (N_46601,N_31141,N_31467);
or U46602 (N_46602,N_38972,N_36280);
nor U46603 (N_46603,N_33403,N_33919);
and U46604 (N_46604,N_34520,N_37868);
or U46605 (N_46605,N_38489,N_32149);
xnor U46606 (N_46606,N_37595,N_35029);
nor U46607 (N_46607,N_37625,N_39405);
nand U46608 (N_46608,N_33722,N_34496);
or U46609 (N_46609,N_34581,N_30864);
nand U46610 (N_46610,N_38875,N_30176);
or U46611 (N_46611,N_34577,N_38322);
and U46612 (N_46612,N_34203,N_30901);
nand U46613 (N_46613,N_31991,N_38259);
xor U46614 (N_46614,N_36989,N_34255);
xnor U46615 (N_46615,N_30786,N_38621);
xor U46616 (N_46616,N_34709,N_33418);
and U46617 (N_46617,N_31434,N_31637);
nand U46618 (N_46618,N_38833,N_32456);
xnor U46619 (N_46619,N_35474,N_39943);
and U46620 (N_46620,N_35413,N_38823);
or U46621 (N_46621,N_34194,N_39158);
or U46622 (N_46622,N_39548,N_34794);
nor U46623 (N_46623,N_35654,N_39069);
nand U46624 (N_46624,N_34417,N_33629);
or U46625 (N_46625,N_39352,N_31293);
or U46626 (N_46626,N_37897,N_33231);
or U46627 (N_46627,N_37073,N_32894);
nor U46628 (N_46628,N_35477,N_35532);
and U46629 (N_46629,N_30812,N_38103);
nand U46630 (N_46630,N_38722,N_32680);
and U46631 (N_46631,N_30044,N_39564);
nand U46632 (N_46632,N_32758,N_38782);
and U46633 (N_46633,N_35861,N_34504);
xnor U46634 (N_46634,N_30012,N_35788);
nor U46635 (N_46635,N_30161,N_30064);
and U46636 (N_46636,N_38026,N_35626);
nand U46637 (N_46637,N_35391,N_34462);
xor U46638 (N_46638,N_32604,N_34916);
xnor U46639 (N_46639,N_31293,N_39814);
nor U46640 (N_46640,N_32450,N_31620);
and U46641 (N_46641,N_30840,N_33650);
xnor U46642 (N_46642,N_35354,N_38396);
and U46643 (N_46643,N_38694,N_36171);
xor U46644 (N_46644,N_33833,N_34910);
nand U46645 (N_46645,N_39834,N_37466);
nand U46646 (N_46646,N_38640,N_39712);
nand U46647 (N_46647,N_33180,N_37729);
xor U46648 (N_46648,N_39451,N_38308);
or U46649 (N_46649,N_30735,N_38614);
or U46650 (N_46650,N_31179,N_32684);
nand U46651 (N_46651,N_36238,N_37130);
and U46652 (N_46652,N_39596,N_30628);
nor U46653 (N_46653,N_33950,N_34795);
nand U46654 (N_46654,N_30074,N_32975);
or U46655 (N_46655,N_39867,N_34385);
nand U46656 (N_46656,N_33624,N_32760);
and U46657 (N_46657,N_32259,N_31462);
xnor U46658 (N_46658,N_35661,N_32334);
nor U46659 (N_46659,N_32567,N_39421);
xor U46660 (N_46660,N_34164,N_30960);
or U46661 (N_46661,N_30070,N_36391);
xnor U46662 (N_46662,N_36323,N_31872);
or U46663 (N_46663,N_38728,N_37946);
nor U46664 (N_46664,N_34586,N_32994);
xnor U46665 (N_46665,N_35740,N_37499);
xnor U46666 (N_46666,N_39617,N_31485);
nand U46667 (N_46667,N_34456,N_31015);
and U46668 (N_46668,N_39780,N_37817);
nand U46669 (N_46669,N_33778,N_35224);
and U46670 (N_46670,N_30886,N_36352);
and U46671 (N_46671,N_39188,N_33807);
xor U46672 (N_46672,N_34453,N_32370);
and U46673 (N_46673,N_38146,N_32259);
nor U46674 (N_46674,N_37148,N_32282);
nor U46675 (N_46675,N_38465,N_33971);
xor U46676 (N_46676,N_39152,N_31903);
xnor U46677 (N_46677,N_32168,N_32839);
nand U46678 (N_46678,N_39652,N_31263);
nor U46679 (N_46679,N_30918,N_35838);
nand U46680 (N_46680,N_36020,N_39689);
and U46681 (N_46681,N_34881,N_36374);
and U46682 (N_46682,N_30621,N_38948);
nor U46683 (N_46683,N_34595,N_36200);
nor U46684 (N_46684,N_39786,N_39810);
nand U46685 (N_46685,N_38929,N_37151);
nor U46686 (N_46686,N_31555,N_39436);
nor U46687 (N_46687,N_39924,N_35845);
or U46688 (N_46688,N_35706,N_38970);
or U46689 (N_46689,N_30238,N_33290);
nand U46690 (N_46690,N_31439,N_33852);
nor U46691 (N_46691,N_34806,N_35875);
xor U46692 (N_46692,N_37390,N_35882);
nor U46693 (N_46693,N_36969,N_30399);
nor U46694 (N_46694,N_34971,N_36936);
xor U46695 (N_46695,N_33424,N_38303);
xnor U46696 (N_46696,N_36069,N_39725);
nand U46697 (N_46697,N_39343,N_32452);
nand U46698 (N_46698,N_39872,N_30975);
nor U46699 (N_46699,N_38306,N_30392);
or U46700 (N_46700,N_34749,N_30726);
and U46701 (N_46701,N_36338,N_39036);
and U46702 (N_46702,N_37858,N_36222);
and U46703 (N_46703,N_34869,N_33148);
nor U46704 (N_46704,N_32505,N_36742);
nor U46705 (N_46705,N_34673,N_34709);
nor U46706 (N_46706,N_32752,N_36547);
or U46707 (N_46707,N_36894,N_35320);
and U46708 (N_46708,N_33257,N_31618);
xor U46709 (N_46709,N_39996,N_38821);
nand U46710 (N_46710,N_39326,N_31694);
nand U46711 (N_46711,N_30303,N_38674);
nand U46712 (N_46712,N_32078,N_38223);
nor U46713 (N_46713,N_30124,N_39452);
and U46714 (N_46714,N_30002,N_33921);
xor U46715 (N_46715,N_34243,N_33147);
xnor U46716 (N_46716,N_36491,N_38036);
or U46717 (N_46717,N_37418,N_39896);
nand U46718 (N_46718,N_34959,N_30606);
nand U46719 (N_46719,N_32686,N_33543);
nand U46720 (N_46720,N_30083,N_33884);
nand U46721 (N_46721,N_31509,N_33545);
nand U46722 (N_46722,N_37183,N_38414);
xnor U46723 (N_46723,N_39600,N_35261);
or U46724 (N_46724,N_30961,N_33566);
nand U46725 (N_46725,N_35431,N_31780);
nand U46726 (N_46726,N_35502,N_39178);
nand U46727 (N_46727,N_36554,N_32109);
nor U46728 (N_46728,N_32434,N_39260);
xnor U46729 (N_46729,N_38637,N_38348);
or U46730 (N_46730,N_34786,N_35372);
and U46731 (N_46731,N_35144,N_39038);
or U46732 (N_46732,N_36090,N_39634);
or U46733 (N_46733,N_35933,N_31783);
xnor U46734 (N_46734,N_39975,N_36958);
nor U46735 (N_46735,N_33719,N_32734);
or U46736 (N_46736,N_34039,N_33209);
xnor U46737 (N_46737,N_38756,N_39775);
and U46738 (N_46738,N_32524,N_34442);
or U46739 (N_46739,N_39029,N_33859);
and U46740 (N_46740,N_38307,N_30999);
nand U46741 (N_46741,N_34279,N_39518);
or U46742 (N_46742,N_36217,N_36553);
xnor U46743 (N_46743,N_38154,N_37563);
or U46744 (N_46744,N_36287,N_37089);
nand U46745 (N_46745,N_37907,N_38560);
xnor U46746 (N_46746,N_38817,N_30965);
nor U46747 (N_46747,N_36225,N_37341);
nor U46748 (N_46748,N_34403,N_37858);
and U46749 (N_46749,N_33045,N_38558);
or U46750 (N_46750,N_35225,N_33753);
xnor U46751 (N_46751,N_35209,N_34893);
nor U46752 (N_46752,N_35077,N_34910);
nor U46753 (N_46753,N_33724,N_34614);
or U46754 (N_46754,N_36270,N_33376);
nand U46755 (N_46755,N_33522,N_31412);
nor U46756 (N_46756,N_31305,N_31223);
and U46757 (N_46757,N_35737,N_37779);
nand U46758 (N_46758,N_35171,N_35735);
nor U46759 (N_46759,N_32438,N_30635);
xor U46760 (N_46760,N_39431,N_32164);
or U46761 (N_46761,N_34827,N_39573);
nand U46762 (N_46762,N_38999,N_39158);
xor U46763 (N_46763,N_32418,N_31932);
xnor U46764 (N_46764,N_38925,N_37359);
nand U46765 (N_46765,N_31977,N_39863);
or U46766 (N_46766,N_32375,N_35768);
nand U46767 (N_46767,N_34926,N_31884);
nor U46768 (N_46768,N_35863,N_35864);
or U46769 (N_46769,N_39462,N_38422);
or U46770 (N_46770,N_33764,N_38129);
nor U46771 (N_46771,N_32459,N_37489);
or U46772 (N_46772,N_32383,N_31297);
and U46773 (N_46773,N_33622,N_34732);
nor U46774 (N_46774,N_39735,N_37953);
xnor U46775 (N_46775,N_33253,N_32471);
nand U46776 (N_46776,N_39630,N_30356);
or U46777 (N_46777,N_39295,N_36571);
nor U46778 (N_46778,N_34586,N_35904);
nor U46779 (N_46779,N_38038,N_36207);
or U46780 (N_46780,N_32466,N_31526);
and U46781 (N_46781,N_30515,N_36114);
xor U46782 (N_46782,N_38520,N_37401);
and U46783 (N_46783,N_31782,N_39846);
or U46784 (N_46784,N_33353,N_38555);
and U46785 (N_46785,N_32310,N_34296);
or U46786 (N_46786,N_31218,N_34121);
nor U46787 (N_46787,N_33750,N_30309);
and U46788 (N_46788,N_31558,N_30928);
or U46789 (N_46789,N_34202,N_39696);
or U46790 (N_46790,N_38243,N_33508);
xnor U46791 (N_46791,N_36587,N_33031);
or U46792 (N_46792,N_39310,N_37371);
nor U46793 (N_46793,N_33285,N_34310);
nor U46794 (N_46794,N_33214,N_39007);
nand U46795 (N_46795,N_39708,N_30793);
or U46796 (N_46796,N_32065,N_35303);
and U46797 (N_46797,N_33636,N_31270);
xnor U46798 (N_46798,N_33239,N_39560);
xor U46799 (N_46799,N_39367,N_37783);
or U46800 (N_46800,N_30844,N_33177);
and U46801 (N_46801,N_34448,N_30762);
nand U46802 (N_46802,N_34395,N_39914);
and U46803 (N_46803,N_34450,N_38896);
xor U46804 (N_46804,N_30228,N_35071);
xor U46805 (N_46805,N_36600,N_39785);
nor U46806 (N_46806,N_38302,N_30216);
nand U46807 (N_46807,N_32706,N_39843);
xor U46808 (N_46808,N_35539,N_33546);
nor U46809 (N_46809,N_30892,N_30417);
or U46810 (N_46810,N_37920,N_36267);
and U46811 (N_46811,N_33026,N_33983);
or U46812 (N_46812,N_35421,N_37259);
and U46813 (N_46813,N_35962,N_38019);
or U46814 (N_46814,N_32888,N_33218);
or U46815 (N_46815,N_38440,N_38118);
nand U46816 (N_46816,N_37451,N_37226);
and U46817 (N_46817,N_33284,N_39617);
or U46818 (N_46818,N_38033,N_39878);
nand U46819 (N_46819,N_32605,N_37910);
or U46820 (N_46820,N_37073,N_36572);
nor U46821 (N_46821,N_36744,N_37239);
xnor U46822 (N_46822,N_31712,N_36072);
nor U46823 (N_46823,N_36910,N_34936);
nand U46824 (N_46824,N_35212,N_37931);
or U46825 (N_46825,N_31103,N_33400);
xor U46826 (N_46826,N_31174,N_38413);
and U46827 (N_46827,N_38444,N_31932);
or U46828 (N_46828,N_37577,N_39710);
or U46829 (N_46829,N_35228,N_35923);
and U46830 (N_46830,N_33857,N_37455);
xnor U46831 (N_46831,N_32201,N_31068);
nand U46832 (N_46832,N_39105,N_32305);
nor U46833 (N_46833,N_37672,N_39076);
and U46834 (N_46834,N_38771,N_39198);
xnor U46835 (N_46835,N_39360,N_36073);
xnor U46836 (N_46836,N_31996,N_33917);
xnor U46837 (N_46837,N_32177,N_39452);
nand U46838 (N_46838,N_34160,N_32815);
nor U46839 (N_46839,N_35975,N_34762);
nor U46840 (N_46840,N_31888,N_34592);
xnor U46841 (N_46841,N_33207,N_33597);
xnor U46842 (N_46842,N_35832,N_36766);
or U46843 (N_46843,N_34966,N_30912);
nand U46844 (N_46844,N_33843,N_35773);
or U46845 (N_46845,N_31082,N_31134);
nand U46846 (N_46846,N_31875,N_36977);
and U46847 (N_46847,N_39411,N_36625);
nand U46848 (N_46848,N_37676,N_37764);
or U46849 (N_46849,N_35726,N_34558);
nand U46850 (N_46850,N_31520,N_32590);
and U46851 (N_46851,N_37286,N_30224);
and U46852 (N_46852,N_32062,N_35779);
nand U46853 (N_46853,N_32253,N_34150);
nand U46854 (N_46854,N_32271,N_32951);
nand U46855 (N_46855,N_38830,N_36329);
nand U46856 (N_46856,N_31098,N_39390);
or U46857 (N_46857,N_35041,N_38703);
xnor U46858 (N_46858,N_30425,N_39635);
and U46859 (N_46859,N_39054,N_30315);
nand U46860 (N_46860,N_36850,N_38386);
and U46861 (N_46861,N_35798,N_37532);
nor U46862 (N_46862,N_38801,N_34520);
nand U46863 (N_46863,N_31095,N_33817);
nand U46864 (N_46864,N_30316,N_33911);
nand U46865 (N_46865,N_36516,N_33135);
nor U46866 (N_46866,N_33759,N_35598);
nor U46867 (N_46867,N_36669,N_35571);
and U46868 (N_46868,N_37717,N_39945);
nand U46869 (N_46869,N_38841,N_34167);
and U46870 (N_46870,N_30477,N_32741);
or U46871 (N_46871,N_38007,N_33054);
nand U46872 (N_46872,N_30458,N_36196);
and U46873 (N_46873,N_33774,N_33846);
nor U46874 (N_46874,N_39501,N_31450);
and U46875 (N_46875,N_30869,N_30092);
xnor U46876 (N_46876,N_34744,N_30315);
nand U46877 (N_46877,N_33019,N_33063);
and U46878 (N_46878,N_31836,N_35869);
and U46879 (N_46879,N_38572,N_32388);
nand U46880 (N_46880,N_35546,N_33883);
nor U46881 (N_46881,N_37330,N_38686);
nor U46882 (N_46882,N_34950,N_38931);
and U46883 (N_46883,N_30162,N_37785);
or U46884 (N_46884,N_37146,N_33436);
nand U46885 (N_46885,N_35861,N_39913);
or U46886 (N_46886,N_31138,N_36231);
nand U46887 (N_46887,N_30534,N_35668);
or U46888 (N_46888,N_33437,N_30610);
or U46889 (N_46889,N_36580,N_32703);
and U46890 (N_46890,N_38053,N_36421);
nor U46891 (N_46891,N_36004,N_33619);
and U46892 (N_46892,N_38611,N_35453);
and U46893 (N_46893,N_35314,N_33508);
nor U46894 (N_46894,N_35170,N_35275);
nor U46895 (N_46895,N_32407,N_37113);
nor U46896 (N_46896,N_33859,N_30650);
xor U46897 (N_46897,N_36969,N_32008);
or U46898 (N_46898,N_38715,N_39989);
or U46899 (N_46899,N_39202,N_39827);
and U46900 (N_46900,N_35590,N_37868);
and U46901 (N_46901,N_39586,N_32299);
or U46902 (N_46902,N_30764,N_37584);
and U46903 (N_46903,N_37648,N_30856);
xor U46904 (N_46904,N_31269,N_34676);
or U46905 (N_46905,N_36462,N_35485);
nor U46906 (N_46906,N_35019,N_38593);
and U46907 (N_46907,N_36445,N_31435);
xnor U46908 (N_46908,N_33460,N_39472);
and U46909 (N_46909,N_38943,N_37682);
nor U46910 (N_46910,N_35204,N_39038);
xor U46911 (N_46911,N_33198,N_33294);
and U46912 (N_46912,N_37037,N_34140);
or U46913 (N_46913,N_39709,N_38227);
nor U46914 (N_46914,N_35373,N_30400);
or U46915 (N_46915,N_32413,N_37136);
nand U46916 (N_46916,N_34600,N_31986);
or U46917 (N_46917,N_31957,N_36178);
and U46918 (N_46918,N_39712,N_38000);
or U46919 (N_46919,N_33065,N_34000);
nand U46920 (N_46920,N_31366,N_34752);
and U46921 (N_46921,N_31633,N_31881);
nand U46922 (N_46922,N_31464,N_30468);
or U46923 (N_46923,N_39324,N_37342);
xor U46924 (N_46924,N_37228,N_36163);
and U46925 (N_46925,N_39564,N_39325);
and U46926 (N_46926,N_39534,N_34244);
or U46927 (N_46927,N_39472,N_32341);
nor U46928 (N_46928,N_33833,N_35749);
xor U46929 (N_46929,N_30366,N_32934);
and U46930 (N_46930,N_38281,N_36564);
nor U46931 (N_46931,N_35993,N_37586);
or U46932 (N_46932,N_37013,N_32361);
or U46933 (N_46933,N_34488,N_36393);
or U46934 (N_46934,N_36270,N_31598);
and U46935 (N_46935,N_34810,N_39253);
nor U46936 (N_46936,N_37875,N_30591);
nand U46937 (N_46937,N_35488,N_37552);
nor U46938 (N_46938,N_37197,N_32171);
and U46939 (N_46939,N_32781,N_33100);
xnor U46940 (N_46940,N_39684,N_31747);
nand U46941 (N_46941,N_37193,N_39849);
nand U46942 (N_46942,N_31320,N_33143);
nand U46943 (N_46943,N_33280,N_37691);
nor U46944 (N_46944,N_31351,N_36295);
nand U46945 (N_46945,N_31828,N_37314);
xnor U46946 (N_46946,N_30386,N_34183);
nor U46947 (N_46947,N_33591,N_37560);
and U46948 (N_46948,N_30345,N_33334);
nor U46949 (N_46949,N_39056,N_31350);
nand U46950 (N_46950,N_35639,N_36605);
and U46951 (N_46951,N_31097,N_33991);
or U46952 (N_46952,N_30730,N_36571);
or U46953 (N_46953,N_39027,N_37718);
and U46954 (N_46954,N_37864,N_30227);
nand U46955 (N_46955,N_36835,N_32560);
nand U46956 (N_46956,N_35333,N_39818);
xor U46957 (N_46957,N_38068,N_39769);
xnor U46958 (N_46958,N_31247,N_39355);
nor U46959 (N_46959,N_38101,N_34394);
or U46960 (N_46960,N_38249,N_33061);
and U46961 (N_46961,N_31829,N_37597);
nand U46962 (N_46962,N_36427,N_33144);
or U46963 (N_46963,N_36353,N_33736);
nand U46964 (N_46964,N_39095,N_36243);
and U46965 (N_46965,N_38848,N_35172);
nand U46966 (N_46966,N_39072,N_38225);
xnor U46967 (N_46967,N_38684,N_39752);
nor U46968 (N_46968,N_31560,N_39232);
or U46969 (N_46969,N_32251,N_33351);
xnor U46970 (N_46970,N_30258,N_37289);
xor U46971 (N_46971,N_32638,N_30211);
or U46972 (N_46972,N_39474,N_36189);
nand U46973 (N_46973,N_31912,N_34516);
nor U46974 (N_46974,N_33105,N_39400);
or U46975 (N_46975,N_32980,N_37051);
nor U46976 (N_46976,N_33299,N_38649);
xnor U46977 (N_46977,N_39198,N_31279);
and U46978 (N_46978,N_36951,N_30356);
and U46979 (N_46979,N_35913,N_35402);
or U46980 (N_46980,N_30414,N_32147);
or U46981 (N_46981,N_36069,N_33964);
or U46982 (N_46982,N_38448,N_39158);
and U46983 (N_46983,N_36945,N_30327);
nand U46984 (N_46984,N_31387,N_32999);
xnor U46985 (N_46985,N_34047,N_37004);
or U46986 (N_46986,N_36350,N_38664);
xor U46987 (N_46987,N_39381,N_34213);
and U46988 (N_46988,N_32275,N_35816);
xnor U46989 (N_46989,N_37147,N_31114);
or U46990 (N_46990,N_37098,N_38711);
nor U46991 (N_46991,N_37824,N_39642);
xnor U46992 (N_46992,N_31827,N_34722);
and U46993 (N_46993,N_33007,N_30803);
nand U46994 (N_46994,N_32407,N_32096);
nand U46995 (N_46995,N_38229,N_36201);
and U46996 (N_46996,N_39997,N_35678);
nor U46997 (N_46997,N_36870,N_36239);
nor U46998 (N_46998,N_35224,N_32279);
nand U46999 (N_46999,N_33697,N_31172);
nand U47000 (N_47000,N_33646,N_33432);
nand U47001 (N_47001,N_37422,N_39304);
or U47002 (N_47002,N_30866,N_32602);
xor U47003 (N_47003,N_31807,N_30186);
and U47004 (N_47004,N_34094,N_30168);
and U47005 (N_47005,N_32492,N_35110);
nand U47006 (N_47006,N_31157,N_37782);
xor U47007 (N_47007,N_30599,N_30558);
and U47008 (N_47008,N_32241,N_36839);
xor U47009 (N_47009,N_31290,N_33751);
xor U47010 (N_47010,N_34714,N_34552);
nor U47011 (N_47011,N_37130,N_39628);
and U47012 (N_47012,N_39207,N_36694);
xor U47013 (N_47013,N_34761,N_38888);
nor U47014 (N_47014,N_37654,N_31817);
nor U47015 (N_47015,N_31393,N_31675);
nor U47016 (N_47016,N_39553,N_36181);
and U47017 (N_47017,N_33230,N_39535);
nor U47018 (N_47018,N_32488,N_37815);
or U47019 (N_47019,N_34082,N_37113);
or U47020 (N_47020,N_33783,N_31124);
nand U47021 (N_47021,N_30410,N_39356);
and U47022 (N_47022,N_35049,N_32345);
nor U47023 (N_47023,N_34281,N_31959);
nor U47024 (N_47024,N_34794,N_32740);
or U47025 (N_47025,N_32478,N_30283);
nand U47026 (N_47026,N_37092,N_37062);
nand U47027 (N_47027,N_34328,N_37040);
nor U47028 (N_47028,N_34316,N_32125);
nand U47029 (N_47029,N_30355,N_35352);
or U47030 (N_47030,N_32181,N_34755);
or U47031 (N_47031,N_32577,N_33963);
nor U47032 (N_47032,N_34564,N_39017);
or U47033 (N_47033,N_37420,N_38834);
xor U47034 (N_47034,N_33825,N_37711);
nor U47035 (N_47035,N_38704,N_34327);
or U47036 (N_47036,N_37865,N_36963);
nor U47037 (N_47037,N_34657,N_33220);
nand U47038 (N_47038,N_37484,N_38490);
and U47039 (N_47039,N_36356,N_32028);
or U47040 (N_47040,N_38204,N_35892);
and U47041 (N_47041,N_32998,N_32988);
nand U47042 (N_47042,N_35562,N_35876);
xnor U47043 (N_47043,N_38525,N_36623);
and U47044 (N_47044,N_39959,N_37154);
nor U47045 (N_47045,N_32789,N_38138);
or U47046 (N_47046,N_35383,N_38051);
and U47047 (N_47047,N_38671,N_33954);
or U47048 (N_47048,N_39814,N_39494);
nand U47049 (N_47049,N_35865,N_38344);
xnor U47050 (N_47050,N_35925,N_39880);
nand U47051 (N_47051,N_38041,N_39656);
or U47052 (N_47052,N_33058,N_32173);
nor U47053 (N_47053,N_36940,N_37303);
xor U47054 (N_47054,N_34443,N_31144);
nand U47055 (N_47055,N_34780,N_31807);
or U47056 (N_47056,N_36934,N_35469);
xor U47057 (N_47057,N_37469,N_37268);
nor U47058 (N_47058,N_33838,N_34431);
xnor U47059 (N_47059,N_39264,N_36199);
and U47060 (N_47060,N_33884,N_38164);
or U47061 (N_47061,N_30994,N_33547);
and U47062 (N_47062,N_32898,N_31898);
xnor U47063 (N_47063,N_36364,N_33402);
nand U47064 (N_47064,N_37242,N_33610);
or U47065 (N_47065,N_33047,N_31334);
nor U47066 (N_47066,N_34653,N_34121);
or U47067 (N_47067,N_33287,N_31288);
or U47068 (N_47068,N_31612,N_31644);
or U47069 (N_47069,N_36576,N_34180);
and U47070 (N_47070,N_34901,N_36157);
and U47071 (N_47071,N_34096,N_33887);
and U47072 (N_47072,N_38181,N_34376);
nand U47073 (N_47073,N_33906,N_39031);
and U47074 (N_47074,N_39746,N_36753);
nand U47075 (N_47075,N_34661,N_33545);
nand U47076 (N_47076,N_32903,N_37053);
nand U47077 (N_47077,N_38031,N_32508);
and U47078 (N_47078,N_36387,N_31439);
xnor U47079 (N_47079,N_34893,N_34558);
or U47080 (N_47080,N_37059,N_36367);
nand U47081 (N_47081,N_39092,N_31265);
and U47082 (N_47082,N_31530,N_36599);
or U47083 (N_47083,N_38808,N_30354);
and U47084 (N_47084,N_31370,N_35035);
xor U47085 (N_47085,N_38993,N_36821);
or U47086 (N_47086,N_31854,N_35809);
or U47087 (N_47087,N_35069,N_36746);
xor U47088 (N_47088,N_37080,N_34364);
nor U47089 (N_47089,N_35687,N_37352);
and U47090 (N_47090,N_38212,N_35753);
xor U47091 (N_47091,N_38274,N_33936);
nand U47092 (N_47092,N_34142,N_37909);
xnor U47093 (N_47093,N_30613,N_30894);
nor U47094 (N_47094,N_31605,N_31283);
xor U47095 (N_47095,N_32986,N_34582);
nor U47096 (N_47096,N_30102,N_38158);
xor U47097 (N_47097,N_34076,N_33704);
nand U47098 (N_47098,N_31599,N_32032);
nand U47099 (N_47099,N_36982,N_35383);
nor U47100 (N_47100,N_36455,N_37901);
nor U47101 (N_47101,N_30411,N_30327);
or U47102 (N_47102,N_36988,N_33085);
or U47103 (N_47103,N_38904,N_33655);
and U47104 (N_47104,N_36540,N_38343);
nand U47105 (N_47105,N_35930,N_38339);
and U47106 (N_47106,N_38385,N_39632);
nor U47107 (N_47107,N_32150,N_33724);
nand U47108 (N_47108,N_36033,N_37583);
xnor U47109 (N_47109,N_34133,N_35948);
or U47110 (N_47110,N_30467,N_36268);
xnor U47111 (N_47111,N_33564,N_34463);
xor U47112 (N_47112,N_31767,N_34843);
and U47113 (N_47113,N_39722,N_30634);
or U47114 (N_47114,N_35114,N_38151);
nor U47115 (N_47115,N_30139,N_39464);
nor U47116 (N_47116,N_32985,N_36408);
xor U47117 (N_47117,N_32016,N_36539);
nand U47118 (N_47118,N_36547,N_32699);
nor U47119 (N_47119,N_33805,N_31444);
nand U47120 (N_47120,N_31341,N_33238);
nor U47121 (N_47121,N_33846,N_38294);
nor U47122 (N_47122,N_39140,N_37192);
nand U47123 (N_47123,N_37102,N_30423);
or U47124 (N_47124,N_39047,N_36738);
xor U47125 (N_47125,N_37034,N_33360);
and U47126 (N_47126,N_35017,N_37902);
or U47127 (N_47127,N_32119,N_36397);
or U47128 (N_47128,N_33558,N_33715);
and U47129 (N_47129,N_34857,N_33687);
nor U47130 (N_47130,N_34673,N_33924);
nand U47131 (N_47131,N_33896,N_32848);
or U47132 (N_47132,N_36734,N_37991);
and U47133 (N_47133,N_34025,N_31285);
and U47134 (N_47134,N_34326,N_34308);
xnor U47135 (N_47135,N_32618,N_35772);
nand U47136 (N_47136,N_30952,N_33340);
nand U47137 (N_47137,N_30584,N_32375);
nor U47138 (N_47138,N_33961,N_38881);
nand U47139 (N_47139,N_33908,N_31415);
xor U47140 (N_47140,N_37186,N_30574);
nor U47141 (N_47141,N_39101,N_36207);
and U47142 (N_47142,N_32301,N_37016);
and U47143 (N_47143,N_33604,N_36243);
xor U47144 (N_47144,N_31514,N_39084);
or U47145 (N_47145,N_36308,N_37038);
and U47146 (N_47146,N_38981,N_37185);
and U47147 (N_47147,N_31013,N_35399);
nor U47148 (N_47148,N_38614,N_32930);
xnor U47149 (N_47149,N_31977,N_37364);
and U47150 (N_47150,N_37535,N_30746);
xnor U47151 (N_47151,N_38390,N_31832);
nor U47152 (N_47152,N_39853,N_34515);
or U47153 (N_47153,N_34587,N_35083);
xor U47154 (N_47154,N_35270,N_38464);
nand U47155 (N_47155,N_34990,N_31717);
xnor U47156 (N_47156,N_39767,N_34787);
and U47157 (N_47157,N_32481,N_36257);
and U47158 (N_47158,N_39051,N_35465);
xnor U47159 (N_47159,N_38883,N_35750);
or U47160 (N_47160,N_35060,N_35118);
xor U47161 (N_47161,N_36669,N_33170);
or U47162 (N_47162,N_31742,N_34225);
xnor U47163 (N_47163,N_32944,N_31857);
xnor U47164 (N_47164,N_34650,N_38201);
xor U47165 (N_47165,N_39364,N_34818);
and U47166 (N_47166,N_32179,N_31121);
or U47167 (N_47167,N_31592,N_34662);
and U47168 (N_47168,N_32400,N_31957);
nor U47169 (N_47169,N_38788,N_32560);
xnor U47170 (N_47170,N_30108,N_30500);
nand U47171 (N_47171,N_37879,N_32989);
or U47172 (N_47172,N_36011,N_34263);
nand U47173 (N_47173,N_35979,N_34927);
or U47174 (N_47174,N_30019,N_31741);
or U47175 (N_47175,N_32940,N_34400);
nor U47176 (N_47176,N_31275,N_31981);
nand U47177 (N_47177,N_32527,N_34735);
or U47178 (N_47178,N_35345,N_37415);
nand U47179 (N_47179,N_33951,N_31780);
nor U47180 (N_47180,N_35500,N_32304);
xnor U47181 (N_47181,N_34532,N_39633);
or U47182 (N_47182,N_32371,N_38611);
nor U47183 (N_47183,N_33741,N_31728);
and U47184 (N_47184,N_31883,N_38741);
and U47185 (N_47185,N_33866,N_37511);
and U47186 (N_47186,N_36552,N_39261);
nor U47187 (N_47187,N_30281,N_38762);
nor U47188 (N_47188,N_33585,N_30972);
and U47189 (N_47189,N_34209,N_34642);
and U47190 (N_47190,N_35740,N_33625);
and U47191 (N_47191,N_37450,N_35569);
or U47192 (N_47192,N_34591,N_36835);
xor U47193 (N_47193,N_34036,N_31462);
nor U47194 (N_47194,N_30623,N_36454);
nand U47195 (N_47195,N_36205,N_39347);
or U47196 (N_47196,N_34429,N_31990);
nand U47197 (N_47197,N_32399,N_33802);
nand U47198 (N_47198,N_30446,N_32709);
nor U47199 (N_47199,N_33152,N_34735);
xnor U47200 (N_47200,N_31241,N_34031);
and U47201 (N_47201,N_31359,N_35250);
nor U47202 (N_47202,N_33037,N_36134);
nand U47203 (N_47203,N_33030,N_37787);
or U47204 (N_47204,N_32580,N_34670);
xor U47205 (N_47205,N_32866,N_37319);
nand U47206 (N_47206,N_37899,N_35858);
xor U47207 (N_47207,N_32758,N_39361);
nor U47208 (N_47208,N_37252,N_30372);
and U47209 (N_47209,N_33146,N_31151);
nor U47210 (N_47210,N_36062,N_38773);
or U47211 (N_47211,N_34103,N_38020);
nor U47212 (N_47212,N_39556,N_32154);
and U47213 (N_47213,N_34112,N_30975);
or U47214 (N_47214,N_34475,N_36965);
and U47215 (N_47215,N_39098,N_37232);
nor U47216 (N_47216,N_30435,N_37804);
nand U47217 (N_47217,N_38445,N_34726);
or U47218 (N_47218,N_33642,N_38142);
xor U47219 (N_47219,N_37443,N_37652);
or U47220 (N_47220,N_33242,N_39583);
nor U47221 (N_47221,N_36442,N_38232);
xor U47222 (N_47222,N_32866,N_37904);
nor U47223 (N_47223,N_38663,N_30056);
nand U47224 (N_47224,N_36215,N_37097);
nand U47225 (N_47225,N_30055,N_35496);
nand U47226 (N_47226,N_37425,N_30308);
nand U47227 (N_47227,N_35860,N_37149);
and U47228 (N_47228,N_34718,N_38557);
nand U47229 (N_47229,N_30236,N_34265);
xor U47230 (N_47230,N_31717,N_33438);
nor U47231 (N_47231,N_36918,N_32986);
nand U47232 (N_47232,N_35010,N_37729);
nand U47233 (N_47233,N_33424,N_39670);
nand U47234 (N_47234,N_31998,N_31364);
and U47235 (N_47235,N_33450,N_35447);
and U47236 (N_47236,N_30830,N_34600);
and U47237 (N_47237,N_35319,N_39206);
and U47238 (N_47238,N_31593,N_35173);
nand U47239 (N_47239,N_32131,N_34162);
and U47240 (N_47240,N_33004,N_34571);
and U47241 (N_47241,N_39862,N_30255);
or U47242 (N_47242,N_30643,N_34538);
or U47243 (N_47243,N_36579,N_33462);
nand U47244 (N_47244,N_38572,N_31305);
nor U47245 (N_47245,N_37755,N_34731);
nand U47246 (N_47246,N_38178,N_32984);
nand U47247 (N_47247,N_34088,N_35239);
nor U47248 (N_47248,N_33191,N_32121);
nor U47249 (N_47249,N_32526,N_36165);
and U47250 (N_47250,N_33271,N_38612);
and U47251 (N_47251,N_37278,N_38501);
xor U47252 (N_47252,N_31778,N_31053);
nand U47253 (N_47253,N_33990,N_32293);
xnor U47254 (N_47254,N_37756,N_38324);
and U47255 (N_47255,N_30120,N_32888);
or U47256 (N_47256,N_36261,N_33064);
and U47257 (N_47257,N_35697,N_31529);
and U47258 (N_47258,N_31599,N_35275);
and U47259 (N_47259,N_32177,N_38046);
or U47260 (N_47260,N_33116,N_35465);
nand U47261 (N_47261,N_31366,N_37517);
xnor U47262 (N_47262,N_30245,N_37638);
nor U47263 (N_47263,N_39735,N_36033);
and U47264 (N_47264,N_33339,N_30078);
xor U47265 (N_47265,N_35205,N_31960);
nand U47266 (N_47266,N_32398,N_38634);
nand U47267 (N_47267,N_30650,N_39711);
and U47268 (N_47268,N_36637,N_30111);
nor U47269 (N_47269,N_30115,N_39446);
xor U47270 (N_47270,N_32061,N_32471);
xor U47271 (N_47271,N_33960,N_37575);
or U47272 (N_47272,N_36994,N_34240);
nor U47273 (N_47273,N_36025,N_31192);
and U47274 (N_47274,N_32514,N_39412);
and U47275 (N_47275,N_38834,N_33904);
nor U47276 (N_47276,N_38817,N_31084);
and U47277 (N_47277,N_37590,N_30996);
xnor U47278 (N_47278,N_33102,N_34455);
nor U47279 (N_47279,N_37316,N_32984);
xor U47280 (N_47280,N_38416,N_37863);
and U47281 (N_47281,N_39967,N_36765);
and U47282 (N_47282,N_36269,N_30072);
or U47283 (N_47283,N_34255,N_30790);
nand U47284 (N_47284,N_34641,N_39294);
xnor U47285 (N_47285,N_31848,N_31188);
and U47286 (N_47286,N_30893,N_38281);
nor U47287 (N_47287,N_36039,N_31739);
nor U47288 (N_47288,N_39846,N_36864);
or U47289 (N_47289,N_34273,N_39181);
xnor U47290 (N_47290,N_32812,N_35648);
nand U47291 (N_47291,N_35000,N_37958);
and U47292 (N_47292,N_32309,N_30107);
and U47293 (N_47293,N_38758,N_37434);
xor U47294 (N_47294,N_34266,N_36085);
nor U47295 (N_47295,N_36716,N_38342);
and U47296 (N_47296,N_36285,N_35269);
xor U47297 (N_47297,N_30071,N_35969);
nand U47298 (N_47298,N_34441,N_36781);
and U47299 (N_47299,N_32597,N_37607);
or U47300 (N_47300,N_35836,N_31693);
or U47301 (N_47301,N_33194,N_34725);
or U47302 (N_47302,N_37365,N_34460);
and U47303 (N_47303,N_32750,N_33918);
and U47304 (N_47304,N_38885,N_38428);
nor U47305 (N_47305,N_35229,N_31247);
xor U47306 (N_47306,N_30571,N_39599);
xnor U47307 (N_47307,N_34620,N_34230);
xnor U47308 (N_47308,N_30902,N_34191);
nand U47309 (N_47309,N_31268,N_35122);
nand U47310 (N_47310,N_39410,N_34616);
nor U47311 (N_47311,N_38948,N_35211);
and U47312 (N_47312,N_31506,N_35346);
or U47313 (N_47313,N_34962,N_30953);
xor U47314 (N_47314,N_34529,N_35038);
or U47315 (N_47315,N_37788,N_33848);
nor U47316 (N_47316,N_33841,N_39022);
and U47317 (N_47317,N_36879,N_37293);
and U47318 (N_47318,N_33652,N_36171);
and U47319 (N_47319,N_38542,N_32853);
nand U47320 (N_47320,N_30177,N_37973);
nor U47321 (N_47321,N_31969,N_39640);
nand U47322 (N_47322,N_30317,N_34662);
nor U47323 (N_47323,N_37238,N_38952);
nor U47324 (N_47324,N_33160,N_33925);
and U47325 (N_47325,N_30402,N_35802);
nor U47326 (N_47326,N_35460,N_30468);
nor U47327 (N_47327,N_39986,N_34989);
nand U47328 (N_47328,N_32276,N_31946);
and U47329 (N_47329,N_34018,N_37372);
or U47330 (N_47330,N_32956,N_36962);
nand U47331 (N_47331,N_39012,N_39517);
or U47332 (N_47332,N_35571,N_38656);
or U47333 (N_47333,N_32266,N_30171);
xor U47334 (N_47334,N_31984,N_37035);
xnor U47335 (N_47335,N_38702,N_37760);
nand U47336 (N_47336,N_38440,N_30714);
or U47337 (N_47337,N_35440,N_31547);
nor U47338 (N_47338,N_35899,N_35209);
and U47339 (N_47339,N_37451,N_32537);
or U47340 (N_47340,N_32359,N_38771);
nor U47341 (N_47341,N_34802,N_33533);
and U47342 (N_47342,N_34205,N_31053);
or U47343 (N_47343,N_38290,N_30057);
nor U47344 (N_47344,N_33960,N_34833);
or U47345 (N_47345,N_32561,N_38269);
nor U47346 (N_47346,N_34758,N_35626);
nor U47347 (N_47347,N_33579,N_35589);
and U47348 (N_47348,N_37354,N_31787);
nand U47349 (N_47349,N_35919,N_30726);
nor U47350 (N_47350,N_39246,N_31251);
or U47351 (N_47351,N_33958,N_34829);
nor U47352 (N_47352,N_32173,N_30996);
xnor U47353 (N_47353,N_33257,N_30944);
and U47354 (N_47354,N_36520,N_39266);
nand U47355 (N_47355,N_31826,N_39690);
and U47356 (N_47356,N_39347,N_33580);
and U47357 (N_47357,N_33195,N_30859);
xnor U47358 (N_47358,N_33254,N_36619);
and U47359 (N_47359,N_32916,N_30235);
xnor U47360 (N_47360,N_35325,N_32271);
xor U47361 (N_47361,N_34096,N_34461);
xnor U47362 (N_47362,N_39418,N_30620);
and U47363 (N_47363,N_38718,N_38373);
or U47364 (N_47364,N_33453,N_36335);
xnor U47365 (N_47365,N_35506,N_38602);
or U47366 (N_47366,N_37763,N_33430);
nand U47367 (N_47367,N_30652,N_39152);
and U47368 (N_47368,N_30307,N_38095);
nor U47369 (N_47369,N_32838,N_31997);
or U47370 (N_47370,N_30258,N_39172);
nand U47371 (N_47371,N_31028,N_36851);
and U47372 (N_47372,N_31988,N_37534);
or U47373 (N_47373,N_30029,N_39879);
nor U47374 (N_47374,N_38863,N_33530);
and U47375 (N_47375,N_38122,N_32414);
nand U47376 (N_47376,N_36809,N_35511);
nand U47377 (N_47377,N_38569,N_33610);
nand U47378 (N_47378,N_32007,N_39642);
and U47379 (N_47379,N_38820,N_33700);
nor U47380 (N_47380,N_30201,N_33373);
nor U47381 (N_47381,N_36718,N_31285);
and U47382 (N_47382,N_38018,N_39557);
xnor U47383 (N_47383,N_38007,N_34715);
nor U47384 (N_47384,N_33203,N_31114);
or U47385 (N_47385,N_39499,N_32100);
nand U47386 (N_47386,N_31382,N_35260);
nor U47387 (N_47387,N_34003,N_33770);
or U47388 (N_47388,N_36254,N_31895);
or U47389 (N_47389,N_33100,N_32510);
nand U47390 (N_47390,N_30923,N_32414);
nand U47391 (N_47391,N_35113,N_36993);
xor U47392 (N_47392,N_38197,N_39489);
nand U47393 (N_47393,N_32268,N_30477);
and U47394 (N_47394,N_33556,N_32131);
xor U47395 (N_47395,N_37646,N_39992);
or U47396 (N_47396,N_34289,N_35504);
and U47397 (N_47397,N_33440,N_31643);
nor U47398 (N_47398,N_37384,N_35870);
nand U47399 (N_47399,N_38193,N_36031);
nand U47400 (N_47400,N_34658,N_38631);
or U47401 (N_47401,N_33356,N_39100);
xnor U47402 (N_47402,N_37215,N_31269);
or U47403 (N_47403,N_38897,N_30729);
nor U47404 (N_47404,N_39088,N_38055);
or U47405 (N_47405,N_36247,N_30836);
or U47406 (N_47406,N_34672,N_32166);
nor U47407 (N_47407,N_38506,N_39271);
nand U47408 (N_47408,N_34583,N_30914);
nor U47409 (N_47409,N_39746,N_30930);
or U47410 (N_47410,N_35761,N_32066);
and U47411 (N_47411,N_39743,N_36465);
nor U47412 (N_47412,N_36116,N_35921);
and U47413 (N_47413,N_34630,N_32054);
nand U47414 (N_47414,N_30434,N_33772);
or U47415 (N_47415,N_32749,N_38640);
and U47416 (N_47416,N_36099,N_36413);
xor U47417 (N_47417,N_33113,N_32354);
and U47418 (N_47418,N_33309,N_37935);
or U47419 (N_47419,N_33193,N_39756);
xnor U47420 (N_47420,N_34214,N_36982);
nand U47421 (N_47421,N_38642,N_36541);
or U47422 (N_47422,N_39907,N_38447);
nor U47423 (N_47423,N_31611,N_35352);
or U47424 (N_47424,N_31234,N_35404);
nor U47425 (N_47425,N_38451,N_36699);
nand U47426 (N_47426,N_30588,N_30081);
nand U47427 (N_47427,N_35078,N_32426);
or U47428 (N_47428,N_30399,N_35361);
and U47429 (N_47429,N_39859,N_31514);
or U47430 (N_47430,N_37461,N_35264);
xor U47431 (N_47431,N_38086,N_37303);
or U47432 (N_47432,N_34208,N_36219);
nor U47433 (N_47433,N_38376,N_38492);
and U47434 (N_47434,N_38221,N_36415);
nor U47435 (N_47435,N_36126,N_33294);
or U47436 (N_47436,N_30574,N_33640);
and U47437 (N_47437,N_32790,N_35210);
nand U47438 (N_47438,N_30798,N_36723);
and U47439 (N_47439,N_36621,N_37949);
nand U47440 (N_47440,N_39512,N_32859);
nor U47441 (N_47441,N_31054,N_30734);
or U47442 (N_47442,N_39172,N_37097);
and U47443 (N_47443,N_34463,N_30779);
or U47444 (N_47444,N_33511,N_31707);
nand U47445 (N_47445,N_36888,N_33267);
or U47446 (N_47446,N_31114,N_38924);
nor U47447 (N_47447,N_39339,N_34945);
nand U47448 (N_47448,N_30401,N_35567);
xnor U47449 (N_47449,N_31561,N_38369);
nand U47450 (N_47450,N_33283,N_32865);
xor U47451 (N_47451,N_39349,N_33372);
or U47452 (N_47452,N_34758,N_36308);
and U47453 (N_47453,N_38439,N_35463);
nor U47454 (N_47454,N_33753,N_39266);
nand U47455 (N_47455,N_38622,N_34941);
or U47456 (N_47456,N_31109,N_35448);
and U47457 (N_47457,N_33587,N_36695);
or U47458 (N_47458,N_36444,N_30775);
nor U47459 (N_47459,N_34133,N_30938);
or U47460 (N_47460,N_31013,N_37250);
xnor U47461 (N_47461,N_39540,N_37753);
xnor U47462 (N_47462,N_30111,N_34673);
nand U47463 (N_47463,N_37130,N_34953);
nor U47464 (N_47464,N_34860,N_36746);
and U47465 (N_47465,N_30306,N_38315);
xnor U47466 (N_47466,N_30338,N_38904);
xnor U47467 (N_47467,N_33237,N_37451);
and U47468 (N_47468,N_37370,N_36757);
xnor U47469 (N_47469,N_36336,N_39019);
nand U47470 (N_47470,N_32457,N_34409);
nand U47471 (N_47471,N_31553,N_32160);
or U47472 (N_47472,N_30390,N_35453);
xor U47473 (N_47473,N_30626,N_32935);
or U47474 (N_47474,N_37922,N_31208);
or U47475 (N_47475,N_31678,N_39876);
nor U47476 (N_47476,N_38307,N_35841);
xor U47477 (N_47477,N_32854,N_37686);
and U47478 (N_47478,N_36478,N_32728);
nor U47479 (N_47479,N_39162,N_36641);
or U47480 (N_47480,N_31462,N_37351);
xor U47481 (N_47481,N_39956,N_35367);
nand U47482 (N_47482,N_31945,N_39519);
nor U47483 (N_47483,N_38521,N_33507);
or U47484 (N_47484,N_37257,N_34659);
or U47485 (N_47485,N_33728,N_35791);
nand U47486 (N_47486,N_34177,N_31682);
nand U47487 (N_47487,N_33650,N_32959);
nand U47488 (N_47488,N_38047,N_36803);
and U47489 (N_47489,N_38664,N_36745);
nand U47490 (N_47490,N_38736,N_36446);
and U47491 (N_47491,N_30181,N_36673);
or U47492 (N_47492,N_38979,N_35829);
nand U47493 (N_47493,N_39933,N_30637);
xnor U47494 (N_47494,N_32098,N_36981);
or U47495 (N_47495,N_39990,N_34201);
nand U47496 (N_47496,N_39227,N_35597);
or U47497 (N_47497,N_37086,N_30318);
nor U47498 (N_47498,N_38631,N_31925);
nand U47499 (N_47499,N_32176,N_38913);
or U47500 (N_47500,N_32426,N_34691);
and U47501 (N_47501,N_37867,N_36761);
xor U47502 (N_47502,N_39201,N_34449);
nor U47503 (N_47503,N_33848,N_36769);
nor U47504 (N_47504,N_39611,N_32660);
nor U47505 (N_47505,N_35638,N_31074);
nand U47506 (N_47506,N_36361,N_30456);
nand U47507 (N_47507,N_35150,N_33873);
or U47508 (N_47508,N_34308,N_38153);
nand U47509 (N_47509,N_37840,N_36986);
and U47510 (N_47510,N_37911,N_30807);
nand U47511 (N_47511,N_39550,N_37054);
and U47512 (N_47512,N_36076,N_30504);
or U47513 (N_47513,N_35691,N_34723);
nor U47514 (N_47514,N_31250,N_30717);
nor U47515 (N_47515,N_32239,N_32761);
nand U47516 (N_47516,N_37303,N_36009);
nor U47517 (N_47517,N_31773,N_34971);
nor U47518 (N_47518,N_34503,N_38640);
nor U47519 (N_47519,N_33284,N_36096);
and U47520 (N_47520,N_33842,N_33373);
and U47521 (N_47521,N_37244,N_30512);
or U47522 (N_47522,N_39785,N_35118);
xor U47523 (N_47523,N_33476,N_39202);
and U47524 (N_47524,N_39553,N_32747);
nor U47525 (N_47525,N_30753,N_39647);
xor U47526 (N_47526,N_30956,N_33682);
nor U47527 (N_47527,N_39886,N_34226);
or U47528 (N_47528,N_34499,N_38679);
or U47529 (N_47529,N_35731,N_34273);
xnor U47530 (N_47530,N_36674,N_32732);
nand U47531 (N_47531,N_32019,N_33891);
xor U47532 (N_47532,N_35093,N_38578);
or U47533 (N_47533,N_31193,N_30779);
xor U47534 (N_47534,N_33977,N_36700);
or U47535 (N_47535,N_33192,N_39897);
and U47536 (N_47536,N_36467,N_37538);
or U47537 (N_47537,N_37695,N_39655);
and U47538 (N_47538,N_37570,N_32750);
nand U47539 (N_47539,N_31983,N_33129);
nand U47540 (N_47540,N_35528,N_32539);
nand U47541 (N_47541,N_35369,N_31413);
nor U47542 (N_47542,N_37379,N_30280);
nand U47543 (N_47543,N_39997,N_38407);
nor U47544 (N_47544,N_33962,N_37719);
nor U47545 (N_47545,N_39550,N_30300);
or U47546 (N_47546,N_30765,N_31405);
and U47547 (N_47547,N_31541,N_35794);
and U47548 (N_47548,N_38404,N_38359);
nand U47549 (N_47549,N_32890,N_36882);
and U47550 (N_47550,N_32426,N_39020);
or U47551 (N_47551,N_32718,N_35866);
xnor U47552 (N_47552,N_39549,N_38276);
nor U47553 (N_47553,N_30057,N_36469);
nand U47554 (N_47554,N_36607,N_37744);
nand U47555 (N_47555,N_35349,N_37210);
nor U47556 (N_47556,N_38080,N_36890);
nor U47557 (N_47557,N_34119,N_32636);
or U47558 (N_47558,N_30714,N_31791);
or U47559 (N_47559,N_34192,N_30794);
xor U47560 (N_47560,N_33223,N_34915);
or U47561 (N_47561,N_31335,N_30983);
and U47562 (N_47562,N_35145,N_38370);
nand U47563 (N_47563,N_30902,N_39372);
and U47564 (N_47564,N_32554,N_31035);
nor U47565 (N_47565,N_32589,N_32538);
or U47566 (N_47566,N_30527,N_35697);
nor U47567 (N_47567,N_39939,N_31761);
xnor U47568 (N_47568,N_33805,N_38031);
nand U47569 (N_47569,N_32891,N_35584);
nor U47570 (N_47570,N_33124,N_31582);
nand U47571 (N_47571,N_39022,N_36283);
nor U47572 (N_47572,N_39328,N_32154);
xnor U47573 (N_47573,N_36862,N_35753);
nand U47574 (N_47574,N_31343,N_33859);
nand U47575 (N_47575,N_37989,N_30788);
or U47576 (N_47576,N_31659,N_39989);
nand U47577 (N_47577,N_36596,N_35609);
nand U47578 (N_47578,N_34138,N_33018);
or U47579 (N_47579,N_37172,N_31470);
and U47580 (N_47580,N_37699,N_35073);
xor U47581 (N_47581,N_35541,N_37436);
xnor U47582 (N_47582,N_38716,N_38060);
xnor U47583 (N_47583,N_33277,N_31118);
or U47584 (N_47584,N_38061,N_38405);
and U47585 (N_47585,N_33650,N_35428);
nor U47586 (N_47586,N_37383,N_39514);
xnor U47587 (N_47587,N_31664,N_31182);
nor U47588 (N_47588,N_36926,N_38984);
nand U47589 (N_47589,N_30714,N_37676);
or U47590 (N_47590,N_33840,N_32005);
nor U47591 (N_47591,N_31140,N_35430);
or U47592 (N_47592,N_30993,N_39448);
or U47593 (N_47593,N_37174,N_36409);
or U47594 (N_47594,N_33349,N_35521);
and U47595 (N_47595,N_30939,N_38859);
or U47596 (N_47596,N_34616,N_31868);
xor U47597 (N_47597,N_39063,N_30983);
and U47598 (N_47598,N_37129,N_36372);
or U47599 (N_47599,N_35847,N_38355);
xor U47600 (N_47600,N_38745,N_39021);
nand U47601 (N_47601,N_30830,N_38008);
or U47602 (N_47602,N_31196,N_33061);
or U47603 (N_47603,N_32790,N_33714);
nand U47604 (N_47604,N_32914,N_35251);
and U47605 (N_47605,N_31883,N_37431);
or U47606 (N_47606,N_30736,N_30895);
nand U47607 (N_47607,N_31182,N_32711);
nor U47608 (N_47608,N_35318,N_38092);
xor U47609 (N_47609,N_34048,N_33493);
or U47610 (N_47610,N_34198,N_38204);
nand U47611 (N_47611,N_39622,N_30437);
or U47612 (N_47612,N_31564,N_31149);
and U47613 (N_47613,N_30296,N_35756);
xor U47614 (N_47614,N_38111,N_31297);
xor U47615 (N_47615,N_37983,N_39919);
nand U47616 (N_47616,N_30685,N_37770);
nand U47617 (N_47617,N_38549,N_32885);
nor U47618 (N_47618,N_36339,N_39720);
and U47619 (N_47619,N_34980,N_31603);
nand U47620 (N_47620,N_33422,N_37168);
and U47621 (N_47621,N_34891,N_31638);
nor U47622 (N_47622,N_32135,N_33590);
and U47623 (N_47623,N_39311,N_34543);
or U47624 (N_47624,N_39876,N_37109);
nand U47625 (N_47625,N_33624,N_33351);
or U47626 (N_47626,N_37374,N_34367);
nor U47627 (N_47627,N_33475,N_35353);
nand U47628 (N_47628,N_31755,N_39718);
nor U47629 (N_47629,N_32983,N_36426);
nor U47630 (N_47630,N_36083,N_31912);
and U47631 (N_47631,N_35586,N_34729);
nor U47632 (N_47632,N_34822,N_39484);
and U47633 (N_47633,N_39398,N_38393);
xor U47634 (N_47634,N_32617,N_32252);
nand U47635 (N_47635,N_30941,N_39638);
nand U47636 (N_47636,N_37252,N_31587);
and U47637 (N_47637,N_34793,N_39968);
nand U47638 (N_47638,N_35686,N_30198);
nand U47639 (N_47639,N_36810,N_38033);
nor U47640 (N_47640,N_37077,N_38473);
and U47641 (N_47641,N_38909,N_30214);
nand U47642 (N_47642,N_32619,N_36176);
nand U47643 (N_47643,N_31994,N_34778);
nor U47644 (N_47644,N_31016,N_38198);
xnor U47645 (N_47645,N_34157,N_38754);
nor U47646 (N_47646,N_38411,N_34584);
nor U47647 (N_47647,N_36423,N_33285);
xor U47648 (N_47648,N_32077,N_37482);
xor U47649 (N_47649,N_32541,N_38819);
or U47650 (N_47650,N_34811,N_38956);
and U47651 (N_47651,N_32814,N_37496);
xor U47652 (N_47652,N_39078,N_30105);
nand U47653 (N_47653,N_38226,N_36580);
and U47654 (N_47654,N_35940,N_37903);
nand U47655 (N_47655,N_34646,N_36451);
nor U47656 (N_47656,N_36662,N_32725);
xor U47657 (N_47657,N_37950,N_39786);
xnor U47658 (N_47658,N_31419,N_39403);
xor U47659 (N_47659,N_33133,N_33970);
and U47660 (N_47660,N_31824,N_32876);
nand U47661 (N_47661,N_31666,N_31139);
or U47662 (N_47662,N_39997,N_31405);
and U47663 (N_47663,N_30429,N_38825);
xor U47664 (N_47664,N_38971,N_30916);
and U47665 (N_47665,N_32769,N_33999);
and U47666 (N_47666,N_32974,N_30073);
or U47667 (N_47667,N_30305,N_34247);
and U47668 (N_47668,N_35090,N_34459);
nand U47669 (N_47669,N_34285,N_32907);
and U47670 (N_47670,N_32985,N_33374);
or U47671 (N_47671,N_33098,N_35166);
or U47672 (N_47672,N_35707,N_30741);
xor U47673 (N_47673,N_35792,N_39107);
nor U47674 (N_47674,N_31353,N_39406);
and U47675 (N_47675,N_31593,N_32380);
xor U47676 (N_47676,N_30224,N_38294);
or U47677 (N_47677,N_30326,N_30816);
nor U47678 (N_47678,N_31995,N_38665);
nand U47679 (N_47679,N_32002,N_35447);
xnor U47680 (N_47680,N_32020,N_39052);
xor U47681 (N_47681,N_36723,N_39188);
and U47682 (N_47682,N_38991,N_32009);
nor U47683 (N_47683,N_34302,N_33556);
and U47684 (N_47684,N_33328,N_31496);
xor U47685 (N_47685,N_37234,N_39414);
or U47686 (N_47686,N_38325,N_37955);
xor U47687 (N_47687,N_32641,N_39023);
or U47688 (N_47688,N_32672,N_35382);
and U47689 (N_47689,N_33405,N_38152);
and U47690 (N_47690,N_30544,N_36822);
xnor U47691 (N_47691,N_32593,N_31886);
nor U47692 (N_47692,N_31986,N_37531);
nand U47693 (N_47693,N_39194,N_31070);
nand U47694 (N_47694,N_32858,N_37831);
xor U47695 (N_47695,N_37039,N_39927);
or U47696 (N_47696,N_39178,N_38211);
nor U47697 (N_47697,N_30973,N_36815);
and U47698 (N_47698,N_33989,N_31551);
xor U47699 (N_47699,N_38880,N_36398);
xor U47700 (N_47700,N_33771,N_39340);
nor U47701 (N_47701,N_30061,N_30228);
nor U47702 (N_47702,N_39485,N_34290);
nand U47703 (N_47703,N_35337,N_34626);
and U47704 (N_47704,N_34585,N_34259);
and U47705 (N_47705,N_39574,N_30129);
and U47706 (N_47706,N_32547,N_39907);
nand U47707 (N_47707,N_34585,N_36513);
xor U47708 (N_47708,N_34592,N_35867);
xnor U47709 (N_47709,N_36004,N_33925);
nor U47710 (N_47710,N_39198,N_32300);
and U47711 (N_47711,N_36652,N_31202);
xnor U47712 (N_47712,N_39895,N_39131);
nor U47713 (N_47713,N_32723,N_36939);
xor U47714 (N_47714,N_38026,N_33798);
and U47715 (N_47715,N_36093,N_36811);
xor U47716 (N_47716,N_32700,N_33335);
xnor U47717 (N_47717,N_30763,N_32417);
nor U47718 (N_47718,N_35651,N_31419);
and U47719 (N_47719,N_31874,N_37726);
and U47720 (N_47720,N_33263,N_32673);
xnor U47721 (N_47721,N_33674,N_35417);
nor U47722 (N_47722,N_35112,N_32921);
or U47723 (N_47723,N_38597,N_35990);
xor U47724 (N_47724,N_33941,N_30871);
xnor U47725 (N_47725,N_33762,N_38746);
xor U47726 (N_47726,N_34526,N_34259);
nor U47727 (N_47727,N_30295,N_32490);
and U47728 (N_47728,N_31731,N_32669);
and U47729 (N_47729,N_34512,N_38305);
and U47730 (N_47730,N_30536,N_36337);
nor U47731 (N_47731,N_31281,N_38372);
or U47732 (N_47732,N_35538,N_30688);
nand U47733 (N_47733,N_35244,N_37617);
nand U47734 (N_47734,N_38844,N_35837);
or U47735 (N_47735,N_38646,N_31755);
or U47736 (N_47736,N_30524,N_38407);
nor U47737 (N_47737,N_39250,N_32061);
nand U47738 (N_47738,N_38940,N_31787);
xor U47739 (N_47739,N_38576,N_31603);
xnor U47740 (N_47740,N_38467,N_39230);
nor U47741 (N_47741,N_32196,N_32048);
nor U47742 (N_47742,N_35961,N_33082);
and U47743 (N_47743,N_35673,N_31902);
or U47744 (N_47744,N_38372,N_36032);
xnor U47745 (N_47745,N_37086,N_38990);
or U47746 (N_47746,N_31642,N_37847);
nand U47747 (N_47747,N_35131,N_31058);
and U47748 (N_47748,N_32271,N_39853);
xor U47749 (N_47749,N_38166,N_33491);
or U47750 (N_47750,N_38346,N_31483);
nor U47751 (N_47751,N_37256,N_32406);
nor U47752 (N_47752,N_36099,N_33642);
or U47753 (N_47753,N_32925,N_38231);
and U47754 (N_47754,N_34620,N_30999);
nor U47755 (N_47755,N_30165,N_32514);
xnor U47756 (N_47756,N_39889,N_34638);
and U47757 (N_47757,N_39974,N_34873);
xnor U47758 (N_47758,N_32563,N_34183);
xnor U47759 (N_47759,N_35641,N_38023);
xnor U47760 (N_47760,N_34927,N_33001);
xor U47761 (N_47761,N_35382,N_39293);
and U47762 (N_47762,N_33953,N_38044);
or U47763 (N_47763,N_39348,N_32587);
or U47764 (N_47764,N_39539,N_31542);
or U47765 (N_47765,N_36448,N_39143);
nand U47766 (N_47766,N_38301,N_33532);
and U47767 (N_47767,N_35819,N_33466);
nand U47768 (N_47768,N_35109,N_30732);
nand U47769 (N_47769,N_32417,N_39735);
nor U47770 (N_47770,N_31858,N_38066);
nand U47771 (N_47771,N_33560,N_30348);
or U47772 (N_47772,N_37361,N_36243);
nand U47773 (N_47773,N_37191,N_38679);
and U47774 (N_47774,N_39931,N_39400);
and U47775 (N_47775,N_30487,N_30951);
xor U47776 (N_47776,N_36417,N_30049);
and U47777 (N_47777,N_39899,N_34509);
or U47778 (N_47778,N_31926,N_31265);
nand U47779 (N_47779,N_34342,N_31992);
or U47780 (N_47780,N_31897,N_38630);
nand U47781 (N_47781,N_30063,N_36945);
and U47782 (N_47782,N_30968,N_39145);
and U47783 (N_47783,N_37761,N_39928);
xnor U47784 (N_47784,N_33020,N_33066);
xnor U47785 (N_47785,N_32821,N_33037);
nor U47786 (N_47786,N_32713,N_37852);
nand U47787 (N_47787,N_32297,N_36364);
and U47788 (N_47788,N_38296,N_37649);
xor U47789 (N_47789,N_30130,N_35478);
nor U47790 (N_47790,N_38488,N_30242);
xnor U47791 (N_47791,N_39346,N_32235);
xnor U47792 (N_47792,N_31143,N_37813);
and U47793 (N_47793,N_37459,N_32760);
nor U47794 (N_47794,N_35130,N_34829);
xor U47795 (N_47795,N_35820,N_30045);
nor U47796 (N_47796,N_30929,N_30754);
or U47797 (N_47797,N_33092,N_36386);
nand U47798 (N_47798,N_34778,N_38724);
nand U47799 (N_47799,N_37545,N_31886);
or U47800 (N_47800,N_30054,N_30789);
xnor U47801 (N_47801,N_39246,N_31431);
xor U47802 (N_47802,N_30608,N_30721);
xor U47803 (N_47803,N_34100,N_36844);
nand U47804 (N_47804,N_34574,N_39312);
nand U47805 (N_47805,N_38770,N_37790);
or U47806 (N_47806,N_32507,N_32326);
and U47807 (N_47807,N_31515,N_39498);
or U47808 (N_47808,N_39375,N_30675);
or U47809 (N_47809,N_36001,N_39822);
nand U47810 (N_47810,N_30890,N_34522);
xnor U47811 (N_47811,N_36206,N_30783);
nand U47812 (N_47812,N_36926,N_30420);
or U47813 (N_47813,N_39431,N_37132);
or U47814 (N_47814,N_38376,N_30836);
nor U47815 (N_47815,N_31422,N_31300);
or U47816 (N_47816,N_35254,N_32203);
or U47817 (N_47817,N_37170,N_39987);
and U47818 (N_47818,N_31125,N_35401);
nor U47819 (N_47819,N_30820,N_33719);
and U47820 (N_47820,N_32628,N_31591);
and U47821 (N_47821,N_35246,N_38218);
nand U47822 (N_47822,N_37838,N_30009);
or U47823 (N_47823,N_38714,N_37721);
nand U47824 (N_47824,N_35678,N_34083);
xor U47825 (N_47825,N_35143,N_34297);
or U47826 (N_47826,N_33816,N_32583);
nor U47827 (N_47827,N_31755,N_32172);
or U47828 (N_47828,N_37320,N_38761);
nor U47829 (N_47829,N_38096,N_39466);
xnor U47830 (N_47830,N_31476,N_37323);
xnor U47831 (N_47831,N_37373,N_32146);
xor U47832 (N_47832,N_35200,N_36816);
nor U47833 (N_47833,N_31096,N_30416);
xnor U47834 (N_47834,N_36796,N_34936);
or U47835 (N_47835,N_32874,N_38186);
nor U47836 (N_47836,N_36162,N_34241);
or U47837 (N_47837,N_34073,N_32839);
or U47838 (N_47838,N_32893,N_31998);
or U47839 (N_47839,N_36978,N_33318);
or U47840 (N_47840,N_31704,N_39254);
nor U47841 (N_47841,N_39257,N_35253);
nor U47842 (N_47842,N_35611,N_31550);
and U47843 (N_47843,N_39337,N_38131);
xor U47844 (N_47844,N_35611,N_30186);
xnor U47845 (N_47845,N_39181,N_33892);
nand U47846 (N_47846,N_32998,N_38495);
or U47847 (N_47847,N_36636,N_32054);
xor U47848 (N_47848,N_36511,N_34978);
xor U47849 (N_47849,N_35815,N_39209);
nor U47850 (N_47850,N_30887,N_35727);
nor U47851 (N_47851,N_36451,N_38980);
nand U47852 (N_47852,N_30008,N_32832);
xor U47853 (N_47853,N_30432,N_35118);
and U47854 (N_47854,N_32920,N_39102);
xnor U47855 (N_47855,N_32061,N_33748);
and U47856 (N_47856,N_39888,N_30767);
xnor U47857 (N_47857,N_32964,N_39289);
nor U47858 (N_47858,N_32924,N_36507);
or U47859 (N_47859,N_31388,N_38329);
or U47860 (N_47860,N_35581,N_37738);
nand U47861 (N_47861,N_35449,N_30685);
xor U47862 (N_47862,N_39027,N_36660);
nand U47863 (N_47863,N_36419,N_34821);
and U47864 (N_47864,N_37508,N_31322);
xor U47865 (N_47865,N_34161,N_35690);
nand U47866 (N_47866,N_37370,N_39631);
xnor U47867 (N_47867,N_30714,N_31692);
nor U47868 (N_47868,N_36095,N_32303);
or U47869 (N_47869,N_34549,N_30371);
nor U47870 (N_47870,N_36809,N_33458);
and U47871 (N_47871,N_37316,N_31453);
nand U47872 (N_47872,N_33909,N_33062);
nor U47873 (N_47873,N_39689,N_38167);
nand U47874 (N_47874,N_37986,N_31932);
and U47875 (N_47875,N_31373,N_32059);
or U47876 (N_47876,N_30782,N_33970);
nand U47877 (N_47877,N_32037,N_36792);
and U47878 (N_47878,N_35838,N_39548);
nor U47879 (N_47879,N_33865,N_32035);
and U47880 (N_47880,N_30193,N_30799);
nand U47881 (N_47881,N_38440,N_35412);
and U47882 (N_47882,N_30083,N_31687);
nor U47883 (N_47883,N_33698,N_31031);
nand U47884 (N_47884,N_34776,N_31920);
or U47885 (N_47885,N_32353,N_36686);
xor U47886 (N_47886,N_31695,N_31426);
nor U47887 (N_47887,N_38044,N_32451);
or U47888 (N_47888,N_30707,N_33142);
and U47889 (N_47889,N_35923,N_37146);
xnor U47890 (N_47890,N_39144,N_38888);
nor U47891 (N_47891,N_35336,N_36274);
or U47892 (N_47892,N_38145,N_37621);
or U47893 (N_47893,N_30470,N_36986);
and U47894 (N_47894,N_34541,N_34844);
and U47895 (N_47895,N_34964,N_33502);
nand U47896 (N_47896,N_34313,N_31376);
xnor U47897 (N_47897,N_34525,N_36996);
nor U47898 (N_47898,N_32106,N_37665);
and U47899 (N_47899,N_31522,N_35225);
or U47900 (N_47900,N_31579,N_33070);
nor U47901 (N_47901,N_39232,N_31361);
and U47902 (N_47902,N_31816,N_32447);
nand U47903 (N_47903,N_39890,N_39321);
nand U47904 (N_47904,N_34760,N_36509);
or U47905 (N_47905,N_37237,N_33962);
and U47906 (N_47906,N_30987,N_31576);
nand U47907 (N_47907,N_33373,N_32755);
nand U47908 (N_47908,N_35742,N_37581);
nor U47909 (N_47909,N_38567,N_35076);
and U47910 (N_47910,N_30050,N_34328);
nor U47911 (N_47911,N_37613,N_37579);
xor U47912 (N_47912,N_31380,N_37681);
and U47913 (N_47913,N_35559,N_30651);
nor U47914 (N_47914,N_35863,N_32672);
and U47915 (N_47915,N_33857,N_33098);
and U47916 (N_47916,N_37675,N_33726);
xor U47917 (N_47917,N_39137,N_33852);
nor U47918 (N_47918,N_36293,N_32056);
nand U47919 (N_47919,N_37594,N_38383);
and U47920 (N_47920,N_38429,N_31011);
nor U47921 (N_47921,N_39755,N_36246);
xor U47922 (N_47922,N_36939,N_36940);
or U47923 (N_47923,N_35060,N_33835);
and U47924 (N_47924,N_39881,N_32532);
or U47925 (N_47925,N_38329,N_33986);
or U47926 (N_47926,N_34096,N_31642);
nand U47927 (N_47927,N_38844,N_34267);
or U47928 (N_47928,N_32884,N_31515);
or U47929 (N_47929,N_32800,N_31784);
nand U47930 (N_47930,N_31643,N_32367);
nor U47931 (N_47931,N_36053,N_32833);
nand U47932 (N_47932,N_32037,N_38241);
nor U47933 (N_47933,N_33348,N_35334);
xor U47934 (N_47934,N_35526,N_30017);
nor U47935 (N_47935,N_35009,N_31873);
nand U47936 (N_47936,N_32012,N_36087);
or U47937 (N_47937,N_37279,N_30269);
nor U47938 (N_47938,N_32648,N_30810);
xor U47939 (N_47939,N_36463,N_37415);
or U47940 (N_47940,N_39597,N_33912);
or U47941 (N_47941,N_33908,N_30764);
nand U47942 (N_47942,N_33077,N_33618);
nor U47943 (N_47943,N_33388,N_37861);
xnor U47944 (N_47944,N_35849,N_33966);
nor U47945 (N_47945,N_36197,N_36022);
nand U47946 (N_47946,N_31529,N_36954);
nand U47947 (N_47947,N_34202,N_37626);
and U47948 (N_47948,N_34781,N_39176);
nand U47949 (N_47949,N_37506,N_30253);
nand U47950 (N_47950,N_36761,N_35035);
or U47951 (N_47951,N_35055,N_33787);
nand U47952 (N_47952,N_30108,N_39540);
and U47953 (N_47953,N_34807,N_32014);
and U47954 (N_47954,N_33416,N_39398);
or U47955 (N_47955,N_36610,N_38256);
and U47956 (N_47956,N_30567,N_36916);
and U47957 (N_47957,N_34337,N_33964);
nand U47958 (N_47958,N_32350,N_36276);
nand U47959 (N_47959,N_39329,N_34989);
and U47960 (N_47960,N_39327,N_32891);
nor U47961 (N_47961,N_36092,N_31751);
nor U47962 (N_47962,N_31253,N_30471);
nand U47963 (N_47963,N_37051,N_39067);
nand U47964 (N_47964,N_30835,N_34420);
and U47965 (N_47965,N_37316,N_38352);
nor U47966 (N_47966,N_32453,N_38740);
and U47967 (N_47967,N_37625,N_33617);
and U47968 (N_47968,N_30183,N_39619);
or U47969 (N_47969,N_37695,N_34005);
nand U47970 (N_47970,N_33972,N_34661);
or U47971 (N_47971,N_33007,N_38231);
nor U47972 (N_47972,N_31710,N_34356);
nand U47973 (N_47973,N_36608,N_32834);
nor U47974 (N_47974,N_34162,N_30754);
nand U47975 (N_47975,N_31883,N_35871);
xor U47976 (N_47976,N_32866,N_33559);
and U47977 (N_47977,N_33748,N_39825);
and U47978 (N_47978,N_39996,N_33803);
xor U47979 (N_47979,N_37660,N_32643);
xor U47980 (N_47980,N_30002,N_33251);
nor U47981 (N_47981,N_32600,N_34273);
and U47982 (N_47982,N_30339,N_35058);
or U47983 (N_47983,N_37812,N_33428);
nand U47984 (N_47984,N_33505,N_33973);
nand U47985 (N_47985,N_36161,N_32343);
nand U47986 (N_47986,N_35448,N_35478);
xnor U47987 (N_47987,N_39521,N_33874);
nand U47988 (N_47988,N_38038,N_35182);
nor U47989 (N_47989,N_35066,N_34452);
or U47990 (N_47990,N_35005,N_36957);
nand U47991 (N_47991,N_33220,N_38208);
or U47992 (N_47992,N_35863,N_31548);
and U47993 (N_47993,N_35007,N_30463);
xnor U47994 (N_47994,N_37918,N_37892);
xnor U47995 (N_47995,N_37308,N_32932);
or U47996 (N_47996,N_38614,N_39575);
or U47997 (N_47997,N_32085,N_34384);
nor U47998 (N_47998,N_32390,N_33668);
and U47999 (N_47999,N_37358,N_31438);
xnor U48000 (N_48000,N_35039,N_36993);
nand U48001 (N_48001,N_32172,N_39477);
nand U48002 (N_48002,N_38852,N_31809);
and U48003 (N_48003,N_38738,N_39460);
nand U48004 (N_48004,N_38770,N_38567);
and U48005 (N_48005,N_31824,N_36067);
or U48006 (N_48006,N_36903,N_30980);
and U48007 (N_48007,N_34740,N_32523);
nor U48008 (N_48008,N_30347,N_34464);
nor U48009 (N_48009,N_38539,N_35304);
nand U48010 (N_48010,N_30807,N_39872);
nand U48011 (N_48011,N_34905,N_37513);
nand U48012 (N_48012,N_34011,N_32193);
or U48013 (N_48013,N_39969,N_39927);
and U48014 (N_48014,N_30116,N_37077);
nand U48015 (N_48015,N_37046,N_37277);
nor U48016 (N_48016,N_37564,N_35897);
xnor U48017 (N_48017,N_37896,N_30390);
xor U48018 (N_48018,N_32203,N_39385);
nor U48019 (N_48019,N_39373,N_30866);
nand U48020 (N_48020,N_37150,N_31782);
nor U48021 (N_48021,N_36768,N_30972);
nor U48022 (N_48022,N_37219,N_38483);
or U48023 (N_48023,N_35095,N_30333);
nor U48024 (N_48024,N_38814,N_36525);
nand U48025 (N_48025,N_34777,N_30953);
nor U48026 (N_48026,N_38207,N_39260);
and U48027 (N_48027,N_39485,N_32723);
and U48028 (N_48028,N_37958,N_34960);
nor U48029 (N_48029,N_39675,N_34582);
or U48030 (N_48030,N_35919,N_32164);
and U48031 (N_48031,N_36651,N_37325);
nor U48032 (N_48032,N_33114,N_32928);
xor U48033 (N_48033,N_30537,N_33180);
nor U48034 (N_48034,N_34191,N_39066);
and U48035 (N_48035,N_39549,N_33763);
nand U48036 (N_48036,N_39372,N_31042);
nand U48037 (N_48037,N_35381,N_38962);
nand U48038 (N_48038,N_34826,N_39355);
xnor U48039 (N_48039,N_35232,N_30466);
and U48040 (N_48040,N_32128,N_36074);
and U48041 (N_48041,N_32049,N_38572);
nand U48042 (N_48042,N_35982,N_39278);
nand U48043 (N_48043,N_35581,N_34333);
nand U48044 (N_48044,N_34444,N_38805);
and U48045 (N_48045,N_39505,N_39111);
or U48046 (N_48046,N_38796,N_39379);
xnor U48047 (N_48047,N_30207,N_36363);
nand U48048 (N_48048,N_37069,N_38441);
or U48049 (N_48049,N_36680,N_38439);
or U48050 (N_48050,N_32533,N_39788);
and U48051 (N_48051,N_36906,N_38616);
nor U48052 (N_48052,N_39072,N_31276);
and U48053 (N_48053,N_36535,N_35925);
nand U48054 (N_48054,N_38917,N_39536);
nand U48055 (N_48055,N_38480,N_34853);
or U48056 (N_48056,N_37979,N_31400);
and U48057 (N_48057,N_37092,N_35235);
or U48058 (N_48058,N_30227,N_37522);
xnor U48059 (N_48059,N_39082,N_32363);
and U48060 (N_48060,N_34388,N_32178);
nor U48061 (N_48061,N_30808,N_37383);
nor U48062 (N_48062,N_36210,N_33531);
and U48063 (N_48063,N_31829,N_33331);
and U48064 (N_48064,N_37685,N_31801);
nor U48065 (N_48065,N_35444,N_32610);
and U48066 (N_48066,N_31852,N_36623);
nand U48067 (N_48067,N_37644,N_36576);
nor U48068 (N_48068,N_35187,N_30474);
nor U48069 (N_48069,N_36427,N_35075);
xnor U48070 (N_48070,N_38314,N_32487);
and U48071 (N_48071,N_33161,N_31213);
nand U48072 (N_48072,N_37318,N_34045);
and U48073 (N_48073,N_32556,N_30762);
and U48074 (N_48074,N_32722,N_37670);
and U48075 (N_48075,N_39542,N_33690);
xor U48076 (N_48076,N_33714,N_34312);
nand U48077 (N_48077,N_37704,N_37435);
and U48078 (N_48078,N_39881,N_32702);
or U48079 (N_48079,N_30676,N_31768);
nand U48080 (N_48080,N_31085,N_36257);
nand U48081 (N_48081,N_30596,N_31106);
or U48082 (N_48082,N_35051,N_38894);
nor U48083 (N_48083,N_32149,N_39354);
and U48084 (N_48084,N_31941,N_33457);
and U48085 (N_48085,N_33831,N_30742);
and U48086 (N_48086,N_34400,N_36738);
xor U48087 (N_48087,N_35457,N_31822);
nand U48088 (N_48088,N_34323,N_32618);
nor U48089 (N_48089,N_30372,N_34246);
and U48090 (N_48090,N_36403,N_30208);
or U48091 (N_48091,N_37505,N_35791);
or U48092 (N_48092,N_38821,N_35513);
nand U48093 (N_48093,N_31632,N_33154);
xor U48094 (N_48094,N_31383,N_31534);
and U48095 (N_48095,N_38666,N_30747);
or U48096 (N_48096,N_39956,N_34671);
nand U48097 (N_48097,N_34479,N_37823);
xnor U48098 (N_48098,N_34688,N_39952);
nor U48099 (N_48099,N_33467,N_37633);
nand U48100 (N_48100,N_37835,N_36328);
nand U48101 (N_48101,N_39409,N_32989);
or U48102 (N_48102,N_36649,N_35050);
or U48103 (N_48103,N_37749,N_30020);
xnor U48104 (N_48104,N_35086,N_39788);
nand U48105 (N_48105,N_31249,N_38225);
and U48106 (N_48106,N_37456,N_33178);
nor U48107 (N_48107,N_34386,N_31164);
or U48108 (N_48108,N_32412,N_37750);
nand U48109 (N_48109,N_33542,N_38060);
and U48110 (N_48110,N_38185,N_32580);
or U48111 (N_48111,N_32836,N_37158);
and U48112 (N_48112,N_35029,N_31313);
and U48113 (N_48113,N_32686,N_32938);
or U48114 (N_48114,N_35473,N_30517);
xor U48115 (N_48115,N_33470,N_39540);
or U48116 (N_48116,N_35348,N_36076);
nor U48117 (N_48117,N_38397,N_36605);
xor U48118 (N_48118,N_31371,N_38328);
nand U48119 (N_48119,N_37015,N_31949);
and U48120 (N_48120,N_31033,N_39242);
or U48121 (N_48121,N_35655,N_34219);
xnor U48122 (N_48122,N_33308,N_36794);
and U48123 (N_48123,N_31815,N_30638);
xor U48124 (N_48124,N_36480,N_36774);
or U48125 (N_48125,N_38735,N_33332);
nor U48126 (N_48126,N_32944,N_39865);
nor U48127 (N_48127,N_38607,N_38648);
xnor U48128 (N_48128,N_34807,N_32582);
nor U48129 (N_48129,N_39400,N_39675);
xor U48130 (N_48130,N_37960,N_36584);
nor U48131 (N_48131,N_36223,N_31350);
or U48132 (N_48132,N_31342,N_34557);
and U48133 (N_48133,N_30073,N_38898);
nor U48134 (N_48134,N_37753,N_30397);
xor U48135 (N_48135,N_32093,N_39958);
and U48136 (N_48136,N_39958,N_39927);
and U48137 (N_48137,N_37493,N_38771);
nand U48138 (N_48138,N_37500,N_31131);
nand U48139 (N_48139,N_32515,N_37416);
xnor U48140 (N_48140,N_38178,N_37771);
and U48141 (N_48141,N_36795,N_32319);
nor U48142 (N_48142,N_39378,N_37794);
and U48143 (N_48143,N_30913,N_36261);
and U48144 (N_48144,N_32368,N_31902);
xor U48145 (N_48145,N_38767,N_31631);
or U48146 (N_48146,N_33329,N_39514);
xnor U48147 (N_48147,N_37327,N_36360);
nor U48148 (N_48148,N_38116,N_31571);
and U48149 (N_48149,N_34384,N_39910);
nor U48150 (N_48150,N_33203,N_31309);
nand U48151 (N_48151,N_38773,N_33885);
xnor U48152 (N_48152,N_30559,N_30279);
or U48153 (N_48153,N_37359,N_30827);
nand U48154 (N_48154,N_36840,N_31529);
or U48155 (N_48155,N_31461,N_32320);
and U48156 (N_48156,N_33008,N_39715);
and U48157 (N_48157,N_37533,N_32924);
nand U48158 (N_48158,N_33490,N_38693);
and U48159 (N_48159,N_35870,N_37469);
nor U48160 (N_48160,N_31048,N_39265);
nand U48161 (N_48161,N_36015,N_31927);
or U48162 (N_48162,N_38612,N_34993);
xnor U48163 (N_48163,N_36963,N_32222);
nand U48164 (N_48164,N_34015,N_39821);
and U48165 (N_48165,N_34592,N_33251);
or U48166 (N_48166,N_38274,N_30852);
nor U48167 (N_48167,N_35558,N_31493);
nor U48168 (N_48168,N_38268,N_31809);
and U48169 (N_48169,N_32120,N_39786);
nand U48170 (N_48170,N_33845,N_39431);
nor U48171 (N_48171,N_30914,N_39744);
nor U48172 (N_48172,N_34195,N_31561);
xnor U48173 (N_48173,N_39814,N_30457);
nand U48174 (N_48174,N_33576,N_39915);
nor U48175 (N_48175,N_39965,N_31591);
and U48176 (N_48176,N_37055,N_30578);
xor U48177 (N_48177,N_32784,N_37999);
nand U48178 (N_48178,N_33265,N_34466);
xnor U48179 (N_48179,N_34344,N_37188);
nor U48180 (N_48180,N_37125,N_35005);
or U48181 (N_48181,N_34832,N_36818);
or U48182 (N_48182,N_36361,N_38638);
nor U48183 (N_48183,N_37453,N_35532);
or U48184 (N_48184,N_34938,N_34399);
or U48185 (N_48185,N_32250,N_37515);
nand U48186 (N_48186,N_32523,N_34262);
xor U48187 (N_48187,N_30312,N_38081);
nor U48188 (N_48188,N_31805,N_35848);
nand U48189 (N_48189,N_32766,N_39306);
nand U48190 (N_48190,N_32455,N_30559);
xnor U48191 (N_48191,N_39355,N_36309);
nor U48192 (N_48192,N_33416,N_31307);
nand U48193 (N_48193,N_31040,N_33571);
nand U48194 (N_48194,N_35043,N_31803);
nor U48195 (N_48195,N_32012,N_32851);
or U48196 (N_48196,N_37105,N_35823);
nor U48197 (N_48197,N_34533,N_32626);
xor U48198 (N_48198,N_33824,N_35042);
nand U48199 (N_48199,N_36327,N_32294);
nor U48200 (N_48200,N_32045,N_39794);
nand U48201 (N_48201,N_36840,N_35451);
and U48202 (N_48202,N_34606,N_35987);
nand U48203 (N_48203,N_30444,N_34069);
xnor U48204 (N_48204,N_35019,N_34473);
and U48205 (N_48205,N_36774,N_39034);
or U48206 (N_48206,N_39025,N_38243);
or U48207 (N_48207,N_38917,N_35253);
and U48208 (N_48208,N_37639,N_37412);
and U48209 (N_48209,N_38309,N_36543);
or U48210 (N_48210,N_30179,N_36320);
xor U48211 (N_48211,N_36169,N_34275);
nand U48212 (N_48212,N_32074,N_35781);
xnor U48213 (N_48213,N_33128,N_32543);
and U48214 (N_48214,N_34626,N_34878);
nand U48215 (N_48215,N_38528,N_33172);
or U48216 (N_48216,N_30958,N_36051);
or U48217 (N_48217,N_38678,N_37167);
and U48218 (N_48218,N_30687,N_35888);
nand U48219 (N_48219,N_30751,N_35571);
and U48220 (N_48220,N_33547,N_38278);
nand U48221 (N_48221,N_36906,N_39244);
xnor U48222 (N_48222,N_34685,N_30755);
xor U48223 (N_48223,N_30236,N_31399);
nor U48224 (N_48224,N_30920,N_36024);
nor U48225 (N_48225,N_30284,N_31562);
xor U48226 (N_48226,N_31467,N_39196);
xor U48227 (N_48227,N_31616,N_33563);
nand U48228 (N_48228,N_34994,N_35607);
or U48229 (N_48229,N_35201,N_39541);
nand U48230 (N_48230,N_31384,N_31572);
nor U48231 (N_48231,N_34174,N_34962);
nand U48232 (N_48232,N_31528,N_37376);
and U48233 (N_48233,N_34454,N_30652);
nand U48234 (N_48234,N_39284,N_34040);
and U48235 (N_48235,N_32399,N_36692);
or U48236 (N_48236,N_35011,N_38830);
or U48237 (N_48237,N_38434,N_39189);
or U48238 (N_48238,N_31629,N_38595);
xnor U48239 (N_48239,N_34087,N_33387);
nor U48240 (N_48240,N_34261,N_37424);
and U48241 (N_48241,N_30482,N_33647);
nand U48242 (N_48242,N_33533,N_37839);
xnor U48243 (N_48243,N_31092,N_33445);
nor U48244 (N_48244,N_39371,N_35148);
xnor U48245 (N_48245,N_36439,N_39693);
or U48246 (N_48246,N_32056,N_39265);
and U48247 (N_48247,N_33313,N_32599);
xor U48248 (N_48248,N_33860,N_32569);
nand U48249 (N_48249,N_31576,N_31436);
xor U48250 (N_48250,N_31478,N_32694);
nand U48251 (N_48251,N_39872,N_35411);
xnor U48252 (N_48252,N_39145,N_33758);
xor U48253 (N_48253,N_30330,N_39656);
nor U48254 (N_48254,N_31469,N_36679);
nor U48255 (N_48255,N_33406,N_32393);
nand U48256 (N_48256,N_35175,N_39242);
nand U48257 (N_48257,N_31087,N_33113);
xor U48258 (N_48258,N_37308,N_37933);
nor U48259 (N_48259,N_36424,N_34679);
nand U48260 (N_48260,N_34236,N_37042);
xnor U48261 (N_48261,N_31007,N_39129);
or U48262 (N_48262,N_31688,N_31878);
or U48263 (N_48263,N_37863,N_35599);
and U48264 (N_48264,N_39069,N_39009);
nor U48265 (N_48265,N_31034,N_38424);
and U48266 (N_48266,N_38516,N_38999);
nand U48267 (N_48267,N_33866,N_34725);
nand U48268 (N_48268,N_39190,N_30351);
xnor U48269 (N_48269,N_33456,N_32775);
xor U48270 (N_48270,N_35668,N_31529);
nand U48271 (N_48271,N_37596,N_32736);
nor U48272 (N_48272,N_30054,N_36989);
xor U48273 (N_48273,N_36584,N_31710);
and U48274 (N_48274,N_32574,N_36574);
or U48275 (N_48275,N_37337,N_32820);
xor U48276 (N_48276,N_30638,N_30735);
nor U48277 (N_48277,N_37669,N_36143);
xor U48278 (N_48278,N_32635,N_32613);
nand U48279 (N_48279,N_32390,N_34795);
or U48280 (N_48280,N_39986,N_35292);
or U48281 (N_48281,N_32260,N_39161);
nor U48282 (N_48282,N_31562,N_38770);
xnor U48283 (N_48283,N_30509,N_38697);
or U48284 (N_48284,N_33771,N_34741);
or U48285 (N_48285,N_34793,N_32106);
xnor U48286 (N_48286,N_39646,N_32820);
and U48287 (N_48287,N_37041,N_37655);
nand U48288 (N_48288,N_39130,N_31625);
nor U48289 (N_48289,N_33693,N_31051);
nor U48290 (N_48290,N_39420,N_36776);
or U48291 (N_48291,N_30281,N_31406);
nand U48292 (N_48292,N_39652,N_35530);
xor U48293 (N_48293,N_30626,N_32783);
nand U48294 (N_48294,N_31648,N_39857);
and U48295 (N_48295,N_36645,N_39860);
nand U48296 (N_48296,N_38135,N_31349);
nor U48297 (N_48297,N_31241,N_38866);
nor U48298 (N_48298,N_32264,N_31793);
nor U48299 (N_48299,N_31197,N_30691);
xnor U48300 (N_48300,N_39783,N_31951);
nand U48301 (N_48301,N_30260,N_32397);
and U48302 (N_48302,N_39091,N_30421);
nor U48303 (N_48303,N_33844,N_32055);
or U48304 (N_48304,N_33546,N_30878);
or U48305 (N_48305,N_38268,N_32536);
or U48306 (N_48306,N_36709,N_34374);
nor U48307 (N_48307,N_33284,N_38201);
nor U48308 (N_48308,N_38995,N_38053);
xnor U48309 (N_48309,N_34256,N_36311);
xor U48310 (N_48310,N_33212,N_32726);
nor U48311 (N_48311,N_39460,N_38060);
nor U48312 (N_48312,N_31013,N_36664);
nor U48313 (N_48313,N_37068,N_39817);
nor U48314 (N_48314,N_36660,N_35541);
or U48315 (N_48315,N_37256,N_37302);
or U48316 (N_48316,N_31327,N_38125);
or U48317 (N_48317,N_33602,N_38780);
or U48318 (N_48318,N_34144,N_33514);
xor U48319 (N_48319,N_30772,N_34631);
or U48320 (N_48320,N_33468,N_31165);
nand U48321 (N_48321,N_34103,N_35352);
xnor U48322 (N_48322,N_31335,N_30880);
or U48323 (N_48323,N_31879,N_36165);
nor U48324 (N_48324,N_34164,N_33508);
nand U48325 (N_48325,N_30997,N_31531);
xor U48326 (N_48326,N_37463,N_30434);
or U48327 (N_48327,N_36367,N_34016);
and U48328 (N_48328,N_32827,N_32159);
nand U48329 (N_48329,N_37394,N_30639);
and U48330 (N_48330,N_33907,N_31265);
or U48331 (N_48331,N_30759,N_34695);
or U48332 (N_48332,N_36660,N_33088);
or U48333 (N_48333,N_30848,N_39719);
nor U48334 (N_48334,N_38809,N_39512);
or U48335 (N_48335,N_33541,N_37593);
or U48336 (N_48336,N_39502,N_30939);
or U48337 (N_48337,N_38101,N_39191);
and U48338 (N_48338,N_39742,N_37442);
nor U48339 (N_48339,N_37197,N_35311);
nand U48340 (N_48340,N_35512,N_38358);
and U48341 (N_48341,N_30381,N_33676);
nor U48342 (N_48342,N_33283,N_38758);
nand U48343 (N_48343,N_35839,N_37505);
or U48344 (N_48344,N_35957,N_31727);
and U48345 (N_48345,N_32561,N_36891);
nor U48346 (N_48346,N_37807,N_35509);
nor U48347 (N_48347,N_35659,N_35196);
and U48348 (N_48348,N_38447,N_32292);
xnor U48349 (N_48349,N_35833,N_35029);
and U48350 (N_48350,N_36972,N_30356);
xnor U48351 (N_48351,N_37015,N_30958);
nor U48352 (N_48352,N_39985,N_34547);
or U48353 (N_48353,N_35087,N_35177);
nor U48354 (N_48354,N_36331,N_36539);
or U48355 (N_48355,N_36908,N_37585);
nor U48356 (N_48356,N_33449,N_33162);
or U48357 (N_48357,N_39718,N_33283);
xnor U48358 (N_48358,N_37238,N_32577);
or U48359 (N_48359,N_34335,N_37471);
xnor U48360 (N_48360,N_36290,N_36112);
nand U48361 (N_48361,N_37297,N_33949);
nor U48362 (N_48362,N_39747,N_38561);
nand U48363 (N_48363,N_32333,N_37352);
xnor U48364 (N_48364,N_39660,N_32161);
nand U48365 (N_48365,N_34462,N_30584);
and U48366 (N_48366,N_35516,N_30722);
or U48367 (N_48367,N_32623,N_32728);
or U48368 (N_48368,N_39703,N_35388);
nor U48369 (N_48369,N_39834,N_33376);
nand U48370 (N_48370,N_35821,N_39303);
nand U48371 (N_48371,N_36143,N_33945);
nor U48372 (N_48372,N_38943,N_34926);
xnor U48373 (N_48373,N_38221,N_38075);
nor U48374 (N_48374,N_38776,N_32951);
and U48375 (N_48375,N_33780,N_31239);
xor U48376 (N_48376,N_34604,N_35493);
nor U48377 (N_48377,N_31244,N_30379);
nand U48378 (N_48378,N_35658,N_37739);
xnor U48379 (N_48379,N_31278,N_33081);
or U48380 (N_48380,N_31174,N_32690);
xor U48381 (N_48381,N_30776,N_32950);
nor U48382 (N_48382,N_39526,N_33393);
or U48383 (N_48383,N_34861,N_31388);
nand U48384 (N_48384,N_33201,N_31511);
and U48385 (N_48385,N_34132,N_33887);
xnor U48386 (N_48386,N_34338,N_35457);
xor U48387 (N_48387,N_31561,N_32947);
nor U48388 (N_48388,N_39677,N_30594);
nand U48389 (N_48389,N_38443,N_32239);
xor U48390 (N_48390,N_39017,N_35179);
xor U48391 (N_48391,N_30026,N_38847);
nor U48392 (N_48392,N_33201,N_35470);
nand U48393 (N_48393,N_36128,N_39307);
nand U48394 (N_48394,N_34711,N_30977);
xor U48395 (N_48395,N_35294,N_33118);
nor U48396 (N_48396,N_35821,N_31533);
and U48397 (N_48397,N_32094,N_35495);
nand U48398 (N_48398,N_34690,N_35124);
and U48399 (N_48399,N_38362,N_33344);
nand U48400 (N_48400,N_32076,N_36549);
or U48401 (N_48401,N_38720,N_35382);
nor U48402 (N_48402,N_37908,N_36149);
nand U48403 (N_48403,N_33314,N_32848);
or U48404 (N_48404,N_37687,N_31580);
and U48405 (N_48405,N_32690,N_31427);
and U48406 (N_48406,N_36765,N_34614);
and U48407 (N_48407,N_36790,N_37163);
nand U48408 (N_48408,N_36907,N_30084);
nand U48409 (N_48409,N_30499,N_31710);
and U48410 (N_48410,N_33334,N_36483);
nand U48411 (N_48411,N_30962,N_33099);
and U48412 (N_48412,N_32633,N_32706);
nor U48413 (N_48413,N_33294,N_31370);
and U48414 (N_48414,N_36492,N_33169);
and U48415 (N_48415,N_32875,N_36052);
xnor U48416 (N_48416,N_39109,N_34580);
nand U48417 (N_48417,N_38660,N_35235);
and U48418 (N_48418,N_32477,N_37849);
or U48419 (N_48419,N_39230,N_34891);
nand U48420 (N_48420,N_33393,N_33613);
xnor U48421 (N_48421,N_39116,N_36535);
xor U48422 (N_48422,N_35494,N_38911);
nor U48423 (N_48423,N_37651,N_32553);
xnor U48424 (N_48424,N_34962,N_35135);
or U48425 (N_48425,N_38636,N_35631);
xor U48426 (N_48426,N_35303,N_37801);
and U48427 (N_48427,N_36898,N_32553);
or U48428 (N_48428,N_32095,N_32253);
and U48429 (N_48429,N_31611,N_33088);
or U48430 (N_48430,N_37836,N_35942);
nand U48431 (N_48431,N_35149,N_37515);
or U48432 (N_48432,N_39647,N_35690);
xnor U48433 (N_48433,N_31602,N_39393);
nor U48434 (N_48434,N_30982,N_30182);
and U48435 (N_48435,N_33977,N_33310);
and U48436 (N_48436,N_31541,N_33820);
or U48437 (N_48437,N_31402,N_33222);
nor U48438 (N_48438,N_33953,N_38687);
nor U48439 (N_48439,N_36774,N_34193);
xnor U48440 (N_48440,N_35001,N_30576);
nor U48441 (N_48441,N_37033,N_30456);
nand U48442 (N_48442,N_31493,N_33605);
nand U48443 (N_48443,N_39379,N_39480);
nand U48444 (N_48444,N_35014,N_33250);
nor U48445 (N_48445,N_37185,N_36537);
nand U48446 (N_48446,N_33714,N_36421);
or U48447 (N_48447,N_30801,N_36976);
xor U48448 (N_48448,N_37655,N_32864);
and U48449 (N_48449,N_34873,N_36496);
or U48450 (N_48450,N_34136,N_35693);
or U48451 (N_48451,N_36065,N_32088);
and U48452 (N_48452,N_36297,N_39631);
xnor U48453 (N_48453,N_38476,N_33603);
or U48454 (N_48454,N_30401,N_30353);
or U48455 (N_48455,N_36055,N_31467);
or U48456 (N_48456,N_38548,N_31208);
nor U48457 (N_48457,N_30736,N_36932);
and U48458 (N_48458,N_36730,N_39304);
xnor U48459 (N_48459,N_30878,N_31513);
nand U48460 (N_48460,N_34363,N_34742);
xor U48461 (N_48461,N_37339,N_30724);
nand U48462 (N_48462,N_37325,N_39349);
nor U48463 (N_48463,N_33204,N_38496);
and U48464 (N_48464,N_33591,N_30167);
nor U48465 (N_48465,N_31037,N_36490);
nand U48466 (N_48466,N_37148,N_32739);
nand U48467 (N_48467,N_31479,N_34520);
nand U48468 (N_48468,N_35998,N_39831);
nor U48469 (N_48469,N_34007,N_39211);
and U48470 (N_48470,N_33778,N_36938);
nor U48471 (N_48471,N_35973,N_32072);
nand U48472 (N_48472,N_37238,N_39562);
nor U48473 (N_48473,N_33376,N_31703);
and U48474 (N_48474,N_30273,N_36882);
xor U48475 (N_48475,N_37765,N_30772);
and U48476 (N_48476,N_39959,N_34545);
or U48477 (N_48477,N_31112,N_33379);
xnor U48478 (N_48478,N_31631,N_39352);
nand U48479 (N_48479,N_37407,N_38405);
xnor U48480 (N_48480,N_34708,N_33605);
or U48481 (N_48481,N_30821,N_37106);
or U48482 (N_48482,N_34722,N_34063);
and U48483 (N_48483,N_35259,N_36928);
or U48484 (N_48484,N_39349,N_35388);
xnor U48485 (N_48485,N_32698,N_34612);
nor U48486 (N_48486,N_30685,N_36679);
and U48487 (N_48487,N_34245,N_38304);
xor U48488 (N_48488,N_37008,N_31535);
or U48489 (N_48489,N_39822,N_36388);
nand U48490 (N_48490,N_39348,N_37213);
nand U48491 (N_48491,N_31198,N_33877);
or U48492 (N_48492,N_35974,N_36663);
xnor U48493 (N_48493,N_31481,N_35002);
or U48494 (N_48494,N_38676,N_32998);
nor U48495 (N_48495,N_35658,N_38319);
xor U48496 (N_48496,N_33149,N_35992);
nor U48497 (N_48497,N_34562,N_39436);
nor U48498 (N_48498,N_34294,N_36823);
and U48499 (N_48499,N_38679,N_32641);
and U48500 (N_48500,N_30084,N_30730);
xnor U48501 (N_48501,N_39313,N_39778);
or U48502 (N_48502,N_34109,N_34833);
nand U48503 (N_48503,N_36878,N_30504);
nand U48504 (N_48504,N_35541,N_31787);
nor U48505 (N_48505,N_38811,N_31263);
and U48506 (N_48506,N_32928,N_37163);
nor U48507 (N_48507,N_35212,N_38658);
nand U48508 (N_48508,N_34437,N_36211);
and U48509 (N_48509,N_31314,N_39215);
and U48510 (N_48510,N_36963,N_31461);
xnor U48511 (N_48511,N_38199,N_38957);
xor U48512 (N_48512,N_34288,N_31117);
and U48513 (N_48513,N_35000,N_33752);
nand U48514 (N_48514,N_36910,N_37062);
nand U48515 (N_48515,N_38244,N_34109);
or U48516 (N_48516,N_38984,N_33273);
and U48517 (N_48517,N_30757,N_35233);
and U48518 (N_48518,N_34004,N_35069);
xnor U48519 (N_48519,N_36122,N_39032);
nand U48520 (N_48520,N_38110,N_38035);
nor U48521 (N_48521,N_36481,N_34617);
nand U48522 (N_48522,N_35795,N_37654);
nand U48523 (N_48523,N_37870,N_35380);
nor U48524 (N_48524,N_34682,N_34121);
nor U48525 (N_48525,N_36044,N_35697);
xnor U48526 (N_48526,N_35959,N_37324);
nand U48527 (N_48527,N_39422,N_30252);
and U48528 (N_48528,N_32871,N_38326);
and U48529 (N_48529,N_37698,N_32211);
and U48530 (N_48530,N_36234,N_36859);
or U48531 (N_48531,N_31300,N_35470);
nand U48532 (N_48532,N_37285,N_33843);
nand U48533 (N_48533,N_33565,N_37349);
nor U48534 (N_48534,N_33919,N_39942);
or U48535 (N_48535,N_35232,N_36337);
xor U48536 (N_48536,N_34599,N_39604);
nand U48537 (N_48537,N_31101,N_34271);
nand U48538 (N_48538,N_34536,N_36773);
and U48539 (N_48539,N_33790,N_30756);
and U48540 (N_48540,N_35323,N_39642);
or U48541 (N_48541,N_36107,N_31647);
nor U48542 (N_48542,N_36261,N_36949);
and U48543 (N_48543,N_39893,N_32536);
nand U48544 (N_48544,N_38557,N_31096);
xor U48545 (N_48545,N_39891,N_35787);
nand U48546 (N_48546,N_32398,N_36108);
nor U48547 (N_48547,N_32888,N_30824);
xnor U48548 (N_48548,N_31816,N_34628);
nand U48549 (N_48549,N_39895,N_31428);
nand U48550 (N_48550,N_32352,N_30391);
nand U48551 (N_48551,N_33848,N_36620);
nand U48552 (N_48552,N_34819,N_39165);
or U48553 (N_48553,N_35961,N_38887);
nand U48554 (N_48554,N_34126,N_32544);
xnor U48555 (N_48555,N_30207,N_35860);
nor U48556 (N_48556,N_36245,N_36799);
xor U48557 (N_48557,N_31635,N_35666);
nand U48558 (N_48558,N_38719,N_35169);
nand U48559 (N_48559,N_36021,N_38096);
nand U48560 (N_48560,N_38749,N_31056);
nand U48561 (N_48561,N_30614,N_36086);
nor U48562 (N_48562,N_37032,N_39821);
nor U48563 (N_48563,N_37609,N_38509);
xnor U48564 (N_48564,N_39817,N_37785);
nand U48565 (N_48565,N_35195,N_30995);
nand U48566 (N_48566,N_31263,N_36431);
nand U48567 (N_48567,N_33725,N_33575);
and U48568 (N_48568,N_38734,N_32585);
and U48569 (N_48569,N_31598,N_31386);
and U48570 (N_48570,N_39774,N_31520);
nor U48571 (N_48571,N_36620,N_33361);
nor U48572 (N_48572,N_31311,N_39671);
nor U48573 (N_48573,N_33749,N_34889);
nor U48574 (N_48574,N_34110,N_37481);
xor U48575 (N_48575,N_38232,N_39605);
nor U48576 (N_48576,N_35300,N_30880);
or U48577 (N_48577,N_31611,N_39105);
xor U48578 (N_48578,N_32441,N_31741);
nor U48579 (N_48579,N_32177,N_30946);
nor U48580 (N_48580,N_37426,N_39132);
xnor U48581 (N_48581,N_37172,N_36879);
xnor U48582 (N_48582,N_31586,N_38918);
and U48583 (N_48583,N_37547,N_36302);
nand U48584 (N_48584,N_34338,N_30014);
and U48585 (N_48585,N_32773,N_37096);
xnor U48586 (N_48586,N_37466,N_31366);
xor U48587 (N_48587,N_36270,N_32596);
or U48588 (N_48588,N_38270,N_36019);
and U48589 (N_48589,N_35254,N_37692);
nand U48590 (N_48590,N_32873,N_31103);
or U48591 (N_48591,N_36482,N_34684);
and U48592 (N_48592,N_32296,N_32676);
and U48593 (N_48593,N_35716,N_32913);
and U48594 (N_48594,N_37268,N_37914);
or U48595 (N_48595,N_30000,N_39925);
or U48596 (N_48596,N_32426,N_30189);
nand U48597 (N_48597,N_37530,N_36240);
nor U48598 (N_48598,N_39887,N_30177);
and U48599 (N_48599,N_35427,N_39219);
or U48600 (N_48600,N_38919,N_38415);
nand U48601 (N_48601,N_37217,N_39441);
xor U48602 (N_48602,N_31424,N_39522);
or U48603 (N_48603,N_30776,N_37006);
and U48604 (N_48604,N_35485,N_32064);
and U48605 (N_48605,N_31765,N_33439);
nor U48606 (N_48606,N_36231,N_34088);
or U48607 (N_48607,N_36465,N_37976);
or U48608 (N_48608,N_39980,N_36303);
nor U48609 (N_48609,N_39394,N_38879);
and U48610 (N_48610,N_32333,N_33141);
and U48611 (N_48611,N_39446,N_34422);
nor U48612 (N_48612,N_32874,N_39197);
nand U48613 (N_48613,N_38625,N_30642);
xor U48614 (N_48614,N_37451,N_31180);
and U48615 (N_48615,N_34088,N_33446);
nor U48616 (N_48616,N_35097,N_39184);
xor U48617 (N_48617,N_33919,N_38742);
nand U48618 (N_48618,N_36527,N_39961);
nor U48619 (N_48619,N_35262,N_36154);
or U48620 (N_48620,N_36362,N_37278);
nor U48621 (N_48621,N_35070,N_39830);
nor U48622 (N_48622,N_31061,N_39662);
xnor U48623 (N_48623,N_39423,N_38233);
nor U48624 (N_48624,N_32243,N_30285);
or U48625 (N_48625,N_33351,N_30894);
and U48626 (N_48626,N_35899,N_35411);
and U48627 (N_48627,N_33342,N_30106);
xnor U48628 (N_48628,N_31974,N_38625);
or U48629 (N_48629,N_38024,N_36670);
nor U48630 (N_48630,N_36505,N_36185);
nor U48631 (N_48631,N_36086,N_38276);
nor U48632 (N_48632,N_37952,N_35602);
nor U48633 (N_48633,N_30385,N_34173);
or U48634 (N_48634,N_39765,N_32848);
xnor U48635 (N_48635,N_30248,N_31469);
and U48636 (N_48636,N_33608,N_36466);
or U48637 (N_48637,N_30282,N_38952);
or U48638 (N_48638,N_30493,N_35009);
or U48639 (N_48639,N_31605,N_30242);
nand U48640 (N_48640,N_35529,N_31398);
xor U48641 (N_48641,N_33264,N_31032);
and U48642 (N_48642,N_31172,N_38077);
or U48643 (N_48643,N_35508,N_31691);
nor U48644 (N_48644,N_36820,N_39891);
nand U48645 (N_48645,N_32283,N_34217);
nor U48646 (N_48646,N_34770,N_38447);
or U48647 (N_48647,N_34810,N_30093);
nand U48648 (N_48648,N_31617,N_31583);
or U48649 (N_48649,N_31265,N_35160);
or U48650 (N_48650,N_32491,N_37094);
and U48651 (N_48651,N_32240,N_33859);
nor U48652 (N_48652,N_36263,N_36122);
nand U48653 (N_48653,N_37640,N_32980);
xnor U48654 (N_48654,N_38765,N_39009);
xnor U48655 (N_48655,N_38092,N_31435);
or U48656 (N_48656,N_38022,N_34347);
xor U48657 (N_48657,N_34881,N_37716);
xnor U48658 (N_48658,N_38518,N_31790);
xor U48659 (N_48659,N_39639,N_32935);
xor U48660 (N_48660,N_33963,N_30526);
nand U48661 (N_48661,N_31482,N_33444);
and U48662 (N_48662,N_34757,N_35902);
or U48663 (N_48663,N_34409,N_33270);
nor U48664 (N_48664,N_33642,N_33379);
or U48665 (N_48665,N_32751,N_35300);
and U48666 (N_48666,N_35584,N_30473);
xnor U48667 (N_48667,N_30679,N_37965);
nand U48668 (N_48668,N_32096,N_39994);
xnor U48669 (N_48669,N_31014,N_39470);
nand U48670 (N_48670,N_30971,N_38226);
nand U48671 (N_48671,N_36720,N_39564);
xor U48672 (N_48672,N_37049,N_38514);
nor U48673 (N_48673,N_35035,N_30382);
nand U48674 (N_48674,N_38018,N_30519);
nor U48675 (N_48675,N_38983,N_39056);
nor U48676 (N_48676,N_33178,N_37812);
and U48677 (N_48677,N_31767,N_30830);
nor U48678 (N_48678,N_32277,N_33588);
nand U48679 (N_48679,N_38500,N_38705);
nand U48680 (N_48680,N_31033,N_30667);
nor U48681 (N_48681,N_32772,N_34385);
nand U48682 (N_48682,N_31102,N_37243);
nor U48683 (N_48683,N_38498,N_34819);
or U48684 (N_48684,N_32079,N_34179);
nand U48685 (N_48685,N_36905,N_35654);
and U48686 (N_48686,N_35135,N_35002);
nand U48687 (N_48687,N_35936,N_39472);
xnor U48688 (N_48688,N_31532,N_30856);
or U48689 (N_48689,N_37778,N_39708);
nor U48690 (N_48690,N_36875,N_38257);
and U48691 (N_48691,N_30812,N_35415);
or U48692 (N_48692,N_33213,N_32930);
or U48693 (N_48693,N_36674,N_32286);
or U48694 (N_48694,N_39411,N_34905);
or U48695 (N_48695,N_31757,N_35880);
or U48696 (N_48696,N_30763,N_31029);
or U48697 (N_48697,N_39280,N_31808);
nor U48698 (N_48698,N_33704,N_31578);
or U48699 (N_48699,N_30589,N_32849);
nor U48700 (N_48700,N_31400,N_39276);
nand U48701 (N_48701,N_35452,N_32106);
xor U48702 (N_48702,N_30263,N_30340);
and U48703 (N_48703,N_31729,N_34457);
or U48704 (N_48704,N_32267,N_37354);
or U48705 (N_48705,N_35780,N_36997);
nand U48706 (N_48706,N_31495,N_36216);
nand U48707 (N_48707,N_33030,N_39673);
xnor U48708 (N_48708,N_31070,N_32915);
and U48709 (N_48709,N_39930,N_33647);
or U48710 (N_48710,N_39220,N_33615);
nor U48711 (N_48711,N_39220,N_31206);
nor U48712 (N_48712,N_32980,N_35944);
nand U48713 (N_48713,N_30852,N_39970);
xor U48714 (N_48714,N_35363,N_39007);
or U48715 (N_48715,N_35741,N_35986);
and U48716 (N_48716,N_35687,N_38847);
and U48717 (N_48717,N_39527,N_39024);
xor U48718 (N_48718,N_39300,N_34795);
and U48719 (N_48719,N_31810,N_32880);
nand U48720 (N_48720,N_32674,N_36164);
nor U48721 (N_48721,N_35435,N_38878);
nand U48722 (N_48722,N_32794,N_37361);
xor U48723 (N_48723,N_36004,N_33990);
nand U48724 (N_48724,N_32086,N_33895);
nand U48725 (N_48725,N_32619,N_37586);
nand U48726 (N_48726,N_36839,N_36890);
and U48727 (N_48727,N_37157,N_36668);
nor U48728 (N_48728,N_38063,N_35392);
or U48729 (N_48729,N_37106,N_36030);
nor U48730 (N_48730,N_30973,N_34624);
and U48731 (N_48731,N_38291,N_30774);
xnor U48732 (N_48732,N_34496,N_37048);
and U48733 (N_48733,N_37119,N_35598);
xnor U48734 (N_48734,N_35829,N_36494);
nor U48735 (N_48735,N_36946,N_30024);
nand U48736 (N_48736,N_39051,N_32098);
xor U48737 (N_48737,N_33084,N_32911);
or U48738 (N_48738,N_31608,N_38162);
or U48739 (N_48739,N_37370,N_36365);
nor U48740 (N_48740,N_39109,N_38801);
xor U48741 (N_48741,N_35361,N_31974);
nor U48742 (N_48742,N_39281,N_33402);
nand U48743 (N_48743,N_34787,N_37567);
nand U48744 (N_48744,N_39635,N_36593);
xor U48745 (N_48745,N_35342,N_32139);
or U48746 (N_48746,N_35420,N_38471);
xor U48747 (N_48747,N_39251,N_34347);
or U48748 (N_48748,N_39736,N_37692);
nand U48749 (N_48749,N_33455,N_37914);
nor U48750 (N_48750,N_30162,N_36701);
xnor U48751 (N_48751,N_38556,N_39514);
or U48752 (N_48752,N_33386,N_33522);
nor U48753 (N_48753,N_39022,N_35367);
nand U48754 (N_48754,N_33505,N_30221);
nand U48755 (N_48755,N_35498,N_35154);
nor U48756 (N_48756,N_30912,N_35524);
nor U48757 (N_48757,N_39463,N_33562);
nand U48758 (N_48758,N_32665,N_31200);
nor U48759 (N_48759,N_38593,N_34013);
nor U48760 (N_48760,N_32782,N_30020);
nor U48761 (N_48761,N_32363,N_33815);
xnor U48762 (N_48762,N_38996,N_34675);
nor U48763 (N_48763,N_33803,N_34059);
xor U48764 (N_48764,N_35923,N_38109);
nor U48765 (N_48765,N_34226,N_37074);
nand U48766 (N_48766,N_33204,N_33072);
or U48767 (N_48767,N_37387,N_36489);
and U48768 (N_48768,N_39954,N_37001);
nand U48769 (N_48769,N_32624,N_39178);
or U48770 (N_48770,N_32381,N_38877);
nand U48771 (N_48771,N_33672,N_30988);
and U48772 (N_48772,N_31996,N_33866);
nor U48773 (N_48773,N_35938,N_30398);
nor U48774 (N_48774,N_36312,N_38959);
nand U48775 (N_48775,N_33413,N_37577);
or U48776 (N_48776,N_30702,N_39368);
and U48777 (N_48777,N_35866,N_34835);
xnor U48778 (N_48778,N_38735,N_37418);
nand U48779 (N_48779,N_34788,N_35088);
or U48780 (N_48780,N_37463,N_34186);
and U48781 (N_48781,N_30700,N_32285);
nor U48782 (N_48782,N_32399,N_38098);
nor U48783 (N_48783,N_35533,N_30586);
xnor U48784 (N_48784,N_32159,N_31743);
nand U48785 (N_48785,N_32860,N_38938);
nor U48786 (N_48786,N_38364,N_38652);
or U48787 (N_48787,N_33391,N_31140);
nor U48788 (N_48788,N_35864,N_36379);
nor U48789 (N_48789,N_35256,N_34246);
nor U48790 (N_48790,N_31881,N_36323);
and U48791 (N_48791,N_34391,N_30354);
and U48792 (N_48792,N_31403,N_36093);
nand U48793 (N_48793,N_33502,N_33997);
nand U48794 (N_48794,N_31383,N_31336);
and U48795 (N_48795,N_34997,N_34976);
xor U48796 (N_48796,N_30839,N_35734);
nand U48797 (N_48797,N_36266,N_39574);
and U48798 (N_48798,N_30092,N_34675);
and U48799 (N_48799,N_35680,N_31873);
and U48800 (N_48800,N_32140,N_31950);
and U48801 (N_48801,N_35250,N_39085);
nand U48802 (N_48802,N_35455,N_35718);
xnor U48803 (N_48803,N_36920,N_32977);
and U48804 (N_48804,N_30939,N_32979);
xor U48805 (N_48805,N_30943,N_36591);
nor U48806 (N_48806,N_39235,N_33886);
and U48807 (N_48807,N_33173,N_37796);
xor U48808 (N_48808,N_39242,N_33181);
or U48809 (N_48809,N_34864,N_37069);
or U48810 (N_48810,N_31923,N_38760);
xor U48811 (N_48811,N_32935,N_35985);
xor U48812 (N_48812,N_36503,N_38599);
and U48813 (N_48813,N_33818,N_37726);
xnor U48814 (N_48814,N_34681,N_31831);
nor U48815 (N_48815,N_35385,N_36038);
or U48816 (N_48816,N_38643,N_38950);
xor U48817 (N_48817,N_31514,N_37359);
nand U48818 (N_48818,N_33237,N_39835);
or U48819 (N_48819,N_31020,N_33116);
or U48820 (N_48820,N_36898,N_38629);
nor U48821 (N_48821,N_34312,N_38165);
xor U48822 (N_48822,N_37662,N_38307);
nor U48823 (N_48823,N_38903,N_31290);
nand U48824 (N_48824,N_30994,N_38731);
xor U48825 (N_48825,N_37475,N_32254);
xor U48826 (N_48826,N_39271,N_30164);
xor U48827 (N_48827,N_30177,N_37603);
xor U48828 (N_48828,N_32277,N_33468);
xor U48829 (N_48829,N_38923,N_35084);
nor U48830 (N_48830,N_32296,N_31329);
nand U48831 (N_48831,N_38038,N_37283);
xnor U48832 (N_48832,N_36994,N_36341);
nand U48833 (N_48833,N_33659,N_37267);
nand U48834 (N_48834,N_32739,N_37566);
xor U48835 (N_48835,N_37371,N_37217);
or U48836 (N_48836,N_37703,N_38903);
or U48837 (N_48837,N_39281,N_32740);
xor U48838 (N_48838,N_34863,N_39451);
and U48839 (N_48839,N_37148,N_38456);
nor U48840 (N_48840,N_31416,N_38677);
nor U48841 (N_48841,N_38954,N_39815);
xnor U48842 (N_48842,N_38830,N_38202);
and U48843 (N_48843,N_32282,N_34902);
xor U48844 (N_48844,N_30310,N_39187);
and U48845 (N_48845,N_38804,N_30645);
nand U48846 (N_48846,N_36733,N_31315);
xor U48847 (N_48847,N_34893,N_33828);
nand U48848 (N_48848,N_36793,N_30892);
nand U48849 (N_48849,N_35421,N_38215);
nand U48850 (N_48850,N_34154,N_36594);
or U48851 (N_48851,N_33197,N_36268);
xnor U48852 (N_48852,N_32972,N_33085);
nor U48853 (N_48853,N_33650,N_30959);
nand U48854 (N_48854,N_37725,N_31643);
xor U48855 (N_48855,N_37048,N_31835);
nor U48856 (N_48856,N_38004,N_35177);
nand U48857 (N_48857,N_37285,N_34184);
or U48858 (N_48858,N_30412,N_34604);
xnor U48859 (N_48859,N_32391,N_39158);
and U48860 (N_48860,N_39614,N_34412);
nand U48861 (N_48861,N_38548,N_30997);
xnor U48862 (N_48862,N_30288,N_34017);
nand U48863 (N_48863,N_32131,N_32712);
or U48864 (N_48864,N_34704,N_34326);
or U48865 (N_48865,N_34177,N_32741);
or U48866 (N_48866,N_39294,N_37949);
and U48867 (N_48867,N_33935,N_30549);
and U48868 (N_48868,N_37393,N_32800);
nor U48869 (N_48869,N_34692,N_37508);
nor U48870 (N_48870,N_34719,N_32545);
or U48871 (N_48871,N_33500,N_37247);
and U48872 (N_48872,N_37007,N_38784);
or U48873 (N_48873,N_33575,N_37367);
and U48874 (N_48874,N_32442,N_39889);
xor U48875 (N_48875,N_38708,N_30442);
and U48876 (N_48876,N_38204,N_37736);
nor U48877 (N_48877,N_33713,N_35135);
and U48878 (N_48878,N_31483,N_37067);
nand U48879 (N_48879,N_33812,N_34236);
xnor U48880 (N_48880,N_36159,N_33884);
nor U48881 (N_48881,N_34671,N_33378);
and U48882 (N_48882,N_33030,N_38124);
nand U48883 (N_48883,N_38761,N_37758);
and U48884 (N_48884,N_35168,N_33173);
or U48885 (N_48885,N_36504,N_39162);
and U48886 (N_48886,N_31576,N_37630);
and U48887 (N_48887,N_36320,N_34451);
nor U48888 (N_48888,N_33792,N_38569);
and U48889 (N_48889,N_34847,N_39325);
and U48890 (N_48890,N_35180,N_31040);
or U48891 (N_48891,N_38163,N_39201);
nor U48892 (N_48892,N_39443,N_33634);
nor U48893 (N_48893,N_39718,N_30696);
and U48894 (N_48894,N_39596,N_35693);
xor U48895 (N_48895,N_38704,N_32652);
xor U48896 (N_48896,N_32484,N_37385);
or U48897 (N_48897,N_37927,N_38201);
and U48898 (N_48898,N_31239,N_30987);
nor U48899 (N_48899,N_34215,N_34200);
and U48900 (N_48900,N_39479,N_39692);
xor U48901 (N_48901,N_36920,N_37352);
nand U48902 (N_48902,N_31937,N_36135);
xnor U48903 (N_48903,N_30248,N_32537);
xor U48904 (N_48904,N_34801,N_35172);
or U48905 (N_48905,N_38853,N_36898);
xnor U48906 (N_48906,N_32661,N_38004);
xnor U48907 (N_48907,N_30315,N_35430);
xnor U48908 (N_48908,N_39897,N_30707);
and U48909 (N_48909,N_38435,N_39291);
nor U48910 (N_48910,N_38775,N_38065);
nand U48911 (N_48911,N_33583,N_36116);
xor U48912 (N_48912,N_30208,N_32256);
nor U48913 (N_48913,N_31079,N_30547);
nand U48914 (N_48914,N_31871,N_35650);
or U48915 (N_48915,N_32128,N_34563);
or U48916 (N_48916,N_30978,N_33215);
xnor U48917 (N_48917,N_35609,N_35031);
nor U48918 (N_48918,N_37501,N_35501);
xor U48919 (N_48919,N_36112,N_35157);
xor U48920 (N_48920,N_36985,N_31354);
or U48921 (N_48921,N_30428,N_36332);
or U48922 (N_48922,N_38541,N_32278);
nand U48923 (N_48923,N_36141,N_31857);
and U48924 (N_48924,N_38546,N_32856);
nor U48925 (N_48925,N_35885,N_39596);
or U48926 (N_48926,N_30198,N_30840);
nor U48927 (N_48927,N_37308,N_39529);
nand U48928 (N_48928,N_31102,N_34767);
nor U48929 (N_48929,N_35561,N_30466);
nand U48930 (N_48930,N_38783,N_35359);
xor U48931 (N_48931,N_39243,N_31371);
nor U48932 (N_48932,N_32705,N_34367);
and U48933 (N_48933,N_32363,N_37551);
and U48934 (N_48934,N_37023,N_32445);
and U48935 (N_48935,N_34960,N_32817);
or U48936 (N_48936,N_30269,N_32420);
nand U48937 (N_48937,N_39177,N_33485);
nor U48938 (N_48938,N_38096,N_31325);
and U48939 (N_48939,N_34700,N_30824);
xor U48940 (N_48940,N_35351,N_30970);
or U48941 (N_48941,N_30353,N_33365);
and U48942 (N_48942,N_38569,N_35637);
or U48943 (N_48943,N_38490,N_34519);
and U48944 (N_48944,N_39790,N_36754);
and U48945 (N_48945,N_31257,N_38780);
xnor U48946 (N_48946,N_31105,N_39219);
nor U48947 (N_48947,N_36795,N_30885);
or U48948 (N_48948,N_33124,N_33356);
and U48949 (N_48949,N_37696,N_37098);
xnor U48950 (N_48950,N_37150,N_39441);
nand U48951 (N_48951,N_35360,N_30614);
nand U48952 (N_48952,N_32647,N_31937);
nor U48953 (N_48953,N_33257,N_31338);
nand U48954 (N_48954,N_35489,N_33643);
and U48955 (N_48955,N_39950,N_31684);
xnor U48956 (N_48956,N_37563,N_34299);
or U48957 (N_48957,N_32213,N_37739);
nor U48958 (N_48958,N_33739,N_36623);
and U48959 (N_48959,N_34934,N_33040);
or U48960 (N_48960,N_39438,N_31145);
xnor U48961 (N_48961,N_32159,N_35704);
xor U48962 (N_48962,N_33108,N_31151);
and U48963 (N_48963,N_35561,N_30668);
nand U48964 (N_48964,N_37491,N_34928);
nor U48965 (N_48965,N_30959,N_33483);
and U48966 (N_48966,N_30866,N_36175);
xor U48967 (N_48967,N_36756,N_30859);
nand U48968 (N_48968,N_37766,N_35677);
or U48969 (N_48969,N_32421,N_38221);
and U48970 (N_48970,N_35937,N_33671);
nor U48971 (N_48971,N_36656,N_30122);
nor U48972 (N_48972,N_39766,N_36217);
xor U48973 (N_48973,N_36949,N_33141);
and U48974 (N_48974,N_37674,N_36317);
or U48975 (N_48975,N_38938,N_32327);
nand U48976 (N_48976,N_31763,N_39650);
xnor U48977 (N_48977,N_31531,N_35691);
xnor U48978 (N_48978,N_35130,N_31276);
nand U48979 (N_48979,N_33834,N_35895);
and U48980 (N_48980,N_37284,N_38826);
nor U48981 (N_48981,N_31133,N_39767);
xnor U48982 (N_48982,N_33904,N_30488);
or U48983 (N_48983,N_31524,N_33585);
or U48984 (N_48984,N_34395,N_32569);
or U48985 (N_48985,N_33324,N_38718);
nand U48986 (N_48986,N_30653,N_34851);
nor U48987 (N_48987,N_31680,N_31782);
xnor U48988 (N_48988,N_37316,N_36443);
and U48989 (N_48989,N_37971,N_33762);
nor U48990 (N_48990,N_36228,N_32140);
nand U48991 (N_48991,N_38386,N_31866);
xor U48992 (N_48992,N_31649,N_30804);
xor U48993 (N_48993,N_39632,N_37243);
and U48994 (N_48994,N_39724,N_39496);
nor U48995 (N_48995,N_37401,N_39051);
or U48996 (N_48996,N_32969,N_35068);
nor U48997 (N_48997,N_33303,N_38153);
nand U48998 (N_48998,N_38300,N_34596);
or U48999 (N_48999,N_33850,N_31312);
and U49000 (N_49000,N_31928,N_32403);
and U49001 (N_49001,N_30166,N_34789);
nand U49002 (N_49002,N_31636,N_37416);
or U49003 (N_49003,N_33456,N_31986);
or U49004 (N_49004,N_35673,N_38440);
xor U49005 (N_49005,N_38140,N_35115);
xnor U49006 (N_49006,N_39460,N_34275);
and U49007 (N_49007,N_35470,N_37032);
or U49008 (N_49008,N_38409,N_34500);
nor U49009 (N_49009,N_36025,N_33636);
xnor U49010 (N_49010,N_31881,N_33222);
nand U49011 (N_49011,N_32481,N_33615);
or U49012 (N_49012,N_36721,N_35248);
nand U49013 (N_49013,N_30645,N_38786);
and U49014 (N_49014,N_38619,N_39180);
or U49015 (N_49015,N_36385,N_39596);
or U49016 (N_49016,N_32868,N_37133);
nor U49017 (N_49017,N_30303,N_30964);
nand U49018 (N_49018,N_30923,N_30895);
xor U49019 (N_49019,N_34353,N_33892);
nor U49020 (N_49020,N_31593,N_38973);
xor U49021 (N_49021,N_32296,N_30298);
nand U49022 (N_49022,N_39713,N_32390);
nand U49023 (N_49023,N_35478,N_32194);
and U49024 (N_49024,N_32917,N_35438);
nand U49025 (N_49025,N_34026,N_32492);
nor U49026 (N_49026,N_33020,N_30037);
nand U49027 (N_49027,N_36021,N_33741);
and U49028 (N_49028,N_35391,N_32899);
xnor U49029 (N_49029,N_30336,N_31170);
nor U49030 (N_49030,N_31382,N_38842);
or U49031 (N_49031,N_32497,N_33867);
or U49032 (N_49032,N_36465,N_36130);
nor U49033 (N_49033,N_33813,N_37713);
nand U49034 (N_49034,N_35311,N_36510);
xnor U49035 (N_49035,N_36122,N_39502);
xnor U49036 (N_49036,N_39416,N_37677);
nand U49037 (N_49037,N_39897,N_39561);
or U49038 (N_49038,N_35331,N_35386);
and U49039 (N_49039,N_30353,N_37961);
and U49040 (N_49040,N_35946,N_30053);
nor U49041 (N_49041,N_30629,N_31594);
nand U49042 (N_49042,N_35851,N_39173);
and U49043 (N_49043,N_39604,N_39706);
and U49044 (N_49044,N_33220,N_38090);
xor U49045 (N_49045,N_39243,N_32865);
xor U49046 (N_49046,N_39175,N_38807);
nand U49047 (N_49047,N_30921,N_35073);
nand U49048 (N_49048,N_37829,N_35822);
and U49049 (N_49049,N_36379,N_30717);
nor U49050 (N_49050,N_36005,N_39422);
nor U49051 (N_49051,N_31647,N_38252);
nor U49052 (N_49052,N_35632,N_30995);
and U49053 (N_49053,N_37995,N_35083);
or U49054 (N_49054,N_31565,N_38371);
nand U49055 (N_49055,N_38466,N_35744);
nor U49056 (N_49056,N_31645,N_34691);
and U49057 (N_49057,N_37086,N_33799);
xor U49058 (N_49058,N_32261,N_38913);
nand U49059 (N_49059,N_39975,N_36289);
nor U49060 (N_49060,N_36458,N_39606);
nor U49061 (N_49061,N_36255,N_37338);
xor U49062 (N_49062,N_33973,N_37851);
xor U49063 (N_49063,N_39449,N_32549);
xnor U49064 (N_49064,N_32035,N_38081);
xnor U49065 (N_49065,N_34926,N_31367);
and U49066 (N_49066,N_34577,N_39668);
nor U49067 (N_49067,N_36383,N_33958);
xnor U49068 (N_49068,N_31479,N_32087);
nor U49069 (N_49069,N_34162,N_34232);
nand U49070 (N_49070,N_30929,N_32024);
xor U49071 (N_49071,N_37119,N_35025);
and U49072 (N_49072,N_35213,N_39018);
nor U49073 (N_49073,N_39961,N_32249);
nand U49074 (N_49074,N_32497,N_34830);
nor U49075 (N_49075,N_30282,N_33691);
nor U49076 (N_49076,N_35340,N_37953);
or U49077 (N_49077,N_39950,N_35749);
nor U49078 (N_49078,N_31051,N_38568);
nor U49079 (N_49079,N_30292,N_37769);
or U49080 (N_49080,N_31345,N_38751);
and U49081 (N_49081,N_36818,N_34512);
nand U49082 (N_49082,N_34504,N_36295);
nor U49083 (N_49083,N_30966,N_37598);
nand U49084 (N_49084,N_39618,N_36311);
nand U49085 (N_49085,N_33771,N_36137);
nand U49086 (N_49086,N_32396,N_39324);
or U49087 (N_49087,N_35408,N_39422);
or U49088 (N_49088,N_32302,N_38682);
xor U49089 (N_49089,N_34602,N_39860);
xor U49090 (N_49090,N_31534,N_31958);
and U49091 (N_49091,N_35106,N_34381);
and U49092 (N_49092,N_32732,N_35959);
or U49093 (N_49093,N_37038,N_32152);
xor U49094 (N_49094,N_39040,N_32080);
and U49095 (N_49095,N_32044,N_34532);
nor U49096 (N_49096,N_37045,N_37589);
nor U49097 (N_49097,N_37017,N_33154);
xnor U49098 (N_49098,N_39969,N_35219);
nand U49099 (N_49099,N_32431,N_34088);
nor U49100 (N_49100,N_34971,N_33206);
nor U49101 (N_49101,N_35762,N_33500);
and U49102 (N_49102,N_39571,N_34854);
xnor U49103 (N_49103,N_30617,N_30600);
nor U49104 (N_49104,N_37367,N_30939);
nand U49105 (N_49105,N_38031,N_36316);
and U49106 (N_49106,N_30239,N_31323);
xor U49107 (N_49107,N_38577,N_31074);
and U49108 (N_49108,N_32796,N_35149);
and U49109 (N_49109,N_34029,N_35480);
or U49110 (N_49110,N_34798,N_31511);
and U49111 (N_49111,N_35664,N_38703);
xor U49112 (N_49112,N_31332,N_34879);
and U49113 (N_49113,N_35117,N_38107);
nor U49114 (N_49114,N_36090,N_37925);
or U49115 (N_49115,N_37253,N_33654);
xor U49116 (N_49116,N_34769,N_30654);
and U49117 (N_49117,N_30240,N_31668);
or U49118 (N_49118,N_35814,N_34706);
nand U49119 (N_49119,N_31307,N_34288);
nor U49120 (N_49120,N_30516,N_30960);
xnor U49121 (N_49121,N_30416,N_31656);
nand U49122 (N_49122,N_32293,N_35662);
or U49123 (N_49123,N_33799,N_35741);
or U49124 (N_49124,N_39162,N_36806);
nand U49125 (N_49125,N_38092,N_38510);
xor U49126 (N_49126,N_36161,N_31299);
nand U49127 (N_49127,N_35073,N_32468);
xor U49128 (N_49128,N_36601,N_35940);
nor U49129 (N_49129,N_33343,N_34816);
nor U49130 (N_49130,N_37948,N_34369);
or U49131 (N_49131,N_37454,N_36701);
nor U49132 (N_49132,N_30923,N_35917);
nand U49133 (N_49133,N_33877,N_35602);
and U49134 (N_49134,N_39097,N_30064);
nor U49135 (N_49135,N_30218,N_33087);
and U49136 (N_49136,N_37086,N_38106);
xor U49137 (N_49137,N_36337,N_35227);
and U49138 (N_49138,N_34499,N_37263);
nor U49139 (N_49139,N_33177,N_34578);
or U49140 (N_49140,N_33486,N_34261);
and U49141 (N_49141,N_31414,N_39605);
nand U49142 (N_49142,N_37040,N_32372);
xnor U49143 (N_49143,N_36399,N_35126);
nand U49144 (N_49144,N_35767,N_37886);
or U49145 (N_49145,N_37472,N_38539);
nor U49146 (N_49146,N_35442,N_33393);
nor U49147 (N_49147,N_36019,N_34361);
xor U49148 (N_49148,N_36724,N_39845);
xor U49149 (N_49149,N_36914,N_36930);
and U49150 (N_49150,N_32310,N_34523);
xor U49151 (N_49151,N_36760,N_32563);
nor U49152 (N_49152,N_39132,N_34429);
nand U49153 (N_49153,N_30302,N_35590);
nor U49154 (N_49154,N_33073,N_30946);
or U49155 (N_49155,N_37959,N_35356);
nand U49156 (N_49156,N_38309,N_34790);
nor U49157 (N_49157,N_36815,N_35941);
nor U49158 (N_49158,N_38157,N_38640);
nor U49159 (N_49159,N_32365,N_31640);
nor U49160 (N_49160,N_30944,N_38604);
or U49161 (N_49161,N_33677,N_39905);
xnor U49162 (N_49162,N_33555,N_35425);
and U49163 (N_49163,N_33405,N_39333);
nor U49164 (N_49164,N_31734,N_34836);
xnor U49165 (N_49165,N_37701,N_37964);
xor U49166 (N_49166,N_37280,N_35077);
and U49167 (N_49167,N_32407,N_37136);
nand U49168 (N_49168,N_36083,N_34288);
nand U49169 (N_49169,N_33713,N_32105);
nor U49170 (N_49170,N_36445,N_31822);
nor U49171 (N_49171,N_35514,N_35434);
xnor U49172 (N_49172,N_34037,N_34436);
or U49173 (N_49173,N_35880,N_33187);
xnor U49174 (N_49174,N_38459,N_30242);
xnor U49175 (N_49175,N_32951,N_39223);
and U49176 (N_49176,N_32462,N_33143);
xnor U49177 (N_49177,N_39794,N_34231);
xor U49178 (N_49178,N_30601,N_31216);
xnor U49179 (N_49179,N_38520,N_31353);
or U49180 (N_49180,N_33356,N_31473);
and U49181 (N_49181,N_38436,N_31281);
xnor U49182 (N_49182,N_31715,N_33620);
or U49183 (N_49183,N_33323,N_34102);
or U49184 (N_49184,N_32352,N_30620);
nor U49185 (N_49185,N_31709,N_33908);
xor U49186 (N_49186,N_32673,N_36336);
and U49187 (N_49187,N_39716,N_37082);
nand U49188 (N_49188,N_31191,N_37925);
or U49189 (N_49189,N_35335,N_37853);
nand U49190 (N_49190,N_35343,N_35218);
nand U49191 (N_49191,N_36722,N_31268);
nand U49192 (N_49192,N_34447,N_37461);
or U49193 (N_49193,N_34706,N_35174);
nand U49194 (N_49194,N_37671,N_36776);
nand U49195 (N_49195,N_31854,N_33976);
nor U49196 (N_49196,N_32526,N_37303);
or U49197 (N_49197,N_39568,N_36858);
xnor U49198 (N_49198,N_39215,N_35981);
xor U49199 (N_49199,N_31064,N_38387);
xor U49200 (N_49200,N_38094,N_37929);
nand U49201 (N_49201,N_32590,N_37799);
and U49202 (N_49202,N_37733,N_35435);
nand U49203 (N_49203,N_36634,N_33943);
xor U49204 (N_49204,N_30001,N_34373);
or U49205 (N_49205,N_39793,N_34464);
and U49206 (N_49206,N_30734,N_39185);
xnor U49207 (N_49207,N_38555,N_31609);
xnor U49208 (N_49208,N_35448,N_33177);
and U49209 (N_49209,N_35389,N_37193);
xnor U49210 (N_49210,N_34649,N_37368);
and U49211 (N_49211,N_37133,N_37537);
nor U49212 (N_49212,N_37235,N_39575);
nand U49213 (N_49213,N_39029,N_37873);
and U49214 (N_49214,N_31753,N_30176);
nand U49215 (N_49215,N_39035,N_39883);
xor U49216 (N_49216,N_33638,N_39319);
nor U49217 (N_49217,N_39586,N_37628);
and U49218 (N_49218,N_34448,N_39881);
or U49219 (N_49219,N_39675,N_34480);
xnor U49220 (N_49220,N_39086,N_34060);
nand U49221 (N_49221,N_37257,N_36780);
or U49222 (N_49222,N_39437,N_37489);
and U49223 (N_49223,N_38406,N_39914);
and U49224 (N_49224,N_37531,N_34256);
nor U49225 (N_49225,N_33021,N_36916);
or U49226 (N_49226,N_32961,N_39397);
nand U49227 (N_49227,N_32868,N_30931);
nand U49228 (N_49228,N_38003,N_32263);
nand U49229 (N_49229,N_32690,N_31896);
or U49230 (N_49230,N_35723,N_38156);
xnor U49231 (N_49231,N_33800,N_33451);
nand U49232 (N_49232,N_37617,N_38260);
nand U49233 (N_49233,N_30433,N_39925);
and U49234 (N_49234,N_30405,N_32743);
xor U49235 (N_49235,N_36224,N_34013);
xor U49236 (N_49236,N_36705,N_36238);
nand U49237 (N_49237,N_35670,N_39541);
or U49238 (N_49238,N_30685,N_30331);
nor U49239 (N_49239,N_30245,N_34110);
nor U49240 (N_49240,N_30981,N_39232);
nor U49241 (N_49241,N_34830,N_31807);
xor U49242 (N_49242,N_31184,N_34974);
nor U49243 (N_49243,N_35817,N_36284);
and U49244 (N_49244,N_33741,N_37040);
or U49245 (N_49245,N_34423,N_36420);
or U49246 (N_49246,N_32647,N_31966);
nand U49247 (N_49247,N_35873,N_34142);
and U49248 (N_49248,N_36568,N_39542);
nor U49249 (N_49249,N_38599,N_39852);
and U49250 (N_49250,N_30540,N_31777);
nand U49251 (N_49251,N_34811,N_35822);
or U49252 (N_49252,N_35765,N_34371);
nand U49253 (N_49253,N_34602,N_35572);
xnor U49254 (N_49254,N_39187,N_36588);
xnor U49255 (N_49255,N_38139,N_38893);
nor U49256 (N_49256,N_37074,N_38234);
xnor U49257 (N_49257,N_38296,N_35308);
xor U49258 (N_49258,N_31455,N_36770);
nor U49259 (N_49259,N_37484,N_31684);
nand U49260 (N_49260,N_32149,N_39866);
or U49261 (N_49261,N_37016,N_30388);
or U49262 (N_49262,N_32057,N_37968);
nor U49263 (N_49263,N_32390,N_34064);
xor U49264 (N_49264,N_31069,N_31752);
nand U49265 (N_49265,N_37076,N_38566);
nand U49266 (N_49266,N_39305,N_37452);
nor U49267 (N_49267,N_35749,N_36454);
nand U49268 (N_49268,N_36060,N_39726);
xnor U49269 (N_49269,N_39247,N_39956);
nor U49270 (N_49270,N_37808,N_31797);
or U49271 (N_49271,N_39581,N_35565);
nand U49272 (N_49272,N_36082,N_35825);
nor U49273 (N_49273,N_36716,N_39355);
nor U49274 (N_49274,N_33671,N_38954);
or U49275 (N_49275,N_35574,N_31886);
or U49276 (N_49276,N_32579,N_33330);
xnor U49277 (N_49277,N_37416,N_39055);
nand U49278 (N_49278,N_38105,N_32242);
nand U49279 (N_49279,N_38740,N_38048);
and U49280 (N_49280,N_39267,N_34914);
or U49281 (N_49281,N_33074,N_30335);
nor U49282 (N_49282,N_34278,N_35029);
nand U49283 (N_49283,N_38451,N_38640);
nand U49284 (N_49284,N_33392,N_39045);
nor U49285 (N_49285,N_39414,N_35257);
or U49286 (N_49286,N_31683,N_39466);
xor U49287 (N_49287,N_37099,N_35714);
xor U49288 (N_49288,N_36093,N_37944);
or U49289 (N_49289,N_37588,N_31947);
nand U49290 (N_49290,N_37455,N_39631);
nand U49291 (N_49291,N_35766,N_34838);
or U49292 (N_49292,N_34699,N_31033);
nand U49293 (N_49293,N_36169,N_31164);
and U49294 (N_49294,N_32104,N_31601);
xnor U49295 (N_49295,N_35055,N_38631);
or U49296 (N_49296,N_32684,N_31948);
or U49297 (N_49297,N_33374,N_30211);
nand U49298 (N_49298,N_38594,N_34550);
nor U49299 (N_49299,N_33125,N_38674);
and U49300 (N_49300,N_34464,N_36684);
and U49301 (N_49301,N_37196,N_37870);
or U49302 (N_49302,N_31058,N_35727);
nor U49303 (N_49303,N_33290,N_39357);
nand U49304 (N_49304,N_38471,N_32169);
nand U49305 (N_49305,N_37612,N_30756);
and U49306 (N_49306,N_33074,N_30090);
nor U49307 (N_49307,N_32038,N_32095);
and U49308 (N_49308,N_35186,N_33394);
and U49309 (N_49309,N_36636,N_31633);
or U49310 (N_49310,N_30745,N_30005);
nand U49311 (N_49311,N_31604,N_34966);
nand U49312 (N_49312,N_38641,N_31478);
nor U49313 (N_49313,N_36858,N_36451);
nor U49314 (N_49314,N_34583,N_30568);
xor U49315 (N_49315,N_39341,N_34955);
nand U49316 (N_49316,N_37674,N_33086);
nand U49317 (N_49317,N_33216,N_30191);
nor U49318 (N_49318,N_34450,N_35522);
or U49319 (N_49319,N_32244,N_32654);
and U49320 (N_49320,N_32760,N_37093);
and U49321 (N_49321,N_34056,N_31991);
or U49322 (N_49322,N_39357,N_36769);
nor U49323 (N_49323,N_36487,N_37407);
nand U49324 (N_49324,N_36688,N_34842);
and U49325 (N_49325,N_34294,N_35800);
or U49326 (N_49326,N_38908,N_36472);
nand U49327 (N_49327,N_35983,N_32865);
and U49328 (N_49328,N_34797,N_30144);
nand U49329 (N_49329,N_30210,N_38784);
and U49330 (N_49330,N_34431,N_34955);
nor U49331 (N_49331,N_31691,N_33272);
xor U49332 (N_49332,N_33290,N_39713);
and U49333 (N_49333,N_38782,N_39604);
or U49334 (N_49334,N_38658,N_37073);
xor U49335 (N_49335,N_39330,N_34048);
and U49336 (N_49336,N_39240,N_37036);
and U49337 (N_49337,N_38681,N_34561);
and U49338 (N_49338,N_37720,N_39899);
and U49339 (N_49339,N_34728,N_32382);
and U49340 (N_49340,N_36197,N_34255);
nor U49341 (N_49341,N_39777,N_33562);
nor U49342 (N_49342,N_31613,N_36738);
or U49343 (N_49343,N_31184,N_32112);
and U49344 (N_49344,N_35661,N_32790);
or U49345 (N_49345,N_34155,N_33720);
xor U49346 (N_49346,N_34766,N_39784);
nor U49347 (N_49347,N_35509,N_38488);
or U49348 (N_49348,N_32601,N_39098);
and U49349 (N_49349,N_39198,N_31586);
or U49350 (N_49350,N_32206,N_37498);
or U49351 (N_49351,N_33859,N_32729);
or U49352 (N_49352,N_32177,N_32189);
or U49353 (N_49353,N_35160,N_37933);
and U49354 (N_49354,N_31549,N_31373);
and U49355 (N_49355,N_38451,N_33285);
nor U49356 (N_49356,N_35408,N_34857);
and U49357 (N_49357,N_33330,N_30943);
nor U49358 (N_49358,N_33915,N_30205);
xor U49359 (N_49359,N_37266,N_30918);
and U49360 (N_49360,N_31739,N_36933);
and U49361 (N_49361,N_38596,N_35772);
and U49362 (N_49362,N_32535,N_39416);
nor U49363 (N_49363,N_36864,N_39423);
or U49364 (N_49364,N_33785,N_37560);
and U49365 (N_49365,N_35038,N_33764);
nand U49366 (N_49366,N_33742,N_32971);
and U49367 (N_49367,N_36819,N_37687);
nor U49368 (N_49368,N_36700,N_30491);
xor U49369 (N_49369,N_33807,N_32852);
nor U49370 (N_49370,N_34331,N_39035);
and U49371 (N_49371,N_32813,N_30696);
or U49372 (N_49372,N_37670,N_39088);
or U49373 (N_49373,N_35307,N_31772);
nand U49374 (N_49374,N_36300,N_36197);
xnor U49375 (N_49375,N_33577,N_38498);
xor U49376 (N_49376,N_34562,N_32130);
nand U49377 (N_49377,N_38678,N_32655);
or U49378 (N_49378,N_36266,N_39713);
nor U49379 (N_49379,N_37358,N_37572);
or U49380 (N_49380,N_33030,N_30431);
xor U49381 (N_49381,N_32325,N_32971);
nand U49382 (N_49382,N_36264,N_30846);
xnor U49383 (N_49383,N_36553,N_36774);
nor U49384 (N_49384,N_34917,N_35978);
or U49385 (N_49385,N_39068,N_35251);
xnor U49386 (N_49386,N_30422,N_38989);
or U49387 (N_49387,N_35498,N_30653);
or U49388 (N_49388,N_30580,N_30812);
or U49389 (N_49389,N_32323,N_31367);
nor U49390 (N_49390,N_31985,N_35403);
or U49391 (N_49391,N_36643,N_35913);
or U49392 (N_49392,N_39090,N_30325);
xor U49393 (N_49393,N_37157,N_38976);
nand U49394 (N_49394,N_33498,N_38199);
nand U49395 (N_49395,N_30503,N_32324);
nand U49396 (N_49396,N_34735,N_30945);
nand U49397 (N_49397,N_33758,N_33824);
or U49398 (N_49398,N_34373,N_31768);
or U49399 (N_49399,N_37413,N_34234);
or U49400 (N_49400,N_31808,N_35720);
and U49401 (N_49401,N_35284,N_36858);
xor U49402 (N_49402,N_34745,N_38031);
xnor U49403 (N_49403,N_35863,N_30174);
xor U49404 (N_49404,N_33250,N_35648);
nand U49405 (N_49405,N_34722,N_30670);
and U49406 (N_49406,N_32234,N_35360);
xnor U49407 (N_49407,N_30845,N_32192);
nor U49408 (N_49408,N_31885,N_36877);
and U49409 (N_49409,N_38644,N_31716);
or U49410 (N_49410,N_30837,N_39826);
nand U49411 (N_49411,N_37183,N_30859);
or U49412 (N_49412,N_37428,N_36025);
or U49413 (N_49413,N_30668,N_35786);
nand U49414 (N_49414,N_37379,N_31115);
or U49415 (N_49415,N_34154,N_36245);
or U49416 (N_49416,N_38703,N_32321);
nor U49417 (N_49417,N_39038,N_31950);
and U49418 (N_49418,N_39090,N_31728);
nand U49419 (N_49419,N_38526,N_31705);
xnor U49420 (N_49420,N_36623,N_30358);
xnor U49421 (N_49421,N_36893,N_37657);
or U49422 (N_49422,N_39009,N_36378);
and U49423 (N_49423,N_39521,N_36541);
or U49424 (N_49424,N_32220,N_37971);
nor U49425 (N_49425,N_37792,N_39064);
or U49426 (N_49426,N_35251,N_35982);
or U49427 (N_49427,N_35344,N_35503);
nand U49428 (N_49428,N_39123,N_38876);
xnor U49429 (N_49429,N_39254,N_37230);
xor U49430 (N_49430,N_38562,N_33870);
nor U49431 (N_49431,N_39630,N_39283);
nor U49432 (N_49432,N_38547,N_30982);
and U49433 (N_49433,N_30829,N_32272);
nor U49434 (N_49434,N_30003,N_30035);
and U49435 (N_49435,N_31426,N_32486);
nor U49436 (N_49436,N_39982,N_37999);
or U49437 (N_49437,N_35134,N_36815);
and U49438 (N_49438,N_39980,N_30967);
and U49439 (N_49439,N_37157,N_37723);
xor U49440 (N_49440,N_35307,N_33570);
nor U49441 (N_49441,N_33648,N_39213);
xor U49442 (N_49442,N_34683,N_35934);
nand U49443 (N_49443,N_31026,N_35540);
and U49444 (N_49444,N_36571,N_32327);
and U49445 (N_49445,N_38631,N_32073);
xor U49446 (N_49446,N_33954,N_39072);
and U49447 (N_49447,N_32189,N_34076);
nand U49448 (N_49448,N_33830,N_31187);
or U49449 (N_49449,N_33564,N_35916);
xor U49450 (N_49450,N_36788,N_37424);
or U49451 (N_49451,N_35917,N_37905);
nand U49452 (N_49452,N_31024,N_38975);
or U49453 (N_49453,N_39814,N_34178);
and U49454 (N_49454,N_35210,N_36118);
nand U49455 (N_49455,N_34870,N_39054);
or U49456 (N_49456,N_37548,N_35015);
or U49457 (N_49457,N_38727,N_31261);
nor U49458 (N_49458,N_37297,N_35643);
and U49459 (N_49459,N_31236,N_39246);
xnor U49460 (N_49460,N_32762,N_31286);
nand U49461 (N_49461,N_37067,N_31491);
nor U49462 (N_49462,N_33718,N_35459);
or U49463 (N_49463,N_38929,N_33739);
nand U49464 (N_49464,N_32599,N_35399);
xor U49465 (N_49465,N_31824,N_31291);
nor U49466 (N_49466,N_32806,N_35813);
nand U49467 (N_49467,N_37152,N_34209);
and U49468 (N_49468,N_31159,N_30453);
nor U49469 (N_49469,N_32004,N_34432);
and U49470 (N_49470,N_31631,N_35535);
xnor U49471 (N_49471,N_33278,N_33149);
nand U49472 (N_49472,N_39514,N_37167);
xor U49473 (N_49473,N_31594,N_35620);
or U49474 (N_49474,N_38064,N_36441);
xnor U49475 (N_49475,N_32688,N_39120);
xor U49476 (N_49476,N_33572,N_37073);
nor U49477 (N_49477,N_30272,N_36603);
nor U49478 (N_49478,N_35484,N_34694);
and U49479 (N_49479,N_31591,N_31075);
xor U49480 (N_49480,N_39852,N_32461);
or U49481 (N_49481,N_37940,N_30642);
and U49482 (N_49482,N_35635,N_38351);
or U49483 (N_49483,N_39945,N_35460);
nor U49484 (N_49484,N_32601,N_31444);
and U49485 (N_49485,N_37503,N_31129);
nand U49486 (N_49486,N_30763,N_35596);
xor U49487 (N_49487,N_38644,N_36350);
xor U49488 (N_49488,N_34039,N_32475);
or U49489 (N_49489,N_38668,N_31175);
or U49490 (N_49490,N_31512,N_34727);
nor U49491 (N_49491,N_36455,N_33601);
xnor U49492 (N_49492,N_32087,N_38463);
nand U49493 (N_49493,N_35253,N_32037);
nor U49494 (N_49494,N_33012,N_31880);
or U49495 (N_49495,N_32286,N_39423);
and U49496 (N_49496,N_32659,N_35560);
xnor U49497 (N_49497,N_34440,N_35325);
xnor U49498 (N_49498,N_33676,N_36429);
xnor U49499 (N_49499,N_32027,N_39929);
xnor U49500 (N_49500,N_32305,N_34361);
or U49501 (N_49501,N_33692,N_36764);
xnor U49502 (N_49502,N_32838,N_38254);
or U49503 (N_49503,N_37026,N_36256);
nand U49504 (N_49504,N_39875,N_39566);
nand U49505 (N_49505,N_33487,N_38134);
nand U49506 (N_49506,N_30282,N_30441);
and U49507 (N_49507,N_34761,N_36418);
nand U49508 (N_49508,N_34002,N_33785);
xnor U49509 (N_49509,N_38506,N_37090);
and U49510 (N_49510,N_31184,N_33889);
nand U49511 (N_49511,N_31300,N_39669);
or U49512 (N_49512,N_32364,N_34538);
xor U49513 (N_49513,N_38867,N_30138);
xor U49514 (N_49514,N_31401,N_36510);
xor U49515 (N_49515,N_30898,N_38324);
nand U49516 (N_49516,N_34141,N_38439);
xnor U49517 (N_49517,N_39114,N_34196);
xnor U49518 (N_49518,N_31077,N_30229);
or U49519 (N_49519,N_36969,N_30245);
xor U49520 (N_49520,N_39924,N_35789);
and U49521 (N_49521,N_37385,N_35072);
nor U49522 (N_49522,N_37574,N_33252);
nor U49523 (N_49523,N_34220,N_38375);
and U49524 (N_49524,N_37349,N_39436);
or U49525 (N_49525,N_30751,N_30211);
and U49526 (N_49526,N_37220,N_36061);
nor U49527 (N_49527,N_35126,N_32765);
or U49528 (N_49528,N_36488,N_31240);
nand U49529 (N_49529,N_36927,N_39109);
and U49530 (N_49530,N_35369,N_32290);
and U49531 (N_49531,N_31008,N_32679);
or U49532 (N_49532,N_34233,N_37707);
nand U49533 (N_49533,N_33645,N_30409);
nor U49534 (N_49534,N_31166,N_37126);
xnor U49535 (N_49535,N_37217,N_34045);
and U49536 (N_49536,N_35296,N_32147);
nand U49537 (N_49537,N_33994,N_39416);
or U49538 (N_49538,N_33684,N_30927);
xnor U49539 (N_49539,N_39758,N_33914);
nor U49540 (N_49540,N_37859,N_33258);
nor U49541 (N_49541,N_36060,N_33362);
and U49542 (N_49542,N_39529,N_38701);
nand U49543 (N_49543,N_38278,N_38684);
and U49544 (N_49544,N_39095,N_32173);
nor U49545 (N_49545,N_37311,N_39646);
nand U49546 (N_49546,N_39448,N_34731);
and U49547 (N_49547,N_39650,N_36060);
or U49548 (N_49548,N_32207,N_32495);
nand U49549 (N_49549,N_37049,N_30667);
nand U49550 (N_49550,N_30270,N_38166);
or U49551 (N_49551,N_31230,N_33680);
nand U49552 (N_49552,N_39649,N_38305);
nand U49553 (N_49553,N_33379,N_33286);
or U49554 (N_49554,N_39716,N_34268);
and U49555 (N_49555,N_37138,N_37490);
xnor U49556 (N_49556,N_30795,N_30199);
xnor U49557 (N_49557,N_31555,N_34174);
nand U49558 (N_49558,N_33535,N_32049);
and U49559 (N_49559,N_38069,N_35595);
xor U49560 (N_49560,N_33353,N_34292);
xor U49561 (N_49561,N_31578,N_34989);
nor U49562 (N_49562,N_36784,N_34219);
nand U49563 (N_49563,N_31416,N_38002);
and U49564 (N_49564,N_39145,N_36238);
nand U49565 (N_49565,N_39272,N_38174);
nand U49566 (N_49566,N_33954,N_31610);
xnor U49567 (N_49567,N_36814,N_30951);
nand U49568 (N_49568,N_38603,N_39072);
or U49569 (N_49569,N_30987,N_37292);
and U49570 (N_49570,N_33910,N_35914);
or U49571 (N_49571,N_30208,N_36521);
or U49572 (N_49572,N_39617,N_35811);
and U49573 (N_49573,N_33010,N_36814);
nand U49574 (N_49574,N_35101,N_30525);
and U49575 (N_49575,N_31356,N_36005);
xnor U49576 (N_49576,N_39500,N_33883);
or U49577 (N_49577,N_37029,N_35651);
nor U49578 (N_49578,N_34436,N_39924);
xor U49579 (N_49579,N_37749,N_32914);
and U49580 (N_49580,N_34760,N_36633);
xor U49581 (N_49581,N_32929,N_33638);
nor U49582 (N_49582,N_32115,N_31947);
nand U49583 (N_49583,N_34205,N_36256);
nand U49584 (N_49584,N_35228,N_35352);
or U49585 (N_49585,N_38942,N_32630);
xor U49586 (N_49586,N_36928,N_33498);
or U49587 (N_49587,N_30886,N_33196);
and U49588 (N_49588,N_33759,N_38850);
nor U49589 (N_49589,N_30302,N_32550);
nor U49590 (N_49590,N_31326,N_35202);
nor U49591 (N_49591,N_34381,N_38821);
nor U49592 (N_49592,N_39268,N_35111);
nor U49593 (N_49593,N_39165,N_30231);
and U49594 (N_49594,N_36847,N_36050);
nor U49595 (N_49595,N_31102,N_38264);
or U49596 (N_49596,N_35402,N_38129);
or U49597 (N_49597,N_39401,N_39497);
and U49598 (N_49598,N_37418,N_38706);
and U49599 (N_49599,N_31665,N_31127);
nand U49600 (N_49600,N_36120,N_38484);
nand U49601 (N_49601,N_37377,N_34763);
and U49602 (N_49602,N_39200,N_35293);
nor U49603 (N_49603,N_39779,N_31134);
and U49604 (N_49604,N_30407,N_39800);
nor U49605 (N_49605,N_35726,N_38266);
or U49606 (N_49606,N_37172,N_35758);
nand U49607 (N_49607,N_33618,N_33390);
or U49608 (N_49608,N_31777,N_30349);
nor U49609 (N_49609,N_35584,N_33459);
and U49610 (N_49610,N_37658,N_38686);
and U49611 (N_49611,N_31795,N_30358);
and U49612 (N_49612,N_33195,N_37161);
nand U49613 (N_49613,N_36666,N_32838);
and U49614 (N_49614,N_30188,N_32331);
nor U49615 (N_49615,N_31407,N_31099);
or U49616 (N_49616,N_36658,N_34687);
xor U49617 (N_49617,N_36799,N_36660);
nor U49618 (N_49618,N_36457,N_38409);
nor U49619 (N_49619,N_34881,N_39221);
xor U49620 (N_49620,N_32787,N_30815);
xnor U49621 (N_49621,N_34919,N_35154);
or U49622 (N_49622,N_33237,N_38103);
nor U49623 (N_49623,N_38430,N_39804);
or U49624 (N_49624,N_32841,N_31202);
or U49625 (N_49625,N_36074,N_39325);
or U49626 (N_49626,N_38381,N_33243);
nand U49627 (N_49627,N_32557,N_34133);
or U49628 (N_49628,N_37130,N_32069);
nor U49629 (N_49629,N_37006,N_34367);
and U49630 (N_49630,N_34661,N_38502);
and U49631 (N_49631,N_31172,N_39154);
nor U49632 (N_49632,N_36649,N_39622);
xnor U49633 (N_49633,N_32471,N_31300);
or U49634 (N_49634,N_32996,N_31386);
and U49635 (N_49635,N_38136,N_39190);
and U49636 (N_49636,N_39919,N_37560);
and U49637 (N_49637,N_37652,N_37361);
nor U49638 (N_49638,N_30575,N_34055);
and U49639 (N_49639,N_30330,N_36457);
xnor U49640 (N_49640,N_37373,N_37998);
nand U49641 (N_49641,N_35076,N_31170);
nor U49642 (N_49642,N_36839,N_35299);
nor U49643 (N_49643,N_31834,N_32479);
nand U49644 (N_49644,N_35225,N_34606);
or U49645 (N_49645,N_34852,N_35819);
nor U49646 (N_49646,N_35470,N_31352);
nor U49647 (N_49647,N_30649,N_38643);
nand U49648 (N_49648,N_38365,N_36888);
nor U49649 (N_49649,N_31011,N_35189);
nor U49650 (N_49650,N_33500,N_35523);
nand U49651 (N_49651,N_30873,N_38331);
or U49652 (N_49652,N_33612,N_33604);
xnor U49653 (N_49653,N_34343,N_36943);
xnor U49654 (N_49654,N_31050,N_32797);
and U49655 (N_49655,N_32017,N_34519);
xor U49656 (N_49656,N_36981,N_35962);
and U49657 (N_49657,N_32551,N_39252);
or U49658 (N_49658,N_32029,N_31540);
xnor U49659 (N_49659,N_31685,N_38675);
nand U49660 (N_49660,N_32207,N_34409);
xnor U49661 (N_49661,N_39448,N_38156);
and U49662 (N_49662,N_31235,N_39644);
xnor U49663 (N_49663,N_36293,N_33801);
and U49664 (N_49664,N_34496,N_39466);
xor U49665 (N_49665,N_30763,N_34514);
nor U49666 (N_49666,N_35681,N_37735);
nor U49667 (N_49667,N_30869,N_38926);
or U49668 (N_49668,N_32884,N_32162);
xor U49669 (N_49669,N_38702,N_39059);
or U49670 (N_49670,N_35553,N_36501);
xor U49671 (N_49671,N_32023,N_35360);
nor U49672 (N_49672,N_39969,N_35864);
nor U49673 (N_49673,N_38638,N_38722);
or U49674 (N_49674,N_35728,N_38931);
nand U49675 (N_49675,N_30135,N_39114);
nor U49676 (N_49676,N_36882,N_31838);
xnor U49677 (N_49677,N_31157,N_34144);
xor U49678 (N_49678,N_34503,N_34727);
nor U49679 (N_49679,N_31096,N_37484);
or U49680 (N_49680,N_32745,N_31361);
xnor U49681 (N_49681,N_30641,N_37739);
nor U49682 (N_49682,N_38637,N_34003);
and U49683 (N_49683,N_31224,N_31665);
nand U49684 (N_49684,N_36380,N_35183);
nor U49685 (N_49685,N_38809,N_39252);
xor U49686 (N_49686,N_33843,N_32753);
nor U49687 (N_49687,N_36649,N_38351);
xnor U49688 (N_49688,N_32412,N_35198);
and U49689 (N_49689,N_30144,N_31516);
nor U49690 (N_49690,N_36206,N_33819);
nor U49691 (N_49691,N_38360,N_31337);
xor U49692 (N_49692,N_35461,N_36813);
nand U49693 (N_49693,N_37759,N_32487);
nand U49694 (N_49694,N_30658,N_31906);
nor U49695 (N_49695,N_35913,N_37403);
nand U49696 (N_49696,N_39594,N_36579);
xnor U49697 (N_49697,N_32614,N_36215);
or U49698 (N_49698,N_33243,N_31894);
xor U49699 (N_49699,N_35495,N_36958);
nand U49700 (N_49700,N_36630,N_35298);
xor U49701 (N_49701,N_33055,N_33981);
and U49702 (N_49702,N_32181,N_30511);
or U49703 (N_49703,N_38547,N_39250);
xnor U49704 (N_49704,N_38583,N_39087);
and U49705 (N_49705,N_34135,N_30169);
nand U49706 (N_49706,N_39712,N_36777);
xor U49707 (N_49707,N_38211,N_37134);
nor U49708 (N_49708,N_36134,N_39721);
nor U49709 (N_49709,N_33573,N_34056);
or U49710 (N_49710,N_30123,N_39682);
or U49711 (N_49711,N_36085,N_33213);
and U49712 (N_49712,N_30422,N_39938);
nor U49713 (N_49713,N_37409,N_31206);
or U49714 (N_49714,N_37730,N_38125);
and U49715 (N_49715,N_33267,N_34098);
or U49716 (N_49716,N_31650,N_30871);
nand U49717 (N_49717,N_31740,N_37153);
nor U49718 (N_49718,N_34121,N_39694);
or U49719 (N_49719,N_32218,N_31223);
and U49720 (N_49720,N_37610,N_34578);
and U49721 (N_49721,N_32684,N_39718);
and U49722 (N_49722,N_39504,N_36045);
xnor U49723 (N_49723,N_34312,N_30679);
xnor U49724 (N_49724,N_35703,N_35166);
and U49725 (N_49725,N_32315,N_33315);
and U49726 (N_49726,N_34377,N_38786);
or U49727 (N_49727,N_32345,N_33628);
xor U49728 (N_49728,N_35472,N_34147);
and U49729 (N_49729,N_33804,N_36196);
and U49730 (N_49730,N_32061,N_37409);
or U49731 (N_49731,N_35233,N_30558);
nand U49732 (N_49732,N_38650,N_35129);
and U49733 (N_49733,N_31812,N_39482);
nor U49734 (N_49734,N_39204,N_30160);
nor U49735 (N_49735,N_36484,N_31772);
nor U49736 (N_49736,N_37129,N_35858);
nand U49737 (N_49737,N_32453,N_38799);
or U49738 (N_49738,N_35658,N_31879);
and U49739 (N_49739,N_30714,N_31977);
nand U49740 (N_49740,N_31076,N_32981);
nor U49741 (N_49741,N_35790,N_38530);
or U49742 (N_49742,N_34179,N_30336);
nand U49743 (N_49743,N_37252,N_35644);
xor U49744 (N_49744,N_37124,N_33173);
xor U49745 (N_49745,N_38782,N_33271);
nor U49746 (N_49746,N_35587,N_38375);
nor U49747 (N_49747,N_33014,N_34365);
nor U49748 (N_49748,N_39908,N_36882);
nor U49749 (N_49749,N_37884,N_31412);
nor U49750 (N_49750,N_34885,N_34264);
xor U49751 (N_49751,N_32469,N_36269);
nand U49752 (N_49752,N_39612,N_34663);
nor U49753 (N_49753,N_32666,N_38869);
nand U49754 (N_49754,N_30543,N_32517);
and U49755 (N_49755,N_30263,N_35557);
and U49756 (N_49756,N_36356,N_39306);
nand U49757 (N_49757,N_37408,N_34297);
nand U49758 (N_49758,N_33998,N_32087);
or U49759 (N_49759,N_35511,N_30920);
nand U49760 (N_49760,N_38648,N_35761);
nand U49761 (N_49761,N_31143,N_31938);
and U49762 (N_49762,N_32013,N_34091);
and U49763 (N_49763,N_35959,N_37598);
xor U49764 (N_49764,N_38089,N_35955);
xnor U49765 (N_49765,N_37954,N_37584);
and U49766 (N_49766,N_38745,N_38760);
or U49767 (N_49767,N_30757,N_34501);
or U49768 (N_49768,N_37635,N_31313);
or U49769 (N_49769,N_32530,N_39614);
nor U49770 (N_49770,N_33083,N_37864);
nor U49771 (N_49771,N_39896,N_30715);
or U49772 (N_49772,N_33117,N_35748);
xor U49773 (N_49773,N_37077,N_31680);
nand U49774 (N_49774,N_37716,N_35116);
and U49775 (N_49775,N_33970,N_37786);
or U49776 (N_49776,N_30704,N_32840);
and U49777 (N_49777,N_32150,N_37733);
xor U49778 (N_49778,N_33944,N_39122);
and U49779 (N_49779,N_33534,N_32333);
or U49780 (N_49780,N_33945,N_33357);
nand U49781 (N_49781,N_36125,N_35930);
nor U49782 (N_49782,N_31430,N_34708);
or U49783 (N_49783,N_39450,N_37445);
or U49784 (N_49784,N_38444,N_36188);
nor U49785 (N_49785,N_36553,N_33027);
and U49786 (N_49786,N_34471,N_33397);
nor U49787 (N_49787,N_34228,N_36659);
nand U49788 (N_49788,N_39457,N_37349);
nor U49789 (N_49789,N_32275,N_36444);
and U49790 (N_49790,N_32573,N_30413);
and U49791 (N_49791,N_36727,N_38599);
or U49792 (N_49792,N_36786,N_32928);
and U49793 (N_49793,N_36657,N_37784);
or U49794 (N_49794,N_38667,N_38275);
xnor U49795 (N_49795,N_34374,N_34189);
and U49796 (N_49796,N_36152,N_32155);
and U49797 (N_49797,N_34505,N_37078);
and U49798 (N_49798,N_36970,N_34463);
nor U49799 (N_49799,N_33707,N_35893);
and U49800 (N_49800,N_38115,N_39149);
and U49801 (N_49801,N_38026,N_36299);
xnor U49802 (N_49802,N_39704,N_38289);
and U49803 (N_49803,N_33150,N_39943);
nor U49804 (N_49804,N_33208,N_32469);
nor U49805 (N_49805,N_31775,N_36850);
nor U49806 (N_49806,N_38990,N_38008);
nand U49807 (N_49807,N_36977,N_31148);
nor U49808 (N_49808,N_35983,N_35993);
and U49809 (N_49809,N_37983,N_35871);
nand U49810 (N_49810,N_37926,N_35175);
and U49811 (N_49811,N_36131,N_33789);
nand U49812 (N_49812,N_30450,N_35982);
and U49813 (N_49813,N_35376,N_35782);
or U49814 (N_49814,N_35163,N_36011);
nor U49815 (N_49815,N_36264,N_37124);
and U49816 (N_49816,N_39230,N_30122);
xnor U49817 (N_49817,N_34410,N_39848);
nand U49818 (N_49818,N_39378,N_36218);
nand U49819 (N_49819,N_32421,N_32913);
and U49820 (N_49820,N_30539,N_34116);
or U49821 (N_49821,N_31144,N_38589);
or U49822 (N_49822,N_30394,N_37305);
or U49823 (N_49823,N_38893,N_34646);
xnor U49824 (N_49824,N_36785,N_36853);
or U49825 (N_49825,N_36126,N_32961);
xnor U49826 (N_49826,N_36194,N_37848);
and U49827 (N_49827,N_33787,N_38273);
or U49828 (N_49828,N_32401,N_30391);
nor U49829 (N_49829,N_34787,N_33640);
nor U49830 (N_49830,N_37276,N_30458);
xor U49831 (N_49831,N_38965,N_33341);
nor U49832 (N_49832,N_35754,N_36082);
nand U49833 (N_49833,N_31628,N_35629);
or U49834 (N_49834,N_32375,N_38267);
xnor U49835 (N_49835,N_33478,N_37198);
nor U49836 (N_49836,N_30920,N_38958);
nor U49837 (N_49837,N_30810,N_32566);
nand U49838 (N_49838,N_35990,N_34194);
nor U49839 (N_49839,N_37747,N_31891);
or U49840 (N_49840,N_37859,N_37449);
or U49841 (N_49841,N_31374,N_35549);
xor U49842 (N_49842,N_33922,N_32534);
nor U49843 (N_49843,N_39540,N_32805);
and U49844 (N_49844,N_32449,N_38372);
nor U49845 (N_49845,N_37504,N_38676);
or U49846 (N_49846,N_33879,N_33331);
xnor U49847 (N_49847,N_37192,N_35392);
and U49848 (N_49848,N_30369,N_33757);
nand U49849 (N_49849,N_38045,N_31190);
nor U49850 (N_49850,N_30144,N_39114);
nor U49851 (N_49851,N_38830,N_30425);
and U49852 (N_49852,N_32170,N_34508);
or U49853 (N_49853,N_37637,N_38351);
and U49854 (N_49854,N_39049,N_37389);
xnor U49855 (N_49855,N_33887,N_37693);
nor U49856 (N_49856,N_33246,N_36136);
or U49857 (N_49857,N_36760,N_32744);
or U49858 (N_49858,N_34104,N_34988);
and U49859 (N_49859,N_38203,N_39813);
xnor U49860 (N_49860,N_35710,N_39390);
nand U49861 (N_49861,N_33402,N_36074);
nand U49862 (N_49862,N_31115,N_38500);
xnor U49863 (N_49863,N_37047,N_37571);
nor U49864 (N_49864,N_33323,N_31533);
xor U49865 (N_49865,N_36742,N_37288);
xnor U49866 (N_49866,N_34307,N_30976);
and U49867 (N_49867,N_33648,N_37684);
xnor U49868 (N_49868,N_35460,N_30140);
nand U49869 (N_49869,N_33994,N_31521);
nand U49870 (N_49870,N_30721,N_36847);
nor U49871 (N_49871,N_34336,N_37960);
xnor U49872 (N_49872,N_30302,N_36641);
and U49873 (N_49873,N_38436,N_32215);
nor U49874 (N_49874,N_35466,N_32792);
or U49875 (N_49875,N_32518,N_39627);
xor U49876 (N_49876,N_30291,N_30283);
nand U49877 (N_49877,N_36255,N_32404);
or U49878 (N_49878,N_37956,N_36446);
xor U49879 (N_49879,N_35767,N_30653);
and U49880 (N_49880,N_35346,N_38165);
xor U49881 (N_49881,N_30365,N_30259);
nand U49882 (N_49882,N_31280,N_33500);
or U49883 (N_49883,N_34446,N_38282);
xor U49884 (N_49884,N_33927,N_33756);
and U49885 (N_49885,N_38056,N_31127);
nor U49886 (N_49886,N_35438,N_32724);
nor U49887 (N_49887,N_36672,N_37733);
and U49888 (N_49888,N_36126,N_32693);
nand U49889 (N_49889,N_39548,N_38269);
xor U49890 (N_49890,N_37592,N_39252);
or U49891 (N_49891,N_36259,N_37894);
or U49892 (N_49892,N_39823,N_39085);
nor U49893 (N_49893,N_39468,N_37152);
nand U49894 (N_49894,N_34443,N_33040);
nor U49895 (N_49895,N_39184,N_38019);
nor U49896 (N_49896,N_34068,N_33722);
xor U49897 (N_49897,N_36127,N_39300);
nor U49898 (N_49898,N_38604,N_38066);
nand U49899 (N_49899,N_36702,N_38946);
xnor U49900 (N_49900,N_38071,N_33456);
xor U49901 (N_49901,N_35900,N_33967);
xnor U49902 (N_49902,N_31069,N_38356);
and U49903 (N_49903,N_31266,N_35981);
nor U49904 (N_49904,N_31814,N_33008);
xnor U49905 (N_49905,N_30605,N_32519);
and U49906 (N_49906,N_36910,N_37061);
and U49907 (N_49907,N_34237,N_30493);
nand U49908 (N_49908,N_36597,N_36836);
nand U49909 (N_49909,N_33841,N_31903);
nor U49910 (N_49910,N_39091,N_36364);
xnor U49911 (N_49911,N_31174,N_33803);
and U49912 (N_49912,N_30410,N_35650);
nor U49913 (N_49913,N_37279,N_35561);
xor U49914 (N_49914,N_32779,N_39082);
xor U49915 (N_49915,N_37744,N_35959);
nand U49916 (N_49916,N_38370,N_34513);
nor U49917 (N_49917,N_33670,N_39801);
nor U49918 (N_49918,N_31559,N_37475);
nand U49919 (N_49919,N_34706,N_37490);
nand U49920 (N_49920,N_33431,N_31708);
nor U49921 (N_49921,N_35115,N_32660);
nand U49922 (N_49922,N_33172,N_39374);
nor U49923 (N_49923,N_38933,N_35775);
or U49924 (N_49924,N_38534,N_39269);
nand U49925 (N_49925,N_38067,N_38875);
nand U49926 (N_49926,N_31943,N_35016);
or U49927 (N_49927,N_32414,N_34753);
and U49928 (N_49928,N_38582,N_34818);
or U49929 (N_49929,N_37832,N_30729);
and U49930 (N_49930,N_30326,N_33673);
xnor U49931 (N_49931,N_37640,N_32911);
and U49932 (N_49932,N_31577,N_34220);
or U49933 (N_49933,N_38031,N_31396);
nor U49934 (N_49934,N_37394,N_35233);
and U49935 (N_49935,N_32875,N_34794);
nand U49936 (N_49936,N_31125,N_33636);
or U49937 (N_49937,N_38588,N_32890);
xnor U49938 (N_49938,N_35810,N_36310);
and U49939 (N_49939,N_39893,N_36139);
and U49940 (N_49940,N_37652,N_39527);
xor U49941 (N_49941,N_37521,N_37776);
nand U49942 (N_49942,N_30217,N_33065);
and U49943 (N_49943,N_33652,N_34502);
nor U49944 (N_49944,N_30793,N_30510);
nand U49945 (N_49945,N_33609,N_37988);
xor U49946 (N_49946,N_38595,N_39390);
and U49947 (N_49947,N_35988,N_31447);
nand U49948 (N_49948,N_39421,N_37152);
and U49949 (N_49949,N_31901,N_32982);
or U49950 (N_49950,N_38921,N_34764);
nand U49951 (N_49951,N_32961,N_31163);
and U49952 (N_49952,N_36982,N_31007);
and U49953 (N_49953,N_32789,N_38052);
and U49954 (N_49954,N_38098,N_37358);
xnor U49955 (N_49955,N_30063,N_33179);
or U49956 (N_49956,N_34384,N_30015);
xor U49957 (N_49957,N_39350,N_38398);
and U49958 (N_49958,N_33941,N_38251);
nor U49959 (N_49959,N_34610,N_37419);
and U49960 (N_49960,N_35019,N_31375);
xor U49961 (N_49961,N_32102,N_30574);
nor U49962 (N_49962,N_32262,N_33479);
and U49963 (N_49963,N_38912,N_30667);
xor U49964 (N_49964,N_31844,N_30635);
xor U49965 (N_49965,N_34468,N_32266);
and U49966 (N_49966,N_36640,N_33290);
and U49967 (N_49967,N_39253,N_35023);
nor U49968 (N_49968,N_36410,N_37258);
nor U49969 (N_49969,N_38626,N_31176);
nor U49970 (N_49970,N_39732,N_33347);
and U49971 (N_49971,N_34221,N_38142);
and U49972 (N_49972,N_34040,N_37542);
xnor U49973 (N_49973,N_33719,N_38663);
and U49974 (N_49974,N_31525,N_30670);
nand U49975 (N_49975,N_34124,N_33977);
or U49976 (N_49976,N_35036,N_39695);
and U49977 (N_49977,N_33744,N_30173);
nand U49978 (N_49978,N_33253,N_37400);
nor U49979 (N_49979,N_36911,N_39259);
nand U49980 (N_49980,N_35403,N_37819);
nand U49981 (N_49981,N_33413,N_36908);
nor U49982 (N_49982,N_37599,N_35572);
nor U49983 (N_49983,N_34675,N_30561);
xnor U49984 (N_49984,N_32839,N_38865);
xnor U49985 (N_49985,N_39245,N_33344);
or U49986 (N_49986,N_36147,N_31321);
nand U49987 (N_49987,N_38511,N_30246);
or U49988 (N_49988,N_37891,N_33703);
or U49989 (N_49989,N_33626,N_33476);
nand U49990 (N_49990,N_33018,N_34566);
nor U49991 (N_49991,N_32278,N_39743);
nand U49992 (N_49992,N_38551,N_30905);
nand U49993 (N_49993,N_36749,N_32625);
nand U49994 (N_49994,N_31690,N_37774);
nor U49995 (N_49995,N_33993,N_37487);
nor U49996 (N_49996,N_38844,N_37304);
xnor U49997 (N_49997,N_38148,N_37188);
and U49998 (N_49998,N_31761,N_33716);
nand U49999 (N_49999,N_32692,N_38571);
xor UO_0 (O_0,N_46747,N_41949);
nor UO_1 (O_1,N_43843,N_40286);
or UO_2 (O_2,N_42521,N_44063);
nand UO_3 (O_3,N_46301,N_45980);
or UO_4 (O_4,N_47673,N_45519);
nand UO_5 (O_5,N_49264,N_45248);
or UO_6 (O_6,N_47794,N_44600);
or UO_7 (O_7,N_45263,N_47972);
xor UO_8 (O_8,N_46298,N_49029);
nor UO_9 (O_9,N_41868,N_45262);
nand UO_10 (O_10,N_43967,N_46876);
nand UO_11 (O_11,N_41016,N_43154);
and UO_12 (O_12,N_40499,N_47613);
and UO_13 (O_13,N_47158,N_49953);
xor UO_14 (O_14,N_48842,N_47577);
and UO_15 (O_15,N_47333,N_46801);
or UO_16 (O_16,N_41800,N_48690);
and UO_17 (O_17,N_48064,N_48532);
xnor UO_18 (O_18,N_46192,N_49521);
nor UO_19 (O_19,N_45373,N_42864);
and UO_20 (O_20,N_45331,N_45634);
and UO_21 (O_21,N_40422,N_42891);
nor UO_22 (O_22,N_40373,N_44033);
and UO_23 (O_23,N_41456,N_47006);
nor UO_24 (O_24,N_45848,N_49403);
nand UO_25 (O_25,N_45729,N_48958);
and UO_26 (O_26,N_42036,N_43890);
nand UO_27 (O_27,N_42425,N_46935);
xor UO_28 (O_28,N_41341,N_45659);
xor UO_29 (O_29,N_44912,N_42576);
nor UO_30 (O_30,N_47290,N_48676);
nor UO_31 (O_31,N_40088,N_47220);
and UO_32 (O_32,N_43150,N_40254);
nor UO_33 (O_33,N_49528,N_41429);
or UO_34 (O_34,N_41746,N_42393);
nor UO_35 (O_35,N_40262,N_42434);
nor UO_36 (O_36,N_45432,N_46536);
nand UO_37 (O_37,N_48406,N_47259);
nor UO_38 (O_38,N_48513,N_42384);
and UO_39 (O_39,N_40869,N_49415);
nor UO_40 (O_40,N_47833,N_46116);
nand UO_41 (O_41,N_44779,N_46916);
nor UO_42 (O_42,N_41097,N_45922);
and UO_43 (O_43,N_49249,N_47084);
xor UO_44 (O_44,N_46158,N_44003);
and UO_45 (O_45,N_40123,N_42059);
xnor UO_46 (O_46,N_49676,N_48651);
and UO_47 (O_47,N_47987,N_44897);
and UO_48 (O_48,N_46091,N_42267);
or UO_49 (O_49,N_48557,N_48585);
xnor UO_50 (O_50,N_40953,N_48685);
nor UO_51 (O_51,N_48621,N_47885);
and UO_52 (O_52,N_48200,N_40457);
nand UO_53 (O_53,N_48490,N_42728);
nand UO_54 (O_54,N_45523,N_41108);
and UO_55 (O_55,N_43585,N_48365);
xor UO_56 (O_56,N_43750,N_49305);
or UO_57 (O_57,N_40031,N_48259);
nor UO_58 (O_58,N_41845,N_44174);
or UO_59 (O_59,N_48859,N_47891);
or UO_60 (O_60,N_40363,N_48874);
and UO_61 (O_61,N_44958,N_40926);
xnor UO_62 (O_62,N_44244,N_49153);
or UO_63 (O_63,N_42895,N_48765);
nor UO_64 (O_64,N_47732,N_40583);
nor UO_65 (O_65,N_42751,N_45626);
nor UO_66 (O_66,N_47371,N_45058);
nand UO_67 (O_67,N_42913,N_47432);
nor UO_68 (O_68,N_47976,N_44368);
or UO_69 (O_69,N_47664,N_49369);
and UO_70 (O_70,N_40812,N_49072);
nor UO_71 (O_71,N_41044,N_44420);
and UO_72 (O_72,N_45055,N_40862);
xnor UO_73 (O_73,N_45942,N_41435);
nand UO_74 (O_74,N_48216,N_43897);
xnor UO_75 (O_75,N_42577,N_46558);
or UO_76 (O_76,N_41767,N_43020);
nor UO_77 (O_77,N_40098,N_43477);
and UO_78 (O_78,N_40823,N_49398);
and UO_79 (O_79,N_41506,N_48312);
nor UO_80 (O_80,N_49485,N_48840);
xnor UO_81 (O_81,N_48622,N_43718);
nor UO_82 (O_82,N_48148,N_48361);
nand UO_83 (O_83,N_46338,N_49447);
xor UO_84 (O_84,N_43816,N_40671);
nor UO_85 (O_85,N_41961,N_42667);
nor UO_86 (O_86,N_40389,N_40785);
nand UO_87 (O_87,N_42572,N_45095);
xnor UO_88 (O_88,N_44142,N_40309);
and UO_89 (O_89,N_49284,N_48531);
xor UO_90 (O_90,N_41295,N_45304);
or UO_91 (O_91,N_44122,N_42987);
and UO_92 (O_92,N_46760,N_45667);
nor UO_93 (O_93,N_43151,N_47043);
or UO_94 (O_94,N_41137,N_46003);
nand UO_95 (O_95,N_47124,N_40106);
and UO_96 (O_96,N_42021,N_46417);
nor UO_97 (O_97,N_41737,N_46596);
nand UO_98 (O_98,N_43971,N_42827);
nor UO_99 (O_99,N_42096,N_48659);
nor UO_100 (O_100,N_48561,N_43470);
and UO_101 (O_101,N_40220,N_46339);
xor UO_102 (O_102,N_49156,N_47007);
xor UO_103 (O_103,N_46734,N_47199);
and UO_104 (O_104,N_42790,N_47139);
xor UO_105 (O_105,N_43430,N_48845);
nor UO_106 (O_106,N_49690,N_49625);
xor UO_107 (O_107,N_47479,N_41934);
xor UO_108 (O_108,N_48113,N_40094);
nor UO_109 (O_109,N_41714,N_44443);
or UO_110 (O_110,N_46279,N_46441);
xnor UO_111 (O_111,N_48174,N_49203);
nor UO_112 (O_112,N_45982,N_40626);
xor UO_113 (O_113,N_41136,N_45146);
xnor UO_114 (O_114,N_47424,N_41696);
nor UO_115 (O_115,N_44963,N_48494);
xor UO_116 (O_116,N_41959,N_43507);
nor UO_117 (O_117,N_44373,N_40804);
and UO_118 (O_118,N_49991,N_48227);
xnor UO_119 (O_119,N_44127,N_41417);
nor UO_120 (O_120,N_40034,N_49514);
nand UO_121 (O_121,N_43252,N_44238);
nor UO_122 (O_122,N_41885,N_45839);
or UO_123 (O_123,N_48796,N_44009);
nor UO_124 (O_124,N_41870,N_43370);
or UO_125 (O_125,N_40784,N_40663);
or UO_126 (O_126,N_46459,N_40864);
nor UO_127 (O_127,N_43058,N_40623);
and UO_128 (O_128,N_49071,N_47496);
xor UO_129 (O_129,N_44018,N_45727);
and UO_130 (O_130,N_42280,N_41884);
and UO_131 (O_131,N_42832,N_41778);
or UO_132 (O_132,N_47046,N_49258);
nor UO_133 (O_133,N_42848,N_40121);
nand UO_134 (O_134,N_42009,N_43156);
nand UO_135 (O_135,N_43451,N_40568);
or UO_136 (O_136,N_40291,N_45970);
nor UO_137 (O_137,N_44894,N_41586);
and UO_138 (O_138,N_40246,N_49509);
and UO_139 (O_139,N_49764,N_48588);
nand UO_140 (O_140,N_47018,N_44223);
xnor UO_141 (O_141,N_41279,N_46885);
nor UO_142 (O_142,N_40680,N_41265);
nor UO_143 (O_143,N_43070,N_45567);
xnor UO_144 (O_144,N_48534,N_47246);
xnor UO_145 (O_145,N_46645,N_46130);
nand UO_146 (O_146,N_46684,N_43371);
nand UO_147 (O_147,N_43413,N_40496);
nand UO_148 (O_148,N_49235,N_46141);
and UO_149 (O_149,N_48605,N_44278);
or UO_150 (O_150,N_41469,N_46763);
nor UO_151 (O_151,N_40004,N_49667);
and UO_152 (O_152,N_49252,N_46103);
xor UO_153 (O_153,N_45305,N_41851);
xnor UO_154 (O_154,N_41346,N_49129);
and UO_155 (O_155,N_40005,N_45930);
xnor UO_156 (O_156,N_45206,N_47791);
and UO_157 (O_157,N_47473,N_40381);
nand UO_158 (O_158,N_42729,N_44441);
nor UO_159 (O_159,N_46065,N_42998);
nand UO_160 (O_160,N_45228,N_42918);
or UO_161 (O_161,N_42432,N_41250);
and UO_162 (O_162,N_41660,N_49705);
nor UO_163 (O_163,N_49355,N_46863);
nor UO_164 (O_164,N_46328,N_45684);
nand UO_165 (O_165,N_43355,N_42121);
nor UO_166 (O_166,N_43796,N_45489);
or UO_167 (O_167,N_40155,N_43386);
nand UO_168 (O_168,N_44212,N_46968);
xor UO_169 (O_169,N_49401,N_42072);
xnor UO_170 (O_170,N_45669,N_43431);
nand UO_171 (O_171,N_48853,N_46131);
or UO_172 (O_172,N_49886,N_40150);
and UO_173 (O_173,N_48748,N_43429);
xor UO_174 (O_174,N_45525,N_46648);
xor UO_175 (O_175,N_43561,N_48817);
xnor UO_176 (O_176,N_49316,N_40024);
or UO_177 (O_177,N_48180,N_41434);
xnor UO_178 (O_178,N_42307,N_46292);
or UO_179 (O_179,N_47841,N_48145);
and UO_180 (O_180,N_42725,N_47513);
or UO_181 (O_181,N_49775,N_45301);
and UO_182 (O_182,N_42006,N_49651);
and UO_183 (O_183,N_41128,N_44467);
xnor UO_184 (O_184,N_48545,N_41757);
and UO_185 (O_185,N_45874,N_49973);
xnor UO_186 (O_186,N_43590,N_41794);
nand UO_187 (O_187,N_40701,N_41518);
nand UO_188 (O_188,N_49839,N_42246);
nor UO_189 (O_189,N_48291,N_49826);
nand UO_190 (O_190,N_46206,N_44437);
xor UO_191 (O_191,N_49281,N_40257);
nor UO_192 (O_192,N_43069,N_43683);
nor UO_193 (O_193,N_40739,N_48429);
nand UO_194 (O_194,N_47497,N_49917);
nand UO_195 (O_195,N_40048,N_45786);
or UO_196 (O_196,N_46939,N_44339);
or UO_197 (O_197,N_46644,N_40641);
or UO_198 (O_198,N_47416,N_47089);
nand UO_199 (O_199,N_44218,N_44959);
or UO_200 (O_200,N_48344,N_43062);
nor UO_201 (O_201,N_49282,N_45165);
nand UO_202 (O_202,N_48844,N_45425);
nand UO_203 (O_203,N_49456,N_41410);
or UO_204 (O_204,N_47950,N_43652);
and UO_205 (O_205,N_48527,N_48354);
or UO_206 (O_206,N_46910,N_46403);
and UO_207 (O_207,N_48186,N_42919);
xnor UO_208 (O_208,N_40541,N_47332);
nor UO_209 (O_209,N_45779,N_43742);
nor UO_210 (O_210,N_44667,N_45385);
or UO_211 (O_211,N_43792,N_40225);
nor UO_212 (O_212,N_47681,N_49773);
nand UO_213 (O_213,N_44906,N_40915);
and UO_214 (O_214,N_40311,N_49923);
or UO_215 (O_215,N_47666,N_40352);
nand UO_216 (O_216,N_43516,N_44439);
nand UO_217 (O_217,N_49116,N_49726);
nor UO_218 (O_218,N_47422,N_41678);
and UO_219 (O_219,N_48956,N_47847);
xor UO_220 (O_220,N_46210,N_45148);
and UO_221 (O_221,N_41997,N_41613);
or UO_222 (O_222,N_44322,N_45998);
xor UO_223 (O_223,N_43949,N_40921);
nand UO_224 (O_224,N_44501,N_41647);
nor UO_225 (O_225,N_41713,N_46211);
and UO_226 (O_226,N_48203,N_42361);
xor UO_227 (O_227,N_46147,N_40022);
nand UO_228 (O_228,N_44341,N_49094);
xnor UO_229 (O_229,N_41652,N_41088);
or UO_230 (O_230,N_46543,N_47689);
or UO_231 (O_231,N_47337,N_47340);
xor UO_232 (O_232,N_49050,N_48266);
nor UO_233 (O_233,N_41705,N_47739);
nor UO_234 (O_234,N_45946,N_41217);
xor UO_235 (O_235,N_45676,N_47492);
nor UO_236 (O_236,N_45989,N_43807);
xor UO_237 (O_237,N_44287,N_46025);
xor UO_238 (O_238,N_41760,N_44440);
xor UO_239 (O_239,N_43562,N_44048);
nand UO_240 (O_240,N_49961,N_40718);
nor UO_241 (O_241,N_41658,N_44862);
and UO_242 (O_242,N_48977,N_43342);
xnor UO_243 (O_243,N_42933,N_47152);
xor UO_244 (O_244,N_42260,N_41228);
and UO_245 (O_245,N_48637,N_41569);
or UO_246 (O_246,N_46392,N_45109);
xor UO_247 (O_247,N_47128,N_44343);
xor UO_248 (O_248,N_44252,N_45064);
nand UO_249 (O_249,N_49935,N_41723);
nor UO_250 (O_250,N_48394,N_48386);
nand UO_251 (O_251,N_48525,N_42516);
nor UO_252 (O_252,N_40191,N_40971);
nand UO_253 (O_253,N_45414,N_45155);
nand UO_254 (O_254,N_46945,N_40833);
xnor UO_255 (O_255,N_45149,N_43110);
nor UO_256 (O_256,N_40614,N_44586);
xnor UO_257 (O_257,N_45108,N_41966);
and UO_258 (O_258,N_40282,N_48517);
xnor UO_259 (O_259,N_48787,N_46432);
and UO_260 (O_260,N_49925,N_47501);
and UO_261 (O_261,N_47583,N_43075);
and UO_262 (O_262,N_47247,N_46401);
or UO_263 (O_263,N_47395,N_49580);
nand UO_264 (O_264,N_45466,N_46109);
nor UO_265 (O_265,N_46256,N_48319);
nand UO_266 (O_266,N_42198,N_40194);
xor UO_267 (O_267,N_40930,N_49617);
nand UO_268 (O_268,N_45313,N_45352);
or UO_269 (O_269,N_41474,N_41283);
xnor UO_270 (O_270,N_49997,N_43390);
nor UO_271 (O_271,N_45001,N_41130);
nand UO_272 (O_272,N_43818,N_44742);
nand UO_273 (O_273,N_44309,N_47462);
and UO_274 (O_274,N_41880,N_45390);
nor UO_275 (O_275,N_45871,N_43400);
or UO_276 (O_276,N_43489,N_40876);
nor UO_277 (O_277,N_44685,N_47161);
and UO_278 (O_278,N_42371,N_48812);
and UO_279 (O_279,N_43501,N_46611);
xor UO_280 (O_280,N_44548,N_48478);
and UO_281 (O_281,N_46132,N_48360);
xnor UO_282 (O_282,N_42589,N_40416);
xor UO_283 (O_283,N_42302,N_42395);
xnor UO_284 (O_284,N_45721,N_48761);
xor UO_285 (O_285,N_49658,N_45560);
nand UO_286 (O_286,N_44325,N_41132);
or UO_287 (O_287,N_40516,N_48431);
nor UO_288 (O_288,N_41095,N_49957);
nand UO_289 (O_289,N_49654,N_49965);
or UO_290 (O_290,N_46124,N_40749);
nor UO_291 (O_291,N_41267,N_43523);
or UO_292 (O_292,N_41914,N_40440);
xnor UO_293 (O_293,N_42561,N_41724);
nand UO_294 (O_294,N_44762,N_48719);
or UO_295 (O_295,N_47646,N_43613);
and UO_296 (O_296,N_40333,N_40115);
and UO_297 (O_297,N_49783,N_41837);
nor UO_298 (O_298,N_46212,N_48711);
xnor UO_299 (O_299,N_40454,N_42124);
and UO_300 (O_300,N_43222,N_48419);
nor UO_301 (O_301,N_44353,N_47721);
or UO_302 (O_302,N_48795,N_43705);
nor UO_303 (O_303,N_49150,N_43077);
and UO_304 (O_304,N_45972,N_42607);
nand UO_305 (O_305,N_41030,N_42999);
nand UO_306 (O_306,N_41353,N_49739);
or UO_307 (O_307,N_43436,N_40838);
nor UO_308 (O_308,N_43254,N_46613);
xor UO_309 (O_309,N_42496,N_48648);
nor UO_310 (O_310,N_44002,N_43977);
or UO_311 (O_311,N_44391,N_41994);
or UO_312 (O_312,N_46531,N_46208);
and UO_313 (O_313,N_47218,N_48393);
and UO_314 (O_314,N_42031,N_40125);
xnor UO_315 (O_315,N_48348,N_46080);
xor UO_316 (O_316,N_42671,N_43831);
nor UO_317 (O_317,N_49732,N_46357);
or UO_318 (O_318,N_48677,N_46873);
nor UO_319 (O_319,N_44691,N_46033);
nand UO_320 (O_320,N_45944,N_40528);
nand UO_321 (O_321,N_49426,N_40062);
and UO_322 (O_322,N_41350,N_45298);
xnor UO_323 (O_323,N_42167,N_47323);
and UO_324 (O_324,N_41588,N_45921);
and UO_325 (O_325,N_48582,N_46845);
or UO_326 (O_326,N_42265,N_49397);
and UO_327 (O_327,N_44527,N_40636);
nand UO_328 (O_328,N_43969,N_46302);
nand UO_329 (O_329,N_47939,N_42878);
nor UO_330 (O_330,N_49104,N_48882);
or UO_331 (O_331,N_43951,N_40321);
xnor UO_332 (O_332,N_48978,N_44715);
nand UO_333 (O_333,N_46469,N_45620);
nor UO_334 (O_334,N_43822,N_44173);
xor UO_335 (O_335,N_41929,N_44964);
xor UO_336 (O_336,N_41960,N_43617);
nand UO_337 (O_337,N_49537,N_42764);
or UO_338 (O_338,N_43310,N_40806);
xnor UO_339 (O_339,N_42957,N_48427);
nor UO_340 (O_340,N_45285,N_41415);
nor UO_341 (O_341,N_46694,N_47927);
nand UO_342 (O_342,N_45925,N_46126);
and UO_343 (O_343,N_44793,N_49010);
and UO_344 (O_344,N_42346,N_42378);
xnor UO_345 (O_345,N_49868,N_46673);
nand UO_346 (O_346,N_42883,N_46060);
nand UO_347 (O_347,N_42882,N_41319);
xnor UO_348 (O_348,N_42931,N_40430);
nor UO_349 (O_349,N_46841,N_43934);
nand UO_350 (O_350,N_42842,N_43698);
nand UO_351 (O_351,N_45975,N_46796);
and UO_352 (O_352,N_44180,N_47085);
and UO_353 (O_353,N_47398,N_40402);
xnor UO_354 (O_354,N_44610,N_40145);
nor UO_355 (O_355,N_46638,N_41742);
and UO_356 (O_356,N_47115,N_44492);
xnor UO_357 (O_357,N_40283,N_40772);
nor UO_358 (O_358,N_41286,N_47499);
xnor UO_359 (O_359,N_45476,N_42812);
nor UO_360 (O_360,N_48104,N_48586);
xnor UO_361 (O_361,N_47077,N_49612);
nand UO_362 (O_362,N_48320,N_44929);
and UO_363 (O_363,N_43763,N_45123);
nor UO_364 (O_364,N_43495,N_41911);
or UO_365 (O_365,N_41318,N_40845);
and UO_366 (O_366,N_41974,N_48678);
nor UO_367 (O_367,N_42180,N_40134);
or UO_368 (O_368,N_41863,N_41933);
nand UO_369 (O_369,N_48265,N_43601);
and UO_370 (O_370,N_42161,N_43502);
nand UO_371 (O_371,N_45565,N_41094);
nand UO_372 (O_372,N_43553,N_40375);
and UO_373 (O_373,N_44045,N_42118);
nor UO_374 (O_374,N_45900,N_49268);
xnor UO_375 (O_375,N_48165,N_43106);
nor UO_376 (O_376,N_45494,N_44799);
nor UO_377 (O_377,N_43088,N_40944);
nand UO_378 (O_378,N_40289,N_42801);
and UO_379 (O_379,N_43434,N_49662);
or UO_380 (O_380,N_41601,N_43910);
nor UO_381 (O_381,N_45910,N_40305);
and UO_382 (O_382,N_45954,N_40172);
and UO_383 (O_383,N_40198,N_40387);
xnor UO_384 (O_384,N_43506,N_49055);
or UO_385 (O_385,N_44794,N_49440);
nor UO_386 (O_386,N_41198,N_46642);
and UO_387 (O_387,N_46405,N_42774);
and UO_388 (O_388,N_47862,N_41873);
or UO_389 (O_389,N_48182,N_49367);
or UO_390 (O_390,N_44810,N_49360);
and UO_391 (O_391,N_47286,N_44461);
nor UO_392 (O_392,N_48797,N_44747);
and UO_393 (O_393,N_46426,N_49200);
xor UO_394 (O_394,N_48595,N_41395);
nor UO_395 (O_395,N_48405,N_44999);
or UO_396 (O_396,N_46846,N_44328);
nand UO_397 (O_397,N_45844,N_40977);
and UO_398 (O_398,N_44901,N_44696);
or UO_399 (O_399,N_40835,N_47904);
xor UO_400 (O_400,N_40312,N_45100);
xor UO_401 (O_401,N_45470,N_40193);
nor UO_402 (O_402,N_49901,N_46385);
and UO_403 (O_403,N_49309,N_49986);
xor UO_404 (O_404,N_48773,N_40510);
or UO_405 (O_405,N_48157,N_49417);
and UO_406 (O_406,N_41042,N_47508);
and UO_407 (O_407,N_44875,N_44458);
and UO_408 (O_408,N_44323,N_41572);
and UO_409 (O_409,N_49405,N_48957);
or UO_410 (O_410,N_47980,N_47532);
and UO_411 (O_411,N_43024,N_41962);
and UO_412 (O_412,N_44512,N_47676);
nor UO_413 (O_413,N_48069,N_48336);
nor UO_414 (O_414,N_43820,N_46599);
xnor UO_415 (O_415,N_43804,N_46979);
nor UO_416 (O_416,N_47835,N_47546);
nor UO_417 (O_417,N_45022,N_45950);
or UO_418 (O_418,N_42558,N_45703);
xnor UO_419 (O_419,N_48376,N_47790);
xor UO_420 (O_420,N_41551,N_41796);
and UO_421 (O_421,N_46566,N_48967);
nor UO_422 (O_422,N_42550,N_46398);
nand UO_423 (O_423,N_40859,N_48865);
nor UO_424 (O_424,N_43122,N_47551);
xor UO_425 (O_425,N_42670,N_44583);
and UO_426 (O_426,N_43673,N_47470);
nor UO_427 (O_427,N_40315,N_47641);
or UO_428 (O_428,N_44874,N_44593);
xor UO_429 (O_429,N_41202,N_43900);
xor UO_430 (O_430,N_40162,N_42416);
nor UO_431 (O_431,N_45736,N_45651);
xnor UO_432 (O_432,N_48068,N_45314);
and UO_433 (O_433,N_45734,N_41244);
xor UO_434 (O_434,N_46413,N_41045);
and UO_435 (O_435,N_45086,N_42387);
nor UO_436 (O_436,N_44481,N_46275);
xnor UO_437 (O_437,N_47617,N_49076);
xor UO_438 (O_438,N_40975,N_44159);
nor UO_439 (O_439,N_44395,N_40501);
or UO_440 (O_440,N_43009,N_44326);
nand UO_441 (O_441,N_44188,N_48655);
xnor UO_442 (O_442,N_48700,N_43650);
nor UO_443 (O_443,N_42544,N_42174);
xor UO_444 (O_444,N_41151,N_49984);
xnor UO_445 (O_445,N_44637,N_42681);
nor UO_446 (O_446,N_48099,N_47691);
and UO_447 (O_447,N_41816,N_49444);
xor UO_448 (O_448,N_43779,N_41928);
and UO_449 (O_449,N_43493,N_43903);
nor UO_450 (O_450,N_45564,N_43060);
or UO_451 (O_451,N_42983,N_47491);
xor UO_452 (O_452,N_42741,N_45034);
xor UO_453 (O_453,N_44296,N_43684);
and UO_454 (O_454,N_43678,N_49911);
nor UO_455 (O_455,N_45723,N_47030);
nand UO_456 (O_456,N_49494,N_45202);
xor UO_457 (O_457,N_40295,N_41858);
xnor UO_458 (O_458,N_42892,N_48495);
xnor UO_459 (O_459,N_48725,N_45653);
xnor UO_460 (O_460,N_47142,N_45914);
xnor UO_461 (O_461,N_49766,N_45321);
nor UO_462 (O_462,N_40451,N_40133);
nand UO_463 (O_463,N_41232,N_44888);
nand UO_464 (O_464,N_47949,N_46114);
or UO_465 (O_465,N_44152,N_44352);
nor UO_466 (O_466,N_41908,N_45908);
xor UO_467 (O_467,N_48734,N_45290);
nand UO_468 (O_468,N_49269,N_44498);
nor UO_469 (O_469,N_49208,N_44735);
or UO_470 (O_470,N_41508,N_49413);
xnor UO_471 (O_471,N_47243,N_42247);
nand UO_472 (O_472,N_44460,N_44262);
nand UO_473 (O_473,N_47278,N_46349);
nand UO_474 (O_474,N_48019,N_40775);
xor UO_475 (O_475,N_45329,N_46180);
nand UO_476 (O_476,N_40367,N_43455);
xor UO_477 (O_477,N_41637,N_48553);
xnor UO_478 (O_478,N_47683,N_42904);
or UO_479 (O_479,N_49280,N_42769);
xor UO_480 (O_480,N_49409,N_43886);
xor UO_481 (O_481,N_42792,N_45945);
xnor UO_482 (O_482,N_43496,N_42492);
or UO_483 (O_483,N_40588,N_45846);
nor UO_484 (O_484,N_44050,N_49263);
or UO_485 (O_485,N_42746,N_49382);
and UO_486 (O_486,N_49803,N_48116);
nor UO_487 (O_487,N_47934,N_46537);
or UO_488 (O_488,N_43427,N_45306);
and UO_489 (O_489,N_49758,N_46585);
nand UO_490 (O_490,N_40654,N_46711);
nor UO_491 (O_491,N_47754,N_43819);
nand UO_492 (O_492,N_41877,N_48022);
nor UO_493 (O_493,N_44197,N_48201);
or UO_494 (O_494,N_46410,N_44387);
xnor UO_495 (O_495,N_49013,N_47592);
and UO_496 (O_496,N_45880,N_42109);
nor UO_497 (O_497,N_48277,N_46356);
and UO_498 (O_498,N_40043,N_48417);
xor UO_499 (O_499,N_44927,N_48256);
xnor UO_500 (O_500,N_43757,N_43793);
and UO_501 (O_501,N_44949,N_40638);
xnor UO_502 (O_502,N_47114,N_40712);
nor UO_503 (O_503,N_47425,N_40032);
nor UO_504 (O_504,N_47849,N_47778);
nand UO_505 (O_505,N_41105,N_44843);
and UO_506 (O_506,N_42909,N_46709);
nand UO_507 (O_507,N_45357,N_45084);
or UO_508 (O_508,N_42949,N_43898);
nor UO_509 (O_509,N_44051,N_46187);
nor UO_510 (O_510,N_42171,N_43000);
and UO_511 (O_511,N_44733,N_41401);
and UO_512 (O_512,N_41302,N_43269);
xor UO_513 (O_513,N_49696,N_48581);
or UO_514 (O_514,N_40059,N_41703);
and UO_515 (O_515,N_40374,N_41538);
or UO_516 (O_516,N_44237,N_47020);
nor UO_517 (O_517,N_47866,N_42207);
or UO_518 (O_518,N_47565,N_46564);
and UO_519 (O_519,N_47705,N_47304);
nor UO_520 (O_520,N_44543,N_49647);
and UO_521 (O_521,N_45127,N_42011);
xor UO_522 (O_522,N_42078,N_43557);
or UO_523 (O_523,N_40625,N_47380);
and UO_524 (O_524,N_49428,N_43103);
nor UO_525 (O_525,N_41986,N_42144);
nor UO_526 (O_526,N_47952,N_41623);
and UO_527 (O_527,N_46964,N_48824);
and UO_528 (O_528,N_46012,N_43513);
xnor UO_529 (O_529,N_41197,N_43713);
nor UO_530 (O_530,N_45718,N_47621);
or UO_531 (O_531,N_48308,N_42798);
nor UO_532 (O_532,N_43243,N_40467);
and UO_533 (O_533,N_44084,N_43795);
nand UO_534 (O_534,N_48556,N_49210);
xnor UO_535 (O_535,N_47153,N_48960);
nand UO_536 (O_536,N_40347,N_41051);
nor UO_537 (O_537,N_48672,N_49025);
nand UO_538 (O_538,N_45337,N_42581);
nand UO_539 (O_539,N_41513,N_45196);
or UO_540 (O_540,N_45184,N_43926);
nand UO_541 (O_541,N_46038,N_48663);
or UO_542 (O_542,N_42810,N_48854);
and UO_543 (O_543,N_49340,N_41470);
xor UO_544 (O_544,N_46295,N_40970);
nor UO_545 (O_545,N_44179,N_46972);
nor UO_546 (O_546,N_48804,N_47227);
nand UO_547 (O_547,N_49715,N_45728);
and UO_548 (O_548,N_46318,N_47907);
xor UO_549 (O_549,N_47585,N_41383);
and UO_550 (O_550,N_48503,N_46904);
or UO_551 (O_551,N_49220,N_46000);
xor UO_552 (O_552,N_45744,N_42173);
nor UO_553 (O_553,N_48215,N_49898);
nand UO_554 (O_554,N_40941,N_47931);
and UO_555 (O_555,N_48929,N_41304);
or UO_556 (O_556,N_45464,N_48018);
nand UO_557 (O_557,N_40856,N_48591);
xnor UO_558 (O_558,N_43641,N_41412);
xnor UO_559 (O_559,N_40007,N_49663);
nor UO_560 (O_560,N_41409,N_41688);
and UO_561 (O_561,N_43084,N_43653);
and UO_562 (O_562,N_48350,N_43865);
xnor UO_563 (O_563,N_48996,N_48138);
xnor UO_564 (O_564,N_47553,N_43207);
xor UO_565 (O_565,N_48645,N_46553);
nor UO_566 (O_566,N_43339,N_45490);
nand UO_567 (O_567,N_46818,N_45956);
nor UO_568 (O_568,N_48964,N_49553);
xnor UO_569 (O_569,N_44571,N_42329);
and UO_570 (O_570,N_46829,N_45791);
and UO_571 (O_571,N_42944,N_48543);
xnor UO_572 (O_572,N_46927,N_46023);
nor UO_573 (O_573,N_49038,N_45045);
nand UO_574 (O_574,N_43550,N_42534);
nor UO_575 (O_575,N_44101,N_47351);
or UO_576 (O_576,N_41773,N_43605);
xnor UO_577 (O_577,N_48643,N_47257);
and UO_578 (O_578,N_41213,N_40782);
xor UO_579 (O_579,N_40721,N_44947);
nand UO_580 (O_580,N_41615,N_48183);
nor UO_581 (O_581,N_49515,N_49684);
nand UO_582 (O_582,N_45941,N_41664);
and UO_583 (O_583,N_42279,N_43878);
nand UO_584 (O_584,N_40353,N_48511);
xor UO_585 (O_585,N_41721,N_45832);
nor UO_586 (O_586,N_48131,N_45081);
nor UO_587 (O_587,N_46358,N_41315);
xnor UO_588 (O_588,N_47076,N_47378);
or UO_589 (O_589,N_47645,N_44471);
xor UO_590 (O_590,N_49634,N_48806);
nor UO_591 (O_591,N_42794,N_42320);
and UO_592 (O_592,N_45961,N_40660);
xor UO_593 (O_593,N_47531,N_45143);
nor UO_594 (O_594,N_47764,N_41203);
and UO_595 (O_595,N_42219,N_43130);
xor UO_596 (O_596,N_41840,N_49279);
nor UO_597 (O_597,N_43860,N_48910);
or UO_598 (O_598,N_47765,N_48392);
nand UO_599 (O_599,N_42023,N_47397);
and UO_600 (O_600,N_47578,N_48580);
and UO_601 (O_601,N_49479,N_43581);
and UO_602 (O_602,N_49670,N_48850);
and UO_603 (O_603,N_47977,N_46175);
and UO_604 (O_604,N_45829,N_41352);
and UO_605 (O_605,N_45467,N_40476);
nor UO_606 (O_606,N_45053,N_45719);
and UO_607 (O_607,N_40727,N_42196);
nor UO_608 (O_608,N_40961,N_49633);
nor UO_609 (O_609,N_40637,N_44021);
xor UO_610 (O_610,N_44090,N_41651);
nand UO_611 (O_611,N_43338,N_49334);
or UO_612 (O_612,N_40991,N_48056);
nor UO_613 (O_613,N_48382,N_46627);
and UO_614 (O_614,N_47784,N_40208);
or UO_615 (O_615,N_43064,N_41686);
nand UO_616 (O_616,N_42711,N_44082);
nand UO_617 (O_617,N_41822,N_49148);
and UO_618 (O_618,N_49278,N_40627);
and UO_619 (O_619,N_45236,N_42407);
or UO_620 (O_620,N_49934,N_48254);
or UO_621 (O_621,N_40351,N_47879);
nand UO_622 (O_622,N_46728,N_46161);
nor UO_623 (O_623,N_43169,N_49788);
nand UO_624 (O_624,N_43978,N_46164);
or UO_625 (O_625,N_43097,N_41391);
xor UO_626 (O_626,N_42615,N_43535);
or UO_627 (O_627,N_42584,N_40204);
nor UO_628 (O_628,N_46182,N_43001);
nand UO_629 (O_629,N_49324,N_49870);
xnor UO_630 (O_630,N_40673,N_43574);
and UO_631 (O_631,N_45558,N_46353);
or UO_632 (O_632,N_49889,N_48708);
nor UO_633 (O_633,N_40453,N_48597);
and UO_634 (O_634,N_49061,N_43994);
or UO_635 (O_635,N_40651,N_48999);
xor UO_636 (O_636,N_47929,N_49712);
nand UO_637 (O_637,N_44627,N_47959);
nor UO_638 (O_638,N_49169,N_41930);
or UO_639 (O_639,N_47864,N_44786);
xor UO_640 (O_640,N_44030,N_48414);
and UO_641 (O_641,N_42722,N_42692);
or UO_642 (O_642,N_42102,N_46982);
nand UO_643 (O_643,N_43234,N_42483);
or UO_644 (O_644,N_43834,N_41835);
xnor UO_645 (O_645,N_43902,N_49586);
or UO_646 (O_646,N_43866,N_40951);
xor UO_647 (O_647,N_49073,N_45741);
or UO_648 (O_648,N_47094,N_49037);
or UO_649 (O_649,N_46730,N_49691);
or UO_650 (O_650,N_45689,N_43531);
and UO_651 (O_651,N_47321,N_43419);
nor UO_652 (O_652,N_49018,N_45088);
xnor UO_653 (O_653,N_44243,N_44930);
or UO_654 (O_654,N_49217,N_48587);
nand UO_655 (O_655,N_40558,N_41238);
xnor UO_656 (O_656,N_42977,N_48689);
and UO_657 (O_657,N_43462,N_41817);
xor UO_658 (O_658,N_49608,N_42037);
nor UO_659 (O_659,N_49604,N_48261);
and UO_660 (O_660,N_45983,N_41299);
nor UO_661 (O_661,N_47644,N_42879);
and UO_662 (O_662,N_49801,N_45847);
or UO_663 (O_663,N_40773,N_46949);
or UO_664 (O_664,N_49837,N_49668);
xnor UO_665 (O_665,N_43249,N_49242);
or UO_666 (O_666,N_45500,N_42352);
xnor UO_667 (O_667,N_49865,N_42940);
nand UO_668 (O_668,N_44438,N_49103);
and UO_669 (O_669,N_44890,N_42438);
nor UO_670 (O_670,N_42923,N_47634);
or UO_671 (O_671,N_46928,N_42762);
nand UO_672 (O_672,N_40793,N_44074);
or UO_673 (O_673,N_45246,N_42458);
and UO_674 (O_674,N_43519,N_49070);
and UO_675 (O_675,N_41495,N_48447);
or UO_676 (O_676,N_49824,N_44835);
or UO_677 (O_677,N_49455,N_43196);
nor UO_678 (O_678,N_48328,N_46860);
nor UO_679 (O_679,N_46359,N_45003);
or UO_680 (O_680,N_41749,N_40732);
nand UO_681 (O_681,N_48943,N_45250);
xnor UO_682 (O_682,N_45214,N_42528);
or UO_683 (O_683,N_40399,N_40154);
or UO_684 (O_684,N_46277,N_48502);
and UO_685 (O_685,N_49026,N_47041);
xnor UO_686 (O_686,N_41779,N_41195);
nand UO_687 (O_687,N_42934,N_49113);
or UO_688 (O_688,N_41511,N_44028);
and UO_689 (O_689,N_49044,N_44775);
nand UO_690 (O_690,N_42975,N_41022);
and UO_691 (O_691,N_47755,N_41740);
or UO_692 (O_692,N_40912,N_45642);
xor UO_693 (O_693,N_44091,N_41983);
and UO_694 (O_694,N_45563,N_40596);
nand UO_695 (O_695,N_41990,N_42319);
and UO_696 (O_696,N_47579,N_46427);
xor UO_697 (O_697,N_43671,N_42222);
xnor UO_698 (O_698,N_46878,N_45090);
or UO_699 (O_699,N_45597,N_41440);
and UO_700 (O_700,N_44468,N_45753);
nor UO_701 (O_701,N_44800,N_48317);
nand UO_702 (O_702,N_46978,N_47832);
nor UO_703 (O_703,N_46591,N_47828);
or UO_704 (O_704,N_44604,N_49543);
and UO_705 (O_705,N_43287,N_46938);
xor UO_706 (O_706,N_42554,N_41301);
nor UO_707 (O_707,N_42200,N_45367);
and UO_708 (O_708,N_46776,N_46196);
nor UO_709 (O_709,N_44705,N_44631);
xor UO_710 (O_710,N_47469,N_42253);
nor UO_711 (O_711,N_49285,N_41888);
or UO_712 (O_712,N_47600,N_43346);
and UO_713 (O_713,N_46081,N_44950);
nand UO_714 (O_714,N_45809,N_48398);
nor UO_715 (O_715,N_49059,N_41476);
nand UO_716 (O_716,N_48514,N_42327);
nand UO_717 (O_717,N_47517,N_48792);
xor UO_718 (O_718,N_47178,N_49504);
and UO_719 (O_719,N_45798,N_43883);
xor UO_720 (O_720,N_43263,N_43711);
nor UO_721 (O_721,N_42134,N_41579);
and UO_722 (O_722,N_46918,N_47825);
nor UO_723 (O_723,N_41679,N_49759);
and UO_724 (O_724,N_49949,N_41512);
or UO_725 (O_725,N_42551,N_46871);
nand UO_726 (O_726,N_49630,N_46842);
nand UO_727 (O_727,N_46572,N_47675);
nor UO_728 (O_728,N_48949,N_42707);
or UO_729 (O_729,N_43676,N_42693);
and UO_730 (O_730,N_41099,N_46544);
and UO_731 (O_731,N_47031,N_46119);
or UO_732 (O_732,N_48086,N_40815);
xnor UO_733 (O_733,N_48306,N_40140);
nand UO_734 (O_734,N_42168,N_42178);
nand UO_735 (O_735,N_45661,N_41193);
and UO_736 (O_736,N_43937,N_42342);
and UO_737 (O_737,N_41158,N_40271);
and UO_738 (O_738,N_43090,N_49536);
nor UO_739 (O_739,N_42152,N_40526);
nor UO_740 (O_740,N_41861,N_45516);
nor UO_741 (O_741,N_47026,N_43312);
nor UO_742 (O_742,N_42424,N_47215);
nor UO_743 (O_743,N_45804,N_40195);
nand UO_744 (O_744,N_48687,N_48292);
or UO_745 (O_745,N_48346,N_47401);
and UO_746 (O_746,N_49915,N_47305);
xnor UO_747 (O_747,N_43025,N_40016);
nor UO_748 (O_748,N_41642,N_49468);
and UO_749 (O_749,N_44880,N_48716);
or UO_750 (O_750,N_44530,N_45951);
nor UO_751 (O_751,N_43260,N_42549);
and UO_752 (O_752,N_47767,N_45455);
and UO_753 (O_753,N_42429,N_47342);
and UO_754 (O_754,N_42136,N_48746);
nand UO_755 (O_755,N_41079,N_47965);
nand UO_756 (O_756,N_40227,N_47694);
nand UO_757 (O_757,N_40667,N_45231);
and UO_758 (O_758,N_41611,N_40503);
nor UO_759 (O_759,N_43662,N_48992);
nand UO_760 (O_760,N_44430,N_47780);
nor UO_761 (O_761,N_41754,N_42742);
or UO_762 (O_762,N_46281,N_46569);
xnor UO_763 (O_763,N_46856,N_44661);
nand UO_764 (O_764,N_44726,N_49247);
and UO_765 (O_765,N_41114,N_49386);
nor UO_766 (O_766,N_46600,N_45172);
nor UO_767 (O_767,N_49218,N_40947);
and UO_768 (O_768,N_41117,N_49004);
xnor UO_769 (O_769,N_42417,N_48178);
nand UO_770 (O_770,N_42449,N_48089);
nand UO_771 (O_771,N_46423,N_40792);
nand UO_772 (O_772,N_40030,N_42761);
or UO_773 (O_773,N_45785,N_47010);
nor UO_774 (O_774,N_45662,N_49351);
xnor UO_775 (O_775,N_44566,N_47024);
nor UO_776 (O_776,N_44815,N_42829);
nor UO_777 (O_777,N_40053,N_43172);
nor UO_778 (O_778,N_45918,N_40828);
nor UO_779 (O_779,N_49721,N_40794);
or UO_780 (O_780,N_44257,N_41691);
and UO_781 (O_781,N_40662,N_43255);
and UO_782 (O_782,N_48271,N_43232);
and UO_783 (O_783,N_48075,N_47320);
xnor UO_784 (O_784,N_40743,N_43826);
xor UO_785 (O_785,N_46953,N_45079);
nor UO_786 (O_786,N_43944,N_40746);
and UO_787 (O_787,N_43670,N_41663);
and UO_788 (O_788,N_47774,N_48323);
or UO_789 (O_789,N_47576,N_45907);
and UO_790 (O_790,N_40585,N_43615);
nor UO_791 (O_791,N_46016,N_46909);
xnor UO_792 (O_792,N_48297,N_46958);
nor UO_793 (O_793,N_41168,N_43998);
nor UO_794 (O_794,N_49137,N_40813);
and UO_795 (O_795,N_49406,N_49441);
nand UO_796 (O_796,N_44109,N_42863);
and UO_797 (O_797,N_44057,N_47805);
xor UO_798 (O_798,N_46399,N_49112);
and UO_799 (O_799,N_47724,N_47151);
or UO_800 (O_800,N_45343,N_44823);
and UO_801 (O_801,N_48692,N_49561);
nand UO_802 (O_802,N_45586,N_41972);
nand UO_803 (O_803,N_42042,N_42022);
and UO_804 (O_804,N_41249,N_41124);
and UO_805 (O_805,N_45855,N_46501);
xnor UO_806 (O_806,N_49809,N_41482);
and UO_807 (O_807,N_45748,N_43247);
and UO_808 (O_808,N_42560,N_44677);
nor UO_809 (O_809,N_48664,N_45356);
nor UO_810 (O_810,N_43600,N_48101);
nor UO_811 (O_811,N_48562,N_43783);
nor UO_812 (O_812,N_47896,N_42765);
nor UO_813 (O_813,N_42095,N_48852);
nand UO_814 (O_814,N_47883,N_42947);
nand UO_815 (O_815,N_44638,N_40836);
xor UO_816 (O_816,N_48154,N_45522);
nand UO_817 (O_817,N_46688,N_45166);
nor UO_818 (O_818,N_44957,N_42445);
nor UO_819 (O_819,N_49724,N_48062);
nand UO_820 (O_820,N_46621,N_48704);
nor UO_821 (O_821,N_45582,N_48839);
nand UO_822 (O_822,N_47878,N_45595);
xnor UO_823 (O_823,N_46744,N_46507);
or UO_824 (O_824,N_46500,N_43661);
xor UO_825 (O_825,N_49627,N_44067);
and UO_826 (O_826,N_40308,N_47344);
nand UO_827 (O_827,N_49637,N_44967);
or UO_828 (O_828,N_47221,N_41481);
or UO_829 (O_829,N_49225,N_45328);
nand UO_830 (O_830,N_43908,N_47075);
nor UO_831 (O_831,N_43668,N_44416);
nand UO_832 (O_832,N_49424,N_45534);
nand UO_833 (O_833,N_49121,N_49046);
or UO_834 (O_834,N_41402,N_43203);
and UO_835 (O_835,N_47941,N_40709);
xor UO_836 (O_836,N_44504,N_43952);
nor UO_837 (O_837,N_40409,N_45318);
nand UO_838 (O_838,N_42868,N_47236);
or UO_839 (O_839,N_44166,N_42073);
or UO_840 (O_840,N_43824,N_43007);
nor UO_841 (O_841,N_45843,N_45457);
xor UO_842 (O_842,N_40984,N_46510);
and UO_843 (O_843,N_42446,N_44859);
or UO_844 (O_844,N_43225,N_41744);
xor UO_845 (O_845,N_43587,N_41798);
or UO_846 (O_846,N_40731,N_45372);
nor UO_847 (O_847,N_46263,N_41593);
nor UO_848 (O_848,N_41562,N_45157);
nand UO_849 (O_849,N_49466,N_43782);
and UO_850 (O_850,N_49596,N_41189);
or UO_851 (O_851,N_42601,N_43778);
xor UO_852 (O_852,N_46954,N_45976);
or UO_853 (O_853,N_45981,N_48058);
nor UO_854 (O_854,N_42103,N_44358);
nor UO_855 (O_855,N_47757,N_43353);
or UO_856 (O_856,N_41147,N_47314);
xnor UO_857 (O_857,N_47029,N_43766);
xor UO_858 (O_858,N_40986,N_40717);
or UO_859 (O_859,N_43664,N_46465);
or UO_860 (O_860,N_42694,N_45247);
nand UO_861 (O_861,N_48369,N_47147);
and UO_862 (O_862,N_40497,N_41140);
nor UO_863 (O_863,N_45218,N_47581);
nor UO_864 (O_864,N_40067,N_47990);
xor UO_865 (O_865,N_48437,N_45713);
or UO_866 (O_866,N_41056,N_43879);
xnor UO_867 (O_867,N_45978,N_41371);
and UO_868 (O_868,N_42899,N_46681);
nor UO_869 (O_869,N_41890,N_40357);
xnor UO_870 (O_870,N_47792,N_40345);
nand UO_871 (O_871,N_48814,N_47045);
nand UO_872 (O_872,N_43918,N_43956);
nand UO_873 (O_873,N_43014,N_49288);
nor UO_874 (O_874,N_43838,N_49573);
xnor UO_875 (O_875,N_44797,N_41058);
nand UO_876 (O_876,N_46986,N_49755);
nand UO_877 (O_877,N_47213,N_43847);
and UO_878 (O_878,N_40821,N_47873);
or UO_879 (O_879,N_46861,N_48401);
or UO_880 (O_880,N_49304,N_48463);
nand UO_881 (O_881,N_43738,N_41215);
nand UO_882 (O_882,N_45665,N_40916);
nor UO_883 (O_883,N_49215,N_41297);
and UO_884 (O_884,N_45625,N_48894);
and UO_885 (O_885,N_40078,N_44876);
nand UO_886 (O_886,N_45389,N_47132);
nor UO_887 (O_887,N_41071,N_47375);
xnor UO_888 (O_888,N_49233,N_43118);
and UO_889 (O_889,N_45374,N_44139);
or UO_890 (O_890,N_45768,N_43665);
or UO_891 (O_891,N_40327,N_46485);
nand UO_892 (O_892,N_48234,N_44160);
or UO_893 (O_893,N_47022,N_45424);
and UO_894 (O_894,N_49777,N_40421);
and UO_895 (O_895,N_45769,N_47353);
and UO_896 (O_896,N_42183,N_48434);
xnor UO_897 (O_897,N_41519,N_49980);
nor UO_898 (O_898,N_45851,N_45420);
and UO_899 (O_899,N_49041,N_43938);
nor UO_900 (O_900,N_48530,N_44678);
or UO_901 (O_901,N_47296,N_44364);
xnor UO_902 (O_902,N_49084,N_44813);
and UO_903 (O_903,N_43148,N_45535);
nor UO_904 (O_904,N_47300,N_45775);
nand UO_905 (O_905,N_44156,N_45350);
or UO_906 (O_906,N_47136,N_42663);
xor UO_907 (O_907,N_41004,N_40028);
or UO_908 (O_908,N_49259,N_45261);
nor UO_909 (O_909,N_43548,N_45232);
xor UO_910 (O_910,N_40085,N_42444);
nor UO_911 (O_911,N_48487,N_48536);
xnor UO_912 (O_912,N_42695,N_42426);
and UO_913 (O_913,N_43560,N_48343);
and UO_914 (O_914,N_45600,N_48479);
nor UO_915 (O_915,N_49863,N_40388);
and UO_916 (O_916,N_40397,N_40089);
and UO_917 (O_917,N_47586,N_44062);
and UO_918 (O_918,N_44654,N_44073);
nand UO_919 (O_919,N_48031,N_41995);
or UO_920 (O_920,N_44980,N_40014);
xnor UO_921 (O_921,N_43739,N_49593);
and UO_922 (O_922,N_44007,N_47225);
and UO_923 (O_923,N_45102,N_49727);
nand UO_924 (O_924,N_46237,N_45587);
xnor UO_925 (O_925,N_49887,N_44038);
and UO_926 (O_926,N_47882,N_47438);
nand UO_927 (O_927,N_42323,N_40425);
and UO_928 (O_928,N_42143,N_46123);
nor UO_929 (O_929,N_46559,N_45738);
xnor UO_930 (O_930,N_44905,N_43828);
nor UO_931 (O_931,N_42517,N_47065);
and UO_932 (O_932,N_45649,N_49167);
or UO_933 (O_933,N_47212,N_49375);
xor UO_934 (O_934,N_40268,N_46150);
nor UO_935 (O_935,N_41673,N_42494);
nor UO_936 (O_936,N_43005,N_43642);
xnor UO_937 (O_937,N_44255,N_45111);
and UO_938 (O_938,N_44374,N_40410);
xor UO_939 (O_939,N_41181,N_43466);
xnor UO_940 (O_940,N_44791,N_49080);
or UO_941 (O_941,N_43266,N_47736);
xor UO_942 (O_942,N_41277,N_48541);
xor UO_943 (O_943,N_46374,N_49699);
nor UO_944 (O_944,N_46475,N_41732);
or UO_945 (O_945,N_48469,N_40364);
or UO_946 (O_946,N_40293,N_49928);
or UO_947 (O_947,N_41978,N_45381);
xor UO_948 (O_948,N_46865,N_45688);
or UO_949 (O_949,N_47093,N_43091);
and UO_950 (O_950,N_42129,N_40494);
nand UO_951 (O_951,N_40911,N_40918);
nand UO_952 (O_952,N_47599,N_47399);
xnor UO_953 (O_953,N_41521,N_40619);
xnor UO_954 (O_954,N_41214,N_40554);
and UO_955 (O_955,N_43540,N_44217);
or UO_956 (O_956,N_40959,N_43803);
xor UO_957 (O_957,N_42740,N_44131);
xnor UO_958 (O_958,N_41871,N_45119);
xor UO_959 (O_959,N_43475,N_44191);
nor UO_960 (O_960,N_48396,N_43993);
or UO_961 (O_961,N_45746,N_48675);
xnor UO_962 (O_962,N_49951,N_43679);
xor UO_963 (O_963,N_48188,N_45427);
nor UO_964 (O_964,N_42131,N_44619);
nand UO_965 (O_965,N_40628,N_46063);
and UO_966 (O_966,N_41810,N_43894);
or UO_967 (O_967,N_40748,N_49452);
nor UO_968 (O_968,N_47545,N_46552);
and UO_969 (O_969,N_47905,N_48489);
nor UO_970 (O_970,N_43161,N_40480);
nor UO_971 (O_971,N_45234,N_46090);
nor UO_972 (O_972,N_49110,N_43930);
nor UO_973 (O_973,N_40000,N_49213);
or UO_974 (O_974,N_45273,N_48504);
and UO_975 (O_975,N_41554,N_41735);
or UO_976 (O_976,N_49792,N_43397);
nor UO_977 (O_977,N_41734,N_49097);
or UO_978 (O_978,N_45767,N_47262);
nor UO_979 (O_979,N_43216,N_49327);
xnor UO_980 (O_980,N_41846,N_40752);
or UO_981 (O_981,N_48442,N_47647);
nor UO_982 (O_982,N_44860,N_48665);
nand UO_983 (O_983,N_42745,N_45032);
nand UO_984 (O_984,N_44266,N_42850);
nor UO_985 (O_985,N_45935,N_40307);
nand UO_986 (O_986,N_48025,N_48214);
or UO_987 (O_987,N_40486,N_45144);
xor UO_988 (O_988,N_40670,N_40163);
and UO_989 (O_989,N_45230,N_46022);
nor UO_990 (O_990,N_49130,N_44277);
xnor UO_991 (O_991,N_42588,N_45926);
nor UO_992 (O_992,N_43578,N_42256);
nor UO_993 (O_993,N_40617,N_48661);
or UO_994 (O_994,N_43059,N_49131);
nor UO_995 (O_995,N_49107,N_43019);
xnor UO_996 (O_996,N_42020,N_41493);
nor UO_997 (O_997,N_48721,N_49655);
and UO_998 (O_998,N_42813,N_49946);
or UO_999 (O_999,N_42195,N_44946);
xor UO_1000 (O_1000,N_47019,N_46108);
nor UO_1001 (O_1001,N_43211,N_45287);
nor UO_1002 (O_1002,N_45437,N_45216);
nor UO_1003 (O_1003,N_44475,N_47855);
or UO_1004 (O_1004,N_47025,N_40111);
and UO_1005 (O_1005,N_42281,N_49226);
and UO_1006 (O_1006,N_45249,N_43309);
or UO_1007 (O_1007,N_43931,N_42574);
and UO_1008 (O_1008,N_49944,N_43935);
or UO_1009 (O_1009,N_47533,N_44206);
nand UO_1010 (O_1010,N_48070,N_49877);
nor UO_1011 (O_1011,N_44632,N_48327);
and UO_1012 (O_1012,N_47110,N_44419);
or UO_1013 (O_1013,N_41537,N_46649);
xnor UO_1014 (O_1014,N_42964,N_45224);
xnor UO_1015 (O_1015,N_45813,N_44106);
or UO_1016 (O_1016,N_46825,N_43135);
nand UO_1017 (O_1017,N_42939,N_43691);
nand UO_1018 (O_1018,N_49250,N_49377);
and UO_1019 (O_1019,N_46551,N_44170);
xor UO_1020 (O_1020,N_43198,N_42989);
xor UO_1021 (O_1021,N_48924,N_45542);
and UO_1022 (O_1022,N_48378,N_40733);
and UO_1023 (O_1023,N_41433,N_40761);
nor UO_1024 (O_1024,N_45209,N_41109);
or UO_1025 (O_1025,N_48061,N_43306);
or UO_1026 (O_1026,N_49866,N_42811);
nor UO_1027 (O_1027,N_48626,N_49910);
nand UO_1028 (O_1028,N_44248,N_49735);
nand UO_1029 (O_1029,N_46926,N_46616);
nor UO_1030 (O_1030,N_44283,N_46646);
xor UO_1031 (O_1031,N_46612,N_41076);
and UO_1032 (O_1032,N_44647,N_41358);
xor UO_1033 (O_1033,N_46526,N_46095);
nor UO_1034 (O_1034,N_48617,N_41989);
and UO_1035 (O_1035,N_45610,N_43021);
xor UO_1036 (O_1036,N_43268,N_42140);
nand UO_1037 (O_1037,N_48507,N_49907);
nand UO_1038 (O_1038,N_45187,N_43304);
xnor UO_1039 (O_1039,N_42520,N_45693);
or UO_1040 (O_1040,N_48816,N_46793);
or UO_1041 (O_1041,N_47522,N_47156);
nand UO_1042 (O_1042,N_43728,N_41865);
nand UO_1043 (O_1043,N_45334,N_46913);
xnor UO_1044 (O_1044,N_43703,N_47216);
or UO_1045 (O_1045,N_41387,N_45774);
nand UO_1046 (O_1046,N_49371,N_45601);
and UO_1047 (O_1047,N_46083,N_44612);
nor UO_1048 (O_1048,N_44663,N_43635);
nand UO_1049 (O_1049,N_49337,N_41271);
xnor UO_1050 (O_1050,N_46951,N_48160);
and UO_1051 (O_1051,N_49419,N_45276);
and UO_1052 (O_1052,N_40504,N_42783);
or UO_1053 (O_1053,N_46833,N_45436);
or UO_1054 (O_1054,N_46959,N_42618);
xnor UO_1055 (O_1055,N_42250,N_46774);
nand UO_1056 (O_1056,N_49533,N_43286);
or UO_1057 (O_1057,N_42608,N_43345);
or UO_1058 (O_1058,N_40841,N_47017);
or UO_1059 (O_1059,N_40759,N_47155);
and UO_1060 (O_1060,N_49632,N_42251);
and UO_1061 (O_1061,N_42123,N_41499);
nand UO_1062 (O_1062,N_41820,N_40105);
nor UO_1063 (O_1063,N_43823,N_40012);
xnor UO_1064 (O_1064,N_41747,N_42405);
nor UO_1065 (O_1065,N_45308,N_40173);
nand UO_1066 (O_1066,N_45853,N_45583);
xnor UO_1067 (O_1067,N_43374,N_41782);
nand UO_1068 (O_1068,N_45724,N_41384);
nand UO_1069 (O_1069,N_49209,N_41365);
or UO_1070 (O_1070,N_41034,N_40071);
and UO_1071 (O_1071,N_43010,N_43547);
nor UO_1072 (O_1072,N_48912,N_44904);
or UO_1073 (O_1073,N_43233,N_40207);
nand UO_1074 (O_1074,N_41950,N_48811);
nor UO_1075 (O_1075,N_47919,N_47317);
nor UO_1076 (O_1076,N_40957,N_47051);
nor UO_1077 (O_1077,N_49689,N_40674);
nand UO_1078 (O_1078,N_43511,N_49971);
or UO_1079 (O_1079,N_48008,N_43715);
or UO_1080 (O_1080,N_42531,N_41739);
or UO_1081 (O_1081,N_41066,N_48212);
or UO_1082 (O_1082,N_49086,N_49797);
and UO_1083 (O_1083,N_41235,N_48081);
and UO_1084 (O_1084,N_40672,N_42887);
and UO_1085 (O_1085,N_49892,N_41420);
and UO_1086 (O_1086,N_41419,N_44915);
or UO_1087 (O_1087,N_46369,N_44850);
and UO_1088 (O_1088,N_41480,N_49488);
nor UO_1089 (O_1089,N_42814,N_41578);
nand UO_1090 (O_1090,N_44936,N_44968);
nor UO_1091 (O_1091,N_41183,N_46011);
or UO_1092 (O_1092,N_43454,N_44989);
nand UO_1093 (O_1093,N_43463,N_42217);
and UO_1094 (O_1094,N_44484,N_47238);
or UO_1095 (O_1095,N_42100,N_40557);
and UO_1096 (O_1096,N_43794,N_44665);
and UO_1097 (O_1097,N_46434,N_47231);
xnor UO_1098 (O_1098,N_49396,N_43051);
nand UO_1099 (O_1099,N_41199,N_47441);
xnor UO_1100 (O_1100,N_48834,N_42295);
xor UO_1101 (O_1101,N_46484,N_43810);
and UO_1102 (O_1102,N_49831,N_49240);
nand UO_1103 (O_1103,N_47711,N_48278);
nand UO_1104 (O_1104,N_40384,N_49313);
nand UO_1105 (O_1105,N_46291,N_47095);
or UO_1106 (O_1106,N_46189,N_48920);
xnor UO_1107 (O_1107,N_46367,N_49972);
xor UO_1108 (O_1108,N_41676,N_41609);
xor UO_1109 (O_1109,N_49067,N_49636);
xor UO_1110 (O_1110,N_49142,N_45365);
or UO_1111 (O_1111,N_46194,N_42858);
nand UO_1112 (O_1112,N_40406,N_48714);
xor UO_1113 (O_1113,N_42860,N_43853);
nand UO_1114 (O_1114,N_43246,N_40726);
nand UO_1115 (O_1115,N_47390,N_49354);
or UO_1116 (O_1116,N_47083,N_45599);
xor UO_1117 (O_1117,N_46032,N_46678);
nand UO_1118 (O_1118,N_48052,N_48533);
or UO_1119 (O_1119,N_41657,N_47734);
xnor UO_1120 (O_1120,N_44914,N_40632);
nor UO_1121 (O_1121,N_45613,N_44114);
xor UO_1122 (O_1122,N_48082,N_40800);
nand UO_1123 (O_1123,N_48111,N_40849);
xor UO_1124 (O_1124,N_43768,N_45811);
and UO_1125 (O_1125,N_45513,N_42077);
or UO_1126 (O_1126,N_44424,N_45377);
xnor UO_1127 (O_1127,N_46152,N_44095);
and UO_1128 (O_1128,N_45405,N_42296);
or UO_1129 (O_1129,N_48971,N_41364);
nor UO_1130 (O_1130,N_49140,N_43954);
nor UO_1131 (O_1131,N_43899,N_43284);
nor UO_1132 (O_1132,N_43146,N_46470);
nor UO_1133 (O_1133,N_41338,N_46354);
or UO_1134 (O_1134,N_45580,N_42155);
nand UO_1135 (O_1135,N_45191,N_48938);
nand UO_1136 (O_1136,N_41324,N_42967);
nand UO_1137 (O_1137,N_44863,N_42888);
and UO_1138 (O_1138,N_47731,N_49600);
or UO_1139 (O_1139,N_48552,N_46815);
or UO_1140 (O_1140,N_45134,N_48830);
xor UO_1141 (O_1141,N_48059,N_43817);
and UO_1142 (O_1142,N_48800,N_42127);
nand UO_1143 (O_1143,N_46908,N_47021);
nand UO_1144 (O_1144,N_47487,N_49581);
nor UO_1145 (O_1145,N_47070,N_41789);
nand UO_1146 (O_1146,N_46561,N_45120);
nor UO_1147 (O_1147,N_42926,N_48410);
xnor UO_1148 (O_1148,N_47654,N_49197);
nor UO_1149 (O_1149,N_49332,N_44662);
xor UO_1150 (O_1150,N_48300,N_45278);
xor UO_1151 (O_1151,N_48866,N_42797);
nand UO_1152 (O_1152,N_49314,N_47505);
or UO_1153 (O_1153,N_41594,N_48757);
or UO_1154 (O_1154,N_42089,N_42902);
nor UO_1155 (O_1155,N_40531,N_48829);
nand UO_1156 (O_1156,N_48399,N_47237);
nor UO_1157 (O_1157,N_48237,N_41307);
or UO_1158 (O_1158,N_44000,N_40675);
nand UO_1159 (O_1159,N_45524,N_46733);
nand UO_1160 (O_1160,N_45340,N_42441);
nor UO_1161 (O_1161,N_47590,N_42590);
nand UO_1162 (O_1162,N_43109,N_48535);
or UO_1163 (O_1163,N_43583,N_45526);
or UO_1164 (O_1164,N_49404,N_47009);
nor UO_1165 (O_1165,N_42718,N_49021);
nand UO_1166 (O_1166,N_46270,N_46293);
or UO_1167 (O_1167,N_47145,N_46215);
nor UO_1168 (O_1168,N_48202,N_46303);
or UO_1169 (O_1169,N_46538,N_43789);
or UO_1170 (O_1170,N_48616,N_46168);
nor UO_1171 (O_1171,N_45537,N_40735);
xor UO_1172 (O_1172,N_45966,N_47538);
and UO_1173 (O_1173,N_48837,N_41368);
xor UO_1174 (O_1174,N_49064,N_47365);
or UO_1175 (O_1175,N_41200,N_41841);
or UO_1176 (O_1176,N_43307,N_46517);
and UO_1177 (O_1177,N_47055,N_43162);
or UO_1178 (O_1178,N_45969,N_40127);
nor UO_1179 (O_1179,N_42942,N_46494);
and UO_1180 (O_1180,N_47570,N_47637);
xor UO_1181 (O_1181,N_42855,N_47358);
nand UO_1182 (O_1182,N_46993,N_49579);
nor UO_1183 (O_1183,N_41895,N_40372);
and UO_1184 (O_1184,N_45576,N_42793);
and UO_1185 (O_1185,N_44711,N_44372);
and UO_1186 (O_1186,N_41644,N_41536);
or UO_1187 (O_1187,N_41316,N_42529);
xnor UO_1188 (O_1188,N_48908,N_47803);
xnor UO_1189 (O_1189,N_40689,N_45743);
nor UO_1190 (O_1190,N_47890,N_40586);
xor UO_1191 (O_1191,N_48841,N_45819);
and UO_1192 (O_1192,N_44892,N_41306);
and UO_1193 (O_1193,N_49260,N_48143);
nor UO_1194 (O_1194,N_46002,N_40002);
xnor UO_1195 (O_1195,N_49074,N_43943);
xor UO_1196 (O_1196,N_42971,N_42442);
or UO_1197 (O_1197,N_47793,N_45488);
or UO_1198 (O_1198,N_41981,N_42500);
nand UO_1199 (O_1199,N_41500,N_45484);
nor UO_1200 (O_1200,N_44994,N_44852);
xor UO_1201 (O_1201,N_40277,N_42686);
nand UO_1202 (O_1202,N_40143,N_43354);
xor UO_1203 (O_1203,N_45319,N_49913);
or UO_1204 (O_1204,N_47588,N_42732);
nor UO_1205 (O_1205,N_45933,N_42803);
nor UO_1206 (O_1206,N_49544,N_42853);
xor UO_1207 (O_1207,N_42478,N_45042);
xnor UO_1208 (O_1208,N_41012,N_44006);
nand UO_1209 (O_1209,N_48745,N_43381);
nand UO_1210 (O_1210,N_49181,N_40058);
or UO_1211 (O_1211,N_49717,N_47354);
nor UO_1212 (O_1212,N_43031,N_40972);
nor UO_1213 (O_1213,N_44624,N_42840);
or UO_1214 (O_1214,N_41060,N_40233);
and UO_1215 (O_1215,N_45979,N_41639);
nor UO_1216 (O_1216,N_41261,N_46400);
nor UO_1217 (O_1217,N_47769,N_48257);
nand UO_1218 (O_1218,N_49695,N_43147);
and UO_1219 (O_1219,N_42257,N_47279);
xor UO_1220 (O_1220,N_45512,N_41743);
and UO_1221 (O_1221,N_40652,N_41112);
and UO_1222 (O_1222,N_41013,N_46610);
and UO_1223 (O_1223,N_45764,N_46532);
nor UO_1224 (O_1224,N_40591,N_40536);
and UO_1225 (O_1225,N_47986,N_43517);
nand UO_1226 (O_1226,N_47685,N_46242);
xor UO_1227 (O_1227,N_42111,N_48289);
xnor UO_1228 (O_1228,N_45444,N_41245);
xnor UO_1229 (O_1229,N_43228,N_46625);
xnor UO_1230 (O_1230,N_44054,N_47626);
or UO_1231 (O_1231,N_40037,N_41649);
and UO_1232 (O_1232,N_46770,N_49350);
or UO_1233 (O_1233,N_47964,N_47662);
nor UO_1234 (O_1234,N_46653,N_42451);
xnor UO_1235 (O_1235,N_48717,N_43871);
xor UO_1236 (O_1236,N_46077,N_47211);
or UO_1237 (O_1237,N_48253,N_40232);
nor UO_1238 (O_1238,N_49082,N_44567);
nand UO_1239 (O_1239,N_48798,N_40398);
or UO_1240 (O_1240,N_46872,N_49492);
nand UO_1241 (O_1241,N_48385,N_49201);
nor UO_1242 (O_1242,N_48989,N_41312);
nor UO_1243 (O_1243,N_40462,N_49642);
nor UO_1244 (O_1244,N_41287,N_42359);
and UO_1245 (O_1245,N_41719,N_47909);
nand UO_1246 (O_1246,N_44759,N_47503);
or UO_1247 (O_1247,N_41612,N_40465);
nor UO_1248 (O_1248,N_42991,N_47126);
nand UO_1249 (O_1249,N_45480,N_42175);
xor UO_1250 (O_1250,N_47811,N_40931);
and UO_1251 (O_1251,N_45623,N_46641);
nand UO_1252 (O_1252,N_48205,N_48055);
and UO_1253 (O_1253,N_44154,N_46522);
and UO_1254 (O_1254,N_41278,N_43166);
nor UO_1255 (O_1255,N_43634,N_43663);
xnor UO_1256 (O_1256,N_45251,N_46635);
nor UO_1257 (O_1257,N_41115,N_47111);
or UO_1258 (O_1258,N_45360,N_42714);
nor UO_1259 (O_1259,N_41212,N_46787);
or UO_1260 (O_1260,N_40361,N_42086);
nand UO_1261 (O_1261,N_46587,N_46259);
and UO_1262 (O_1262,N_40720,N_46145);
nand UO_1263 (O_1263,N_45912,N_44592);
nand UO_1264 (O_1264,N_44289,N_46937);
or UO_1265 (O_1265,N_43892,N_45037);
nor UO_1266 (O_1266,N_43973,N_48239);
nand UO_1267 (O_1267,N_42929,N_45238);
or UO_1268 (O_1268,N_48657,N_45296);
nor UO_1269 (O_1269,N_48072,N_49549);
or UO_1270 (O_1270,N_48474,N_41795);
or UO_1271 (O_1271,N_43175,N_48280);
or UO_1272 (O_1272,N_44845,N_49628);
nor UO_1273 (O_1273,N_48032,N_40335);
nand UO_1274 (O_1274,N_49254,N_42193);
and UO_1275 (O_1275,N_41624,N_49501);
nor UO_1276 (O_1276,N_49394,N_44670);
and UO_1277 (O_1277,N_40656,N_43316);
or UO_1278 (O_1278,N_49292,N_49231);
nand UO_1279 (O_1279,N_48044,N_44079);
nand UO_1280 (O_1280,N_46319,N_40261);
or UO_1281 (O_1281,N_41717,N_41141);
nor UO_1282 (O_1282,N_46445,N_44652);
nand UO_1283 (O_1283,N_47707,N_41709);
nor UO_1284 (O_1284,N_42316,N_44193);
xor UO_1285 (O_1285,N_46960,N_47663);
xor UO_1286 (O_1286,N_47817,N_40703);
and UO_1287 (O_1287,N_48383,N_40574);
xnor UO_1288 (O_1288,N_44182,N_42471);
nor UO_1289 (O_1289,N_47530,N_41447);
nand UO_1290 (O_1290,N_44298,N_48461);
nor UO_1291 (O_1291,N_42337,N_45474);
nor UO_1292 (O_1292,N_47785,N_45833);
nand UO_1293 (O_1293,N_46037,N_46323);
nor UO_1294 (O_1294,N_40489,N_40495);
or UO_1295 (O_1295,N_41096,N_47349);
and UO_1296 (O_1296,N_44187,N_48696);
nor UO_1297 (O_1297,N_40883,N_48825);
xnor UO_1298 (O_1298,N_42331,N_46171);
nand UO_1299 (O_1299,N_48620,N_41457);
nand UO_1300 (O_1300,N_46064,N_45893);
xor UO_1301 (O_1301,N_47456,N_41730);
nor UO_1302 (O_1302,N_45557,N_44392);
nand UO_1303 (O_1303,N_47806,N_40724);
and UO_1304 (O_1304,N_41460,N_46820);
nand UO_1305 (O_1305,N_47429,N_44029);
nand UO_1306 (O_1306,N_41430,N_42484);
nand UO_1307 (O_1307,N_46264,N_44801);
or UO_1308 (O_1308,N_45507,N_40610);
nand UO_1309 (O_1309,N_44599,N_42787);
or UO_1310 (O_1310,N_48359,N_47865);
nand UO_1311 (O_1311,N_45189,N_49619);
xnor UO_1312 (O_1312,N_45828,N_41763);
nor UO_1313 (O_1313,N_41081,N_40329);
nand UO_1314 (O_1314,N_42889,N_48268);
nor UO_1315 (O_1315,N_40607,N_42391);
nand UO_1316 (O_1316,N_47704,N_49245);
and UO_1317 (O_1317,N_47143,N_44210);
nor UO_1318 (O_1318,N_46528,N_45416);
and UO_1319 (O_1319,N_46067,N_47746);
xnor UO_1320 (O_1320,N_41804,N_45031);
xor UO_1321 (O_1321,N_42511,N_41894);
and UO_1322 (O_1322,N_40832,N_40551);
or UO_1323 (O_1323,N_41535,N_44442);
and UO_1324 (O_1324,N_48349,N_48140);
or UO_1325 (O_1325,N_44040,N_41426);
or UO_1326 (O_1326,N_42988,N_49851);
or UO_1327 (O_1327,N_47779,N_43011);
nand UO_1328 (O_1328,N_48262,N_42350);
or UO_1329 (O_1329,N_43524,N_46692);
or UO_1330 (O_1330,N_41120,N_47867);
nor UO_1331 (O_1331,N_42474,N_49318);
nor UO_1332 (O_1332,N_48860,N_44587);
nand UO_1333 (O_1333,N_41019,N_43404);
nand UO_1334 (O_1334,N_43746,N_45359);
nand UO_1335 (O_1335,N_43543,N_40790);
nor UO_1336 (O_1336,N_44335,N_45793);
and UO_1337 (O_1337,N_42629,N_42229);
nand UO_1338 (O_1338,N_44898,N_44660);
and UO_1339 (O_1339,N_46004,N_45906);
nand UO_1340 (O_1340,N_49968,N_48316);
and UO_1341 (O_1341,N_46807,N_42334);
nor UO_1342 (O_1342,N_44072,N_40952);
or UO_1343 (O_1343,N_47564,N_47723);
or UO_1344 (O_1344,N_43756,N_44754);
nand UO_1345 (O_1345,N_49346,N_42872);
and UO_1346 (O_1346,N_47367,N_47935);
or UO_1347 (O_1347,N_48564,N_48857);
xnor UO_1348 (O_1348,N_44849,N_45293);
nor UO_1349 (O_1349,N_49361,N_44986);
nand UO_1350 (O_1350,N_46098,N_48220);
and UO_1351 (O_1351,N_48753,N_49385);
xor UO_1352 (O_1352,N_40511,N_40713);
xnor UO_1353 (O_1353,N_42739,N_41957);
nor UO_1354 (O_1354,N_45934,N_42404);
or UO_1355 (O_1355,N_46601,N_48911);
and UO_1356 (O_1356,N_43453,N_48037);
and UO_1357 (O_1357,N_43442,N_49960);
and UO_1358 (O_1358,N_49932,N_44769);
or UO_1359 (O_1359,N_44455,N_43500);
nand UO_1360 (O_1360,N_46102,N_43720);
and UO_1361 (O_1361,N_41541,N_43751);
nand UO_1362 (O_1362,N_49793,N_49212);
and UO_1363 (O_1363,N_42276,N_44041);
nor UO_1364 (O_1364,N_41670,N_48199);
nand UO_1365 (O_1365,N_45548,N_43054);
and UO_1366 (O_1366,N_44396,N_46163);
and UO_1367 (O_1367,N_41159,N_45699);
and UO_1368 (O_1368,N_46335,N_45107);
nor UO_1369 (O_1369,N_44393,N_46105);
xor UO_1370 (O_1370,N_42014,N_43868);
nand UO_1371 (O_1371,N_42298,N_48928);
nand UO_1372 (O_1372,N_41712,N_48638);
xor UO_1373 (O_1373,N_47940,N_49380);
or UO_1374 (O_1374,N_40243,N_47598);
xor UO_1375 (O_1375,N_40190,N_41557);
or UO_1376 (O_1376,N_48871,N_43050);
xnor UO_1377 (O_1377,N_47870,N_49620);
nand UO_1378 (O_1378,N_40223,N_48007);
xnor UO_1379 (O_1379,N_43633,N_48526);
nor UO_1380 (O_1380,N_45027,N_46589);
or UO_1381 (O_1381,N_49697,N_43426);
nand UO_1382 (O_1382,N_44414,N_43808);
nor UO_1383 (O_1383,N_41326,N_40996);
or UO_1384 (O_1384,N_42258,N_40993);
nand UO_1385 (O_1385,N_40400,N_47742);
nand UO_1386 (O_1386,N_42912,N_48235);
xor UO_1387 (O_1387,N_44645,N_40290);
nand UO_1388 (O_1388,N_45063,N_48732);
nor UO_1389 (O_1389,N_48445,N_41229);
or UO_1390 (O_1390,N_43666,N_44087);
nor UO_1391 (O_1391,N_49606,N_43460);
or UO_1392 (O_1392,N_42877,N_42841);
xor UO_1393 (O_1393,N_43880,N_45581);
and UO_1394 (O_1394,N_47850,N_40744);
nor UO_1395 (O_1395,N_42382,N_42976);
nand UO_1396 (O_1396,N_46759,N_44987);
nand UO_1397 (O_1397,N_46980,N_44861);
xnor UO_1398 (O_1398,N_46371,N_42463);
or UO_1399 (O_1399,N_46198,N_44432);
or UO_1400 (O_1400,N_48522,N_48411);
xnor UO_1401 (O_1401,N_42580,N_40702);
xnor UO_1402 (O_1402,N_40294,N_43610);
xor UO_1403 (O_1403,N_43349,N_47892);
or UO_1404 (O_1404,N_49559,N_41167);
nor UO_1405 (O_1405,N_41163,N_44185);
and UO_1406 (O_1406,N_40553,N_41062);
nor UO_1407 (O_1407,N_45923,N_45097);
or UO_1408 (O_1408,N_40314,N_41072);
xor UO_1409 (O_1409,N_45608,N_42553);
xor UO_1410 (O_1410,N_49912,N_45802);
nor UO_1411 (O_1411,N_44857,N_46343);
and UO_1412 (O_1412,N_46169,N_49368);
or UO_1413 (O_1413,N_46144,N_41702);
nor UO_1414 (O_1414,N_41874,N_42459);
or UO_1415 (O_1415,N_46605,N_40736);
xor UO_1416 (O_1416,N_41549,N_44398);
or UO_1417 (O_1417,N_48409,N_49329);
xor UO_1418 (O_1418,N_44541,N_43522);
xor UO_1419 (O_1419,N_48904,N_47502);
nand UO_1420 (O_1420,N_40281,N_45527);
or UO_1421 (O_1421,N_45303,N_49890);
nor UO_1422 (O_1422,N_46388,N_41765);
or UO_1423 (O_1423,N_47232,N_49816);
or UO_1424 (O_1424,N_45445,N_40900);
and UO_1425 (O_1425,N_45014,N_42373);
or UO_1426 (O_1426,N_49188,N_41534);
nor UO_1427 (O_1427,N_40605,N_42418);
and UO_1428 (O_1428,N_40882,N_44044);
xor UO_1429 (O_1429,N_44259,N_43497);
xor UO_1430 (O_1430,N_47614,N_48168);
or UO_1431 (O_1431,N_45787,N_45875);
or UO_1432 (O_1432,N_44751,N_44750);
nor UO_1433 (O_1433,N_40500,N_41814);
and UO_1434 (O_1434,N_46499,N_41061);
xor UO_1435 (O_1435,N_41886,N_45849);
nand UO_1436 (O_1436,N_43248,N_47753);
nand UO_1437 (O_1437,N_42880,N_47615);
xor UO_1438 (O_1438,N_49999,N_49843);
and UO_1439 (O_1439,N_47222,N_48861);
and UO_1440 (O_1440,N_45167,N_45654);
nor UO_1441 (O_1441,N_43099,N_46862);
nor UO_1442 (O_1442,N_44136,N_48248);
or UO_1443 (O_1443,N_40490,N_48654);
and UO_1444 (O_1444,N_41262,N_40529);
xor UO_1445 (O_1445,N_43364,N_45220);
or UO_1446 (O_1446,N_44774,N_44589);
nor UO_1447 (O_1447,N_42322,N_40562);
nand UO_1448 (O_1448,N_40824,N_43564);
and UO_1449 (O_1449,N_43458,N_46847);
xor UO_1450 (O_1450,N_47403,N_44572);
nand UO_1451 (O_1451,N_45265,N_45316);
nand UO_1452 (O_1452,N_40330,N_45754);
xnor UO_1453 (O_1453,N_43707,N_45277);
xor UO_1454 (O_1454,N_45593,N_43512);
nor UO_1455 (O_1455,N_43209,N_47355);
nand UO_1456 (O_1456,N_41343,N_45417);
and UO_1457 (O_1457,N_45332,N_47559);
nand UO_1458 (O_1458,N_49985,N_42605);
and UO_1459 (O_1459,N_45940,N_44657);
nand UO_1460 (O_1460,N_46296,N_44719);
nand UO_1461 (O_1461,N_43335,N_44910);
xnor UO_1462 (O_1462,N_40902,N_43549);
nor UO_1463 (O_1463,N_42756,N_44562);
nor UO_1464 (O_1464,N_45093,N_40978);
and UO_1465 (O_1465,N_46727,N_41545);
and UO_1466 (O_1466,N_44207,N_40810);
and UO_1467 (O_1467,N_49740,N_48339);
xor UO_1468 (O_1468,N_45468,N_45223);
xor UO_1469 (O_1469,N_47756,N_45025);
or UO_1470 (O_1470,N_45643,N_41374);
xor UO_1471 (O_1471,N_41221,N_41958);
and UO_1472 (O_1472,N_49173,N_43646);
nor UO_1473 (O_1473,N_42915,N_45379);
nor UO_1474 (O_1474,N_42870,N_40693);
or UO_1475 (O_1475,N_44961,N_48951);
nand UO_1476 (O_1476,N_41831,N_44524);
nor UO_1477 (O_1477,N_46352,N_47557);
nor UO_1478 (O_1478,N_43227,N_43628);
or UO_1479 (O_1479,N_45668,N_43594);
or UO_1480 (O_1480,N_45784,N_47783);
nor UO_1481 (O_1481,N_49578,N_47490);
and UO_1482 (O_1482,N_43301,N_40041);
and UO_1483 (O_1483,N_49132,N_40460);
nand UO_1484 (O_1484,N_48071,N_43539);
or UO_1485 (O_1485,N_48039,N_46155);
nand UO_1486 (O_1486,N_44617,N_43473);
nor UO_1487 (O_1487,N_48029,N_48990);
nand UO_1488 (O_1488,N_48102,N_47625);
and UO_1489 (O_1489,N_47804,N_45219);
and UO_1490 (O_1490,N_47461,N_43815);
nand UO_1491 (O_1491,N_40569,N_46735);
and UO_1492 (O_1492,N_42332,N_43712);
or UO_1493 (O_1493,N_43389,N_48133);
and UO_1494 (O_1494,N_43752,N_49066);
xor UO_1495 (O_1495,N_40723,N_43392);
nand UO_1496 (O_1496,N_41850,N_45375);
nand UO_1497 (O_1497,N_43573,N_42613);
and UO_1498 (O_1498,N_45637,N_48098);
or UO_1499 (O_1499,N_41074,N_41561);
or UO_1500 (O_1500,N_48953,N_49883);
nand UO_1501 (O_1501,N_48726,N_46698);
xor UO_1502 (O_1502,N_42412,N_47068);
nor UO_1503 (O_1503,N_45245,N_47271);
xnor UO_1504 (O_1504,N_48004,N_43274);
xor UO_1505 (O_1505,N_40572,N_40038);
nor UO_1506 (O_1506,N_45854,N_46280);
and UO_1507 (O_1507,N_41769,N_41396);
nor UO_1508 (O_1508,N_42491,N_42866);
or UO_1509 (O_1509,N_41190,N_44149);
and UO_1510 (O_1510,N_46683,N_43264);
xor UO_1511 (O_1511,N_48166,N_42844);
nor UO_1512 (O_1512,N_42800,N_46084);
or UO_1513 (O_1513,N_47534,N_44881);
and UO_1514 (O_1514,N_46351,N_40237);
xnor UO_1515 (O_1515,N_41164,N_40408);
nor UO_1516 (O_1516,N_47131,N_40860);
nand UO_1517 (O_1517,N_48402,N_41067);
and UO_1518 (O_1518,N_47834,N_46824);
nor UO_1519 (O_1519,N_45289,N_46984);
and UO_1520 (O_1520,N_44035,N_44584);
nand UO_1521 (O_1521,N_46009,N_46715);
and UO_1522 (O_1522,N_43724,N_48013);
or UO_1523 (O_1523,N_48876,N_44215);
or UO_1524 (O_1524,N_49448,N_41378);
or UO_1525 (O_1525,N_45776,N_49798);
and UO_1526 (O_1526,N_47795,N_47957);
and UO_1527 (O_1527,N_49666,N_42522);
and UO_1528 (O_1528,N_49853,N_47328);
nand UO_1529 (O_1529,N_42910,N_45307);
nor UO_1530 (O_1530,N_49299,N_45761);
xnor UO_1531 (O_1531,N_49343,N_46148);
or UO_1532 (O_1532,N_46069,N_48932);
and UO_1533 (O_1533,N_41807,N_46617);
nand UO_1534 (O_1534,N_49813,N_40929);
xnor UO_1535 (O_1535,N_46705,N_41891);
xnor UO_1536 (O_1536,N_42893,N_44580);
and UO_1537 (O_1537,N_41427,N_46795);
and UO_1538 (O_1538,N_49880,N_49075);
xnor UO_1539 (O_1539,N_42433,N_45647);
nand UO_1540 (O_1540,N_44826,N_48954);
or UO_1541 (O_1541,N_41903,N_43325);
and UO_1542 (O_1542,N_48770,N_43811);
xnor UO_1543 (O_1543,N_47766,N_40288);
or UO_1544 (O_1544,N_40522,N_48710);
or UO_1545 (O_1545,N_43872,N_42240);
and UO_1546 (O_1546,N_49817,N_45105);
xnor UO_1547 (O_1547,N_43155,N_41631);
nand UO_1548 (O_1548,N_46001,N_48666);
xnor UO_1549 (O_1549,N_43485,N_46869);
xnor UO_1550 (O_1550,N_45423,N_41359);
nor UO_1551 (O_1551,N_46920,N_45555);
and UO_1552 (O_1552,N_47106,N_41969);
xor UO_1553 (O_1553,N_49974,N_40561);
nand UO_1554 (O_1554,N_43632,N_48893);
nor UO_1555 (O_1555,N_47449,N_40818);
and UO_1556 (O_1556,N_40767,N_41918);
nand UO_1557 (O_1557,N_44515,N_41240);
nor UO_1558 (O_1558,N_45735,N_48937);
xor UO_1559 (O_1559,N_45605,N_46624);
or UO_1560 (O_1560,N_48780,N_48225);
nor UO_1561 (O_1561,N_42974,N_46257);
or UO_1562 (O_1562,N_42981,N_48925);
nor UO_1563 (O_1563,N_47733,N_42936);
or UO_1564 (O_1564,N_49506,N_40634);
and UO_1565 (O_1565,N_49694,N_49565);
or UO_1566 (O_1566,N_44830,N_42340);
nand UO_1567 (O_1567,N_45780,N_46397);
nand UO_1568 (O_1568,N_45322,N_48363);
and UO_1569 (O_1569,N_47857,N_45556);
nor UO_1570 (O_1570,N_48607,N_49782);
or UO_1571 (O_1571,N_48615,N_49750);
or UO_1572 (O_1572,N_48529,N_45505);
nand UO_1573 (O_1573,N_45885,N_40266);
and UO_1574 (O_1574,N_41628,N_48843);
xnor UO_1575 (O_1575,N_45609,N_45150);
nand UO_1576 (O_1576,N_47998,N_45823);
xnor UO_1577 (O_1577,N_40844,N_42408);
nand UO_1578 (O_1578,N_41488,N_45991);
xor UO_1579 (O_1579,N_41591,N_45392);
nand UO_1580 (O_1580,N_49672,N_40622);
xnor UO_1581 (O_1581,N_49358,N_45075);
xor UO_1582 (O_1582,N_41247,N_40579);
or UO_1583 (O_1583,N_44032,N_45763);
nand UO_1584 (O_1584,N_49860,N_46516);
nor UO_1585 (O_1585,N_43686,N_43947);
or UO_1586 (O_1586,N_45051,N_48739);
nor UO_1587 (O_1587,N_41671,N_41828);
or UO_1588 (O_1588,N_41802,N_46040);
or UO_1589 (O_1589,N_40934,N_42034);
and UO_1590 (O_1590,N_48688,N_48551);
and UO_1591 (O_1591,N_44679,N_40348);
nor UO_1592 (O_1592,N_43201,N_44200);
or UO_1593 (O_1593,N_43486,N_44394);
and UO_1594 (O_1594,N_44509,N_43323);
and UO_1595 (O_1595,N_42205,N_41321);
nand UO_1596 (O_1596,N_42816,N_42818);
or UO_1597 (O_1597,N_47515,N_45499);
or UO_1598 (O_1598,N_48249,N_44102);
nor UO_1599 (O_1599,N_42390,N_48754);
xor UO_1600 (O_1600,N_44588,N_49769);
nand UO_1601 (O_1601,N_43375,N_41812);
or UO_1602 (O_1602,N_45831,N_46075);
or UO_1603 (O_1603,N_44585,N_40129);
or UO_1604 (O_1604,N_45428,N_40003);
xnor UO_1605 (O_1605,N_40754,N_46013);
nor UO_1606 (O_1606,N_49736,N_47639);
and UO_1607 (O_1607,N_44075,N_47341);
nand UO_1608 (O_1608,N_42497,N_41510);
and UO_1609 (O_1609,N_43527,N_41370);
and UO_1610 (O_1610,N_49538,N_48430);
and UO_1611 (O_1611,N_45205,N_45836);
nor UO_1612 (O_1612,N_42710,N_48126);
nor UO_1613 (O_1613,N_40879,N_49205);
nor UO_1614 (O_1614,N_40788,N_45905);
or UO_1615 (O_1615,N_40234,N_44128);
or UO_1616 (O_1616,N_47104,N_40415);
nand UO_1617 (O_1617,N_48823,N_49391);
nor UO_1618 (O_1618,N_45766,N_44143);
nor UO_1619 (O_1619,N_41372,N_48043);
and UO_1620 (O_1620,N_40050,N_48965);
or UO_1621 (O_1621,N_46042,N_46487);
and UO_1622 (O_1622,N_43773,N_42447);
xnor UO_1623 (O_1623,N_42030,N_46555);
and UO_1624 (O_1624,N_48123,N_47445);
nor UO_1625 (O_1625,N_45098,N_46073);
or UO_1626 (O_1626,N_45861,N_42024);
nor UO_1627 (O_1627,N_45339,N_40263);
xnor UO_1628 (O_1628,N_49320,N_42184);
and UO_1629 (O_1629,N_45592,N_47575);
xor UO_1630 (O_1630,N_41629,N_48741);
nor UO_1631 (O_1631,N_49267,N_47382);
nor UO_1632 (O_1632,N_49722,N_41920);
nor UO_1633 (O_1633,N_43039,N_44053);
xnor UO_1634 (O_1634,N_45147,N_40196);
and UO_1635 (O_1635,N_43120,N_47899);
xor UO_1636 (O_1636,N_46849,N_41113);
xnor UO_1637 (O_1637,N_48686,N_45730);
xnor UO_1638 (O_1638,N_45272,N_40349);
xnor UO_1639 (O_1639,N_47191,N_43812);
nand UO_1640 (O_1640,N_46720,N_44836);
nand UO_1641 (O_1641,N_46623,N_47750);
or UO_1642 (O_1642,N_45125,N_45039);
xor UO_1643 (O_1643,N_41272,N_49429);
or UO_1644 (O_1644,N_42065,N_47844);
xor UO_1645 (O_1645,N_41507,N_45739);
xor UO_1646 (O_1646,N_49065,N_40008);
or UO_1647 (O_1647,N_43352,N_47269);
nand UO_1648 (O_1648,N_49317,N_47423);
and UO_1649 (O_1649,N_46973,N_46101);
or UO_1650 (O_1650,N_40437,N_45269);
xnor UO_1651 (O_1651,N_48311,N_43693);
or UO_1652 (O_1652,N_48995,N_48749);
xnor UO_1653 (O_1653,N_42188,N_43369);
nor UO_1654 (O_1654,N_48077,N_47768);
nor UO_1655 (O_1655,N_46365,N_44272);
and UO_1656 (O_1656,N_41424,N_46817);
nor UO_1657 (O_1657,N_42865,N_40235);
nor UO_1658 (O_1658,N_46074,N_45711);
xnor UO_1659 (O_1659,N_49648,N_42317);
xnor UO_1660 (O_1660,N_45056,N_42487);
or UO_1661 (O_1661,N_40119,N_48599);
or UO_1662 (O_1662,N_47005,N_42233);
or UO_1663 (O_1663,N_48751,N_48164);
nor UO_1664 (O_1664,N_47511,N_46047);
and UO_1665 (O_1665,N_41288,N_47593);
nand UO_1666 (O_1666,N_42288,N_40956);
or UO_1667 (O_1667,N_49089,N_49952);
xor UO_1668 (O_1668,N_44485,N_47568);
nand UO_1669 (O_1669,N_47944,N_47897);
nor UO_1670 (O_1670,N_47815,N_45635);
nor UO_1671 (O_1671,N_40575,N_43911);
nand UO_1672 (O_1672,N_46545,N_48987);
nand UO_1673 (O_1673,N_48269,N_40011);
and UO_1674 (O_1674,N_46437,N_49510);
or UO_1675 (O_1675,N_46781,N_48642);
or UO_1676 (O_1676,N_48197,N_43238);
nand UO_1677 (O_1677,N_40340,N_49470);
and UO_1678 (O_1678,N_40236,N_45685);
xor UO_1679 (O_1679,N_48287,N_43326);
nor UO_1680 (O_1680,N_43760,N_42153);
nor UO_1681 (O_1681,N_49085,N_44312);
nand UO_1682 (O_1682,N_48428,N_42345);
or UO_1683 (O_1683,N_49879,N_43191);
nor UO_1684 (O_1684,N_45826,N_44664);
or UO_1685 (O_1685,N_49096,N_40170);
xnor UO_1686 (O_1686,N_40853,N_43749);
nand UO_1687 (O_1687,N_45777,N_45521);
or UO_1688 (O_1688,N_42768,N_45121);
nand UO_1689 (O_1689,N_49195,N_42784);
nor UO_1690 (O_1690,N_41300,N_43777);
or UO_1691 (O_1691,N_41733,N_47146);
and UO_1692 (O_1692,N_46021,N_44564);
xnor UO_1693 (O_1693,N_45017,N_44250);
nor UO_1694 (O_1694,N_47809,N_47836);
nor UO_1695 (O_1695,N_42776,N_47960);
and UO_1696 (O_1696,N_41205,N_44216);
xor UO_1697 (O_1697,N_41777,N_40395);
nand UO_1698 (O_1698,N_49381,N_40391);
or UO_1699 (O_1699,N_44974,N_40707);
xor UO_1700 (O_1700,N_40910,N_47971);
nand UO_1701 (O_1701,N_41620,N_46819);
nor UO_1702 (O_1702,N_40264,N_44626);
or UO_1703 (O_1703,N_48913,N_43285);
nor UO_1704 (O_1704,N_43315,N_43688);
xnor UO_1705 (O_1705,N_42396,N_49955);
and UO_1706 (O_1706,N_42157,N_41597);
nor UO_1707 (O_1707,N_46435,N_42680);
nand UO_1708 (O_1708,N_47536,N_41640);
nand UO_1709 (O_1709,N_42403,N_49039);
and UO_1710 (O_1710,N_49931,N_49163);
or UO_1711 (O_1711,N_41892,N_44228);
xnor UO_1712 (O_1712,N_44943,N_41526);
nor UO_1713 (O_1713,N_48251,N_49256);
xnor UO_1714 (O_1714,N_42328,N_49791);
or UO_1715 (O_1715,N_41446,N_43416);
nand UO_1716 (O_1716,N_42847,N_47851);
or UO_1717 (O_1717,N_43981,N_46379);
xnor UO_1718 (O_1718,N_43061,N_42364);
or UO_1719 (O_1719,N_40664,N_48550);
nand UO_1720 (O_1720,N_44844,N_44042);
xnor UO_1721 (O_1721,N_49844,N_44704);
nand UO_1722 (O_1722,N_47895,N_40392);
or UO_1723 (O_1723,N_45040,N_41046);
xnor UO_1724 (O_1724,N_40251,N_48547);
or UO_1725 (O_1725,N_46415,N_45471);
xnor UO_1726 (O_1726,N_47379,N_44789);
or UO_1727 (O_1727,N_46443,N_45348);
xnor UO_1728 (O_1728,N_47101,N_41766);
nor UO_1729 (O_1729,N_43343,N_42282);
nor UO_1730 (O_1730,N_47347,N_41565);
nor UO_1731 (O_1731,N_42513,N_43241);
nor UO_1732 (O_1732,N_45323,N_47194);
nand UO_1733 (O_1733,N_47267,N_44107);
nor UO_1734 (O_1734,N_45937,N_43565);
or UO_1735 (O_1735,N_48905,N_49287);
nor UO_1736 (O_1736,N_48786,N_48653);
nand UO_1737 (O_1737,N_49483,N_40550);
nand UO_1738 (O_1738,N_44917,N_46578);
xor UO_1739 (O_1739,N_40433,N_40188);
xor UO_1740 (O_1740,N_45660,N_44521);
and UO_1741 (O_1741,N_42082,N_41801);
and UO_1742 (O_1742,N_44321,N_40447);
nor UO_1743 (O_1743,N_49451,N_40895);
nor UO_1744 (O_1744,N_49679,N_41432);
nor UO_1745 (O_1745,N_49325,N_47996);
nor UO_1746 (O_1746,N_47061,N_42495);
nor UO_1747 (O_1747,N_49502,N_40502);
xor UO_1748 (O_1748,N_45702,N_41182);
nor UO_1749 (O_1749,N_41206,N_46190);
nor UO_1750 (O_1750,N_46406,N_42611);
xnor UO_1751 (O_1751,N_45268,N_47049);
nand UO_1752 (O_1752,N_47229,N_40213);
xor UO_1753 (O_1753,N_41089,N_47058);
and UO_1754 (O_1754,N_41025,N_44718);
or UO_1755 (O_1755,N_48024,N_41204);
nand UO_1756 (O_1756,N_46844,N_42488);
or UO_1757 (O_1757,N_45126,N_43479);
nand UO_1758 (O_1758,N_42476,N_46311);
nor UO_1759 (O_1759,N_48347,N_40492);
and UO_1760 (O_1760,N_48766,N_42696);
or UO_1761 (O_1761,N_47822,N_48425);
or UO_1762 (O_1762,N_41043,N_49639);
xor UO_1763 (O_1763,N_42804,N_42016);
nand UO_1764 (O_1764,N_47252,N_47303);
xnor UO_1765 (O_1765,N_45361,N_41191);
and UO_1766 (O_1766,N_49372,N_42876);
and UO_1767 (O_1767,N_40446,N_43576);
and UO_1768 (O_1768,N_45087,N_49102);
and UO_1769 (O_1769,N_40382,N_46768);
nor UO_1770 (O_1770,N_44303,N_42428);
or UO_1771 (O_1771,N_46890,N_45971);
or UO_1772 (O_1772,N_42533,N_49199);
xnor UO_1773 (O_1773,N_46329,N_45138);
nor UO_1774 (O_1774,N_43324,N_45398);
xnor UO_1775 (O_1775,N_40768,N_42499);
nor UO_1776 (O_1776,N_48210,N_43190);
or UO_1777 (O_1777,N_41599,N_41451);
and UO_1778 (O_1778,N_48390,N_48152);
nor UO_1779 (O_1779,N_40563,N_40249);
and UO_1780 (O_1780,N_48481,N_40524);
and UO_1781 (O_1781,N_46782,N_46199);
and UO_1782 (O_1782,N_49582,N_44764);
nor UO_1783 (O_1783,N_47430,N_41905);
nand UO_1784 (O_1784,N_47846,N_48326);
xnor UO_1785 (O_1785,N_46915,N_45714);
nor UO_1786 (O_1786,N_47129,N_40151);
or UO_1787 (O_1787,N_40863,N_46418);
nor UO_1788 (O_1788,N_45492,N_49149);
and UO_1789 (O_1789,N_40699,N_46957);
xnor UO_1790 (O_1790,N_46146,N_40242);
and UO_1791 (O_1791,N_45007,N_48810);
or UO_1792 (O_1792,N_44231,N_41924);
nor UO_1793 (O_1793,N_48454,N_48088);
and UO_1794 (O_1794,N_43657,N_40909);
nand UO_1795 (O_1795,N_47185,N_45115);
and UO_1796 (O_1796,N_46093,N_49347);
nand UO_1797 (O_1797,N_40218,N_49192);
or UO_1798 (O_1798,N_43112,N_43682);
and UO_1799 (O_1799,N_45886,N_45835);
and UO_1800 (O_1800,N_43857,N_41127);
xor UO_1801 (O_1801,N_46808,N_41956);
nand UO_1802 (O_1802,N_41982,N_48779);
nand UO_1803 (O_1803,N_48432,N_41225);
or UO_1804 (O_1804,N_46449,N_41131);
and UO_1805 (O_1805,N_40571,N_43873);
xor UO_1806 (O_1806,N_43852,N_45732);
or UO_1807 (O_1807,N_46567,N_40710);
nand UO_1808 (O_1808,N_44549,N_47100);
and UO_1809 (O_1809,N_47605,N_48926);
nand UO_1810 (O_1810,N_48185,N_42759);
nor UO_1811 (O_1811,N_49942,N_46439);
and UO_1812 (O_1812,N_46372,N_46748);
nor UO_1813 (O_1813,N_45656,N_46533);
nand UO_1814 (O_1814,N_41922,N_49926);
or UO_1815 (O_1815,N_45430,N_44951);
xor UO_1816 (O_1816,N_48794,N_43604);
nor UO_1817 (O_1817,N_43074,N_41442);
or UO_1818 (O_1818,N_43672,N_47408);
and UO_1819 (O_1819,N_47028,N_48935);
or UO_1820 (O_1820,N_42465,N_45834);
nor UO_1821 (O_1821,N_42325,N_40449);
xor UO_1822 (O_1822,N_41398,N_46496);
and UO_1823 (O_1823,N_49077,N_41954);
xnor UO_1824 (O_1824,N_44899,N_42469);
nor UO_1825 (O_1825,N_44085,N_46127);
xnor UO_1826 (O_1826,N_44175,N_41872);
xnor UO_1827 (O_1827,N_42911,N_49388);
and UO_1828 (O_1828,N_48276,N_40950);
xnor UO_1829 (O_1829,N_47859,N_44563);
or UO_1830 (O_1830,N_46481,N_48598);
nand UO_1831 (O_1831,N_44757,N_47079);
xnor UO_1832 (O_1832,N_45185,N_43735);
nor UO_1833 (O_1833,N_49585,N_49179);
nor UO_1834 (O_1834,N_47518,N_45451);
and UO_1835 (O_1835,N_48217,N_41823);
and UO_1836 (O_1836,N_49293,N_44838);
nor UO_1837 (O_1837,N_42430,N_40640);
xnor UO_1838 (O_1838,N_43748,N_45909);
or UO_1839 (O_1839,N_47900,N_41720);
and UO_1840 (O_1840,N_46843,N_43079);
nor UO_1841 (O_1841,N_40339,N_49547);
and UO_1842 (O_1842,N_45443,N_47798);
or UO_1843 (O_1843,N_41563,N_46976);
xor UO_1844 (O_1844,N_40781,N_45680);
and UO_1845 (O_1845,N_41110,N_41394);
nand UO_1846 (O_1846,N_45801,N_46850);
and UO_1847 (O_1847,N_41825,N_42819);
or UO_1848 (O_1848,N_42648,N_49744);
and UO_1849 (O_1849,N_43282,N_43045);
and UO_1850 (O_1850,N_41627,N_40697);
nor UO_1851 (O_1851,N_46350,N_48836);
nor UO_1852 (O_1852,N_42894,N_44760);
nand UO_1853 (O_1853,N_49602,N_40276);
or UO_1854 (O_1854,N_45133,N_46260);
or UO_1855 (O_1855,N_44565,N_45281);
or UO_1856 (O_1856,N_44105,N_42453);
or UO_1857 (O_1857,N_46345,N_45816);
nand UO_1858 (O_1858,N_41907,N_43848);
nor UO_1859 (O_1859,N_47643,N_42973);
or UO_1860 (O_1860,N_49119,N_41552);
xor UO_1861 (O_1861,N_42555,N_40259);
or UO_1862 (O_1862,N_49622,N_47120);
nor UO_1863 (O_1863,N_44274,N_44165);
nor UO_1864 (O_1864,N_40624,N_49594);
xnor UO_1865 (O_1865,N_44700,N_46203);
nor UO_1866 (O_1866,N_48085,N_48568);
xnor UO_1867 (O_1867,N_44656,N_44245);
xnor UO_1868 (O_1868,N_44251,N_41748);
or UO_1869 (O_1869,N_40023,N_44294);
or UO_1870 (O_1870,N_49248,N_45132);
nand UO_1871 (O_1871,N_41118,N_48315);
or UO_1872 (O_1872,N_44752,N_47242);
nor UO_1873 (O_1873,N_41661,N_48984);
nand UO_1874 (O_1874,N_45520,N_46110);
or UO_1875 (O_1875,N_41553,N_46690);
nor UO_1876 (O_1876,N_46106,N_43215);
nand UO_1877 (O_1877,N_40616,N_49516);
xor UO_1878 (O_1878,N_49427,N_40448);
and UO_1879 (O_1879,N_48194,N_47967);
or UO_1880 (O_1880,N_45069,N_45845);
and UO_1881 (O_1881,N_47050,N_43595);
or UO_1882 (O_1882,N_47459,N_40404);
xnor UO_1883 (O_1883,N_43450,N_40156);
or UO_1884 (O_1884,N_44495,N_48818);
xnor UO_1885 (O_1885,N_43754,N_41543);
and UO_1886 (O_1886,N_44713,N_48362);
nor UO_1887 (O_1887,N_40987,N_44578);
xor UO_1888 (O_1888,N_42056,N_43412);
nand UO_1889 (O_1889,N_42747,N_47339);
nor UO_1890 (O_1890,N_46340,N_44756);
xor UO_1891 (O_1891,N_45579,N_43801);
xor UO_1892 (O_1892,N_47015,N_48015);
and UO_1893 (O_1893,N_49328,N_48255);
nor UO_1894 (O_1894,N_44405,N_41362);
nor UO_1895 (O_1895,N_42515,N_42773);
or UO_1896 (O_1896,N_44093,N_46515);
or UO_1897 (O_1897,N_43962,N_48471);
xor UO_1898 (O_1898,N_43508,N_40525);
nor UO_1899 (O_1899,N_44839,N_49487);
nor UO_1900 (O_1900,N_44976,N_47635);
nor UO_1901 (O_1901,N_49588,N_43152);
xor UO_1902 (O_1902,N_48028,N_41175);
nand UO_1903 (O_1903,N_40267,N_44380);
nor UO_1904 (O_1904,N_48465,N_40063);
and UO_1905 (O_1905,N_42230,N_41220);
or UO_1906 (O_1906,N_49958,N_42996);
or UO_1907 (O_1907,N_42003,N_43805);
nand UO_1908 (O_1908,N_41296,N_41201);
or UO_1909 (O_1909,N_46940,N_42733);
xor UO_1910 (O_1910,N_48092,N_45865);
nor UO_1911 (O_1911,N_43290,N_40211);
nand UO_1912 (O_1912,N_46043,N_45282);
nor UO_1913 (O_1913,N_42622,N_44956);
nor UO_1914 (O_1914,N_45169,N_43685);
xnor UO_1915 (O_1915,N_47638,N_49881);
nand UO_1916 (O_1916,N_43492,N_49718);
and UO_1917 (O_1917,N_43208,N_44574);
nand UO_1918 (O_1918,N_44275,N_46360);
xor UO_1919 (O_1919,N_44960,N_40992);
and UO_1920 (O_1920,N_47302,N_43185);
nand UO_1921 (O_1921,N_40549,N_42435);
nand UO_1922 (O_1922,N_43881,N_49230);
nand UO_1923 (O_1923,N_42871,N_48438);
nand UO_1924 (O_1924,N_49650,N_46595);
and UO_1925 (O_1925,N_41580,N_41952);
nor UO_1926 (O_1926,N_43096,N_46586);
and UO_1927 (O_1927,N_49091,N_49555);
and UO_1928 (O_1928,N_43478,N_48144);
nor UO_1929 (O_1929,N_46661,N_43907);
and UO_1930 (O_1930,N_47442,N_41738);
or UO_1931 (O_1931,N_44695,N_46492);
nor UO_1932 (O_1932,N_49014,N_44698);
or UO_1933 (O_1933,N_43845,N_41484);
nor UO_1934 (O_1934,N_46087,N_47071);
nand UO_1935 (O_1935,N_43385,N_45402);
nand UO_1936 (O_1936,N_46201,N_41208);
xnor UO_1937 (O_1937,N_42706,N_43418);
and UO_1938 (O_1938,N_47081,N_42537);
and UO_1939 (O_1939,N_41598,N_42301);
or UO_1940 (O_1940,N_49432,N_47608);
nand UO_1941 (O_1941,N_48699,N_45815);
and UO_1942 (O_1942,N_40990,N_46179);
nor UO_1943 (O_1943,N_48444,N_43329);
or UO_1944 (O_1944,N_48038,N_46971);
nor UO_1945 (O_1945,N_42921,N_43537);
or UO_1946 (O_1946,N_48464,N_46429);
nand UO_1947 (O_1947,N_44680,N_46221);
nand UO_1948 (O_1948,N_43598,N_46523);
nand UO_1949 (O_1949,N_49512,N_44295);
or UO_1950 (O_1950,N_47485,N_42035);
xor UO_1951 (O_1951,N_40928,N_46085);
and UO_1952 (O_1952,N_44744,N_46704);
or UO_1953 (O_1953,N_44681,N_44347);
xnor UO_1954 (O_1954,N_49527,N_43482);
nand UO_1955 (O_1955,N_42146,N_44477);
xnor UO_1956 (O_1956,N_40068,N_49105);
or UO_1957 (O_1957,N_42924,N_47419);
and UO_1958 (O_1958,N_40045,N_42849);
or UO_1959 (O_1959,N_43081,N_45566);
xor UO_1960 (O_1960,N_47173,N_42162);
nand UO_1961 (O_1961,N_40945,N_49180);
xnor UO_1962 (O_1962,N_46944,N_40260);
nor UO_1963 (O_1963,N_42185,N_43770);
or UO_1964 (O_1964,N_44895,N_47343);
or UO_1965 (O_1965,N_43821,N_47868);
xor UO_1966 (O_1966,N_46308,N_43275);
nand UO_1967 (O_1967,N_40542,N_40949);
or UO_1968 (O_1968,N_44317,N_42614);
nand UO_1969 (O_1969,N_40167,N_49858);
or UO_1970 (O_1970,N_41985,N_46276);
nor UO_1971 (O_1971,N_45241,N_43916);
or UO_1972 (O_1972,N_42672,N_41793);
nor UO_1973 (O_1973,N_40884,N_48611);
xor UO_1974 (O_1974,N_46070,N_49950);
or UO_1975 (O_1975,N_46453,N_40493);
or UO_1976 (O_1976,N_48892,N_40517);
or UO_1977 (O_1977,N_42851,N_41472);
and UO_1978 (O_1978,N_40546,N_47702);
nand UO_1979 (O_1979,N_49056,N_46639);
or UO_1980 (O_1980,N_43970,N_45253);
or UO_1981 (O_1981,N_41498,N_45611);
xor UO_1982 (O_1982,N_41192,N_47195);
nand UO_1983 (O_1983,N_42066,N_45997);
or UO_1984 (O_1984,N_40661,N_48897);
nand UO_1985 (O_1985,N_44311,N_42593);
nor UO_1986 (O_1986,N_45137,N_43896);
xor UO_1987 (O_1987,N_40555,N_47902);
and UO_1988 (O_1988,N_47272,N_49276);
xor UO_1989 (O_1989,N_46722,N_49977);
and UO_1990 (O_1990,N_42540,N_42235);
or UO_1991 (O_1991,N_49551,N_48902);
nand UO_1992 (O_1992,N_44517,N_48631);
and UO_1993 (O_1993,N_47275,N_41587);
and UO_1994 (O_1994,N_48803,N_44559);
and UO_1995 (O_1995,N_46988,N_44853);
nand UO_1996 (O_1996,N_41454,N_48998);
nor UO_1997 (O_1997,N_46699,N_48633);
nor UO_1998 (O_1998,N_46746,N_47406);
nand UO_1999 (O_1999,N_46205,N_40894);
nor UO_2000 (O_2000,N_42216,N_49590);
nor UO_2001 (O_2001,N_48040,N_45508);
nand UO_2002 (O_2002,N_47903,N_42509);
nand UO_2003 (O_2003,N_44753,N_43200);
or UO_2004 (O_2004,N_49335,N_45594);
or UO_2005 (O_2005,N_41020,N_45640);
and UO_2006 (O_2006,N_40592,N_42091);
nand UO_2007 (O_2007,N_47932,N_48084);
nand UO_2008 (O_2008,N_43534,N_41178);
or UO_2009 (O_2009,N_41813,N_44130);
xor UO_2010 (O_2010,N_41925,N_44996);
nand UO_2011 (O_2011,N_47525,N_44871);
nor UO_2012 (O_2012,N_47561,N_47241);
or UO_2013 (O_2013,N_49795,N_41539);
nand UO_2014 (O_2014,N_45479,N_43567);
nand UO_2015 (O_2015,N_41759,N_47169);
and UO_2016 (O_2016,N_48542,N_41050);
xnor UO_2017 (O_2017,N_42379,N_47273);
nor UO_2018 (O_2018,N_40948,N_42419);
or UO_2019 (O_2019,N_48694,N_46121);
or UO_2020 (O_2020,N_43929,N_47170);
xor UO_2021 (O_2021,N_48883,N_47946);
or UO_2022 (O_2022,N_46031,N_47175);
nor UO_2023 (O_2023,N_43361,N_46227);
nand UO_2024 (O_2024,N_44634,N_49239);
or UO_2025 (O_2025,N_43643,N_49450);
xnor UO_2026 (O_2026,N_40692,N_48671);
nand UO_2027 (O_2027,N_43884,N_45536);
xor UO_2028 (O_2028,N_47369,N_45897);
and UO_2029 (O_2029,N_44724,N_44969);
nand UO_2030 (O_2030,N_49216,N_42209);
nor UO_2031 (O_2031,N_41977,N_45096);
or UO_2032 (O_2032,N_46018,N_43833);
nor UO_2033 (O_2033,N_47436,N_43382);
nor UO_2034 (O_2034,N_44239,N_44299);
or UO_2035 (O_2035,N_41945,N_44412);
or UO_2036 (O_2036,N_41698,N_49948);
xor UO_2037 (O_2037,N_43915,N_41669);
nand UO_2038 (O_2038,N_45362,N_41505);
or UO_2039 (O_2039,N_42427,N_46912);
nand UO_2040 (O_2040,N_46230,N_47853);
and UO_2041 (O_2041,N_44308,N_47234);
nor UO_2042 (O_2042,N_40279,N_45550);
and UO_2043 (O_2043,N_42214,N_40878);
or UO_2044 (O_2044,N_40734,N_45283);
or UO_2045 (O_2045,N_42807,N_47943);
or UO_2046 (O_2046,N_43202,N_49653);
or UO_2047 (O_2047,N_41542,N_40870);
and UO_2048 (O_2048,N_41941,N_46225);
and UO_2049 (O_2049,N_40650,N_43317);
nand UO_2050 (O_2050,N_42239,N_49572);
and UO_2051 (O_2051,N_47642,N_46300);
or UO_2052 (O_2052,N_44300,N_47251);
and UO_2053 (O_2053,N_43518,N_43446);
nor UO_2054 (O_2054,N_42564,N_48554);
or UO_2055 (O_2055,N_40797,N_40189);
nor UO_2056 (O_2056,N_44459,N_42351);
xnor UO_2057 (O_2057,N_40513,N_43464);
nand UO_2058 (O_2058,N_44646,N_46828);
or UO_2059 (O_2059,N_46666,N_47063);
or UO_2060 (O_2060,N_49747,N_44052);
or UO_2061 (O_2061,N_41604,N_46556);
nand UO_2062 (O_2062,N_42468,N_46286);
and UO_2063 (O_2063,N_41251,N_41281);
and UO_2064 (O_2064,N_46364,N_44596);
and UO_2065 (O_2065,N_49344,N_42368);
and UO_2066 (O_2066,N_48777,N_40590);
or UO_2067 (O_2067,N_42330,N_44060);
xnor UO_2068 (O_2068,N_44390,N_47773);
and UO_2069 (O_2069,N_40700,N_41263);
xnor UO_2070 (O_2070,N_49296,N_47726);
or UO_2071 (O_2071,N_43692,N_46797);
nand UO_2072 (O_2072,N_41899,N_46030);
xnor UO_2073 (O_2073,N_49322,N_46891);
nand UO_2074 (O_2074,N_49257,N_47610);
nand UO_2075 (O_2075,N_45538,N_47601);
nor UO_2076 (O_2076,N_40229,N_48712);
nor UO_2077 (O_2077,N_48521,N_44058);
and UO_2078 (O_2078,N_48540,N_48768);
nor UO_2079 (O_2079,N_49389,N_42786);
and UO_2080 (O_2080,N_44126,N_48724);
nor UO_2081 (O_2081,N_44825,N_44407);
and UO_2082 (O_2082,N_45747,N_41677);
xnor UO_2083 (O_2083,N_45235,N_49182);
or UO_2084 (O_2084,N_49339,N_47718);
nor UO_2085 (O_2085,N_44225,N_41912);
or UO_2086 (O_2086,N_42835,N_47918);
or UO_2087 (O_2087,N_47901,N_41126);
or UO_2088 (O_2088,N_43697,N_46907);
nor UO_2089 (O_2089,N_44616,N_45049);
nand UO_2090 (O_2090,N_45141,N_45486);
xnor UO_2091 (O_2091,N_46696,N_43599);
or UO_2092 (O_2092,N_47715,N_40791);
and UO_2093 (O_2093,N_44436,N_47447);
and UO_2094 (O_2094,N_41264,N_43127);
and UO_2095 (O_2095,N_41258,N_41256);
or UO_2096 (O_2096,N_43870,N_43424);
nor UO_2097 (O_2097,N_44319,N_45562);
and UO_2098 (O_2098,N_40649,N_44008);
and UO_2099 (O_2099,N_40029,N_42703);
and UO_2100 (O_2100,N_41174,N_47747);
nor UO_2101 (O_2101,N_49943,N_46444);
and UO_2102 (O_2102,N_44036,N_41423);
nor UO_2103 (O_2103,N_42676,N_41459);
or UO_2104 (O_2104,N_47324,N_45406);
and UO_2105 (O_2105,N_40789,N_41349);
or UO_2106 (O_2106,N_44902,N_42661);
nand UO_2107 (O_2107,N_43360,N_43153);
nor UO_2108 (O_2108,N_43946,N_46738);
nand UO_2109 (O_2109,N_40803,N_40714);
xnor UO_2110 (O_2110,N_49214,N_44017);
xnor UO_2111 (O_2111,N_43432,N_47444);
or UO_2112 (O_2112,N_43586,N_42439);
xor UO_2113 (O_2113,N_48802,N_48400);
nand UO_2114 (O_2114,N_42206,N_43622);
xor UO_2115 (O_2115,N_40230,N_41993);
nor UO_2116 (O_2116,N_43188,N_43509);
nand UO_2117 (O_2117,N_47712,N_49875);
nor UO_2118 (O_2118,N_44046,N_48134);
nand UO_2119 (O_2119,N_49503,N_45291);
xor UO_2120 (O_2120,N_40535,N_40099);
xor UO_2121 (O_2121,N_44077,N_42898);
xnor UO_2122 (O_2122,N_47752,N_40851);
or UO_2123 (O_2123,N_41585,N_46017);
nor UO_2124 (O_2124,N_48294,N_47144);
xor UO_2125 (O_2125,N_44342,N_47800);
xnor UO_2126 (O_2126,N_48713,N_48738);
and UO_2127 (O_2127,N_46568,N_46457);
xnor UO_2128 (O_2128,N_45615,N_44767);
nor UO_2129 (O_2129,N_45048,N_45574);
and UO_2130 (O_2130,N_40963,N_44824);
and UO_2131 (O_2131,N_43199,N_42901);
nand UO_2132 (O_2132,N_46430,N_49583);
nor UO_2133 (O_2133,N_40890,N_47226);
nand UO_2134 (O_2134,N_46620,N_49458);
and UO_2135 (O_2135,N_48674,N_41729);
or UO_2136 (O_2136,N_47537,N_44349);
or UO_2137 (O_2137,N_44693,N_41636);
nor UO_2138 (O_2138,N_41479,N_48209);
nor UO_2139 (O_2139,N_48003,N_49265);
or UO_2140 (O_2140,N_43341,N_43940);
or UO_2141 (O_2141,N_41913,N_40047);
and UO_2142 (O_2142,N_48575,N_46574);
and UO_2143 (O_2143,N_49161,N_44447);
nor UO_2144 (O_2144,N_45633,N_42628);
nor UO_2145 (O_2145,N_47141,N_42536);
nor UO_2146 (O_2146,N_43328,N_45336);
nor UO_2147 (O_2147,N_48583,N_43067);
and UO_2148 (O_2148,N_40337,N_45895);
nor UO_2149 (O_2149,N_46503,N_49366);
or UO_2150 (O_2150,N_48512,N_48388);
xnor UO_2151 (O_2151,N_45570,N_45622);
xnor UO_2152 (O_2152,N_45514,N_40117);
nor UO_2153 (O_2153,N_45518,N_47268);
and UO_2154 (O_2154,N_40275,N_44707);
or UO_2155 (O_2155,N_40149,N_49987);
or UO_2156 (O_2156,N_41328,N_43022);
and UO_2157 (O_2157,N_48577,N_40197);
nand UO_2158 (O_2158,N_49020,N_42012);
nand UO_2159 (O_2159,N_49310,N_49507);
or UO_2160 (O_2160,N_48868,N_48146);
xnor UO_2161 (O_2161,N_46273,N_46769);
xor UO_2162 (O_2162,N_45530,N_47528);
nor UO_2163 (O_2163,N_41233,N_48662);
nor UO_2164 (O_2164,N_47789,N_47713);
and UO_2165 (O_2165,N_45092,N_49656);
or UO_2166 (O_2166,N_41082,N_48310);
and UO_2167 (O_2167,N_43403,N_48668);
xor UO_2168 (O_2168,N_41783,N_41142);
and UO_2169 (O_2169,N_40049,N_45817);
xnor UO_2170 (O_2170,N_44233,N_48737);
nor UO_2171 (O_2171,N_49023,N_42335);
or UO_2172 (O_2172,N_42657,N_49035);
nand UO_2173 (O_2173,N_49135,N_40210);
and UO_2174 (O_2174,N_41833,N_44855);
or UO_2175 (O_2175,N_46628,N_48238);
xor UO_2176 (O_2176,N_45947,N_48073);
and UO_2177 (O_2177,N_42284,N_42138);
and UO_2178 (O_2178,N_43456,N_45797);
and UO_2179 (O_2179,N_45509,N_46866);
nand UO_2180 (O_2180,N_46877,N_47054);
nor UO_2181 (O_2181,N_49008,N_45429);
or UO_2182 (O_2182,N_41965,N_41471);
and UO_2183 (O_2183,N_40377,N_46058);
or UO_2184 (O_2184,N_42743,N_48391);
xor UO_2185 (O_2185,N_41826,N_47948);
or UO_2186 (O_2186,N_40618,N_44333);
or UO_2187 (O_2187,N_47082,N_46786);
or UO_2188 (O_2188,N_43957,N_42005);
nand UO_2189 (O_2189,N_45382,N_46414);
xor UO_2190 (O_2190,N_44535,N_46883);
xor UO_2191 (O_2191,N_49246,N_42318);
or UO_2192 (O_2192,N_45210,N_44979);
nor UO_2193 (O_2193,N_41408,N_45639);
xnor UO_2194 (O_2194,N_46288,N_44782);
nor UO_2195 (O_2195,N_40924,N_40560);
nand UO_2196 (O_2196,N_43989,N_44972);
nor UO_2197 (O_2197,N_42980,N_44688);
xor UO_2198 (O_2198,N_45631,N_44415);
nand UO_2199 (O_2199,N_40342,N_43901);
or UO_2200 (O_2200,N_49918,N_44340);
nand UO_2201 (O_2201,N_47962,N_46322);
and UO_2202 (O_2202,N_47563,N_43558);
xnor UO_2203 (O_2203,N_47483,N_42324);
xnor UO_2204 (O_2204,N_43141,N_46742);
nand UO_2205 (O_2205,N_49895,N_46079);
and UO_2206 (O_2206,N_48877,N_44434);
or UO_2207 (O_2207,N_46495,N_48980);
and UO_2208 (O_2208,N_42338,N_40141);
and UO_2209 (O_2209,N_45650,N_40848);
or UO_2210 (O_2210,N_44118,N_46336);
and UO_2211 (O_2211,N_46864,N_41856);
or UO_2212 (O_2212,N_44265,N_42541);
nand UO_2213 (O_2213,N_43800,N_47629);
nand UO_2214 (O_2214,N_46540,N_46631);
and UO_2215 (O_2215,N_40184,N_43555);
or UO_2216 (O_2216,N_43922,N_44803);
nand UO_2217 (O_2217,N_48563,N_46534);
and UO_2218 (O_2218,N_42044,N_41086);
xnor UO_2219 (O_2219,N_40192,N_49550);
or UO_2220 (O_2220,N_48107,N_43105);
nor UO_2221 (O_2221,N_47426,N_49529);
and UO_2222 (O_2222,N_48176,N_43013);
and UO_2223 (O_2223,N_46408,N_43277);
xnor UO_2224 (O_2224,N_43034,N_41774);
or UO_2225 (O_2225,N_42623,N_43699);
or UO_2226 (O_2226,N_43480,N_43961);
and UO_2227 (O_2227,N_45026,N_44537);
or UO_2228 (O_2228,N_47656,N_49505);
xor UO_2229 (O_2229,N_41397,N_49125);
nand UO_2230 (O_2230,N_44332,N_41583);
and UO_2231 (O_2231,N_45122,N_48191);
and UO_2232 (O_2232,N_40455,N_48501);
and UO_2233 (O_2233,N_48709,N_47669);
nor UO_2234 (O_2234,N_41951,N_45252);
nand UO_2235 (O_2235,N_43472,N_49700);
xnor UO_2236 (O_2236,N_46142,N_43769);
and UO_2237 (O_2237,N_44171,N_44478);
xnor UO_2238 (O_2238,N_45694,N_46387);
and UO_2239 (O_2239,N_43965,N_46122);
or UO_2240 (O_2240,N_48198,N_40552);
xor UO_2241 (O_2241,N_41443,N_46245);
and UO_2242 (O_2242,N_45383,N_45569);
nand UO_2243 (O_2243,N_47383,N_49713);
nor UO_2244 (O_2244,N_41226,N_48558);
or UO_2245 (O_2245,N_45888,N_48848);
and UO_2246 (O_2246,N_42922,N_43976);
or UO_2247 (O_2247,N_41827,N_43399);
or UO_2248 (O_2248,N_45317,N_40519);
or UO_2249 (O_2249,N_40567,N_48975);
xor UO_2250 (O_2250,N_47233,N_44431);
and UO_2251 (O_2251,N_42986,N_41449);
and UO_2252 (O_2252,N_48567,N_44292);
nand UO_2253 (O_2253,N_41806,N_40426);
or UO_2254 (O_2254,N_48118,N_47067);
xnor UO_2255 (O_2255,N_42033,N_42208);
and UO_2256 (O_2256,N_49442,N_46594);
and UO_2257 (O_2257,N_48458,N_43101);
or UO_2258 (O_2258,N_49083,N_41340);
nor UO_2259 (O_2259,N_44648,N_44010);
nand UO_2260 (O_2260,N_45869,N_49170);
and UO_2261 (O_2261,N_48313,N_41006);
or UO_2262 (O_2262,N_43471,N_40073);
nand UO_2263 (O_2263,N_47407,N_42172);
and UO_2264 (O_2264,N_44785,N_44306);
nor UO_2265 (O_2265,N_42409,N_46593);
nor UO_2266 (O_2266,N_45614,N_48213);
and UO_2267 (O_2267,N_47098,N_43596);
or UO_2268 (O_2268,N_45129,N_41119);
and UO_2269 (O_2269,N_46513,N_40538);
nor UO_2270 (O_2270,N_40355,N_47062);
and UO_2271 (O_2271,N_43437,N_44361);
or UO_2272 (O_2272,N_49862,N_44702);
nor UO_2273 (O_2273,N_43714,N_48485);
and UO_2274 (O_2274,N_49283,N_41310);
xnor UO_2275 (O_2275,N_48413,N_41144);
xnor UO_2276 (O_2276,N_45666,N_44222);
xor UO_2277 (O_2277,N_45501,N_45000);
nand UO_2278 (O_2278,N_42660,N_42959);
and UO_2279 (O_2279,N_46115,N_46592);
xor UO_2280 (O_2280,N_43895,N_45325);
nand UO_2281 (O_2281,N_43221,N_40807);
nor UO_2282 (O_2282,N_40922,N_41336);
or UO_2283 (O_2283,N_47720,N_46669);
nor UO_2284 (O_2284,N_41385,N_43322);
or UO_2285 (O_2285,N_41403,N_46224);
and UO_2286 (O_2286,N_40146,N_40609);
nor UO_2287 (O_2287,N_47366,N_47818);
nor UO_2288 (O_2288,N_41188,N_49407);
or UO_2289 (O_2289,N_44614,N_49053);
or UO_2290 (O_2290,N_49990,N_48115);
nand UO_2291 (O_2291,N_47942,N_41942);
nor UO_2292 (O_2292,N_49229,N_45541);
or UO_2293 (O_2293,N_46324,N_43300);
or UO_2294 (O_2294,N_48747,N_41348);
or UO_2295 (O_2295,N_43483,N_48762);
nand UO_2296 (O_2296,N_44305,N_40595);
or UO_2297 (O_2297,N_42311,N_43359);
nor UO_2298 (O_2298,N_40298,N_47312);
xor UO_2299 (O_2299,N_47313,N_49781);
nor UO_2300 (O_2300,N_40417,N_42413);
nand UO_2301 (O_2301,N_40964,N_41716);
xor UO_2302 (O_2302,N_48559,N_47460);
or UO_2303 (O_2303,N_47087,N_41576);
xor UO_2304 (O_2304,N_43924,N_44701);
and UO_2305 (O_2305,N_40370,N_41567);
nor UO_2306 (O_2306,N_44697,N_41490);
nor UO_2307 (O_2307,N_48952,N_41634);
or UO_2308 (O_2308,N_49289,N_45686);
or UO_2309 (O_2309,N_40485,N_44983);
nor UO_2310 (O_2310,N_48263,N_47640);
nor UO_2311 (O_2311,N_48635,N_49454);
nand UO_2312 (O_2312,N_48423,N_49601);
nand UO_2313 (O_2313,N_40927,N_44226);
nand UO_2314 (O_2314,N_44290,N_42530);
nand UO_2315 (O_2315,N_46086,N_44740);
xor UO_2316 (O_2316,N_44199,N_48207);
and UO_2317 (O_2317,N_43213,N_44425);
and UO_2318 (O_2318,N_48863,N_48885);
xnor UO_2319 (O_2319,N_41575,N_42727);
and UO_2320 (O_2320,N_48452,N_43484);
nor UO_2321 (O_2321,N_48735,N_47529);
nand UO_2322 (O_2322,N_45943,N_41750);
xor UO_2323 (O_2323,N_42150,N_42300);
and UO_2324 (O_2324,N_44877,N_47869);
nand UO_2325 (O_2325,N_48658,N_44066);
and UO_2326 (O_2326,N_45320,N_40253);
or UO_2327 (O_2327,N_41829,N_43240);
and UO_2328 (O_2328,N_45052,N_49688);
nand UO_2329 (O_2329,N_46436,N_48372);
or UO_2330 (O_2330,N_48946,N_49805);
nor UO_2331 (O_2331,N_41194,N_44891);
xnor UO_2332 (O_2332,N_47157,N_44513);
and UO_2333 (O_2333,N_44435,N_45692);
or UO_2334 (O_2334,N_42599,N_49819);
nand UO_2335 (O_2335,N_40341,N_40527);
nand UO_2336 (O_2336,N_40969,N_49846);
nand UO_2337 (O_2337,N_41002,N_43651);
nand UO_2338 (O_2338,N_49657,N_43377);
or UO_2339 (O_2339,N_43487,N_42048);
xor UO_2340 (O_2340,N_46675,N_48574);
and UO_2341 (O_2341,N_45094,N_45810);
nor UO_2342 (O_2342,N_45475,N_45082);
and UO_2343 (O_2343,N_45394,N_49198);
or UO_2344 (O_2344,N_47827,N_42007);
or UO_2345 (O_2345,N_43914,N_42148);
nand UO_2346 (O_2346,N_41842,N_49687);
nor UO_2347 (O_2347,N_49353,N_40613);
nand UO_2348 (O_2348,N_43592,N_45346);
nand UO_2349 (O_2349,N_46034,N_49238);
nand UO_2350 (O_2350,N_40319,N_49467);
or UO_2351 (O_2351,N_44453,N_48252);
and UO_2352 (O_2352,N_41838,N_45857);
nand UO_2353 (O_2353,N_44169,N_43076);
xor UO_2354 (O_2354,N_48808,N_49126);
nand UO_2355 (O_2355,N_43979,N_44409);
nand UO_2356 (O_2356,N_42662,N_47150);
xor UO_2357 (O_2357,N_44819,N_49495);
and UO_2358 (O_2358,N_42339,N_41755);
and UO_2359 (O_2359,N_41478,N_46213);
nand UO_2360 (O_2360,N_41528,N_44240);
nand UO_2361 (O_2361,N_49562,N_48764);
or UO_2362 (O_2362,N_43987,N_46967);
nor UO_2363 (O_2363,N_43842,N_46362);
or UO_2364 (O_2364,N_48880,N_43142);
or UO_2365 (O_2365,N_47887,N_40054);
xor UO_2366 (O_2366,N_44313,N_46477);
nor UO_2367 (O_2367,N_46716,N_48519);
or UO_2368 (O_2368,N_49261,N_47032);
nand UO_2369 (O_2369,N_47064,N_48613);
nand UO_2370 (O_2370,N_44694,N_44140);
and UO_2371 (O_2371,N_47714,N_48159);
nor UO_2372 (O_2372,N_43503,N_41266);
xnor UO_2373 (O_2373,N_44597,N_43827);
and UO_2374 (O_2374,N_45168,N_43706);
xor UO_2375 (O_2375,N_40096,N_45197);
nor UO_2376 (O_2376,N_44997,N_46514);
nand UO_2377 (O_2377,N_41646,N_44314);
xor UO_2378 (O_2378,N_40923,N_42480);
nand UO_2379 (O_2379,N_45099,N_44723);
and UO_2380 (O_2380,N_44658,N_44708);
or UO_2381 (O_2381,N_43219,N_41939);
or UO_2382 (O_2382,N_41014,N_49478);
or UO_2383 (O_2383,N_45221,N_49323);
nor UO_2384 (O_2384,N_40866,N_45716);
nor UO_2385 (O_2385,N_42815,N_44444);
xnor UO_2386 (O_2386,N_45636,N_48218);
nand UO_2387 (O_2387,N_48314,N_44147);
nand UO_2388 (O_2388,N_49185,N_43376);
and UO_2389 (O_2389,N_43608,N_41369);
and UO_2390 (O_2390,N_46299,N_48105);
nor UO_2391 (O_2391,N_42147,N_48100);
nand UO_2392 (O_2392,N_40324,N_44301);
or UO_2393 (O_2393,N_48468,N_48627);
nor UO_2394 (O_2394,N_48302,N_44024);
or UO_2395 (O_2395,N_40974,N_42503);
or UO_2396 (O_2396,N_45481,N_49078);
or UO_2397 (O_2397,N_45065,N_42966);
or UO_2398 (O_2398,N_49966,N_48610);
or UO_2399 (O_2399,N_40885,N_46752);
and UO_2400 (O_2400,N_49392,N_44622);
nor UO_2401 (O_2401,N_44676,N_44577);
nand UO_2402 (O_2402,N_40056,N_49311);
nand UO_2403 (O_2403,N_42821,N_43836);
and UO_2404 (O_2404,N_45433,N_43589);
nor UO_2405 (O_2405,N_46078,N_40730);
xor UO_2406 (O_2406,N_40780,N_40255);
nand UO_2407 (O_2407,N_44078,N_42595);
nor UO_2408 (O_2408,N_47558,N_40228);
xor UO_2409 (O_2409,N_47427,N_49571);
or UO_2410 (O_2410,N_43078,N_43055);
or UO_2411 (O_2411,N_42928,N_43689);
nand UO_2412 (O_2412,N_48873,N_44146);
or UO_2413 (O_2413,N_41185,N_46488);
xor UO_2414 (O_2414,N_42738,N_40566);
or UO_2415 (O_2415,N_42063,N_48404);
and UO_2416 (O_2416,N_42885,N_46717);
or UO_2417 (O_2417,N_42908,N_43844);
or UO_2418 (O_2418,N_45453,N_46511);
and UO_2419 (O_2419,N_47624,N_41157);
and UO_2420 (O_2420,N_42691,N_40795);
and UO_2421 (O_2421,N_48377,N_44474);
and UO_2422 (O_2422,N_47433,N_44812);
or UO_2423 (O_2423,N_46602,N_44476);
xnor UO_2424 (O_2424,N_43731,N_43046);
or UO_2425 (O_2425,N_48914,N_48163);
nand UO_2426 (O_2426,N_47263,N_43830);
and UO_2427 (O_2427,N_40142,N_40899);
nor UO_2428 (O_2428,N_40597,N_43139);
xor UO_2429 (O_2429,N_48900,N_45182);
and UO_2430 (O_2430,N_42380,N_45421);
nor UO_2431 (O_2431,N_44922,N_44510);
or UO_2432 (O_2432,N_45949,N_42224);
nand UO_2433 (O_2433,N_41465,N_48412);
xor UO_2434 (O_2434,N_41332,N_40424);
nor UO_2435 (O_2435,N_42271,N_49779);
xor UO_2436 (O_2436,N_40385,N_44621);
and UO_2437 (O_2437,N_46491,N_45646);
nor UO_2438 (O_2438,N_45029,N_46767);
or UO_2439 (O_2439,N_43701,N_41027);
or UO_2440 (O_2440,N_40774,N_42519);
nand UO_2441 (O_2441,N_43785,N_48371);
xor UO_2442 (O_2442,N_47283,N_47135);
xnor UO_2443 (O_2443,N_42713,N_41211);
nand UO_2444 (O_2444,N_40097,N_49682);
nand UO_2445 (O_2445,N_47751,N_43033);
xor UO_2446 (O_2446,N_42305,N_47443);
nor UO_2447 (O_2447,N_49273,N_46925);
xor UO_2448 (O_2448,N_48443,N_46498);
or UO_2449 (O_2449,N_49045,N_44993);
nor UO_2450 (O_2450,N_42105,N_49298);
and UO_2451 (O_2451,N_43092,N_41606);
nand UO_2452 (O_2452,N_46581,N_45837);
xor UO_2453 (O_2453,N_47239,N_48483);
nand UO_2454 (O_2454,N_46766,N_43837);
and UO_2455 (O_2455,N_46560,N_48014);
xor UO_2456 (O_2456,N_46792,N_48293);
or UO_2457 (O_2457,N_40764,N_41489);
or UO_2458 (O_2458,N_42049,N_47489);
nand UO_2459 (O_2459,N_40178,N_48887);
nand UO_2460 (O_2460,N_46464,N_49204);
nand UO_2461 (O_2461,N_43026,N_49677);
nand UO_2462 (O_2462,N_49753,N_44519);
or UO_2463 (O_2463,N_42749,N_40334);
and UO_2464 (O_2464,N_45181,N_46039);
or UO_2465 (O_2465,N_40646,N_49134);
nor UO_2466 (O_2466,N_45742,N_48142);
nand UO_2467 (O_2467,N_40463,N_44547);
and UO_2468 (O_2468,N_49034,N_47122);
and UO_2469 (O_2469,N_40132,N_44649);
xnor UO_2470 (O_2470,N_48270,N_41031);
nand UO_2471 (O_2471,N_41860,N_48325);
and UO_2472 (O_2472,N_49365,N_48624);
nor UO_2473 (O_2473,N_46249,N_46798);
nor UO_2474 (O_2474,N_47573,N_49737);
xnor UO_2475 (O_2475,N_44083,N_47413);
and UO_2476 (O_2476,N_49587,N_42585);
or UO_2477 (O_2477,N_46762,N_49189);
nor UO_2478 (O_2478,N_44858,N_40412);
nand UO_2479 (O_2479,N_45364,N_43137);
and UO_2480 (O_2480,N_41083,N_44348);
nand UO_2481 (O_2481,N_49659,N_46082);
or UO_2482 (O_2482,N_46402,N_47056);
and UO_2483 (O_2483,N_43775,N_49812);
nand UO_2484 (O_2484,N_47596,N_46176);
xnor UO_2485 (O_2485,N_47839,N_41756);
or UO_2486 (O_2486,N_41039,N_42582);
xor UO_2487 (O_2487,N_46008,N_41063);
and UO_2488 (O_2488,N_40865,N_46630);
and UO_2489 (O_2489,N_42884,N_43037);
xor UO_2490 (O_2490,N_46905,N_45783);
xor UO_2491 (O_2491,N_49693,N_47189);
nor UO_2492 (O_2492,N_48045,N_45708);
nor UO_2493 (O_2493,N_43302,N_46721);
and UO_2494 (O_2494,N_46107,N_46812);
nor UO_2495 (O_2495,N_42591,N_43912);
nand UO_2496 (O_2496,N_40886,N_41413);
or UO_2497 (O_2497,N_44582,N_44653);
nand UO_2498 (O_2498,N_49251,N_43829);
nand UO_2499 (O_2499,N_49160,N_43281);
and UO_2500 (O_2500,N_47925,N_43117);
and UO_2501 (O_2501,N_43457,N_40897);
xor UO_2502 (O_2502,N_40687,N_46659);
nand UO_2503 (O_2503,N_41875,N_44903);
nand UO_2504 (O_2504,N_44615,N_41943);
and UO_2505 (O_2505,N_44362,N_46810);
and UO_2506 (O_2506,N_40698,N_43582);
or UO_2507 (O_2507,N_47912,N_48449);
nand UO_2508 (O_2508,N_43145,N_42154);
and UO_2509 (O_2509,N_48537,N_42782);
nor UO_2510 (O_2510,N_42970,N_48441);
or UO_2511 (O_2511,N_44137,N_44158);
xnor UO_2512 (O_2512,N_49802,N_46740);
nand UO_2513 (O_2513,N_49069,N_45709);
nand UO_2514 (O_2514,N_40362,N_45770);
or UO_2515 (O_2515,N_45617,N_48236);
or UO_2516 (O_2516,N_40239,N_49963);
or UO_2517 (O_2517,N_42113,N_42081);
and UO_2518 (O_2518,N_43559,N_47510);
or UO_2519 (O_2519,N_40407,N_48451);
nor UO_2520 (O_2520,N_41848,N_49878);
xnor UO_2521 (O_2521,N_48114,N_41494);
xor UO_2522 (O_2522,N_44689,N_43630);
xnor UO_2523 (O_2523,N_40414,N_43708);
or UO_2524 (O_2524,N_46111,N_40484);
xnor UO_2525 (O_2525,N_44247,N_47861);
or UO_2526 (O_2526,N_41009,N_43410);
nand UO_2527 (O_2527,N_41073,N_45806);
nand UO_2528 (O_2528,N_44633,N_41699);
nor UO_2529 (O_2529,N_41603,N_46827);
xor UO_2530 (O_2530,N_43438,N_45953);
nand UO_2531 (O_2531,N_43721,N_45632);
or UO_2532 (O_2532,N_45180,N_49475);
or UO_2533 (O_2533,N_46672,N_48771);
nand UO_2534 (O_2534,N_40620,N_40356);
or UO_2535 (O_2535,N_46676,N_49742);
nand UO_2536 (O_2536,N_41237,N_41005);
or UO_2537 (O_2537,N_40937,N_44932);
nand UO_2538 (O_2538,N_47450,N_44886);
and UO_2539 (O_2539,N_48544,N_49818);
nand UO_2540 (O_2540,N_49120,N_43296);
nand UO_2541 (O_2541,N_43170,N_41166);
nand UO_2542 (O_2542,N_40982,N_49698);
or UO_2543 (O_2543,N_47548,N_47631);
and UO_2544 (O_2544,N_41224,N_44737);
and UO_2545 (O_2545,N_42526,N_43441);
nor UO_2546 (O_2546,N_46020,N_49983);
nor UO_2547 (O_2547,N_44837,N_45036);
or UO_2548 (O_2548,N_46239,N_47539);
and UO_2549 (O_2549,N_47926,N_44482);
or UO_2550 (O_2550,N_45288,N_40846);
nand UO_2551 (O_2551,N_40471,N_41107);
and UO_2552 (O_2552,N_44020,N_45577);
xnor UO_2553 (O_2553,N_41269,N_48878);
xnor UO_2554 (O_2554,N_41187,N_48435);
nand UO_2555 (O_2555,N_42950,N_45737);
xor UO_2556 (O_2556,N_41638,N_45266);
or UO_2557 (O_2557,N_41937,N_40114);
nand UO_2558 (O_2558,N_40742,N_48933);
nand UO_2559 (O_2559,N_46154,N_48793);
nor UO_2560 (O_2560,N_45544,N_40507);
nand UO_2561 (O_2561,N_44772,N_41666);
nor UO_2562 (O_2562,N_48334,N_47310);
xor UO_2563 (O_2563,N_49079,N_46320);
xor UO_2564 (O_2564,N_48679,N_41784);
and UO_2565 (O_2565,N_44985,N_48272);
or UO_2566 (O_2566,N_43292,N_41728);
nor UO_2567 (O_2567,N_40183,N_48063);
nand UO_2568 (O_2568,N_45838,N_42932);
xor UO_2569 (O_2569,N_47172,N_49854);
or UO_2570 (O_2570,N_49449,N_41799);
nor UO_2571 (O_2571,N_47471,N_44788);
nand UO_2572 (O_2572,N_41662,N_48181);
or UO_2573 (O_2573,N_48728,N_49924);
nor UO_2574 (O_2574,N_42750,N_41600);
and UO_2575 (O_2575,N_43602,N_44809);
nand UO_2576 (O_2576,N_40061,N_40310);
or UO_2577 (O_2577,N_44418,N_42504);
nand UO_2578 (O_2578,N_43176,N_47924);
xnor UO_2579 (O_2579,N_48614,N_46120);
nand UO_2580 (O_2580,N_44280,N_44781);
nand UO_2581 (O_2581,N_49300,N_49569);
or UO_2582 (O_2582,N_47886,N_45894);
xor UO_2583 (O_2583,N_47289,N_48267);
nor UO_2584 (O_2584,N_40318,N_47554);
or UO_2585 (O_2585,N_42177,N_45002);
nand UO_2586 (O_2586,N_44081,N_49888);
or UO_2587 (O_2587,N_45066,N_44406);
nand UO_2588 (O_2588,N_45604,N_41334);
nor UO_2589 (O_2589,N_49128,N_48548);
nor UO_2590 (O_2590,N_44092,N_49789);
or UO_2591 (O_2591,N_43293,N_40365);
and UO_2592 (O_2592,N_46882,N_41259);
and UO_2593 (O_2593,N_48010,N_46128);
nand UO_2594 (O_2594,N_40185,N_47484);
nand UO_2595 (O_2595,N_44450,N_42636);
nor UO_2596 (O_2596,N_45023,N_46283);
or UO_2597 (O_2597,N_43452,N_45110);
and UO_2598 (O_2598,N_41980,N_46134);
and UO_2599 (O_2599,N_45447,N_43927);
nor UO_2600 (O_2600,N_47961,N_41026);
and UO_2601 (O_2601,N_45573,N_44832);
or UO_2602 (O_2602,N_47775,N_49108);
xnor UO_2603 (O_2603,N_42191,N_41555);
and UO_2604 (O_2604,N_40443,N_48352);
nand UO_2605 (O_2605,N_48775,N_40512);
or UO_2606 (O_2606,N_44338,N_44181);
and UO_2607 (O_2607,N_41155,N_43447);
xor UO_2608 (O_2608,N_41053,N_45043);
and UO_2609 (O_2609,N_46424,N_48720);
or UO_2610 (O_2610,N_40545,N_47258);
and UO_2611 (O_2611,N_49616,N_41125);
and UO_2612 (O_2612,N_44457,N_49015);
xnor UO_2613 (O_2613,N_43276,N_46216);
and UO_2614 (O_2614,N_47287,N_44848);
nand UO_2615 (O_2615,N_40481,N_41616);
xnor UO_2616 (O_2616,N_48408,N_47409);
and UO_2617 (O_2617,N_45788,N_40366);
or UO_2618 (O_2618,N_42873,N_46133);
nand UO_2619 (O_2619,N_43411,N_46549);
nor UO_2620 (O_2620,N_44766,N_45020);
or UO_2621 (O_2621,N_42852,N_44401);
and UO_2622 (O_2622,N_44606,N_47840);
nand UO_2623 (O_2623,N_46057,N_48733);
and UO_2624 (O_2624,N_40893,N_46758);
and UO_2625 (O_2625,N_49568,N_45091);
nand UO_2626 (O_2626,N_43928,N_45349);
or UO_2627 (O_2627,N_49423,N_42392);
nand UO_2628 (O_2628,N_45183,N_49532);
xor UO_2629 (O_2629,N_44771,N_48050);
xor UO_2630 (O_2630,N_49410,N_41992);
nand UO_2631 (O_2631,N_46902,N_47316);
xnor UO_2632 (O_2632,N_43966,N_47816);
nand UO_2633 (O_2633,N_49425,N_44841);
xnor UO_2634 (O_2634,N_47012,N_45005);
nor UO_2635 (O_2635,N_49603,N_49723);
nor UO_2636 (O_2636,N_40688,N_48367);
nand UO_2637 (O_2637,N_41963,N_48226);
nand UO_2638 (O_2638,N_45395,N_42721);
xnor UO_2639 (O_2639,N_43991,N_42047);
nor UO_2640 (O_2640,N_45578,N_45670);
nor UO_2641 (O_2641,N_48110,N_48147);
nand UO_2642 (O_2642,N_48150,N_47274);
nor UO_2643 (O_2643,N_48727,N_48087);
and UO_2644 (O_2644,N_46541,N_48609);
or UO_2645 (O_2645,N_41450,N_41253);
xnor UO_2646 (O_2646,N_49418,N_40153);
or UO_2647 (O_2647,N_43294,N_43365);
and UO_2648 (O_2648,N_41503,N_44167);
xnor UO_2649 (O_2649,N_48815,N_48791);
and UO_2650 (O_2650,N_42789,N_40587);
nor UO_2651 (O_2651,N_44428,N_40757);
or UO_2652 (O_2652,N_44070,N_44687);
nor UO_2653 (O_2653,N_44076,N_45201);
and UO_2654 (O_2654,N_46519,N_44384);
and UO_2655 (O_2655,N_49049,N_44263);
nand UO_2656 (O_2656,N_47695,N_47648);
or UO_2657 (O_2657,N_41909,N_47102);
nand UO_2658 (O_2658,N_48167,N_46287);
and UO_2659 (O_2659,N_46266,N_43591);
or UO_2660 (O_2660,N_48355,N_40187);
xnor UO_2661 (O_2661,N_49146,N_49525);
or UO_2662 (O_2662,N_46749,N_40874);
xor UO_2663 (O_2663,N_47743,N_45690);
and UO_2664 (O_2664,N_42542,N_42834);
nor UO_2665 (O_2665,N_43656,N_42720);
and UO_2666 (O_2666,N_49028,N_42552);
nor UO_2667 (O_2667,N_47008,N_41988);
and UO_2668 (O_2668,N_49613,N_47113);
and UO_2669 (O_2669,N_46438,N_40758);
or UO_2670 (O_2670,N_46731,N_46775);
nand UO_2671 (O_2671,N_42514,N_43764);
xnor UO_2672 (O_2672,N_49566,N_45877);
and UO_2673 (O_2673,N_46832,N_41881);
or UO_2674 (O_2674,N_44743,N_44377);
and UO_2675 (O_2675,N_44268,N_43846);
or UO_2676 (O_2676,N_44923,N_42984);
nand UO_2677 (O_2677,N_45720,N_40548);
nand UO_2678 (O_2678,N_40118,N_47749);
or UO_2679 (O_2679,N_48380,N_40107);
nor UO_2680 (O_2680,N_42972,N_49534);
nand UO_2681 (O_2681,N_49412,N_41399);
nand UO_2682 (O_2682,N_40131,N_41121);
and UO_2683 (O_2683,N_45192,N_48875);
and UO_2684 (O_2684,N_41438,N_45824);
nand UO_2685 (O_2685,N_47858,N_45418);
xnor UO_2686 (O_2686,N_47466,N_48838);
xor UO_2687 (O_2687,N_47745,N_40518);
and UO_2688 (O_2688,N_40919,N_48983);
nand UO_2689 (O_2689,N_45113,N_49211);
and UO_2690 (O_2690,N_48298,N_49772);
xor UO_2691 (O_2691,N_48332,N_47819);
or UO_2692 (O_2692,N_43932,N_42398);
and UO_2693 (O_2693,N_48993,N_44717);
nor UO_2694 (O_2694,N_44641,N_49842);
nor UO_2695 (O_2695,N_40491,N_44576);
xnor UO_2696 (O_2696,N_40130,N_41049);
nor UO_2697 (O_2697,N_48493,N_48976);
xor UO_2698 (O_2698,N_43123,N_44579);
nand UO_2699 (O_2699,N_45549,N_42767);
nor UO_2700 (O_2700,N_42204,N_40082);
nand UO_2701 (O_2701,N_44229,N_45456);
xnor UO_2702 (O_2702,N_44019,N_40906);
or UO_2703 (O_2703,N_43696,N_44015);
or UO_2704 (O_2704,N_40822,N_46671);
nand UO_2705 (O_2705,N_47266,N_43734);
or UO_2706 (O_2706,N_41084,N_49006);
and UO_2707 (O_2707,N_41685,N_46710);
or UO_2708 (O_2708,N_43626,N_47618);
and UO_2709 (O_2709,N_46467,N_46218);
nand UO_2710 (O_2710,N_48054,N_46777);
and UO_2711 (O_2711,N_49835,N_45275);
or UO_2712 (O_2712,N_47295,N_47123);
nor UO_2713 (O_2713,N_43849,N_40722);
and UO_2714 (O_2714,N_45195,N_42861);
nand UO_2715 (O_2715,N_42285,N_49665);
xnor UO_2716 (O_2716,N_41172,N_40776);
nand UO_2717 (O_2717,N_45695,N_43239);
xor UO_2718 (O_2718,N_45363,N_41887);
nand UO_2719 (O_2719,N_42046,N_46051);
or UO_2720 (O_2720,N_42360,N_46267);
nand UO_2721 (O_2721,N_48053,N_42261);
and UO_2722 (O_2722,N_48189,N_46044);
or UO_2723 (O_2723,N_46006,N_43181);
nor UO_2724 (O_2724,N_43521,N_40968);
and UO_2725 (O_2725,N_46892,N_42101);
nor UO_2726 (O_2726,N_45757,N_43270);
xor UO_2727 (O_2727,N_46442,N_40202);
and UO_2728 (O_2728,N_41683,N_46370);
or UO_2729 (O_2729,N_42780,N_45131);
nand UO_2730 (O_2730,N_40576,N_42038);
nor UO_2731 (O_2731,N_40072,N_45211);
and UO_2732 (O_2732,N_44866,N_40705);
and UO_2733 (O_2733,N_40396,N_41711);
or UO_2734 (O_2734,N_40122,N_49058);
xor UO_2735 (O_2735,N_46202,N_46380);
xnor UO_2736 (O_2736,N_44327,N_46193);
and UO_2737 (O_2737,N_41581,N_42149);
nand UO_2738 (O_2738,N_41068,N_48931);
or UO_2739 (O_2739,N_49517,N_40304);
or UO_2740 (O_2740,N_42401,N_40171);
or UO_2741 (O_2741,N_47978,N_47678);
or UO_2742 (O_2742,N_44727,N_49290);
or UO_2743 (O_2743,N_49822,N_41351);
and UO_2744 (O_2744,N_43491,N_40026);
nor UO_2745 (O_2745,N_42385,N_48986);
xnor UO_2746 (O_2746,N_46821,N_47387);
nand UO_2747 (O_2747,N_46460,N_43814);
nand UO_2748 (O_2748,N_48358,N_40301);
or UO_2749 (O_2749,N_48641,N_49815);
and UO_2750 (O_2750,N_42656,N_49326);
or UO_2751 (O_2751,N_42286,N_48065);
and UO_2752 (O_2752,N_43018,N_48161);
and UO_2753 (O_2753,N_44928,N_45068);
and UO_2754 (O_2754,N_42304,N_42093);
xor UO_2755 (O_2755,N_42737,N_42510);
or UO_2756 (O_2756,N_47655,N_42525);
and UO_2757 (O_2757,N_40648,N_42869);
nor UO_2758 (O_2758,N_40514,N_43283);
nand UO_2759 (O_2759,N_48296,N_47244);
nand UO_2760 (O_2760,N_43941,N_47632);
xor UO_2761 (O_2761,N_49370,N_47820);
nor UO_2762 (O_2762,N_40612,N_44190);
xor UO_2763 (O_2763,N_47048,N_42394);
or UO_2764 (O_2764,N_46297,N_49400);
nor UO_2765 (O_2765,N_41548,N_47042);
and UO_2766 (O_2766,N_41111,N_48169);
nand UO_2767 (O_2767,N_47609,N_40328);
or UO_2768 (O_2768,N_44644,N_44675);
nand UO_2769 (O_2769,N_47730,N_48496);
nor UO_2770 (O_2770,N_49234,N_45469);
xnor UO_2771 (O_2771,N_47154,N_47393);
and UO_2772 (O_2772,N_43640,N_42697);
and UO_2773 (O_2773,N_42709,N_41491);
xnor UO_2774 (O_2774,N_43536,N_42268);
xnor UO_2775 (O_2775,N_49749,N_48467);
xor UO_2776 (O_2776,N_45315,N_49978);
nor UO_2777 (O_2777,N_41882,N_44745);
and UO_2778 (O_2778,N_42376,N_41919);
xor UO_2779 (O_2779,N_49101,N_42806);
nand UO_2780 (O_2780,N_48669,N_44777);
nor UO_2781 (O_2781,N_47787,N_44867);
and UO_2782 (O_2782,N_48538,N_45274);
xnor UO_2783 (O_2783,N_41849,N_47845);
nand UO_2784 (O_2784,N_42569,N_41055);
or UO_2785 (O_2785,N_48606,N_40905);
nor UO_2786 (O_2786,N_49707,N_44049);
nor UO_2787 (O_2787,N_47270,N_44014);
and UO_2788 (O_2788,N_44037,N_44975);
xnor UO_2789 (O_2789,N_47288,N_43569);
and UO_2790 (O_2790,N_45190,N_43744);
xor UO_2791 (O_2791,N_43709,N_43177);
nand UO_2792 (O_2792,N_45717,N_43393);
xnor UO_2793 (O_2793,N_41976,N_47597);
nor UO_2794 (O_2794,N_43044,N_43173);
nor UO_2795 (O_2795,N_42649,N_43351);
nor UO_2796 (O_2796,N_43363,N_47035);
xor UO_2797 (O_2797,N_42678,N_49903);
xnor UO_2798 (O_2798,N_41305,N_49331);
nand UO_2799 (O_2799,N_41339,N_41219);
and UO_2800 (O_2800,N_40887,N_43694);
and UO_2801 (O_2801,N_43571,N_44569);
and UO_2802 (O_2802,N_47078,N_44148);
xor UO_2803 (O_2803,N_47716,N_45795);
nand UO_2804 (O_2804,N_49087,N_40939);
or UO_2805 (O_2805,N_44962,N_43261);
or UO_2806 (O_2806,N_47697,N_42805);
and UO_2807 (O_2807,N_41317,N_48715);
nor UO_2808 (O_2808,N_48170,N_48281);
nand UO_2809 (O_2809,N_47327,N_47761);
nand UO_2810 (O_2810,N_42462,N_46450);
nor UO_2811 (O_2811,N_45254,N_40580);
xnor UO_2812 (O_2812,N_47760,N_44331);
xor UO_2813 (O_2813,N_44500,N_45103);
xor UO_2814 (O_2814,N_48407,N_42308);
nand UO_2815 (O_2815,N_49202,N_43541);
xor UO_2816 (O_2816,N_46071,N_48060);
xnor UO_2817 (O_2817,N_47357,N_48486);
and UO_2818 (O_2818,N_44209,N_42372);
nor UO_2819 (O_2819,N_45158,N_40633);
nand UO_2820 (O_2820,N_42708,N_41210);
and UO_2821 (O_2821,N_45059,N_43002);
xnor UO_2822 (O_2822,N_48042,N_42017);
or UO_2823 (O_2823,N_40829,N_46919);
and UO_2824 (O_2824,N_49828,N_43271);
nor UO_2825 (O_2825,N_47034,N_41897);
and UO_2826 (O_2826,N_48422,N_46315);
nand UO_2827 (O_2827,N_48862,N_47521);
xnor UO_2828 (O_2828,N_40946,N_44172);
and UO_2829 (O_2829,N_43702,N_41418);
nand UO_2830 (O_2830,N_49054,N_43776);
or UO_2831 (O_2831,N_46756,N_44783);
or UO_2832 (O_2832,N_45929,N_41901);
nand UO_2833 (O_2833,N_45627,N_44168);
nor UO_2834 (O_2834,N_48736,N_45152);
or UO_2835 (O_2835,N_46262,N_41483);
xnor UO_2836 (O_2836,N_46138,N_49785);
and UO_2837 (O_2837,N_45866,N_45446);
nor UO_2838 (O_2838,N_45551,N_49099);
or UO_2839 (O_2839,N_46404,N_44595);
nand UO_2840 (O_2840,N_43624,N_48460);
nor UO_2841 (O_2841,N_49154,N_47235);
and UO_2842 (O_2842,N_43875,N_41329);
or UO_2843 (O_2843,N_49673,N_45391);
nand UO_2844 (O_2844,N_44768,N_40747);
nor UO_2845 (O_2845,N_41139,N_44383);
or UO_2846 (O_2846,N_49321,N_47205);
or UO_2847 (O_2847,N_49477,N_49387);
xor UO_2848 (O_2848,N_49433,N_43068);
and UO_2849 (O_2849,N_46911,N_43461);
or UO_2850 (O_2850,N_48566,N_46028);
nand UO_2851 (O_2851,N_47930,N_45057);
or UO_2852 (O_2852,N_46867,N_41787);
nand UO_2853 (O_2853,N_46396,N_42824);
and UO_2854 (O_2854,N_48994,N_41768);
or UO_2855 (O_2855,N_47872,N_40801);
nand UO_2856 (O_2856,N_45233,N_44749);
xnor UO_2857 (O_2857,N_44375,N_44153);
nand UO_2858 (O_2858,N_44628,N_43964);
and UO_2859 (O_2859,N_45762,N_46836);
or UO_2860 (O_2860,N_40010,N_45931);
nand UO_2861 (O_2861,N_49499,N_44846);
and UO_2862 (O_2862,N_48619,N_47284);
and UO_2863 (O_2863,N_46271,N_45628);
nor UO_2864 (O_2864,N_44878,N_40643);
and UO_2865 (O_2865,N_43974,N_49408);
nand UO_2866 (O_2866,N_43588,N_48420);
and UO_2867 (O_2867,N_41007,N_45458);
or UO_2868 (O_2868,N_41893,N_44100);
nand UO_2869 (O_2869,N_46054,N_49855);
xnor UO_2870 (O_2870,N_47854,N_44055);
xor UO_2871 (O_2871,N_43245,N_40368);
or UO_2872 (O_2872,N_40303,N_40850);
nor UO_2873 (O_2873,N_40831,N_44088);
and UO_2874 (O_2874,N_42001,N_49166);
or UO_2875 (O_2875,N_46874,N_41693);
nand UO_2876 (O_2876,N_47121,N_42029);
nor UO_2877 (O_2877,N_49830,N_44636);
and UO_2878 (O_2878,N_42071,N_47956);
xnor UO_2879 (O_2879,N_41154,N_45917);
or UO_2880 (O_2880,N_46886,N_48498);
xor UO_2881 (O_2881,N_49164,N_49443);
or UO_2882 (O_2882,N_45913,N_47658);
or UO_2883 (O_2883,N_49438,N_41650);
or UO_2884 (O_2884,N_48847,N_45529);
xor UO_2885 (O_2885,N_46654,N_42715);
and UO_2886 (O_2886,N_42236,N_41917);
nand UO_2887 (O_2887,N_46826,N_42348);
nand UO_2888 (O_2888,N_46066,N_49133);
nand UO_2889 (O_2889,N_40827,N_49302);
xnor UO_2890 (O_2890,N_41883,N_49994);
xor UO_2891 (O_2891,N_40478,N_47014);
nand UO_2892 (O_2892,N_42309,N_42139);
nor UO_2893 (O_2893,N_41935,N_43939);
or UO_2894 (O_2894,N_48969,N_49838);
and UO_2895 (O_2895,N_47788,N_43116);
nand UO_2896 (O_2896,N_46677,N_48035);
and UO_2897 (O_2897,N_46471,N_49352);
or UO_2898 (O_2898,N_45388,N_45450);
nor UO_2899 (O_2899,N_42353,N_47569);
nor UO_2900 (O_2900,N_47514,N_49000);
and UO_2901 (O_2901,N_46922,N_47555);
nor UO_2902 (O_2902,N_44522,N_42002);
and UO_2903 (O_2903,N_40383,N_46851);
xnor UO_2904 (O_2904,N_43774,N_46342);
or UO_2905 (O_2905,N_44761,N_42060);
or UO_2906 (O_2906,N_40606,N_48809);
xor UO_2907 (O_2907,N_45222,N_44208);
and UO_2908 (O_2908,N_40602,N_46036);
and UO_2909 (O_2909,N_42057,N_45638);
or UO_2910 (O_2910,N_46389,N_48373);
and UO_2911 (O_2911,N_42212,N_49864);
nand UO_2912 (O_2912,N_40544,N_42277);
or UO_2913 (O_2913,N_49357,N_44982);
nor UO_2914 (O_2914,N_46700,N_41866);
xnor UO_2915 (O_2915,N_40292,N_40051);
or UO_2916 (O_2916,N_44683,N_43373);
or UO_2917 (O_2917,N_45511,N_48518);
and UO_2918 (O_2918,N_46447,N_45911);
and UO_2919 (O_2919,N_41248,N_46382);
nor UO_2920 (O_2920,N_49057,N_40840);
or UO_2921 (O_2921,N_46325,N_46219);
nor UO_2922 (O_2922,N_46046,N_46732);
nor UO_2923 (O_2923,N_40025,N_49937);
nand UO_2924 (O_2924,N_43985,N_40737);
or UO_2925 (O_2925,N_40052,N_42064);
or UO_2926 (O_2926,N_42128,N_47797);
and UO_2927 (O_2927,N_40679,N_40427);
xnor UO_2928 (O_2928,N_43736,N_48636);
or UO_2929 (O_2929,N_48602,N_41436);
xnor UO_2930 (O_2930,N_43784,N_48333);
nand UO_2931 (O_2931,N_46337,N_45672);
xor UO_2932 (O_2932,N_40540,N_45705);
xnor UO_2933 (O_2933,N_44096,N_49869);
and UO_2934 (O_2934,N_45585,N_46284);
and UO_2935 (O_2935,N_41718,N_41830);
nor UO_2936 (O_2936,N_43378,N_48693);
nand UO_2937 (O_2937,N_48729,N_44462);
nor UO_2938 (O_2938,N_41522,N_44104);
xnor UO_2939 (O_2939,N_41781,N_44720);
or UO_2940 (O_2940,N_48979,N_42490);
xnor UO_2941 (O_2941,N_40676,N_44205);
xnor UO_2942 (O_2942,N_41303,N_42092);
nand UO_2943 (O_2943,N_41129,N_49787);
nand UO_2944 (O_2944,N_47719,N_46104);
nor UO_2945 (O_2945,N_48950,N_45080);
or UO_2946 (O_2946,N_49274,N_42273);
nor UO_2947 (O_2947,N_43859,N_45860);
and UO_2948 (O_2948,N_42935,N_49303);
or UO_2949 (O_2949,N_44254,N_46573);
nand UO_2950 (O_2950,N_43733,N_40336);
nand UO_2951 (O_2951,N_44746,N_41252);
xnor UO_2952 (O_2952,N_49671,N_44086);
and UO_2953 (O_2953,N_44802,N_45477);
nand UO_2954 (O_2954,N_43725,N_45657);
nand UO_2955 (O_2955,N_47696,N_46950);
or UO_2956 (O_2956,N_40027,N_41694);
or UO_2957 (O_2957,N_49100,N_48629);
and UO_2958 (O_2958,N_44080,N_43660);
nor UO_2959 (O_2959,N_46368,N_46062);
nand UO_2960 (O_2960,N_47464,N_48612);
or UO_2961 (O_2961,N_46056,N_45380);
xor UO_2962 (O_2962,N_49599,N_46223);
or UO_2963 (O_2963,N_42900,N_46197);
or UO_2964 (O_2964,N_44739,N_44721);
and UO_2965 (O_2965,N_40483,N_41143);
or UO_2966 (O_2966,N_41284,N_43490);
or UO_2967 (O_2967,N_42760,N_45967);
and UO_2968 (O_2968,N_42455,N_43913);
xnor UO_2969 (O_2969,N_45358,N_43893);
nand UO_2970 (O_2970,N_45554,N_47346);
and UO_2971 (O_2971,N_49872,N_42854);
nor UO_2972 (O_2972,N_47428,N_49905);
xnor UO_2973 (O_2973,N_46664,N_43053);
or UO_2974 (O_2974,N_44413,N_42925);
nand UO_2975 (O_2975,N_43422,N_42112);
nor UO_2976 (O_2976,N_46881,N_45575);
or UO_2977 (O_2977,N_40875,N_40436);
xnor UO_2978 (O_2978,N_42724,N_49738);
and UO_2979 (O_2979,N_42640,N_49646);
or UO_2980 (O_2980,N_44189,N_47572);
xnor UO_2981 (O_2981,N_48389,N_49011);
nand UO_2982 (O_2982,N_40017,N_44344);
or UO_2983 (O_2983,N_41101,N_48784);
xor UO_2984 (O_2984,N_45994,N_42719);
nand UO_2985 (O_2985,N_43107,N_42655);
nor UO_2986 (O_2986,N_48337,N_43984);
or UO_2987 (O_2987,N_42248,N_42547);
xnor UO_2988 (O_2988,N_44094,N_41577);
or UO_2989 (O_2989,N_47995,N_46482);
nand UO_2990 (O_2990,N_43909,N_40287);
xor UO_2991 (O_2991,N_40346,N_49005);
or UO_2992 (O_2992,N_48230,N_40808);
xnor UO_2993 (O_2993,N_49221,N_45440);
or UO_2994 (O_2994,N_42830,N_46546);
xnor UO_2995 (O_2995,N_45745,N_46952);
or UO_2996 (O_2996,N_48630,N_49243);
or UO_2997 (O_2997,N_42639,N_46508);
nor UO_2998 (O_2998,N_47520,N_42000);
xnor UO_2999 (O_2999,N_49060,N_42993);
nand UO_3000 (O_3000,N_48660,N_40217);
nand UO_3001 (O_3001,N_40629,N_47297);
nand UO_3002 (O_3002,N_49374,N_47674);
and UO_3003 (O_3003,N_44807,N_49138);
nand UO_3004 (O_3004,N_47188,N_42050);
xnor UO_3005 (O_3005,N_40021,N_44651);
or UO_3006 (O_3006,N_44787,N_40039);
or UO_3007 (O_3007,N_45217,N_48827);
nand UO_3008 (O_3008,N_48681,N_43758);
nor UO_3009 (O_3009,N_46041,N_40908);
xor UO_3010 (O_3010,N_40763,N_48864);
xor UO_3011 (O_3011,N_43111,N_42704);
or UO_3012 (O_3012,N_49771,N_41152);
nor UO_3013 (O_3013,N_42084,N_41626);
nand UO_3014 (O_3014,N_49373,N_49253);
xnor UO_3015 (O_3015,N_47394,N_40881);
or UO_3016 (O_3016,N_46840,N_46518);
nor UO_3017 (O_3017,N_41150,N_45701);
nor UO_3018 (O_3018,N_47177,N_47201);
or UO_3019 (O_3019,N_40871,N_42961);
or UO_3020 (O_3020,N_45559,N_47708);
and UO_3021 (O_3021,N_43115,N_40250);
xor UO_3022 (O_3022,N_43023,N_44099);
xnor UO_3023 (O_3023,N_44920,N_48584);
and UO_3024 (O_3024,N_48821,N_42201);
xnor UO_3025 (O_3025,N_43006,N_42400);
nand UO_3026 (O_3026,N_44479,N_43259);
and UO_3027 (O_3027,N_45952,N_41405);
nand UO_3028 (O_3028,N_49746,N_48290);
or UO_3029 (O_3029,N_43043,N_40796);
or UO_3030 (O_3030,N_45928,N_41314);
and UO_3031 (O_3031,N_44942,N_46914);
or UO_3032 (O_3032,N_46870,N_46035);
and UO_3033 (O_3033,N_40543,N_49241);
and UO_3034 (O_3034,N_42506,N_46936);
xor UO_3035 (O_3035,N_42960,N_43556);
or UO_3036 (O_3036,N_42431,N_42061);
or UO_3037 (O_3037,N_45959,N_48473);
nor UO_3038 (O_3038,N_47190,N_47735);
xor UO_3039 (O_3039,N_40696,N_49796);
nor UO_3040 (O_3040,N_44966,N_46214);
and UO_3041 (O_3041,N_42578,N_48981);
or UO_3042 (O_3042,N_45173,N_41968);
or UO_3043 (O_3043,N_41393,N_42452);
nor UO_3044 (O_3044,N_49363,N_48318);
nand UO_3045 (O_3045,N_48697,N_47013);
nand UO_3046 (O_3046,N_48516,N_45434);
xor UO_3047 (O_3047,N_48177,N_43700);
and UO_3048 (O_3048,N_49493,N_48279);
xor UO_3049 (O_3049,N_41797,N_40547);
nor UO_3050 (O_3050,N_44273,N_48184);
nand UO_3051 (O_3051,N_44796,N_41681);
nand UO_3052 (O_3052,N_40852,N_40891);
nor UO_3053 (O_3053,N_42620,N_41052);
nand UO_3054 (O_3054,N_46486,N_42532);
and UO_3055 (O_3055,N_48955,N_48482);
nand UO_3056 (O_3056,N_43165,N_46702);
nor UO_3057 (O_3057,N_47360,N_42748);
or UO_3058 (O_3058,N_47088,N_43906);
or UO_3059 (O_3059,N_40998,N_42040);
and UO_3060 (O_3060,N_47504,N_45497);
xor UO_3061 (O_3061,N_42979,N_41270);
nand UO_3062 (O_3062,N_45664,N_48813);
nand UO_3063 (O_3063,N_41123,N_45899);
and UO_3064 (O_3064,N_49223,N_44472);
or UO_3065 (O_3065,N_41944,N_40647);
nor UO_3066 (O_3066,N_41406,N_46794);
or UO_3067 (O_3067,N_47325,N_44731);
or UO_3068 (O_3068,N_45448,N_47915);
xnor UO_3069 (O_3069,N_48079,N_41461);
nor UO_3070 (O_3070,N_42638,N_45825);
nand UO_3071 (O_3071,N_42039,N_43311);
and UO_3072 (O_3072,N_46900,N_44686);
and UO_3073 (O_3073,N_46272,N_44714);
and UO_3074 (O_3074,N_48942,N_44061);
and UO_3075 (O_3075,N_42651,N_40925);
nand UO_3076 (O_3076,N_45707,N_48030);
nand UO_3077 (O_3077,N_43347,N_47331);
nor UO_3078 (O_3078,N_41695,N_42464);
and UO_3079 (O_3079,N_48944,N_43113);
nand UO_3080 (O_3080,N_49867,N_41923);
nand UO_3081 (O_3081,N_44497,N_48922);
nand UO_3082 (O_3082,N_43057,N_46941);
xnor UO_3083 (O_3083,N_47701,N_46480);
xor UO_3084 (O_3084,N_47376,N_46837);
nand UO_3085 (O_3085,N_42291,N_48722);
xnor UO_3086 (O_3086,N_48135,N_41592);
xnor UO_3087 (O_3087,N_42108,N_43394);
nor UO_3088 (O_3088,N_43262,N_44163);
xor UO_3089 (O_3089,N_43747,N_47385);
nand UO_3090 (O_3090,N_47260,N_49940);
and UO_3091 (O_3091,N_47665,N_44538);
nor UO_3092 (O_3092,N_41556,N_42785);
or UO_3093 (O_3093,N_42644,N_42358);
xor UO_3094 (O_3094,N_46027,N_40076);
or UO_3095 (O_3095,N_49730,N_45591);
or UO_3096 (O_3096,N_49421,N_43648);
nor UO_3097 (O_3097,N_44449,N_46562);
nand UO_3098 (O_3098,N_41138,N_46094);
xor UO_3099 (O_3099,N_49845,N_43415);
xnor UO_3100 (O_3100,N_49836,N_49435);
or UO_3101 (O_3101,N_49219,N_49711);
xor UO_3102 (O_3102,N_48499,N_45396);
nand UO_3103 (O_3103,N_48125,N_45015);
and UO_3104 (O_3104,N_47291,N_48243);
xor UO_3105 (O_3105,N_43333,N_46923);
and UO_3106 (O_3106,N_49927,N_44410);
or UO_3107 (O_3107,N_41280,N_45546);
nor UO_3108 (O_3108,N_48057,N_48634);
nand UO_3109 (O_3109,N_46160,N_45156);
nand UO_3110 (O_3110,N_40805,N_42772);
and UO_3111 (O_3111,N_48936,N_40615);
nand UO_3112 (O_3112,N_40837,N_45973);
or UO_3113 (O_3113,N_40006,N_46723);
and UO_3114 (O_3114,N_41276,N_40354);
xor UO_3115 (O_3115,N_48421,N_45498);
nand UO_3116 (O_3116,N_48106,N_48046);
nand UO_3117 (O_3117,N_47781,N_48011);
nor UO_3118 (O_3118,N_46363,N_41057);
nor UO_3119 (O_3119,N_41455,N_46691);
or UO_3120 (O_3120,N_40461,N_40603);
nor UO_3121 (O_3121,N_44001,N_40359);
and UO_3122 (O_3122,N_45072,N_43839);
and UO_3123 (O_3123,N_42647,N_43723);
and UO_3124 (O_3124,N_48509,N_40769);
nor UO_3125 (O_3125,N_43498,N_42249);
and UO_3126 (O_3126,N_47728,N_48416);
xnor UO_3127 (O_3127,N_41497,N_43631);
nand UO_3128 (O_3128,N_49481,N_43958);
xor UO_3129 (O_3129,N_49605,N_44532);
or UO_3130 (O_3130,N_49804,N_44659);
and UO_3131 (O_3131,N_41710,N_45603);
or UO_3132 (O_3132,N_48909,N_45435);
nand UO_3133 (O_3133,N_40432,N_45873);
and UO_3134 (O_3134,N_46789,N_45267);
xnor UO_3135 (O_3135,N_40245,N_43716);
or UO_3136 (O_3136,N_40215,N_48090);
and UO_3137 (O_3137,N_42802,N_46455);
nor UO_3138 (O_3138,N_47876,N_47562);
nand UO_3139 (O_3139,N_44068,N_48224);
nor UO_3140 (O_3140,N_40040,N_47003);
nand UO_3141 (O_3141,N_47294,N_46889);
or UO_3142 (O_3142,N_46468,N_48774);
nor UO_3143 (O_3143,N_48649,N_46989);
nand UO_3144 (O_3144,N_45047,N_42862);
and UO_3145 (O_3145,N_48433,N_42995);
nor UO_3146 (O_3146,N_44729,N_45619);
or UO_3147 (O_3147,N_41697,N_48851);
xor UO_3148 (O_3148,N_43704,N_41731);
nor UO_3149 (O_3149,N_46899,N_46393);
and UO_3150 (O_3150,N_44371,N_45645);
or UO_3151 (O_3151,N_40888,N_42557);
and UO_3152 (O_3152,N_47981,N_47699);
and UO_3153 (O_3153,N_40144,N_43476);
xor UO_3154 (O_3154,N_41028,N_49825);
nor UO_3155 (O_3155,N_44684,N_46755);
nand UO_3156 (O_3156,N_40997,N_47326);
nor UO_3157 (O_3157,N_47318,N_48939);
xnor UO_3158 (O_3158,N_44446,N_46376);
nand UO_3159 (O_3159,N_46879,N_48988);
nor UO_3160 (O_3160,N_40498,N_46149);
nand UO_3161 (O_3161,N_43168,N_44411);
xor UO_3162 (O_3162,N_43230,N_41862);
xnor UO_3163 (O_3163,N_45996,N_43087);
nand UO_3164 (O_3164,N_46476,N_48497);
or UO_3165 (O_3165,N_45078,N_45404);
or UO_3166 (O_3166,N_48305,N_44404);
nand UO_3167 (O_3167,N_41308,N_46917);
nor UO_3168 (O_3168,N_45089,N_46857);
and UO_3169 (O_3169,N_41590,N_44369);
or UO_3170 (O_3170,N_45675,N_43644);
xnor UO_3171 (O_3171,N_40694,N_41386);
and UO_3172 (O_3172,N_45792,N_46088);
nor UO_3173 (O_3173,N_47500,N_42245);
xnor UO_3174 (O_3174,N_44242,N_43167);
and UO_3175 (O_3175,N_40630,N_49768);
and UO_3176 (O_3176,N_44144,N_43236);
or UO_3177 (O_3177,N_49333,N_49861);
nor UO_3178 (O_3178,N_49191,N_40843);
xor UO_3179 (O_3179,N_40102,N_45118);
or UO_3180 (O_3180,N_41345,N_45465);
nand UO_3181 (O_3181,N_45771,N_49402);
and UO_3182 (O_3182,N_43193,N_46525);
and UO_3183 (O_3183,N_40168,N_41947);
xor UO_3184 (O_3184,N_48221,N_40401);
nand UO_3185 (O_3185,N_48127,N_45256);
nand UO_3186 (O_3186,N_45758,N_43035);
nand UO_3187 (O_3187,N_47388,N_42809);
and UO_3188 (O_3188,N_41955,N_46231);
nor UO_3189 (O_3189,N_44570,N_46670);
nor UO_3190 (O_3190,N_43840,N_44264);
nand UO_3191 (O_3191,N_42460,N_45213);
or UO_3192 (O_3192,N_42501,N_47116);
nand UO_3193 (O_3193,N_40967,N_40601);
nor UO_3194 (O_3194,N_45704,N_40976);
xnor UO_3195 (O_3195,N_43925,N_45194);
nor UO_3196 (O_3196,N_49584,N_40214);
xor UO_3197 (O_3197,N_40611,N_46992);
or UO_3198 (O_3198,N_42179,N_45145);
xnor UO_3199 (O_3199,N_49908,N_49936);
or UO_3200 (O_3200,N_47230,N_45883);
xor UO_3201 (O_3201,N_45641,N_45292);
nor UO_3202 (O_3202,N_45992,N_41160);
nand UO_3203 (O_3203,N_46725,N_46334);
nand UO_3204 (O_3204,N_42190,N_45598);
xor UO_3205 (O_3205,N_43417,N_43288);
or UO_3206 (O_3206,N_44913,N_47361);
and UO_3207 (O_3207,N_45722,N_43344);
or UO_3208 (O_3208,N_47744,N_48901);
nand UO_3209 (O_3209,N_44031,N_46456);
nor UO_3210 (O_3210,N_42051,N_47560);
or UO_3211 (O_3211,N_49597,N_43348);
nor UO_3212 (O_3212,N_45503,N_47630);
nor UO_3213 (O_3213,N_44921,N_40139);
nor UO_3214 (O_3214,N_42259,N_45715);
and UO_3215 (O_3215,N_43621,N_41608);
nor UO_3216 (O_3216,N_42717,N_43953);
xnor UO_3217 (O_3217,N_48158,N_42079);
or UO_3218 (O_3218,N_46703,N_48639);
or UO_3219 (O_3219,N_49660,N_40055);
nor UO_3220 (O_3220,N_47911,N_43072);
nor UO_3221 (O_3221,N_43955,N_42027);
xnor UO_3222 (O_3222,N_45260,N_48930);
xnor UO_3223 (O_3223,N_41889,N_46858);
nor UO_3224 (O_3224,N_40445,N_40556);
nand UO_3225 (O_3225,N_40323,N_42616);
xnor UO_3226 (O_3226,N_46136,N_47512);
and UO_3227 (O_3227,N_40199,N_42596);
and UO_3228 (O_3228,N_45400,N_46055);
and UO_3229 (O_3229,N_47894,N_43405);
xnor UO_3230 (O_3230,N_49017,N_48258);
and UO_3231 (O_3231,N_48805,N_45887);
xnor UO_3232 (O_3232,N_45532,N_43008);
nor UO_3233 (O_3233,N_40108,N_47881);
nand UO_3234 (O_3234,N_48023,N_44192);
nor UO_3235 (O_3235,N_44423,N_40248);
nand UO_3236 (O_3236,N_41815,N_48759);
or UO_3237 (O_3237,N_47074,N_48572);
nand UO_3238 (O_3238,N_49531,N_47293);
xor UO_3239 (O_3239,N_40112,N_41242);
and UO_3240 (O_3240,N_45399,N_40064);
nor UO_3241 (O_3241,N_41855,N_49520);
and UO_3242 (O_3242,N_44016,N_47187);
nor UO_3243 (O_3243,N_48321,N_42568);
xor UO_3244 (O_3244,N_43256,N_42938);
and UO_3245 (O_3245,N_48819,N_42758);
nand UO_3246 (O_3246,N_40639,N_44909);
nor UO_3247 (O_3247,N_47415,N_44355);
xnor UO_3248 (O_3248,N_43042,N_43210);
xnor UO_3249 (O_3249,N_46712,N_48370);
xor UO_3250 (O_3250,N_42507,N_45648);
xnor UO_3251 (O_3251,N_49463,N_42674);
or UO_3252 (O_3252,N_40472,N_43303);
xor UO_3253 (O_3253,N_46451,N_42470);
nand UO_3254 (O_3254,N_43439,N_44847);
and UO_3255 (O_3255,N_40252,N_45658);
nand UO_3256 (O_3256,N_42355,N_45781);
and UO_3257 (O_3257,N_42952,N_49683);
xor UO_3258 (O_3258,N_46165,N_44196);
nor UO_3259 (O_3259,N_48846,N_41643);
xnor UO_3260 (O_3260,N_48706,N_43004);
nor UO_3261 (O_3261,N_48684,N_47826);
nor UO_3262 (O_3262,N_46994,N_44360);
and UO_3263 (O_3263,N_49979,N_44590);
xor UO_3264 (O_3264,N_48187,N_43638);
xor UO_3265 (O_3265,N_41360,N_49674);
xnor UO_3266 (O_3266,N_44971,N_41762);
xor UO_3267 (O_3267,N_42753,N_43171);
xor UO_3268 (O_3268,N_49266,N_46312);
nand UO_3269 (O_3269,N_42189,N_45116);
nand UO_3270 (O_3270,N_43730,N_41772);
xor UO_3271 (O_3271,N_44123,N_47690);
and UO_3272 (O_3272,N_44267,N_44456);
nor UO_3273 (O_3273,N_48799,N_44176);
and UO_3274 (O_3274,N_47963,N_43036);
and UO_3275 (O_3275,N_46505,N_40378);
nand UO_3276 (O_3276,N_49376,N_47982);
nor UO_3277 (O_3277,N_43138,N_47362);
nand UO_3278 (O_3278,N_44487,N_46420);
nor UO_3279 (O_3279,N_42546,N_43395);
nand UO_3280 (O_3280,N_48895,N_49093);
and UO_3281 (O_3281,N_43048,N_42646);
or UO_3282 (O_3282,N_46663,N_47197);
xnor UO_3283 (O_3283,N_42946,N_41656);
nand UO_3284 (O_3284,N_44494,N_47823);
nor UO_3285 (O_3285,N_49564,N_47848);
or UO_3286 (O_3286,N_41311,N_40273);
and UO_3287 (O_3287,N_48242,N_42545);
and UO_3288 (O_3288,N_47799,N_44773);
and UO_3289 (O_3289,N_44526,N_40867);
nor UO_3290 (O_3290,N_49692,N_43855);
or UO_3291 (O_3291,N_48881,N_47506);
and UO_3292 (O_3292,N_44429,N_45410);
nand UO_3293 (O_3293,N_47285,N_43272);
and UO_3294 (O_3294,N_49906,N_42985);
nor UO_3295 (O_3295,N_43433,N_42795);
or UO_3296 (O_3296,N_47994,N_48171);
xnor UO_3297 (O_3297,N_49414,N_45188);
nor UO_3298 (O_3298,N_45237,N_42423);
nor UO_3299 (O_3299,N_44939,N_41416);
or UO_3300 (O_3300,N_43132,N_47801);
or UO_3301 (O_3301,N_47250,N_46473);
nand UO_3302 (O_3302,N_43968,N_46167);
nor UO_3303 (O_3303,N_49558,N_47808);
xor UO_3304 (O_3304,N_45203,N_48966);
nand UO_3305 (O_3305,N_48923,N_40716);
xnor UO_3306 (O_3306,N_41431,N_42436);
xnor UO_3307 (O_3307,N_48756,N_48455);
or UO_3308 (O_3308,N_44047,N_47649);
nand UO_3309 (O_3309,N_46344,N_42867);
xnor UO_3310 (O_3310,N_47391,N_46588);
or UO_3311 (O_3311,N_45902,N_42094);
or UO_3312 (O_3312,N_44198,N_49052);
nor UO_3313 (O_3313,N_44316,N_43515);
nor UO_3314 (O_3314,N_46633,N_40711);
xnor UO_3315 (O_3315,N_47249,N_47661);
xor UO_3316 (O_3316,N_43358,N_47396);
and UO_3317 (O_3317,N_49118,N_43687);
xor UO_3318 (O_3318,N_40060,N_49885);
xnor UO_3319 (O_3319,N_41065,N_44776);
nand UO_3320 (O_3320,N_49472,N_48524);
nor UO_3321 (O_3321,N_48982,N_45242);
or UO_3322 (O_3322,N_44249,N_44613);
and UO_3323 (O_3323,N_46331,N_41632);
nor UO_3324 (O_3324,N_45749,N_45083);
or UO_3325 (O_3325,N_41463,N_42402);
nor UO_3326 (O_3326,N_41008,N_41687);
or UO_3327 (O_3327,N_47400,N_44552);
xor UO_3328 (O_3328,N_43690,N_42604);
or UO_3329 (O_3329,N_47913,N_49526);
nand UO_3330 (O_3330,N_43357,N_43525);
nor UO_3331 (O_3331,N_49598,N_48156);
nor UO_3332 (O_3332,N_48066,N_46780);
or UO_3333 (O_3333,N_42058,N_47210);
nand UO_3334 (O_3334,N_43124,N_40814);
and UO_3335 (O_3335,N_41040,N_47160);
nor UO_3336 (O_3336,N_45270,N_43134);
or UO_3337 (O_3337,N_45789,N_49165);
or UO_3338 (O_3338,N_42194,N_41309);
nand UO_3339 (O_3339,N_44071,N_47454);
nand UO_3340 (O_3340,N_48223,N_47066);
xnor UO_3341 (O_3341,N_48356,N_47315);
xnor UO_3342 (O_3342,N_42312,N_44232);
or UO_3343 (O_3343,N_41375,N_41092);
xnor UO_3344 (O_3344,N_46278,N_44703);
nand UO_3345 (O_3345,N_42757,N_41645);
nand UO_3346 (O_3346,N_40035,N_47955);
xor UO_3347 (O_3347,N_40690,N_40128);
xnor UO_3348 (O_3348,N_49145,N_46583);
xor UO_3349 (O_3349,N_46316,N_43367);
nor UO_3350 (O_3350,N_47000,N_49498);
xor UO_3351 (O_3351,N_48179,N_42903);
nand UO_3352 (O_3352,N_46461,N_45531);
nand UO_3353 (O_3353,N_47740,N_45821);
nor UO_3354 (O_3354,N_44607,N_44557);
and UO_3355 (O_3355,N_40306,N_44558);
nor UO_3356 (O_3356,N_40598,N_45153);
or UO_3357 (O_3357,N_46029,N_40581);
xnor UO_3358 (O_3358,N_44491,N_40681);
xnor UO_3359 (O_3359,N_49998,N_40216);
or UO_3360 (O_3360,N_45028,N_47992);
nand UO_3361 (O_3361,N_47812,N_47574);
and UO_3362 (O_3362,N_42414,N_46421);
or UO_3363 (O_3363,N_46785,N_48963);
and UO_3364 (O_3364,N_49048,N_46921);
xnor UO_3365 (O_3365,N_48462,N_45606);
or UO_3366 (O_3366,N_42699,N_44896);
nand UO_3367 (O_3367,N_40704,N_43114);
or UO_3368 (O_3368,N_41811,N_48097);
nor UO_3369 (O_3369,N_43695,N_47254);
xor UO_3370 (O_3370,N_42388,N_41103);
nor UO_3371 (O_3371,N_43809,N_46159);
xor UO_3372 (O_3372,N_49763,N_46788);
or UO_3373 (O_3373,N_47350,N_45161);
nand UO_3374 (O_3374,N_47176,N_46512);
nor UO_3375 (O_3375,N_49524,N_41087);
xor UO_3376 (O_3376,N_47217,N_40369);
nor UO_3377 (O_3377,N_45411,N_42969);
xnor UO_3378 (O_3378,N_47359,N_49291);
nand UO_3379 (O_3379,N_45009,N_42019);
or UO_3380 (O_3380,N_48299,N_41641);
nor UO_3381 (O_3381,N_46428,N_42635);
nand UO_3382 (O_3382,N_43797,N_43616);
nand UO_3383 (O_3383,N_49393,N_46542);
and UO_3384 (O_3384,N_44023,N_43755);
or UO_3385 (O_3385,N_49295,N_44865);
nand UO_3386 (O_3386,N_41869,N_40338);
nor UO_3387 (O_3387,N_44546,N_44623);
or UO_3388 (O_3388,N_44261,N_47080);
nand UO_3389 (O_3389,N_43197,N_48076);
or UO_3390 (O_3390,N_46765,N_44977);
nand UO_3391 (O_3391,N_49945,N_41701);
and UO_3392 (O_3392,N_41327,N_42685);
xnor UO_3393 (O_3393,N_42817,N_45449);
xnor UO_3394 (O_3394,N_48755,N_43164);
or UO_3395 (O_3395,N_41173,N_46773);
nand UO_3396 (O_3396,N_40403,N_46153);
nor UO_3397 (O_3397,N_43612,N_49652);
or UO_3398 (O_3398,N_45840,N_42771);
nand UO_3399 (O_3399,N_42633,N_46550);
nand UO_3400 (O_3400,N_42228,N_41834);
or UO_3401 (O_3401,N_48192,N_48889);
and UO_3402 (O_3402,N_44611,N_47059);
nor UO_3403 (O_3403,N_43566,N_41975);
and UO_3404 (O_3404,N_45884,N_41243);
nor UO_3405 (O_3405,N_45799,N_41260);
nand UO_3406 (O_3406,N_44630,N_49486);
or UO_3407 (O_3407,N_43220,N_42631);
xnor UO_3408 (O_3408,N_42698,N_47524);
nand UO_3409 (O_3409,N_47908,N_41859);
and UO_3410 (O_3410,N_49345,N_44356);
nor UO_3411 (O_3411,N_49829,N_41605);
or UO_3412 (O_3412,N_42958,N_45889);
and UO_3413 (O_3413,N_42159,N_44253);
nand UO_3414 (O_3414,N_49832,N_40669);
and UO_3415 (O_3415,N_47475,N_49306);
nor UO_3416 (O_3416,N_40873,N_43016);
nor UO_3417 (O_3417,N_41024,N_49115);
nor UO_3418 (O_3418,N_48275,N_42347);
and UO_3419 (O_3419,N_42527,N_45663);
nand UO_3420 (O_3420,N_49482,N_45644);
nand UO_3421 (O_3421,N_49338,N_46333);
nor UO_3422 (O_3422,N_41906,N_48424);
and UO_3423 (O_3423,N_47651,N_42070);
and UO_3424 (O_3424,N_48972,N_43869);
nor UO_3425 (O_3425,N_41246,N_44790);
nor UO_3426 (O_3426,N_41153,N_44069);
nand UO_3427 (O_3427,N_48397,N_48919);
or UO_3428 (O_3428,N_49124,N_40182);
xnor UO_3429 (O_3429,N_43467,N_49151);
nor UO_3430 (O_3430,N_45384,N_47824);
or UO_3431 (O_3431,N_41223,N_41411);
xor UO_3432 (O_3432,N_45671,N_49933);
nor UO_3433 (O_3433,N_40917,N_46479);
or UO_3434 (O_3434,N_43862,N_43136);
nor UO_3435 (O_3435,N_48329,N_44241);
xor UO_3436 (O_3436,N_41854,N_46622);
and UO_3437 (O_3437,N_47336,N_41617);
xnor UO_3438 (O_3438,N_40666,N_46997);
and UO_3439 (O_3439,N_47099,N_45302);
nand UO_3440 (O_3440,N_40226,N_46373);
nor UO_3441 (O_3441,N_42238,N_41102);
and UO_3442 (O_3442,N_42621,N_46814);
or UO_3443 (O_3443,N_40973,N_40434);
and UO_3444 (O_3444,N_45422,N_45602);
or UO_3445 (O_3445,N_44941,N_49123);
or UO_3446 (O_3446,N_48867,N_43187);
nor UO_3447 (O_3447,N_48457,N_46274);
and UO_3448 (O_3448,N_44833,N_42642);
and UO_3449 (O_3449,N_44204,N_47167);
xnor UO_3450 (O_3450,N_47468,N_40521);
and UO_3451 (O_3451,N_47368,N_41927);
nand UO_3452 (O_3452,N_49174,N_44004);
nand UO_3453 (O_3453,N_43618,N_48884);
nand UO_3454 (O_3454,N_40994,N_45054);
nand UO_3455 (O_3455,N_49893,N_44710);
and UO_3456 (O_3456,N_49236,N_45790);
and UO_3457 (O_3457,N_44937,N_48026);
nor UO_3458 (O_3458,N_46390,N_47776);
nor UO_3459 (O_3459,N_45572,N_41290);
nor UO_3460 (O_3460,N_40176,N_45397);
and UO_3461 (O_3461,N_40683,N_46848);
xnor UO_3462 (O_3462,N_48232,N_44201);
xor UO_3463 (O_3463,N_45862,N_44765);
nor UO_3464 (O_3464,N_44012,N_42575);
nor UO_3465 (O_3465,N_47448,N_41354);
or UO_3466 (O_3466,N_48012,N_41630);
nand UO_3467 (O_3467,N_41452,N_42723);
xor UO_3468 (O_3468,N_49462,N_43047);
nand UO_3469 (O_3469,N_40979,N_44706);
nand UO_3470 (O_3470,N_48985,N_41844);
and UO_3471 (O_3471,N_44889,N_46888);
nand UO_3472 (O_3472,N_45616,N_40160);
nor UO_3473 (O_3473,N_41770,N_46802);
or UO_3474 (O_3474,N_49975,N_43015);
nand UO_3475 (O_3475,N_45988,N_45179);
or UO_3476 (O_3476,N_47777,N_44124);
nor UO_3477 (O_3477,N_47137,N_42907);
and UO_3478 (O_3478,N_44692,N_44814);
xnor UO_3479 (O_3479,N_47168,N_40901);
or UO_3480 (O_3480,N_45030,N_48592);
xor UO_3481 (O_3481,N_45892,N_43743);
nor UO_3482 (O_3482,N_43184,N_48335);
xor UO_3483 (O_3483,N_42099,N_42705);
nor UO_3484 (O_3484,N_47807,N_43806);
nor UO_3485 (O_3485,N_43997,N_45441);
nor UO_3486 (O_3486,N_41527,N_45229);
nand UO_3487 (O_3487,N_48510,N_48731);
and UO_3488 (O_3488,N_47863,N_46609);
nor UO_3489 (O_3489,N_48288,N_41916);
or UO_3490 (O_3490,N_49806,N_44403);
xor UO_3491 (O_3491,N_47224,N_45898);
or UO_3492 (O_3492,N_40080,N_46754);
and UO_3493 (O_3493,N_42132,N_46893);
and UO_3494 (O_3494,N_49383,N_45726);
nand UO_3495 (O_3495,N_42779,N_44214);
nor UO_3496 (O_3496,N_44934,N_48041);
nor UO_3497 (O_3497,N_48120,N_41171);
and UO_3498 (O_3498,N_44421,N_40983);
nor UO_3499 (O_3499,N_41382,N_46151);
and UO_3500 (O_3500,N_47633,N_44573);
nor UO_3501 (O_3501,N_41207,N_48600);
xor UO_3502 (O_3502,N_45882,N_49664);
and UO_3503 (O_3503,N_44490,N_43372);
and UO_3504 (O_3504,N_42254,N_45186);
or UO_3505 (O_3505,N_49640,N_44856);
or UO_3506 (O_3506,N_43160,N_44385);
or UO_3507 (O_3507,N_43607,N_49761);
and UO_3508 (O_3508,N_44027,N_44236);
nand UO_3509 (O_3509,N_44556,N_46024);
xor UO_3510 (O_3510,N_45004,N_40350);
xnor UO_3511 (O_3511,N_43936,N_49611);
and UO_3512 (O_3512,N_41546,N_46049);
and UO_3513 (O_3513,N_43802,N_42953);
or UO_3514 (O_3514,N_49624,N_48801);
xnor UO_3515 (O_3515,N_40087,N_49461);
xnor UO_3516 (O_3516,N_40376,N_44103);
nor UO_3517 (O_3517,N_49954,N_48730);
or UO_3518 (O_3518,N_43063,N_46962);
nor UO_3519 (O_3519,N_49016,N_40584);
and UO_3520 (O_3520,N_45193,N_46970);
nor UO_3521 (O_3521,N_48769,N_41792);
xnor UO_3522 (O_3522,N_48384,N_46811);
and UO_3523 (O_3523,N_44227,N_44804);
and UO_3524 (O_3524,N_49513,N_44186);
xor UO_3525 (O_3525,N_43321,N_43787);
nor UO_3526 (O_3526,N_47679,N_44916);
nor UO_3527 (O_3527,N_44400,N_43861);
xor UO_3528 (O_3528,N_40892,N_48301);
xor UO_3529 (O_3529,N_49530,N_41879);
and UO_3530 (O_3530,N_49237,N_49909);
nand UO_3531 (O_3531,N_41363,N_41234);
nand UO_3532 (O_3532,N_45496,N_46172);
nor UO_3533 (O_3533,N_47345,N_42679);
nand UO_3534 (O_3534,N_45473,N_49874);
or UO_3535 (O_3535,N_41824,N_45140);
and UO_3536 (O_3536,N_41533,N_43528);
xnor UO_3537 (O_3537,N_44981,N_47653);
nor UO_3538 (O_3538,N_43575,N_49919);
or UO_3539 (O_3539,N_40505,N_44005);
or UO_3540 (O_3540,N_47282,N_40539);
and UO_3541 (O_3541,N_46251,N_43798);
nor UO_3542 (O_3542,N_45504,N_45800);
or UO_3543 (O_3543,N_41530,N_46377);
and UO_3544 (O_3544,N_45401,N_46348);
nand UO_3545 (O_3545,N_43530,N_45061);
xnor UO_3546 (O_3546,N_48330,N_49430);
xnor UO_3547 (O_3547,N_41672,N_49540);
and UO_3548 (O_3548,N_46859,N_47951);
nand UO_3549 (O_3549,N_44955,N_42489);
and UO_3550 (O_3550,N_44755,N_44285);
nand UO_3551 (O_3551,N_46640,N_47002);
and UO_3552 (O_3552,N_40938,N_46726);
and UO_3553 (O_3553,N_48601,N_46502);
and UO_3554 (O_3554,N_46771,N_46289);
nor UO_3555 (O_3555,N_46741,N_44157);
nor UO_3556 (O_3556,N_45019,N_40113);
xor UO_3557 (O_3557,N_45927,N_45710);
xor UO_3558 (O_3558,N_48331,N_49959);
nor UO_3559 (O_3559,N_49535,N_45198);
or UO_3560 (O_3560,N_49162,N_47580);
nand UO_3561 (O_3561,N_46961,N_48573);
or UO_3562 (O_3562,N_44806,N_40537);
and UO_3563 (O_3563,N_44882,N_42583);
or UO_3564 (O_3564,N_43030,N_48650);
nand UO_3565 (O_3565,N_42083,N_44381);
xor UO_3566 (O_3566,N_46576,N_49714);
or UO_3567 (O_3567,N_45955,N_43387);
and UO_3568 (O_3568,N_40046,N_41618);
and UO_3569 (O_3569,N_49227,N_44864);
nor UO_3570 (O_3570,N_45818,N_44672);
nand UO_3571 (O_3571,N_46637,N_43366);
nor UO_3572 (O_3572,N_44926,N_47223);
or UO_3573 (O_3573,N_45796,N_41257);
xnor UO_3574 (O_3574,N_47698,N_47107);
nor UO_3575 (O_3575,N_45778,N_46524);
or UO_3576 (O_3576,N_49708,N_40083);
nor UO_3577 (O_3577,N_42990,N_46217);
or UO_3578 (O_3578,N_44516,N_42906);
nor UO_3579 (O_3579,N_41015,N_45366);
and UO_3580 (O_3580,N_40244,N_42770);
nor UO_3581 (O_3581,N_43609,N_48723);
and UO_3582 (O_3582,N_44138,N_44868);
or UO_3583 (O_3583,N_45901,N_47898);
or UO_3584 (O_3584,N_45915,N_47159);
or UO_3585 (O_3585,N_45033,N_47091);
or UO_3586 (O_3586,N_47414,N_41582);
xnor UO_3587 (O_3587,N_44945,N_40842);
nand UO_3588 (O_3588,N_41180,N_44065);
nand UO_3589 (O_3589,N_41771,N_46682);
xnor UO_3590 (O_3590,N_43402,N_48211);
nor UO_3591 (O_3591,N_48742,N_49168);
and UO_3592 (O_3592,N_44351,N_47958);
and UO_3593 (O_3593,N_46290,N_47657);
and UO_3594 (O_3594,N_43066,N_41970);
nand UO_3595 (O_3595,N_46181,N_48628);
nand UO_3596 (O_3596,N_49186,N_44350);
nor UO_3597 (O_3597,N_48139,N_49416);
or UO_3598 (O_3598,N_42399,N_40509);
or UO_3599 (O_3599,N_40092,N_40322);
or UO_3600 (O_3600,N_43637,N_40231);
or UO_3601 (O_3601,N_48594,N_43636);
and UO_3602 (O_3602,N_47984,N_47979);
and UO_3603 (O_3603,N_43065,N_42579);
xnor UO_3604 (O_3604,N_40018,N_42169);
nor UO_3605 (O_3605,N_44115,N_41786);
nand UO_3606 (O_3606,N_42943,N_49778);
and UO_3607 (O_3607,N_45341,N_45333);
or UO_3608 (O_3608,N_46618,N_45226);
xor UO_3609 (O_3609,N_46903,N_42571);
nor UO_3610 (O_3610,N_40559,N_46719);
xnor UO_3611 (O_3611,N_46615,N_45756);
and UO_3612 (O_3612,N_49976,N_47603);
xor UO_3613 (O_3613,N_43680,N_44417);
or UO_3614 (O_3614,N_47871,N_40756);
xnor UO_3615 (O_3615,N_49841,N_48644);
nor UO_3616 (O_3616,N_42106,N_45312);
xnor UO_3617 (O_3617,N_40564,N_46529);
and UO_3618 (O_3618,N_47988,N_45870);
xnor UO_3619 (O_3619,N_43425,N_43729);
nand UO_3620 (O_3620,N_48570,N_40169);
nor UO_3621 (O_3621,N_44608,N_40965);
xnor UO_3622 (O_3622,N_46736,N_44422);
nand UO_3623 (O_3623,N_47659,N_46597);
xnor UO_3624 (O_3624,N_42135,N_44887);
or UO_3625 (O_3625,N_41509,N_48915);
or UO_3626 (O_3626,N_47622,N_45483);
and UO_3627 (O_3627,N_49941,N_44271);
or UO_3628 (O_3628,N_46089,N_46255);
nand UO_3629 (O_3629,N_47103,N_41373);
or UO_3630 (O_3630,N_42479,N_47472);
xnor UO_3631 (O_3631,N_47057,N_47455);
or UO_3632 (O_3632,N_42567,N_49720);
nor UO_3633 (O_3633,N_43762,N_47281);
xor UO_3634 (O_3634,N_44741,N_49262);
nand UO_3635 (O_3635,N_45330,N_43620);
or UO_3636 (O_3636,N_43649,N_42232);
or UO_3637 (O_3637,N_42791,N_44671);
nand UO_3638 (O_3638,N_41659,N_46652);
nand UO_3639 (O_3639,N_40955,N_49840);
xnor UO_3640 (O_3640,N_49607,N_40645);
xor UO_3641 (O_3641,N_42321,N_41458);
nand UO_3642 (O_3642,N_41003,N_42366);
nand UO_3643 (O_3643,N_47928,N_44550);
nor UO_3644 (O_3644,N_40297,N_45805);
and UO_3645 (O_3645,N_44712,N_46170);
nor UO_3646 (O_3646,N_48124,N_43224);
or UO_3647 (O_3647,N_44811,N_46045);
nor UO_3648 (O_3648,N_43629,N_49745);
or UO_3649 (O_3649,N_45977,N_43645);
or UO_3650 (O_3650,N_49277,N_42262);
and UO_3651 (O_3651,N_43449,N_44402);
and UO_3652 (O_3652,N_46347,N_49092);
nand UO_3653 (O_3653,N_46839,N_49307);
xor UO_3654 (O_3654,N_45999,N_43178);
xnor UO_3655 (O_3655,N_46932,N_40468);
nor UO_3656 (O_3656,N_49995,N_49873);
or UO_3657 (O_3657,N_47917,N_45309);
xor UO_3658 (O_3658,N_48005,N_41241);
nand UO_3659 (O_3659,N_42074,N_47652);
or UO_3660 (O_3660,N_45674,N_44162);
and UO_3661 (O_3661,N_48921,N_45482);
and UO_3662 (O_3662,N_40166,N_41780);
and UO_3663 (O_3663,N_46191,N_41520);
xor UO_3664 (O_3664,N_43623,N_41790);
nand UO_3665 (O_3665,N_45487,N_43639);
or UO_3666 (O_3666,N_43726,N_42397);
nor UO_3667 (O_3667,N_44674,N_41282);
nor UO_3668 (O_3668,N_41654,N_46285);
or UO_3669 (O_3669,N_41222,N_49556);
or UO_3670 (O_3670,N_47526,N_46739);
nand UO_3671 (O_3671,N_47758,N_40238);
nor UO_3672 (O_3672,N_40771,N_45919);
nor UO_3673 (O_3673,N_46416,N_46005);
xor UO_3674 (O_3674,N_43856,N_40783);
and UO_3675 (O_3675,N_43157,N_42467);
or UO_3676 (O_3676,N_49342,N_41953);
and UO_3677 (O_3677,N_48917,N_42369);
xnor UO_3678 (O_3678,N_48820,N_48927);
nor UO_3679 (O_3679,N_41380,N_44763);
nand UO_3680 (O_3680,N_48246,N_46658);
or UO_3681 (O_3681,N_48625,N_41726);
xor UO_3682 (O_3682,N_41333,N_40751);
nand UO_3683 (O_3683,N_47207,N_42566);
nor UO_3684 (O_3684,N_41355,N_42641);
or UO_3685 (O_3685,N_47877,N_45491);
nand UO_3686 (O_3686,N_44873,N_42354);
nor UO_3687 (O_3687,N_41230,N_43597);
nand UO_3688 (O_3688,N_46822,N_45154);
and UO_3689 (O_3689,N_42377,N_48190);
xnor UO_3690 (O_3690,N_41573,N_44346);
xnor UO_3691 (O_3691,N_40371,N_49554);
and UO_3692 (O_3692,N_41525,N_46854);
or UO_3693 (O_3693,N_42466,N_44625);
xor UO_3694 (O_3694,N_44818,N_46539);
xnor UO_3695 (O_3695,N_44525,N_48009);
xor UO_3696 (O_3696,N_46220,N_47381);
and UO_3697 (O_3697,N_41357,N_41690);
nand UO_3698 (O_3698,N_47181,N_47628);
xnor UO_3699 (O_3699,N_42297,N_46598);
nand UO_3700 (O_3700,N_49704,N_48448);
and UO_3701 (O_3701,N_47594,N_42116);
and UO_3702 (O_3702,N_47933,N_48240);
or UO_3703 (O_3703,N_40766,N_45890);
nand UO_3704 (O_3704,N_47363,N_42450);
nand UO_3705 (O_3705,N_48743,N_42313);
or UO_3706 (O_3706,N_48576,N_47127);
nor UO_3707 (O_3707,N_42293,N_46929);
and UO_3708 (O_3708,N_48646,N_45442);
or UO_3709 (O_3709,N_47480,N_40186);
xnor UO_3710 (O_3710,N_43614,N_45438);
or UO_3711 (O_3711,N_44464,N_49719);
nand UO_3712 (O_3712,N_40036,N_47544);
or UO_3713 (O_3713,N_42052,N_42965);
nor UO_3714 (O_3714,N_42675,N_44293);
and UO_3715 (O_3715,N_43465,N_40506);
or UO_3716 (O_3716,N_45859,N_43028);
xnor UO_3717 (O_3717,N_44108,N_48450);
nand UO_3718 (O_3718,N_43579,N_43414);
xor UO_3719 (O_3719,N_46687,N_40981);
xnor UO_3720 (O_3720,N_43174,N_41788);
xor UO_3721 (O_3721,N_49297,N_42406);
xor UO_3722 (O_3722,N_47248,N_46253);
nor UO_3723 (O_3723,N_45842,N_47162);
nor UO_3724 (O_3724,N_49589,N_46697);
nor UO_3725 (O_3725,N_45175,N_47004);
nand UO_3726 (O_3726,N_42272,N_45584);
and UO_3727 (O_3727,N_43206,N_45903);
xor UO_3728 (O_3728,N_44211,N_48973);
or UO_3729 (O_3729,N_49631,N_40695);
xor UO_3730 (O_3730,N_45335,N_40589);
nor UO_3731 (O_3731,N_49117,N_48492);
and UO_3732 (O_3732,N_43093,N_41625);
nand UO_3733 (O_3733,N_47446,N_49244);
and UO_3734 (O_3734,N_47208,N_44732);
xnor UO_3735 (O_3735,N_44639,N_40428);
nand UO_3736 (O_3736,N_42315,N_44544);
nand UO_3737 (O_3737,N_40920,N_43554);
nor UO_3738 (O_3738,N_41984,N_47523);
or UO_3739 (O_3739,N_40684,N_41078);
xor UO_3740 (O_3740,N_45696,N_48264);
xor UO_3741 (O_3741,N_42237,N_43835);
and UO_3742 (O_3742,N_49030,N_46412);
and UO_3743 (O_3743,N_41821,N_48426);
nand UO_3744 (O_3744,N_48229,N_47540);
xor UO_3745 (O_3745,N_47402,N_44034);
nor UO_3746 (O_3746,N_41090,N_41021);
and UO_3747 (O_3747,N_46714,N_41425);
xnor UO_3748 (O_3748,N_43904,N_47636);
and UO_3749 (O_3749,N_41485,N_40578);
nand UO_3750 (O_3750,N_40256,N_42363);
or UO_3751 (O_3751,N_43278,N_44900);
nor UO_3752 (O_3752,N_43388,N_46125);
xor UO_3753 (O_3753,N_41857,N_42890);
and UO_3754 (O_3754,N_43488,N_41428);
xnor UO_3755 (O_3755,N_47417,N_45528);
nand UO_3756 (O_3756,N_45750,N_46686);
xor UO_3757 (O_3757,N_48896,N_48879);
xor UO_3758 (O_3758,N_45074,N_43753);
nor UO_3759 (O_3759,N_40896,N_44666);
and UO_3760 (O_3760,N_42659,N_45067);
nor UO_3761 (O_3761,N_41322,N_45062);
and UO_3762 (O_3762,N_46474,N_40332);
nand UO_3763 (O_3763,N_43223,N_42156);
or UO_3764 (O_3764,N_42731,N_48204);
nand UO_3765 (O_3765,N_48667,N_43027);
nor UO_3766 (O_3766,N_42164,N_40065);
or UO_3767 (O_3767,N_42231,N_41381);
nand UO_3768 (O_3768,N_40765,N_46584);
and UO_3769 (O_3769,N_48941,N_47527);
nor UO_3770 (O_3770,N_48112,N_47814);
nand UO_3771 (O_3771,N_46184,N_48831);
xor UO_3772 (O_3772,N_46713,N_46614);
and UO_3773 (O_3773,N_45510,N_41468);
and UO_3774 (O_3774,N_42437,N_45012);
and UO_3775 (O_3775,N_47420,N_43745);
and UO_3776 (O_3776,N_44508,N_46135);
or UO_3777 (O_3777,N_42627,N_45760);
and UO_3778 (O_3778,N_42778,N_45794);
or UO_3779 (O_3779,N_46112,N_40738);
nor UO_3780 (O_3780,N_43983,N_44669);
nand UO_3781 (O_3781,N_43832,N_46248);
or UO_3782 (O_3782,N_40077,N_42422);
nor UO_3783 (O_3783,N_41106,N_47796);
or UO_3784 (O_3784,N_44829,N_45993);
and UO_3785 (O_3785,N_45279,N_42192);
or UO_3786 (O_3786,N_44129,N_43677);
nor UO_3787 (O_3787,N_44805,N_44496);
xnor UO_3788 (O_3788,N_47725,N_48466);
and UO_3789 (O_3789,N_45164,N_45517);
nor UO_3790 (O_3790,N_43182,N_49330);
nand UO_3791 (O_3791,N_41291,N_47140);
nand UO_3792 (O_3792,N_40444,N_46162);
xor UO_3793 (O_3793,N_46996,N_40872);
xor UO_3794 (O_3794,N_48446,N_48381);
xor UO_3795 (O_3795,N_49807,N_43242);
nor UO_3796 (O_3796,N_46431,N_46137);
and UO_3797 (O_3797,N_44365,N_42107);
nor UO_3798 (O_3798,N_41938,N_46693);
nor UO_3799 (O_3799,N_49471,N_42828);
nor UO_3800 (O_3800,N_46059,N_47037);
xor UO_3801 (O_3801,N_43945,N_49068);
or UO_3802 (O_3802,N_44155,N_45986);
nor UO_3803 (O_3803,N_47509,N_47405);
nor UO_3804 (O_3804,N_49675,N_41540);
nor UO_3805 (O_3805,N_48219,N_47481);
nand UO_3806 (O_3806,N_42687,N_45354);
xor UO_3807 (O_3807,N_41466,N_46969);
and UO_3808 (O_3808,N_47667,N_46458);
or UO_3809 (O_3809,N_49702,N_47377);
and UO_3810 (O_3810,N_40093,N_41335);
nor UO_3811 (O_3811,N_40777,N_49894);
and UO_3812 (O_3812,N_42087,N_49272);
nor UO_3813 (O_3813,N_46258,N_45011);
or UO_3814 (O_3814,N_43073,N_40658);
or UO_3815 (O_3815,N_43253,N_44113);
nor UO_3816 (O_3816,N_49348,N_40442);
or UO_3817 (O_3817,N_45378,N_46118);
nand UO_3818 (O_3818,N_49519,N_42734);
and UO_3819 (O_3819,N_47999,N_49319);
xnor UO_3820 (O_3820,N_43917,N_49609);
xor UO_3821 (O_3821,N_43772,N_43986);
nor UO_3822 (O_3822,N_42461,N_42026);
nand UO_3823 (O_3823,N_45071,N_42130);
or UO_3824 (O_3824,N_45327,N_40360);
xnor UO_3825 (O_3825,N_46174,N_40889);
and UO_3826 (O_3826,N_46530,N_42822);
nand UO_3827 (O_3827,N_44919,N_41010);
nor UO_3828 (O_3828,N_42415,N_48375);
nor UO_3829 (O_3829,N_49762,N_41293);
nor UO_3830 (O_3830,N_47541,N_49158);
or UO_3831 (O_3831,N_41971,N_42218);
nor UO_3832 (O_3832,N_45240,N_41550);
or UO_3833 (O_3833,N_42242,N_40070);
nand UO_3834 (O_3834,N_46157,N_47688);
nor UO_3835 (O_3835,N_47786,N_42808);
xnor UO_3836 (O_3836,N_41568,N_42374);
nor UO_3837 (O_3837,N_47668,N_47914);
xor UO_3838 (O_3838,N_41161,N_42839);
or UO_3839 (O_3839,N_47595,N_47969);
xor UO_3840 (O_3840,N_49859,N_46634);
nand UO_3841 (O_3841,N_43083,N_46521);
or UO_3842 (O_3842,N_44427,N_49748);
nor UO_3843 (O_3843,N_42278,N_45852);
xor UO_3844 (O_3844,N_48790,N_44454);
and UO_3845 (O_3845,N_47616,N_43920);
nor UO_3846 (O_3846,N_42158,N_45271);
xor UO_3847 (O_3847,N_49144,N_42223);
or UO_3848 (O_3848,N_46050,N_47437);
nand UO_3849 (O_3849,N_46321,N_49850);
or UO_3850 (O_3850,N_43995,N_49725);
and UO_3851 (O_3851,N_46805,N_48604);
nand UO_3852 (O_3852,N_45725,N_49970);
nor UO_3853 (O_3853,N_41325,N_42186);
nor UO_3854 (O_3854,N_49638,N_42090);
nand UO_3855 (O_3855,N_44995,N_41706);
nor UO_3856 (O_3856,N_49139,N_47060);
nand UO_3857 (O_3857,N_49743,N_46974);
nor UO_3858 (O_3858,N_48891,N_43251);
and UO_3859 (O_3859,N_41902,N_43864);
nand UO_3860 (O_3860,N_47039,N_49445);
nor UO_3861 (O_3861,N_48528,N_49459);
xor UO_3862 (O_3862,N_49956,N_43468);
nand UO_3863 (O_3863,N_49823,N_46235);
and UO_3864 (O_3864,N_49155,N_43854);
nand UO_3865 (O_3865,N_49904,N_47467);
and UO_3866 (O_3866,N_43140,N_45677);
or UO_3867 (O_3867,N_45207,N_47821);
nand UO_3868 (O_3868,N_42226,N_41176);
or UO_3869 (O_3869,N_43428,N_46254);
nor UO_3870 (O_3870,N_44336,N_47953);
nor UO_3871 (O_3871,N_43291,N_45112);
and UO_3872 (O_3872,N_43781,N_47684);
xnor UO_3873 (O_3873,N_40219,N_49484);
or UO_3874 (O_3874,N_49800,N_43330);
and UO_3875 (O_3875,N_46983,N_44690);
nand UO_3876 (O_3876,N_46226,N_43885);
nand UO_3877 (O_3877,N_45948,N_48826);
and UO_3878 (O_3878,N_48027,N_47299);
and UO_3879 (O_3879,N_49557,N_45070);
or UO_3880 (O_3880,N_48506,N_42028);
or UO_3881 (O_3881,N_43568,N_41998);
xor UO_3882 (O_3882,N_46178,N_45177);
and UO_3883 (O_3883,N_42381,N_48515);
and UO_3884 (O_3884,N_40816,N_49896);
or UO_3885 (O_3885,N_41595,N_44507);
and UO_3886 (O_3886,N_43279,N_46579);
nor UO_3887 (O_3887,N_40103,N_44673);
xor UO_3888 (O_3888,N_44389,N_47888);
xnor UO_3889 (O_3889,N_48945,N_49575);
or UO_3890 (O_3890,N_42630,N_49756);
or UO_3891 (O_3891,N_40745,N_40933);
nand UO_3892 (O_3892,N_46228,N_43420);
nor UO_3893 (O_3893,N_44097,N_47298);
nand UO_3894 (O_3894,N_49595,N_48117);
nor UO_3895 (O_3895,N_49577,N_41492);
xor UO_3896 (O_3896,N_45376,N_42068);
and UO_3897 (O_3897,N_40270,N_43144);
xor UO_3898 (O_3898,N_42410,N_49741);
xnor UO_3899 (O_3899,N_42781,N_43481);
xnor UO_3900 (O_3900,N_47535,N_44469);
and UO_3901 (O_3901,N_43121,N_48141);
nand UO_3902 (O_3902,N_43975,N_46977);
nor UO_3903 (O_3903,N_46607,N_44978);
and UO_3904 (O_3904,N_42962,N_41239);
xnor UO_3905 (O_3905,N_43727,N_45878);
or UO_3906 (O_3906,N_48208,N_45174);
nor UO_3907 (O_3907,N_49833,N_46835);
xor UO_3908 (O_3908,N_44213,N_49063);
or UO_3909 (O_3909,N_46831,N_43435);
nand UO_3910 (O_3910,N_45460,N_43179);
or UO_3911 (O_3911,N_40212,N_40877);
and UO_3912 (O_3912,N_45472,N_45850);
or UO_3913 (O_3913,N_42886,N_47036);
nor UO_3914 (O_3914,N_49476,N_40995);
and UO_3915 (O_3915,N_49680,N_46186);
nand UO_3916 (O_3916,N_45041,N_42948);
xnor UO_3917 (O_3917,N_45629,N_42411);
nand UO_3918 (O_3918,N_42587,N_44043);
nand UO_3919 (O_3919,N_49031,N_41342);
nand UO_3920 (O_3920,N_41330,N_49645);
or UO_3921 (O_3921,N_45812,N_49774);
nand UO_3922 (O_3922,N_48122,N_46246);
and UO_3923 (O_3923,N_46252,N_40962);
xor UO_3924 (O_3924,N_45960,N_43858);
and UO_3925 (O_3925,N_46548,N_47276);
xor UO_3926 (O_3926,N_48196,N_44382);
xor UO_3927 (O_3927,N_48546,N_45114);
or UO_3928 (O_3928,N_49122,N_40770);
xnor UO_3929 (O_3929,N_40450,N_49312);
and UO_3930 (O_3930,N_43298,N_47612);
and UO_3931 (O_3931,N_44520,N_48500);
nor UO_3932 (O_3932,N_46378,N_47741);
nand UO_3933 (O_3933,N_43336,N_46440);
and UO_3934 (O_3934,N_47770,N_47261);
nor UO_3935 (O_3935,N_48565,N_46751);
or UO_3936 (O_3936,N_41404,N_41836);
xnor UO_3937 (O_3937,N_43771,N_45712);
nor UO_3938 (O_3938,N_42333,N_43741);
xnor UO_3939 (O_3939,N_44908,N_40405);
and UO_3940 (O_3940,N_43504,N_42982);
and UO_3941 (O_3941,N_40124,N_41069);
xnor UO_3942 (O_3942,N_46965,N_49508);
nand UO_3943 (O_3943,N_42535,N_42688);
nand UO_3944 (O_3944,N_42951,N_45691);
nand UO_3945 (O_3945,N_47920,N_45506);
nor UO_3946 (O_3946,N_44379,N_44629);
or UO_3947 (O_3947,N_42712,N_40778);
and UO_3948 (O_3948,N_42683,N_46007);
nand UO_3949 (O_3949,N_48000,N_49411);
nor UO_3950 (O_3950,N_45673,N_47384);
nand UO_3951 (O_3951,N_46783,N_47392);
nor UO_3952 (O_3952,N_48095,N_47412);
or UO_3953 (O_3953,N_40470,N_41936);
nor UO_3954 (O_3954,N_49709,N_42244);
or UO_3955 (O_3955,N_49228,N_42264);
or UO_3956 (O_3956,N_41584,N_43603);
xnor UO_3957 (O_3957,N_46099,N_47202);
or UO_3958 (O_3958,N_41029,N_40222);
or UO_3959 (O_3959,N_48763,N_46433);
nor UO_3960 (O_3960,N_40464,N_47373);
nand UO_3961 (O_3961,N_43767,N_40741);
or UO_3962 (O_3962,N_45408,N_46466);
and UO_3963 (O_3963,N_48453,N_44821);
and UO_3964 (O_3964,N_47180,N_43545);
or UO_3965 (O_3965,N_42831,N_45024);
xnor UO_3966 (O_3966,N_41931,N_49183);
or UO_3967 (O_3967,N_47352,N_40631);
xor UO_3968 (O_3968,N_49270,N_45596);
nand UO_3969 (O_3969,N_46072,N_44643);
xor UO_3970 (O_3970,N_40520,N_43759);
xor UO_3971 (O_3971,N_46963,N_47495);
and UO_3972 (O_3972,N_48036,N_46753);
and UO_3973 (O_3973,N_46261,N_40594);
nand UO_3974 (O_3974,N_46304,N_41847);
or UO_3975 (O_3975,N_44386,N_44533);
xnor UO_3976 (O_3976,N_43737,N_42666);
nand UO_3977 (O_3977,N_42097,N_40224);
nor UO_3978 (O_3978,N_42213,N_48934);
or UO_3979 (O_3979,N_43520,N_40179);
and UO_3980 (O_3980,N_49891,N_46853);
and UO_3981 (O_3981,N_42837,N_41035);
nand UO_3982 (O_3982,N_48172,N_43980);
or UO_3983 (O_3983,N_44337,N_43052);
xor UO_3984 (O_3984,N_48778,N_46346);
xnor UO_3985 (O_3985,N_40109,N_42702);
xnor UO_3986 (O_3986,N_44954,N_44465);
and UO_3987 (O_3987,N_47072,N_49939);
nor UO_3988 (O_3988,N_49574,N_45199);
and UO_3989 (O_3989,N_43514,N_47463);
and UO_3990 (O_3990,N_44953,N_40181);
xor UO_3991 (O_3991,N_41148,N_45159);
and UO_3992 (O_3992,N_47607,N_46779);
nand UO_3993 (O_3993,N_40936,N_49184);
xor UO_3994 (O_3994,N_49794,N_49539);
nor UO_3995 (O_3995,N_40075,N_44235);
nor UO_3996 (O_3996,N_42440,N_45808);
nor UO_3997 (O_3997,N_42252,N_40138);
xnor UO_3998 (O_3998,N_43318,N_49729);
or UO_3999 (O_3999,N_48789,N_40599);
or UO_4000 (O_4000,N_43327,N_40009);
nand UO_4001 (O_4001,N_44151,N_48997);
nand UO_4002 (O_4002,N_40419,N_41758);
or UO_4003 (O_4003,N_45135,N_48283);
xnor UO_4004 (O_4004,N_45344,N_42963);
xor UO_4005 (O_4005,N_46326,N_49464);
nand UO_4006 (O_4006,N_45353,N_47023);
and UO_4007 (O_4007,N_46244,N_47306);
and UO_4008 (O_4008,N_43082,N_42160);
nor UO_4009 (O_4009,N_45478,N_44778);
xnor UO_4010 (O_4010,N_45050,N_41289);
or UO_4011 (O_4011,N_41753,N_42054);
and UO_4012 (O_4012,N_47179,N_47033);
xor UO_4013 (O_4013,N_40811,N_43012);
nand UO_4014 (O_4014,N_45876,N_42673);
nor UO_4015 (O_4015,N_40147,N_42556);
or UO_4016 (O_4016,N_49095,N_41610);
xnor UO_4017 (O_4017,N_44935,N_48016);
nand UO_4018 (O_4018,N_42634,N_43086);
and UO_4019 (O_4019,N_42274,N_46626);
nand UO_4020 (O_4020,N_43533,N_42799);
nor UO_4021 (O_4021,N_41574,N_44872);
nand UO_4022 (O_4022,N_42539,N_41700);
and UO_4023 (O_4023,N_45814,N_43180);
nor UO_4024 (O_4024,N_47329,N_44540);
xnor UO_4025 (O_4025,N_43003,N_49088);
xor UO_4026 (O_4026,N_42677,N_47334);
nor UO_4027 (O_4027,N_46504,N_48093);
xnor UO_4028 (O_4028,N_41444,N_49222);
and UO_4029 (O_4029,N_48822,N_44555);
and UO_4030 (O_4030,N_44918,N_40469);
nand UO_4031 (O_4031,N_46606,N_40855);
and UO_4032 (O_4032,N_45101,N_47974);
nor UO_4033 (O_4033,N_40435,N_47090);
nor UO_4034 (O_4034,N_45974,N_46660);
nand UO_4035 (O_4035,N_40706,N_47119);
nand UO_4036 (O_4036,N_40069,N_43250);
or UO_4037 (O_4037,N_40861,N_42843);
xor UO_4038 (O_4038,N_45827,N_49106);
xor UO_4039 (O_4039,N_40817,N_44399);
xnor UO_4040 (O_4040,N_49649,N_40411);
nor UO_4041 (O_4041,N_42612,N_47478);
nor UO_4042 (O_4042,N_46314,N_42142);
nand UO_4043 (O_4043,N_46701,N_40913);
nand UO_4044 (O_4044,N_42597,N_45351);
nor UO_4045 (O_4045,N_44304,N_44281);
xor UO_4046 (O_4046,N_47435,N_45879);
and UO_4047 (O_4047,N_46076,N_45533);
nand UO_4048 (O_4048,N_46269,N_47476);
nand UO_4049 (O_4049,N_46166,N_40604);
nor UO_4050 (O_4050,N_48578,N_41011);
or UO_4051 (O_4051,N_43732,N_41867);
nor UO_4052 (O_4052,N_48898,N_47165);
or UO_4053 (O_4053,N_43040,N_42775);
nor UO_4054 (O_4054,N_41146,N_47138);
and UO_4055 (O_4055,N_43799,N_49062);
or UO_4056 (O_4056,N_47047,N_44998);
and UO_4057 (O_4057,N_47973,N_48078);
and UO_4058 (O_4058,N_48017,N_45773);
nor UO_4059 (O_4059,N_45077,N_44178);
xor UO_4060 (O_4060,N_43950,N_47457);
xor UO_4061 (O_4061,N_41532,N_44297);
nand UO_4062 (O_4062,N_46478,N_48233);
nand UO_4063 (O_4063,N_49921,N_45462);
nor UO_4064 (O_4064,N_44064,N_46655);
xnor UO_4065 (O_4065,N_42008,N_49206);
or UO_4066 (O_4066,N_40265,N_41196);
nor UO_4067 (O_4067,N_43882,N_44135);
or UO_4068 (O_4068,N_41843,N_45485);
xnor UO_4069 (O_4069,N_44133,N_44269);
xor UO_4070 (O_4070,N_47771,N_43675);
nand UO_4071 (O_4071,N_44116,N_41559);
nor UO_4072 (O_4072,N_41337,N_41100);
or UO_4073 (O_4073,N_43786,N_48788);
nor UO_4074 (O_4074,N_45697,N_48247);
nand UO_4075 (O_4075,N_40487,N_49511);
nand UO_4076 (O_4076,N_47717,N_45733);
and UO_4077 (O_4077,N_48440,N_45117);
and UO_4078 (O_4078,N_45765,N_45920);
or UO_4079 (O_4079,N_45652,N_49592);
nor UO_4080 (O_4080,N_47910,N_47670);
and UO_4081 (O_4081,N_42654,N_49359);
and UO_4082 (O_4082,N_48094,N_47453);
or UO_4083 (O_4083,N_40779,N_44940);
xnor UO_4084 (O_4084,N_49090,N_44822);
or UO_4085 (O_4085,N_45076,N_48357);
xor UO_4086 (O_4086,N_40175,N_44938);
or UO_4087 (O_4087,N_47112,N_47938);
and UO_4088 (O_4088,N_49614,N_45021);
and UO_4089 (O_4089,N_47311,N_44722);
and UO_4090 (O_4090,N_47584,N_40086);
and UO_4091 (O_4091,N_41689,N_41356);
xnor UO_4092 (O_4092,N_48129,N_42598);
nand UO_4093 (O_4093,N_41077,N_48436);
or UO_4094 (O_4094,N_41392,N_40834);
or UO_4095 (O_4095,N_42336,N_45355);
or UO_4096 (O_4096,N_40164,N_45212);
nand UO_4097 (O_4097,N_46019,N_46966);
xnor UO_4098 (O_4098,N_40750,N_48886);
nor UO_4099 (O_4099,N_42682,N_41515);
or UO_4100 (O_4100,N_45225,N_48034);
and UO_4101 (O_4101,N_42518,N_49552);
nor UO_4102 (O_4102,N_44931,N_44132);
xnor UO_4103 (O_4103,N_49685,N_47519);
or UO_4104 (O_4104,N_46097,N_43133);
nand UO_4105 (O_4105,N_47186,N_42653);
nand UO_4106 (O_4106,N_45700,N_49548);
xor UO_4107 (O_4107,N_48484,N_40317);
or UO_4108 (O_4108,N_42176,N_46185);
or UO_4109 (O_4109,N_48132,N_41818);
nand UO_4110 (O_4110,N_40159,N_46791);
xnor UO_4111 (O_4111,N_41896,N_47214);
and UO_4112 (O_4112,N_47183,N_49036);
nor UO_4113 (O_4113,N_47516,N_45409);
nor UO_4114 (O_4114,N_40278,N_47970);
and UO_4115 (O_4115,N_41048,N_44893);
nor UO_4116 (O_4116,N_45938,N_47997);
xnor UO_4117 (O_4117,N_47240,N_45215);
nand UO_4118 (O_4118,N_41741,N_44536);
nand UO_4119 (O_4119,N_40999,N_45326);
or UO_4120 (O_4120,N_41285,N_42225);
nor UO_4121 (O_4121,N_49989,N_41344);
or UO_4122 (O_4122,N_43244,N_41516);
and UO_4123 (O_4123,N_45495,N_40090);
or UO_4124 (O_4124,N_44784,N_45426);
nor UO_4125 (O_4125,N_47301,N_45299);
and UO_4126 (O_4126,N_41607,N_41504);
nor UO_4127 (O_4127,N_46139,N_46806);
xnor UO_4128 (O_4128,N_45239,N_41104);
xnor UO_4129 (O_4129,N_48245,N_48244);
or UO_4130 (O_4130,N_47759,N_42375);
or UO_4131 (O_4131,N_42602,N_49446);
nand UO_4132 (O_4132,N_43625,N_43186);
or UO_4133 (O_4133,N_43459,N_41422);
or UO_4134 (O_4134,N_48849,N_48067);
xnor UO_4135 (O_4135,N_40532,N_43790);
or UO_4136 (O_4136,N_46942,N_42203);
and UO_4137 (O_4137,N_48618,N_44480);
and UO_4138 (O_4138,N_43674,N_46619);
or UO_4139 (O_4139,N_47411,N_46309);
and UO_4140 (O_4140,N_49497,N_44605);
nand UO_4141 (O_4141,N_48589,N_47134);
nand UO_4142 (O_4142,N_47852,N_43029);
and UO_4143 (O_4143,N_49757,N_43299);
or UO_4144 (O_4144,N_45493,N_40989);
nor UO_4145 (O_4145,N_40091,N_45106);
or UO_4146 (O_4146,N_42098,N_47682);
nand UO_4147 (O_4147,N_46238,N_47486);
nor UO_4148 (O_4148,N_43237,N_46535);
and UO_4149 (O_4149,N_41361,N_48488);
and UO_4150 (O_4150,N_48760,N_44834);
and UO_4151 (O_4151,N_40508,N_43874);
nor UO_4152 (O_4152,N_44161,N_44792);
xnor UO_4153 (O_4153,N_43258,N_41564);
nor UO_4154 (O_4154,N_48021,N_43297);
and UO_4155 (O_4155,N_41751,N_45142);
or UO_4156 (O_4156,N_41692,N_48109);
nand UO_4157 (O_4157,N_45431,N_42896);
and UO_4158 (O_4158,N_44366,N_46243);
or UO_4159 (O_4159,N_49751,N_45136);
nor UO_4160 (O_4160,N_46448,N_41991);
xor UO_4161 (O_4161,N_47196,N_48130);
or UO_4162 (O_4162,N_42215,N_47602);
or UO_4163 (O_4163,N_49686,N_47916);
or UO_4164 (O_4164,N_42166,N_42573);
nor UO_4165 (O_4165,N_40020,N_41122);
nor UO_4166 (O_4166,N_47166,N_43189);
or UO_4167 (O_4167,N_44635,N_47837);
or UO_4168 (O_4168,N_45985,N_46053);
xor UO_4169 (O_4169,N_41292,N_42617);
or UO_4170 (O_4170,N_45243,N_42299);
nor UO_4171 (O_4171,N_47256,N_49902);
or UO_4172 (O_4172,N_45822,N_49780);
nor UO_4173 (O_4173,N_49009,N_49232);
nand UO_4174 (O_4174,N_45369,N_47118);
or UO_4175 (O_4175,N_48656,N_47133);
nor UO_4176 (O_4176,N_42523,N_41170);
and UO_4177 (O_4177,N_45655,N_47308);
nand UO_4178 (O_4178,N_42454,N_47418);
nand UO_4179 (O_4179,N_44448,N_42080);
nor UO_4180 (O_4180,N_43129,N_45881);
nor UO_4181 (O_4181,N_47404,N_41093);
and UO_4182 (O_4182,N_47687,N_45016);
nand UO_4183 (O_4183,N_43877,N_43532);
nor UO_4184 (O_4184,N_45297,N_48153);
and UO_4185 (O_4185,N_47906,N_46943);
or UO_4186 (O_4186,N_41531,N_46665);
nand UO_4187 (O_4187,N_41864,N_47922);
nand UO_4188 (O_4188,N_45924,N_49899);
xnor UO_4189 (O_4189,N_49152,N_46803);
and UO_4190 (O_4190,N_49821,N_48870);
or UO_4191 (O_4191,N_49964,N_47763);
and UO_4192 (O_4192,N_45258,N_41407);
nand UO_4193 (O_4193,N_49900,N_40819);
nand UO_4194 (O_4194,N_44378,N_41033);
nor UO_4195 (O_4195,N_49969,N_42210);
and UO_4196 (O_4196,N_46520,N_42956);
xnor UO_4197 (O_4197,N_41571,N_42754);
nand UO_4198 (O_4198,N_42994,N_47936);
or UO_4199 (O_4199,N_44561,N_42562);
xnor UO_4200 (O_4200,N_48403,N_47989);
xor UO_4201 (O_4201,N_43988,N_43408);
and UO_4202 (O_4202,N_41876,N_45759);
nand UO_4203 (O_4203,N_49733,N_47322);
and UO_4204 (O_4204,N_49799,N_45965);
nand UO_4205 (O_4205,N_49884,N_44164);
nand UO_4206 (O_4206,N_43257,N_45130);
or UO_4207 (O_4207,N_49143,N_48520);
and UO_4208 (O_4208,N_41135,N_44952);
nand UO_4209 (O_4209,N_49457,N_49560);
or UO_4210 (O_4210,N_42625,N_43850);
nor UO_4211 (O_4211,N_48571,N_48783);
nor UO_4212 (O_4212,N_45740,N_49929);
nor UO_4213 (O_4213,N_42920,N_42664);
nor UO_4214 (O_4214,N_44486,N_40659);
and UO_4215 (O_4215,N_48772,N_41653);
nand UO_4216 (O_4216,N_48345,N_48549);
nor UO_4217 (O_4217,N_49157,N_44433);
xnor UO_4218 (O_4218,N_44345,N_43032);
or UO_4219 (O_4219,N_44320,N_46366);
nor UO_4220 (O_4220,N_42163,N_41274);
nand UO_4221 (O_4221,N_45621,N_45311);
and UO_4222 (O_4222,N_42314,N_44869);
or UO_4223 (O_4223,N_40057,N_41926);
and UO_4224 (O_4224,N_41001,N_43887);
nor UO_4225 (O_4225,N_49922,N_42306);
xor UO_4226 (O_4226,N_41149,N_44988);
nand UO_4227 (O_4227,N_45936,N_49081);
and UO_4228 (O_4228,N_42266,N_43611);
nor UO_4229 (O_4229,N_48121,N_45038);
or UO_4230 (O_4230,N_47677,N_48872);
xnor UO_4231 (O_4231,N_48608,N_42859);
nor UO_4232 (O_4232,N_40331,N_40269);
xor UO_4233 (O_4233,N_44542,N_48750);
and UO_4234 (O_4234,N_41665,N_46934);
xor UO_4235 (O_4235,N_41400,N_42117);
nand UO_4236 (O_4236,N_46425,N_41414);
and UO_4237 (O_4237,N_46092,N_49042);
or UO_4238 (O_4238,N_49194,N_40326);
xor UO_4239 (O_4239,N_44554,N_44089);
xor UO_4240 (O_4240,N_46330,N_43085);
and UO_4241 (O_4241,N_44840,N_40325);
nand UO_4242 (O_4242,N_46571,N_49171);
or UO_4243 (O_4243,N_40296,N_44451);
xnor UO_4244 (O_4244,N_40725,N_46236);
or UO_4245 (O_4245,N_40418,N_40358);
nor UO_4246 (O_4246,N_47706,N_46991);
and UO_4247 (O_4247,N_45553,N_41570);
xor UO_4248 (O_4248,N_40441,N_46590);
nor UO_4249 (O_4249,N_42668,N_40523);
nand UO_4250 (O_4250,N_43217,N_46411);
or UO_4251 (O_4251,N_43423,N_47606);
or UO_4252 (O_4252,N_43265,N_49947);
or UO_4253 (O_4253,N_48907,N_40858);
xor UO_4254 (O_4254,N_46497,N_45035);
nor UO_4255 (O_4255,N_47452,N_49474);
nor UO_4256 (O_4256,N_48918,N_41036);
xor UO_4257 (O_4257,N_40577,N_43095);
nor UO_4258 (O_4258,N_49341,N_44601);
xnor UO_4259 (O_4259,N_49701,N_44370);
nand UO_4260 (O_4260,N_47889,N_46580);
nor UO_4261 (O_4261,N_45731,N_46924);
nor UO_4262 (O_4262,N_46509,N_44511);
and UO_4263 (O_4263,N_47552,N_45841);
xnor UO_4264 (O_4264,N_41487,N_44256);
and UO_4265 (O_4265,N_42220,N_43717);
nor UO_4266 (O_4266,N_46361,N_47182);
nor UO_4267 (O_4267,N_46947,N_40459);
nor UO_4268 (O_4268,N_47543,N_49635);
nor UO_4269 (O_4269,N_48888,N_43391);
and UO_4270 (O_4270,N_40809,N_49938);
or UO_4271 (O_4271,N_49681,N_43308);
xnor UO_4272 (O_4272,N_43235,N_41032);
or UO_4273 (O_4273,N_44655,N_48307);
nand UO_4274 (O_4274,N_49051,N_49176);
nor UO_4275 (O_4275,N_45415,N_47494);
nor UO_4276 (O_4276,N_41979,N_40177);
nand UO_4277 (O_4277,N_43350,N_43572);
and UO_4278 (O_4278,N_46188,N_41635);
nand UO_4279 (O_4279,N_47498,N_46100);
xnor UO_4280 (O_4280,N_42941,N_49623);
xnor UO_4281 (O_4281,N_41017,N_43289);
xor UO_4282 (O_4282,N_49993,N_49641);
and UO_4283 (O_4283,N_43131,N_47109);
or UO_4284 (O_4284,N_45963,N_42502);
nand UO_4285 (O_4285,N_49728,N_47038);
nor UO_4286 (O_4286,N_45073,N_47097);
or UO_4287 (O_4287,N_47125,N_49190);
and UO_4288 (O_4288,N_42088,N_49308);
nor UO_4289 (O_4289,N_40515,N_49897);
xor UO_4290 (O_4290,N_40221,N_45259);
xnor UO_4291 (O_4291,N_41059,N_47810);
or UO_4292 (O_4292,N_45872,N_45461);
xnor UO_4293 (O_4293,N_49992,N_41254);
nor UO_4294 (O_4294,N_47831,N_47542);
xor UO_4295 (O_4295,N_43580,N_48074);
and UO_4296 (O_4296,N_40452,N_46317);
and UO_4297 (O_4297,N_44990,N_40608);
or UO_4298 (O_4298,N_41655,N_48758);
nand UO_4299 (O_4299,N_40439,N_40954);
nor UO_4300 (O_4300,N_40343,N_43889);
and UO_4301 (O_4301,N_40137,N_41809);
xor UO_4302 (O_4302,N_42744,N_42665);
nand UO_4303 (O_4303,N_43143,N_48222);
nand UO_4304 (O_4304,N_44594,N_48137);
nand UO_4305 (O_4305,N_46026,N_46383);
nor UO_4306 (O_4306,N_40668,N_43905);
or UO_4307 (O_4307,N_47947,N_49136);
nor UO_4308 (O_4308,N_48149,N_45257);
nor UO_4309 (O_4309,N_46689,N_41209);
and UO_4310 (O_4310,N_45013,N_49621);
or UO_4311 (O_4311,N_46232,N_49567);
and UO_4312 (O_4312,N_42726,N_47921);
or UO_4313 (O_4313,N_41948,N_47556);
nand UO_4314 (O_4314,N_44827,N_44924);
nand UO_4315 (O_4315,N_43529,N_46987);
or UO_4316 (O_4316,N_49996,N_45459);
and UO_4317 (O_4317,N_40600,N_45681);
nand UO_4318 (O_4318,N_43295,N_48703);
nor UO_4319 (O_4319,N_40985,N_47130);
nor UO_4320 (O_4320,N_47672,N_45163);
and UO_4321 (O_4321,N_43440,N_48555);
nor UO_4322 (O_4322,N_49002,N_43379);
and UO_4323 (O_4323,N_47842,N_47829);
nand UO_4324 (O_4324,N_49849,N_49834);
nand UO_4325 (O_4325,N_47108,N_46990);
and UO_4326 (O_4326,N_41707,N_42370);
nand UO_4327 (O_4327,N_43851,N_44286);
and UO_4328 (O_4328,N_42570,N_47985);
xor UO_4329 (O_4329,N_47073,N_46772);
nor UO_4330 (O_4330,N_49706,N_46729);
or UO_4331 (O_4331,N_47105,N_43218);
nand UO_4332 (O_4332,N_46563,N_46830);
nor UO_4333 (O_4333,N_46068,N_43192);
or UO_4334 (O_4334,N_44518,N_48603);
and UO_4335 (O_4335,N_45896,N_41973);
or UO_4336 (O_4336,N_40635,N_46355);
xor UO_4337 (O_4337,N_47374,N_43982);
nor UO_4338 (O_4338,N_42508,N_41177);
nor UO_4339 (O_4339,N_44545,N_40904);
nor UO_4340 (O_4340,N_43510,N_42609);
or UO_4341 (O_4341,N_44948,N_40475);
nand UO_4342 (O_4342,N_40760,N_49496);
and UO_4343 (O_4343,N_43384,N_48835);
nand UO_4344 (O_4344,N_42004,N_46884);
nor UO_4345 (O_4345,N_46750,N_48282);
and UO_4346 (O_4346,N_44445,N_45208);
xor UO_4347 (O_4347,N_43921,N_44150);
xor UO_4348 (O_4348,N_45412,N_45403);
nand UO_4349 (O_4349,N_49159,N_46894);
nand UO_4350 (O_4350,N_42548,N_40302);
nor UO_4351 (O_4351,N_48702,N_49716);
or UO_4352 (O_4352,N_46493,N_44528);
nand UO_4353 (O_4353,N_47451,N_42119);
xnor UO_4354 (O_4354,N_49301,N_44598);
nand UO_4355 (O_4355,N_42141,N_47782);
or UO_4356 (O_4356,N_42524,N_42181);
nand UO_4357 (O_4357,N_48767,N_47410);
and UO_4358 (O_4358,N_46395,N_46887);
or UO_4359 (O_4359,N_40101,N_41803);
nand UO_4360 (O_4360,N_46265,N_45984);
or UO_4361 (O_4361,N_41839,N_44502);
xor UO_4362 (O_4362,N_42897,N_48948);
or UO_4363 (O_4363,N_47117,N_49615);
and UO_4364 (O_4364,N_47945,N_46490);
xnor UO_4365 (O_4365,N_45863,N_43100);
and UO_4366 (O_4366,N_44260,N_46575);
and UO_4367 (O_4367,N_49294,N_49752);
nand UO_4368 (O_4368,N_48303,N_47884);
nor UO_4369 (O_4369,N_44119,N_43383);
or UO_4370 (O_4370,N_41523,N_42448);
xnor UO_4371 (O_4371,N_48476,N_48782);
or UO_4372 (O_4372,N_43681,N_49019);
nor UO_4373 (O_4373,N_48539,N_42881);
or UO_4374 (O_4374,N_40943,N_48705);
and UO_4375 (O_4375,N_47053,N_40394);
xor UO_4376 (O_4376,N_44748,N_48456);
nand UO_4377 (O_4377,N_42303,N_46565);
nand UO_4378 (O_4378,N_41047,N_43999);
or UO_4379 (O_4379,N_48033,N_48640);
and UO_4380 (O_4380,N_48364,N_41745);
or UO_4381 (O_4381,N_42619,N_42563);
or UO_4382 (O_4382,N_44933,N_42367);
xor UO_4383 (O_4383,N_46173,N_46061);
or UO_4384 (O_4384,N_44795,N_42846);
and UO_4385 (O_4385,N_45588,N_42457);
and UO_4386 (O_4386,N_44730,N_46778);
or UO_4387 (O_4387,N_40474,N_46657);
and UO_4388 (O_4388,N_47389,N_49920);
nand UO_4389 (O_4389,N_44134,N_47477);
xor UO_4390 (O_4390,N_41775,N_46679);
and UO_4391 (O_4391,N_44603,N_49827);
or UO_4392 (O_4392,N_46662,N_43658);
nor UO_4393 (O_4393,N_41388,N_41091);
or UO_4394 (O_4394,N_49626,N_45755);
nor UO_4395 (O_4395,N_49848,N_41064);
nand UO_4396 (O_4396,N_48858,N_40799);
nand UO_4397 (O_4397,N_40653,N_46419);
nand UO_4398 (O_4398,N_42110,N_47096);
xor UO_4399 (O_4399,N_49981,N_43791);
and UO_4400 (O_4400,N_42341,N_40284);
and UO_4401 (O_4401,N_47338,N_48899);
or UO_4402 (O_4402,N_44270,N_44376);
xnor UO_4403 (O_4403,N_49916,N_44194);
nand UO_4404 (O_4404,N_43923,N_46764);
xnor UO_4405 (O_4405,N_41376,N_43876);
and UO_4406 (O_4406,N_45772,N_46608);
nor UO_4407 (O_4407,N_47874,N_49820);
xnor UO_4408 (O_4408,N_49196,N_45987);
nand UO_4409 (O_4409,N_40802,N_43659);
nor UO_4410 (O_4410,N_45820,N_49007);
nand UO_4411 (O_4411,N_46554,N_40316);
and UO_4412 (O_4412,N_48752,N_40285);
nor UO_4413 (O_4413,N_42766,N_49871);
or UO_4414 (O_4414,N_44246,N_42594);
nand UO_4415 (O_4415,N_41441,N_46737);
nand UO_4416 (O_4416,N_40013,N_47092);
nor UO_4417 (O_4417,N_44334,N_49047);
xor UO_4418 (O_4418,N_47421,N_48304);
nand UO_4419 (O_4419,N_46868,N_48508);
xnor UO_4420 (O_4420,N_41218,N_47474);
nor UO_4421 (O_4421,N_40907,N_41502);
and UO_4422 (O_4422,N_47619,N_46816);
xnor UO_4423 (O_4423,N_48340,N_44145);
or UO_4424 (O_4424,N_42905,N_41379);
nor UO_4425 (O_4425,N_41544,N_41389);
xnor UO_4426 (O_4426,N_46985,N_41674);
nand UO_4427 (O_4427,N_47245,N_46489);
xor UO_4428 (O_4428,N_40798,N_45590);
nor UO_4429 (O_4429,N_48002,N_48632);
xor UO_4430 (O_4430,N_42151,N_40958);
xnor UO_4431 (O_4431,N_42475,N_43126);
nor UO_4432 (O_4432,N_43080,N_46685);
nor UO_4433 (O_4433,N_45413,N_48683);
xnor UO_4434 (O_4434,N_42624,N_41145);
nand UO_4435 (O_4435,N_47016,N_48959);
nor UO_4436 (O_4436,N_49431,N_46310);
or UO_4437 (O_4437,N_47589,N_44609);
xor UO_4438 (O_4438,N_48173,N_41320);
or UO_4439 (O_4439,N_40657,N_49364);
and UO_4440 (O_4440,N_45439,N_40825);
nor UO_4441 (O_4441,N_46222,N_40932);
nor UO_4442 (O_4442,N_41999,N_40390);
or UO_4443 (O_4443,N_47228,N_42115);
nor UO_4444 (O_4444,N_45342,N_42085);
nor UO_4445 (O_4445,N_44282,N_42287);
and UO_4446 (O_4446,N_46674,N_47431);
xnor UO_4447 (O_4447,N_44121,N_42874);
xor UO_4448 (O_4448,N_43959,N_48374);
nand UO_4449 (O_4449,N_44539,N_46799);
nor UO_4450 (O_4450,N_43667,N_49610);
nor UO_4451 (O_4451,N_42165,N_41070);
nand UO_4452 (O_4452,N_48286,N_46784);
and UO_4453 (O_4453,N_46901,N_40079);
or UO_4454 (O_4454,N_48260,N_46680);
nor UO_4455 (O_4455,N_43867,N_41558);
or UO_4456 (O_4456,N_49790,N_49629);
nand UO_4457 (O_4457,N_42310,N_42255);
or UO_4458 (O_4458,N_49967,N_43194);
xor UO_4459 (O_4459,N_44780,N_49286);
and UO_4460 (O_4460,N_42062,N_41791);
nand UO_4461 (O_4461,N_41832,N_41852);
nor UO_4462 (O_4462,N_48395,N_46391);
or UO_4463 (O_4463,N_40033,N_46695);
nand UO_4464 (O_4464,N_49177,N_44620);
or UO_4465 (O_4465,N_42736,N_41566);
xnor UO_4466 (O_4466,N_42978,N_43320);
nor UO_4467 (O_4467,N_47991,N_44728);
or UO_4468 (O_4468,N_46809,N_49224);
xnor UO_4469 (O_4469,N_43195,N_40830);
nor UO_4470 (O_4470,N_43368,N_43474);
nor UO_4471 (O_4471,N_47709,N_48155);
nand UO_4472 (O_4472,N_45624,N_40174);
or UO_4473 (O_4473,N_45463,N_42645);
xnor UO_4474 (O_4474,N_47253,N_44808);
nand UO_4475 (O_4475,N_44056,N_41156);
xor UO_4476 (O_4476,N_48505,N_42326);
and UO_4477 (O_4477,N_40148,N_42592);
or UO_4478 (O_4478,N_43570,N_46632);
and UO_4479 (O_4479,N_46096,N_42125);
nor UO_4480 (O_4480,N_49644,N_42133);
nor UO_4481 (O_4481,N_40621,N_42075);
xor UO_4482 (O_4482,N_44330,N_40582);
xnor UO_4483 (O_4483,N_46233,N_47192);
and UO_4484 (O_4484,N_47762,N_45807);
and UO_4485 (O_4485,N_45151,N_41736);
xor UO_4486 (O_4486,N_49336,N_40839);
and UO_4487 (O_4487,N_48906,N_44310);
xor UO_4488 (O_4488,N_44581,N_41529);
nand UO_4489 (O_4489,N_43056,N_40854);
or UO_4490 (O_4490,N_48048,N_47493);
nor UO_4491 (O_4491,N_42637,N_42700);
nor UO_4492 (O_4492,N_44318,N_47319);
nand UO_4493 (O_4493,N_41453,N_49570);
nand UO_4494 (O_4494,N_46381,N_42344);
and UO_4495 (O_4495,N_44307,N_42690);
or UO_4496 (O_4496,N_48241,N_44842);
or UO_4497 (O_4497,N_48273,N_41633);
nor UO_4498 (O_4498,N_41085,N_46229);
nor UO_4499 (O_4499,N_46454,N_48051);
and UO_4500 (O_4500,N_43273,N_43765);
nand UO_4501 (O_4501,N_42263,N_43443);
nor UO_4502 (O_4502,N_46577,N_45227);
and UO_4503 (O_4503,N_47203,N_43102);
and UO_4504 (O_4504,N_44184,N_40126);
and UO_4505 (O_4505,N_40708,N_40988);
or UO_4506 (O_4506,N_49808,N_49591);
nand UO_4507 (O_4507,N_42836,N_43305);
xor UO_4508 (O_4508,N_45044,N_41000);
and UO_4509 (O_4509,N_43891,N_41727);
nand UO_4510 (O_4510,N_44817,N_41268);
nand UO_4511 (O_4511,N_42227,N_43788);
and UO_4512 (O_4512,N_44925,N_49436);
and UO_4513 (O_4513,N_41255,N_43041);
nand UO_4514 (O_4514,N_46898,N_42015);
nand UO_4515 (O_4515,N_45589,N_49857);
xnor UO_4516 (O_4516,N_48418,N_42875);
nor UO_4517 (O_4517,N_48869,N_49545);
or UO_4518 (O_4518,N_47219,N_43619);
nor UO_4519 (O_4519,N_42992,N_44560);
nand UO_4520 (O_4520,N_44112,N_40042);
nor UO_4521 (O_4521,N_48856,N_42586);
xnor UO_4522 (O_4522,N_41560,N_46113);
or UO_4523 (O_4523,N_46629,N_47200);
nor UO_4524 (O_4524,N_44709,N_41668);
nand UO_4525 (O_4525,N_41940,N_40379);
and UO_4526 (O_4526,N_40685,N_40740);
and UO_4527 (O_4527,N_42716,N_40380);
or UO_4528 (O_4528,N_48128,N_48274);
and UO_4529 (O_4529,N_43406,N_45891);
xnor UO_4530 (O_4530,N_48195,N_41619);
or UO_4531 (O_4531,N_40431,N_44098);
nand UO_4532 (O_4532,N_42120,N_49111);
nand UO_4533 (O_4533,N_41501,N_46117);
xnor UO_4534 (O_4534,N_45006,N_41445);
nand UO_4535 (O_4535,N_46946,N_44884);
or UO_4536 (O_4536,N_40135,N_41179);
nor UO_4537 (O_4537,N_41910,N_46604);
nor UO_4538 (O_4538,N_47587,N_42292);
or UO_4539 (O_4539,N_46603,N_49003);
xnor UO_4540 (O_4540,N_41298,N_49643);
and UO_4541 (O_4541,N_43229,N_41116);
or UO_4542 (O_4542,N_42735,N_40320);
xor UO_4543 (O_4543,N_47611,N_46875);
nand UO_4544 (O_4544,N_43544,N_40787);
nand UO_4545 (O_4545,N_45386,N_43780);
nand UO_4546 (O_4546,N_48569,N_42930);
nor UO_4547 (O_4547,N_48439,N_41038);
xor UO_4548 (O_4548,N_41514,N_45552);
or UO_4549 (O_4549,N_44141,N_40247);
xor UO_4550 (O_4550,N_44183,N_47264);
and UO_4551 (O_4551,N_43331,N_43538);
nor UO_4552 (O_4552,N_48647,N_48776);
and UO_4553 (O_4553,N_47983,N_41216);
or UO_4554 (O_4554,N_47680,N_48991);
and UO_4555 (O_4555,N_44668,N_44013);
or UO_4556 (O_4556,N_44324,N_49349);
xnor UO_4557 (O_4557,N_40280,N_40753);
xnor UO_4558 (O_4558,N_40095,N_45324);
nand UO_4559 (O_4559,N_46143,N_47627);
nor UO_4560 (O_4560,N_44026,N_49399);
nand UO_4561 (O_4561,N_46341,N_42443);
nand UO_4562 (O_4562,N_49914,N_40914);
and UO_4563 (O_4563,N_40161,N_46930);
nor UO_4564 (O_4564,N_40755,N_41904);
nand UO_4565 (O_4565,N_43469,N_49811);
and UO_4566 (O_4566,N_47860,N_44984);
or UO_4567 (O_4567,N_40762,N_46506);
xor UO_4568 (O_4568,N_46656,N_40110);
nand UO_4569 (O_4569,N_41477,N_48175);
xnor UO_4570 (O_4570,N_45706,N_47206);
xor UO_4571 (O_4571,N_42652,N_48491);
xnor UO_4572 (O_4572,N_44716,N_42606);
xnor UO_4573 (O_4573,N_40857,N_42270);
nor UO_4574 (O_4574,N_48231,N_43996);
nor UO_4575 (O_4575,N_45046,N_45864);
and UO_4576 (O_4576,N_41367,N_40691);
xnor UO_4577 (O_4577,N_44397,N_46446);
or UO_4578 (O_4578,N_45682,N_46015);
xor UO_4579 (O_4579,N_41169,N_46955);
nor UO_4580 (O_4580,N_47571,N_40205);
or UO_4581 (O_4581,N_40458,N_43396);
or UO_4582 (O_4582,N_45618,N_42477);
and UO_4583 (O_4583,N_49109,N_40158);
xor UO_4584 (O_4584,N_45904,N_41996);
nand UO_4585 (O_4585,N_43863,N_45962);
and UO_4586 (O_4586,N_41764,N_46234);
or UO_4587 (O_4587,N_40241,N_47386);
nor UO_4588 (O_4588,N_42485,N_49473);
nand UO_4589 (O_4589,N_42025,N_49001);
and UO_4590 (O_4590,N_45968,N_47052);
and UO_4591 (O_4591,N_41602,N_48832);
and UO_4592 (O_4592,N_49856,N_44367);
nand UO_4593 (O_4593,N_47843,N_46906);
nand UO_4594 (O_4594,N_44329,N_42945);
nand UO_4595 (O_4595,N_48968,N_44025);
nor UO_4596 (O_4596,N_43825,N_41023);
or UO_4597 (O_4597,N_41347,N_48020);
nand UO_4598 (O_4598,N_46570,N_40665);
and UO_4599 (O_4599,N_40201,N_42043);
and UO_4600 (O_4600,N_46282,N_44854);
nor UO_4601 (O_4601,N_49469,N_40729);
and UO_4602 (O_4602,N_48379,N_40935);
or UO_4603 (O_4603,N_42968,N_45264);
nor UO_4604 (O_4604,N_40686,N_43017);
nand UO_4605 (O_4605,N_42197,N_47566);
or UO_4606 (O_4606,N_42838,N_48285);
or UO_4607 (O_4607,N_48080,N_45295);
and UO_4608 (O_4608,N_47703,N_40728);
xor UO_4609 (O_4609,N_43094,N_40677);
or UO_4610 (O_4610,N_42241,N_48691);
or UO_4611 (O_4611,N_44618,N_46204);
or UO_4612 (O_4612,N_41018,N_49518);
nand UO_4613 (O_4613,N_43563,N_48701);
nand UO_4614 (O_4614,N_43163,N_40152);
xor UO_4615 (O_4615,N_47710,N_42937);
and UO_4616 (O_4616,N_44117,N_40104);
or UO_4617 (O_4617,N_49379,N_47086);
nand UO_4618 (O_4618,N_43654,N_47307);
nor UO_4619 (O_4619,N_42610,N_42603);
and UO_4620 (O_4620,N_46931,N_49490);
and UO_4621 (O_4621,N_47966,N_44452);
or UO_4622 (O_4622,N_47488,N_45698);
nand UO_4623 (O_4623,N_45176,N_41294);
or UO_4624 (O_4624,N_40477,N_45939);
nor UO_4625 (O_4625,N_47567,N_48206);
or UO_4626 (O_4626,N_41273,N_47620);
and UO_4627 (O_4627,N_48387,N_47440);
xor UO_4628 (O_4628,N_49882,N_46981);
nor UO_4629 (O_4629,N_40868,N_41227);
nor UO_4630 (O_4630,N_46527,N_45868);
xnor UO_4631 (O_4631,N_48623,N_44224);
and UO_4632 (O_4632,N_48366,N_43313);
xnor UO_4633 (O_4633,N_46209,N_42796);
or UO_4634 (O_4634,N_47686,N_49453);
nand UO_4635 (O_4635,N_43972,N_41853);
xnor UO_4636 (O_4636,N_45310,N_44816);
nor UO_4637 (O_4637,N_48083,N_40482);
nor UO_4638 (O_4638,N_40570,N_46247);
and UO_4639 (O_4639,N_44640,N_45803);
nor UO_4640 (O_4640,N_44725,N_42137);
nor UO_4641 (O_4641,N_43108,N_45345);
nand UO_4642 (O_4642,N_44110,N_41037);
nor UO_4643 (O_4643,N_49541,N_47830);
xor UO_4644 (O_4644,N_49356,N_44363);
xnor UO_4645 (O_4645,N_45255,N_46834);
and UO_4646 (O_4646,N_43963,N_47069);
and UO_4647 (O_4647,N_46804,N_41439);
and UO_4648 (O_4648,N_41184,N_43125);
nand UO_4649 (O_4649,N_42114,N_45547);
and UO_4650 (O_4650,N_45958,N_42104);
xor UO_4651 (O_4651,N_46838,N_49776);
or UO_4652 (O_4652,N_42356,N_42076);
nand UO_4653 (O_4653,N_42626,N_49315);
nand UO_4654 (O_4654,N_47171,N_42269);
nor UO_4655 (O_4655,N_48593,N_41596);
nand UO_4656 (O_4656,N_47149,N_45830);
and UO_4657 (O_4657,N_46852,N_47729);
and UO_4658 (O_4658,N_44488,N_49141);
or UO_4659 (O_4659,N_42856,N_47364);
nor UO_4660 (O_4660,N_48470,N_47040);
nor UO_4661 (O_4661,N_46452,N_43089);
nor UO_4662 (O_4662,N_42013,N_45454);
and UO_4663 (O_4663,N_47348,N_44426);
xor UO_4664 (O_4664,N_43593,N_40980);
and UO_4665 (O_4665,N_42182,N_48475);
nor UO_4666 (O_4666,N_44944,N_40682);
nand UO_4667 (O_4667,N_46790,N_44820);
nand UO_4668 (O_4668,N_40429,N_49271);
nand UO_4669 (O_4669,N_49178,N_48560);
nor UO_4670 (O_4670,N_45540,N_43356);
nor UO_4671 (O_4671,N_47727,N_46332);
or UO_4672 (O_4672,N_46463,N_44466);
nand UO_4673 (O_4673,N_43362,N_49522);
nand UO_4674 (O_4674,N_43448,N_43183);
xnor UO_4675 (O_4675,N_47292,N_45612);
nor UO_4676 (O_4676,N_45085,N_40044);
nand UO_4677 (O_4677,N_42559,N_43719);
or UO_4678 (O_4678,N_45957,N_47458);
or UO_4679 (O_4679,N_46156,N_41964);
or UO_4680 (O_4680,N_45607,N_45571);
or UO_4681 (O_4681,N_46995,N_42482);
nand UO_4682 (O_4682,N_41752,N_43380);
and UO_4683 (O_4683,N_40533,N_47813);
xor UO_4684 (O_4684,N_40203,N_48353);
nor UO_4685 (O_4685,N_44234,N_41437);
nor UO_4686 (O_4686,N_47650,N_42481);
nand UO_4687 (O_4687,N_42689,N_42294);
xor UO_4688 (O_4688,N_47370,N_47722);
nand UO_4689 (O_4689,N_48903,N_49434);
or UO_4690 (O_4690,N_49187,N_45170);
xnor UO_4691 (O_4691,N_48523,N_41898);
nand UO_4692 (O_4692,N_44489,N_45543);
xnor UO_4693 (O_4693,N_41785,N_47923);
nor UO_4694 (O_4694,N_40438,N_41098);
and UO_4695 (O_4695,N_49546,N_47937);
and UO_4696 (O_4696,N_44758,N_44011);
and UO_4697 (O_4697,N_49576,N_41366);
nor UO_4698 (O_4698,N_47802,N_41377);
nor UO_4699 (O_4699,N_40966,N_42283);
nand UO_4700 (O_4700,N_41946,N_44575);
nand UO_4701 (O_4701,N_46999,N_43627);
nand UO_4702 (O_4702,N_43546,N_46933);
and UO_4703 (O_4703,N_48916,N_45683);
xnor UO_4704 (O_4704,N_44992,N_49767);
xnor UO_4705 (O_4705,N_46650,N_49786);
and UO_4706 (O_4706,N_45867,N_47309);
xor UO_4707 (O_4707,N_42954,N_41932);
xor UO_4708 (O_4708,N_46706,N_41921);
nor UO_4709 (O_4709,N_45916,N_42067);
or UO_4710 (O_4710,N_47255,N_45124);
nand UO_4711 (O_4711,N_47482,N_42055);
nand UO_4712 (O_4712,N_43407,N_42600);
nor UO_4713 (O_4713,N_46757,N_45371);
and UO_4714 (O_4714,N_46268,N_46800);
nor UO_4715 (O_4715,N_44591,N_43332);
or UO_4716 (O_4716,N_46998,N_40466);
nor UO_4717 (O_4717,N_44483,N_48833);
or UO_4718 (O_4718,N_41517,N_47738);
xnor UO_4719 (O_4719,N_43204,N_46582);
or UO_4720 (O_4720,N_40274,N_40344);
nand UO_4721 (O_4721,N_42916,N_45286);
or UO_4722 (O_4722,N_41915,N_49127);
xor UO_4723 (O_4723,N_41547,N_47671);
and UO_4724 (O_4724,N_42777,N_48341);
nor UO_4725 (O_4725,N_45419,N_41236);
xnor UO_4726 (O_4726,N_47148,N_47737);
nor UO_4727 (O_4727,N_45782,N_43337);
xor UO_4728 (O_4728,N_41486,N_44770);
or UO_4729 (O_4729,N_49422,N_42833);
nand UO_4730 (O_4730,N_42917,N_42826);
and UO_4731 (O_4731,N_48415,N_41133);
nand UO_4732 (O_4732,N_48047,N_47693);
xnor UO_4733 (O_4733,N_48673,N_49040);
nor UO_4734 (O_4734,N_48855,N_45545);
and UO_4735 (O_4735,N_46823,N_48342);
or UO_4736 (O_4736,N_46241,N_41390);
nor UO_4737 (O_4737,N_46855,N_47011);
nand UO_4738 (O_4738,N_42486,N_40299);
nor UO_4739 (O_4739,N_42927,N_44851);
or UO_4740 (O_4740,N_44970,N_41715);
xor UO_4741 (O_4741,N_42187,N_43421);
nand UO_4742 (O_4742,N_48228,N_49175);
and UO_4743 (O_4743,N_45679,N_42825);
nand UO_4744 (O_4744,N_43722,N_43551);
or UO_4745 (O_4745,N_44736,N_42069);
or UO_4746 (O_4746,N_46306,N_46643);
xor UO_4747 (O_4747,N_48477,N_47692);
nor UO_4748 (O_4748,N_41421,N_45280);
xnor UO_4749 (O_4749,N_49172,N_40081);
nand UO_4750 (O_4750,N_47280,N_40206);
and UO_4751 (O_4751,N_40120,N_45407);
and UO_4752 (O_4752,N_40719,N_43231);
or UO_4753 (O_4753,N_47893,N_42997);
or UO_4754 (O_4754,N_45990,N_40180);
nor UO_4755 (O_4755,N_44493,N_42290);
nand UO_4756 (O_4756,N_42538,N_41722);
or UO_4757 (O_4757,N_46667,N_43398);
and UO_4758 (O_4758,N_42643,N_40413);
nand UO_4759 (O_4759,N_46327,N_47001);
and UO_4760 (O_4760,N_48091,N_40530);
xnor UO_4761 (O_4761,N_45568,N_45502);
or UO_4762 (O_4762,N_46195,N_40165);
or UO_4763 (O_4763,N_42045,N_41805);
nand UO_4764 (O_4764,N_44965,N_45284);
nor UO_4765 (O_4765,N_46718,N_41589);
nand UO_4766 (O_4766,N_46743,N_41462);
nand UO_4767 (O_4767,N_46375,N_48119);
and UO_4768 (O_4768,N_49710,N_46384);
or UO_4769 (O_4769,N_40066,N_47604);
nor UO_4770 (O_4770,N_48049,N_45244);
or UO_4771 (O_4771,N_43340,N_43119);
or UO_4772 (O_4772,N_46707,N_44534);
xor UO_4773 (O_4773,N_42032,N_40960);
or UO_4774 (O_4774,N_48970,N_49043);
and UO_4775 (O_4775,N_43444,N_41684);
nor UO_4776 (O_4776,N_43159,N_40456);
xnor UO_4777 (O_4777,N_42126,N_44276);
nor UO_4778 (O_4778,N_49754,N_44359);
and UO_4779 (O_4779,N_44738,N_48480);
nand UO_4780 (O_4780,N_42684,N_49480);
xnor UO_4781 (O_4781,N_44302,N_44831);
nor UO_4782 (O_4782,N_42755,N_40019);
or UO_4783 (O_4783,N_49661,N_44221);
and UO_4784 (O_4784,N_42365,N_48596);
nor UO_4785 (O_4785,N_45393,N_42456);
or UO_4786 (O_4786,N_46177,N_40116);
nor UO_4787 (O_4787,N_42122,N_49032);
or UO_4788 (O_4788,N_47330,N_45300);
xnor UO_4789 (O_4789,N_49033,N_49852);
nand UO_4790 (O_4790,N_48682,N_40942);
and UO_4791 (O_4791,N_43128,N_42498);
and UO_4792 (O_4792,N_40573,N_46472);
nor UO_4793 (O_4793,N_40940,N_46207);
nand UO_4794 (O_4794,N_44220,N_42820);
xnor UO_4795 (O_4795,N_46052,N_43942);
nand UO_4796 (O_4796,N_42421,N_48001);
nor UO_4797 (O_4797,N_47856,N_46708);
or UO_4798 (O_4798,N_40593,N_46250);
and UO_4799 (O_4799,N_44529,N_40084);
or UO_4800 (O_4800,N_44650,N_47434);
or UO_4801 (O_4801,N_41808,N_48103);
nor UO_4802 (O_4802,N_44354,N_48785);
or UO_4803 (O_4803,N_43813,N_45856);
nor UO_4804 (O_4804,N_42234,N_46557);
xnor UO_4805 (O_4805,N_42362,N_41186);
or UO_4806 (O_4806,N_42420,N_48351);
or UO_4807 (O_4807,N_45171,N_43038);
or UO_4808 (O_4808,N_42383,N_44408);
and UO_4809 (O_4809,N_49618,N_44315);
xnor UO_4810 (O_4810,N_48309,N_46386);
xnor UO_4811 (O_4811,N_45452,N_44514);
or UO_4812 (O_4812,N_45630,N_45751);
nor UO_4813 (O_4813,N_41667,N_48108);
nand UO_4814 (O_4814,N_41725,N_42493);
xor UO_4815 (O_4815,N_43280,N_47507);
nand UO_4816 (O_4816,N_40898,N_43104);
and UO_4817 (O_4817,N_48890,N_49439);
nand UO_4818 (O_4818,N_41524,N_48459);
nor UO_4819 (O_4819,N_47174,N_41680);
xor UO_4820 (O_4820,N_49390,N_40313);
and UO_4821 (O_4821,N_49207,N_49012);
nor UO_4822 (O_4822,N_48940,N_49930);
and UO_4823 (O_4823,N_41967,N_40786);
xnor UO_4824 (O_4824,N_49362,N_49098);
nor UO_4825 (O_4825,N_48322,N_40300);
nand UO_4826 (O_4826,N_40258,N_49022);
and UO_4827 (O_4827,N_44039,N_42275);
nor UO_4828 (O_4828,N_43214,N_40001);
nand UO_4829 (O_4829,N_47875,N_42343);
or UO_4830 (O_4830,N_40565,N_49420);
or UO_4831 (O_4831,N_44798,N_49460);
xor UO_4832 (O_4832,N_41323,N_44388);
xnor UO_4833 (O_4833,N_45200,N_46668);
nand UO_4834 (O_4834,N_49814,N_41621);
xnor UO_4835 (O_4835,N_46240,N_45387);
and UO_4836 (O_4836,N_44883,N_45060);
and UO_4837 (O_4837,N_45338,N_45515);
or UO_4838 (O_4838,N_43226,N_47209);
nand UO_4839 (O_4839,N_48338,N_40272);
nor UO_4840 (O_4840,N_47772,N_44125);
nor UO_4841 (O_4841,N_45162,N_46880);
nand UO_4842 (O_4842,N_45858,N_40903);
and UO_4843 (O_4843,N_47880,N_40100);
and UO_4844 (O_4844,N_44602,N_49876);
xnor UO_4845 (O_4845,N_44230,N_47975);
xnor UO_4846 (O_4846,N_43992,N_45539);
xor UO_4847 (O_4847,N_48472,N_43526);
and UO_4848 (O_4848,N_40880,N_49542);
and UO_4849 (O_4849,N_40136,N_42199);
nor UO_4850 (O_4850,N_44734,N_47582);
or UO_4851 (O_4851,N_43740,N_42202);
and UO_4852 (O_4852,N_42145,N_40847);
xnor UO_4853 (O_4853,N_45128,N_44828);
nor UO_4854 (O_4854,N_44177,N_40820);
xnor UO_4855 (O_4855,N_46200,N_46651);
xnor UO_4856 (O_4856,N_45104,N_40678);
nor UO_4857 (O_4857,N_48698,N_40534);
nor UO_4858 (O_4858,N_45932,N_41075);
or UO_4859 (O_4859,N_41165,N_48828);
nand UO_4860 (O_4860,N_48695,N_41708);
nor UO_4861 (O_4861,N_41467,N_49193);
nor UO_4862 (O_4862,N_47954,N_44219);
nor UO_4863 (O_4863,N_43445,N_49770);
nor UO_4864 (O_4864,N_48670,N_43584);
nand UO_4865 (O_4865,N_40644,N_45995);
xnor UO_4866 (O_4866,N_43960,N_47184);
or UO_4867 (O_4867,N_41041,N_43606);
nor UO_4868 (O_4868,N_44473,N_48250);
xnor UO_4869 (O_4869,N_43505,N_44568);
or UO_4870 (O_4870,N_44523,N_40488);
nand UO_4871 (O_4871,N_49523,N_45010);
and UO_4872 (O_4872,N_47356,N_43494);
nand UO_4873 (O_4873,N_49395,N_42658);
nor UO_4874 (O_4874,N_41162,N_41878);
and UO_4875 (O_4875,N_42914,N_45294);
and UO_4876 (O_4876,N_45139,N_46896);
nor UO_4877 (O_4877,N_49255,N_49378);
nor UO_4878 (O_4878,N_44870,N_48136);
or UO_4879 (O_4879,N_42505,N_42386);
and UO_4880 (O_4880,N_47193,N_46294);
nor UO_4881 (O_4881,N_45687,N_43499);
nand UO_4882 (O_4882,N_42701,N_48193);
or UO_4883 (O_4883,N_49784,N_44120);
xor UO_4884 (O_4884,N_41080,N_41614);
or UO_4885 (O_4885,N_44022,N_46813);
and UO_4886 (O_4886,N_44642,N_48324);
or UO_4887 (O_4887,N_42845,N_41675);
xnor UO_4888 (O_4888,N_46647,N_42170);
or UO_4889 (O_4889,N_44279,N_46313);
or UO_4890 (O_4890,N_47163,N_42763);
xnor UO_4891 (O_4891,N_44258,N_46407);
xor UO_4892 (O_4892,N_44991,N_40200);
nand UO_4893 (O_4893,N_49027,N_47549);
xor UO_4894 (O_4894,N_45561,N_42053);
xor UO_4895 (O_4895,N_41900,N_43267);
xor UO_4896 (O_4896,N_49500,N_46048);
or UO_4897 (O_4897,N_45204,N_40393);
or UO_4898 (O_4898,N_48961,N_47204);
nand UO_4899 (O_4899,N_46745,N_41987);
and UO_4900 (O_4900,N_44111,N_46895);
and UO_4901 (O_4901,N_47027,N_43049);
nand UO_4902 (O_4902,N_42823,N_41496);
and UO_4903 (O_4903,N_47748,N_42565);
nand UO_4904 (O_4904,N_40826,N_46724);
or UO_4905 (O_4905,N_49678,N_48740);
nand UO_4906 (O_4906,N_47550,N_45752);
and UO_4907 (O_4907,N_43401,N_46897);
nor UO_4908 (O_4908,N_48590,N_48368);
xnor UO_4909 (O_4909,N_44357,N_41331);
or UO_4910 (O_4910,N_49847,N_48652);
and UO_4911 (O_4911,N_44203,N_45008);
or UO_4912 (O_4912,N_42221,N_41275);
nand UO_4913 (O_4913,N_43919,N_42955);
nor UO_4914 (O_4914,N_47439,N_48807);
nand UO_4915 (O_4915,N_41622,N_44682);
or UO_4916 (O_4916,N_45347,N_44553);
xnor UO_4917 (O_4917,N_43647,N_44907);
nand UO_4918 (O_4918,N_42632,N_41682);
nand UO_4919 (O_4919,N_43158,N_43655);
or UO_4920 (O_4920,N_44506,N_41776);
nor UO_4921 (O_4921,N_47265,N_44911);
or UO_4922 (O_4922,N_40642,N_48707);
xnor UO_4923 (O_4923,N_47465,N_40209);
nor UO_4924 (O_4924,N_46305,N_44288);
nor UO_4925 (O_4925,N_43841,N_48744);
xnor UO_4926 (O_4926,N_46183,N_42669);
nor UO_4927 (O_4927,N_41134,N_41761);
xor UO_4928 (O_4928,N_44973,N_40240);
or UO_4929 (O_4929,N_48295,N_40423);
and UO_4930 (O_4930,N_40479,N_41704);
and UO_4931 (O_4931,N_44531,N_49489);
xor UO_4932 (O_4932,N_43761,N_46129);
nor UO_4933 (O_4933,N_40473,N_49384);
xor UO_4934 (O_4934,N_42788,N_45678);
or UO_4935 (O_4935,N_47335,N_42543);
nor UO_4936 (O_4936,N_45018,N_42472);
nor UO_4937 (O_4937,N_49731,N_45964);
nor UO_4938 (O_4938,N_47198,N_49147);
nor UO_4939 (O_4939,N_46409,N_43071);
or UO_4940 (O_4940,N_46483,N_48579);
or UO_4941 (O_4941,N_44463,N_49703);
nand UO_4942 (O_4942,N_49962,N_46394);
and UO_4943 (O_4943,N_41475,N_47700);
or UO_4944 (O_4944,N_42041,N_49765);
nor UO_4945 (O_4945,N_41648,N_43409);
nor UO_4946 (O_4946,N_48718,N_46010);
and UO_4947 (O_4947,N_49734,N_43098);
and UO_4948 (O_4948,N_43710,N_42857);
nor UO_4949 (O_4949,N_42357,N_41448);
xnor UO_4950 (O_4950,N_48162,N_48096);
xnor UO_4951 (O_4951,N_41819,N_45178);
xnor UO_4952 (O_4952,N_43212,N_40074);
nand UO_4953 (O_4953,N_48962,N_42650);
and UO_4954 (O_4954,N_46956,N_48974);
xor UO_4955 (O_4955,N_42289,N_42243);
or UO_4956 (O_4956,N_46547,N_42473);
nor UO_4957 (O_4957,N_43948,N_43314);
nand UO_4958 (O_4958,N_40420,N_49810);
xnor UO_4959 (O_4959,N_47044,N_40655);
nand UO_4960 (O_4960,N_47968,N_44699);
xnor UO_4961 (O_4961,N_42730,N_42752);
nand UO_4962 (O_4962,N_49437,N_44195);
nand UO_4963 (O_4963,N_44503,N_43577);
xor UO_4964 (O_4964,N_47993,N_49024);
nand UO_4965 (O_4965,N_43888,N_44291);
nand UO_4966 (O_4966,N_41054,N_43990);
xor UO_4967 (O_4967,N_49988,N_42211);
and UO_4968 (O_4968,N_43205,N_46307);
and UO_4969 (O_4969,N_41313,N_43149);
nor UO_4970 (O_4970,N_40157,N_44202);
nor UO_4971 (O_4971,N_43334,N_40386);
or UO_4972 (O_4972,N_48680,N_48947);
xnor UO_4973 (O_4973,N_44505,N_44284);
nand UO_4974 (O_4974,N_40715,N_47372);
nor UO_4975 (O_4975,N_47591,N_46975);
or UO_4976 (O_4976,N_49760,N_46636);
or UO_4977 (O_4977,N_42349,N_49491);
and UO_4978 (O_4978,N_47164,N_46140);
and UO_4979 (O_4979,N_45370,N_42512);
or UO_4980 (O_4980,N_44470,N_41464);
nand UO_4981 (O_4981,N_44879,N_43552);
and UO_4982 (O_4982,N_46422,N_47838);
xor UO_4983 (O_4983,N_48151,N_41473);
xnor UO_4984 (O_4984,N_48284,N_43933);
nor UO_4985 (O_4985,N_49982,N_46014);
nor UO_4986 (O_4986,N_44885,N_48006);
xnor UO_4987 (O_4987,N_46948,N_49114);
nor UO_4988 (O_4988,N_43669,N_44499);
and UO_4989 (O_4989,N_43319,N_49669);
nor UO_4990 (O_4990,N_47660,N_42010);
and UO_4991 (O_4991,N_46761,N_47547);
and UO_4992 (O_4992,N_47623,N_45160);
nand UO_4993 (O_4993,N_44551,N_49275);
nor UO_4994 (O_4994,N_46462,N_48781);
and UO_4995 (O_4995,N_49563,N_40015);
nor UO_4996 (O_4996,N_47277,N_45368);
or UO_4997 (O_4997,N_43542,N_42389);
or UO_4998 (O_4998,N_44059,N_49465);
nand UO_4999 (O_4999,N_42018,N_41231);
endmodule