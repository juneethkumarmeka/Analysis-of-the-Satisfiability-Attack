module basic_1500_15000_2000_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1190,In_1438);
or U1 (N_1,In_825,In_786);
nor U2 (N_2,In_1155,In_608);
and U3 (N_3,In_762,In_595);
or U4 (N_4,In_534,In_85);
or U5 (N_5,In_943,In_1430);
nand U6 (N_6,In_927,In_1004);
and U7 (N_7,In_620,In_1020);
or U8 (N_8,In_1059,In_1393);
nor U9 (N_9,In_1118,In_430);
nand U10 (N_10,In_143,In_326);
nor U11 (N_11,In_1209,In_1019);
xnor U12 (N_12,In_156,In_310);
nand U13 (N_13,In_767,In_533);
or U14 (N_14,In_1226,In_1062);
nor U15 (N_15,In_94,In_72);
nor U16 (N_16,In_850,In_37);
and U17 (N_17,In_493,In_538);
nand U18 (N_18,In_868,In_59);
nand U19 (N_19,In_983,In_33);
or U20 (N_20,In_691,In_1409);
nand U21 (N_21,In_295,In_11);
or U22 (N_22,In_896,In_886);
and U23 (N_23,In_1424,In_1367);
and U24 (N_24,In_75,In_1244);
and U25 (N_25,In_1181,In_700);
or U26 (N_26,In_734,In_346);
xnor U27 (N_27,In_340,In_571);
xor U28 (N_28,In_1414,In_139);
or U29 (N_29,In_1324,In_1405);
nor U30 (N_30,In_1309,In_677);
nor U31 (N_31,In_584,In_628);
nand U32 (N_32,In_312,In_31);
nand U33 (N_33,In_502,In_759);
nand U34 (N_34,In_205,In_427);
nor U35 (N_35,In_409,In_758);
nor U36 (N_36,In_577,In_977);
nand U37 (N_37,In_806,In_875);
nand U38 (N_38,In_1386,In_1021);
or U39 (N_39,In_275,In_802);
or U40 (N_40,In_1453,In_258);
and U41 (N_41,In_58,In_1331);
nand U42 (N_42,In_36,In_711);
nor U43 (N_43,In_385,In_589);
nand U44 (N_44,In_1216,In_892);
and U45 (N_45,In_261,In_622);
or U46 (N_46,In_1197,In_764);
and U47 (N_47,In_1379,In_1033);
nand U48 (N_48,In_390,In_352);
or U49 (N_49,In_551,In_1345);
nand U50 (N_50,In_980,In_387);
or U51 (N_51,In_226,In_720);
or U52 (N_52,In_173,In_1201);
or U53 (N_53,In_463,In_138);
or U54 (N_54,In_1093,In_997);
nand U55 (N_55,In_922,In_1317);
xor U56 (N_56,In_154,In_467);
and U57 (N_57,In_1225,In_1032);
and U58 (N_58,In_456,In_280);
and U59 (N_59,In_1422,In_1109);
xnor U60 (N_60,In_1352,In_547);
xor U61 (N_61,In_626,In_634);
nor U62 (N_62,In_1389,In_1227);
nand U63 (N_63,In_313,In_130);
and U64 (N_64,In_640,In_871);
or U65 (N_65,In_1494,In_214);
xnor U66 (N_66,In_747,In_650);
and U67 (N_67,In_392,In_837);
xnor U68 (N_68,In_350,In_1192);
or U69 (N_69,In_245,In_1290);
or U70 (N_70,In_1125,In_457);
and U71 (N_71,In_207,In_356);
xnor U72 (N_72,In_1465,In_1314);
nor U73 (N_73,In_1188,In_100);
xor U74 (N_74,In_241,In_916);
or U75 (N_75,In_972,In_1497);
xnor U76 (N_76,In_57,In_1126);
nor U77 (N_77,In_317,In_1428);
and U78 (N_78,In_1463,In_674);
or U79 (N_79,In_729,In_1137);
nand U80 (N_80,In_632,In_668);
or U81 (N_81,In_363,In_482);
and U82 (N_82,In_591,In_775);
nor U83 (N_83,In_655,In_1274);
or U84 (N_84,In_150,In_1307);
or U85 (N_85,In_1236,In_103);
or U86 (N_86,In_498,In_675);
and U87 (N_87,In_1408,In_598);
nor U88 (N_88,In_600,In_856);
or U89 (N_89,In_670,In_869);
or U90 (N_90,In_1083,In_530);
xnor U91 (N_91,In_88,In_158);
nand U92 (N_92,In_707,In_216);
nor U93 (N_93,In_889,In_21);
or U94 (N_94,In_905,In_1316);
nor U95 (N_95,In_987,In_953);
xor U96 (N_96,In_1143,In_259);
or U97 (N_97,In_680,In_681);
or U98 (N_98,In_172,In_1281);
and U99 (N_99,In_779,In_135);
nand U100 (N_100,In_426,In_781);
or U101 (N_101,In_208,In_958);
nor U102 (N_102,In_537,In_903);
nand U103 (N_103,In_257,In_243);
and U104 (N_104,In_1454,In_564);
nor U105 (N_105,In_4,In_318);
xnor U106 (N_106,In_1223,In_1270);
nor U107 (N_107,In_1182,In_726);
nand U108 (N_108,In_1241,In_1253);
xor U109 (N_109,In_1427,In_851);
or U110 (N_110,In_126,In_353);
and U111 (N_111,In_1263,In_1466);
and U112 (N_112,In_1363,In_422);
or U113 (N_113,In_247,In_1206);
or U114 (N_114,In_204,In_1346);
and U115 (N_115,In_1392,In_177);
and U116 (N_116,In_1005,In_855);
nor U117 (N_117,In_1296,In_1355);
nor U118 (N_118,In_455,In_512);
nand U119 (N_119,In_1339,In_671);
xnor U120 (N_120,In_236,In_448);
nor U121 (N_121,In_828,In_760);
xor U122 (N_122,In_1458,In_82);
nor U123 (N_123,In_937,In_1249);
xnor U124 (N_124,In_840,In_113);
xor U125 (N_125,In_1370,In_813);
and U126 (N_126,In_1315,In_1174);
or U127 (N_127,In_296,In_203);
or U128 (N_128,In_466,In_1057);
nand U129 (N_129,In_266,In_900);
xor U130 (N_130,In_516,In_1031);
or U131 (N_131,In_1202,In_80);
nand U132 (N_132,In_894,In_933);
or U133 (N_133,In_612,In_646);
xnor U134 (N_134,In_787,In_473);
xor U135 (N_135,In_104,In_685);
xor U136 (N_136,In_1425,In_215);
and U137 (N_137,In_507,In_1383);
nand U138 (N_138,In_1489,In_106);
nor U139 (N_139,In_348,In_1419);
and U140 (N_140,In_543,In_621);
nor U141 (N_141,In_879,In_490);
nand U142 (N_142,In_489,In_1158);
nor U143 (N_143,In_400,In_1230);
and U144 (N_144,In_1015,In_220);
nor U145 (N_145,In_1377,In_234);
xnor U146 (N_146,In_238,In_157);
nor U147 (N_147,In_1113,In_1374);
or U148 (N_148,In_952,In_240);
nand U149 (N_149,In_1306,In_373);
or U150 (N_150,In_223,In_785);
and U151 (N_151,In_664,In_1473);
and U152 (N_152,In_1495,In_374);
or U153 (N_153,In_1037,In_845);
xnor U154 (N_154,In_487,In_1214);
or U155 (N_155,In_847,In_102);
nand U156 (N_156,In_239,In_1455);
nor U157 (N_157,In_349,In_1237);
or U158 (N_158,In_594,In_1282);
xnor U159 (N_159,In_343,In_221);
nor U160 (N_160,In_960,In_1287);
or U161 (N_161,In_1448,In_1283);
nor U162 (N_162,In_553,In_155);
nor U163 (N_163,In_185,In_1433);
or U164 (N_164,In_123,In_829);
nand U165 (N_165,In_627,In_1268);
nand U166 (N_166,In_48,In_599);
xor U167 (N_167,In_225,In_902);
or U168 (N_168,In_6,In_345);
xnor U169 (N_169,In_527,In_311);
nand U170 (N_170,In_1360,In_504);
nor U171 (N_171,In_1293,In_890);
nor U172 (N_172,In_125,In_1299);
nand U173 (N_173,In_464,In_909);
or U174 (N_174,In_830,In_1395);
or U175 (N_175,In_821,In_1243);
nand U176 (N_176,In_302,In_590);
nor U177 (N_177,In_1161,In_34);
or U178 (N_178,In_818,In_1460);
nor U179 (N_179,In_682,In_919);
nand U180 (N_180,In_633,In_605);
and U181 (N_181,In_791,In_1277);
nor U182 (N_182,In_683,In_1080);
and U183 (N_183,In_437,In_1045);
xor U184 (N_184,In_406,In_950);
xnor U185 (N_185,In_925,In_478);
xor U186 (N_186,In_74,In_801);
and U187 (N_187,In_1272,In_961);
xnor U188 (N_188,In_1084,In_462);
xor U189 (N_189,In_279,In_1029);
xnor U190 (N_190,In_64,In_66);
or U191 (N_191,In_784,In_1251);
xnor U192 (N_192,In_1207,In_1476);
nor U193 (N_193,In_248,In_63);
nor U194 (N_194,In_260,In_942);
nor U195 (N_195,In_1075,In_141);
nand U196 (N_196,In_1050,In_792);
or U197 (N_197,In_1099,In_1325);
nor U198 (N_198,In_938,In_1341);
nor U199 (N_199,In_1239,In_964);
nand U200 (N_200,In_607,In_486);
nand U201 (N_201,In_1337,In_330);
xnor U202 (N_202,In_81,In_982);
xnor U203 (N_203,In_1364,In_32);
and U204 (N_204,In_0,In_440);
or U205 (N_205,In_1009,In_454);
nor U206 (N_206,In_853,In_1036);
and U207 (N_207,In_689,In_558);
xnor U208 (N_208,In_630,In_403);
nand U209 (N_209,In_857,In_99);
nand U210 (N_210,In_283,In_841);
and U211 (N_211,In_272,In_1231);
or U212 (N_212,In_69,In_1179);
or U213 (N_213,In_499,In_494);
nand U214 (N_214,In_877,In_53);
or U215 (N_215,In_575,In_1399);
and U216 (N_216,In_93,In_859);
and U217 (N_217,In_39,In_610);
or U218 (N_218,In_1396,In_218);
nor U219 (N_219,In_67,In_996);
nor U220 (N_220,In_290,In_323);
and U221 (N_221,In_1048,In_1087);
xor U222 (N_222,In_415,In_271);
or U223 (N_223,In_539,In_649);
xor U224 (N_224,In_265,In_1280);
or U225 (N_225,In_528,In_1413);
nand U226 (N_226,In_1065,In_965);
xor U227 (N_227,In_524,In_1159);
xnor U228 (N_228,In_966,In_161);
or U229 (N_229,In_1139,In_366);
or U230 (N_230,In_705,In_1432);
and U231 (N_231,In_227,In_1286);
xor U232 (N_232,In_1248,In_926);
xnor U233 (N_233,In_321,In_397);
nand U234 (N_234,In_865,In_1371);
or U235 (N_235,In_749,In_56);
nor U236 (N_236,In_181,In_1211);
nand U237 (N_237,In_242,In_176);
nor U238 (N_238,In_453,In_105);
xor U239 (N_239,In_1491,In_957);
nor U240 (N_240,In_255,In_1081);
nor U241 (N_241,In_842,In_274);
xor U242 (N_242,In_1238,In_1097);
nand U243 (N_243,In_95,In_287);
and U244 (N_244,In_1441,In_412);
nor U245 (N_245,In_624,In_885);
xnor U246 (N_246,In_1166,In_1496);
xor U247 (N_247,In_1017,In_369);
and U248 (N_248,In_951,In_219);
nand U249 (N_249,In_96,In_550);
or U250 (N_250,In_424,In_1499);
nand U251 (N_251,In_656,In_128);
xnor U252 (N_252,In_289,In_167);
or U253 (N_253,In_1487,In_755);
xnor U254 (N_254,In_780,In_906);
nor U255 (N_255,In_393,In_924);
xnor U256 (N_256,In_581,In_134);
nor U257 (N_257,In_179,In_1146);
or U258 (N_258,In_1305,In_120);
xor U259 (N_259,In_1298,In_1028);
xor U260 (N_260,In_1076,In_793);
or U261 (N_261,In_79,In_619);
and U262 (N_262,In_20,In_505);
nor U263 (N_263,In_688,In_631);
xor U264 (N_264,In_552,In_963);
or U265 (N_265,In_1149,In_526);
or U266 (N_266,In_1429,In_583);
nor U267 (N_267,In_998,In_519);
nor U268 (N_268,In_77,In_1132);
nor U269 (N_269,In_928,In_800);
nor U270 (N_270,In_1024,In_481);
nand U271 (N_271,In_618,In_693);
xor U272 (N_272,In_1129,In_824);
xor U273 (N_273,In_202,In_1416);
and U274 (N_274,In_1043,In_46);
xor U275 (N_275,In_669,In_1077);
nand U276 (N_276,In_663,In_1276);
or U277 (N_277,In_1407,In_477);
and U278 (N_278,In_1481,In_1189);
nand U279 (N_279,In_285,In_864);
and U280 (N_280,In_1030,In_122);
nand U281 (N_281,In_999,In_70);
nor U282 (N_282,In_661,In_144);
xor U283 (N_283,In_1108,In_1347);
xnor U284 (N_284,In_410,In_1417);
nor U285 (N_285,In_1074,In_1204);
nor U286 (N_286,In_145,In_38);
nand U287 (N_287,In_1470,In_962);
or U288 (N_288,In_485,In_402);
nand U289 (N_289,In_1275,In_1058);
nor U290 (N_290,In_1185,In_362);
and U291 (N_291,In_133,In_573);
and U292 (N_292,In_217,In_382);
nand U293 (N_293,In_338,In_291);
nand U294 (N_294,In_913,In_30);
xor U295 (N_295,In_186,In_1400);
nor U296 (N_296,In_1397,In_1044);
and U297 (N_297,In_1250,In_1119);
and U298 (N_298,In_344,In_1328);
xnor U299 (N_299,In_1114,In_1122);
and U300 (N_300,In_1382,In_375);
or U301 (N_301,In_1456,In_954);
xor U302 (N_302,In_1426,In_1078);
and U303 (N_303,In_1098,In_665);
nand U304 (N_304,In_835,In_1047);
nand U305 (N_305,In_629,In_183);
and U306 (N_306,In_182,In_956);
nand U307 (N_307,In_1449,In_1369);
and U308 (N_308,In_1172,In_1111);
and U309 (N_309,In_1135,In_770);
nand U310 (N_310,In_572,In_672);
and U311 (N_311,In_460,In_833);
nand U312 (N_312,In_267,In_132);
nand U313 (N_313,In_147,In_1040);
and U314 (N_314,In_1421,In_506);
and U315 (N_315,In_1054,In_662);
xnor U316 (N_316,In_191,In_946);
xnor U317 (N_317,In_1284,In_1224);
and U318 (N_318,In_1168,In_1213);
xnor U319 (N_319,In_1349,In_1485);
xor U320 (N_320,In_1008,In_118);
nand U321 (N_321,In_433,In_1488);
xnor U322 (N_322,In_1361,In_1320);
or U323 (N_323,In_615,In_262);
nor U324 (N_324,In_873,In_920);
xnor U325 (N_325,In_399,In_654);
nor U326 (N_326,In_2,In_480);
and U327 (N_327,In_532,In_1138);
xnor U328 (N_328,In_119,In_1215);
xor U329 (N_329,In_394,In_468);
nor U330 (N_330,In_199,In_1252);
nand U331 (N_331,In_1010,In_1235);
nor U332 (N_332,In_163,In_1469);
nor U333 (N_333,In_673,In_389);
nand U334 (N_334,In_587,In_848);
xnor U335 (N_335,In_50,In_1165);
and U336 (N_336,In_423,In_1096);
nor U337 (N_337,In_435,In_1411);
nor U338 (N_338,In_979,In_1447);
nand U339 (N_339,In_1265,In_1060);
and U340 (N_340,In_934,In_153);
nand U341 (N_341,In_372,In_772);
nor U342 (N_342,In_171,In_1141);
or U343 (N_343,In_1446,In_1035);
and U344 (N_344,In_1340,In_1094);
nand U345 (N_345,In_1200,In_503);
and U346 (N_346,In_807,In_686);
xor U347 (N_347,In_1354,In_1356);
and U348 (N_348,In_948,In_1359);
xor U349 (N_349,In_929,In_763);
xnor U350 (N_350,In_836,In_708);
nor U351 (N_351,In_636,In_1082);
or U352 (N_352,In_1203,In_333);
and U353 (N_353,In_798,In_544);
and U354 (N_354,In_395,In_578);
and U355 (N_355,In_783,In_1329);
nand U356 (N_356,In_520,In_1368);
nand U357 (N_357,In_332,In_574);
nand U358 (N_358,In_880,In_593);
nor U359 (N_359,In_174,In_898);
nor U360 (N_360,In_1170,In_12);
and U361 (N_361,In_560,In_131);
and U362 (N_362,In_1333,In_71);
nand U363 (N_363,In_1457,In_55);
nand U364 (N_364,In_442,In_771);
xor U365 (N_365,In_211,In_1480);
nand U366 (N_366,In_715,In_613);
nand U367 (N_367,In_18,In_276);
and U368 (N_368,In_769,In_1003);
nor U369 (N_369,In_107,In_449);
and U370 (N_370,In_178,In_536);
nor U371 (N_371,In_854,In_1343);
or U372 (N_372,In_1322,In_89);
nor U373 (N_373,In_334,In_1388);
or U374 (N_374,In_597,In_367);
xnor U375 (N_375,In_1154,In_495);
and U376 (N_376,In_391,In_730);
nor U377 (N_377,In_315,In_1066);
and U378 (N_378,In_1210,In_244);
or U379 (N_379,In_229,In_1101);
or U380 (N_380,In_418,In_884);
and U381 (N_381,In_405,In_743);
and U382 (N_382,In_557,In_1266);
nor U383 (N_383,In_230,In_774);
nor U384 (N_384,In_465,In_166);
or U385 (N_385,In_434,In_623);
xor U386 (N_386,In_832,In_459);
or U387 (N_387,In_588,In_911);
or U388 (N_388,In_357,In_111);
nor U389 (N_389,In_989,In_320);
or U390 (N_390,In_35,In_509);
xor U391 (N_391,In_701,In_1212);
nand U392 (N_392,In_151,In_510);
nand U393 (N_393,In_1103,In_354);
nand U394 (N_394,In_62,In_1255);
nand U395 (N_395,In_115,In_254);
or U396 (N_396,In_1063,In_1366);
nor U397 (N_397,In_614,In_667);
or U398 (N_398,In_1271,In_1472);
nor U399 (N_399,In_1483,In_1342);
or U400 (N_400,In_136,In_1051);
or U401 (N_401,In_969,In_1171);
xnor U402 (N_402,In_1372,In_168);
or U403 (N_403,In_1150,In_461);
nand U404 (N_404,In_1380,In_531);
xnor U405 (N_405,In_169,In_1326);
xor U406 (N_406,In_149,In_561);
and U407 (N_407,In_1127,In_753);
nor U408 (N_408,In_541,In_947);
or U409 (N_409,In_501,In_1443);
nand U410 (N_410,In_1186,In_407);
xor U411 (N_411,In_562,In_1474);
or U412 (N_412,In_765,In_548);
or U413 (N_413,In_298,In_838);
or U414 (N_414,In_881,In_1313);
or U415 (N_415,In_233,In_192);
or U416 (N_416,In_897,In_1068);
nand U417 (N_417,In_1312,In_1117);
xor U418 (N_418,In_1435,In_728);
and U419 (N_419,In_1398,In_264);
nor U420 (N_420,In_735,In_1319);
nor U421 (N_421,In_224,In_559);
xor U422 (N_422,In_761,In_1195);
nor U423 (N_423,In_907,In_895);
nand U424 (N_424,In_445,In_1387);
or U425 (N_425,In_1144,In_380);
nor U426 (N_426,In_1116,In_1365);
nand U427 (N_427,In_180,In_1440);
or U428 (N_428,In_676,In_336);
or U429 (N_429,In_638,In_794);
and U430 (N_430,In_1431,In_42);
xor U431 (N_431,In_901,In_817);
or U432 (N_432,In_523,In_1471);
nor U433 (N_433,In_849,In_370);
xor U434 (N_434,In_360,In_337);
xor U435 (N_435,In_1136,In_844);
nor U436 (N_436,In_1180,In_1072);
or U437 (N_437,In_827,In_379);
and U438 (N_438,In_1025,In_1308);
nand U439 (N_439,In_251,In_1234);
xnor U440 (N_440,In_732,In_1148);
and U441 (N_441,In_1240,In_250);
and U442 (N_442,In_684,In_874);
nand U443 (N_443,In_371,In_570);
or U444 (N_444,In_1258,In_201);
and U445 (N_445,In_1163,In_307);
nand U446 (N_446,In_910,In_1175);
nand U447 (N_447,In_60,In_1330);
nand U448 (N_448,In_194,In_137);
nor U449 (N_449,In_941,In_1384);
and U450 (N_450,In_1378,In_635);
nand U451 (N_451,In_61,In_811);
nand U452 (N_452,In_1353,In_1436);
nand U453 (N_453,In_441,In_1208);
nand U454 (N_454,In_300,In_1351);
or U455 (N_455,In_44,In_1310);
or U456 (N_456,In_742,In_294);
nand U457 (N_457,In_1285,In_554);
nor U458 (N_458,In_1056,In_1079);
nand U459 (N_459,In_967,In_87);
nand U460 (N_460,In_29,In_1256);
nand U461 (N_461,In_232,In_1478);
and U462 (N_462,In_469,In_757);
xnor U463 (N_463,In_569,In_1198);
or U464 (N_464,In_995,In_696);
and U465 (N_465,In_443,In_1018);
and U466 (N_466,In_648,In_447);
or U467 (N_467,In_8,In_5);
xor U468 (N_468,In_582,In_1022);
and U469 (N_469,In_322,In_789);
and U470 (N_470,In_1042,In_413);
or U471 (N_471,In_1178,In_479);
and U472 (N_472,In_342,In_1162);
nand U473 (N_473,In_117,In_425);
or U474 (N_474,In_1152,In_1145);
or U475 (N_475,In_1402,In_91);
nor U476 (N_476,In_1461,In_1041);
nor U477 (N_477,In_1014,In_450);
and U478 (N_478,In_565,In_1262);
xnor U479 (N_479,In_508,In_316);
and U480 (N_480,In_51,In_994);
xor U481 (N_481,In_1151,In_284);
or U482 (N_482,In_452,In_718);
nor U483 (N_483,In_602,In_973);
xor U484 (N_484,In_745,In_563);
nor U485 (N_485,In_293,In_1247);
nor U486 (N_486,In_808,In_1492);
or U487 (N_487,In_923,In_365);
nor U488 (N_488,In_659,In_883);
nor U489 (N_489,In_1484,In_754);
xor U490 (N_490,In_645,In_568);
nand U491 (N_491,In_603,In_47);
xor U492 (N_492,In_637,In_932);
xor U493 (N_493,In_1477,In_870);
xor U494 (N_494,In_981,In_1067);
and U495 (N_495,In_722,In_1012);
xnor U496 (N_496,In_483,In_992);
nand U497 (N_497,In_347,In_497);
and U498 (N_498,In_709,In_1468);
xnor U499 (N_499,In_1437,In_746);
xor U500 (N_500,In_535,In_1088);
or U501 (N_501,In_1131,In_1112);
nand U502 (N_502,In_10,In_1069);
and U503 (N_503,In_1194,In_488);
xnor U504 (N_504,In_511,In_694);
or U505 (N_505,In_142,In_944);
and U506 (N_506,In_1257,In_1156);
nor U507 (N_507,In_1027,In_1264);
and U508 (N_508,In_97,In_719);
nor U509 (N_509,In_609,In_1311);
and U510 (N_510,In_1090,In_325);
or U511 (N_511,In_1007,In_500);
nand U512 (N_512,In_1157,In_1420);
or U513 (N_513,In_124,In_1321);
or U514 (N_514,In_165,In_852);
nor U515 (N_515,In_329,In_140);
nand U516 (N_516,In_358,In_1376);
nor U517 (N_517,In_384,In_788);
and U518 (N_518,In_175,In_1121);
nand U519 (N_519,In_816,In_1261);
nand U520 (N_520,In_1278,In_304);
nand U521 (N_521,In_1089,In_428);
nor U522 (N_522,In_496,In_1193);
nor U523 (N_523,In_246,In_518);
nor U524 (N_524,In_68,In_1086);
nand U525 (N_525,In_40,In_476);
xnor U526 (N_526,In_1147,In_282);
or U527 (N_527,In_717,In_339);
xnor U528 (N_528,In_23,In_727);
xor U529 (N_529,In_616,In_1184);
or U530 (N_530,In_1301,In_1222);
and U531 (N_531,In_738,In_19);
nand U532 (N_532,In_1292,In_396);
nor U533 (N_533,In_1323,In_1053);
or U534 (N_534,In_699,In_822);
nor U535 (N_535,In_891,In_695);
nand U536 (N_536,In_273,In_1362);
nor U537 (N_537,In_1006,In_1173);
and U538 (N_538,In_408,In_414);
xnor U539 (N_539,In_514,In_733);
or U540 (N_540,In_1100,In_990);
nor U541 (N_541,In_417,In_731);
or U542 (N_542,In_253,In_931);
xor U543 (N_543,In_1073,In_1232);
and U544 (N_544,In_451,In_101);
nand U545 (N_545,In_723,In_839);
or U546 (N_546,In_1196,In_1335);
and U547 (N_547,In_803,In_858);
xnor U548 (N_548,In_268,In_752);
xnor U549 (N_549,In_492,In_567);
or U550 (N_550,In_641,In_692);
nand U551 (N_551,In_739,In_893);
and U552 (N_552,In_796,In_712);
nand U553 (N_553,In_1294,In_741);
xor U554 (N_554,In_585,In_773);
or U555 (N_555,In_22,In_1026);
nor U556 (N_556,In_1260,In_1002);
or U557 (N_557,In_566,In_73);
nor U558 (N_558,In_212,In_474);
nor U559 (N_559,In_15,In_766);
and U560 (N_560,In_1318,In_305);
or U561 (N_561,In_429,In_116);
and U562 (N_562,In_862,In_1442);
nand U563 (N_563,In_197,In_768);
and U564 (N_564,In_127,In_324);
or U565 (N_565,In_1071,In_1479);
nor U566 (N_566,In_431,In_270);
xor U567 (N_567,In_986,In_1183);
and U568 (N_568,In_1085,In_725);
nor U569 (N_569,In_206,In_955);
or U570 (N_570,In_359,In_917);
nor U571 (N_571,In_1242,In_1217);
and U572 (N_572,In_690,In_1273);
xnor U573 (N_573,In_968,In_658);
nor U574 (N_574,In_940,In_866);
nand U575 (N_575,In_878,In_1482);
or U576 (N_576,In_861,In_1344);
nor U577 (N_577,In_41,In_887);
xor U578 (N_578,In_411,In_1358);
nand U579 (N_579,In_625,In_1415);
nor U580 (N_580,In_867,In_1259);
nand U581 (N_581,In_1297,In_912);
nand U582 (N_582,In_388,In_549);
or U583 (N_583,In_3,In_908);
nand U584 (N_584,In_1169,In_1450);
xnor U585 (N_585,In_790,In_200);
or U586 (N_586,In_1475,In_297);
xor U587 (N_587,In_820,In_888);
and U588 (N_588,In_592,In_1038);
nor U589 (N_589,In_596,In_90);
or U590 (N_590,In_930,In_978);
xor U591 (N_591,In_108,In_484);
xor U592 (N_592,In_904,In_1176);
nand U593 (N_593,In_647,In_109);
or U594 (N_594,In_237,In_1115);
or U595 (N_595,In_555,In_1228);
xor U596 (N_596,In_876,In_355);
nor U597 (N_597,In_831,In_446);
nor U598 (N_598,In_28,In_419);
and U599 (N_599,In_642,In_988);
xor U600 (N_600,In_1052,In_1334);
or U601 (N_601,In_1304,In_525);
nor U602 (N_602,In_750,In_309);
xnor U603 (N_603,In_1177,In_744);
and U604 (N_604,In_945,In_1269);
and U605 (N_605,In_1221,In_580);
and U606 (N_606,In_470,In_984);
or U607 (N_607,In_319,In_16);
and U608 (N_608,In_1291,In_7);
or U609 (N_609,In_351,In_1199);
nand U610 (N_610,In_170,In_17);
nand U611 (N_611,In_1034,In_1403);
nor U612 (N_612,In_970,In_834);
xnor U613 (N_613,In_1218,In_991);
xor U614 (N_614,In_1401,In_472);
and U615 (N_615,In_804,In_263);
nor U616 (N_616,In_159,In_809);
nor U617 (N_617,In_1039,In_1046);
xor U618 (N_618,In_601,In_1013);
xnor U619 (N_619,In_1336,In_1061);
nand U620 (N_620,In_1459,In_1357);
or U621 (N_621,In_471,In_1406);
and U622 (N_622,In_1302,In_421);
and U623 (N_623,In_1434,In_328);
xnor U624 (N_624,In_83,In_639);
xnor U625 (N_625,In_439,In_25);
nor U626 (N_626,In_517,In_444);
or U627 (N_627,In_1486,In_756);
nor U628 (N_628,In_196,In_361);
and U629 (N_629,In_935,In_376);
or U630 (N_630,In_160,In_716);
xor U631 (N_631,In_513,In_1153);
xor U632 (N_632,In_529,In_438);
or U633 (N_633,In_974,In_1391);
xnor U634 (N_634,In_1133,In_401);
xor U635 (N_635,In_815,In_235);
or U636 (N_636,In_1464,In_1000);
or U637 (N_637,In_195,In_1160);
xor U638 (N_638,In_914,In_810);
or U639 (N_639,In_281,In_1375);
nor U640 (N_640,In_52,In_1410);
nor U641 (N_641,In_860,In_545);
or U642 (N_642,In_1338,In_846);
nor U643 (N_643,In_737,In_778);
or U644 (N_644,In_1385,In_586);
xor U645 (N_645,In_231,In_1267);
and U646 (N_646,In_331,In_915);
or U647 (N_647,In_651,In_721);
and U648 (N_648,In_1348,In_797);
and U649 (N_649,In_736,In_814);
nand U650 (N_650,In_579,In_706);
nand U651 (N_651,In_985,In_522);
or U652 (N_652,In_92,In_617);
xnor U653 (N_653,In_697,In_1467);
and U654 (N_654,In_776,In_1439);
nor U655 (N_655,In_652,In_187);
nand U656 (N_656,In_1254,In_1);
and U657 (N_657,In_823,In_65);
nand U658 (N_658,In_377,In_26);
or U659 (N_659,In_256,In_740);
or U660 (N_660,In_416,In_54);
nand U661 (N_661,In_43,In_1070);
xor U662 (N_662,In_657,In_611);
nor U663 (N_663,In_209,In_162);
and U664 (N_664,In_278,In_521);
nand U665 (N_665,In_49,In_188);
nand U666 (N_666,In_1102,In_228);
nor U667 (N_667,In_795,In_1219);
or U668 (N_668,In_643,In_378);
xnor U669 (N_669,In_269,In_1493);
and U670 (N_670,In_286,In_1124);
nand U671 (N_671,In_129,In_1300);
nor U672 (N_672,In_1011,In_327);
xnor U673 (N_673,In_1452,In_13);
and U674 (N_674,In_84,In_546);
nor U675 (N_675,In_975,In_1016);
xor U676 (N_676,In_1390,In_404);
xor U677 (N_677,In_1373,In_606);
or U678 (N_678,In_1229,In_899);
nor U679 (N_679,In_198,In_1104);
nor U680 (N_680,In_959,In_812);
or U681 (N_681,In_1220,In_1187);
or U682 (N_682,In_148,In_189);
xor U683 (N_683,In_799,In_515);
and U684 (N_684,In_306,In_704);
and U685 (N_685,In_1327,In_436);
or U686 (N_686,In_491,In_819);
nor U687 (N_687,In_114,In_921);
nand U688 (N_688,In_713,In_1134);
or U689 (N_689,In_301,In_1105);
nor U690 (N_690,In_210,In_1106);
or U691 (N_691,In_303,In_678);
and U692 (N_692,In_213,In_76);
and U693 (N_693,In_653,In_1164);
nand U694 (N_694,In_1490,In_164);
and U695 (N_695,In_748,In_277);
nand U696 (N_696,In_710,In_190);
or U697 (N_697,In_872,In_698);
nor U698 (N_698,In_341,In_1049);
nand U699 (N_699,In_308,In_660);
xnor U700 (N_700,In_381,In_1444);
nand U701 (N_701,In_27,In_1128);
and U702 (N_702,In_540,In_1418);
or U703 (N_703,In_110,In_1303);
and U704 (N_704,In_335,In_1167);
and U705 (N_705,In_936,In_386);
xor U706 (N_706,In_9,In_1289);
or U707 (N_707,In_604,In_777);
or U708 (N_708,In_1123,In_939);
and U709 (N_709,In_1462,In_1110);
or U710 (N_710,In_368,In_971);
nor U711 (N_711,In_1205,In_666);
xnor U712 (N_712,In_863,In_976);
nor U713 (N_713,In_843,In_314);
and U714 (N_714,In_1092,In_98);
nand U715 (N_715,In_1423,In_184);
nand U716 (N_716,In_679,In_805);
and U717 (N_717,In_826,In_1288);
xnor U718 (N_718,In_882,In_1095);
xor U719 (N_719,In_1107,In_1233);
xor U720 (N_720,In_398,In_86);
nor U721 (N_721,In_78,In_687);
and U722 (N_722,In_292,In_724);
and U723 (N_723,In_1451,In_121);
xor U724 (N_724,In_1295,In_1001);
and U725 (N_725,In_364,In_1445);
nand U726 (N_726,In_458,In_576);
xnor U727 (N_727,In_1245,In_432);
nor U728 (N_728,In_383,In_1350);
or U729 (N_729,In_1120,In_45);
nand U730 (N_730,In_24,In_1191);
nor U731 (N_731,In_1412,In_542);
nand U732 (N_732,In_14,In_193);
nor U733 (N_733,In_475,In_1130);
nand U734 (N_734,In_714,In_420);
nor U735 (N_735,In_1498,In_782);
nand U736 (N_736,In_1404,In_1394);
xor U737 (N_737,In_1279,In_1381);
and U738 (N_738,In_644,In_703);
nand U739 (N_739,In_993,In_152);
xor U740 (N_740,In_1091,In_112);
nor U741 (N_741,In_299,In_1140);
nor U742 (N_742,In_751,In_249);
nand U743 (N_743,In_1055,In_288);
nand U744 (N_744,In_1064,In_949);
nand U745 (N_745,In_1332,In_556);
or U746 (N_746,In_702,In_146);
nand U747 (N_747,In_1142,In_918);
or U748 (N_748,In_222,In_1023);
xor U749 (N_749,In_252,In_1246);
xor U750 (N_750,In_1258,In_700);
nand U751 (N_751,In_1037,In_1259);
or U752 (N_752,In_1360,In_511);
and U753 (N_753,In_135,In_1363);
nor U754 (N_754,In_1488,In_571);
or U755 (N_755,In_1069,In_281);
nand U756 (N_756,In_931,In_568);
nand U757 (N_757,In_1329,In_884);
or U758 (N_758,In_517,In_1111);
nor U759 (N_759,In_69,In_340);
nor U760 (N_760,In_6,In_497);
nand U761 (N_761,In_219,In_1050);
or U762 (N_762,In_891,In_964);
nand U763 (N_763,In_1480,In_1044);
or U764 (N_764,In_1198,In_293);
or U765 (N_765,In_476,In_67);
and U766 (N_766,In_725,In_1134);
xor U767 (N_767,In_278,In_438);
xor U768 (N_768,In_13,In_111);
nor U769 (N_769,In_399,In_672);
and U770 (N_770,In_326,In_1481);
and U771 (N_771,In_251,In_1302);
and U772 (N_772,In_714,In_1062);
and U773 (N_773,In_1152,In_1425);
or U774 (N_774,In_953,In_135);
or U775 (N_775,In_780,In_741);
xnor U776 (N_776,In_215,In_1466);
nor U777 (N_777,In_355,In_440);
nor U778 (N_778,In_894,In_297);
nor U779 (N_779,In_68,In_792);
or U780 (N_780,In_48,In_138);
nand U781 (N_781,In_846,In_1223);
nor U782 (N_782,In_1094,In_209);
or U783 (N_783,In_915,In_1267);
or U784 (N_784,In_291,In_189);
nor U785 (N_785,In_433,In_281);
nor U786 (N_786,In_1441,In_1018);
nand U787 (N_787,In_906,In_1171);
nand U788 (N_788,In_1062,In_874);
and U789 (N_789,In_557,In_267);
and U790 (N_790,In_505,In_285);
nor U791 (N_791,In_141,In_102);
nand U792 (N_792,In_933,In_1407);
nand U793 (N_793,In_147,In_974);
or U794 (N_794,In_133,In_167);
xnor U795 (N_795,In_389,In_65);
or U796 (N_796,In_1412,In_1277);
nand U797 (N_797,In_973,In_1365);
nand U798 (N_798,In_453,In_555);
nor U799 (N_799,In_591,In_1218);
nor U800 (N_800,In_312,In_1295);
and U801 (N_801,In_318,In_900);
or U802 (N_802,In_900,In_455);
or U803 (N_803,In_466,In_467);
and U804 (N_804,In_405,In_1256);
xor U805 (N_805,In_1291,In_92);
nand U806 (N_806,In_937,In_71);
nor U807 (N_807,In_564,In_645);
nor U808 (N_808,In_1324,In_1297);
nand U809 (N_809,In_452,In_1331);
and U810 (N_810,In_164,In_1381);
and U811 (N_811,In_937,In_900);
and U812 (N_812,In_899,In_1280);
and U813 (N_813,In_150,In_1410);
nand U814 (N_814,In_359,In_760);
xnor U815 (N_815,In_1160,In_639);
or U816 (N_816,In_460,In_925);
or U817 (N_817,In_567,In_75);
nor U818 (N_818,In_756,In_102);
and U819 (N_819,In_706,In_906);
xor U820 (N_820,In_510,In_44);
nor U821 (N_821,In_1038,In_1362);
nand U822 (N_822,In_851,In_793);
or U823 (N_823,In_195,In_451);
xnor U824 (N_824,In_1224,In_724);
xnor U825 (N_825,In_823,In_1090);
and U826 (N_826,In_78,In_144);
xnor U827 (N_827,In_942,In_1429);
xor U828 (N_828,In_1487,In_1011);
nor U829 (N_829,In_50,In_4);
nor U830 (N_830,In_1278,In_383);
or U831 (N_831,In_550,In_84);
and U832 (N_832,In_1383,In_379);
xnor U833 (N_833,In_92,In_649);
and U834 (N_834,In_1199,In_373);
and U835 (N_835,In_394,In_490);
nand U836 (N_836,In_1356,In_1435);
nor U837 (N_837,In_45,In_817);
nor U838 (N_838,In_400,In_615);
or U839 (N_839,In_164,In_40);
nand U840 (N_840,In_840,In_269);
xnor U841 (N_841,In_413,In_710);
or U842 (N_842,In_64,In_525);
xnor U843 (N_843,In_905,In_332);
nand U844 (N_844,In_391,In_91);
and U845 (N_845,In_421,In_998);
nand U846 (N_846,In_134,In_14);
or U847 (N_847,In_750,In_62);
nor U848 (N_848,In_234,In_1048);
nor U849 (N_849,In_16,In_728);
nor U850 (N_850,In_952,In_328);
xnor U851 (N_851,In_1320,In_512);
nor U852 (N_852,In_942,In_869);
or U853 (N_853,In_799,In_127);
xor U854 (N_854,In_523,In_434);
and U855 (N_855,In_696,In_1153);
nand U856 (N_856,In_363,In_1468);
and U857 (N_857,In_1178,In_1479);
xnor U858 (N_858,In_1244,In_916);
nand U859 (N_859,In_650,In_1452);
or U860 (N_860,In_520,In_751);
xor U861 (N_861,In_236,In_659);
nand U862 (N_862,In_534,In_29);
nand U863 (N_863,In_242,In_1247);
xnor U864 (N_864,In_428,In_1208);
nor U865 (N_865,In_177,In_648);
nand U866 (N_866,In_1141,In_153);
xor U867 (N_867,In_623,In_1046);
xor U868 (N_868,In_85,In_1493);
xnor U869 (N_869,In_2,In_1272);
nor U870 (N_870,In_666,In_1244);
nand U871 (N_871,In_672,In_319);
and U872 (N_872,In_317,In_771);
nand U873 (N_873,In_584,In_25);
xnor U874 (N_874,In_56,In_730);
and U875 (N_875,In_1230,In_285);
and U876 (N_876,In_469,In_507);
nor U877 (N_877,In_645,In_1099);
or U878 (N_878,In_527,In_899);
nand U879 (N_879,In_149,In_1112);
xor U880 (N_880,In_364,In_205);
xnor U881 (N_881,In_654,In_296);
nand U882 (N_882,In_108,In_849);
nor U883 (N_883,In_286,In_1255);
nor U884 (N_884,In_1451,In_514);
nand U885 (N_885,In_1371,In_1355);
or U886 (N_886,In_941,In_185);
nand U887 (N_887,In_630,In_251);
nor U888 (N_888,In_516,In_897);
and U889 (N_889,In_582,In_1080);
and U890 (N_890,In_1092,In_130);
nand U891 (N_891,In_599,In_161);
xor U892 (N_892,In_206,In_535);
or U893 (N_893,In_80,In_525);
nor U894 (N_894,In_1305,In_545);
xnor U895 (N_895,In_1347,In_429);
nand U896 (N_896,In_1065,In_874);
nand U897 (N_897,In_84,In_10);
xnor U898 (N_898,In_1142,In_1450);
and U899 (N_899,In_1262,In_827);
or U900 (N_900,In_1280,In_1155);
or U901 (N_901,In_262,In_648);
nand U902 (N_902,In_319,In_238);
or U903 (N_903,In_446,In_1392);
and U904 (N_904,In_1243,In_532);
and U905 (N_905,In_270,In_615);
and U906 (N_906,In_117,In_369);
xor U907 (N_907,In_1202,In_951);
nand U908 (N_908,In_823,In_1198);
xor U909 (N_909,In_311,In_84);
nand U910 (N_910,In_1466,In_169);
xor U911 (N_911,In_583,In_81);
nand U912 (N_912,In_504,In_1068);
nor U913 (N_913,In_1431,In_841);
nand U914 (N_914,In_841,In_812);
nand U915 (N_915,In_1310,In_757);
nand U916 (N_916,In_763,In_26);
and U917 (N_917,In_40,In_1139);
xnor U918 (N_918,In_234,In_85);
and U919 (N_919,In_1231,In_1121);
xnor U920 (N_920,In_129,In_1428);
nor U921 (N_921,In_1485,In_620);
or U922 (N_922,In_1392,In_915);
nor U923 (N_923,In_1254,In_605);
xnor U924 (N_924,In_393,In_864);
xnor U925 (N_925,In_555,In_604);
and U926 (N_926,In_972,In_327);
and U927 (N_927,In_1494,In_1423);
nor U928 (N_928,In_1353,In_88);
and U929 (N_929,In_538,In_1080);
nor U930 (N_930,In_1253,In_280);
and U931 (N_931,In_394,In_1031);
nand U932 (N_932,In_1071,In_179);
nand U933 (N_933,In_74,In_507);
or U934 (N_934,In_1492,In_627);
nand U935 (N_935,In_137,In_418);
xor U936 (N_936,In_564,In_9);
and U937 (N_937,In_57,In_775);
nor U938 (N_938,In_1181,In_1050);
or U939 (N_939,In_15,In_1471);
nor U940 (N_940,In_696,In_142);
nand U941 (N_941,In_272,In_1447);
and U942 (N_942,In_304,In_682);
and U943 (N_943,In_386,In_1492);
xnor U944 (N_944,In_240,In_19);
xor U945 (N_945,In_1000,In_376);
or U946 (N_946,In_1228,In_358);
and U947 (N_947,In_1390,In_305);
nor U948 (N_948,In_857,In_730);
or U949 (N_949,In_277,In_181);
nand U950 (N_950,In_981,In_465);
and U951 (N_951,In_1340,In_100);
or U952 (N_952,In_437,In_812);
nor U953 (N_953,In_796,In_438);
xor U954 (N_954,In_109,In_826);
or U955 (N_955,In_648,In_509);
xnor U956 (N_956,In_1299,In_910);
nor U957 (N_957,In_983,In_1138);
nor U958 (N_958,In_1063,In_134);
nand U959 (N_959,In_587,In_1179);
nand U960 (N_960,In_238,In_330);
nand U961 (N_961,In_446,In_961);
xor U962 (N_962,In_162,In_1376);
xnor U963 (N_963,In_694,In_542);
and U964 (N_964,In_430,In_1313);
or U965 (N_965,In_678,In_318);
xor U966 (N_966,In_1267,In_1108);
nand U967 (N_967,In_1232,In_712);
nor U968 (N_968,In_225,In_323);
and U969 (N_969,In_1171,In_985);
and U970 (N_970,In_762,In_68);
or U971 (N_971,In_733,In_1089);
nand U972 (N_972,In_100,In_440);
xor U973 (N_973,In_806,In_699);
or U974 (N_974,In_1440,In_906);
xor U975 (N_975,In_491,In_373);
xor U976 (N_976,In_1000,In_185);
and U977 (N_977,In_970,In_951);
xor U978 (N_978,In_1260,In_914);
nand U979 (N_979,In_1405,In_1221);
and U980 (N_980,In_1365,In_1461);
xnor U981 (N_981,In_272,In_810);
and U982 (N_982,In_1196,In_988);
and U983 (N_983,In_55,In_798);
xor U984 (N_984,In_409,In_1267);
or U985 (N_985,In_1204,In_1420);
nand U986 (N_986,In_1045,In_1138);
nand U987 (N_987,In_50,In_1259);
and U988 (N_988,In_1367,In_342);
and U989 (N_989,In_304,In_256);
nand U990 (N_990,In_1315,In_313);
nor U991 (N_991,In_1205,In_778);
and U992 (N_992,In_1214,In_1395);
and U993 (N_993,In_1135,In_94);
xnor U994 (N_994,In_1385,In_627);
nor U995 (N_995,In_826,In_775);
nor U996 (N_996,In_132,In_771);
or U997 (N_997,In_1353,In_588);
nand U998 (N_998,In_1149,In_736);
or U999 (N_999,In_831,In_820);
xor U1000 (N_1000,In_930,In_140);
and U1001 (N_1001,In_23,In_1498);
and U1002 (N_1002,In_528,In_919);
xor U1003 (N_1003,In_861,In_1395);
and U1004 (N_1004,In_425,In_1188);
nor U1005 (N_1005,In_252,In_775);
nand U1006 (N_1006,In_939,In_209);
or U1007 (N_1007,In_1493,In_960);
or U1008 (N_1008,In_1101,In_484);
or U1009 (N_1009,In_880,In_1157);
xor U1010 (N_1010,In_372,In_1267);
xnor U1011 (N_1011,In_693,In_294);
xnor U1012 (N_1012,In_1256,In_547);
or U1013 (N_1013,In_1444,In_1416);
xor U1014 (N_1014,In_435,In_1423);
or U1015 (N_1015,In_477,In_492);
or U1016 (N_1016,In_1184,In_1412);
nand U1017 (N_1017,In_728,In_479);
and U1018 (N_1018,In_1246,In_1401);
or U1019 (N_1019,In_1378,In_314);
nand U1020 (N_1020,In_231,In_758);
xnor U1021 (N_1021,In_580,In_1261);
nor U1022 (N_1022,In_1190,In_1492);
nand U1023 (N_1023,In_1191,In_288);
or U1024 (N_1024,In_1055,In_477);
nand U1025 (N_1025,In_172,In_3);
nor U1026 (N_1026,In_724,In_153);
nand U1027 (N_1027,In_523,In_930);
and U1028 (N_1028,In_1302,In_1429);
xnor U1029 (N_1029,In_1071,In_588);
nand U1030 (N_1030,In_1270,In_199);
xor U1031 (N_1031,In_211,In_96);
xor U1032 (N_1032,In_652,In_345);
nand U1033 (N_1033,In_1200,In_280);
xnor U1034 (N_1034,In_1165,In_1321);
nor U1035 (N_1035,In_1417,In_934);
nor U1036 (N_1036,In_371,In_366);
or U1037 (N_1037,In_308,In_465);
nand U1038 (N_1038,In_584,In_1357);
and U1039 (N_1039,In_1375,In_653);
and U1040 (N_1040,In_969,In_831);
nor U1041 (N_1041,In_621,In_806);
xor U1042 (N_1042,In_1320,In_235);
xnor U1043 (N_1043,In_1036,In_1286);
nand U1044 (N_1044,In_1338,In_1429);
xnor U1045 (N_1045,In_1083,In_1153);
nor U1046 (N_1046,In_255,In_590);
xor U1047 (N_1047,In_714,In_5);
nand U1048 (N_1048,In_1349,In_1393);
nor U1049 (N_1049,In_489,In_1089);
and U1050 (N_1050,In_1265,In_1122);
nor U1051 (N_1051,In_946,In_981);
nand U1052 (N_1052,In_1267,In_422);
nor U1053 (N_1053,In_665,In_960);
nor U1054 (N_1054,In_688,In_1461);
nand U1055 (N_1055,In_1177,In_87);
nand U1056 (N_1056,In_924,In_295);
or U1057 (N_1057,In_368,In_1370);
nand U1058 (N_1058,In_294,In_750);
or U1059 (N_1059,In_1242,In_730);
xnor U1060 (N_1060,In_973,In_690);
and U1061 (N_1061,In_189,In_819);
xnor U1062 (N_1062,In_1108,In_1103);
xor U1063 (N_1063,In_325,In_1430);
and U1064 (N_1064,In_1378,In_59);
and U1065 (N_1065,In_1417,In_294);
or U1066 (N_1066,In_515,In_878);
and U1067 (N_1067,In_194,In_1070);
or U1068 (N_1068,In_1348,In_532);
and U1069 (N_1069,In_1018,In_673);
nand U1070 (N_1070,In_1222,In_696);
nand U1071 (N_1071,In_471,In_1125);
or U1072 (N_1072,In_549,In_947);
nand U1073 (N_1073,In_1096,In_688);
nor U1074 (N_1074,In_1068,In_630);
or U1075 (N_1075,In_1005,In_835);
nor U1076 (N_1076,In_920,In_1373);
nand U1077 (N_1077,In_224,In_1072);
xnor U1078 (N_1078,In_111,In_1412);
or U1079 (N_1079,In_1347,In_966);
xnor U1080 (N_1080,In_200,In_571);
nor U1081 (N_1081,In_941,In_681);
nor U1082 (N_1082,In_479,In_185);
xor U1083 (N_1083,In_935,In_887);
and U1084 (N_1084,In_1314,In_1400);
nor U1085 (N_1085,In_263,In_388);
nand U1086 (N_1086,In_225,In_1207);
nor U1087 (N_1087,In_107,In_1430);
or U1088 (N_1088,In_851,In_291);
nand U1089 (N_1089,In_292,In_1322);
or U1090 (N_1090,In_1174,In_488);
nand U1091 (N_1091,In_907,In_1275);
and U1092 (N_1092,In_1143,In_296);
nand U1093 (N_1093,In_1202,In_687);
or U1094 (N_1094,In_63,In_45);
xor U1095 (N_1095,In_1375,In_332);
nand U1096 (N_1096,In_339,In_598);
nand U1097 (N_1097,In_546,In_486);
nand U1098 (N_1098,In_308,In_385);
xnor U1099 (N_1099,In_150,In_311);
xor U1100 (N_1100,In_1484,In_383);
nor U1101 (N_1101,In_1222,In_192);
nand U1102 (N_1102,In_1,In_1053);
or U1103 (N_1103,In_1416,In_991);
nand U1104 (N_1104,In_1162,In_749);
nor U1105 (N_1105,In_1143,In_686);
and U1106 (N_1106,In_688,In_248);
xor U1107 (N_1107,In_164,In_369);
or U1108 (N_1108,In_992,In_718);
xnor U1109 (N_1109,In_387,In_1380);
xor U1110 (N_1110,In_631,In_203);
and U1111 (N_1111,In_523,In_225);
or U1112 (N_1112,In_607,In_362);
or U1113 (N_1113,In_1381,In_242);
xor U1114 (N_1114,In_859,In_170);
or U1115 (N_1115,In_463,In_486);
nand U1116 (N_1116,In_1315,In_649);
nor U1117 (N_1117,In_224,In_1355);
xnor U1118 (N_1118,In_733,In_301);
and U1119 (N_1119,In_1428,In_673);
xor U1120 (N_1120,In_980,In_775);
xor U1121 (N_1121,In_1075,In_399);
nor U1122 (N_1122,In_406,In_1004);
nand U1123 (N_1123,In_723,In_903);
nand U1124 (N_1124,In_1023,In_1391);
nand U1125 (N_1125,In_185,In_875);
xnor U1126 (N_1126,In_1459,In_552);
xor U1127 (N_1127,In_16,In_873);
nand U1128 (N_1128,In_238,In_410);
xnor U1129 (N_1129,In_1493,In_654);
or U1130 (N_1130,In_193,In_1416);
xor U1131 (N_1131,In_665,In_244);
nor U1132 (N_1132,In_872,In_1002);
nor U1133 (N_1133,In_537,In_1247);
nor U1134 (N_1134,In_824,In_187);
nand U1135 (N_1135,In_1072,In_328);
nand U1136 (N_1136,In_399,In_421);
nand U1137 (N_1137,In_1437,In_663);
xor U1138 (N_1138,In_1227,In_906);
nand U1139 (N_1139,In_451,In_790);
and U1140 (N_1140,In_1135,In_26);
or U1141 (N_1141,In_147,In_1399);
xor U1142 (N_1142,In_1289,In_983);
or U1143 (N_1143,In_830,In_1052);
nand U1144 (N_1144,In_1052,In_1084);
or U1145 (N_1145,In_1382,In_238);
or U1146 (N_1146,In_1350,In_91);
nor U1147 (N_1147,In_184,In_192);
nor U1148 (N_1148,In_1450,In_1079);
nor U1149 (N_1149,In_1323,In_1072);
nand U1150 (N_1150,In_340,In_641);
nand U1151 (N_1151,In_701,In_1365);
nand U1152 (N_1152,In_635,In_730);
nor U1153 (N_1153,In_981,In_1310);
and U1154 (N_1154,In_623,In_1371);
nand U1155 (N_1155,In_464,In_1096);
xnor U1156 (N_1156,In_1093,In_1037);
nor U1157 (N_1157,In_773,In_765);
and U1158 (N_1158,In_479,In_555);
and U1159 (N_1159,In_1104,In_177);
and U1160 (N_1160,In_1028,In_59);
or U1161 (N_1161,In_1110,In_188);
nand U1162 (N_1162,In_1416,In_820);
or U1163 (N_1163,In_147,In_623);
and U1164 (N_1164,In_309,In_1412);
and U1165 (N_1165,In_1120,In_1449);
and U1166 (N_1166,In_427,In_92);
xor U1167 (N_1167,In_191,In_355);
nand U1168 (N_1168,In_636,In_1142);
or U1169 (N_1169,In_598,In_192);
and U1170 (N_1170,In_1150,In_953);
nor U1171 (N_1171,In_124,In_1012);
or U1172 (N_1172,In_507,In_771);
nor U1173 (N_1173,In_175,In_170);
xor U1174 (N_1174,In_1357,In_1320);
nor U1175 (N_1175,In_1359,In_1462);
nor U1176 (N_1176,In_686,In_1408);
nor U1177 (N_1177,In_970,In_794);
and U1178 (N_1178,In_444,In_799);
or U1179 (N_1179,In_873,In_426);
or U1180 (N_1180,In_308,In_189);
xnor U1181 (N_1181,In_265,In_1160);
xor U1182 (N_1182,In_803,In_87);
or U1183 (N_1183,In_286,In_1358);
nand U1184 (N_1184,In_1015,In_984);
nand U1185 (N_1185,In_410,In_1498);
and U1186 (N_1186,In_908,In_729);
nor U1187 (N_1187,In_749,In_1263);
nand U1188 (N_1188,In_204,In_919);
nor U1189 (N_1189,In_112,In_838);
nand U1190 (N_1190,In_287,In_1205);
xor U1191 (N_1191,In_464,In_1025);
or U1192 (N_1192,In_1001,In_704);
or U1193 (N_1193,In_1411,In_429);
xor U1194 (N_1194,In_1220,In_409);
nand U1195 (N_1195,In_875,In_1103);
and U1196 (N_1196,In_880,In_31);
and U1197 (N_1197,In_912,In_1372);
or U1198 (N_1198,In_88,In_1271);
nor U1199 (N_1199,In_58,In_945);
xnor U1200 (N_1200,In_1229,In_447);
nor U1201 (N_1201,In_365,In_1165);
and U1202 (N_1202,In_515,In_742);
or U1203 (N_1203,In_351,In_851);
nand U1204 (N_1204,In_1011,In_62);
or U1205 (N_1205,In_455,In_257);
nand U1206 (N_1206,In_1214,In_613);
or U1207 (N_1207,In_785,In_192);
and U1208 (N_1208,In_457,In_1326);
nor U1209 (N_1209,In_224,In_756);
nand U1210 (N_1210,In_529,In_1000);
and U1211 (N_1211,In_971,In_1291);
or U1212 (N_1212,In_486,In_735);
or U1213 (N_1213,In_1231,In_1175);
xnor U1214 (N_1214,In_225,In_1028);
nor U1215 (N_1215,In_1256,In_748);
or U1216 (N_1216,In_1162,In_30);
or U1217 (N_1217,In_1417,In_1376);
xor U1218 (N_1218,In_777,In_1192);
xor U1219 (N_1219,In_846,In_630);
nand U1220 (N_1220,In_935,In_273);
nand U1221 (N_1221,In_1165,In_1120);
nor U1222 (N_1222,In_473,In_1267);
xor U1223 (N_1223,In_1103,In_955);
nor U1224 (N_1224,In_115,In_663);
nand U1225 (N_1225,In_1373,In_1343);
or U1226 (N_1226,In_916,In_190);
and U1227 (N_1227,In_35,In_581);
nor U1228 (N_1228,In_851,In_893);
xor U1229 (N_1229,In_1364,In_328);
nor U1230 (N_1230,In_476,In_1282);
xor U1231 (N_1231,In_1197,In_217);
and U1232 (N_1232,In_1454,In_799);
and U1233 (N_1233,In_1458,In_459);
nor U1234 (N_1234,In_183,In_1122);
and U1235 (N_1235,In_1157,In_1089);
nand U1236 (N_1236,In_228,In_25);
or U1237 (N_1237,In_265,In_453);
and U1238 (N_1238,In_372,In_367);
xnor U1239 (N_1239,In_322,In_942);
nand U1240 (N_1240,In_1329,In_578);
and U1241 (N_1241,In_822,In_502);
nand U1242 (N_1242,In_1273,In_597);
and U1243 (N_1243,In_1140,In_933);
nor U1244 (N_1244,In_1181,In_1105);
nand U1245 (N_1245,In_1452,In_889);
xor U1246 (N_1246,In_218,In_717);
nand U1247 (N_1247,In_592,In_398);
and U1248 (N_1248,In_434,In_352);
nor U1249 (N_1249,In_1022,In_1184);
nor U1250 (N_1250,In_20,In_1430);
and U1251 (N_1251,In_1298,In_1273);
or U1252 (N_1252,In_1302,In_1037);
nand U1253 (N_1253,In_1109,In_1222);
nand U1254 (N_1254,In_952,In_1187);
or U1255 (N_1255,In_810,In_417);
and U1256 (N_1256,In_336,In_509);
xnor U1257 (N_1257,In_51,In_361);
or U1258 (N_1258,In_595,In_1403);
nand U1259 (N_1259,In_542,In_777);
nand U1260 (N_1260,In_670,In_988);
nor U1261 (N_1261,In_835,In_1384);
nor U1262 (N_1262,In_280,In_412);
nand U1263 (N_1263,In_296,In_44);
nand U1264 (N_1264,In_515,In_368);
nand U1265 (N_1265,In_218,In_892);
nand U1266 (N_1266,In_499,In_711);
xor U1267 (N_1267,In_100,In_872);
nor U1268 (N_1268,In_1175,In_1061);
or U1269 (N_1269,In_1082,In_900);
and U1270 (N_1270,In_1240,In_1273);
xor U1271 (N_1271,In_479,In_1218);
xor U1272 (N_1272,In_365,In_1384);
xor U1273 (N_1273,In_1260,In_162);
or U1274 (N_1274,In_9,In_1195);
nor U1275 (N_1275,In_1344,In_913);
nor U1276 (N_1276,In_519,In_1127);
nand U1277 (N_1277,In_484,In_595);
nor U1278 (N_1278,In_271,In_1353);
nand U1279 (N_1279,In_1477,In_890);
xor U1280 (N_1280,In_596,In_1083);
and U1281 (N_1281,In_25,In_434);
nor U1282 (N_1282,In_496,In_1136);
and U1283 (N_1283,In_1425,In_1174);
or U1284 (N_1284,In_524,In_501);
and U1285 (N_1285,In_682,In_1486);
nor U1286 (N_1286,In_1462,In_673);
or U1287 (N_1287,In_487,In_1381);
or U1288 (N_1288,In_273,In_501);
and U1289 (N_1289,In_283,In_1212);
or U1290 (N_1290,In_1292,In_215);
nor U1291 (N_1291,In_292,In_838);
nand U1292 (N_1292,In_879,In_903);
or U1293 (N_1293,In_129,In_672);
nand U1294 (N_1294,In_1169,In_1496);
and U1295 (N_1295,In_1101,In_52);
nand U1296 (N_1296,In_345,In_238);
or U1297 (N_1297,In_483,In_218);
or U1298 (N_1298,In_521,In_36);
xnor U1299 (N_1299,In_1189,In_506);
or U1300 (N_1300,In_1413,In_1128);
or U1301 (N_1301,In_427,In_924);
and U1302 (N_1302,In_762,In_1105);
and U1303 (N_1303,In_892,In_579);
or U1304 (N_1304,In_1398,In_891);
and U1305 (N_1305,In_889,In_676);
nor U1306 (N_1306,In_1466,In_1087);
xnor U1307 (N_1307,In_1148,In_1279);
and U1308 (N_1308,In_21,In_1060);
and U1309 (N_1309,In_958,In_570);
nor U1310 (N_1310,In_492,In_410);
xnor U1311 (N_1311,In_1369,In_1109);
or U1312 (N_1312,In_928,In_1490);
nand U1313 (N_1313,In_1474,In_275);
nor U1314 (N_1314,In_1332,In_881);
or U1315 (N_1315,In_1224,In_859);
or U1316 (N_1316,In_249,In_384);
and U1317 (N_1317,In_106,In_841);
nand U1318 (N_1318,In_306,In_1288);
xnor U1319 (N_1319,In_244,In_316);
and U1320 (N_1320,In_779,In_1423);
and U1321 (N_1321,In_287,In_1254);
xor U1322 (N_1322,In_1003,In_781);
and U1323 (N_1323,In_1006,In_292);
and U1324 (N_1324,In_533,In_413);
xor U1325 (N_1325,In_203,In_1002);
xor U1326 (N_1326,In_22,In_1441);
xnor U1327 (N_1327,In_350,In_1026);
nor U1328 (N_1328,In_141,In_621);
or U1329 (N_1329,In_839,In_198);
or U1330 (N_1330,In_467,In_794);
nand U1331 (N_1331,In_40,In_1345);
nor U1332 (N_1332,In_359,In_201);
nor U1333 (N_1333,In_719,In_1155);
nand U1334 (N_1334,In_998,In_1130);
xor U1335 (N_1335,In_250,In_918);
nand U1336 (N_1336,In_16,In_1317);
nor U1337 (N_1337,In_119,In_597);
xor U1338 (N_1338,In_61,In_116);
xnor U1339 (N_1339,In_417,In_1316);
nand U1340 (N_1340,In_1338,In_115);
and U1341 (N_1341,In_152,In_862);
and U1342 (N_1342,In_1198,In_526);
nand U1343 (N_1343,In_874,In_188);
or U1344 (N_1344,In_329,In_845);
nand U1345 (N_1345,In_1279,In_1301);
or U1346 (N_1346,In_807,In_1255);
nor U1347 (N_1347,In_1218,In_730);
and U1348 (N_1348,In_674,In_918);
and U1349 (N_1349,In_776,In_470);
and U1350 (N_1350,In_842,In_391);
nand U1351 (N_1351,In_605,In_763);
and U1352 (N_1352,In_74,In_182);
or U1353 (N_1353,In_117,In_1283);
xor U1354 (N_1354,In_1290,In_263);
nand U1355 (N_1355,In_1185,In_54);
and U1356 (N_1356,In_331,In_787);
nand U1357 (N_1357,In_612,In_1069);
and U1358 (N_1358,In_106,In_40);
and U1359 (N_1359,In_114,In_283);
nor U1360 (N_1360,In_504,In_334);
and U1361 (N_1361,In_335,In_1458);
nor U1362 (N_1362,In_860,In_998);
or U1363 (N_1363,In_933,In_156);
and U1364 (N_1364,In_37,In_261);
and U1365 (N_1365,In_1391,In_1308);
nand U1366 (N_1366,In_132,In_264);
nor U1367 (N_1367,In_324,In_738);
xor U1368 (N_1368,In_1029,In_1498);
or U1369 (N_1369,In_967,In_276);
nor U1370 (N_1370,In_1006,In_1083);
nor U1371 (N_1371,In_431,In_6);
or U1372 (N_1372,In_872,In_86);
nor U1373 (N_1373,In_194,In_1243);
or U1374 (N_1374,In_1141,In_36);
or U1375 (N_1375,In_399,In_1318);
or U1376 (N_1376,In_1169,In_1480);
nor U1377 (N_1377,In_600,In_1303);
xnor U1378 (N_1378,In_1215,In_1417);
or U1379 (N_1379,In_285,In_390);
or U1380 (N_1380,In_758,In_1469);
and U1381 (N_1381,In_841,In_58);
nand U1382 (N_1382,In_891,In_482);
xor U1383 (N_1383,In_649,In_926);
or U1384 (N_1384,In_761,In_267);
nor U1385 (N_1385,In_1455,In_373);
nand U1386 (N_1386,In_997,In_287);
xnor U1387 (N_1387,In_115,In_270);
xor U1388 (N_1388,In_851,In_1183);
nor U1389 (N_1389,In_241,In_351);
nand U1390 (N_1390,In_1233,In_355);
and U1391 (N_1391,In_1049,In_902);
nor U1392 (N_1392,In_1378,In_666);
and U1393 (N_1393,In_860,In_1497);
or U1394 (N_1394,In_1119,In_1367);
nand U1395 (N_1395,In_1064,In_995);
nor U1396 (N_1396,In_299,In_553);
or U1397 (N_1397,In_1338,In_1375);
or U1398 (N_1398,In_585,In_312);
xor U1399 (N_1399,In_10,In_236);
and U1400 (N_1400,In_1253,In_1107);
nor U1401 (N_1401,In_819,In_1212);
nand U1402 (N_1402,In_1485,In_533);
nor U1403 (N_1403,In_1383,In_473);
or U1404 (N_1404,In_891,In_1417);
xor U1405 (N_1405,In_15,In_733);
and U1406 (N_1406,In_548,In_1007);
or U1407 (N_1407,In_318,In_1307);
and U1408 (N_1408,In_1489,In_1063);
nand U1409 (N_1409,In_322,In_1055);
and U1410 (N_1410,In_930,In_1474);
nor U1411 (N_1411,In_1292,In_120);
xnor U1412 (N_1412,In_484,In_115);
nor U1413 (N_1413,In_336,In_742);
nand U1414 (N_1414,In_697,In_325);
xnor U1415 (N_1415,In_425,In_359);
xor U1416 (N_1416,In_212,In_248);
or U1417 (N_1417,In_1009,In_1230);
or U1418 (N_1418,In_455,In_388);
nor U1419 (N_1419,In_1146,In_86);
nor U1420 (N_1420,In_213,In_707);
nor U1421 (N_1421,In_937,In_620);
xnor U1422 (N_1422,In_424,In_153);
nand U1423 (N_1423,In_1035,In_1049);
and U1424 (N_1424,In_1355,In_25);
nand U1425 (N_1425,In_1036,In_524);
xnor U1426 (N_1426,In_1116,In_1436);
or U1427 (N_1427,In_220,In_1396);
nand U1428 (N_1428,In_1116,In_1308);
xnor U1429 (N_1429,In_190,In_1420);
and U1430 (N_1430,In_91,In_702);
and U1431 (N_1431,In_1472,In_743);
nor U1432 (N_1432,In_719,In_539);
or U1433 (N_1433,In_1269,In_1069);
nor U1434 (N_1434,In_664,In_693);
or U1435 (N_1435,In_779,In_184);
nand U1436 (N_1436,In_1287,In_845);
nand U1437 (N_1437,In_695,In_1064);
nor U1438 (N_1438,In_1223,In_1096);
nor U1439 (N_1439,In_639,In_308);
nand U1440 (N_1440,In_1371,In_1395);
and U1441 (N_1441,In_1200,In_600);
or U1442 (N_1442,In_1075,In_1395);
nand U1443 (N_1443,In_431,In_89);
or U1444 (N_1444,In_1281,In_1228);
or U1445 (N_1445,In_1481,In_1242);
nor U1446 (N_1446,In_300,In_464);
and U1447 (N_1447,In_969,In_534);
nor U1448 (N_1448,In_634,In_438);
nor U1449 (N_1449,In_1490,In_356);
nand U1450 (N_1450,In_21,In_608);
xor U1451 (N_1451,In_208,In_1474);
nand U1452 (N_1452,In_1162,In_233);
and U1453 (N_1453,In_24,In_899);
nand U1454 (N_1454,In_385,In_1199);
nand U1455 (N_1455,In_1233,In_838);
and U1456 (N_1456,In_445,In_1398);
nor U1457 (N_1457,In_1475,In_1497);
nand U1458 (N_1458,In_177,In_1293);
xor U1459 (N_1459,In_690,In_571);
nand U1460 (N_1460,In_258,In_430);
nand U1461 (N_1461,In_1227,In_664);
xnor U1462 (N_1462,In_1362,In_1405);
nand U1463 (N_1463,In_451,In_1295);
nor U1464 (N_1464,In_973,In_660);
and U1465 (N_1465,In_729,In_1271);
nand U1466 (N_1466,In_165,In_662);
and U1467 (N_1467,In_288,In_1193);
or U1468 (N_1468,In_183,In_1330);
nand U1469 (N_1469,In_57,In_1034);
nand U1470 (N_1470,In_1198,In_1218);
nor U1471 (N_1471,In_518,In_487);
or U1472 (N_1472,In_930,In_116);
or U1473 (N_1473,In_362,In_196);
xnor U1474 (N_1474,In_590,In_790);
xor U1475 (N_1475,In_94,In_751);
xnor U1476 (N_1476,In_907,In_771);
or U1477 (N_1477,In_357,In_1240);
nor U1478 (N_1478,In_919,In_420);
or U1479 (N_1479,In_1279,In_537);
or U1480 (N_1480,In_793,In_769);
or U1481 (N_1481,In_70,In_988);
xor U1482 (N_1482,In_135,In_225);
nand U1483 (N_1483,In_659,In_230);
xnor U1484 (N_1484,In_1493,In_1220);
xnor U1485 (N_1485,In_695,In_560);
nor U1486 (N_1486,In_939,In_565);
nand U1487 (N_1487,In_166,In_447);
nand U1488 (N_1488,In_193,In_6);
nor U1489 (N_1489,In_1200,In_1429);
xor U1490 (N_1490,In_1261,In_1230);
nor U1491 (N_1491,In_151,In_333);
or U1492 (N_1492,In_484,In_1464);
or U1493 (N_1493,In_1366,In_906);
nand U1494 (N_1494,In_1264,In_944);
nor U1495 (N_1495,In_888,In_1428);
and U1496 (N_1496,In_37,In_167);
and U1497 (N_1497,In_281,In_928);
and U1498 (N_1498,In_704,In_426);
nor U1499 (N_1499,In_982,In_1119);
xnor U1500 (N_1500,In_891,In_369);
xor U1501 (N_1501,In_554,In_1033);
nor U1502 (N_1502,In_658,In_786);
and U1503 (N_1503,In_1167,In_1499);
and U1504 (N_1504,In_294,In_181);
nand U1505 (N_1505,In_567,In_245);
xnor U1506 (N_1506,In_547,In_755);
and U1507 (N_1507,In_1246,In_1422);
xor U1508 (N_1508,In_1321,In_92);
and U1509 (N_1509,In_1470,In_161);
xor U1510 (N_1510,In_1381,In_691);
nand U1511 (N_1511,In_668,In_1290);
and U1512 (N_1512,In_842,In_1151);
nor U1513 (N_1513,In_1228,In_346);
or U1514 (N_1514,In_950,In_710);
nor U1515 (N_1515,In_1456,In_1020);
and U1516 (N_1516,In_1181,In_295);
xor U1517 (N_1517,In_48,In_694);
xnor U1518 (N_1518,In_147,In_721);
or U1519 (N_1519,In_646,In_805);
and U1520 (N_1520,In_376,In_805);
or U1521 (N_1521,In_331,In_605);
or U1522 (N_1522,In_1065,In_1443);
xnor U1523 (N_1523,In_88,In_56);
and U1524 (N_1524,In_1477,In_618);
and U1525 (N_1525,In_1274,In_296);
and U1526 (N_1526,In_1083,In_870);
nand U1527 (N_1527,In_493,In_178);
nor U1528 (N_1528,In_1100,In_500);
nand U1529 (N_1529,In_125,In_1092);
xor U1530 (N_1530,In_997,In_685);
xnor U1531 (N_1531,In_374,In_241);
nor U1532 (N_1532,In_1387,In_586);
xnor U1533 (N_1533,In_155,In_248);
xor U1534 (N_1534,In_70,In_561);
nand U1535 (N_1535,In_995,In_1387);
or U1536 (N_1536,In_620,In_1251);
nand U1537 (N_1537,In_318,In_717);
and U1538 (N_1538,In_2,In_423);
xor U1539 (N_1539,In_983,In_55);
and U1540 (N_1540,In_518,In_732);
or U1541 (N_1541,In_1130,In_1430);
nand U1542 (N_1542,In_1010,In_480);
xnor U1543 (N_1543,In_788,In_1271);
and U1544 (N_1544,In_106,In_1221);
nor U1545 (N_1545,In_387,In_593);
xor U1546 (N_1546,In_682,In_1390);
xnor U1547 (N_1547,In_1305,In_1410);
xnor U1548 (N_1548,In_348,In_809);
xor U1549 (N_1549,In_412,In_362);
nand U1550 (N_1550,In_1224,In_124);
and U1551 (N_1551,In_100,In_29);
xor U1552 (N_1552,In_1283,In_889);
and U1553 (N_1553,In_1090,In_1181);
xor U1554 (N_1554,In_1193,In_1421);
nand U1555 (N_1555,In_1055,In_1038);
nand U1556 (N_1556,In_817,In_978);
and U1557 (N_1557,In_1257,In_1297);
and U1558 (N_1558,In_1233,In_583);
xnor U1559 (N_1559,In_1064,In_239);
or U1560 (N_1560,In_549,In_177);
xnor U1561 (N_1561,In_646,In_346);
xnor U1562 (N_1562,In_1378,In_1420);
nand U1563 (N_1563,In_1389,In_50);
nand U1564 (N_1564,In_1384,In_433);
or U1565 (N_1565,In_1112,In_292);
xnor U1566 (N_1566,In_483,In_1406);
xor U1567 (N_1567,In_1282,In_1000);
and U1568 (N_1568,In_231,In_1155);
nand U1569 (N_1569,In_184,In_1476);
xor U1570 (N_1570,In_181,In_1152);
nor U1571 (N_1571,In_1246,In_196);
nor U1572 (N_1572,In_636,In_1202);
nor U1573 (N_1573,In_298,In_305);
xor U1574 (N_1574,In_563,In_134);
nor U1575 (N_1575,In_984,In_1324);
nor U1576 (N_1576,In_195,In_84);
nor U1577 (N_1577,In_832,In_944);
nor U1578 (N_1578,In_1055,In_1268);
and U1579 (N_1579,In_1218,In_871);
xor U1580 (N_1580,In_1471,In_434);
nand U1581 (N_1581,In_813,In_137);
nor U1582 (N_1582,In_558,In_524);
xnor U1583 (N_1583,In_1132,In_624);
and U1584 (N_1584,In_236,In_419);
or U1585 (N_1585,In_1163,In_920);
xor U1586 (N_1586,In_1287,In_1375);
and U1587 (N_1587,In_677,In_1030);
nand U1588 (N_1588,In_766,In_264);
xnor U1589 (N_1589,In_1156,In_884);
nand U1590 (N_1590,In_294,In_597);
nor U1591 (N_1591,In_1424,In_182);
nor U1592 (N_1592,In_1390,In_810);
and U1593 (N_1593,In_261,In_607);
nor U1594 (N_1594,In_195,In_1468);
xnor U1595 (N_1595,In_169,In_2);
nand U1596 (N_1596,In_1464,In_327);
xor U1597 (N_1597,In_821,In_638);
nand U1598 (N_1598,In_247,In_372);
or U1599 (N_1599,In_1166,In_911);
xor U1600 (N_1600,In_1226,In_606);
and U1601 (N_1601,In_380,In_940);
and U1602 (N_1602,In_534,In_994);
and U1603 (N_1603,In_285,In_738);
or U1604 (N_1604,In_1006,In_475);
nand U1605 (N_1605,In_1035,In_380);
nand U1606 (N_1606,In_738,In_96);
xor U1607 (N_1607,In_71,In_655);
nor U1608 (N_1608,In_1351,In_84);
xnor U1609 (N_1609,In_296,In_1123);
xnor U1610 (N_1610,In_918,In_874);
nand U1611 (N_1611,In_51,In_1183);
and U1612 (N_1612,In_773,In_1057);
nand U1613 (N_1613,In_248,In_1400);
xor U1614 (N_1614,In_1159,In_536);
nand U1615 (N_1615,In_129,In_569);
and U1616 (N_1616,In_1343,In_869);
and U1617 (N_1617,In_1152,In_1091);
or U1618 (N_1618,In_165,In_1417);
or U1619 (N_1619,In_1255,In_768);
or U1620 (N_1620,In_1069,In_1228);
and U1621 (N_1621,In_577,In_586);
or U1622 (N_1622,In_0,In_85);
xor U1623 (N_1623,In_984,In_1468);
xor U1624 (N_1624,In_492,In_522);
nand U1625 (N_1625,In_1366,In_803);
and U1626 (N_1626,In_1445,In_614);
xnor U1627 (N_1627,In_733,In_1219);
xor U1628 (N_1628,In_499,In_574);
or U1629 (N_1629,In_235,In_196);
or U1630 (N_1630,In_1054,In_734);
xnor U1631 (N_1631,In_899,In_1055);
nand U1632 (N_1632,In_1092,In_493);
xor U1633 (N_1633,In_648,In_1298);
xnor U1634 (N_1634,In_98,In_1192);
or U1635 (N_1635,In_658,In_160);
nand U1636 (N_1636,In_123,In_692);
xor U1637 (N_1637,In_492,In_1014);
nor U1638 (N_1638,In_153,In_902);
nand U1639 (N_1639,In_548,In_639);
nor U1640 (N_1640,In_990,In_816);
and U1641 (N_1641,In_1336,In_749);
xnor U1642 (N_1642,In_752,In_600);
or U1643 (N_1643,In_118,In_799);
and U1644 (N_1644,In_610,In_1039);
nor U1645 (N_1645,In_1435,In_441);
and U1646 (N_1646,In_5,In_1184);
xor U1647 (N_1647,In_864,In_849);
nor U1648 (N_1648,In_344,In_531);
and U1649 (N_1649,In_1495,In_1097);
nor U1650 (N_1650,In_663,In_289);
and U1651 (N_1651,In_1291,In_1421);
and U1652 (N_1652,In_710,In_1253);
and U1653 (N_1653,In_1072,In_458);
nor U1654 (N_1654,In_1022,In_199);
nor U1655 (N_1655,In_1134,In_115);
nand U1656 (N_1656,In_1214,In_164);
or U1657 (N_1657,In_408,In_413);
nor U1658 (N_1658,In_85,In_1113);
xor U1659 (N_1659,In_830,In_1351);
nor U1660 (N_1660,In_1298,In_294);
xnor U1661 (N_1661,In_824,In_531);
nor U1662 (N_1662,In_787,In_1375);
or U1663 (N_1663,In_1256,In_1341);
nor U1664 (N_1664,In_32,In_498);
nor U1665 (N_1665,In_559,In_1434);
and U1666 (N_1666,In_322,In_379);
nor U1667 (N_1667,In_1410,In_705);
nand U1668 (N_1668,In_1174,In_384);
nand U1669 (N_1669,In_897,In_211);
or U1670 (N_1670,In_1242,In_1354);
nor U1671 (N_1671,In_259,In_11);
and U1672 (N_1672,In_950,In_451);
or U1673 (N_1673,In_1330,In_714);
nor U1674 (N_1674,In_1237,In_610);
xor U1675 (N_1675,In_827,In_540);
nor U1676 (N_1676,In_430,In_1192);
nand U1677 (N_1677,In_686,In_587);
xnor U1678 (N_1678,In_1102,In_130);
nor U1679 (N_1679,In_13,In_1022);
nor U1680 (N_1680,In_1233,In_449);
or U1681 (N_1681,In_1414,In_891);
nor U1682 (N_1682,In_42,In_782);
and U1683 (N_1683,In_170,In_1083);
xor U1684 (N_1684,In_286,In_502);
and U1685 (N_1685,In_470,In_879);
or U1686 (N_1686,In_126,In_612);
nand U1687 (N_1687,In_790,In_746);
nor U1688 (N_1688,In_1204,In_1442);
nor U1689 (N_1689,In_678,In_809);
xnor U1690 (N_1690,In_42,In_1411);
nor U1691 (N_1691,In_75,In_477);
xor U1692 (N_1692,In_94,In_748);
nand U1693 (N_1693,In_584,In_616);
or U1694 (N_1694,In_849,In_567);
and U1695 (N_1695,In_1079,In_883);
nor U1696 (N_1696,In_380,In_628);
or U1697 (N_1697,In_1482,In_587);
nor U1698 (N_1698,In_340,In_36);
nand U1699 (N_1699,In_490,In_1386);
nand U1700 (N_1700,In_554,In_985);
xor U1701 (N_1701,In_1062,In_1273);
nor U1702 (N_1702,In_130,In_1019);
xnor U1703 (N_1703,In_157,In_285);
xnor U1704 (N_1704,In_1089,In_59);
or U1705 (N_1705,In_329,In_1330);
and U1706 (N_1706,In_946,In_291);
xor U1707 (N_1707,In_95,In_1353);
and U1708 (N_1708,In_992,In_1449);
nor U1709 (N_1709,In_307,In_319);
or U1710 (N_1710,In_1478,In_267);
nor U1711 (N_1711,In_987,In_610);
nor U1712 (N_1712,In_782,In_910);
xnor U1713 (N_1713,In_1200,In_1395);
nand U1714 (N_1714,In_132,In_1319);
xor U1715 (N_1715,In_905,In_715);
nor U1716 (N_1716,In_133,In_1413);
or U1717 (N_1717,In_1456,In_493);
nand U1718 (N_1718,In_891,In_745);
or U1719 (N_1719,In_461,In_624);
xor U1720 (N_1720,In_1031,In_28);
or U1721 (N_1721,In_473,In_907);
nor U1722 (N_1722,In_1304,In_1449);
and U1723 (N_1723,In_11,In_110);
or U1724 (N_1724,In_1159,In_1184);
xnor U1725 (N_1725,In_616,In_697);
and U1726 (N_1726,In_476,In_112);
nand U1727 (N_1727,In_561,In_1076);
xnor U1728 (N_1728,In_654,In_1357);
nor U1729 (N_1729,In_190,In_1424);
nand U1730 (N_1730,In_852,In_160);
and U1731 (N_1731,In_1391,In_102);
and U1732 (N_1732,In_334,In_733);
or U1733 (N_1733,In_84,In_593);
xnor U1734 (N_1734,In_1453,In_103);
and U1735 (N_1735,In_155,In_1210);
nor U1736 (N_1736,In_686,In_1436);
or U1737 (N_1737,In_845,In_1304);
and U1738 (N_1738,In_1198,In_128);
or U1739 (N_1739,In_677,In_31);
nand U1740 (N_1740,In_1184,In_742);
nor U1741 (N_1741,In_1313,In_1074);
or U1742 (N_1742,In_499,In_1267);
and U1743 (N_1743,In_176,In_1357);
and U1744 (N_1744,In_1292,In_1359);
nor U1745 (N_1745,In_905,In_81);
or U1746 (N_1746,In_845,In_148);
nor U1747 (N_1747,In_933,In_1307);
and U1748 (N_1748,In_1149,In_504);
nand U1749 (N_1749,In_1094,In_713);
xnor U1750 (N_1750,In_1337,In_33);
and U1751 (N_1751,In_830,In_1492);
and U1752 (N_1752,In_1097,In_1464);
or U1753 (N_1753,In_41,In_1118);
or U1754 (N_1754,In_774,In_1230);
or U1755 (N_1755,In_498,In_1087);
or U1756 (N_1756,In_555,In_1226);
nor U1757 (N_1757,In_53,In_1033);
and U1758 (N_1758,In_735,In_446);
nor U1759 (N_1759,In_197,In_1436);
xnor U1760 (N_1760,In_437,In_1233);
nand U1761 (N_1761,In_1498,In_156);
xnor U1762 (N_1762,In_943,In_150);
or U1763 (N_1763,In_709,In_1105);
or U1764 (N_1764,In_1452,In_878);
nor U1765 (N_1765,In_1105,In_1079);
nor U1766 (N_1766,In_362,In_693);
nand U1767 (N_1767,In_1017,In_818);
xnor U1768 (N_1768,In_1190,In_946);
nor U1769 (N_1769,In_287,In_259);
nor U1770 (N_1770,In_1203,In_892);
or U1771 (N_1771,In_430,In_292);
xor U1772 (N_1772,In_1058,In_1422);
or U1773 (N_1773,In_1319,In_1128);
xor U1774 (N_1774,In_1145,In_1406);
xor U1775 (N_1775,In_1385,In_724);
or U1776 (N_1776,In_426,In_29);
nand U1777 (N_1777,In_917,In_937);
nand U1778 (N_1778,In_448,In_626);
or U1779 (N_1779,In_1431,In_418);
nand U1780 (N_1780,In_134,In_1082);
nor U1781 (N_1781,In_1336,In_1123);
nor U1782 (N_1782,In_1331,In_1386);
nand U1783 (N_1783,In_678,In_372);
and U1784 (N_1784,In_103,In_1385);
nand U1785 (N_1785,In_665,In_1114);
and U1786 (N_1786,In_753,In_1056);
and U1787 (N_1787,In_1451,In_127);
xnor U1788 (N_1788,In_480,In_1280);
or U1789 (N_1789,In_246,In_86);
nor U1790 (N_1790,In_128,In_1115);
and U1791 (N_1791,In_986,In_1149);
or U1792 (N_1792,In_823,In_580);
or U1793 (N_1793,In_836,In_368);
nand U1794 (N_1794,In_77,In_930);
or U1795 (N_1795,In_432,In_292);
xnor U1796 (N_1796,In_104,In_929);
or U1797 (N_1797,In_181,In_360);
nor U1798 (N_1798,In_1416,In_254);
and U1799 (N_1799,In_701,In_1414);
nor U1800 (N_1800,In_1133,In_898);
and U1801 (N_1801,In_129,In_1169);
nor U1802 (N_1802,In_1110,In_332);
nand U1803 (N_1803,In_358,In_1356);
or U1804 (N_1804,In_1394,In_1490);
or U1805 (N_1805,In_65,In_947);
xnor U1806 (N_1806,In_271,In_266);
xnor U1807 (N_1807,In_1462,In_1279);
nand U1808 (N_1808,In_50,In_105);
xor U1809 (N_1809,In_348,In_40);
nor U1810 (N_1810,In_569,In_476);
or U1811 (N_1811,In_459,In_245);
or U1812 (N_1812,In_196,In_298);
nor U1813 (N_1813,In_146,In_156);
or U1814 (N_1814,In_1442,In_1452);
nor U1815 (N_1815,In_1037,In_27);
xnor U1816 (N_1816,In_888,In_360);
and U1817 (N_1817,In_1444,In_717);
nand U1818 (N_1818,In_1485,In_1245);
nor U1819 (N_1819,In_607,In_967);
xor U1820 (N_1820,In_1091,In_1081);
xor U1821 (N_1821,In_1495,In_1485);
xnor U1822 (N_1822,In_1274,In_894);
xor U1823 (N_1823,In_255,In_1349);
nor U1824 (N_1824,In_1450,In_517);
nor U1825 (N_1825,In_344,In_735);
nor U1826 (N_1826,In_541,In_555);
nor U1827 (N_1827,In_175,In_340);
nand U1828 (N_1828,In_131,In_76);
xor U1829 (N_1829,In_615,In_1433);
or U1830 (N_1830,In_1262,In_1086);
or U1831 (N_1831,In_951,In_270);
nor U1832 (N_1832,In_1027,In_1060);
nand U1833 (N_1833,In_62,In_1357);
or U1834 (N_1834,In_416,In_19);
nor U1835 (N_1835,In_548,In_63);
or U1836 (N_1836,In_404,In_1493);
and U1837 (N_1837,In_1328,In_45);
and U1838 (N_1838,In_985,In_174);
nand U1839 (N_1839,In_1466,In_477);
nand U1840 (N_1840,In_322,In_1003);
and U1841 (N_1841,In_559,In_710);
nor U1842 (N_1842,In_685,In_1034);
and U1843 (N_1843,In_322,In_451);
nand U1844 (N_1844,In_1170,In_818);
and U1845 (N_1845,In_930,In_999);
and U1846 (N_1846,In_1483,In_550);
xnor U1847 (N_1847,In_1370,In_1042);
xnor U1848 (N_1848,In_1116,In_262);
and U1849 (N_1849,In_598,In_264);
or U1850 (N_1850,In_1381,In_611);
xor U1851 (N_1851,In_1263,In_1220);
xor U1852 (N_1852,In_1222,In_1499);
or U1853 (N_1853,In_1153,In_387);
nor U1854 (N_1854,In_211,In_18);
and U1855 (N_1855,In_900,In_1106);
or U1856 (N_1856,In_182,In_420);
nor U1857 (N_1857,In_691,In_1330);
or U1858 (N_1858,In_856,In_138);
nor U1859 (N_1859,In_355,In_1241);
or U1860 (N_1860,In_173,In_506);
xor U1861 (N_1861,In_1216,In_1282);
and U1862 (N_1862,In_41,In_611);
nor U1863 (N_1863,In_1406,In_731);
nor U1864 (N_1864,In_62,In_1115);
nor U1865 (N_1865,In_457,In_935);
xnor U1866 (N_1866,In_592,In_424);
nor U1867 (N_1867,In_680,In_699);
nor U1868 (N_1868,In_89,In_524);
nand U1869 (N_1869,In_987,In_1299);
nor U1870 (N_1870,In_36,In_1361);
or U1871 (N_1871,In_129,In_1213);
xor U1872 (N_1872,In_1206,In_645);
nand U1873 (N_1873,In_79,In_981);
nand U1874 (N_1874,In_562,In_298);
xor U1875 (N_1875,In_961,In_1477);
nor U1876 (N_1876,In_647,In_1068);
and U1877 (N_1877,In_461,In_1076);
and U1878 (N_1878,In_1287,In_941);
and U1879 (N_1879,In_1268,In_558);
nor U1880 (N_1880,In_441,In_577);
and U1881 (N_1881,In_551,In_157);
nand U1882 (N_1882,In_88,In_245);
xnor U1883 (N_1883,In_717,In_1318);
and U1884 (N_1884,In_1371,In_79);
nand U1885 (N_1885,In_460,In_291);
nor U1886 (N_1886,In_137,In_380);
nor U1887 (N_1887,In_668,In_319);
nand U1888 (N_1888,In_83,In_526);
and U1889 (N_1889,In_194,In_1060);
or U1890 (N_1890,In_930,In_47);
or U1891 (N_1891,In_1282,In_643);
xor U1892 (N_1892,In_160,In_1181);
or U1893 (N_1893,In_960,In_660);
xor U1894 (N_1894,In_1458,In_1351);
and U1895 (N_1895,In_250,In_178);
and U1896 (N_1896,In_605,In_321);
xor U1897 (N_1897,In_196,In_70);
xor U1898 (N_1898,In_104,In_1188);
nand U1899 (N_1899,In_60,In_831);
nand U1900 (N_1900,In_403,In_491);
or U1901 (N_1901,In_883,In_30);
or U1902 (N_1902,In_109,In_740);
and U1903 (N_1903,In_430,In_336);
xor U1904 (N_1904,In_305,In_842);
xnor U1905 (N_1905,In_539,In_58);
xor U1906 (N_1906,In_34,In_915);
nor U1907 (N_1907,In_23,In_1082);
xor U1908 (N_1908,In_1220,In_491);
nor U1909 (N_1909,In_286,In_1047);
or U1910 (N_1910,In_574,In_1293);
nor U1911 (N_1911,In_843,In_1011);
nand U1912 (N_1912,In_834,In_461);
and U1913 (N_1913,In_124,In_830);
nor U1914 (N_1914,In_1144,In_623);
and U1915 (N_1915,In_531,In_741);
nor U1916 (N_1916,In_1273,In_1274);
nor U1917 (N_1917,In_713,In_749);
or U1918 (N_1918,In_1255,In_267);
or U1919 (N_1919,In_1298,In_1417);
xor U1920 (N_1920,In_869,In_1311);
nor U1921 (N_1921,In_114,In_55);
and U1922 (N_1922,In_1077,In_1409);
and U1923 (N_1923,In_17,In_1325);
and U1924 (N_1924,In_1410,In_1217);
xnor U1925 (N_1925,In_222,In_568);
nor U1926 (N_1926,In_1149,In_1167);
and U1927 (N_1927,In_1051,In_171);
nor U1928 (N_1928,In_1216,In_1127);
or U1929 (N_1929,In_209,In_494);
nor U1930 (N_1930,In_165,In_283);
or U1931 (N_1931,In_923,In_1156);
and U1932 (N_1932,In_928,In_820);
and U1933 (N_1933,In_136,In_1168);
nor U1934 (N_1934,In_1084,In_803);
or U1935 (N_1935,In_673,In_1193);
xnor U1936 (N_1936,In_867,In_102);
nor U1937 (N_1937,In_645,In_1471);
nand U1938 (N_1938,In_180,In_1218);
xnor U1939 (N_1939,In_889,In_67);
xor U1940 (N_1940,In_1198,In_111);
and U1941 (N_1941,In_39,In_1213);
nor U1942 (N_1942,In_557,In_1134);
xnor U1943 (N_1943,In_1219,In_326);
nor U1944 (N_1944,In_6,In_1254);
nand U1945 (N_1945,In_681,In_335);
xnor U1946 (N_1946,In_345,In_671);
or U1947 (N_1947,In_824,In_685);
nand U1948 (N_1948,In_1489,In_228);
xnor U1949 (N_1949,In_248,In_1130);
nand U1950 (N_1950,In_1046,In_586);
xor U1951 (N_1951,In_942,In_1112);
and U1952 (N_1952,In_238,In_1495);
or U1953 (N_1953,In_238,In_567);
and U1954 (N_1954,In_361,In_1301);
xor U1955 (N_1955,In_1102,In_206);
or U1956 (N_1956,In_879,In_148);
nand U1957 (N_1957,In_304,In_1222);
or U1958 (N_1958,In_389,In_1132);
nor U1959 (N_1959,In_577,In_249);
or U1960 (N_1960,In_1410,In_915);
and U1961 (N_1961,In_456,In_256);
or U1962 (N_1962,In_1122,In_127);
xnor U1963 (N_1963,In_101,In_963);
nand U1964 (N_1964,In_644,In_410);
nor U1965 (N_1965,In_735,In_944);
xnor U1966 (N_1966,In_733,In_95);
or U1967 (N_1967,In_1154,In_881);
or U1968 (N_1968,In_999,In_992);
xor U1969 (N_1969,In_89,In_1175);
xnor U1970 (N_1970,In_390,In_978);
nand U1971 (N_1971,In_1270,In_819);
nor U1972 (N_1972,In_903,In_506);
nor U1973 (N_1973,In_600,In_310);
or U1974 (N_1974,In_1424,In_1206);
nor U1975 (N_1975,In_812,In_275);
nor U1976 (N_1976,In_755,In_1209);
and U1977 (N_1977,In_1051,In_1469);
and U1978 (N_1978,In_1075,In_1121);
xnor U1979 (N_1979,In_1075,In_438);
nor U1980 (N_1980,In_21,In_910);
or U1981 (N_1981,In_67,In_1297);
and U1982 (N_1982,In_357,In_1433);
or U1983 (N_1983,In_361,In_200);
nor U1984 (N_1984,In_695,In_770);
nand U1985 (N_1985,In_1138,In_141);
nand U1986 (N_1986,In_777,In_1095);
xnor U1987 (N_1987,In_594,In_1147);
or U1988 (N_1988,In_217,In_879);
nand U1989 (N_1989,In_413,In_1382);
and U1990 (N_1990,In_722,In_802);
nor U1991 (N_1991,In_1458,In_1014);
nor U1992 (N_1992,In_1216,In_1047);
and U1993 (N_1993,In_1303,In_442);
nand U1994 (N_1994,In_1203,In_990);
and U1995 (N_1995,In_1340,In_498);
nand U1996 (N_1996,In_745,In_772);
xor U1997 (N_1997,In_1287,In_619);
and U1998 (N_1998,In_376,In_1006);
nor U1999 (N_1999,In_372,In_244);
xor U2000 (N_2000,In_1163,In_398);
or U2001 (N_2001,In_78,In_735);
and U2002 (N_2002,In_1416,In_1180);
nor U2003 (N_2003,In_12,In_1490);
and U2004 (N_2004,In_932,In_465);
xor U2005 (N_2005,In_90,In_1075);
xor U2006 (N_2006,In_681,In_1079);
xnor U2007 (N_2007,In_1478,In_1445);
or U2008 (N_2008,In_84,In_25);
or U2009 (N_2009,In_198,In_955);
xor U2010 (N_2010,In_1327,In_997);
xor U2011 (N_2011,In_462,In_891);
or U2012 (N_2012,In_210,In_1001);
and U2013 (N_2013,In_1336,In_559);
or U2014 (N_2014,In_333,In_209);
nand U2015 (N_2015,In_1417,In_1482);
or U2016 (N_2016,In_1081,In_701);
xor U2017 (N_2017,In_1342,In_442);
nand U2018 (N_2018,In_312,In_15);
and U2019 (N_2019,In_543,In_223);
nand U2020 (N_2020,In_318,In_824);
nand U2021 (N_2021,In_1100,In_277);
and U2022 (N_2022,In_741,In_1035);
nand U2023 (N_2023,In_888,In_449);
nand U2024 (N_2024,In_961,In_1397);
nand U2025 (N_2025,In_646,In_1066);
nor U2026 (N_2026,In_19,In_1202);
xor U2027 (N_2027,In_1328,In_1114);
nor U2028 (N_2028,In_1053,In_255);
xnor U2029 (N_2029,In_300,In_642);
and U2030 (N_2030,In_1054,In_672);
or U2031 (N_2031,In_446,In_1373);
nand U2032 (N_2032,In_148,In_819);
nand U2033 (N_2033,In_784,In_920);
nor U2034 (N_2034,In_730,In_1480);
nand U2035 (N_2035,In_2,In_658);
or U2036 (N_2036,In_233,In_1177);
nand U2037 (N_2037,In_1228,In_211);
nand U2038 (N_2038,In_808,In_47);
xnor U2039 (N_2039,In_967,In_1255);
and U2040 (N_2040,In_142,In_1047);
nand U2041 (N_2041,In_1384,In_1495);
or U2042 (N_2042,In_1261,In_648);
and U2043 (N_2043,In_1228,In_1337);
xor U2044 (N_2044,In_1063,In_184);
or U2045 (N_2045,In_322,In_1120);
and U2046 (N_2046,In_41,In_148);
nand U2047 (N_2047,In_348,In_1070);
nand U2048 (N_2048,In_879,In_720);
nor U2049 (N_2049,In_896,In_544);
and U2050 (N_2050,In_160,In_104);
nor U2051 (N_2051,In_396,In_428);
and U2052 (N_2052,In_347,In_957);
xnor U2053 (N_2053,In_737,In_403);
and U2054 (N_2054,In_1224,In_1059);
xor U2055 (N_2055,In_1059,In_1167);
and U2056 (N_2056,In_770,In_74);
nor U2057 (N_2057,In_882,In_1215);
nor U2058 (N_2058,In_1290,In_1244);
nand U2059 (N_2059,In_124,In_1126);
or U2060 (N_2060,In_813,In_180);
xor U2061 (N_2061,In_1173,In_897);
nand U2062 (N_2062,In_1454,In_1359);
and U2063 (N_2063,In_654,In_866);
nand U2064 (N_2064,In_368,In_1439);
or U2065 (N_2065,In_652,In_834);
xor U2066 (N_2066,In_1057,In_431);
and U2067 (N_2067,In_463,In_648);
nand U2068 (N_2068,In_659,In_533);
nand U2069 (N_2069,In_1210,In_1094);
nor U2070 (N_2070,In_1432,In_173);
or U2071 (N_2071,In_1435,In_540);
nor U2072 (N_2072,In_46,In_1276);
xor U2073 (N_2073,In_1337,In_297);
nor U2074 (N_2074,In_1361,In_110);
and U2075 (N_2075,In_802,In_1128);
or U2076 (N_2076,In_75,In_383);
xnor U2077 (N_2077,In_129,In_34);
nand U2078 (N_2078,In_1011,In_715);
xor U2079 (N_2079,In_1462,In_1156);
xor U2080 (N_2080,In_205,In_158);
nor U2081 (N_2081,In_1112,In_107);
nand U2082 (N_2082,In_40,In_266);
nand U2083 (N_2083,In_913,In_1192);
or U2084 (N_2084,In_810,In_1116);
nor U2085 (N_2085,In_560,In_620);
or U2086 (N_2086,In_1074,In_606);
nand U2087 (N_2087,In_351,In_140);
or U2088 (N_2088,In_85,In_57);
and U2089 (N_2089,In_73,In_661);
nand U2090 (N_2090,In_163,In_1187);
xnor U2091 (N_2091,In_10,In_1496);
and U2092 (N_2092,In_943,In_1477);
or U2093 (N_2093,In_437,In_400);
nand U2094 (N_2094,In_737,In_1382);
xor U2095 (N_2095,In_818,In_615);
nand U2096 (N_2096,In_53,In_131);
and U2097 (N_2097,In_1077,In_442);
nor U2098 (N_2098,In_208,In_360);
or U2099 (N_2099,In_25,In_107);
xnor U2100 (N_2100,In_1237,In_262);
and U2101 (N_2101,In_311,In_395);
and U2102 (N_2102,In_109,In_1228);
nand U2103 (N_2103,In_1098,In_170);
or U2104 (N_2104,In_1138,In_1467);
nand U2105 (N_2105,In_1260,In_1351);
nor U2106 (N_2106,In_1001,In_900);
xor U2107 (N_2107,In_505,In_408);
or U2108 (N_2108,In_891,In_808);
and U2109 (N_2109,In_1374,In_865);
or U2110 (N_2110,In_545,In_956);
or U2111 (N_2111,In_590,In_1360);
xor U2112 (N_2112,In_634,In_499);
and U2113 (N_2113,In_1291,In_1143);
xor U2114 (N_2114,In_609,In_159);
nand U2115 (N_2115,In_782,In_215);
xnor U2116 (N_2116,In_134,In_1426);
or U2117 (N_2117,In_1478,In_801);
nand U2118 (N_2118,In_651,In_948);
xor U2119 (N_2119,In_837,In_593);
xnor U2120 (N_2120,In_305,In_276);
nor U2121 (N_2121,In_471,In_915);
xor U2122 (N_2122,In_498,In_375);
nand U2123 (N_2123,In_998,In_139);
nand U2124 (N_2124,In_570,In_260);
xnor U2125 (N_2125,In_1219,In_632);
xnor U2126 (N_2126,In_863,In_914);
nand U2127 (N_2127,In_1436,In_470);
or U2128 (N_2128,In_1055,In_479);
xor U2129 (N_2129,In_398,In_152);
nand U2130 (N_2130,In_601,In_1012);
or U2131 (N_2131,In_449,In_441);
nand U2132 (N_2132,In_993,In_1323);
nand U2133 (N_2133,In_1333,In_8);
xor U2134 (N_2134,In_75,In_1252);
and U2135 (N_2135,In_723,In_950);
xnor U2136 (N_2136,In_462,In_1417);
nand U2137 (N_2137,In_385,In_1046);
nand U2138 (N_2138,In_29,In_632);
xor U2139 (N_2139,In_407,In_1404);
and U2140 (N_2140,In_1155,In_1401);
nor U2141 (N_2141,In_636,In_583);
nor U2142 (N_2142,In_1403,In_320);
nand U2143 (N_2143,In_232,In_303);
nand U2144 (N_2144,In_727,In_592);
nor U2145 (N_2145,In_1194,In_1195);
nor U2146 (N_2146,In_1118,In_873);
xnor U2147 (N_2147,In_512,In_920);
and U2148 (N_2148,In_797,In_374);
and U2149 (N_2149,In_327,In_969);
and U2150 (N_2150,In_287,In_288);
nand U2151 (N_2151,In_3,In_430);
or U2152 (N_2152,In_1474,In_1088);
nor U2153 (N_2153,In_989,In_970);
nand U2154 (N_2154,In_1226,In_929);
or U2155 (N_2155,In_896,In_1358);
or U2156 (N_2156,In_1029,In_1480);
and U2157 (N_2157,In_413,In_1468);
and U2158 (N_2158,In_441,In_277);
nand U2159 (N_2159,In_939,In_1356);
or U2160 (N_2160,In_1142,In_707);
nand U2161 (N_2161,In_194,In_531);
and U2162 (N_2162,In_1260,In_1469);
and U2163 (N_2163,In_570,In_729);
nand U2164 (N_2164,In_1341,In_569);
and U2165 (N_2165,In_99,In_840);
or U2166 (N_2166,In_406,In_1287);
xnor U2167 (N_2167,In_1024,In_382);
nand U2168 (N_2168,In_1272,In_1498);
nand U2169 (N_2169,In_776,In_459);
nand U2170 (N_2170,In_1087,In_379);
or U2171 (N_2171,In_402,In_772);
nor U2172 (N_2172,In_665,In_533);
and U2173 (N_2173,In_153,In_449);
and U2174 (N_2174,In_1447,In_217);
nand U2175 (N_2175,In_680,In_413);
nand U2176 (N_2176,In_678,In_1261);
or U2177 (N_2177,In_207,In_494);
xnor U2178 (N_2178,In_488,In_94);
or U2179 (N_2179,In_1330,In_1044);
and U2180 (N_2180,In_760,In_767);
and U2181 (N_2181,In_317,In_484);
and U2182 (N_2182,In_1137,In_6);
nand U2183 (N_2183,In_85,In_975);
xor U2184 (N_2184,In_216,In_730);
and U2185 (N_2185,In_566,In_1397);
and U2186 (N_2186,In_1344,In_453);
nor U2187 (N_2187,In_754,In_6);
or U2188 (N_2188,In_572,In_229);
xnor U2189 (N_2189,In_1356,In_663);
nand U2190 (N_2190,In_918,In_646);
xor U2191 (N_2191,In_562,In_236);
or U2192 (N_2192,In_585,In_482);
and U2193 (N_2193,In_45,In_631);
xnor U2194 (N_2194,In_32,In_712);
nand U2195 (N_2195,In_680,In_808);
or U2196 (N_2196,In_641,In_660);
nor U2197 (N_2197,In_124,In_154);
and U2198 (N_2198,In_1006,In_110);
and U2199 (N_2199,In_1476,In_1326);
nor U2200 (N_2200,In_39,In_1426);
and U2201 (N_2201,In_6,In_1245);
xnor U2202 (N_2202,In_1228,In_608);
or U2203 (N_2203,In_900,In_1497);
xor U2204 (N_2204,In_1021,In_255);
xnor U2205 (N_2205,In_900,In_450);
or U2206 (N_2206,In_500,In_226);
nand U2207 (N_2207,In_558,In_1294);
xor U2208 (N_2208,In_951,In_1251);
nand U2209 (N_2209,In_990,In_306);
xor U2210 (N_2210,In_1069,In_309);
or U2211 (N_2211,In_453,In_1250);
and U2212 (N_2212,In_1138,In_741);
or U2213 (N_2213,In_168,In_1374);
nand U2214 (N_2214,In_313,In_189);
and U2215 (N_2215,In_850,In_21);
xnor U2216 (N_2216,In_208,In_1344);
or U2217 (N_2217,In_419,In_1284);
nand U2218 (N_2218,In_375,In_520);
and U2219 (N_2219,In_338,In_1163);
and U2220 (N_2220,In_843,In_750);
xnor U2221 (N_2221,In_886,In_1395);
nor U2222 (N_2222,In_282,In_1086);
nor U2223 (N_2223,In_725,In_766);
nor U2224 (N_2224,In_284,In_1204);
nor U2225 (N_2225,In_525,In_1158);
or U2226 (N_2226,In_1074,In_1430);
nor U2227 (N_2227,In_450,In_32);
nor U2228 (N_2228,In_1478,In_593);
and U2229 (N_2229,In_1041,In_1453);
nor U2230 (N_2230,In_1050,In_1258);
and U2231 (N_2231,In_1433,In_487);
and U2232 (N_2232,In_129,In_670);
nand U2233 (N_2233,In_363,In_414);
xor U2234 (N_2234,In_946,In_369);
or U2235 (N_2235,In_654,In_546);
nor U2236 (N_2236,In_1293,In_1009);
xnor U2237 (N_2237,In_1345,In_439);
xor U2238 (N_2238,In_561,In_482);
and U2239 (N_2239,In_623,In_339);
and U2240 (N_2240,In_1281,In_1397);
nor U2241 (N_2241,In_535,In_546);
nor U2242 (N_2242,In_1239,In_1443);
and U2243 (N_2243,In_977,In_147);
nand U2244 (N_2244,In_5,In_27);
nand U2245 (N_2245,In_847,In_1016);
xor U2246 (N_2246,In_707,In_1117);
nand U2247 (N_2247,In_619,In_1333);
nor U2248 (N_2248,In_120,In_1265);
and U2249 (N_2249,In_1146,In_760);
nand U2250 (N_2250,In_1106,In_887);
or U2251 (N_2251,In_1203,In_591);
nand U2252 (N_2252,In_789,In_433);
or U2253 (N_2253,In_1094,In_900);
and U2254 (N_2254,In_1078,In_1027);
or U2255 (N_2255,In_257,In_1424);
and U2256 (N_2256,In_319,In_1498);
or U2257 (N_2257,In_1256,In_382);
nor U2258 (N_2258,In_1415,In_1141);
or U2259 (N_2259,In_592,In_1271);
xnor U2260 (N_2260,In_1401,In_413);
and U2261 (N_2261,In_490,In_303);
xnor U2262 (N_2262,In_1161,In_1216);
and U2263 (N_2263,In_304,In_188);
nand U2264 (N_2264,In_478,In_319);
xnor U2265 (N_2265,In_1481,In_692);
nand U2266 (N_2266,In_951,In_774);
xnor U2267 (N_2267,In_478,In_1371);
xor U2268 (N_2268,In_634,In_866);
xnor U2269 (N_2269,In_194,In_721);
or U2270 (N_2270,In_200,In_884);
nor U2271 (N_2271,In_605,In_477);
or U2272 (N_2272,In_1150,In_1177);
or U2273 (N_2273,In_541,In_787);
and U2274 (N_2274,In_1382,In_1417);
xnor U2275 (N_2275,In_816,In_183);
and U2276 (N_2276,In_692,In_1384);
and U2277 (N_2277,In_1141,In_374);
or U2278 (N_2278,In_854,In_1459);
and U2279 (N_2279,In_561,In_1318);
or U2280 (N_2280,In_491,In_397);
xor U2281 (N_2281,In_1317,In_389);
xnor U2282 (N_2282,In_1170,In_1182);
xnor U2283 (N_2283,In_560,In_619);
nand U2284 (N_2284,In_1117,In_61);
or U2285 (N_2285,In_150,In_34);
nor U2286 (N_2286,In_1355,In_1027);
nor U2287 (N_2287,In_1326,In_977);
and U2288 (N_2288,In_519,In_1254);
xor U2289 (N_2289,In_894,In_144);
or U2290 (N_2290,In_833,In_1315);
nand U2291 (N_2291,In_69,In_185);
nand U2292 (N_2292,In_705,In_636);
nand U2293 (N_2293,In_773,In_3);
or U2294 (N_2294,In_911,In_840);
or U2295 (N_2295,In_1317,In_230);
and U2296 (N_2296,In_94,In_1401);
or U2297 (N_2297,In_568,In_1235);
xnor U2298 (N_2298,In_110,In_943);
nor U2299 (N_2299,In_266,In_1205);
nor U2300 (N_2300,In_697,In_36);
xor U2301 (N_2301,In_451,In_44);
nor U2302 (N_2302,In_833,In_1319);
or U2303 (N_2303,In_367,In_860);
nor U2304 (N_2304,In_1300,In_135);
nor U2305 (N_2305,In_835,In_1147);
and U2306 (N_2306,In_1036,In_341);
nor U2307 (N_2307,In_1331,In_1131);
xor U2308 (N_2308,In_702,In_606);
nor U2309 (N_2309,In_1231,In_774);
nand U2310 (N_2310,In_497,In_67);
or U2311 (N_2311,In_1388,In_1232);
nand U2312 (N_2312,In_843,In_541);
nand U2313 (N_2313,In_495,In_301);
xnor U2314 (N_2314,In_1247,In_875);
or U2315 (N_2315,In_1092,In_192);
nor U2316 (N_2316,In_755,In_892);
nand U2317 (N_2317,In_1197,In_87);
nor U2318 (N_2318,In_460,In_1005);
or U2319 (N_2319,In_697,In_235);
xor U2320 (N_2320,In_156,In_1452);
nand U2321 (N_2321,In_731,In_1181);
nor U2322 (N_2322,In_378,In_1102);
xor U2323 (N_2323,In_917,In_567);
nand U2324 (N_2324,In_65,In_834);
and U2325 (N_2325,In_122,In_1156);
nand U2326 (N_2326,In_1430,In_590);
xnor U2327 (N_2327,In_1323,In_1038);
and U2328 (N_2328,In_1442,In_1477);
nor U2329 (N_2329,In_752,In_414);
nand U2330 (N_2330,In_1490,In_1172);
nor U2331 (N_2331,In_1273,In_552);
and U2332 (N_2332,In_144,In_66);
nand U2333 (N_2333,In_427,In_1028);
nor U2334 (N_2334,In_644,In_786);
or U2335 (N_2335,In_93,In_1324);
xnor U2336 (N_2336,In_384,In_987);
or U2337 (N_2337,In_208,In_397);
or U2338 (N_2338,In_826,In_218);
nand U2339 (N_2339,In_1396,In_1450);
xor U2340 (N_2340,In_802,In_1204);
nor U2341 (N_2341,In_1094,In_707);
nor U2342 (N_2342,In_555,In_571);
xnor U2343 (N_2343,In_728,In_929);
and U2344 (N_2344,In_534,In_1282);
nor U2345 (N_2345,In_507,In_613);
nor U2346 (N_2346,In_1041,In_205);
nor U2347 (N_2347,In_40,In_1094);
xor U2348 (N_2348,In_539,In_925);
and U2349 (N_2349,In_278,In_1207);
or U2350 (N_2350,In_88,In_872);
and U2351 (N_2351,In_1047,In_434);
nand U2352 (N_2352,In_1085,In_964);
or U2353 (N_2353,In_1152,In_1424);
nor U2354 (N_2354,In_670,In_924);
nand U2355 (N_2355,In_847,In_839);
nor U2356 (N_2356,In_820,In_1055);
nor U2357 (N_2357,In_976,In_1172);
nor U2358 (N_2358,In_140,In_622);
nand U2359 (N_2359,In_1175,In_351);
and U2360 (N_2360,In_1109,In_1384);
nor U2361 (N_2361,In_1240,In_23);
nor U2362 (N_2362,In_771,In_481);
nor U2363 (N_2363,In_1390,In_1053);
xor U2364 (N_2364,In_547,In_1315);
xnor U2365 (N_2365,In_1274,In_941);
nand U2366 (N_2366,In_571,In_764);
xor U2367 (N_2367,In_824,In_54);
and U2368 (N_2368,In_595,In_487);
xnor U2369 (N_2369,In_503,In_324);
and U2370 (N_2370,In_612,In_1317);
xor U2371 (N_2371,In_1187,In_958);
and U2372 (N_2372,In_466,In_407);
and U2373 (N_2373,In_1456,In_394);
and U2374 (N_2374,In_1052,In_1041);
or U2375 (N_2375,In_1293,In_1262);
and U2376 (N_2376,In_179,In_1438);
nand U2377 (N_2377,In_573,In_825);
nor U2378 (N_2378,In_1059,In_1249);
or U2379 (N_2379,In_435,In_869);
xnor U2380 (N_2380,In_1140,In_1189);
or U2381 (N_2381,In_974,In_957);
nor U2382 (N_2382,In_1446,In_1263);
or U2383 (N_2383,In_55,In_957);
xnor U2384 (N_2384,In_434,In_1230);
xor U2385 (N_2385,In_1162,In_767);
nand U2386 (N_2386,In_270,In_1487);
and U2387 (N_2387,In_797,In_1371);
nand U2388 (N_2388,In_1307,In_524);
nand U2389 (N_2389,In_1149,In_1092);
or U2390 (N_2390,In_846,In_409);
and U2391 (N_2391,In_1371,In_71);
or U2392 (N_2392,In_505,In_1240);
nor U2393 (N_2393,In_604,In_471);
nand U2394 (N_2394,In_864,In_470);
or U2395 (N_2395,In_1103,In_1238);
xnor U2396 (N_2396,In_815,In_1116);
or U2397 (N_2397,In_1108,In_445);
nand U2398 (N_2398,In_479,In_1165);
nor U2399 (N_2399,In_494,In_1421);
or U2400 (N_2400,In_803,In_317);
nand U2401 (N_2401,In_963,In_1470);
xnor U2402 (N_2402,In_1419,In_781);
nor U2403 (N_2403,In_333,In_204);
or U2404 (N_2404,In_397,In_1218);
nor U2405 (N_2405,In_736,In_33);
xnor U2406 (N_2406,In_411,In_555);
nand U2407 (N_2407,In_899,In_554);
and U2408 (N_2408,In_621,In_876);
xnor U2409 (N_2409,In_1362,In_300);
or U2410 (N_2410,In_1486,In_78);
xor U2411 (N_2411,In_873,In_863);
nand U2412 (N_2412,In_639,In_224);
xnor U2413 (N_2413,In_1453,In_1120);
and U2414 (N_2414,In_974,In_1256);
nand U2415 (N_2415,In_1046,In_473);
xnor U2416 (N_2416,In_847,In_732);
and U2417 (N_2417,In_196,In_377);
xnor U2418 (N_2418,In_538,In_57);
or U2419 (N_2419,In_1143,In_509);
and U2420 (N_2420,In_380,In_235);
and U2421 (N_2421,In_780,In_1366);
nor U2422 (N_2422,In_765,In_1039);
nor U2423 (N_2423,In_64,In_1194);
or U2424 (N_2424,In_702,In_485);
nor U2425 (N_2425,In_664,In_1317);
or U2426 (N_2426,In_1180,In_321);
nand U2427 (N_2427,In_474,In_398);
or U2428 (N_2428,In_155,In_694);
and U2429 (N_2429,In_570,In_285);
xnor U2430 (N_2430,In_1498,In_1105);
nor U2431 (N_2431,In_41,In_688);
xnor U2432 (N_2432,In_1090,In_486);
nand U2433 (N_2433,In_483,In_1477);
and U2434 (N_2434,In_1167,In_1129);
nor U2435 (N_2435,In_774,In_1069);
and U2436 (N_2436,In_1409,In_1223);
and U2437 (N_2437,In_193,In_1163);
and U2438 (N_2438,In_1182,In_633);
xnor U2439 (N_2439,In_268,In_1301);
or U2440 (N_2440,In_764,In_1045);
nor U2441 (N_2441,In_546,In_741);
or U2442 (N_2442,In_123,In_42);
nand U2443 (N_2443,In_637,In_957);
or U2444 (N_2444,In_702,In_269);
nor U2445 (N_2445,In_350,In_907);
nand U2446 (N_2446,In_610,In_152);
or U2447 (N_2447,In_108,In_829);
or U2448 (N_2448,In_484,In_187);
nand U2449 (N_2449,In_909,In_881);
nand U2450 (N_2450,In_1049,In_239);
nor U2451 (N_2451,In_1379,In_1041);
nand U2452 (N_2452,In_203,In_581);
and U2453 (N_2453,In_356,In_94);
xnor U2454 (N_2454,In_1301,In_1243);
nand U2455 (N_2455,In_166,In_215);
xor U2456 (N_2456,In_1007,In_622);
nor U2457 (N_2457,In_956,In_1443);
xor U2458 (N_2458,In_309,In_1105);
nor U2459 (N_2459,In_404,In_747);
or U2460 (N_2460,In_195,In_1369);
nand U2461 (N_2461,In_823,In_465);
or U2462 (N_2462,In_1325,In_22);
or U2463 (N_2463,In_1329,In_72);
xor U2464 (N_2464,In_1303,In_501);
or U2465 (N_2465,In_995,In_1065);
xor U2466 (N_2466,In_958,In_836);
xor U2467 (N_2467,In_1139,In_31);
nor U2468 (N_2468,In_1453,In_1067);
xnor U2469 (N_2469,In_177,In_855);
xnor U2470 (N_2470,In_608,In_288);
nor U2471 (N_2471,In_141,In_1060);
xnor U2472 (N_2472,In_957,In_211);
nand U2473 (N_2473,In_1195,In_1163);
or U2474 (N_2474,In_347,In_1125);
and U2475 (N_2475,In_64,In_957);
xor U2476 (N_2476,In_376,In_1377);
xor U2477 (N_2477,In_548,In_518);
and U2478 (N_2478,In_1225,In_138);
nor U2479 (N_2479,In_1119,In_77);
nor U2480 (N_2480,In_343,In_1240);
and U2481 (N_2481,In_743,In_378);
xor U2482 (N_2482,In_454,In_139);
or U2483 (N_2483,In_291,In_624);
nor U2484 (N_2484,In_295,In_555);
xnor U2485 (N_2485,In_1493,In_1081);
or U2486 (N_2486,In_358,In_1263);
nand U2487 (N_2487,In_488,In_1026);
xor U2488 (N_2488,In_436,In_1125);
nor U2489 (N_2489,In_392,In_973);
nand U2490 (N_2490,In_1201,In_521);
nand U2491 (N_2491,In_90,In_119);
or U2492 (N_2492,In_1295,In_472);
nor U2493 (N_2493,In_10,In_446);
nor U2494 (N_2494,In_235,In_523);
xnor U2495 (N_2495,In_722,In_1255);
nor U2496 (N_2496,In_1396,In_865);
or U2497 (N_2497,In_204,In_549);
or U2498 (N_2498,In_1090,In_411);
and U2499 (N_2499,In_94,In_599);
nor U2500 (N_2500,In_863,In_1443);
and U2501 (N_2501,In_535,In_1441);
or U2502 (N_2502,In_815,In_87);
xor U2503 (N_2503,In_256,In_860);
and U2504 (N_2504,In_1260,In_451);
nor U2505 (N_2505,In_1273,In_1282);
or U2506 (N_2506,In_899,In_682);
and U2507 (N_2507,In_1448,In_122);
xnor U2508 (N_2508,In_603,In_439);
or U2509 (N_2509,In_699,In_1035);
nor U2510 (N_2510,In_1347,In_1319);
xnor U2511 (N_2511,In_841,In_861);
or U2512 (N_2512,In_552,In_1220);
nor U2513 (N_2513,In_1174,In_386);
nand U2514 (N_2514,In_1077,In_706);
or U2515 (N_2515,In_158,In_202);
nor U2516 (N_2516,In_937,In_261);
xor U2517 (N_2517,In_1361,In_413);
xor U2518 (N_2518,In_57,In_773);
xnor U2519 (N_2519,In_1193,In_1225);
or U2520 (N_2520,In_456,In_339);
or U2521 (N_2521,In_1113,In_1015);
or U2522 (N_2522,In_31,In_400);
nand U2523 (N_2523,In_863,In_17);
xor U2524 (N_2524,In_1138,In_1395);
nor U2525 (N_2525,In_847,In_1433);
or U2526 (N_2526,In_122,In_792);
xor U2527 (N_2527,In_890,In_728);
nand U2528 (N_2528,In_719,In_748);
and U2529 (N_2529,In_1439,In_144);
xnor U2530 (N_2530,In_635,In_1411);
nand U2531 (N_2531,In_1402,In_116);
xor U2532 (N_2532,In_625,In_535);
or U2533 (N_2533,In_1015,In_734);
or U2534 (N_2534,In_439,In_1334);
and U2535 (N_2535,In_251,In_1414);
nor U2536 (N_2536,In_763,In_226);
xnor U2537 (N_2537,In_1315,In_1267);
or U2538 (N_2538,In_180,In_1430);
nor U2539 (N_2539,In_15,In_1017);
nand U2540 (N_2540,In_902,In_285);
nor U2541 (N_2541,In_872,In_63);
nand U2542 (N_2542,In_1049,In_87);
nand U2543 (N_2543,In_793,In_609);
nor U2544 (N_2544,In_1302,In_344);
nand U2545 (N_2545,In_1064,In_68);
or U2546 (N_2546,In_471,In_1118);
nor U2547 (N_2547,In_97,In_285);
and U2548 (N_2548,In_704,In_1180);
or U2549 (N_2549,In_1492,In_59);
nand U2550 (N_2550,In_340,In_1026);
nor U2551 (N_2551,In_702,In_730);
xnor U2552 (N_2552,In_858,In_1202);
and U2553 (N_2553,In_1456,In_485);
and U2554 (N_2554,In_460,In_413);
nand U2555 (N_2555,In_579,In_1192);
or U2556 (N_2556,In_419,In_1172);
nor U2557 (N_2557,In_192,In_319);
and U2558 (N_2558,In_1200,In_1404);
nand U2559 (N_2559,In_826,In_478);
and U2560 (N_2560,In_1387,In_151);
nor U2561 (N_2561,In_134,In_895);
nor U2562 (N_2562,In_1164,In_464);
nand U2563 (N_2563,In_319,In_967);
or U2564 (N_2564,In_525,In_687);
and U2565 (N_2565,In_1375,In_389);
or U2566 (N_2566,In_1004,In_884);
or U2567 (N_2567,In_1483,In_1215);
nor U2568 (N_2568,In_1322,In_1357);
and U2569 (N_2569,In_1013,In_906);
or U2570 (N_2570,In_184,In_922);
xor U2571 (N_2571,In_738,In_697);
and U2572 (N_2572,In_1423,In_1229);
nor U2573 (N_2573,In_809,In_1470);
xor U2574 (N_2574,In_1007,In_573);
or U2575 (N_2575,In_1199,In_556);
and U2576 (N_2576,In_137,In_1311);
nor U2577 (N_2577,In_885,In_1411);
or U2578 (N_2578,In_1370,In_1455);
nor U2579 (N_2579,In_1346,In_957);
or U2580 (N_2580,In_683,In_1374);
nand U2581 (N_2581,In_74,In_21);
xnor U2582 (N_2582,In_300,In_739);
nand U2583 (N_2583,In_911,In_168);
and U2584 (N_2584,In_861,In_375);
nand U2585 (N_2585,In_991,In_1425);
xor U2586 (N_2586,In_6,In_1206);
nand U2587 (N_2587,In_901,In_716);
nand U2588 (N_2588,In_1490,In_1098);
and U2589 (N_2589,In_75,In_57);
or U2590 (N_2590,In_33,In_1239);
and U2591 (N_2591,In_1472,In_860);
or U2592 (N_2592,In_389,In_897);
nand U2593 (N_2593,In_519,In_1093);
nor U2594 (N_2594,In_1106,In_591);
xnor U2595 (N_2595,In_1045,In_207);
or U2596 (N_2596,In_1464,In_799);
or U2597 (N_2597,In_357,In_270);
xnor U2598 (N_2598,In_1414,In_1187);
and U2599 (N_2599,In_768,In_1428);
and U2600 (N_2600,In_1376,In_1098);
and U2601 (N_2601,In_973,In_338);
and U2602 (N_2602,In_1163,In_667);
xnor U2603 (N_2603,In_356,In_527);
and U2604 (N_2604,In_180,In_770);
and U2605 (N_2605,In_1442,In_856);
xor U2606 (N_2606,In_871,In_840);
and U2607 (N_2607,In_71,In_674);
nor U2608 (N_2608,In_811,In_804);
nand U2609 (N_2609,In_32,In_1080);
xor U2610 (N_2610,In_259,In_1493);
xor U2611 (N_2611,In_33,In_67);
and U2612 (N_2612,In_949,In_1467);
or U2613 (N_2613,In_309,In_1339);
or U2614 (N_2614,In_1133,In_949);
xnor U2615 (N_2615,In_1354,In_313);
or U2616 (N_2616,In_15,In_382);
nand U2617 (N_2617,In_971,In_851);
xor U2618 (N_2618,In_848,In_299);
nor U2619 (N_2619,In_700,In_1266);
and U2620 (N_2620,In_779,In_80);
and U2621 (N_2621,In_137,In_1481);
xor U2622 (N_2622,In_1110,In_1440);
and U2623 (N_2623,In_49,In_649);
nor U2624 (N_2624,In_160,In_335);
xnor U2625 (N_2625,In_682,In_93);
and U2626 (N_2626,In_945,In_1281);
xor U2627 (N_2627,In_1224,In_1299);
nand U2628 (N_2628,In_430,In_830);
nor U2629 (N_2629,In_898,In_894);
xnor U2630 (N_2630,In_1088,In_811);
xnor U2631 (N_2631,In_1164,In_940);
and U2632 (N_2632,In_138,In_1299);
or U2633 (N_2633,In_1164,In_1035);
or U2634 (N_2634,In_717,In_1102);
and U2635 (N_2635,In_690,In_536);
nand U2636 (N_2636,In_839,In_1478);
and U2637 (N_2637,In_1366,In_1112);
and U2638 (N_2638,In_1408,In_363);
xnor U2639 (N_2639,In_1491,In_262);
and U2640 (N_2640,In_803,In_3);
nor U2641 (N_2641,In_915,In_1273);
xnor U2642 (N_2642,In_1321,In_347);
nor U2643 (N_2643,In_992,In_484);
and U2644 (N_2644,In_1146,In_828);
and U2645 (N_2645,In_114,In_550);
xor U2646 (N_2646,In_1120,In_535);
nand U2647 (N_2647,In_1020,In_1359);
xor U2648 (N_2648,In_1101,In_500);
nand U2649 (N_2649,In_1172,In_591);
nor U2650 (N_2650,In_1111,In_569);
nand U2651 (N_2651,In_664,In_403);
and U2652 (N_2652,In_767,In_1163);
nor U2653 (N_2653,In_0,In_638);
or U2654 (N_2654,In_686,In_1174);
and U2655 (N_2655,In_817,In_1359);
nor U2656 (N_2656,In_306,In_801);
nand U2657 (N_2657,In_1244,In_862);
nand U2658 (N_2658,In_430,In_1213);
or U2659 (N_2659,In_781,In_91);
or U2660 (N_2660,In_1271,In_1026);
nand U2661 (N_2661,In_1068,In_1297);
nor U2662 (N_2662,In_1334,In_1484);
nand U2663 (N_2663,In_318,In_1330);
nand U2664 (N_2664,In_661,In_1068);
or U2665 (N_2665,In_546,In_1242);
or U2666 (N_2666,In_629,In_886);
nand U2667 (N_2667,In_766,In_984);
and U2668 (N_2668,In_317,In_520);
nand U2669 (N_2669,In_1446,In_579);
or U2670 (N_2670,In_1288,In_1462);
xor U2671 (N_2671,In_713,In_1246);
nor U2672 (N_2672,In_1027,In_201);
and U2673 (N_2673,In_1284,In_476);
xor U2674 (N_2674,In_164,In_380);
and U2675 (N_2675,In_765,In_935);
and U2676 (N_2676,In_518,In_1125);
or U2677 (N_2677,In_240,In_178);
and U2678 (N_2678,In_325,In_816);
and U2679 (N_2679,In_514,In_977);
or U2680 (N_2680,In_1392,In_675);
nor U2681 (N_2681,In_190,In_601);
and U2682 (N_2682,In_1008,In_1141);
and U2683 (N_2683,In_126,In_597);
nor U2684 (N_2684,In_476,In_629);
nor U2685 (N_2685,In_155,In_1251);
nand U2686 (N_2686,In_356,In_523);
nor U2687 (N_2687,In_981,In_136);
nand U2688 (N_2688,In_778,In_471);
xnor U2689 (N_2689,In_1061,In_249);
nand U2690 (N_2690,In_259,In_439);
nor U2691 (N_2691,In_1416,In_961);
and U2692 (N_2692,In_140,In_1084);
xnor U2693 (N_2693,In_1386,In_706);
nor U2694 (N_2694,In_527,In_462);
and U2695 (N_2695,In_1197,In_473);
or U2696 (N_2696,In_1017,In_95);
and U2697 (N_2697,In_1488,In_758);
xor U2698 (N_2698,In_437,In_764);
and U2699 (N_2699,In_218,In_1066);
xnor U2700 (N_2700,In_393,In_1418);
xnor U2701 (N_2701,In_1232,In_498);
or U2702 (N_2702,In_1251,In_167);
and U2703 (N_2703,In_1246,In_1436);
nand U2704 (N_2704,In_1161,In_79);
xor U2705 (N_2705,In_998,In_890);
nand U2706 (N_2706,In_413,In_355);
or U2707 (N_2707,In_1356,In_821);
and U2708 (N_2708,In_1360,In_786);
and U2709 (N_2709,In_1221,In_1166);
or U2710 (N_2710,In_1402,In_1209);
or U2711 (N_2711,In_487,In_1003);
xnor U2712 (N_2712,In_640,In_1224);
xor U2713 (N_2713,In_1239,In_1122);
and U2714 (N_2714,In_768,In_846);
nor U2715 (N_2715,In_438,In_640);
xnor U2716 (N_2716,In_375,In_75);
and U2717 (N_2717,In_891,In_803);
nor U2718 (N_2718,In_1279,In_619);
nor U2719 (N_2719,In_299,In_1463);
or U2720 (N_2720,In_1467,In_25);
and U2721 (N_2721,In_1176,In_367);
nand U2722 (N_2722,In_680,In_1185);
nand U2723 (N_2723,In_754,In_197);
nor U2724 (N_2724,In_331,In_162);
nor U2725 (N_2725,In_123,In_634);
and U2726 (N_2726,In_703,In_687);
nor U2727 (N_2727,In_778,In_672);
nor U2728 (N_2728,In_429,In_1055);
xnor U2729 (N_2729,In_1059,In_716);
and U2730 (N_2730,In_936,In_624);
or U2731 (N_2731,In_977,In_677);
xor U2732 (N_2732,In_575,In_458);
nor U2733 (N_2733,In_1273,In_251);
or U2734 (N_2734,In_796,In_451);
and U2735 (N_2735,In_1480,In_955);
or U2736 (N_2736,In_708,In_582);
or U2737 (N_2737,In_600,In_542);
xnor U2738 (N_2738,In_588,In_935);
and U2739 (N_2739,In_1207,In_1215);
and U2740 (N_2740,In_13,In_1333);
xnor U2741 (N_2741,In_1045,In_149);
or U2742 (N_2742,In_1127,In_99);
nand U2743 (N_2743,In_294,In_248);
nor U2744 (N_2744,In_699,In_100);
or U2745 (N_2745,In_549,In_1133);
xor U2746 (N_2746,In_631,In_214);
xor U2747 (N_2747,In_714,In_1322);
and U2748 (N_2748,In_789,In_1274);
and U2749 (N_2749,In_1180,In_442);
nand U2750 (N_2750,In_1072,In_1013);
nor U2751 (N_2751,In_1465,In_1163);
nand U2752 (N_2752,In_40,In_610);
or U2753 (N_2753,In_970,In_866);
and U2754 (N_2754,In_941,In_1448);
nor U2755 (N_2755,In_363,In_802);
and U2756 (N_2756,In_1049,In_1397);
or U2757 (N_2757,In_222,In_616);
and U2758 (N_2758,In_888,In_687);
and U2759 (N_2759,In_685,In_476);
nand U2760 (N_2760,In_423,In_1495);
nand U2761 (N_2761,In_598,In_47);
or U2762 (N_2762,In_714,In_1319);
xnor U2763 (N_2763,In_276,In_1070);
xnor U2764 (N_2764,In_1345,In_1144);
and U2765 (N_2765,In_190,In_452);
and U2766 (N_2766,In_279,In_59);
or U2767 (N_2767,In_882,In_548);
nand U2768 (N_2768,In_731,In_1009);
or U2769 (N_2769,In_969,In_1022);
nand U2770 (N_2770,In_1074,In_187);
nand U2771 (N_2771,In_702,In_1385);
nor U2772 (N_2772,In_971,In_459);
and U2773 (N_2773,In_1229,In_69);
and U2774 (N_2774,In_1130,In_668);
nor U2775 (N_2775,In_450,In_19);
or U2776 (N_2776,In_657,In_499);
xor U2777 (N_2777,In_863,In_20);
nand U2778 (N_2778,In_404,In_1335);
xor U2779 (N_2779,In_1054,In_1426);
or U2780 (N_2780,In_1285,In_267);
or U2781 (N_2781,In_1472,In_1284);
or U2782 (N_2782,In_817,In_881);
nand U2783 (N_2783,In_801,In_1407);
xor U2784 (N_2784,In_691,In_865);
and U2785 (N_2785,In_3,In_449);
and U2786 (N_2786,In_287,In_137);
and U2787 (N_2787,In_134,In_72);
nand U2788 (N_2788,In_1145,In_1079);
or U2789 (N_2789,In_572,In_961);
or U2790 (N_2790,In_114,In_68);
xnor U2791 (N_2791,In_1118,In_1186);
nand U2792 (N_2792,In_234,In_1030);
and U2793 (N_2793,In_1387,In_1219);
or U2794 (N_2794,In_246,In_171);
nor U2795 (N_2795,In_404,In_419);
nor U2796 (N_2796,In_1405,In_1432);
and U2797 (N_2797,In_567,In_1199);
or U2798 (N_2798,In_599,In_1458);
xor U2799 (N_2799,In_741,In_1140);
or U2800 (N_2800,In_344,In_839);
xnor U2801 (N_2801,In_1333,In_965);
nor U2802 (N_2802,In_256,In_730);
or U2803 (N_2803,In_657,In_1413);
or U2804 (N_2804,In_1287,In_1465);
or U2805 (N_2805,In_1192,In_960);
nor U2806 (N_2806,In_818,In_1205);
nand U2807 (N_2807,In_1433,In_173);
xor U2808 (N_2808,In_1060,In_181);
and U2809 (N_2809,In_1284,In_649);
nor U2810 (N_2810,In_873,In_872);
nand U2811 (N_2811,In_670,In_507);
xnor U2812 (N_2812,In_1166,In_446);
nand U2813 (N_2813,In_1381,In_158);
nand U2814 (N_2814,In_1169,In_232);
nor U2815 (N_2815,In_1003,In_1314);
and U2816 (N_2816,In_1353,In_1184);
xnor U2817 (N_2817,In_952,In_280);
xor U2818 (N_2818,In_933,In_729);
nor U2819 (N_2819,In_1010,In_387);
nand U2820 (N_2820,In_1085,In_1236);
or U2821 (N_2821,In_165,In_1087);
or U2822 (N_2822,In_668,In_658);
nor U2823 (N_2823,In_616,In_831);
xnor U2824 (N_2824,In_884,In_490);
xor U2825 (N_2825,In_790,In_1205);
and U2826 (N_2826,In_1257,In_336);
and U2827 (N_2827,In_446,In_192);
xnor U2828 (N_2828,In_902,In_871);
xor U2829 (N_2829,In_413,In_1191);
or U2830 (N_2830,In_197,In_1149);
nor U2831 (N_2831,In_1305,In_1157);
xor U2832 (N_2832,In_1091,In_1096);
nor U2833 (N_2833,In_444,In_123);
xor U2834 (N_2834,In_1277,In_768);
or U2835 (N_2835,In_869,In_950);
nor U2836 (N_2836,In_979,In_845);
nand U2837 (N_2837,In_442,In_469);
or U2838 (N_2838,In_1129,In_1398);
nor U2839 (N_2839,In_1414,In_1349);
or U2840 (N_2840,In_457,In_646);
xor U2841 (N_2841,In_80,In_369);
nand U2842 (N_2842,In_452,In_1330);
or U2843 (N_2843,In_1481,In_1440);
and U2844 (N_2844,In_993,In_367);
or U2845 (N_2845,In_1130,In_765);
and U2846 (N_2846,In_1060,In_85);
and U2847 (N_2847,In_887,In_1354);
nor U2848 (N_2848,In_1400,In_9);
nor U2849 (N_2849,In_228,In_1467);
xnor U2850 (N_2850,In_240,In_813);
xor U2851 (N_2851,In_176,In_667);
or U2852 (N_2852,In_11,In_886);
xnor U2853 (N_2853,In_736,In_348);
nand U2854 (N_2854,In_1075,In_1047);
xnor U2855 (N_2855,In_457,In_917);
nand U2856 (N_2856,In_274,In_834);
xnor U2857 (N_2857,In_936,In_949);
xor U2858 (N_2858,In_652,In_1285);
and U2859 (N_2859,In_1438,In_1345);
nor U2860 (N_2860,In_1355,In_234);
nand U2861 (N_2861,In_240,In_275);
xnor U2862 (N_2862,In_1343,In_1457);
xnor U2863 (N_2863,In_519,In_989);
nand U2864 (N_2864,In_957,In_1059);
and U2865 (N_2865,In_1430,In_490);
nand U2866 (N_2866,In_521,In_131);
xnor U2867 (N_2867,In_331,In_565);
and U2868 (N_2868,In_559,In_4);
and U2869 (N_2869,In_1050,In_1372);
or U2870 (N_2870,In_540,In_222);
nand U2871 (N_2871,In_1147,In_146);
nor U2872 (N_2872,In_72,In_636);
nand U2873 (N_2873,In_592,In_1058);
nor U2874 (N_2874,In_151,In_187);
xor U2875 (N_2875,In_175,In_978);
nor U2876 (N_2876,In_792,In_708);
or U2877 (N_2877,In_201,In_1316);
xnor U2878 (N_2878,In_1236,In_1426);
xnor U2879 (N_2879,In_786,In_962);
xor U2880 (N_2880,In_887,In_196);
nor U2881 (N_2881,In_614,In_2);
xor U2882 (N_2882,In_302,In_5);
and U2883 (N_2883,In_635,In_78);
and U2884 (N_2884,In_806,In_960);
nor U2885 (N_2885,In_127,In_931);
and U2886 (N_2886,In_196,In_544);
or U2887 (N_2887,In_773,In_1328);
nor U2888 (N_2888,In_769,In_177);
nor U2889 (N_2889,In_1319,In_851);
xnor U2890 (N_2890,In_336,In_1416);
nor U2891 (N_2891,In_400,In_908);
xor U2892 (N_2892,In_307,In_1125);
xor U2893 (N_2893,In_395,In_924);
or U2894 (N_2894,In_927,In_0);
nand U2895 (N_2895,In_382,In_1238);
xor U2896 (N_2896,In_530,In_1407);
or U2897 (N_2897,In_208,In_972);
and U2898 (N_2898,In_1254,In_822);
xnor U2899 (N_2899,In_425,In_408);
nand U2900 (N_2900,In_482,In_1354);
nand U2901 (N_2901,In_1103,In_1317);
or U2902 (N_2902,In_1284,In_371);
nand U2903 (N_2903,In_1141,In_216);
nor U2904 (N_2904,In_103,In_1147);
nor U2905 (N_2905,In_896,In_1252);
or U2906 (N_2906,In_1237,In_247);
nor U2907 (N_2907,In_961,In_733);
nand U2908 (N_2908,In_1250,In_34);
xnor U2909 (N_2909,In_1421,In_1067);
or U2910 (N_2910,In_897,In_814);
nand U2911 (N_2911,In_1283,In_1453);
xnor U2912 (N_2912,In_893,In_1369);
and U2913 (N_2913,In_588,In_1095);
and U2914 (N_2914,In_1064,In_410);
nor U2915 (N_2915,In_1233,In_1047);
and U2916 (N_2916,In_757,In_1049);
nand U2917 (N_2917,In_1220,In_720);
nand U2918 (N_2918,In_972,In_302);
nor U2919 (N_2919,In_565,In_435);
nor U2920 (N_2920,In_893,In_1284);
xnor U2921 (N_2921,In_371,In_645);
xor U2922 (N_2922,In_1075,In_316);
and U2923 (N_2923,In_19,In_404);
nor U2924 (N_2924,In_62,In_470);
nor U2925 (N_2925,In_3,In_961);
and U2926 (N_2926,In_1082,In_29);
xor U2927 (N_2927,In_1352,In_605);
or U2928 (N_2928,In_1188,In_461);
and U2929 (N_2929,In_1220,In_218);
and U2930 (N_2930,In_1479,In_1208);
nand U2931 (N_2931,In_702,In_1476);
and U2932 (N_2932,In_7,In_641);
nor U2933 (N_2933,In_911,In_206);
nor U2934 (N_2934,In_1473,In_1279);
nand U2935 (N_2935,In_550,In_514);
nand U2936 (N_2936,In_406,In_924);
or U2937 (N_2937,In_1345,In_923);
xor U2938 (N_2938,In_614,In_73);
and U2939 (N_2939,In_241,In_773);
or U2940 (N_2940,In_261,In_1458);
nor U2941 (N_2941,In_128,In_1033);
nand U2942 (N_2942,In_450,In_521);
nor U2943 (N_2943,In_444,In_1117);
nor U2944 (N_2944,In_621,In_829);
or U2945 (N_2945,In_410,In_604);
nor U2946 (N_2946,In_97,In_939);
nor U2947 (N_2947,In_414,In_275);
or U2948 (N_2948,In_835,In_574);
nor U2949 (N_2949,In_332,In_1345);
or U2950 (N_2950,In_1444,In_1078);
nor U2951 (N_2951,In_522,In_427);
nor U2952 (N_2952,In_256,In_1293);
and U2953 (N_2953,In_452,In_1346);
xor U2954 (N_2954,In_335,In_1004);
and U2955 (N_2955,In_501,In_696);
nor U2956 (N_2956,In_336,In_89);
and U2957 (N_2957,In_208,In_326);
and U2958 (N_2958,In_642,In_630);
or U2959 (N_2959,In_269,In_1051);
nand U2960 (N_2960,In_1365,In_1336);
nor U2961 (N_2961,In_274,In_88);
or U2962 (N_2962,In_6,In_42);
nor U2963 (N_2963,In_366,In_213);
or U2964 (N_2964,In_86,In_558);
and U2965 (N_2965,In_468,In_526);
and U2966 (N_2966,In_727,In_960);
nand U2967 (N_2967,In_180,In_301);
and U2968 (N_2968,In_826,In_1099);
nor U2969 (N_2969,In_512,In_1202);
nor U2970 (N_2970,In_1381,In_271);
nor U2971 (N_2971,In_1146,In_797);
or U2972 (N_2972,In_79,In_1081);
or U2973 (N_2973,In_1126,In_1328);
xnor U2974 (N_2974,In_1432,In_890);
and U2975 (N_2975,In_780,In_1355);
nor U2976 (N_2976,In_255,In_176);
and U2977 (N_2977,In_1176,In_570);
xnor U2978 (N_2978,In_306,In_1327);
nand U2979 (N_2979,In_729,In_1300);
nand U2980 (N_2980,In_1034,In_1345);
nand U2981 (N_2981,In_1153,In_259);
nand U2982 (N_2982,In_1212,In_1313);
and U2983 (N_2983,In_59,In_285);
nor U2984 (N_2984,In_1331,In_1191);
or U2985 (N_2985,In_897,In_96);
and U2986 (N_2986,In_437,In_1438);
nand U2987 (N_2987,In_1262,In_590);
xnor U2988 (N_2988,In_1166,In_1344);
and U2989 (N_2989,In_1408,In_977);
nor U2990 (N_2990,In_145,In_1189);
nand U2991 (N_2991,In_513,In_869);
nand U2992 (N_2992,In_1337,In_1206);
or U2993 (N_2993,In_1063,In_345);
or U2994 (N_2994,In_605,In_1432);
nor U2995 (N_2995,In_893,In_1327);
nor U2996 (N_2996,In_337,In_994);
or U2997 (N_2997,In_1319,In_314);
or U2998 (N_2998,In_667,In_244);
or U2999 (N_2999,In_1433,In_1156);
nor U3000 (N_3000,N_1379,N_2162);
or U3001 (N_3001,N_2113,N_1179);
xor U3002 (N_3002,N_26,N_1418);
and U3003 (N_3003,N_1031,N_2972);
and U3004 (N_3004,N_377,N_395);
or U3005 (N_3005,N_689,N_732);
and U3006 (N_3006,N_1820,N_2659);
xor U3007 (N_3007,N_765,N_118);
nor U3008 (N_3008,N_91,N_185);
nand U3009 (N_3009,N_2880,N_133);
xnor U3010 (N_3010,N_772,N_2188);
nand U3011 (N_3011,N_2121,N_626);
xor U3012 (N_3012,N_1568,N_2053);
or U3013 (N_3013,N_2490,N_2349);
or U3014 (N_3014,N_1732,N_969);
and U3015 (N_3015,N_1902,N_679);
or U3016 (N_3016,N_2205,N_2954);
nand U3017 (N_3017,N_2872,N_1480);
and U3018 (N_3018,N_2437,N_50);
xor U3019 (N_3019,N_620,N_1699);
nor U3020 (N_3020,N_863,N_472);
nor U3021 (N_3021,N_1718,N_980);
xor U3022 (N_3022,N_2468,N_173);
nand U3023 (N_3023,N_1071,N_2452);
and U3024 (N_3024,N_1758,N_2409);
xnor U3025 (N_3025,N_2589,N_2673);
nand U3026 (N_3026,N_2364,N_24);
or U3027 (N_3027,N_65,N_1149);
or U3028 (N_3028,N_2712,N_476);
nand U3029 (N_3029,N_1807,N_436);
and U3030 (N_3030,N_2008,N_855);
nor U3031 (N_3031,N_2996,N_2318);
or U3032 (N_3032,N_1714,N_2513);
nor U3033 (N_3033,N_2463,N_1617);
and U3034 (N_3034,N_338,N_825);
and U3035 (N_3035,N_1382,N_149);
or U3036 (N_3036,N_502,N_1402);
and U3037 (N_3037,N_2411,N_1519);
and U3038 (N_3038,N_2765,N_2035);
nand U3039 (N_3039,N_2439,N_1683);
and U3040 (N_3040,N_2789,N_1533);
or U3041 (N_3041,N_2803,N_2685);
xor U3042 (N_3042,N_928,N_1586);
nor U3043 (N_3043,N_1443,N_990);
xnor U3044 (N_3044,N_591,N_1206);
nor U3045 (N_3045,N_77,N_90);
nand U3046 (N_3046,N_831,N_2984);
nand U3047 (N_3047,N_1272,N_2370);
nor U3048 (N_3048,N_2290,N_2948);
and U3049 (N_3049,N_797,N_1589);
and U3050 (N_3050,N_2961,N_2638);
or U3051 (N_3051,N_1906,N_2330);
nand U3052 (N_3052,N_346,N_2316);
nor U3053 (N_3053,N_2098,N_1258);
and U3054 (N_3054,N_849,N_1893);
nor U3055 (N_3055,N_975,N_76);
and U3056 (N_3056,N_1313,N_1774);
and U3057 (N_3057,N_2988,N_2737);
or U3058 (N_3058,N_2271,N_735);
nor U3059 (N_3059,N_2166,N_1090);
nand U3060 (N_3060,N_2197,N_538);
nor U3061 (N_3061,N_36,N_1359);
nor U3062 (N_3062,N_2480,N_2103);
and U3063 (N_3063,N_1394,N_1963);
and U3064 (N_3064,N_1116,N_193);
nor U3065 (N_3065,N_1542,N_456);
and U3066 (N_3066,N_2628,N_1994);
nor U3067 (N_3067,N_2847,N_2857);
nor U3068 (N_3068,N_7,N_867);
nand U3069 (N_3069,N_1596,N_1870);
nor U3070 (N_3070,N_2057,N_957);
nand U3071 (N_3071,N_2598,N_1876);
xor U3072 (N_3072,N_489,N_2011);
nand U3073 (N_3073,N_1932,N_1562);
xor U3074 (N_3074,N_231,N_1161);
nand U3075 (N_3075,N_788,N_2042);
nand U3076 (N_3076,N_2587,N_2667);
and U3077 (N_3077,N_542,N_762);
or U3078 (N_3078,N_1177,N_1500);
or U3079 (N_3079,N_195,N_1559);
xnor U3080 (N_3080,N_2656,N_21);
nor U3081 (N_3081,N_530,N_471);
or U3082 (N_3082,N_2865,N_445);
nand U3083 (N_3083,N_356,N_2753);
xnor U3084 (N_3084,N_1093,N_2939);
and U3085 (N_3085,N_2503,N_1254);
xnor U3086 (N_3086,N_1358,N_1713);
and U3087 (N_3087,N_903,N_2641);
and U3088 (N_3088,N_1777,N_2297);
nand U3089 (N_3089,N_2395,N_194);
or U3090 (N_3090,N_2819,N_135);
or U3091 (N_3091,N_847,N_1340);
nor U3092 (N_3092,N_2822,N_1631);
and U3093 (N_3093,N_1001,N_441);
nand U3094 (N_3094,N_2791,N_1334);
or U3095 (N_3095,N_2029,N_612);
or U3096 (N_3096,N_1776,N_104);
nand U3097 (N_3097,N_2474,N_954);
xnor U3098 (N_3098,N_2666,N_1775);
xnor U3099 (N_3099,N_2684,N_1998);
xnor U3100 (N_3100,N_2894,N_937);
nor U3101 (N_3101,N_1086,N_820);
or U3102 (N_3102,N_1860,N_2698);
nor U3103 (N_3103,N_1499,N_1987);
nand U3104 (N_3104,N_1634,N_1045);
xor U3105 (N_3105,N_1233,N_2112);
nor U3106 (N_3106,N_1951,N_508);
or U3107 (N_3107,N_2921,N_1377);
and U3108 (N_3108,N_1689,N_682);
nor U3109 (N_3109,N_2911,N_1305);
or U3110 (N_3110,N_1407,N_2888);
nor U3111 (N_3111,N_1772,N_2848);
nor U3112 (N_3112,N_2728,N_1386);
nand U3113 (N_3113,N_335,N_386);
or U3114 (N_3114,N_1194,N_659);
nand U3115 (N_3115,N_2385,N_2289);
nor U3116 (N_3116,N_465,N_1761);
xor U3117 (N_3117,N_1320,N_1477);
or U3118 (N_3118,N_1024,N_2863);
xor U3119 (N_3119,N_2623,N_2209);
xor U3120 (N_3120,N_306,N_138);
xnor U3121 (N_3121,N_1770,N_492);
and U3122 (N_3122,N_2640,N_1196);
xor U3123 (N_3123,N_2399,N_1605);
xnor U3124 (N_3124,N_2373,N_2975);
nand U3125 (N_3125,N_527,N_2823);
and U3126 (N_3126,N_1960,N_1250);
xnor U3127 (N_3127,N_2947,N_600);
xor U3128 (N_3128,N_1120,N_2950);
and U3129 (N_3129,N_1434,N_683);
nor U3130 (N_3130,N_948,N_2251);
or U3131 (N_3131,N_1995,N_1773);
and U3132 (N_3132,N_1855,N_731);
xor U3133 (N_3133,N_1041,N_2146);
or U3134 (N_3134,N_2945,N_1642);
or U3135 (N_3135,N_2635,N_1907);
nand U3136 (N_3136,N_2647,N_2);
and U3137 (N_3137,N_1240,N_1370);
or U3138 (N_3138,N_2760,N_1975);
and U3139 (N_3139,N_1084,N_2982);
nand U3140 (N_3140,N_1193,N_434);
and U3141 (N_3141,N_2884,N_1989);
nor U3142 (N_3142,N_1676,N_1174);
and U3143 (N_3143,N_340,N_2683);
nand U3144 (N_3144,N_544,N_866);
nand U3145 (N_3145,N_75,N_1417);
xor U3146 (N_3146,N_1447,N_2198);
or U3147 (N_3147,N_536,N_1208);
or U3148 (N_3148,N_2787,N_1216);
and U3149 (N_3149,N_1278,N_171);
xnor U3150 (N_3150,N_56,N_2481);
or U3151 (N_3151,N_2036,N_2979);
or U3152 (N_3152,N_247,N_2438);
and U3153 (N_3153,N_661,N_1523);
or U3154 (N_3154,N_27,N_1037);
xor U3155 (N_3155,N_1003,N_1551);
nand U3156 (N_3156,N_505,N_2000);
nand U3157 (N_3157,N_42,N_2580);
nor U3158 (N_3158,N_353,N_2958);
and U3159 (N_3159,N_933,N_1748);
and U3160 (N_3160,N_1652,N_47);
or U3161 (N_3161,N_710,N_2799);
nand U3162 (N_3162,N_1114,N_2985);
xnor U3163 (N_3163,N_1362,N_1460);
or U3164 (N_3164,N_2779,N_641);
or U3165 (N_3165,N_303,N_758);
xor U3166 (N_3166,N_1913,N_2875);
nand U3167 (N_3167,N_1481,N_1685);
or U3168 (N_3168,N_981,N_1843);
nand U3169 (N_3169,N_2956,N_1808);
nand U3170 (N_3170,N_1701,N_1673);
xor U3171 (N_3171,N_1124,N_2949);
nand U3172 (N_3172,N_533,N_2167);
xnor U3173 (N_3173,N_1669,N_1482);
and U3174 (N_3174,N_110,N_776);
nor U3175 (N_3175,N_923,N_460);
nand U3176 (N_3176,N_2158,N_2567);
xnor U3177 (N_3177,N_677,N_537);
and U3178 (N_3178,N_501,N_2778);
xnor U3179 (N_3179,N_1075,N_332);
nor U3180 (N_3180,N_1346,N_1502);
nor U3181 (N_3181,N_2601,N_1217);
nand U3182 (N_3182,N_1971,N_1762);
or U3183 (N_3183,N_575,N_2994);
or U3184 (N_3184,N_2187,N_2590);
and U3185 (N_3185,N_385,N_2274);
nand U3186 (N_3186,N_2637,N_917);
and U3187 (N_3187,N_2755,N_1740);
or U3188 (N_3188,N_1841,N_2960);
and U3189 (N_3189,N_187,N_2585);
and U3190 (N_3190,N_1722,N_1328);
and U3191 (N_3191,N_2649,N_410);
and U3192 (N_3192,N_2957,N_1736);
or U3193 (N_3193,N_1092,N_2573);
nand U3194 (N_3194,N_1029,N_918);
xnor U3195 (N_3195,N_1503,N_1743);
nand U3196 (N_3196,N_2471,N_1085);
nor U3197 (N_3197,N_1485,N_2164);
and U3198 (N_3198,N_1224,N_2866);
nor U3199 (N_3199,N_1473,N_2082);
or U3200 (N_3200,N_1663,N_1547);
nor U3201 (N_3201,N_2138,N_2172);
xnor U3202 (N_3202,N_848,N_2804);
xnor U3203 (N_3203,N_657,N_2044);
nor U3204 (N_3204,N_2278,N_163);
or U3205 (N_3205,N_2786,N_1506);
nand U3206 (N_3206,N_159,N_2929);
xnor U3207 (N_3207,N_404,N_1857);
nor U3208 (N_3208,N_794,N_1077);
nand U3209 (N_3209,N_801,N_2296);
and U3210 (N_3210,N_2052,N_2389);
or U3211 (N_3211,N_2615,N_111);
nand U3212 (N_3212,N_771,N_2018);
xnor U3213 (N_3213,N_277,N_2837);
and U3214 (N_3214,N_1815,N_2930);
nor U3215 (N_3215,N_2259,N_580);
nand U3216 (N_3216,N_1046,N_905);
nand U3217 (N_3217,N_275,N_684);
xor U3218 (N_3218,N_1798,N_2361);
nand U3219 (N_3219,N_2340,N_550);
or U3220 (N_3220,N_2499,N_1536);
nor U3221 (N_3221,N_2441,N_930);
or U3222 (N_3222,N_1779,N_2342);
and U3223 (N_3223,N_1170,N_1795);
and U3224 (N_3224,N_1099,N_2379);
nor U3225 (N_3225,N_1865,N_2420);
or U3226 (N_3226,N_1204,N_2719);
or U3227 (N_3227,N_2771,N_642);
or U3228 (N_3228,N_2695,N_2030);
xor U3229 (N_3229,N_1791,N_1323);
and U3230 (N_3230,N_209,N_2506);
nor U3231 (N_3231,N_1164,N_1052);
and U3232 (N_3232,N_941,N_1730);
nor U3233 (N_3233,N_510,N_1577);
or U3234 (N_3234,N_245,N_1805);
xor U3235 (N_3235,N_992,N_2725);
or U3236 (N_3236,N_1273,N_254);
and U3237 (N_3237,N_1212,N_1471);
nand U3238 (N_3238,N_2552,N_2091);
or U3239 (N_3239,N_972,N_1138);
or U3240 (N_3240,N_963,N_2286);
nand U3241 (N_3241,N_1719,N_126);
or U3242 (N_3242,N_973,N_2045);
xnor U3243 (N_3243,N_223,N_1476);
nand U3244 (N_3244,N_2898,N_1988);
and U3245 (N_3245,N_1329,N_2727);
xor U3246 (N_3246,N_2225,N_773);
xnor U3247 (N_3247,N_1575,N_480);
or U3248 (N_3248,N_2969,N_1168);
nor U3249 (N_3249,N_1658,N_705);
or U3250 (N_3250,N_2494,N_541);
and U3251 (N_3251,N_547,N_2536);
and U3252 (N_3252,N_1427,N_1060);
nand U3253 (N_3253,N_2740,N_2015);
nand U3254 (N_3254,N_2636,N_1708);
xnor U3255 (N_3255,N_2242,N_1784);
nor U3256 (N_3256,N_1629,N_2664);
and U3257 (N_3257,N_1432,N_2759);
xnor U3258 (N_3258,N_1842,N_2264);
nand U3259 (N_3259,N_2610,N_1526);
or U3260 (N_3260,N_572,N_287);
or U3261 (N_3261,N_1552,N_1871);
and U3262 (N_3262,N_1896,N_2665);
and U3263 (N_3263,N_674,N_131);
nand U3264 (N_3264,N_2106,N_1429);
nand U3265 (N_3265,N_141,N_74);
xnor U3266 (N_3266,N_217,N_1065);
or U3267 (N_3267,N_152,N_1771);
nor U3268 (N_3268,N_1091,N_802);
and U3269 (N_3269,N_164,N_1826);
xor U3270 (N_3270,N_1211,N_391);
nor U3271 (N_3271,N_2206,N_92);
or U3272 (N_3272,N_1244,N_2696);
xnor U3273 (N_3273,N_2801,N_2566);
or U3274 (N_3274,N_678,N_939);
xor U3275 (N_3275,N_724,N_2191);
xnor U3276 (N_3276,N_886,N_1767);
and U3277 (N_3277,N_162,N_2903);
nor U3278 (N_3278,N_219,N_1438);
nand U3279 (N_3279,N_1919,N_1933);
or U3280 (N_3280,N_2137,N_694);
nand U3281 (N_3281,N_592,N_2055);
and U3282 (N_3282,N_1668,N_2016);
and U3283 (N_3283,N_174,N_2851);
nand U3284 (N_3284,N_419,N_1264);
or U3285 (N_3285,N_1374,N_915);
xnor U3286 (N_3286,N_2764,N_718);
xnor U3287 (N_3287,N_1741,N_2889);
and U3288 (N_3288,N_619,N_321);
nor U3289 (N_3289,N_897,N_2382);
and U3290 (N_3290,N_2990,N_2999);
nor U3291 (N_3291,N_807,N_2159);
xor U3292 (N_3292,N_1293,N_2858);
nor U3293 (N_3293,N_2669,N_1709);
nor U3294 (N_3294,N_339,N_789);
or U3295 (N_3295,N_1588,N_2794);
and U3296 (N_3296,N_1534,N_1508);
xnor U3297 (N_3297,N_1215,N_2149);
nand U3298 (N_3298,N_1005,N_2378);
or U3299 (N_3299,N_1426,N_1404);
nand U3300 (N_3300,N_698,N_2273);
and U3301 (N_3301,N_2428,N_1353);
nand U3302 (N_3302,N_150,N_519);
xor U3303 (N_3303,N_1310,N_876);
nand U3304 (N_3304,N_2504,N_1984);
or U3305 (N_3305,N_979,N_967);
or U3306 (N_3306,N_875,N_2549);
and U3307 (N_3307,N_1228,N_1645);
and U3308 (N_3308,N_38,N_1889);
xnor U3309 (N_3309,N_154,N_148);
nor U3310 (N_3310,N_113,N_2592);
and U3311 (N_3311,N_1366,N_1132);
or U3312 (N_3312,N_0,N_729);
xor U3313 (N_3313,N_146,N_1375);
and U3314 (N_3314,N_1127,N_407);
and U3315 (N_3315,N_2002,N_707);
nand U3316 (N_3316,N_1840,N_2203);
xor U3317 (N_3317,N_2108,N_257);
nor U3318 (N_3318,N_2768,N_2007);
or U3319 (N_3319,N_2432,N_1861);
xnor U3320 (N_3320,N_1449,N_2092);
or U3321 (N_3321,N_37,N_2235);
and U3322 (N_3322,N_1814,N_1096);
nor U3323 (N_3323,N_2498,N_1556);
nand U3324 (N_3324,N_1104,N_669);
xor U3325 (N_3325,N_2981,N_1947);
xor U3326 (N_3326,N_1867,N_1786);
or U3327 (N_3327,N_1517,N_1627);
nand U3328 (N_3328,N_2477,N_1597);
nor U3329 (N_3329,N_934,N_670);
nand U3330 (N_3330,N_1422,N_1678);
xor U3331 (N_3331,N_1461,N_680);
and U3332 (N_3332,N_2953,N_2141);
nand U3333 (N_3333,N_1739,N_242);
nand U3334 (N_3334,N_62,N_746);
nand U3335 (N_3335,N_2562,N_1890);
xor U3336 (N_3336,N_838,N_2261);
nor U3337 (N_3337,N_25,N_1769);
nor U3338 (N_3338,N_1295,N_1760);
or U3339 (N_3339,N_2182,N_2184);
and U3340 (N_3340,N_1553,N_2998);
and U3341 (N_3341,N_1900,N_1868);
nor U3342 (N_3342,N_483,N_1630);
or U3343 (N_3343,N_1043,N_970);
xor U3344 (N_3344,N_2731,N_706);
xnor U3345 (N_3345,N_690,N_2626);
nand U3346 (N_3346,N_2815,N_986);
xnor U3347 (N_3347,N_488,N_2118);
nand U3348 (N_3348,N_1943,N_1409);
or U3349 (N_3349,N_1117,N_295);
nand U3350 (N_3350,N_1512,N_621);
xnor U3351 (N_3351,N_921,N_69);
or U3352 (N_3352,N_1557,N_668);
nor U3353 (N_3353,N_784,N_2747);
or U3354 (N_3354,N_1974,N_6);
or U3355 (N_3355,N_167,N_1756);
xnor U3356 (N_3356,N_1725,N_2588);
nand U3357 (N_3357,N_971,N_2697);
nand U3358 (N_3358,N_2232,N_1800);
nor U3359 (N_3359,N_832,N_2217);
xnor U3360 (N_3360,N_2893,N_2798);
or U3361 (N_3361,N_1569,N_1304);
nor U3362 (N_3362,N_1494,N_940);
nor U3363 (N_3363,N_568,N_123);
nor U3364 (N_3364,N_1296,N_302);
nand U3365 (N_3365,N_2693,N_463);
nand U3366 (N_3366,N_1150,N_2678);
and U3367 (N_3367,N_2927,N_1111);
nand U3368 (N_3368,N_1567,N_1372);
or U3369 (N_3369,N_2124,N_2833);
xor U3370 (N_3370,N_1700,N_271);
nor U3371 (N_3371,N_581,N_1529);
nand U3372 (N_3372,N_2745,N_2069);
xor U3373 (N_3373,N_1875,N_2021);
or U3374 (N_3374,N_80,N_1992);
or U3375 (N_3375,N_2607,N_805);
nand U3376 (N_3376,N_2408,N_108);
nand U3377 (N_3377,N_2024,N_950);
and U3378 (N_3378,N_1235,N_1821);
and U3379 (N_3379,N_1999,N_1192);
or U3380 (N_3380,N_2519,N_579);
xnor U3381 (N_3381,N_1746,N_2028);
nor U3382 (N_3382,N_2078,N_938);
and U3383 (N_3383,N_1591,N_244);
nor U3384 (N_3384,N_1931,N_1146);
xor U3385 (N_3385,N_1269,N_2020);
or U3386 (N_3386,N_1087,N_1133);
nand U3387 (N_3387,N_466,N_2133);
nand U3388 (N_3388,N_1276,N_1082);
and U3389 (N_3389,N_1766,N_310);
xnor U3390 (N_3390,N_352,N_2356);
nand U3391 (N_3391,N_2151,N_363);
or U3392 (N_3392,N_1078,N_1978);
nor U3393 (N_3393,N_1792,N_1119);
nand U3394 (N_3394,N_2565,N_314);
xor U3395 (N_3395,N_1142,N_1498);
nand U3396 (N_3396,N_212,N_2313);
nor U3397 (N_3397,N_951,N_1854);
nor U3398 (N_3398,N_2461,N_1027);
or U3399 (N_3399,N_635,N_2874);
nor U3400 (N_3400,N_474,N_2025);
or U3401 (N_3401,N_2630,N_623);
xor U3402 (N_3402,N_43,N_325);
nor U3403 (N_3403,N_761,N_415);
nand U3404 (N_3404,N_1237,N_213);
nand U3405 (N_3405,N_2951,N_2869);
xnor U3406 (N_3406,N_583,N_2258);
or U3407 (N_3407,N_2572,N_651);
and U3408 (N_3408,N_2013,N_1703);
or U3409 (N_3409,N_2663,N_2938);
nor U3410 (N_3410,N_955,N_2417);
xnor U3411 (N_3411,N_2236,N_1288);
xnor U3412 (N_3412,N_2152,N_479);
and U3413 (N_3413,N_1486,N_978);
nand U3414 (N_3414,N_473,N_85);
xnor U3415 (N_3415,N_570,N_528);
nand U3416 (N_3416,N_2834,N_214);
and U3417 (N_3417,N_1436,N_224);
nand U3418 (N_3418,N_2622,N_1007);
or U3419 (N_3419,N_1303,N_1880);
and U3420 (N_3420,N_999,N_169);
nor U3421 (N_3421,N_422,N_716);
nand U3422 (N_3422,N_1619,N_737);
xnor U3423 (N_3423,N_2897,N_1266);
nor U3424 (N_3424,N_380,N_2976);
nor U3425 (N_3425,N_2321,N_2780);
xor U3426 (N_3426,N_549,N_107);
xor U3427 (N_3427,N_1904,N_87);
and U3428 (N_3428,N_1423,N_1899);
xor U3429 (N_3429,N_1478,N_1153);
and U3430 (N_3430,N_1496,N_1925);
or U3431 (N_3431,N_298,N_861);
and U3432 (N_3432,N_220,N_1845);
and U3433 (N_3433,N_259,N_1459);
nand U3434 (N_3434,N_1381,N_1229);
and U3435 (N_3435,N_1661,N_2776);
or U3436 (N_3436,N_2447,N_1525);
nor U3437 (N_3437,N_839,N_1797);
nor U3438 (N_3438,N_1582,N_4);
and U3439 (N_3439,N_145,N_2129);
nand U3440 (N_3440,N_276,N_879);
or U3441 (N_3441,N_2136,N_1245);
nand U3442 (N_3442,N_2658,N_2234);
and U3443 (N_3443,N_1162,N_2061);
nor U3444 (N_3444,N_1163,N_114);
and U3445 (N_3445,N_631,N_2469);
and U3446 (N_3446,N_1479,N_343);
or U3447 (N_3447,N_478,N_714);
nand U3448 (N_3448,N_1,N_318);
and U3449 (N_3449,N_723,N_2270);
nor U3450 (N_3450,N_2703,N_1284);
xnor U3451 (N_3451,N_2034,N_186);
nand U3452 (N_3452,N_136,N_2102);
or U3453 (N_3453,N_1316,N_1872);
xor U3454 (N_3454,N_1950,N_2966);
or U3455 (N_3455,N_2769,N_2909);
and U3456 (N_3456,N_2292,N_2967);
nor U3457 (N_3457,N_1360,N_2721);
nor U3458 (N_3458,N_1016,N_82);
or U3459 (N_3459,N_618,N_2328);
nand U3460 (N_3460,N_2551,N_2933);
xnor U3461 (N_3461,N_1414,N_362);
xor U3462 (N_3462,N_139,N_850);
nand U3463 (N_3463,N_2180,N_2459);
xor U3464 (N_3464,N_1189,N_402);
or U3465 (N_3465,N_2320,N_3);
nor U3466 (N_3466,N_543,N_1727);
or U3467 (N_3467,N_499,N_1607);
and U3468 (N_3468,N_1910,N_2424);
nor U3469 (N_3469,N_413,N_2691);
xor U3470 (N_3470,N_300,N_359);
xnor U3471 (N_3471,N_234,N_2827);
xor U3472 (N_3472,N_1368,N_222);
xnor U3473 (N_3473,N_882,N_486);
and U3474 (N_3474,N_1696,N_2606);
nor U3475 (N_3475,N_2841,N_1225);
or U3476 (N_3476,N_1232,N_431);
nand U3477 (N_3477,N_1458,N_2767);
nor U3478 (N_3478,N_2609,N_382);
nand U3479 (N_3479,N_726,N_1834);
xnor U3480 (N_3480,N_665,N_1241);
xor U3481 (N_3481,N_1579,N_991);
nor U3482 (N_3482,N_2808,N_2229);
and U3483 (N_3483,N_2742,N_2039);
and U3484 (N_3484,N_1307,N_1641);
or U3485 (N_3485,N_250,N_1892);
nand U3486 (N_3486,N_2563,N_1465);
and U3487 (N_3487,N_17,N_835);
xnor U3488 (N_3488,N_1956,N_34);
and U3489 (N_3489,N_304,N_1935);
or U3490 (N_3490,N_2971,N_889);
xor U3491 (N_3491,N_215,N_988);
nor U3492 (N_3492,N_317,N_365);
or U3493 (N_3493,N_299,N_2375);
or U3494 (N_3494,N_1524,N_1330);
and U3495 (N_3495,N_2047,N_1176);
nand U3496 (N_3496,N_1181,N_2741);
xnor U3497 (N_3497,N_2524,N_1594);
xor U3498 (N_3498,N_2816,N_2632);
nor U3499 (N_3499,N_1603,N_305);
nand U3500 (N_3500,N_686,N_1081);
nor U3501 (N_3501,N_2022,N_2970);
nand U3502 (N_3502,N_2688,N_1564);
nor U3503 (N_3503,N_1986,N_2633);
xnor U3504 (N_3504,N_1306,N_1757);
xnor U3505 (N_3505,N_2281,N_1953);
xor U3506 (N_3506,N_2301,N_1014);
and U3507 (N_3507,N_1321,N_1539);
or U3508 (N_3508,N_1869,N_697);
and U3509 (N_3509,N_578,N_2781);
and U3510 (N_3510,N_1924,N_2305);
or U3511 (N_3511,N_2489,N_673);
nand U3512 (N_3512,N_1022,N_2390);
and U3513 (N_3513,N_559,N_1744);
nor U3514 (N_3514,N_2730,N_1555);
and U3515 (N_3515,N_1692,N_324);
or U3516 (N_3516,N_1812,N_1625);
or U3517 (N_3517,N_2168,N_2879);
xor U3518 (N_3518,N_1231,N_1961);
nor U3519 (N_3519,N_2690,N_2491);
xnor U3520 (N_3520,N_2360,N_573);
nand U3521 (N_3521,N_1497,N_2449);
nand U3522 (N_3522,N_522,N_2299);
xnor U3523 (N_3523,N_1101,N_2702);
nor U3524 (N_3524,N_129,N_2357);
nor U3525 (N_3525,N_640,N_2774);
nand U3526 (N_3526,N_112,N_1356);
xnor U3527 (N_3527,N_2995,N_1159);
nand U3528 (N_3528,N_1723,N_2599);
xnor U3529 (N_3529,N_1421,N_1079);
xor U3530 (N_3530,N_2377,N_2226);
xnor U3531 (N_3531,N_2422,N_2818);
xor U3532 (N_3532,N_2132,N_122);
nor U3533 (N_3533,N_1347,N_1469);
nand U3534 (N_3534,N_2048,N_1822);
nor U3535 (N_3535,N_688,N_2944);
and U3536 (N_3536,N_2277,N_2005);
nor U3537 (N_3537,N_2096,N_1660);
nor U3538 (N_3538,N_253,N_2388);
nor U3539 (N_3539,N_2618,N_2196);
nor U3540 (N_3540,N_1672,N_1350);
xor U3541 (N_3541,N_1702,N_2070);
or U3542 (N_3542,N_2201,N_634);
or U3543 (N_3543,N_2973,N_2051);
nand U3544 (N_3544,N_1887,N_2269);
xor U3545 (N_3545,N_1682,N_2541);
xnor U3546 (N_3546,N_2031,N_2932);
and U3547 (N_3547,N_685,N_1884);
xor U3548 (N_3548,N_2298,N_996);
nor U3549 (N_3549,N_2363,N_1056);
xor U3550 (N_3550,N_2899,N_294);
or U3551 (N_3551,N_2396,N_1712);
nor U3552 (N_3552,N_1018,N_1435);
and U3553 (N_3553,N_770,N_177);
nand U3554 (N_3554,N_2415,N_115);
or U3555 (N_3555,N_2413,N_748);
nand U3556 (N_3556,N_349,N_2579);
xor U3557 (N_3557,N_2294,N_2066);
xor U3558 (N_3558,N_912,N_1352);
nand U3559 (N_3559,N_2306,N_1126);
nor U3560 (N_3560,N_520,N_412);
or U3561 (N_3561,N_319,N_2935);
nand U3562 (N_3562,N_828,N_741);
or U3563 (N_3563,N_1238,N_1369);
and U3564 (N_3564,N_1903,N_2528);
or U3565 (N_3565,N_1268,N_2220);
or U3566 (N_3566,N_795,N_1728);
nand U3567 (N_3567,N_567,N_200);
and U3568 (N_3568,N_1311,N_2716);
nand U3569 (N_3569,N_1622,N_392);
nand U3570 (N_3570,N_511,N_1187);
nor U3571 (N_3571,N_1501,N_233);
or U3572 (N_3572,N_2881,N_808);
or U3573 (N_3573,N_2161,N_2941);
nor U3574 (N_3574,N_83,N_2861);
xor U3575 (N_3575,N_2809,N_2531);
or U3576 (N_3576,N_2896,N_2578);
or U3577 (N_3577,N_920,N_2919);
nand U3578 (N_3578,N_2775,N_671);
nor U3579 (N_3579,N_2813,N_449);
or U3580 (N_3580,N_1681,N_496);
xnor U3581 (N_3581,N_374,N_2123);
nand U3582 (N_3582,N_1612,N_1926);
nand U3583 (N_3583,N_2853,N_1613);
and U3584 (N_3584,N_2105,N_1157);
nor U3585 (N_3585,N_2228,N_1796);
nor U3586 (N_3586,N_2800,N_961);
or U3587 (N_3587,N_475,N_72);
nor U3588 (N_3588,N_806,N_1862);
nand U3589 (N_3589,N_2111,N_1788);
and U3590 (N_3590,N_822,N_1160);
and U3591 (N_3591,N_2165,N_258);
nand U3592 (N_3592,N_2405,N_1537);
nand U3593 (N_3593,N_1484,N_367);
nor U3594 (N_3594,N_2348,N_2777);
nor U3595 (N_3595,N_1028,N_985);
xor U3596 (N_3596,N_2462,N_2868);
nor U3597 (N_3597,N_2761,N_312);
and U3598 (N_3598,N_629,N_1970);
nor U3599 (N_3599,N_814,N_1948);
and U3600 (N_3600,N_5,N_1694);
or U3601 (N_3601,N_1839,N_763);
nand U3602 (N_3602,N_589,N_1034);
and U3603 (N_3603,N_1076,N_1566);
xnor U3604 (N_3604,N_874,N_1637);
nand U3605 (N_3605,N_2131,N_11);
nor U3606 (N_3606,N_2337,N_1580);
nor U3607 (N_3607,N_1643,N_2338);
xnor U3608 (N_3608,N_1518,N_1859);
nand U3609 (N_3609,N_2546,N_2279);
or U3610 (N_3610,N_2247,N_387);
or U3611 (N_3611,N_846,N_400);
and U3612 (N_3612,N_2421,N_1050);
or U3613 (N_3613,N_1333,N_1452);
or U3614 (N_3614,N_2545,N_255);
or U3615 (N_3615,N_1125,N_403);
xor U3616 (N_3616,N_218,N_836);
and U3617 (N_3617,N_1015,N_1399);
or U3618 (N_3618,N_2317,N_1389);
nor U3619 (N_3619,N_908,N_1520);
xor U3620 (N_3620,N_2358,N_1314);
nand U3621 (N_3621,N_790,N_1799);
or U3622 (N_3622,N_896,N_2748);
nand U3623 (N_3623,N_2547,N_30);
nand U3624 (N_3624,N_1136,N_2181);
or U3625 (N_3625,N_2355,N_892);
and U3626 (N_3626,N_261,N_394);
and U3627 (N_3627,N_1008,N_1972);
and U3628 (N_3628,N_2064,N_566);
or U3629 (N_3629,N_834,N_1705);
nor U3630 (N_3630,N_1349,N_2586);
nor U3631 (N_3631,N_1590,N_2918);
and U3632 (N_3632,N_1207,N_2650);
or U3633 (N_3633,N_1033,N_2522);
nor U3634 (N_3634,N_2817,N_2071);
xor U3635 (N_3635,N_2351,N_2176);
nor U3636 (N_3636,N_1653,N_411);
or U3637 (N_3637,N_749,N_59);
and U3638 (N_3638,N_490,N_1558);
nor U3639 (N_3639,N_2826,N_1089);
or U3640 (N_3640,N_1437,N_1973);
xnor U3641 (N_3641,N_1595,N_311);
nor U3642 (N_3642,N_2726,N_1069);
nand U3643 (N_3643,N_482,N_2686);
nor U3644 (N_3644,N_1270,N_638);
nor U3645 (N_3645,N_498,N_1837);
and U3646 (N_3646,N_652,N_1665);
nand U3647 (N_3647,N_1249,N_1068);
or U3648 (N_3648,N_2795,N_221);
or U3649 (N_3649,N_1420,N_1094);
and U3650 (N_3650,N_2457,N_1809);
nor U3651 (N_3651,N_2620,N_2910);
or U3652 (N_3652,N_1764,N_2644);
nand U3653 (N_3653,N_1415,N_891);
and U3654 (N_3654,N_1783,N_2214);
nor U3655 (N_3655,N_1451,N_2877);
nand U3656 (N_3656,N_2308,N_226);
nor U3657 (N_3657,N_2193,N_1095);
or U3658 (N_3658,N_2033,N_190);
nand U3659 (N_3659,N_1794,N_1309);
nor U3660 (N_3660,N_1810,N_901);
or U3661 (N_3661,N_1098,N_2451);
nor U3662 (N_3662,N_1624,N_1532);
nor U3663 (N_3663,N_1711,N_1403);
nand U3664 (N_3664,N_2347,N_2194);
and U3665 (N_3665,N_320,N_35);
nor U3666 (N_3666,N_1491,N_1178);
nor U3667 (N_3667,N_1656,N_931);
nand U3668 (N_3668,N_633,N_627);
xor U3669 (N_3669,N_1921,N_1325);
or U3670 (N_3670,N_288,N_286);
nand U3671 (N_3671,N_2754,N_2104);
or U3672 (N_3672,N_1707,N_2694);
and U3673 (N_3673,N_15,N_2864);
nand U3674 (N_3674,N_2593,N_1010);
xnor U3675 (N_3675,N_109,N_1298);
and U3676 (N_3676,N_2230,N_2386);
or U3677 (N_3677,N_2085,N_1410);
nor U3678 (N_3678,N_2668,N_468);
and U3679 (N_3679,N_610,N_1522);
or U3680 (N_3680,N_1059,N_2521);
nor U3681 (N_3681,N_662,N_399);
nor U3682 (N_3682,N_1747,N_1985);
or U3683 (N_3683,N_134,N_1717);
nand U3684 (N_3684,N_1444,N_2806);
and U3685 (N_3685,N_922,N_2989);
and U3686 (N_3686,N_1874,N_949);
nor U3687 (N_3687,N_1376,N_9);
and U3688 (N_3688,N_2796,N_952);
and U3689 (N_3689,N_1275,N_622);
xor U3690 (N_3690,N_2365,N_1401);
or U3691 (N_3691,N_230,N_2450);
nand U3692 (N_3692,N_1470,N_2574);
or U3693 (N_3693,N_2992,N_426);
xor U3694 (N_3694,N_1934,N_1286);
and U3695 (N_3695,N_2001,N_256);
nor U3696 (N_3696,N_66,N_2614);
or U3697 (N_3697,N_736,N_144);
xor U3698 (N_3698,N_2746,N_1221);
or U3699 (N_3699,N_1930,N_2842);
and U3700 (N_3700,N_333,N_2639);
nand U3701 (N_3701,N_2429,N_1413);
nand U3702 (N_3702,N_2419,N_354);
and U3703 (N_3703,N_347,N_2117);
xnor U3704 (N_3704,N_944,N_58);
nand U3705 (N_3705,N_757,N_1592);
and U3706 (N_3706,N_1521,N_778);
nand U3707 (N_3707,N_1070,N_2516);
xnor U3708 (N_3708,N_2917,N_243);
nor U3709 (N_3709,N_557,N_249);
or U3710 (N_3710,N_2063,N_2525);
nand U3711 (N_3711,N_2605,N_2772);
xor U3712 (N_3712,N_2397,N_1445);
nor U3713 (N_3713,N_2752,N_2445);
or U3714 (N_3714,N_2253,N_2115);
xor U3715 (N_3715,N_1733,N_444);
xor U3716 (N_3716,N_10,N_1549);
xor U3717 (N_3717,N_1103,N_101);
nand U3718 (N_3718,N_2568,N_2502);
xor U3719 (N_3719,N_1246,N_361);
and U3720 (N_3720,N_2237,N_2553);
nor U3721 (N_3721,N_2006,N_1844);
and U3722 (N_3722,N_1324,N_1493);
nor U3723 (N_3723,N_2325,N_2505);
nor U3724 (N_3724,N_2706,N_1688);
and U3725 (N_3725,N_2260,N_709);
xor U3726 (N_3726,N_2488,N_1729);
nand U3727 (N_3727,N_796,N_2770);
or U3728 (N_3728,N_817,N_1543);
nor U3729 (N_3729,N_1019,N_2793);
nand U3730 (N_3730,N_1327,N_791);
and U3731 (N_3731,N_2431,N_157);
nand U3732 (N_3732,N_906,N_608);
and U3733 (N_3733,N_624,N_1055);
and U3734 (N_3734,N_379,N_526);
and U3735 (N_3735,N_1639,N_1632);
and U3736 (N_3736,N_2571,N_1039);
or U3737 (N_3737,N_1662,N_1336);
xor U3738 (N_3738,N_2376,N_2211);
nand U3739 (N_3739,N_1223,N_1186);
xnor U3740 (N_3740,N_2792,N_1628);
or U3741 (N_3741,N_160,N_2095);
nand U3742 (N_3742,N_2475,N_158);
nor U3743 (N_3743,N_296,N_1430);
xor U3744 (N_3744,N_2812,N_1823);
nand U3745 (N_3745,N_987,N_2402);
nand U3746 (N_3746,N_695,N_1049);
nor U3747 (N_3747,N_643,N_1431);
nand U3748 (N_3748,N_216,N_1690);
or U3749 (N_3749,N_119,N_2946);
xnor U3750 (N_3750,N_556,N_1243);
xor U3751 (N_3751,N_998,N_2974);
xnor U3752 (N_3752,N_603,N_1023);
nand U3753 (N_3753,N_650,N_598);
xnor U3754 (N_3754,N_943,N_1490);
nor U3755 (N_3755,N_1380,N_1140);
and U3756 (N_3756,N_2750,N_2501);
or U3757 (N_3757,N_2150,N_653);
nand U3758 (N_3758,N_237,N_1545);
xnor U3759 (N_3759,N_2624,N_2878);
xnor U3760 (N_3760,N_960,N_364);
nand U3761 (N_3761,N_1650,N_1337);
xnor U3762 (N_3762,N_2762,N_18);
xor U3763 (N_3763,N_2178,N_1863);
nand U3764 (N_3764,N_1297,N_628);
nor U3765 (N_3765,N_2336,N_916);
xor U3766 (N_3766,N_1040,N_2179);
xor U3767 (N_3767,N_878,N_1918);
nand U3768 (N_3768,N_2074,N_1287);
nor U3769 (N_3769,N_2401,N_2266);
xor U3770 (N_3770,N_2671,N_265);
or U3771 (N_3771,N_1236,N_974);
xnor U3772 (N_3772,N_548,N_2244);
or U3773 (N_3773,N_2583,N_211);
or U3774 (N_3774,N_2964,N_94);
xnor U3775 (N_3775,N_2241,N_1790);
or U3776 (N_3776,N_2148,N_798);
nor U3777 (N_3777,N_648,N_712);
and U3778 (N_3778,N_1013,N_515);
xnor U3779 (N_3779,N_1198,N_826);
and U3780 (N_3780,N_416,N_611);
and U3781 (N_3781,N_1914,N_2043);
nand U3782 (N_3782,N_739,N_2680);
and U3783 (N_3783,N_997,N_2423);
nor U3784 (N_3784,N_2613,N_595);
xnor U3785 (N_3785,N_2470,N_782);
and U3786 (N_3786,N_1067,N_2559);
nand U3787 (N_3787,N_308,N_143);
nor U3788 (N_3788,N_1222,N_2739);
and U3789 (N_3789,N_481,N_2219);
nor U3790 (N_3790,N_2262,N_1883);
nor U3791 (N_3791,N_2075,N_2440);
or U3792 (N_3792,N_1428,N_2256);
or U3793 (N_3793,N_602,N_1137);
nand U3794 (N_3794,N_1554,N_983);
and U3795 (N_3795,N_540,N_663);
nand U3796 (N_3796,N_2157,N_2537);
or U3797 (N_3797,N_977,N_1516);
xor U3798 (N_3798,N_1749,N_282);
xnor U3799 (N_3799,N_140,N_512);
nor U3800 (N_3800,N_2681,N_1446);
nor U3801 (N_3801,N_389,N_485);
xnor U3802 (N_3802,N_1937,N_2891);
xnor U3803 (N_3803,N_2962,N_646);
or U3804 (N_3804,N_590,N_2192);
nand U3805 (N_3805,N_1183,N_1341);
and U3806 (N_3806,N_647,N_2189);
xor U3807 (N_3807,N_1280,N_1693);
or U3808 (N_3808,N_443,N_760);
nor U3809 (N_3809,N_438,N_274);
xor U3810 (N_3810,N_232,N_1113);
nand U3811 (N_3811,N_285,N_535);
and U3812 (N_3812,N_1818,N_2876);
nor U3813 (N_3813,N_1219,N_1102);
nor U3814 (N_3814,N_2341,N_2084);
xor U3815 (N_3815,N_1393,N_180);
nand U3816 (N_3816,N_368,N_2050);
and U3817 (N_3817,N_366,N_2332);
or U3818 (N_3818,N_430,N_1695);
or U3819 (N_3819,N_2173,N_2856);
and U3820 (N_3820,N_2362,N_1317);
or U3821 (N_3821,N_28,N_1513);
and U3822 (N_3822,N_1509,N_1574);
nor U3823 (N_3823,N_484,N_1123);
nor U3824 (N_3824,N_344,N_2472);
and U3825 (N_3825,N_252,N_1200);
and U3826 (N_3826,N_843,N_48);
and U3827 (N_3827,N_2003,N_2072);
xor U3828 (N_3828,N_2497,N_2602);
or U3829 (N_3829,N_869,N_117);
nand U3830 (N_3830,N_2940,N_2843);
nand U3831 (N_3831,N_2883,N_2544);
or U3832 (N_3832,N_995,N_1466);
xnor U3833 (N_3833,N_281,N_837);
nor U3834 (N_3834,N_830,N_2079);
nand U3835 (N_3835,N_1515,N_125);
nor U3836 (N_3836,N_57,N_1185);
xnor U3837 (N_3837,N_636,N_2067);
and U3838 (N_3838,N_1940,N_14);
xnor U3839 (N_3839,N_956,N_2643);
nand U3840 (N_3840,N_2617,N_2710);
or U3841 (N_3841,N_2090,N_500);
nor U3842 (N_3842,N_676,N_2557);
and U3843 (N_3843,N_1129,N_585);
xnor U3844 (N_3844,N_454,N_263);
xor U3845 (N_3845,N_1959,N_730);
xnor U3846 (N_3846,N_1977,N_1671);
nor U3847 (N_3847,N_1291,N_759);
xnor U3848 (N_3848,N_2621,N_2383);
nand U3849 (N_3849,N_1121,N_334);
xor U3850 (N_3850,N_1687,N_1342);
nor U3851 (N_3851,N_1115,N_2707);
xnor U3852 (N_3852,N_2037,N_2319);
xnor U3853 (N_3853,N_2675,N_2991);
or U3854 (N_3854,N_45,N_1654);
nand U3855 (N_3855,N_2062,N_681);
xnor U3856 (N_3856,N_1938,N_330);
or U3857 (N_3857,N_1047,N_70);
nor U3858 (N_3858,N_201,N_2345);
and U3859 (N_3859,N_202,N_1560);
nand U3860 (N_3860,N_1608,N_672);
nand U3861 (N_3861,N_946,N_2604);
and U3862 (N_3862,N_1724,N_2645);
xor U3863 (N_3863,N_1858,N_1602);
nand U3864 (N_3864,N_2327,N_23);
and U3865 (N_3865,N_189,N_44);
and U3866 (N_3866,N_2394,N_507);
and U3867 (N_3867,N_534,N_1172);
xor U3868 (N_3868,N_1122,N_447);
or U3869 (N_3869,N_2724,N_2380);
nor U3870 (N_3870,N_1234,N_1540);
and U3871 (N_3871,N_1738,N_2353);
xor U3872 (N_3872,N_105,N_1915);
nor U3873 (N_3873,N_584,N_2454);
nand U3874 (N_3874,N_166,N_2916);
or U3875 (N_3875,N_711,N_1155);
nor U3876 (N_3876,N_1544,N_587);
xor U3877 (N_3877,N_2597,N_577);
or U3878 (N_3878,N_73,N_1789);
nor U3879 (N_3879,N_1209,N_2627);
and U3880 (N_3880,N_273,N_2134);
and U3881 (N_3881,N_1983,N_1621);
nand U3882 (N_3882,N_264,N_2177);
xnor U3883 (N_3883,N_96,N_1644);
and U3884 (N_3884,N_2097,N_2248);
and U3885 (N_3885,N_1199,N_1061);
nand U3886 (N_3886,N_1962,N_2384);
nor U3887 (N_3887,N_1110,N_433);
or U3888 (N_3888,N_854,N_1259);
nand U3889 (N_3889,N_2381,N_1946);
nor U3890 (N_3890,N_1604,N_2625);
nor U3891 (N_3891,N_2254,N_2514);
nand U3892 (N_3892,N_1411,N_1367);
nor U3893 (N_3893,N_227,N_1851);
and U3894 (N_3894,N_925,N_241);
and U3895 (N_3895,N_2110,N_787);
or U3896 (N_3896,N_824,N_2955);
and U3897 (N_3897,N_1755,N_1793);
nand U3898 (N_3898,N_1955,N_2523);
nand U3899 (N_3899,N_1279,N_2339);
xnor U3900 (N_3900,N_780,N_370);
nand U3901 (N_3901,N_743,N_1301);
nor U3902 (N_3902,N_1158,N_2444);
and U3903 (N_3903,N_2427,N_1804);
and U3904 (N_3904,N_2718,N_1134);
nand U3905 (N_3905,N_2285,N_2004);
and U3906 (N_3906,N_2993,N_99);
or U3907 (N_3907,N_301,N_2282);
and U3908 (N_3908,N_958,N_1475);
nand U3909 (N_3909,N_1751,N_1464);
xnor U3910 (N_3910,N_2820,N_1939);
xnor U3911 (N_3911,N_2824,N_372);
nand U3912 (N_3912,N_183,N_1895);
nor U3913 (N_3913,N_942,N_192);
xor U3914 (N_3914,N_2311,N_1848);
nand U3915 (N_3915,N_388,N_2968);
xor U3916 (N_3916,N_1051,N_2672);
nand U3917 (N_3917,N_1392,N_783);
and U3918 (N_3918,N_1816,N_328);
or U3919 (N_3919,N_1735,N_2077);
or U3920 (N_3920,N_947,N_1649);
nor U3921 (N_3921,N_2835,N_1097);
nor U3922 (N_3922,N_532,N_1384);
xor U3923 (N_3923,N_2465,N_2453);
or U3924 (N_3924,N_2651,N_342);
nand U3925 (N_3925,N_717,N_2518);
nand U3926 (N_3926,N_2662,N_1787);
nor U3927 (N_3927,N_1167,N_2619);
nand U3928 (N_3928,N_2088,N_2185);
xor U3929 (N_3929,N_1991,N_2127);
or U3930 (N_3930,N_853,N_926);
xnor U3931 (N_3931,N_316,N_1294);
nand U3932 (N_3932,N_864,N_1053);
xnor U3933 (N_3933,N_2443,N_751);
nor U3934 (N_3934,N_103,N_2926);
and U3935 (N_3935,N_1080,N_351);
nor U3936 (N_3936,N_852,N_2611);
nand U3937 (N_3937,N_2797,N_2652);
or U3938 (N_3938,N_1806,N_2280);
xor U3939 (N_3939,N_2555,N_2100);
xnor U3940 (N_3940,N_326,N_2509);
and U3941 (N_3941,N_188,N_1467);
or U3942 (N_3942,N_1252,N_1285);
xnor U3943 (N_3943,N_432,N_2125);
or U3944 (N_3944,N_607,N_1262);
or U3945 (N_3945,N_1396,N_2660);
nand U3946 (N_3946,N_754,N_1184);
nor U3947 (N_3947,N_1292,N_246);
nor U3948 (N_3948,N_378,N_982);
or U3949 (N_3949,N_206,N_2109);
nor U3950 (N_3950,N_870,N_845);
nor U3951 (N_3951,N_1828,N_2595);
nor U3952 (N_3952,N_2272,N_2344);
and U3953 (N_3953,N_283,N_40);
and U3954 (N_3954,N_297,N_1169);
nand U3955 (N_3955,N_446,N_675);
nand U3956 (N_3956,N_614,N_703);
xnor U3957 (N_3957,N_1942,N_1395);
or U3958 (N_3958,N_39,N_1944);
nand U3959 (N_3959,N_1391,N_262);
xnor U3960 (N_3960,N_2315,N_1338);
nor U3961 (N_3961,N_2223,N_1917);
nand U3962 (N_3962,N_79,N_2679);
nor U3963 (N_3963,N_68,N_1778);
nor U3964 (N_3964,N_2154,N_2811);
xor U3965 (N_3965,N_2902,N_1765);
nor U3966 (N_3966,N_2041,N_2059);
and U3967 (N_3967,N_1945,N_2543);
or U3968 (N_3968,N_1954,N_2014);
xnor U3969 (N_3969,N_2486,N_2977);
xor U3970 (N_3970,N_1128,N_2240);
or U3971 (N_3971,N_2527,N_2027);
xnor U3972 (N_3972,N_872,N_2596);
nor U3973 (N_3973,N_2163,N_2838);
nor U3974 (N_3974,N_155,N_1670);
and U3975 (N_3975,N_1378,N_810);
and U3976 (N_3976,N_1626,N_816);
xor U3977 (N_3977,N_1651,N_2268);
and U3978 (N_3978,N_1036,N_98);
xor U3979 (N_3979,N_1242,N_664);
or U3980 (N_3980,N_1267,N_2135);
and U3981 (N_3981,N_1332,N_2393);
xnor U3982 (N_3982,N_375,N_605);
xor U3983 (N_3983,N_976,N_451);
or U3984 (N_3984,N_1106,N_1021);
and U3985 (N_3985,N_1453,N_1355);
and U3986 (N_3986,N_1450,N_2682);
xnor U3987 (N_3987,N_2561,N_1472);
and U3988 (N_3988,N_1213,N_2904);
xnor U3989 (N_3989,N_2406,N_1315);
nor U3990 (N_3990,N_2263,N_327);
or U3991 (N_3991,N_833,N_1000);
and U3992 (N_3992,N_1831,N_1667);
or U3993 (N_3993,N_779,N_1335);
nor U3994 (N_3994,N_1745,N_637);
nor U3995 (N_3995,N_2101,N_197);
nor U3996 (N_3996,N_2140,N_2252);
nor U3997 (N_3997,N_902,N_2860);
xor U3998 (N_3998,N_2403,N_2081);
nor U3999 (N_3999,N_2425,N_1488);
and U4000 (N_4000,N_1424,N_461);
or U4001 (N_4001,N_269,N_1647);
and U4002 (N_4002,N_687,N_1949);
and U4003 (N_4003,N_764,N_2713);
nor U4004 (N_4004,N_2174,N_239);
xor U4005 (N_4005,N_813,N_462);
nand U4006 (N_4006,N_2307,N_2126);
nand U4007 (N_4007,N_2581,N_953);
or U4008 (N_4008,N_20,N_369);
nand U4009 (N_4009,N_2058,N_1599);
or U4010 (N_4010,N_819,N_156);
xor U4011 (N_4011,N_251,N_2446);
and U4012 (N_4012,N_654,N_1609);
and U4013 (N_4013,N_1020,N_175);
xnor U4014 (N_4014,N_450,N_1190);
nor U4015 (N_4015,N_2576,N_290);
nor U4016 (N_4016,N_398,N_1197);
and U4017 (N_4017,N_2026,N_552);
nor U4018 (N_4018,N_1339,N_1528);
or U4019 (N_4019,N_2387,N_491);
nand U4020 (N_4020,N_1017,N_2171);
xnor U4021 (N_4021,N_2122,N_1397);
nor U4022 (N_4022,N_2160,N_1388);
xor U4023 (N_4023,N_127,N_279);
and U4024 (N_4024,N_2906,N_2329);
or U4025 (N_4025,N_1251,N_545);
or U4026 (N_4026,N_1274,N_2416);
nor U4027 (N_4027,N_2560,N_2215);
nor U4028 (N_4028,N_2143,N_1282);
nor U4029 (N_4029,N_424,N_2309);
and U4030 (N_4030,N_1561,N_919);
nand U4031 (N_4031,N_1057,N_1601);
and U4032 (N_4032,N_1408,N_1780);
nand U4033 (N_4033,N_315,N_1610);
nor U4034 (N_4034,N_1143,N_179);
and U4035 (N_4035,N_2153,N_1530);
xnor U4036 (N_4036,N_574,N_777);
nor U4037 (N_4037,N_467,N_1965);
nor U4038 (N_4038,N_2923,N_910);
nand U4039 (N_4039,N_728,N_414);
nor U4040 (N_4040,N_1829,N_721);
nand U4041 (N_4041,N_2997,N_1248);
nor U4042 (N_4042,N_1261,N_1131);
and U4043 (N_4043,N_2540,N_1675);
and U4044 (N_4044,N_523,N_455);
nand U4045 (N_4045,N_2732,N_2128);
nand U4046 (N_4046,N_1721,N_2155);
nor U4047 (N_4047,N_16,N_88);
nor U4048 (N_4048,N_2199,N_13);
xor U4049 (N_4049,N_964,N_914);
nor U4050 (N_4050,N_2495,N_1916);
nor U4051 (N_4051,N_2830,N_823);
or U4052 (N_4052,N_208,N_267);
xor U4053 (N_4053,N_2407,N_1964);
nand U4054 (N_4054,N_2714,N_1171);
or U4055 (N_4055,N_1638,N_1684);
and U4056 (N_4056,N_2517,N_323);
xor U4057 (N_4057,N_1982,N_2788);
xnor U4058 (N_4058,N_336,N_2845);
nor U4059 (N_4059,N_1300,N_2068);
nand U4060 (N_4060,N_2368,N_630);
nand U4061 (N_4061,N_93,N_1659);
or U4062 (N_4062,N_401,N_2116);
nand U4063 (N_4063,N_693,N_1759);
or U4064 (N_4064,N_2019,N_1188);
xnor U4065 (N_4065,N_1898,N_1390);
nand U4066 (N_4066,N_1716,N_1173);
or U4067 (N_4067,N_2782,N_702);
xnor U4068 (N_4068,N_2239,N_196);
nand U4069 (N_4069,N_2766,N_2371);
nor U4070 (N_4070,N_2709,N_859);
and U4071 (N_4071,N_2304,N_767);
or U4072 (N_4072,N_2914,N_1265);
nor U4073 (N_4073,N_1923,N_1441);
xor U4074 (N_4074,N_1873,N_2756);
xor U4075 (N_4075,N_470,N_2200);
or U4076 (N_4076,N_2556,N_2705);
and U4077 (N_4077,N_2743,N_844);
or U4078 (N_4078,N_1996,N_1706);
xnor U4079 (N_4079,N_715,N_2701);
nand U4080 (N_4080,N_78,N_521);
or U4081 (N_4081,N_142,N_235);
xnor U4082 (N_4082,N_427,N_1606);
or U4083 (N_4083,N_2733,N_2221);
nand U4084 (N_4084,N_341,N_442);
and U4085 (N_4085,N_1455,N_1715);
nor U4086 (N_4086,N_51,N_1781);
nor U4087 (N_4087,N_1202,N_55);
or U4088 (N_4088,N_2484,N_719);
nor U4089 (N_4089,N_733,N_2744);
nor U4090 (N_4090,N_1636,N_1483);
nand U4091 (N_4091,N_2831,N_1813);
or U4092 (N_4092,N_1218,N_2009);
nand U4093 (N_4093,N_2119,N_514);
nand U4094 (N_4094,N_1677,N_1405);
or U4095 (N_4095,N_2087,N_1754);
xnor U4096 (N_4096,N_1511,N_2908);
nor U4097 (N_4097,N_1220,N_41);
and U4098 (N_4098,N_1664,N_293);
xnor U4099 (N_4099,N_371,N_2852);
nor U4100 (N_4100,N_803,N_609);
and U4101 (N_4101,N_696,N_1042);
nand U4102 (N_4102,N_1640,N_181);
nand U4103 (N_4103,N_1205,N_596);
nand U4104 (N_4104,N_1398,N_2139);
or U4105 (N_4105,N_2900,N_1803);
and U4106 (N_4106,N_266,N_2548);
or U4107 (N_4107,N_616,N_615);
xor U4108 (N_4108,N_2986,N_851);
nand U4109 (N_4109,N_8,N_2629);
nand U4110 (N_4110,N_2392,N_2616);
or U4111 (N_4111,N_1038,N_2757);
and U4112 (N_4112,N_184,N_2677);
and U4113 (N_4113,N_2825,N_1002);
and U4114 (N_4114,N_2145,N_1958);
or U4115 (N_4115,N_383,N_2335);
nand U4116 (N_4116,N_1928,N_1952);
nor U4117 (N_4117,N_1570,N_420);
and U4118 (N_4118,N_2912,N_421);
and U4119 (N_4119,N_2093,N_2773);
nor U4120 (N_4120,N_1908,N_1618);
nor U4121 (N_4121,N_2821,N_52);
nor U4122 (N_4122,N_2895,N_2550);
nor U4123 (N_4123,N_887,N_1226);
nand U4124 (N_4124,N_1830,N_2169);
nor U4125 (N_4125,N_2634,N_22);
xor U4126 (N_4126,N_203,N_2915);
and U4127 (N_4127,N_2689,N_337);
and U4128 (N_4128,N_818,N_1691);
nor U4129 (N_4129,N_2487,N_1541);
and U4130 (N_4130,N_1456,N_2805);
xor U4131 (N_4131,N_2482,N_1148);
nand U4132 (N_4132,N_1492,N_1593);
or U4133 (N_4133,N_2410,N_1825);
nor U4134 (N_4134,N_569,N_381);
or U4135 (N_4135,N_2114,N_2190);
nand U4136 (N_4136,N_1406,N_2359);
nor U4137 (N_4137,N_89,N_147);
nor U4138 (N_4138,N_2120,N_1852);
and U4139 (N_4139,N_2836,N_2715);
nand U4140 (N_4140,N_936,N_560);
xnor U4141 (N_4141,N_1849,N_1782);
xor U4142 (N_4142,N_1145,N_1731);
or U4143 (N_4143,N_106,N_2699);
nor U4144 (N_4144,N_1514,N_373);
xnor U4145 (N_4145,N_1009,N_1343);
and U4146 (N_4146,N_1912,N_2532);
nand U4147 (N_4147,N_1277,N_1620);
or U4148 (N_4148,N_2711,N_1614);
nor U4149 (N_4149,N_1468,N_2850);
nor U4150 (N_4150,N_509,N_989);
xor U4151 (N_4151,N_2216,N_720);
xor U4152 (N_4152,N_2312,N_1073);
nand U4153 (N_4153,N_2735,N_857);
nand U4154 (N_4154,N_405,N_1387);
nor U4155 (N_4155,N_503,N_2594);
nor U4156 (N_4156,N_2802,N_1538);
and U4157 (N_4157,N_1674,N_428);
nor U4158 (N_4158,N_2284,N_962);
nor U4159 (N_4159,N_1454,N_1646);
and U4160 (N_4160,N_1440,N_1253);
or U4161 (N_4161,N_2558,N_667);
nand U4162 (N_4162,N_655,N_1083);
nor U4163 (N_4163,N_2496,N_63);
and U4164 (N_4164,N_924,N_1030);
or U4165 (N_4165,N_2412,N_2222);
nand U4166 (N_4166,N_2839,N_899);
nand U4167 (N_4167,N_1463,N_747);
or U4168 (N_4168,N_1361,N_877);
nor U4169 (N_4169,N_525,N_613);
or U4170 (N_4170,N_2414,N_700);
and U4171 (N_4171,N_2436,N_768);
nand U4172 (N_4172,N_2204,N_1035);
nor U4173 (N_4173,N_792,N_2534);
and U4174 (N_4174,N_71,N_1201);
or U4175 (N_4175,N_2708,N_868);
nand U4176 (N_4176,N_2473,N_1734);
nor U4177 (N_4177,N_1710,N_268);
or U4178 (N_4178,N_911,N_2374);
nor U4179 (N_4179,N_1419,N_390);
nand U4180 (N_4180,N_2937,N_1331);
and U4181 (N_4181,N_785,N_1905);
xor U4182 (N_4182,N_459,N_885);
nor U4183 (N_4183,N_2073,N_1584);
xor U4184 (N_4184,N_1302,N_2040);
or U4185 (N_4185,N_313,N_1838);
and U4186 (N_4186,N_2653,N_2832);
nand U4187 (N_4187,N_2086,N_1768);
and U4188 (N_4188,N_345,N_60);
or U4189 (N_4189,N_742,N_2400);
xnor U4190 (N_4190,N_1548,N_531);
and U4191 (N_4191,N_860,N_1118);
and U4192 (N_4192,N_2738,N_2350);
or U4193 (N_4193,N_1811,N_2729);
nor U4194 (N_4194,N_1364,N_210);
xnor U4195 (N_4195,N_2460,N_666);
or U4196 (N_4196,N_1527,N_1833);
or U4197 (N_4197,N_2720,N_289);
and U4198 (N_4198,N_842,N_1611);
nand U4199 (N_4199,N_2492,N_2227);
xnor U4200 (N_4200,N_606,N_752);
and U4201 (N_4201,N_2512,N_1345);
or U4202 (N_4202,N_2687,N_604);
and U4203 (N_4203,N_2535,N_2023);
nor U4204 (N_4204,N_1901,N_766);
and U4205 (N_4205,N_292,N_238);
and U4206 (N_4206,N_12,N_168);
or U4207 (N_4207,N_423,N_2455);
xor U4208 (N_4208,N_1054,N_2952);
nor U4209 (N_4209,N_815,N_357);
nor U4210 (N_4210,N_994,N_1565);
xnor U4211 (N_4211,N_1318,N_2810);
or U4212 (N_4212,N_1929,N_713);
xor U4213 (N_4213,N_775,N_2785);
nor U4214 (N_4214,N_360,N_102);
or U4215 (N_4215,N_2511,N_2369);
or U4216 (N_4216,N_793,N_207);
and U4217 (N_4217,N_1135,N_2302);
nand U4218 (N_4218,N_738,N_2483);
xor U4219 (N_4219,N_2038,N_645);
or U4220 (N_4220,N_1351,N_1439);
xor U4221 (N_4221,N_1165,N_1920);
xor U4222 (N_4222,N_1967,N_120);
and U4223 (N_4223,N_469,N_1704);
nand U4224 (N_4224,N_1832,N_1941);
or U4225 (N_4225,N_425,N_439);
nand U4226 (N_4226,N_2885,N_1894);
xnor U4227 (N_4227,N_1344,N_355);
xor U4228 (N_4228,N_350,N_884);
xnor U4229 (N_4229,N_2418,N_81);
or U4230 (N_4230,N_1686,N_1271);
or U4231 (N_4231,N_1817,N_1130);
or U4232 (N_4232,N_809,N_2507);
or U4233 (N_4233,N_1853,N_1064);
nor U4234 (N_4234,N_593,N_495);
nand U4235 (N_4235,N_494,N_1312);
nand U4236 (N_4236,N_1281,N_1072);
nand U4237 (N_4237,N_513,N_1063);
nand U4238 (N_4238,N_1881,N_968);
nor U4239 (N_4239,N_1227,N_2763);
xnor U4240 (N_4240,N_1763,N_2448);
and U4241 (N_4241,N_1801,N_121);
nand U4242 (N_4242,N_408,N_1166);
and U4243 (N_4243,N_2107,N_2334);
nor U4244 (N_4244,N_2584,N_1505);
nand U4245 (N_4245,N_1753,N_576);
nor U4246 (N_4246,N_504,N_406);
or U4247 (N_4247,N_67,N_53);
nor U4248 (N_4248,N_64,N_1531);
xnor U4249 (N_4249,N_1066,N_2430);
nor U4250 (N_4250,N_1263,N_1997);
nor U4251 (N_4251,N_19,N_769);
nand U4252 (N_4252,N_1680,N_1203);
or U4253 (N_4253,N_2717,N_2887);
xnor U4254 (N_4254,N_2295,N_586);
and U4255 (N_4255,N_539,N_458);
nand U4256 (N_4256,N_1885,N_1976);
and U4257 (N_4257,N_2243,N_554);
nand U4258 (N_4258,N_2060,N_660);
nand U4259 (N_4259,N_2433,N_2612);
xor U4260 (N_4260,N_932,N_1633);
and U4261 (N_4261,N_2983,N_1979);
nand U4262 (N_4262,N_966,N_2575);
and U4263 (N_4263,N_457,N_2130);
nor U4264 (N_4264,N_2310,N_744);
nand U4265 (N_4265,N_1144,N_691);
and U4266 (N_4266,N_2807,N_1927);
nor U4267 (N_4267,N_1657,N_1112);
and U4268 (N_4268,N_1357,N_1371);
or U4269 (N_4269,N_2303,N_440);
nor U4270 (N_4270,N_2526,N_1416);
or U4271 (N_4271,N_477,N_1074);
or U4272 (N_4272,N_2882,N_562);
nor U4273 (N_4273,N_1442,N_1210);
nand U4274 (N_4274,N_1966,N_418);
nand U4275 (N_4275,N_1247,N_384);
nand U4276 (N_4276,N_429,N_1578);
and U4277 (N_4277,N_1969,N_2322);
xor U4278 (N_4278,N_881,N_658);
nor U4279 (N_4279,N_1886,N_225);
or U4280 (N_4280,N_1891,N_895);
xor U4281 (N_4281,N_1598,N_2366);
xnor U4282 (N_4282,N_1026,N_1044);
nor U4283 (N_4283,N_128,N_1648);
nor U4284 (N_4284,N_755,N_2346);
xor U4285 (N_4285,N_2784,N_1882);
nand U4286 (N_4286,N_1139,N_1348);
and U4287 (N_4287,N_137,N_1006);
nand U4288 (N_4288,N_898,N_1507);
nor U4289 (N_4289,N_2238,N_1365);
and U4290 (N_4290,N_1425,N_2208);
xor U4291 (N_4291,N_331,N_588);
xnor U4292 (N_4292,N_862,N_1107);
nor U4293 (N_4293,N_2326,N_1864);
and U4294 (N_4294,N_260,N_2467);
nor U4295 (N_4295,N_2291,N_2442);
or U4296 (N_4296,N_2654,N_2255);
xnor U4297 (N_4297,N_811,N_198);
xnor U4298 (N_4298,N_452,N_1457);
xnor U4299 (N_4299,N_2485,N_2582);
nor U4300 (N_4300,N_2539,N_2276);
nor U4301 (N_4301,N_2300,N_1819);
xor U4302 (N_4302,N_2010,N_1846);
and U4303 (N_4303,N_2928,N_913);
and U4304 (N_4304,N_2924,N_722);
nand U4305 (N_4305,N_800,N_1993);
xor U4306 (N_4306,N_625,N_2913);
xor U4307 (N_4307,N_2646,N_2564);
nor U4308 (N_4308,N_601,N_649);
nor U4309 (N_4309,N_644,N_1011);
nand U4310 (N_4310,N_437,N_2147);
and U4311 (N_4311,N_2065,N_1802);
nor U4312 (N_4312,N_2267,N_2943);
xnor U4313 (N_4313,N_904,N_756);
xnor U4314 (N_4314,N_205,N_734);
nor U4315 (N_4315,N_617,N_409);
or U4316 (N_4316,N_1698,N_558);
and U4317 (N_4317,N_561,N_2435);
nor U4318 (N_4318,N_1879,N_2333);
nand U4319 (N_4319,N_2233,N_2175);
nor U4320 (N_4320,N_1850,N_1888);
nor U4321 (N_4321,N_745,N_2963);
and U4322 (N_4322,N_564,N_2978);
nor U4323 (N_4323,N_2570,N_2920);
nor U4324 (N_4324,N_2670,N_1257);
and U4325 (N_4325,N_151,N_2195);
nor U4326 (N_4326,N_2925,N_2367);
nand U4327 (N_4327,N_2202,N_2661);
nor U4328 (N_4328,N_900,N_1100);
xor U4329 (N_4329,N_1726,N_165);
nand U4330 (N_4330,N_2783,N_827);
or U4331 (N_4331,N_841,N_2352);
nor U4332 (N_4332,N_272,N_2987);
and U4333 (N_4333,N_448,N_1936);
and U4334 (N_4334,N_1616,N_1152);
or U4335 (N_4335,N_551,N_506);
and U4336 (N_4336,N_1182,N_2867);
xor U4337 (N_4337,N_2089,N_1877);
nor U4338 (N_4338,N_2907,N_1412);
nand U4339 (N_4339,N_2965,N_2283);
nor U4340 (N_4340,N_1720,N_2959);
and U4341 (N_4341,N_2608,N_516);
nand U4342 (N_4342,N_2464,N_2426);
nor U4343 (N_4343,N_2099,N_1824);
nand U4344 (N_4344,N_2855,N_594);
and U4345 (N_4345,N_799,N_563);
or U4346 (N_4346,N_2529,N_1322);
nor U4347 (N_4347,N_1326,N_1058);
xor U4348 (N_4348,N_2508,N_699);
and U4349 (N_4349,N_1737,N_1968);
nand U4350 (N_4350,N_2083,N_2873);
or U4351 (N_4351,N_2287,N_2676);
or U4352 (N_4352,N_453,N_2862);
or U4353 (N_4353,N_1581,N_2314);
xnor U4354 (N_4354,N_1108,N_2434);
or U4355 (N_4355,N_829,N_2343);
nand U4356 (N_4356,N_2170,N_1878);
nand U4357 (N_4357,N_2372,N_781);
nand U4358 (N_4358,N_2142,N_883);
nand U4359 (N_4359,N_2790,N_2012);
xor U4360 (N_4360,N_1383,N_565);
or U4361 (N_4361,N_1585,N_2212);
nor U4362 (N_4362,N_2934,N_1151);
and U4363 (N_4363,N_116,N_2704);
or U4364 (N_4364,N_2591,N_1827);
or U4365 (N_4365,N_1847,N_727);
xor U4366 (N_4366,N_1922,N_33);
nor U4367 (N_4367,N_2655,N_435);
nand U4368 (N_4368,N_546,N_518);
or U4369 (N_4369,N_1600,N_1156);
xnor U4370 (N_4370,N_2520,N_284);
nand U4371 (N_4371,N_753,N_2642);
or U4372 (N_4372,N_2722,N_31);
and U4373 (N_4373,N_1487,N_2846);
nand U4374 (N_4374,N_1290,N_1785);
nor U4375 (N_4375,N_2404,N_2017);
nand U4376 (N_4376,N_2849,N_280);
nand U4377 (N_4377,N_2749,N_161);
xnor U4378 (N_4378,N_1571,N_821);
or U4379 (N_4379,N_49,N_2054);
nand U4380 (N_4380,N_599,N_1032);
and U4381 (N_4381,N_1012,N_1615);
xnor U4382 (N_4382,N_132,N_2210);
nand U4383 (N_4383,N_291,N_2398);
and U4384 (N_4384,N_1289,N_417);
nand U4385 (N_4385,N_1109,N_2476);
or U4386 (N_4386,N_945,N_2500);
nor U4387 (N_4387,N_2249,N_493);
nor U4388 (N_4388,N_1587,N_248);
or U4389 (N_4389,N_2859,N_2080);
nor U4390 (N_4390,N_1462,N_95);
xor U4391 (N_4391,N_2871,N_2692);
nand U4392 (N_4392,N_182,N_228);
nand U4393 (N_4393,N_2515,N_1535);
or U4394 (N_4394,N_2456,N_2600);
or U4395 (N_4395,N_2324,N_2331);
nand U4396 (N_4396,N_725,N_1856);
nand U4397 (N_4397,N_2479,N_2886);
nand U4398 (N_4398,N_1385,N_1283);
xor U4399 (N_4399,N_804,N_1433);
nand U4400 (N_4400,N_993,N_1897);
xor U4401 (N_4401,N_1260,N_2458);
or U4402 (N_4402,N_464,N_2186);
xnor U4403 (N_4403,N_1909,N_46);
xnor U4404 (N_4404,N_1750,N_2936);
and U4405 (N_4405,N_1742,N_2890);
and U4406 (N_4406,N_130,N_774);
xor U4407 (N_4407,N_750,N_2931);
nor U4408 (N_4408,N_2207,N_888);
xnor U4409 (N_4409,N_1141,N_1299);
nor U4410 (N_4410,N_240,N_1474);
and U4411 (N_4411,N_1147,N_1256);
or U4412 (N_4412,N_1489,N_2542);
or U4413 (N_4413,N_487,N_2569);
or U4414 (N_4414,N_880,N_2056);
nand U4415 (N_4415,N_2213,N_2674);
and U4416 (N_4416,N_2554,N_1911);
nor U4417 (N_4417,N_397,N_786);
or U4418 (N_4418,N_1981,N_2533);
or U4419 (N_4419,N_322,N_348);
and U4420 (N_4420,N_1191,N_1957);
and U4421 (N_4421,N_2980,N_1239);
or U4422 (N_4422,N_704,N_84);
and U4423 (N_4423,N_1354,N_204);
xnor U4424 (N_4424,N_97,N_555);
or U4425 (N_4425,N_2854,N_553);
nor U4426 (N_4426,N_1195,N_2323);
nor U4427 (N_4427,N_1048,N_701);
nor U4428 (N_4428,N_2538,N_2870);
or U4429 (N_4429,N_191,N_2478);
nor U4430 (N_4430,N_100,N_984);
nor U4431 (N_4431,N_1308,N_124);
and U4432 (N_4432,N_1576,N_2577);
nand U4433 (N_4433,N_2391,N_1400);
xnor U4434 (N_4434,N_1583,N_278);
or U4435 (N_4435,N_1666,N_2942);
and U4436 (N_4436,N_2257,N_871);
nor U4437 (N_4437,N_2657,N_571);
nor U4438 (N_4438,N_1004,N_178);
or U4439 (N_4439,N_229,N_708);
xor U4440 (N_4440,N_2224,N_1550);
nand U4441 (N_4441,N_2603,N_692);
nor U4442 (N_4442,N_1495,N_2156);
and U4443 (N_4443,N_2046,N_2828);
or U4444 (N_4444,N_2892,N_2493);
or U4445 (N_4445,N_1623,N_1180);
nand U4446 (N_4446,N_2246,N_396);
xor U4447 (N_4447,N_524,N_517);
or U4448 (N_4448,N_1373,N_1655);
nand U4449 (N_4449,N_1563,N_153);
and U4450 (N_4450,N_1980,N_2510);
and U4451 (N_4451,N_2700,N_86);
nand U4452 (N_4452,N_894,N_2354);
nor U4453 (N_4453,N_2218,N_1025);
nor U4454 (N_4454,N_2231,N_329);
or U4455 (N_4455,N_2144,N_935);
nor U4456 (N_4456,N_2905,N_959);
or U4457 (N_4457,N_1752,N_1088);
nor U4458 (N_4458,N_2723,N_2275);
nor U4459 (N_4459,N_2250,N_929);
xor U4460 (N_4460,N_858,N_172);
and U4461 (N_4461,N_1510,N_2049);
and U4462 (N_4462,N_1105,N_597);
and U4463 (N_4463,N_1062,N_497);
and U4464 (N_4464,N_2094,N_1175);
xnor U4465 (N_4465,N_1255,N_2631);
nand U4466 (N_4466,N_32,N_873);
and U4467 (N_4467,N_909,N_893);
nand U4468 (N_4468,N_2840,N_1214);
or U4469 (N_4469,N_393,N_2829);
xnor U4470 (N_4470,N_2648,N_1154);
xnor U4471 (N_4471,N_29,N_2922);
nor U4472 (N_4472,N_236,N_656);
xnor U4473 (N_4473,N_376,N_927);
or U4474 (N_4474,N_2901,N_2293);
nand U4475 (N_4475,N_1504,N_840);
xor U4476 (N_4476,N_2288,N_582);
or U4477 (N_4477,N_2466,N_1990);
nor U4478 (N_4478,N_907,N_1546);
or U4479 (N_4479,N_307,N_856);
and U4480 (N_4480,N_2032,N_2245);
nor U4481 (N_4481,N_632,N_2076);
and U4482 (N_4482,N_1448,N_1679);
nand U4483 (N_4483,N_965,N_2734);
and U4484 (N_4484,N_1573,N_639);
xnor U4485 (N_4485,N_2736,N_1836);
nor U4486 (N_4486,N_812,N_1635);
xnor U4487 (N_4487,N_1697,N_2758);
and U4488 (N_4488,N_1572,N_1319);
nor U4489 (N_4489,N_54,N_890);
xor U4490 (N_4490,N_1835,N_1866);
or U4491 (N_4491,N_170,N_529);
nand U4492 (N_4492,N_2530,N_2183);
xor U4493 (N_4493,N_2814,N_865);
nor U4494 (N_4494,N_2265,N_358);
or U4495 (N_4495,N_176,N_1363);
nand U4496 (N_4496,N_2844,N_270);
xnor U4497 (N_4497,N_309,N_1230);
xnor U4498 (N_4498,N_740,N_199);
nand U4499 (N_4499,N_2751,N_61);
xnor U4500 (N_4500,N_23,N_1685);
or U4501 (N_4501,N_2562,N_1359);
or U4502 (N_4502,N_1252,N_2832);
nand U4503 (N_4503,N_294,N_1552);
nor U4504 (N_4504,N_2725,N_633);
or U4505 (N_4505,N_1898,N_684);
or U4506 (N_4506,N_2268,N_2346);
nand U4507 (N_4507,N_1597,N_2915);
or U4508 (N_4508,N_289,N_1339);
xor U4509 (N_4509,N_150,N_815);
xnor U4510 (N_4510,N_241,N_2395);
nand U4511 (N_4511,N_8,N_1129);
nor U4512 (N_4512,N_315,N_1438);
xor U4513 (N_4513,N_451,N_1910);
and U4514 (N_4514,N_2734,N_2248);
nor U4515 (N_4515,N_2299,N_930);
nor U4516 (N_4516,N_2487,N_2257);
or U4517 (N_4517,N_2686,N_1624);
nand U4518 (N_4518,N_1438,N_2023);
nor U4519 (N_4519,N_2754,N_1650);
or U4520 (N_4520,N_796,N_1532);
nor U4521 (N_4521,N_2845,N_196);
xnor U4522 (N_4522,N_1924,N_393);
or U4523 (N_4523,N_2614,N_1347);
xor U4524 (N_4524,N_2061,N_1360);
nand U4525 (N_4525,N_2824,N_1457);
xnor U4526 (N_4526,N_2888,N_1190);
nor U4527 (N_4527,N_1704,N_2922);
nand U4528 (N_4528,N_2128,N_2813);
nand U4529 (N_4529,N_833,N_494);
nor U4530 (N_4530,N_221,N_628);
nor U4531 (N_4531,N_1009,N_284);
xnor U4532 (N_4532,N_2821,N_84);
or U4533 (N_4533,N_1722,N_1646);
nor U4534 (N_4534,N_2521,N_2409);
xnor U4535 (N_4535,N_280,N_207);
xnor U4536 (N_4536,N_100,N_1361);
xnor U4537 (N_4537,N_1653,N_2015);
nand U4538 (N_4538,N_2613,N_1721);
nor U4539 (N_4539,N_2475,N_2535);
xnor U4540 (N_4540,N_329,N_341);
and U4541 (N_4541,N_331,N_421);
xnor U4542 (N_4542,N_2941,N_2107);
nand U4543 (N_4543,N_46,N_1205);
nand U4544 (N_4544,N_1087,N_1732);
and U4545 (N_4545,N_2767,N_1042);
nor U4546 (N_4546,N_1465,N_149);
nor U4547 (N_4547,N_1852,N_661);
and U4548 (N_4548,N_2047,N_257);
nor U4549 (N_4549,N_2188,N_1673);
and U4550 (N_4550,N_2660,N_1284);
nor U4551 (N_4551,N_1468,N_2309);
nor U4552 (N_4552,N_1202,N_326);
nor U4553 (N_4553,N_1159,N_2533);
nand U4554 (N_4554,N_2503,N_568);
xor U4555 (N_4555,N_849,N_2999);
and U4556 (N_4556,N_2046,N_417);
and U4557 (N_4557,N_2343,N_1705);
nand U4558 (N_4558,N_390,N_601);
or U4559 (N_4559,N_1548,N_2486);
or U4560 (N_4560,N_1592,N_2362);
or U4561 (N_4561,N_1049,N_2037);
and U4562 (N_4562,N_1802,N_402);
xnor U4563 (N_4563,N_2072,N_1094);
and U4564 (N_4564,N_795,N_718);
and U4565 (N_4565,N_1950,N_2433);
xnor U4566 (N_4566,N_2576,N_2917);
nor U4567 (N_4567,N_2770,N_2678);
and U4568 (N_4568,N_2170,N_2982);
xnor U4569 (N_4569,N_1905,N_636);
nand U4570 (N_4570,N_2994,N_722);
xor U4571 (N_4571,N_1413,N_1172);
and U4572 (N_4572,N_2982,N_2524);
nor U4573 (N_4573,N_328,N_2265);
nor U4574 (N_4574,N_357,N_1772);
and U4575 (N_4575,N_699,N_1183);
nand U4576 (N_4576,N_1759,N_498);
or U4577 (N_4577,N_579,N_620);
nand U4578 (N_4578,N_183,N_1224);
or U4579 (N_4579,N_1400,N_1640);
nor U4580 (N_4580,N_674,N_816);
nor U4581 (N_4581,N_2307,N_415);
and U4582 (N_4582,N_1577,N_296);
or U4583 (N_4583,N_488,N_2155);
or U4584 (N_4584,N_1025,N_271);
xor U4585 (N_4585,N_1423,N_257);
nor U4586 (N_4586,N_44,N_2499);
and U4587 (N_4587,N_2776,N_22);
nor U4588 (N_4588,N_1945,N_1913);
nor U4589 (N_4589,N_1180,N_1937);
or U4590 (N_4590,N_1882,N_1250);
or U4591 (N_4591,N_1423,N_877);
and U4592 (N_4592,N_2637,N_2742);
xor U4593 (N_4593,N_1846,N_1443);
nor U4594 (N_4594,N_943,N_1719);
and U4595 (N_4595,N_2460,N_2500);
or U4596 (N_4596,N_599,N_1112);
nor U4597 (N_4597,N_2432,N_1953);
nand U4598 (N_4598,N_2391,N_1479);
xnor U4599 (N_4599,N_2334,N_2354);
nor U4600 (N_4600,N_2528,N_1313);
and U4601 (N_4601,N_2318,N_2237);
xor U4602 (N_4602,N_491,N_2627);
or U4603 (N_4603,N_1500,N_991);
xor U4604 (N_4604,N_1792,N_32);
nor U4605 (N_4605,N_1167,N_2967);
xor U4606 (N_4606,N_1040,N_784);
or U4607 (N_4607,N_2546,N_811);
and U4608 (N_4608,N_165,N_489);
xnor U4609 (N_4609,N_2472,N_1482);
nor U4610 (N_4610,N_2412,N_2849);
xor U4611 (N_4611,N_2210,N_740);
or U4612 (N_4612,N_778,N_1796);
nor U4613 (N_4613,N_1847,N_2662);
nand U4614 (N_4614,N_795,N_2750);
nor U4615 (N_4615,N_1615,N_2841);
or U4616 (N_4616,N_2467,N_2607);
and U4617 (N_4617,N_2740,N_1954);
nand U4618 (N_4618,N_1124,N_818);
xor U4619 (N_4619,N_1146,N_1079);
or U4620 (N_4620,N_2574,N_140);
nand U4621 (N_4621,N_1482,N_1420);
nor U4622 (N_4622,N_1892,N_617);
and U4623 (N_4623,N_2806,N_1507);
nand U4624 (N_4624,N_522,N_553);
nor U4625 (N_4625,N_77,N_267);
xnor U4626 (N_4626,N_1329,N_442);
nor U4627 (N_4627,N_1083,N_1940);
nand U4628 (N_4628,N_2660,N_2896);
xor U4629 (N_4629,N_2275,N_469);
nand U4630 (N_4630,N_1904,N_679);
or U4631 (N_4631,N_2220,N_2779);
nand U4632 (N_4632,N_2823,N_56);
nor U4633 (N_4633,N_828,N_539);
nand U4634 (N_4634,N_1418,N_2261);
nand U4635 (N_4635,N_2987,N_561);
xnor U4636 (N_4636,N_240,N_344);
and U4637 (N_4637,N_106,N_2712);
nor U4638 (N_4638,N_2688,N_1852);
and U4639 (N_4639,N_2722,N_850);
and U4640 (N_4640,N_1711,N_269);
nand U4641 (N_4641,N_2433,N_572);
and U4642 (N_4642,N_1859,N_684);
nand U4643 (N_4643,N_1361,N_1314);
xor U4644 (N_4644,N_2516,N_742);
or U4645 (N_4645,N_1655,N_296);
nand U4646 (N_4646,N_973,N_1434);
or U4647 (N_4647,N_2245,N_128);
xor U4648 (N_4648,N_223,N_2219);
nor U4649 (N_4649,N_1049,N_1481);
nor U4650 (N_4650,N_2656,N_2182);
nor U4651 (N_4651,N_378,N_1091);
or U4652 (N_4652,N_2038,N_446);
and U4653 (N_4653,N_1114,N_2692);
nor U4654 (N_4654,N_74,N_568);
nor U4655 (N_4655,N_1116,N_781);
xor U4656 (N_4656,N_1167,N_1192);
nand U4657 (N_4657,N_2450,N_1779);
or U4658 (N_4658,N_2797,N_1570);
or U4659 (N_4659,N_645,N_1816);
and U4660 (N_4660,N_1261,N_1915);
nand U4661 (N_4661,N_2705,N_1293);
and U4662 (N_4662,N_488,N_897);
or U4663 (N_4663,N_1158,N_2721);
nand U4664 (N_4664,N_1765,N_206);
nand U4665 (N_4665,N_916,N_1396);
nand U4666 (N_4666,N_230,N_1485);
and U4667 (N_4667,N_719,N_1631);
nor U4668 (N_4668,N_2057,N_1630);
nor U4669 (N_4669,N_1948,N_338);
and U4670 (N_4670,N_2448,N_551);
nand U4671 (N_4671,N_73,N_1665);
nand U4672 (N_4672,N_1603,N_718);
and U4673 (N_4673,N_541,N_859);
xnor U4674 (N_4674,N_1175,N_66);
nor U4675 (N_4675,N_690,N_2363);
xor U4676 (N_4676,N_2908,N_1033);
xnor U4677 (N_4677,N_625,N_2606);
or U4678 (N_4678,N_1510,N_2261);
nor U4679 (N_4679,N_68,N_295);
xnor U4680 (N_4680,N_436,N_585);
nand U4681 (N_4681,N_2746,N_2514);
nor U4682 (N_4682,N_1347,N_18);
or U4683 (N_4683,N_166,N_879);
or U4684 (N_4684,N_1128,N_772);
or U4685 (N_4685,N_1095,N_352);
xnor U4686 (N_4686,N_2926,N_2001);
and U4687 (N_4687,N_1614,N_2665);
or U4688 (N_4688,N_1129,N_1555);
nor U4689 (N_4689,N_1874,N_1032);
nor U4690 (N_4690,N_1060,N_1685);
nand U4691 (N_4691,N_1430,N_1077);
and U4692 (N_4692,N_958,N_1601);
nor U4693 (N_4693,N_605,N_1693);
nand U4694 (N_4694,N_429,N_888);
nor U4695 (N_4695,N_1589,N_1108);
xor U4696 (N_4696,N_2486,N_1195);
nor U4697 (N_4697,N_819,N_1680);
or U4698 (N_4698,N_2423,N_274);
xor U4699 (N_4699,N_1908,N_192);
and U4700 (N_4700,N_758,N_1063);
nor U4701 (N_4701,N_2019,N_2075);
nand U4702 (N_4702,N_1602,N_1659);
and U4703 (N_4703,N_1933,N_735);
or U4704 (N_4704,N_697,N_575);
and U4705 (N_4705,N_859,N_877);
and U4706 (N_4706,N_1139,N_1519);
xnor U4707 (N_4707,N_1377,N_322);
and U4708 (N_4708,N_826,N_1919);
and U4709 (N_4709,N_2947,N_2249);
and U4710 (N_4710,N_1999,N_991);
or U4711 (N_4711,N_902,N_1390);
nand U4712 (N_4712,N_1488,N_1844);
or U4713 (N_4713,N_2065,N_2288);
nor U4714 (N_4714,N_2365,N_927);
xor U4715 (N_4715,N_419,N_24);
or U4716 (N_4716,N_878,N_1022);
and U4717 (N_4717,N_1469,N_740);
nand U4718 (N_4718,N_1440,N_2102);
and U4719 (N_4719,N_2894,N_1072);
nand U4720 (N_4720,N_1278,N_872);
xor U4721 (N_4721,N_1378,N_2809);
nor U4722 (N_4722,N_684,N_1428);
xor U4723 (N_4723,N_18,N_2605);
nand U4724 (N_4724,N_651,N_548);
and U4725 (N_4725,N_1201,N_1157);
nor U4726 (N_4726,N_798,N_2054);
and U4727 (N_4727,N_1049,N_1785);
nor U4728 (N_4728,N_2608,N_1015);
and U4729 (N_4729,N_2083,N_2501);
and U4730 (N_4730,N_938,N_1400);
or U4731 (N_4731,N_1813,N_2951);
or U4732 (N_4732,N_2494,N_1319);
nor U4733 (N_4733,N_1964,N_550);
nand U4734 (N_4734,N_1217,N_1920);
or U4735 (N_4735,N_2169,N_455);
nor U4736 (N_4736,N_1913,N_2858);
nand U4737 (N_4737,N_167,N_1875);
and U4738 (N_4738,N_387,N_2817);
xnor U4739 (N_4739,N_2413,N_578);
nor U4740 (N_4740,N_2626,N_1189);
nor U4741 (N_4741,N_2382,N_310);
xor U4742 (N_4742,N_2181,N_2911);
and U4743 (N_4743,N_237,N_1619);
or U4744 (N_4744,N_1273,N_1978);
nand U4745 (N_4745,N_2809,N_637);
nor U4746 (N_4746,N_852,N_417);
or U4747 (N_4747,N_1003,N_129);
nand U4748 (N_4748,N_161,N_1734);
xor U4749 (N_4749,N_1219,N_2623);
or U4750 (N_4750,N_1201,N_818);
xnor U4751 (N_4751,N_2422,N_2634);
nand U4752 (N_4752,N_185,N_2726);
xor U4753 (N_4753,N_1773,N_1584);
and U4754 (N_4754,N_2104,N_1612);
or U4755 (N_4755,N_1041,N_1215);
nor U4756 (N_4756,N_1444,N_1333);
and U4757 (N_4757,N_2026,N_955);
xor U4758 (N_4758,N_2135,N_1548);
xnor U4759 (N_4759,N_1366,N_880);
nor U4760 (N_4760,N_1167,N_1569);
nor U4761 (N_4761,N_1086,N_1502);
xor U4762 (N_4762,N_1432,N_1655);
nand U4763 (N_4763,N_505,N_836);
xor U4764 (N_4764,N_874,N_2174);
xnor U4765 (N_4765,N_2149,N_2615);
nand U4766 (N_4766,N_9,N_2658);
nand U4767 (N_4767,N_2948,N_239);
nor U4768 (N_4768,N_2719,N_1274);
nand U4769 (N_4769,N_1611,N_1956);
xor U4770 (N_4770,N_1178,N_2261);
nor U4771 (N_4771,N_2902,N_1179);
and U4772 (N_4772,N_13,N_2001);
nor U4773 (N_4773,N_769,N_2971);
and U4774 (N_4774,N_2956,N_2580);
xor U4775 (N_4775,N_386,N_1954);
and U4776 (N_4776,N_1639,N_2682);
xor U4777 (N_4777,N_1185,N_1668);
nor U4778 (N_4778,N_2576,N_1285);
nor U4779 (N_4779,N_1481,N_945);
and U4780 (N_4780,N_1937,N_2579);
and U4781 (N_4781,N_1225,N_137);
or U4782 (N_4782,N_641,N_1888);
xnor U4783 (N_4783,N_288,N_2375);
nand U4784 (N_4784,N_742,N_2360);
nor U4785 (N_4785,N_641,N_699);
nor U4786 (N_4786,N_2034,N_54);
nor U4787 (N_4787,N_961,N_1783);
xor U4788 (N_4788,N_2832,N_2831);
nor U4789 (N_4789,N_1669,N_2540);
and U4790 (N_4790,N_1119,N_195);
nor U4791 (N_4791,N_2975,N_1544);
nand U4792 (N_4792,N_626,N_1547);
and U4793 (N_4793,N_1723,N_1464);
and U4794 (N_4794,N_337,N_927);
and U4795 (N_4795,N_1419,N_1207);
nor U4796 (N_4796,N_2657,N_1948);
xor U4797 (N_4797,N_1165,N_2021);
nor U4798 (N_4798,N_2990,N_340);
nor U4799 (N_4799,N_1480,N_1740);
nand U4800 (N_4800,N_1159,N_2130);
or U4801 (N_4801,N_1779,N_514);
nor U4802 (N_4802,N_90,N_560);
nand U4803 (N_4803,N_846,N_1784);
or U4804 (N_4804,N_1133,N_2316);
and U4805 (N_4805,N_2556,N_2116);
nor U4806 (N_4806,N_1624,N_2159);
or U4807 (N_4807,N_530,N_2553);
or U4808 (N_4808,N_1609,N_1147);
xor U4809 (N_4809,N_1996,N_432);
nor U4810 (N_4810,N_1453,N_2714);
xor U4811 (N_4811,N_2619,N_2939);
nand U4812 (N_4812,N_2176,N_904);
or U4813 (N_4813,N_2042,N_1751);
xor U4814 (N_4814,N_1656,N_2333);
or U4815 (N_4815,N_449,N_1247);
and U4816 (N_4816,N_1511,N_2816);
or U4817 (N_4817,N_793,N_656);
and U4818 (N_4818,N_2834,N_2467);
xnor U4819 (N_4819,N_1285,N_605);
and U4820 (N_4820,N_2243,N_1044);
xnor U4821 (N_4821,N_197,N_436);
or U4822 (N_4822,N_7,N_1168);
or U4823 (N_4823,N_2079,N_746);
nor U4824 (N_4824,N_2077,N_818);
and U4825 (N_4825,N_566,N_1189);
nand U4826 (N_4826,N_327,N_2997);
nor U4827 (N_4827,N_2974,N_852);
xnor U4828 (N_4828,N_2948,N_91);
xnor U4829 (N_4829,N_2694,N_2152);
nand U4830 (N_4830,N_2842,N_2151);
and U4831 (N_4831,N_1131,N_1310);
or U4832 (N_4832,N_2952,N_2127);
xor U4833 (N_4833,N_2767,N_435);
and U4834 (N_4834,N_1113,N_2437);
xnor U4835 (N_4835,N_1065,N_2463);
and U4836 (N_4836,N_1124,N_95);
nand U4837 (N_4837,N_874,N_1743);
xnor U4838 (N_4838,N_2791,N_833);
nor U4839 (N_4839,N_1475,N_1347);
nor U4840 (N_4840,N_2123,N_2749);
and U4841 (N_4841,N_1691,N_2728);
and U4842 (N_4842,N_252,N_607);
nor U4843 (N_4843,N_1698,N_1780);
and U4844 (N_4844,N_1553,N_1361);
and U4845 (N_4845,N_49,N_2167);
nor U4846 (N_4846,N_1824,N_2202);
nor U4847 (N_4847,N_897,N_1529);
or U4848 (N_4848,N_206,N_1131);
nand U4849 (N_4849,N_995,N_1540);
or U4850 (N_4850,N_1772,N_1430);
nor U4851 (N_4851,N_242,N_1550);
and U4852 (N_4852,N_1967,N_2371);
and U4853 (N_4853,N_151,N_672);
nor U4854 (N_4854,N_1548,N_17);
and U4855 (N_4855,N_2142,N_2774);
nor U4856 (N_4856,N_857,N_2843);
nand U4857 (N_4857,N_1737,N_2784);
and U4858 (N_4858,N_1923,N_1389);
or U4859 (N_4859,N_841,N_217);
nor U4860 (N_4860,N_2924,N_2542);
and U4861 (N_4861,N_306,N_2046);
nor U4862 (N_4862,N_1608,N_2197);
xor U4863 (N_4863,N_1859,N_2569);
xnor U4864 (N_4864,N_2915,N_1683);
xor U4865 (N_4865,N_385,N_2969);
nand U4866 (N_4866,N_776,N_1675);
or U4867 (N_4867,N_1262,N_138);
nor U4868 (N_4868,N_1310,N_1252);
or U4869 (N_4869,N_519,N_2449);
and U4870 (N_4870,N_2563,N_1557);
and U4871 (N_4871,N_1536,N_2305);
xor U4872 (N_4872,N_1239,N_279);
or U4873 (N_4873,N_2799,N_824);
nand U4874 (N_4874,N_65,N_706);
or U4875 (N_4875,N_757,N_1300);
xnor U4876 (N_4876,N_625,N_1150);
and U4877 (N_4877,N_278,N_2172);
nand U4878 (N_4878,N_1812,N_992);
nand U4879 (N_4879,N_1829,N_1994);
nor U4880 (N_4880,N_2264,N_482);
nand U4881 (N_4881,N_1261,N_463);
and U4882 (N_4882,N_938,N_405);
and U4883 (N_4883,N_1387,N_2925);
nor U4884 (N_4884,N_1255,N_1037);
nand U4885 (N_4885,N_256,N_1785);
xnor U4886 (N_4886,N_918,N_2790);
nand U4887 (N_4887,N_655,N_2497);
nand U4888 (N_4888,N_507,N_2555);
and U4889 (N_4889,N_985,N_2237);
and U4890 (N_4890,N_922,N_2599);
nor U4891 (N_4891,N_2174,N_971);
nand U4892 (N_4892,N_1081,N_1723);
xnor U4893 (N_4893,N_262,N_1819);
xnor U4894 (N_4894,N_444,N_816);
nor U4895 (N_4895,N_1590,N_2741);
and U4896 (N_4896,N_568,N_2666);
and U4897 (N_4897,N_1751,N_972);
nor U4898 (N_4898,N_803,N_2375);
and U4899 (N_4899,N_2696,N_418);
or U4900 (N_4900,N_973,N_927);
nor U4901 (N_4901,N_1868,N_359);
nand U4902 (N_4902,N_1241,N_1469);
or U4903 (N_4903,N_1843,N_141);
and U4904 (N_4904,N_2196,N_2617);
nor U4905 (N_4905,N_267,N_2138);
nor U4906 (N_4906,N_150,N_2138);
or U4907 (N_4907,N_2797,N_1719);
and U4908 (N_4908,N_88,N_822);
and U4909 (N_4909,N_208,N_2304);
or U4910 (N_4910,N_1610,N_1480);
and U4911 (N_4911,N_1028,N_1423);
nor U4912 (N_4912,N_1986,N_875);
nor U4913 (N_4913,N_151,N_1878);
or U4914 (N_4914,N_2469,N_1391);
xnor U4915 (N_4915,N_837,N_1815);
or U4916 (N_4916,N_1563,N_1773);
and U4917 (N_4917,N_1293,N_699);
xor U4918 (N_4918,N_2260,N_2607);
nand U4919 (N_4919,N_469,N_1763);
nand U4920 (N_4920,N_598,N_41);
nand U4921 (N_4921,N_1071,N_1801);
nor U4922 (N_4922,N_2578,N_2511);
nand U4923 (N_4923,N_1297,N_1498);
and U4924 (N_4924,N_278,N_181);
or U4925 (N_4925,N_1324,N_2128);
nand U4926 (N_4926,N_2650,N_287);
and U4927 (N_4927,N_1368,N_68);
or U4928 (N_4928,N_2997,N_1189);
xor U4929 (N_4929,N_218,N_2248);
or U4930 (N_4930,N_2188,N_319);
and U4931 (N_4931,N_2643,N_2711);
and U4932 (N_4932,N_1036,N_966);
nand U4933 (N_4933,N_576,N_821);
xnor U4934 (N_4934,N_2455,N_916);
and U4935 (N_4935,N_2327,N_287);
or U4936 (N_4936,N_2350,N_556);
and U4937 (N_4937,N_773,N_37);
xor U4938 (N_4938,N_2375,N_1543);
nor U4939 (N_4939,N_378,N_1864);
or U4940 (N_4940,N_2846,N_1536);
nor U4941 (N_4941,N_1722,N_984);
or U4942 (N_4942,N_1150,N_1730);
or U4943 (N_4943,N_590,N_298);
xnor U4944 (N_4944,N_1877,N_2168);
nor U4945 (N_4945,N_2690,N_2218);
xor U4946 (N_4946,N_541,N_623);
or U4947 (N_4947,N_2150,N_2970);
nor U4948 (N_4948,N_677,N_124);
nand U4949 (N_4949,N_657,N_395);
or U4950 (N_4950,N_2058,N_1620);
xnor U4951 (N_4951,N_2682,N_2393);
and U4952 (N_4952,N_2030,N_2484);
nand U4953 (N_4953,N_1977,N_1309);
or U4954 (N_4954,N_1906,N_2524);
nand U4955 (N_4955,N_473,N_1538);
xor U4956 (N_4956,N_2724,N_1171);
nand U4957 (N_4957,N_1502,N_2925);
xnor U4958 (N_4958,N_438,N_1631);
nand U4959 (N_4959,N_604,N_1081);
xnor U4960 (N_4960,N_2498,N_397);
or U4961 (N_4961,N_1409,N_1483);
and U4962 (N_4962,N_999,N_2993);
or U4963 (N_4963,N_1464,N_786);
xnor U4964 (N_4964,N_1333,N_2655);
and U4965 (N_4965,N_2594,N_2208);
and U4966 (N_4966,N_895,N_715);
nand U4967 (N_4967,N_372,N_877);
xor U4968 (N_4968,N_2548,N_464);
xor U4969 (N_4969,N_4,N_2998);
and U4970 (N_4970,N_480,N_1903);
or U4971 (N_4971,N_475,N_1816);
and U4972 (N_4972,N_1393,N_2367);
xnor U4973 (N_4973,N_1889,N_309);
nor U4974 (N_4974,N_1310,N_1795);
nand U4975 (N_4975,N_30,N_597);
nor U4976 (N_4976,N_2150,N_99);
and U4977 (N_4977,N_26,N_2525);
nand U4978 (N_4978,N_1454,N_334);
nand U4979 (N_4979,N_2982,N_2741);
nand U4980 (N_4980,N_1556,N_729);
and U4981 (N_4981,N_1868,N_2702);
and U4982 (N_4982,N_1598,N_248);
and U4983 (N_4983,N_928,N_2308);
or U4984 (N_4984,N_1183,N_1234);
nand U4985 (N_4985,N_1563,N_2706);
nand U4986 (N_4986,N_1521,N_1695);
or U4987 (N_4987,N_1822,N_218);
and U4988 (N_4988,N_1248,N_29);
nor U4989 (N_4989,N_1420,N_1119);
or U4990 (N_4990,N_1899,N_1340);
nand U4991 (N_4991,N_866,N_2466);
xnor U4992 (N_4992,N_1796,N_2742);
or U4993 (N_4993,N_236,N_2263);
nor U4994 (N_4994,N_39,N_794);
nand U4995 (N_4995,N_241,N_2773);
xnor U4996 (N_4996,N_1883,N_1713);
or U4997 (N_4997,N_323,N_983);
nand U4998 (N_4998,N_2464,N_149);
or U4999 (N_4999,N_1439,N_2258);
nor U5000 (N_5000,N_2694,N_1160);
nand U5001 (N_5001,N_319,N_2361);
nor U5002 (N_5002,N_474,N_433);
and U5003 (N_5003,N_1612,N_2795);
nand U5004 (N_5004,N_1735,N_436);
xor U5005 (N_5005,N_820,N_2859);
and U5006 (N_5006,N_243,N_2173);
or U5007 (N_5007,N_472,N_2380);
and U5008 (N_5008,N_34,N_418);
or U5009 (N_5009,N_2153,N_2470);
nand U5010 (N_5010,N_1820,N_2334);
nor U5011 (N_5011,N_347,N_1085);
nor U5012 (N_5012,N_557,N_1013);
nor U5013 (N_5013,N_2478,N_1377);
xor U5014 (N_5014,N_1769,N_961);
and U5015 (N_5015,N_2061,N_1282);
nor U5016 (N_5016,N_42,N_1366);
xor U5017 (N_5017,N_2943,N_2946);
or U5018 (N_5018,N_967,N_2454);
nand U5019 (N_5019,N_1808,N_1768);
or U5020 (N_5020,N_2903,N_1895);
nand U5021 (N_5021,N_928,N_1226);
nand U5022 (N_5022,N_700,N_1135);
nor U5023 (N_5023,N_2635,N_1575);
nor U5024 (N_5024,N_754,N_1475);
xor U5025 (N_5025,N_1637,N_112);
nand U5026 (N_5026,N_268,N_723);
nor U5027 (N_5027,N_2230,N_2197);
nor U5028 (N_5028,N_2064,N_629);
nand U5029 (N_5029,N_739,N_1185);
or U5030 (N_5030,N_64,N_2129);
and U5031 (N_5031,N_1017,N_721);
or U5032 (N_5032,N_1692,N_500);
xor U5033 (N_5033,N_2376,N_1897);
nand U5034 (N_5034,N_2520,N_2438);
and U5035 (N_5035,N_2317,N_1330);
and U5036 (N_5036,N_2795,N_1165);
nand U5037 (N_5037,N_1834,N_1081);
nor U5038 (N_5038,N_2087,N_597);
and U5039 (N_5039,N_161,N_2352);
or U5040 (N_5040,N_71,N_1022);
nor U5041 (N_5041,N_2471,N_2917);
or U5042 (N_5042,N_2233,N_1309);
nand U5043 (N_5043,N_319,N_1460);
nand U5044 (N_5044,N_173,N_2013);
xor U5045 (N_5045,N_1493,N_2675);
and U5046 (N_5046,N_2157,N_2305);
or U5047 (N_5047,N_1794,N_514);
or U5048 (N_5048,N_237,N_1754);
and U5049 (N_5049,N_2927,N_1114);
nand U5050 (N_5050,N_2218,N_1037);
xnor U5051 (N_5051,N_2116,N_934);
and U5052 (N_5052,N_2539,N_2621);
and U5053 (N_5053,N_2101,N_1587);
or U5054 (N_5054,N_1143,N_2877);
xnor U5055 (N_5055,N_789,N_679);
nor U5056 (N_5056,N_1890,N_2019);
nor U5057 (N_5057,N_2152,N_1179);
xnor U5058 (N_5058,N_2419,N_2115);
xor U5059 (N_5059,N_1758,N_707);
and U5060 (N_5060,N_381,N_1392);
xnor U5061 (N_5061,N_1421,N_2852);
xnor U5062 (N_5062,N_2845,N_1826);
xor U5063 (N_5063,N_147,N_297);
xor U5064 (N_5064,N_1230,N_2267);
nor U5065 (N_5065,N_1266,N_2878);
nor U5066 (N_5066,N_1840,N_776);
nand U5067 (N_5067,N_423,N_1339);
nor U5068 (N_5068,N_374,N_1130);
nor U5069 (N_5069,N_1899,N_214);
or U5070 (N_5070,N_2220,N_1155);
and U5071 (N_5071,N_714,N_2597);
xor U5072 (N_5072,N_2863,N_2596);
and U5073 (N_5073,N_2073,N_2220);
xor U5074 (N_5074,N_2410,N_2542);
nor U5075 (N_5075,N_1536,N_525);
and U5076 (N_5076,N_1099,N_2283);
xnor U5077 (N_5077,N_1007,N_2848);
xnor U5078 (N_5078,N_629,N_2053);
nand U5079 (N_5079,N_2532,N_2733);
or U5080 (N_5080,N_1535,N_1210);
xnor U5081 (N_5081,N_2051,N_1996);
or U5082 (N_5082,N_2730,N_1548);
or U5083 (N_5083,N_2942,N_833);
xor U5084 (N_5084,N_2124,N_1044);
nor U5085 (N_5085,N_2922,N_2159);
and U5086 (N_5086,N_458,N_1663);
or U5087 (N_5087,N_2112,N_1475);
nand U5088 (N_5088,N_947,N_1891);
and U5089 (N_5089,N_2276,N_390);
or U5090 (N_5090,N_337,N_2499);
and U5091 (N_5091,N_2901,N_109);
and U5092 (N_5092,N_956,N_2345);
nor U5093 (N_5093,N_1938,N_2250);
and U5094 (N_5094,N_2240,N_768);
xnor U5095 (N_5095,N_493,N_2216);
xor U5096 (N_5096,N_1615,N_1633);
xor U5097 (N_5097,N_483,N_2460);
or U5098 (N_5098,N_855,N_2637);
nand U5099 (N_5099,N_2429,N_2601);
or U5100 (N_5100,N_1462,N_1995);
or U5101 (N_5101,N_2445,N_1545);
nand U5102 (N_5102,N_1209,N_1124);
nand U5103 (N_5103,N_1273,N_1798);
nand U5104 (N_5104,N_2995,N_1182);
or U5105 (N_5105,N_2508,N_450);
and U5106 (N_5106,N_1135,N_2355);
and U5107 (N_5107,N_1025,N_37);
nor U5108 (N_5108,N_558,N_1228);
nand U5109 (N_5109,N_1323,N_2456);
or U5110 (N_5110,N_2687,N_17);
and U5111 (N_5111,N_1781,N_2385);
or U5112 (N_5112,N_1273,N_1143);
and U5113 (N_5113,N_1822,N_538);
nor U5114 (N_5114,N_2302,N_1203);
xnor U5115 (N_5115,N_1771,N_665);
nor U5116 (N_5116,N_2670,N_2662);
nor U5117 (N_5117,N_2501,N_1777);
and U5118 (N_5118,N_2815,N_2003);
nand U5119 (N_5119,N_1731,N_616);
xnor U5120 (N_5120,N_2849,N_608);
and U5121 (N_5121,N_1715,N_793);
nand U5122 (N_5122,N_318,N_958);
and U5123 (N_5123,N_2450,N_2344);
and U5124 (N_5124,N_2945,N_1626);
xnor U5125 (N_5125,N_1305,N_255);
nand U5126 (N_5126,N_133,N_2231);
nor U5127 (N_5127,N_2432,N_1022);
and U5128 (N_5128,N_1866,N_323);
and U5129 (N_5129,N_2959,N_2580);
and U5130 (N_5130,N_1213,N_2254);
xnor U5131 (N_5131,N_951,N_1883);
or U5132 (N_5132,N_328,N_2509);
xor U5133 (N_5133,N_319,N_1035);
nor U5134 (N_5134,N_1430,N_305);
and U5135 (N_5135,N_2157,N_255);
nand U5136 (N_5136,N_2244,N_2535);
nor U5137 (N_5137,N_1618,N_1351);
or U5138 (N_5138,N_1180,N_783);
xor U5139 (N_5139,N_2445,N_1187);
nor U5140 (N_5140,N_1371,N_1959);
or U5141 (N_5141,N_255,N_1009);
or U5142 (N_5142,N_866,N_2151);
nor U5143 (N_5143,N_680,N_2247);
nand U5144 (N_5144,N_1539,N_511);
xor U5145 (N_5145,N_1935,N_525);
or U5146 (N_5146,N_1116,N_2973);
or U5147 (N_5147,N_2536,N_985);
xnor U5148 (N_5148,N_2561,N_945);
nor U5149 (N_5149,N_2096,N_2219);
nand U5150 (N_5150,N_1206,N_2227);
xor U5151 (N_5151,N_1890,N_1622);
and U5152 (N_5152,N_2373,N_867);
nor U5153 (N_5153,N_1051,N_1270);
and U5154 (N_5154,N_1935,N_1303);
or U5155 (N_5155,N_2322,N_2335);
or U5156 (N_5156,N_2525,N_812);
and U5157 (N_5157,N_525,N_1671);
xor U5158 (N_5158,N_796,N_2077);
nand U5159 (N_5159,N_1425,N_1374);
nand U5160 (N_5160,N_914,N_1993);
xnor U5161 (N_5161,N_892,N_1996);
or U5162 (N_5162,N_514,N_2282);
nand U5163 (N_5163,N_590,N_1191);
or U5164 (N_5164,N_929,N_442);
nand U5165 (N_5165,N_2968,N_1719);
xnor U5166 (N_5166,N_2657,N_2906);
or U5167 (N_5167,N_1432,N_808);
and U5168 (N_5168,N_652,N_2632);
nand U5169 (N_5169,N_2407,N_2934);
and U5170 (N_5170,N_234,N_1714);
and U5171 (N_5171,N_888,N_2336);
and U5172 (N_5172,N_2698,N_2577);
nor U5173 (N_5173,N_2610,N_2813);
and U5174 (N_5174,N_1747,N_2116);
xnor U5175 (N_5175,N_1349,N_299);
nand U5176 (N_5176,N_2907,N_1235);
or U5177 (N_5177,N_911,N_2261);
and U5178 (N_5178,N_948,N_1181);
nand U5179 (N_5179,N_421,N_2060);
xnor U5180 (N_5180,N_1891,N_2155);
or U5181 (N_5181,N_2568,N_2941);
and U5182 (N_5182,N_2063,N_2602);
xor U5183 (N_5183,N_1351,N_2982);
xnor U5184 (N_5184,N_1694,N_29);
nor U5185 (N_5185,N_288,N_2189);
nor U5186 (N_5186,N_2646,N_2020);
nor U5187 (N_5187,N_1699,N_2207);
nor U5188 (N_5188,N_2954,N_2721);
nor U5189 (N_5189,N_1139,N_2667);
nand U5190 (N_5190,N_2946,N_1936);
nor U5191 (N_5191,N_2255,N_2647);
nor U5192 (N_5192,N_2732,N_100);
nor U5193 (N_5193,N_2172,N_1020);
and U5194 (N_5194,N_282,N_201);
and U5195 (N_5195,N_2388,N_1352);
nand U5196 (N_5196,N_2922,N_844);
nand U5197 (N_5197,N_1707,N_1804);
or U5198 (N_5198,N_232,N_609);
or U5199 (N_5199,N_1505,N_2427);
or U5200 (N_5200,N_1288,N_334);
xnor U5201 (N_5201,N_1650,N_1310);
nand U5202 (N_5202,N_1511,N_730);
nand U5203 (N_5203,N_41,N_1193);
or U5204 (N_5204,N_2125,N_2471);
or U5205 (N_5205,N_2733,N_333);
and U5206 (N_5206,N_795,N_1354);
or U5207 (N_5207,N_2978,N_1365);
and U5208 (N_5208,N_2086,N_1115);
and U5209 (N_5209,N_1049,N_2768);
xnor U5210 (N_5210,N_706,N_2347);
or U5211 (N_5211,N_453,N_2824);
xor U5212 (N_5212,N_676,N_2714);
or U5213 (N_5213,N_2152,N_1282);
or U5214 (N_5214,N_2305,N_2531);
nor U5215 (N_5215,N_2279,N_1647);
xnor U5216 (N_5216,N_2479,N_2743);
or U5217 (N_5217,N_1441,N_2178);
nor U5218 (N_5218,N_1238,N_930);
or U5219 (N_5219,N_2450,N_511);
nor U5220 (N_5220,N_103,N_361);
nor U5221 (N_5221,N_1749,N_2085);
nor U5222 (N_5222,N_2218,N_164);
xnor U5223 (N_5223,N_412,N_2007);
or U5224 (N_5224,N_456,N_2337);
or U5225 (N_5225,N_451,N_1728);
nor U5226 (N_5226,N_1793,N_193);
and U5227 (N_5227,N_1767,N_1620);
nand U5228 (N_5228,N_107,N_838);
nand U5229 (N_5229,N_2159,N_1459);
nor U5230 (N_5230,N_617,N_1483);
nor U5231 (N_5231,N_1724,N_2460);
or U5232 (N_5232,N_1024,N_2141);
xnor U5233 (N_5233,N_2288,N_1002);
and U5234 (N_5234,N_714,N_1558);
and U5235 (N_5235,N_1924,N_1153);
nor U5236 (N_5236,N_2042,N_473);
nor U5237 (N_5237,N_2887,N_1528);
and U5238 (N_5238,N_1994,N_765);
xor U5239 (N_5239,N_420,N_2476);
and U5240 (N_5240,N_2979,N_1573);
xnor U5241 (N_5241,N_1657,N_2339);
nor U5242 (N_5242,N_2661,N_1654);
or U5243 (N_5243,N_1094,N_2302);
xor U5244 (N_5244,N_1189,N_187);
and U5245 (N_5245,N_1943,N_556);
or U5246 (N_5246,N_2922,N_260);
nor U5247 (N_5247,N_1935,N_297);
and U5248 (N_5248,N_2771,N_1387);
xnor U5249 (N_5249,N_1770,N_1143);
nand U5250 (N_5250,N_1315,N_2894);
nor U5251 (N_5251,N_943,N_770);
xor U5252 (N_5252,N_1025,N_2392);
nand U5253 (N_5253,N_604,N_2832);
or U5254 (N_5254,N_327,N_1265);
nor U5255 (N_5255,N_1492,N_415);
nand U5256 (N_5256,N_1163,N_2204);
and U5257 (N_5257,N_2235,N_35);
and U5258 (N_5258,N_2384,N_874);
xor U5259 (N_5259,N_932,N_277);
xnor U5260 (N_5260,N_1389,N_477);
or U5261 (N_5261,N_1019,N_1354);
xnor U5262 (N_5262,N_415,N_1229);
nand U5263 (N_5263,N_387,N_555);
or U5264 (N_5264,N_514,N_2232);
nand U5265 (N_5265,N_919,N_2245);
nand U5266 (N_5266,N_1139,N_2152);
and U5267 (N_5267,N_768,N_517);
and U5268 (N_5268,N_1391,N_787);
nor U5269 (N_5269,N_2871,N_1143);
nor U5270 (N_5270,N_423,N_2862);
nor U5271 (N_5271,N_1060,N_2168);
nand U5272 (N_5272,N_915,N_2428);
nor U5273 (N_5273,N_2179,N_1924);
nor U5274 (N_5274,N_735,N_2899);
or U5275 (N_5275,N_751,N_1156);
and U5276 (N_5276,N_614,N_500);
or U5277 (N_5277,N_1090,N_1545);
or U5278 (N_5278,N_1610,N_1212);
nor U5279 (N_5279,N_2346,N_766);
nand U5280 (N_5280,N_808,N_384);
or U5281 (N_5281,N_1998,N_419);
and U5282 (N_5282,N_701,N_2642);
and U5283 (N_5283,N_1081,N_2605);
nand U5284 (N_5284,N_1490,N_2681);
nand U5285 (N_5285,N_1533,N_965);
nand U5286 (N_5286,N_1391,N_1988);
or U5287 (N_5287,N_2909,N_53);
or U5288 (N_5288,N_2851,N_2200);
or U5289 (N_5289,N_1113,N_2944);
xor U5290 (N_5290,N_2065,N_1703);
nand U5291 (N_5291,N_586,N_354);
nand U5292 (N_5292,N_2857,N_310);
nor U5293 (N_5293,N_1609,N_1234);
nor U5294 (N_5294,N_755,N_1713);
and U5295 (N_5295,N_2459,N_1935);
or U5296 (N_5296,N_1478,N_1463);
xor U5297 (N_5297,N_2360,N_331);
xor U5298 (N_5298,N_739,N_1663);
or U5299 (N_5299,N_849,N_602);
nand U5300 (N_5300,N_2225,N_38);
and U5301 (N_5301,N_2120,N_2495);
or U5302 (N_5302,N_2604,N_2589);
and U5303 (N_5303,N_1389,N_2044);
xor U5304 (N_5304,N_2666,N_916);
nand U5305 (N_5305,N_538,N_198);
and U5306 (N_5306,N_834,N_559);
xnor U5307 (N_5307,N_2671,N_1782);
nand U5308 (N_5308,N_1213,N_1148);
nor U5309 (N_5309,N_2289,N_2066);
nor U5310 (N_5310,N_1507,N_2766);
xor U5311 (N_5311,N_580,N_444);
and U5312 (N_5312,N_496,N_2430);
nand U5313 (N_5313,N_1046,N_1326);
nand U5314 (N_5314,N_825,N_2667);
nor U5315 (N_5315,N_1030,N_74);
xnor U5316 (N_5316,N_95,N_540);
nand U5317 (N_5317,N_60,N_960);
or U5318 (N_5318,N_1756,N_1709);
nand U5319 (N_5319,N_1975,N_403);
or U5320 (N_5320,N_2630,N_1930);
xnor U5321 (N_5321,N_1458,N_260);
nor U5322 (N_5322,N_2620,N_2234);
nor U5323 (N_5323,N_377,N_2414);
nand U5324 (N_5324,N_1012,N_1032);
nor U5325 (N_5325,N_2207,N_2558);
nand U5326 (N_5326,N_2582,N_1537);
nand U5327 (N_5327,N_1601,N_1701);
nand U5328 (N_5328,N_154,N_1344);
or U5329 (N_5329,N_671,N_1526);
nor U5330 (N_5330,N_1842,N_2800);
nor U5331 (N_5331,N_1170,N_1196);
xor U5332 (N_5332,N_1364,N_2168);
xor U5333 (N_5333,N_1544,N_410);
and U5334 (N_5334,N_1208,N_217);
xor U5335 (N_5335,N_790,N_467);
or U5336 (N_5336,N_1254,N_175);
nand U5337 (N_5337,N_1777,N_745);
nand U5338 (N_5338,N_2354,N_139);
xnor U5339 (N_5339,N_987,N_1239);
xnor U5340 (N_5340,N_2298,N_2730);
and U5341 (N_5341,N_1748,N_1051);
xor U5342 (N_5342,N_1341,N_834);
nand U5343 (N_5343,N_1376,N_2854);
nor U5344 (N_5344,N_1093,N_604);
nand U5345 (N_5345,N_747,N_387);
xor U5346 (N_5346,N_1851,N_2678);
and U5347 (N_5347,N_2746,N_100);
nor U5348 (N_5348,N_2284,N_1884);
nor U5349 (N_5349,N_2037,N_533);
or U5350 (N_5350,N_2332,N_286);
or U5351 (N_5351,N_1947,N_1840);
and U5352 (N_5352,N_557,N_2600);
or U5353 (N_5353,N_917,N_2378);
xnor U5354 (N_5354,N_552,N_1651);
nor U5355 (N_5355,N_117,N_2133);
nor U5356 (N_5356,N_566,N_1851);
xor U5357 (N_5357,N_922,N_2394);
or U5358 (N_5358,N_226,N_1923);
nor U5359 (N_5359,N_579,N_1320);
xnor U5360 (N_5360,N_1146,N_2577);
xnor U5361 (N_5361,N_2277,N_2024);
and U5362 (N_5362,N_263,N_312);
or U5363 (N_5363,N_764,N_1300);
xnor U5364 (N_5364,N_860,N_728);
and U5365 (N_5365,N_1819,N_727);
xor U5366 (N_5366,N_652,N_1603);
nand U5367 (N_5367,N_1020,N_185);
nand U5368 (N_5368,N_1068,N_1123);
nand U5369 (N_5369,N_1101,N_2852);
xnor U5370 (N_5370,N_377,N_2490);
or U5371 (N_5371,N_880,N_1484);
nand U5372 (N_5372,N_2068,N_2909);
xnor U5373 (N_5373,N_327,N_977);
and U5374 (N_5374,N_2204,N_1871);
xor U5375 (N_5375,N_682,N_2965);
and U5376 (N_5376,N_1140,N_1262);
xor U5377 (N_5377,N_1081,N_2742);
nand U5378 (N_5378,N_1033,N_592);
or U5379 (N_5379,N_132,N_2966);
xor U5380 (N_5380,N_1842,N_1358);
xnor U5381 (N_5381,N_903,N_2146);
or U5382 (N_5382,N_1181,N_1292);
or U5383 (N_5383,N_1450,N_2395);
or U5384 (N_5384,N_2044,N_1273);
nor U5385 (N_5385,N_1534,N_2036);
xor U5386 (N_5386,N_2906,N_1202);
and U5387 (N_5387,N_623,N_521);
xnor U5388 (N_5388,N_914,N_1325);
nor U5389 (N_5389,N_2034,N_785);
nor U5390 (N_5390,N_1899,N_1283);
or U5391 (N_5391,N_706,N_2982);
nand U5392 (N_5392,N_2472,N_1308);
nand U5393 (N_5393,N_1847,N_1518);
nor U5394 (N_5394,N_1114,N_2607);
and U5395 (N_5395,N_2028,N_659);
nor U5396 (N_5396,N_2194,N_2781);
nand U5397 (N_5397,N_1916,N_2451);
or U5398 (N_5398,N_2220,N_987);
or U5399 (N_5399,N_1399,N_1071);
xnor U5400 (N_5400,N_2834,N_2735);
nand U5401 (N_5401,N_1243,N_1860);
xor U5402 (N_5402,N_2274,N_115);
or U5403 (N_5403,N_682,N_1863);
or U5404 (N_5404,N_2022,N_2351);
and U5405 (N_5405,N_2802,N_399);
xor U5406 (N_5406,N_1409,N_1105);
nand U5407 (N_5407,N_2455,N_210);
nor U5408 (N_5408,N_783,N_2493);
xor U5409 (N_5409,N_1020,N_1978);
xnor U5410 (N_5410,N_484,N_296);
nand U5411 (N_5411,N_790,N_1467);
nor U5412 (N_5412,N_212,N_2001);
or U5413 (N_5413,N_1951,N_286);
xnor U5414 (N_5414,N_1194,N_1766);
or U5415 (N_5415,N_383,N_185);
nand U5416 (N_5416,N_911,N_560);
or U5417 (N_5417,N_1352,N_726);
or U5418 (N_5418,N_2514,N_302);
and U5419 (N_5419,N_2194,N_2698);
nor U5420 (N_5420,N_2938,N_322);
and U5421 (N_5421,N_1788,N_854);
nand U5422 (N_5422,N_230,N_1011);
nor U5423 (N_5423,N_2557,N_1621);
or U5424 (N_5424,N_885,N_2898);
xor U5425 (N_5425,N_1753,N_2288);
or U5426 (N_5426,N_648,N_1709);
and U5427 (N_5427,N_2563,N_1691);
or U5428 (N_5428,N_2255,N_2832);
and U5429 (N_5429,N_1495,N_2385);
nor U5430 (N_5430,N_2638,N_748);
xnor U5431 (N_5431,N_1623,N_2492);
nor U5432 (N_5432,N_2197,N_311);
nor U5433 (N_5433,N_1086,N_1701);
or U5434 (N_5434,N_834,N_2892);
and U5435 (N_5435,N_411,N_1320);
or U5436 (N_5436,N_1166,N_767);
nor U5437 (N_5437,N_2493,N_1070);
nand U5438 (N_5438,N_114,N_597);
or U5439 (N_5439,N_2555,N_1837);
nand U5440 (N_5440,N_2877,N_2611);
nor U5441 (N_5441,N_706,N_2529);
or U5442 (N_5442,N_135,N_878);
nand U5443 (N_5443,N_2719,N_1141);
nand U5444 (N_5444,N_2234,N_1359);
nor U5445 (N_5445,N_373,N_254);
nand U5446 (N_5446,N_2093,N_2890);
nor U5447 (N_5447,N_1142,N_1979);
or U5448 (N_5448,N_1043,N_2649);
nand U5449 (N_5449,N_1754,N_2988);
nor U5450 (N_5450,N_712,N_2157);
and U5451 (N_5451,N_1802,N_480);
or U5452 (N_5452,N_2370,N_1495);
or U5453 (N_5453,N_1042,N_1683);
nor U5454 (N_5454,N_2302,N_2319);
nand U5455 (N_5455,N_2945,N_687);
xor U5456 (N_5456,N_1503,N_2969);
or U5457 (N_5457,N_2034,N_1409);
and U5458 (N_5458,N_756,N_2026);
xnor U5459 (N_5459,N_2446,N_1309);
xor U5460 (N_5460,N_27,N_563);
xor U5461 (N_5461,N_1051,N_1327);
or U5462 (N_5462,N_1597,N_352);
nor U5463 (N_5463,N_1845,N_558);
nand U5464 (N_5464,N_358,N_626);
and U5465 (N_5465,N_2299,N_2507);
xnor U5466 (N_5466,N_1623,N_1113);
xor U5467 (N_5467,N_497,N_2325);
and U5468 (N_5468,N_2314,N_2282);
and U5469 (N_5469,N_1719,N_2065);
or U5470 (N_5470,N_1744,N_811);
or U5471 (N_5471,N_2738,N_1452);
and U5472 (N_5472,N_2294,N_2596);
nand U5473 (N_5473,N_1624,N_823);
xnor U5474 (N_5474,N_1917,N_2460);
nor U5475 (N_5475,N_940,N_2766);
or U5476 (N_5476,N_8,N_1701);
and U5477 (N_5477,N_2024,N_2267);
xnor U5478 (N_5478,N_1077,N_674);
nand U5479 (N_5479,N_2855,N_1729);
nand U5480 (N_5480,N_808,N_1602);
xor U5481 (N_5481,N_2931,N_1130);
or U5482 (N_5482,N_2508,N_1303);
nand U5483 (N_5483,N_2273,N_1938);
and U5484 (N_5484,N_188,N_1775);
and U5485 (N_5485,N_1867,N_591);
nor U5486 (N_5486,N_223,N_864);
nor U5487 (N_5487,N_1248,N_2340);
xnor U5488 (N_5488,N_280,N_683);
nand U5489 (N_5489,N_1838,N_2495);
nor U5490 (N_5490,N_1902,N_1867);
or U5491 (N_5491,N_1484,N_2194);
xor U5492 (N_5492,N_2092,N_2621);
nand U5493 (N_5493,N_1944,N_2772);
or U5494 (N_5494,N_2313,N_2845);
and U5495 (N_5495,N_729,N_2541);
and U5496 (N_5496,N_2510,N_1776);
nand U5497 (N_5497,N_614,N_993);
or U5498 (N_5498,N_2323,N_649);
nor U5499 (N_5499,N_1510,N_2389);
nor U5500 (N_5500,N_1778,N_555);
xnor U5501 (N_5501,N_2068,N_668);
or U5502 (N_5502,N_286,N_2072);
xor U5503 (N_5503,N_1240,N_1922);
or U5504 (N_5504,N_505,N_2963);
and U5505 (N_5505,N_1202,N_1493);
or U5506 (N_5506,N_2380,N_1565);
xor U5507 (N_5507,N_1591,N_676);
and U5508 (N_5508,N_2229,N_1280);
nand U5509 (N_5509,N_2209,N_1678);
and U5510 (N_5510,N_2991,N_1009);
xor U5511 (N_5511,N_1525,N_1309);
xor U5512 (N_5512,N_2978,N_2240);
nor U5513 (N_5513,N_1734,N_1379);
xnor U5514 (N_5514,N_1429,N_571);
or U5515 (N_5515,N_1749,N_1247);
nor U5516 (N_5516,N_1530,N_2590);
nor U5517 (N_5517,N_2593,N_2825);
xor U5518 (N_5518,N_977,N_2597);
xor U5519 (N_5519,N_2867,N_1456);
xnor U5520 (N_5520,N_1134,N_962);
or U5521 (N_5521,N_1522,N_2383);
and U5522 (N_5522,N_1189,N_2164);
nor U5523 (N_5523,N_2774,N_1937);
and U5524 (N_5524,N_1986,N_2150);
or U5525 (N_5525,N_2734,N_352);
nor U5526 (N_5526,N_1441,N_838);
nand U5527 (N_5527,N_1603,N_143);
and U5528 (N_5528,N_2299,N_1796);
or U5529 (N_5529,N_2504,N_2587);
nand U5530 (N_5530,N_718,N_49);
and U5531 (N_5531,N_447,N_2897);
nor U5532 (N_5532,N_1828,N_1172);
nor U5533 (N_5533,N_2696,N_1707);
or U5534 (N_5534,N_2456,N_2472);
nand U5535 (N_5535,N_405,N_1127);
nor U5536 (N_5536,N_2603,N_462);
xnor U5537 (N_5537,N_851,N_700);
nor U5538 (N_5538,N_2502,N_2192);
xnor U5539 (N_5539,N_1966,N_1395);
or U5540 (N_5540,N_265,N_2297);
nand U5541 (N_5541,N_268,N_2671);
nand U5542 (N_5542,N_2663,N_191);
and U5543 (N_5543,N_2609,N_1913);
and U5544 (N_5544,N_1825,N_2212);
nor U5545 (N_5545,N_2092,N_1207);
nor U5546 (N_5546,N_520,N_361);
nand U5547 (N_5547,N_75,N_627);
xnor U5548 (N_5548,N_605,N_1869);
xnor U5549 (N_5549,N_1981,N_2874);
and U5550 (N_5550,N_2533,N_1818);
nor U5551 (N_5551,N_1396,N_1016);
xor U5552 (N_5552,N_520,N_1123);
and U5553 (N_5553,N_2340,N_2706);
and U5554 (N_5554,N_1232,N_1377);
or U5555 (N_5555,N_2087,N_934);
xnor U5556 (N_5556,N_446,N_1190);
and U5557 (N_5557,N_884,N_1631);
and U5558 (N_5558,N_2421,N_1961);
xnor U5559 (N_5559,N_2718,N_463);
or U5560 (N_5560,N_2097,N_2556);
and U5561 (N_5561,N_1676,N_890);
nor U5562 (N_5562,N_1961,N_1667);
nand U5563 (N_5563,N_1715,N_2447);
nand U5564 (N_5564,N_116,N_1804);
and U5565 (N_5565,N_919,N_853);
xnor U5566 (N_5566,N_1995,N_521);
nand U5567 (N_5567,N_1626,N_2462);
nor U5568 (N_5568,N_183,N_1590);
xnor U5569 (N_5569,N_961,N_541);
nor U5570 (N_5570,N_442,N_2406);
xor U5571 (N_5571,N_1444,N_2761);
and U5572 (N_5572,N_2103,N_222);
xnor U5573 (N_5573,N_2295,N_2883);
xor U5574 (N_5574,N_1977,N_2313);
or U5575 (N_5575,N_530,N_2862);
xnor U5576 (N_5576,N_2063,N_860);
xnor U5577 (N_5577,N_183,N_1037);
xnor U5578 (N_5578,N_2921,N_2810);
nand U5579 (N_5579,N_173,N_212);
nor U5580 (N_5580,N_1286,N_2932);
nand U5581 (N_5581,N_1381,N_2271);
and U5582 (N_5582,N_574,N_641);
or U5583 (N_5583,N_436,N_1177);
nand U5584 (N_5584,N_2591,N_1654);
nand U5585 (N_5585,N_2975,N_1633);
or U5586 (N_5586,N_2703,N_2505);
nor U5587 (N_5587,N_2650,N_2882);
nand U5588 (N_5588,N_1347,N_2838);
and U5589 (N_5589,N_249,N_1100);
nor U5590 (N_5590,N_351,N_1788);
nand U5591 (N_5591,N_122,N_1234);
nand U5592 (N_5592,N_1552,N_2291);
xor U5593 (N_5593,N_753,N_2444);
xor U5594 (N_5594,N_1268,N_1995);
and U5595 (N_5595,N_2603,N_536);
nor U5596 (N_5596,N_247,N_336);
and U5597 (N_5597,N_1186,N_2747);
xnor U5598 (N_5598,N_979,N_1119);
or U5599 (N_5599,N_749,N_1308);
or U5600 (N_5600,N_2310,N_1521);
and U5601 (N_5601,N_2272,N_1545);
nand U5602 (N_5602,N_115,N_2138);
xnor U5603 (N_5603,N_1038,N_1247);
xnor U5604 (N_5604,N_1454,N_1185);
nand U5605 (N_5605,N_1753,N_2977);
and U5606 (N_5606,N_160,N_2115);
and U5607 (N_5607,N_740,N_554);
xor U5608 (N_5608,N_2067,N_1584);
nor U5609 (N_5609,N_568,N_1554);
and U5610 (N_5610,N_1572,N_296);
or U5611 (N_5611,N_1769,N_132);
nand U5612 (N_5612,N_2947,N_963);
nand U5613 (N_5613,N_394,N_2134);
and U5614 (N_5614,N_2237,N_138);
nand U5615 (N_5615,N_423,N_1329);
xnor U5616 (N_5616,N_2407,N_381);
or U5617 (N_5617,N_361,N_1960);
xnor U5618 (N_5618,N_2494,N_2490);
and U5619 (N_5619,N_2492,N_216);
and U5620 (N_5620,N_1091,N_695);
and U5621 (N_5621,N_498,N_1141);
nand U5622 (N_5622,N_1359,N_1033);
nand U5623 (N_5623,N_2705,N_773);
xnor U5624 (N_5624,N_905,N_1033);
xnor U5625 (N_5625,N_889,N_2228);
xor U5626 (N_5626,N_108,N_2638);
nand U5627 (N_5627,N_1878,N_528);
nor U5628 (N_5628,N_1540,N_2929);
nor U5629 (N_5629,N_1389,N_2647);
nor U5630 (N_5630,N_195,N_1685);
or U5631 (N_5631,N_70,N_2665);
nor U5632 (N_5632,N_840,N_281);
or U5633 (N_5633,N_865,N_945);
nand U5634 (N_5634,N_1107,N_1985);
or U5635 (N_5635,N_438,N_898);
xor U5636 (N_5636,N_1402,N_923);
nand U5637 (N_5637,N_2600,N_153);
and U5638 (N_5638,N_2239,N_951);
nand U5639 (N_5639,N_2395,N_1806);
xnor U5640 (N_5640,N_527,N_1257);
and U5641 (N_5641,N_636,N_52);
or U5642 (N_5642,N_1993,N_2275);
and U5643 (N_5643,N_2979,N_2940);
xor U5644 (N_5644,N_2007,N_2810);
or U5645 (N_5645,N_871,N_934);
nor U5646 (N_5646,N_282,N_1146);
nor U5647 (N_5647,N_1830,N_976);
xor U5648 (N_5648,N_130,N_1602);
or U5649 (N_5649,N_2523,N_2597);
nor U5650 (N_5650,N_893,N_2143);
or U5651 (N_5651,N_1377,N_1024);
xor U5652 (N_5652,N_850,N_1445);
xnor U5653 (N_5653,N_2070,N_342);
xor U5654 (N_5654,N_2450,N_287);
or U5655 (N_5655,N_863,N_2428);
xnor U5656 (N_5656,N_2378,N_20);
nor U5657 (N_5657,N_1171,N_415);
xor U5658 (N_5658,N_1271,N_2797);
nor U5659 (N_5659,N_1210,N_502);
nand U5660 (N_5660,N_2806,N_2711);
nand U5661 (N_5661,N_384,N_1018);
and U5662 (N_5662,N_2100,N_670);
and U5663 (N_5663,N_2293,N_1715);
xnor U5664 (N_5664,N_656,N_1243);
nor U5665 (N_5665,N_352,N_371);
and U5666 (N_5666,N_62,N_673);
and U5667 (N_5667,N_2393,N_1975);
and U5668 (N_5668,N_2691,N_2727);
or U5669 (N_5669,N_239,N_1377);
xor U5670 (N_5670,N_2000,N_874);
nand U5671 (N_5671,N_1515,N_840);
or U5672 (N_5672,N_2146,N_979);
nor U5673 (N_5673,N_176,N_345);
and U5674 (N_5674,N_139,N_1273);
and U5675 (N_5675,N_1919,N_2935);
or U5676 (N_5676,N_1070,N_161);
xor U5677 (N_5677,N_119,N_295);
nand U5678 (N_5678,N_106,N_2722);
and U5679 (N_5679,N_1272,N_465);
xnor U5680 (N_5680,N_158,N_17);
nand U5681 (N_5681,N_1898,N_2864);
nand U5682 (N_5682,N_2141,N_2331);
xor U5683 (N_5683,N_1994,N_1993);
nand U5684 (N_5684,N_2181,N_2771);
xor U5685 (N_5685,N_563,N_938);
and U5686 (N_5686,N_2983,N_2952);
nand U5687 (N_5687,N_2221,N_1716);
and U5688 (N_5688,N_1105,N_1717);
xor U5689 (N_5689,N_349,N_2314);
nand U5690 (N_5690,N_345,N_1018);
or U5691 (N_5691,N_92,N_568);
and U5692 (N_5692,N_1381,N_1181);
or U5693 (N_5693,N_1787,N_1838);
nand U5694 (N_5694,N_858,N_713);
nor U5695 (N_5695,N_1233,N_2831);
nor U5696 (N_5696,N_2021,N_284);
or U5697 (N_5697,N_206,N_257);
nand U5698 (N_5698,N_1560,N_1785);
nor U5699 (N_5699,N_954,N_2045);
nor U5700 (N_5700,N_1072,N_1841);
or U5701 (N_5701,N_487,N_1344);
nand U5702 (N_5702,N_88,N_1738);
xor U5703 (N_5703,N_60,N_487);
nor U5704 (N_5704,N_1056,N_1222);
xnor U5705 (N_5705,N_2361,N_2692);
nor U5706 (N_5706,N_2678,N_273);
or U5707 (N_5707,N_2654,N_434);
or U5708 (N_5708,N_724,N_246);
and U5709 (N_5709,N_2346,N_1663);
nor U5710 (N_5710,N_1477,N_1988);
nor U5711 (N_5711,N_2386,N_2974);
xor U5712 (N_5712,N_2651,N_1494);
or U5713 (N_5713,N_1575,N_1455);
and U5714 (N_5714,N_1652,N_2688);
xor U5715 (N_5715,N_2007,N_823);
xor U5716 (N_5716,N_456,N_2028);
xor U5717 (N_5717,N_20,N_947);
and U5718 (N_5718,N_657,N_2210);
nand U5719 (N_5719,N_1952,N_2493);
nor U5720 (N_5720,N_3,N_269);
nor U5721 (N_5721,N_1636,N_2490);
nor U5722 (N_5722,N_2660,N_2375);
and U5723 (N_5723,N_2424,N_969);
nor U5724 (N_5724,N_2634,N_1873);
nor U5725 (N_5725,N_1151,N_103);
nor U5726 (N_5726,N_1524,N_387);
and U5727 (N_5727,N_2542,N_247);
or U5728 (N_5728,N_2452,N_2696);
xnor U5729 (N_5729,N_2400,N_2416);
or U5730 (N_5730,N_391,N_2298);
nor U5731 (N_5731,N_2077,N_2153);
nand U5732 (N_5732,N_2169,N_192);
nor U5733 (N_5733,N_574,N_2360);
nand U5734 (N_5734,N_2570,N_2631);
nor U5735 (N_5735,N_479,N_1045);
nand U5736 (N_5736,N_232,N_1610);
nor U5737 (N_5737,N_189,N_412);
nand U5738 (N_5738,N_1408,N_2373);
nor U5739 (N_5739,N_2797,N_1940);
and U5740 (N_5740,N_2783,N_880);
xnor U5741 (N_5741,N_937,N_2637);
or U5742 (N_5742,N_1585,N_1309);
nand U5743 (N_5743,N_757,N_1648);
and U5744 (N_5744,N_1213,N_1015);
nor U5745 (N_5745,N_2278,N_2796);
xor U5746 (N_5746,N_170,N_2719);
or U5747 (N_5747,N_2847,N_1908);
or U5748 (N_5748,N_1654,N_2459);
nor U5749 (N_5749,N_726,N_920);
and U5750 (N_5750,N_1192,N_2992);
or U5751 (N_5751,N_1576,N_2265);
nand U5752 (N_5752,N_2945,N_1740);
or U5753 (N_5753,N_1509,N_2154);
nor U5754 (N_5754,N_1719,N_1204);
and U5755 (N_5755,N_2568,N_529);
xnor U5756 (N_5756,N_2678,N_775);
xnor U5757 (N_5757,N_2264,N_1237);
xor U5758 (N_5758,N_2160,N_1472);
xor U5759 (N_5759,N_1725,N_1858);
or U5760 (N_5760,N_2440,N_2148);
nor U5761 (N_5761,N_275,N_506);
nor U5762 (N_5762,N_88,N_1708);
nor U5763 (N_5763,N_2018,N_2723);
nor U5764 (N_5764,N_2777,N_2183);
nand U5765 (N_5765,N_2300,N_1577);
or U5766 (N_5766,N_974,N_1987);
nor U5767 (N_5767,N_104,N_1575);
nand U5768 (N_5768,N_2389,N_88);
and U5769 (N_5769,N_2722,N_2687);
or U5770 (N_5770,N_1844,N_2441);
nor U5771 (N_5771,N_644,N_1405);
nand U5772 (N_5772,N_2816,N_1622);
and U5773 (N_5773,N_1073,N_1235);
or U5774 (N_5774,N_1241,N_1369);
xnor U5775 (N_5775,N_76,N_1449);
or U5776 (N_5776,N_2582,N_1084);
nor U5777 (N_5777,N_1908,N_2646);
and U5778 (N_5778,N_2609,N_554);
or U5779 (N_5779,N_1124,N_2325);
and U5780 (N_5780,N_2001,N_1625);
or U5781 (N_5781,N_1378,N_1163);
nand U5782 (N_5782,N_406,N_225);
nand U5783 (N_5783,N_2720,N_581);
nor U5784 (N_5784,N_1172,N_1806);
or U5785 (N_5785,N_1364,N_860);
nand U5786 (N_5786,N_474,N_2488);
or U5787 (N_5787,N_1915,N_1852);
or U5788 (N_5788,N_2915,N_2380);
xnor U5789 (N_5789,N_1288,N_1322);
and U5790 (N_5790,N_1569,N_1161);
nand U5791 (N_5791,N_1172,N_1148);
nor U5792 (N_5792,N_2025,N_962);
xor U5793 (N_5793,N_2650,N_2023);
nand U5794 (N_5794,N_2413,N_2786);
nor U5795 (N_5795,N_455,N_2587);
or U5796 (N_5796,N_1101,N_382);
or U5797 (N_5797,N_98,N_733);
and U5798 (N_5798,N_1777,N_2053);
or U5799 (N_5799,N_1272,N_183);
nor U5800 (N_5800,N_50,N_2121);
xnor U5801 (N_5801,N_15,N_933);
nand U5802 (N_5802,N_559,N_1393);
nor U5803 (N_5803,N_1339,N_2264);
or U5804 (N_5804,N_1310,N_2380);
nand U5805 (N_5805,N_1981,N_715);
xnor U5806 (N_5806,N_2719,N_1133);
and U5807 (N_5807,N_1107,N_176);
nand U5808 (N_5808,N_1036,N_277);
nand U5809 (N_5809,N_1144,N_292);
nor U5810 (N_5810,N_2440,N_252);
xnor U5811 (N_5811,N_2293,N_2656);
xor U5812 (N_5812,N_291,N_2116);
nand U5813 (N_5813,N_2607,N_1423);
nor U5814 (N_5814,N_2138,N_1528);
nor U5815 (N_5815,N_525,N_414);
nor U5816 (N_5816,N_0,N_363);
and U5817 (N_5817,N_113,N_1968);
nor U5818 (N_5818,N_169,N_2989);
or U5819 (N_5819,N_1971,N_1138);
or U5820 (N_5820,N_2821,N_2346);
and U5821 (N_5821,N_2846,N_1719);
nand U5822 (N_5822,N_1009,N_649);
and U5823 (N_5823,N_2643,N_2030);
nor U5824 (N_5824,N_865,N_2095);
xnor U5825 (N_5825,N_1119,N_992);
nand U5826 (N_5826,N_1616,N_1945);
or U5827 (N_5827,N_2735,N_2951);
nor U5828 (N_5828,N_1307,N_1159);
xor U5829 (N_5829,N_1360,N_1765);
xnor U5830 (N_5830,N_2670,N_1799);
xnor U5831 (N_5831,N_1285,N_941);
or U5832 (N_5832,N_2603,N_469);
nand U5833 (N_5833,N_110,N_1338);
nand U5834 (N_5834,N_184,N_2627);
nor U5835 (N_5835,N_1788,N_649);
and U5836 (N_5836,N_2415,N_16);
and U5837 (N_5837,N_2145,N_1276);
nor U5838 (N_5838,N_394,N_2022);
nand U5839 (N_5839,N_2925,N_2492);
nor U5840 (N_5840,N_816,N_1255);
xor U5841 (N_5841,N_2123,N_1957);
and U5842 (N_5842,N_102,N_1893);
nor U5843 (N_5843,N_1827,N_2874);
or U5844 (N_5844,N_2778,N_1923);
and U5845 (N_5845,N_1650,N_383);
and U5846 (N_5846,N_2970,N_877);
nor U5847 (N_5847,N_2350,N_565);
and U5848 (N_5848,N_727,N_591);
xnor U5849 (N_5849,N_2984,N_1619);
and U5850 (N_5850,N_38,N_1081);
nor U5851 (N_5851,N_2498,N_2357);
and U5852 (N_5852,N_1568,N_1962);
nand U5853 (N_5853,N_1302,N_2292);
nand U5854 (N_5854,N_579,N_1633);
xnor U5855 (N_5855,N_96,N_184);
nor U5856 (N_5856,N_2802,N_2808);
or U5857 (N_5857,N_994,N_593);
nand U5858 (N_5858,N_1521,N_2380);
and U5859 (N_5859,N_1637,N_2475);
nand U5860 (N_5860,N_2083,N_370);
xor U5861 (N_5861,N_282,N_2310);
nor U5862 (N_5862,N_1412,N_2467);
nand U5863 (N_5863,N_1028,N_609);
or U5864 (N_5864,N_265,N_2534);
nor U5865 (N_5865,N_2425,N_2889);
xnor U5866 (N_5866,N_139,N_944);
or U5867 (N_5867,N_495,N_2382);
nor U5868 (N_5868,N_962,N_354);
xor U5869 (N_5869,N_397,N_2430);
and U5870 (N_5870,N_2574,N_2784);
or U5871 (N_5871,N_81,N_2258);
xor U5872 (N_5872,N_954,N_1746);
xor U5873 (N_5873,N_2564,N_2258);
nand U5874 (N_5874,N_847,N_2855);
or U5875 (N_5875,N_2566,N_1735);
nand U5876 (N_5876,N_2313,N_768);
xor U5877 (N_5877,N_1046,N_758);
nor U5878 (N_5878,N_767,N_2440);
nor U5879 (N_5879,N_930,N_2524);
xor U5880 (N_5880,N_2897,N_2526);
xor U5881 (N_5881,N_553,N_228);
nor U5882 (N_5882,N_1024,N_1843);
xnor U5883 (N_5883,N_2730,N_968);
xor U5884 (N_5884,N_1793,N_2897);
and U5885 (N_5885,N_176,N_181);
and U5886 (N_5886,N_2620,N_298);
and U5887 (N_5887,N_89,N_848);
nand U5888 (N_5888,N_409,N_440);
nor U5889 (N_5889,N_149,N_2895);
nor U5890 (N_5890,N_455,N_1079);
xor U5891 (N_5891,N_2942,N_1463);
nand U5892 (N_5892,N_0,N_2263);
and U5893 (N_5893,N_950,N_1720);
xnor U5894 (N_5894,N_2484,N_1860);
xnor U5895 (N_5895,N_648,N_1796);
nor U5896 (N_5896,N_531,N_2101);
nor U5897 (N_5897,N_710,N_2803);
and U5898 (N_5898,N_814,N_775);
nor U5899 (N_5899,N_2010,N_2267);
and U5900 (N_5900,N_2873,N_656);
nand U5901 (N_5901,N_635,N_2853);
or U5902 (N_5902,N_1240,N_2498);
nand U5903 (N_5903,N_1829,N_503);
xor U5904 (N_5904,N_1417,N_1614);
nor U5905 (N_5905,N_2737,N_1400);
nand U5906 (N_5906,N_68,N_2034);
and U5907 (N_5907,N_2481,N_1809);
and U5908 (N_5908,N_739,N_513);
xor U5909 (N_5909,N_1936,N_1738);
and U5910 (N_5910,N_675,N_2285);
xor U5911 (N_5911,N_2519,N_1720);
and U5912 (N_5912,N_2943,N_468);
xor U5913 (N_5913,N_1443,N_270);
nor U5914 (N_5914,N_2647,N_56);
xnor U5915 (N_5915,N_2005,N_1935);
nand U5916 (N_5916,N_1347,N_498);
or U5917 (N_5917,N_2125,N_2005);
nor U5918 (N_5918,N_1169,N_2265);
or U5919 (N_5919,N_2134,N_1929);
nand U5920 (N_5920,N_652,N_163);
nand U5921 (N_5921,N_965,N_2517);
or U5922 (N_5922,N_1804,N_532);
xnor U5923 (N_5923,N_2098,N_729);
or U5924 (N_5924,N_2062,N_1310);
nand U5925 (N_5925,N_566,N_1630);
nand U5926 (N_5926,N_2060,N_180);
and U5927 (N_5927,N_642,N_1718);
nor U5928 (N_5928,N_1064,N_991);
or U5929 (N_5929,N_2801,N_2539);
nand U5930 (N_5930,N_1591,N_24);
or U5931 (N_5931,N_2792,N_2312);
xor U5932 (N_5932,N_2520,N_368);
or U5933 (N_5933,N_1782,N_1995);
nand U5934 (N_5934,N_1129,N_2181);
or U5935 (N_5935,N_2334,N_1458);
nor U5936 (N_5936,N_1199,N_2779);
and U5937 (N_5937,N_910,N_2167);
or U5938 (N_5938,N_1231,N_2750);
nor U5939 (N_5939,N_766,N_25);
or U5940 (N_5940,N_773,N_1710);
and U5941 (N_5941,N_961,N_2696);
nand U5942 (N_5942,N_1054,N_915);
xnor U5943 (N_5943,N_1650,N_35);
xnor U5944 (N_5944,N_1746,N_262);
and U5945 (N_5945,N_2262,N_1331);
nand U5946 (N_5946,N_564,N_628);
xor U5947 (N_5947,N_2774,N_123);
xor U5948 (N_5948,N_44,N_134);
nor U5949 (N_5949,N_863,N_1332);
and U5950 (N_5950,N_435,N_1275);
xnor U5951 (N_5951,N_2334,N_631);
nand U5952 (N_5952,N_2712,N_2630);
and U5953 (N_5953,N_1159,N_2689);
or U5954 (N_5954,N_2758,N_569);
or U5955 (N_5955,N_412,N_2807);
or U5956 (N_5956,N_2,N_1373);
nand U5957 (N_5957,N_238,N_1067);
nor U5958 (N_5958,N_89,N_1007);
nor U5959 (N_5959,N_386,N_38);
xnor U5960 (N_5960,N_1472,N_2861);
and U5961 (N_5961,N_171,N_2214);
xor U5962 (N_5962,N_1387,N_470);
nor U5963 (N_5963,N_1405,N_2584);
nand U5964 (N_5964,N_1756,N_2264);
xor U5965 (N_5965,N_1092,N_1964);
and U5966 (N_5966,N_68,N_764);
or U5967 (N_5967,N_2227,N_1643);
nor U5968 (N_5968,N_69,N_1874);
or U5969 (N_5969,N_1654,N_2727);
nor U5970 (N_5970,N_232,N_1962);
xnor U5971 (N_5971,N_782,N_2321);
xnor U5972 (N_5972,N_2619,N_1365);
and U5973 (N_5973,N_1332,N_2486);
nor U5974 (N_5974,N_2026,N_2781);
or U5975 (N_5975,N_2106,N_628);
and U5976 (N_5976,N_1332,N_311);
or U5977 (N_5977,N_1903,N_1388);
and U5978 (N_5978,N_1977,N_1967);
nand U5979 (N_5979,N_2245,N_1663);
and U5980 (N_5980,N_2216,N_1714);
or U5981 (N_5981,N_2448,N_2098);
nor U5982 (N_5982,N_152,N_1354);
or U5983 (N_5983,N_804,N_1351);
xnor U5984 (N_5984,N_2065,N_1189);
nor U5985 (N_5985,N_48,N_1471);
or U5986 (N_5986,N_1611,N_1118);
xor U5987 (N_5987,N_84,N_2893);
and U5988 (N_5988,N_2976,N_295);
and U5989 (N_5989,N_516,N_1224);
or U5990 (N_5990,N_297,N_1732);
and U5991 (N_5991,N_2479,N_1208);
and U5992 (N_5992,N_1914,N_1234);
nand U5993 (N_5993,N_1080,N_2263);
nor U5994 (N_5994,N_2129,N_1690);
nor U5995 (N_5995,N_2582,N_1307);
nor U5996 (N_5996,N_1658,N_1224);
xnor U5997 (N_5997,N_524,N_603);
or U5998 (N_5998,N_454,N_2942);
nand U5999 (N_5999,N_268,N_2283);
xnor U6000 (N_6000,N_5201,N_5368);
or U6001 (N_6001,N_3849,N_4530);
and U6002 (N_6002,N_3758,N_5782);
nor U6003 (N_6003,N_5329,N_4739);
and U6004 (N_6004,N_3401,N_3426);
and U6005 (N_6005,N_4776,N_3938);
nor U6006 (N_6006,N_4856,N_3738);
and U6007 (N_6007,N_4577,N_4235);
or U6008 (N_6008,N_4278,N_4765);
nor U6009 (N_6009,N_4712,N_5557);
nand U6010 (N_6010,N_3271,N_3334);
xor U6011 (N_6011,N_4689,N_5966);
xnor U6012 (N_6012,N_4506,N_4870);
xor U6013 (N_6013,N_5730,N_5976);
and U6014 (N_6014,N_4289,N_3070);
and U6015 (N_6015,N_3330,N_3836);
or U6016 (N_6016,N_3056,N_3850);
xnor U6017 (N_6017,N_3593,N_3711);
nand U6018 (N_6018,N_4077,N_5977);
and U6019 (N_6019,N_5099,N_3717);
or U6020 (N_6020,N_4324,N_3153);
nand U6021 (N_6021,N_4848,N_4967);
and U6022 (N_6022,N_5781,N_3398);
and U6023 (N_6023,N_3287,N_4238);
and U6024 (N_6024,N_5550,N_5942);
nand U6025 (N_6025,N_3897,N_5186);
or U6026 (N_6026,N_3822,N_3756);
xor U6027 (N_6027,N_3504,N_4194);
nand U6028 (N_6028,N_5635,N_4729);
xor U6029 (N_6029,N_3356,N_5842);
nor U6030 (N_6030,N_3073,N_3256);
xnor U6031 (N_6031,N_4040,N_3257);
or U6032 (N_6032,N_5930,N_4624);
nor U6033 (N_6033,N_3441,N_3116);
nor U6034 (N_6034,N_3828,N_3485);
and U6035 (N_6035,N_5658,N_5462);
xor U6036 (N_6036,N_5137,N_3808);
or U6037 (N_6037,N_5642,N_3408);
and U6038 (N_6038,N_5364,N_3164);
nor U6039 (N_6039,N_4604,N_5480);
and U6040 (N_6040,N_3264,N_4627);
and U6041 (N_6041,N_3418,N_3643);
xnor U6042 (N_6042,N_5307,N_3963);
or U6043 (N_6043,N_5523,N_4834);
nor U6044 (N_6044,N_3099,N_4212);
nand U6045 (N_6045,N_3678,N_4590);
nand U6046 (N_6046,N_3660,N_5379);
and U6047 (N_6047,N_3252,N_5048);
nor U6048 (N_6048,N_4178,N_5237);
nand U6049 (N_6049,N_4231,N_5469);
xnor U6050 (N_6050,N_3361,N_4626);
xnor U6051 (N_6051,N_3674,N_3102);
or U6052 (N_6052,N_3241,N_5773);
xor U6053 (N_6053,N_5770,N_3682);
xnor U6054 (N_6054,N_5270,N_4353);
xor U6055 (N_6055,N_4159,N_5793);
nand U6056 (N_6056,N_4386,N_3284);
nor U6057 (N_6057,N_5470,N_3618);
nand U6058 (N_6058,N_4520,N_5356);
nand U6059 (N_6059,N_5820,N_4602);
or U6060 (N_6060,N_5583,N_4912);
nand U6061 (N_6061,N_5290,N_3596);
nand U6062 (N_6062,N_5626,N_5592);
nand U6063 (N_6063,N_5315,N_3087);
and U6064 (N_6064,N_4163,N_3825);
nand U6065 (N_6065,N_4688,N_4217);
nor U6066 (N_6066,N_3658,N_3174);
nand U6067 (N_6067,N_3251,N_3795);
nor U6068 (N_6068,N_3857,N_5042);
or U6069 (N_6069,N_4575,N_5141);
xor U6070 (N_6070,N_4989,N_4828);
xnor U6071 (N_6071,N_3824,N_3886);
or U6072 (N_6072,N_4678,N_4871);
or U6073 (N_6073,N_5938,N_3097);
xor U6074 (N_6074,N_3629,N_4204);
and U6075 (N_6075,N_4378,N_3659);
xnor U6076 (N_6076,N_5325,N_4424);
and U6077 (N_6077,N_5674,N_4770);
and U6078 (N_6078,N_4334,N_3704);
and U6079 (N_6079,N_3422,N_5828);
and U6080 (N_6080,N_4079,N_5920);
nand U6081 (N_6081,N_3123,N_5323);
or U6082 (N_6082,N_4693,N_3166);
xnor U6083 (N_6083,N_5296,N_4019);
xor U6084 (N_6084,N_3156,N_3013);
xnor U6085 (N_6085,N_3992,N_5958);
xnor U6086 (N_6086,N_3407,N_4321);
nor U6087 (N_6087,N_5444,N_5016);
or U6088 (N_6088,N_4850,N_4682);
nand U6089 (N_6089,N_4705,N_3798);
nand U6090 (N_6090,N_5433,N_4941);
or U6091 (N_6091,N_3909,N_5413);
or U6092 (N_6092,N_3293,N_5490);
nor U6093 (N_6093,N_4366,N_3213);
nor U6094 (N_6094,N_4843,N_5401);
and U6095 (N_6095,N_3845,N_3957);
or U6096 (N_6096,N_4262,N_5381);
nand U6097 (N_6097,N_4412,N_3910);
nand U6098 (N_6098,N_3433,N_5407);
xor U6099 (N_6099,N_3809,N_4781);
and U6100 (N_6100,N_3332,N_4084);
nor U6101 (N_6101,N_5984,N_3238);
or U6102 (N_6102,N_3577,N_4860);
and U6103 (N_6103,N_3096,N_4697);
xnor U6104 (N_6104,N_4182,N_5590);
and U6105 (N_6105,N_4096,N_5617);
or U6106 (N_6106,N_3453,N_5351);
nor U6107 (N_6107,N_3242,N_5151);
or U6108 (N_6108,N_4890,N_5182);
xor U6109 (N_6109,N_4645,N_4883);
or U6110 (N_6110,N_4960,N_3805);
or U6111 (N_6111,N_3090,N_3871);
and U6112 (N_6112,N_4229,N_5352);
and U6113 (N_6113,N_5508,N_3765);
nand U6114 (N_6114,N_3145,N_3172);
or U6115 (N_6115,N_4582,N_4001);
or U6116 (N_6116,N_5265,N_3377);
or U6117 (N_6117,N_3313,N_4186);
xor U6118 (N_6118,N_5372,N_5481);
and U6119 (N_6119,N_3892,N_4901);
and U6120 (N_6120,N_4949,N_3564);
nand U6121 (N_6121,N_3576,N_3616);
and U6122 (N_6122,N_3733,N_4181);
and U6123 (N_6123,N_4296,N_4075);
nor U6124 (N_6124,N_5403,N_3894);
nand U6125 (N_6125,N_5675,N_4025);
nand U6126 (N_6126,N_4862,N_4662);
and U6127 (N_6127,N_4256,N_5205);
nand U6128 (N_6128,N_3322,N_4793);
nand U6129 (N_6129,N_4674,N_5108);
nor U6130 (N_6130,N_3788,N_3709);
xnor U6131 (N_6131,N_3880,N_3180);
and U6132 (N_6132,N_5327,N_5259);
nor U6133 (N_6133,N_3051,N_5349);
nand U6134 (N_6134,N_5094,N_3866);
and U6135 (N_6135,N_3868,N_4690);
nor U6136 (N_6136,N_5535,N_3112);
and U6137 (N_6137,N_5267,N_3980);
xor U6138 (N_6138,N_3011,N_3445);
and U6139 (N_6139,N_3667,N_5247);
or U6140 (N_6140,N_3403,N_5563);
nand U6141 (N_6141,N_4006,N_5233);
nor U6142 (N_6142,N_4291,N_4320);
and U6143 (N_6143,N_5025,N_3675);
and U6144 (N_6144,N_5892,N_4101);
xnor U6145 (N_6145,N_4701,N_4885);
nor U6146 (N_6146,N_3951,N_3666);
nor U6147 (N_6147,N_3904,N_3955);
xor U6148 (N_6148,N_5377,N_3695);
and U6149 (N_6149,N_4827,N_4655);
and U6150 (N_6150,N_5880,N_4005);
and U6151 (N_6151,N_3353,N_3608);
nand U6152 (N_6152,N_5740,N_3728);
xor U6153 (N_6153,N_3454,N_4823);
xnor U6154 (N_6154,N_4195,N_3231);
nand U6155 (N_6155,N_5593,N_5418);
xnor U6156 (N_6156,N_3571,N_5121);
nor U6157 (N_6157,N_5074,N_3829);
and U6158 (N_6158,N_5900,N_4027);
xor U6159 (N_6159,N_4640,N_5672);
nand U6160 (N_6160,N_4389,N_3954);
and U6161 (N_6161,N_4868,N_4493);
xnor U6162 (N_6162,N_3589,N_5609);
xor U6163 (N_6163,N_3160,N_4628);
or U6164 (N_6164,N_3442,N_4600);
and U6165 (N_6165,N_4302,N_5985);
nand U6166 (N_6166,N_5514,N_4936);
and U6167 (N_6167,N_3518,N_5556);
nand U6168 (N_6168,N_4149,N_4166);
xor U6169 (N_6169,N_5117,N_5622);
and U6170 (N_6170,N_5638,N_5402);
and U6171 (N_6171,N_5603,N_3583);
and U6172 (N_6172,N_5494,N_5560);
and U6173 (N_6173,N_4659,N_5571);
nand U6174 (N_6174,N_3797,N_4984);
nor U6175 (N_6175,N_4753,N_5037);
xor U6176 (N_6176,N_4292,N_3713);
nand U6177 (N_6177,N_3131,N_3902);
xor U6178 (N_6178,N_4847,N_3721);
nand U6179 (N_6179,N_4034,N_4191);
nand U6180 (N_6180,N_4436,N_4259);
or U6181 (N_6181,N_4432,N_3423);
nand U6182 (N_6182,N_5066,N_3137);
nor U6183 (N_6183,N_3872,N_4916);
and U6184 (N_6184,N_3295,N_3029);
or U6185 (N_6185,N_5471,N_3997);
nand U6186 (N_6186,N_4831,N_4316);
nor U6187 (N_6187,N_3889,N_4341);
and U6188 (N_6188,N_3705,N_5572);
and U6189 (N_6189,N_3911,N_4350);
and U6190 (N_6190,N_4309,N_5071);
nand U6191 (N_6191,N_3383,N_4650);
or U6192 (N_6192,N_4286,N_5055);
nand U6193 (N_6193,N_4709,N_4997);
and U6194 (N_6194,N_4018,N_5858);
nand U6195 (N_6195,N_4450,N_3919);
nor U6196 (N_6196,N_3336,N_4728);
nand U6197 (N_6197,N_3609,N_4932);
nand U6198 (N_6198,N_5673,N_4263);
xor U6199 (N_6199,N_3155,N_4784);
or U6200 (N_6200,N_5595,N_5095);
and U6201 (N_6201,N_5419,N_3098);
and U6202 (N_6202,N_3842,N_5623);
nand U6203 (N_6203,N_4087,N_5125);
and U6204 (N_6204,N_5335,N_5221);
and U6205 (N_6205,N_3806,N_5276);
and U6206 (N_6206,N_3091,N_5559);
xor U6207 (N_6207,N_3368,N_4507);
xnor U6208 (N_6208,N_5499,N_4447);
nand U6209 (N_6209,N_3104,N_3501);
and U6210 (N_6210,N_5657,N_4955);
and U6211 (N_6211,N_3050,N_4536);
nand U6212 (N_6212,N_5519,N_3509);
nand U6213 (N_6213,N_5359,N_5032);
or U6214 (N_6214,N_4009,N_5637);
nor U6215 (N_6215,N_4406,N_3127);
nor U6216 (N_6216,N_3223,N_5823);
and U6217 (N_6217,N_4511,N_3823);
and U6218 (N_6218,N_4400,N_4239);
nand U6219 (N_6219,N_5809,N_3025);
nor U6220 (N_6220,N_4060,N_5734);
nor U6221 (N_6221,N_4428,N_5131);
xor U6222 (N_6222,N_5751,N_4319);
xnor U6223 (N_6223,N_3010,N_4934);
and U6224 (N_6224,N_5870,N_5532);
and U6225 (N_6225,N_3597,N_5273);
and U6226 (N_6226,N_3663,N_4852);
nor U6227 (N_6227,N_4151,N_4171);
nand U6228 (N_6228,N_5033,N_3723);
nor U6229 (N_6229,N_4363,N_5780);
xnor U6230 (N_6230,N_5999,N_5453);
nand U6231 (N_6231,N_4008,N_3452);
nand U6232 (N_6232,N_4702,N_3740);
xor U6233 (N_6233,N_3005,N_5891);
or U6234 (N_6234,N_5811,N_3652);
xor U6235 (N_6235,N_4703,N_4517);
xnor U6236 (N_6236,N_5175,N_4260);
and U6237 (N_6237,N_5456,N_3323);
or U6238 (N_6238,N_3048,N_5241);
or U6239 (N_6239,N_3458,N_4268);
nor U6240 (N_6240,N_4724,N_3266);
xor U6241 (N_6241,N_5040,N_3744);
nor U6242 (N_6242,N_3425,N_5901);
and U6243 (N_6243,N_4158,N_3531);
or U6244 (N_6244,N_3272,N_4156);
xor U6245 (N_6245,N_5973,N_3890);
nor U6246 (N_6246,N_5946,N_3664);
nor U6247 (N_6247,N_4535,N_3060);
nand U6248 (N_6248,N_5846,N_3516);
nor U6249 (N_6249,N_4824,N_4494);
nor U6250 (N_6250,N_3631,N_4240);
nor U6251 (N_6251,N_5876,N_4359);
nor U6252 (N_6252,N_3141,N_5395);
and U6253 (N_6253,N_3676,N_5669);
xor U6254 (N_6254,N_4094,N_5929);
nor U6255 (N_6255,N_5813,N_3354);
nor U6256 (N_6256,N_4617,N_3170);
nand U6257 (N_6257,N_3369,N_5990);
nor U6258 (N_6258,N_4462,N_5786);
nand U6259 (N_6259,N_5597,N_5361);
or U6260 (N_6260,N_3128,N_3157);
or U6261 (N_6261,N_3668,N_5173);
and U6262 (N_6262,N_3562,N_4095);
nor U6263 (N_6263,N_3396,N_3497);
and U6264 (N_6264,N_4656,N_3639);
nand U6265 (N_6265,N_3685,N_3249);
and U6266 (N_6266,N_5878,N_3535);
xnor U6267 (N_6267,N_5646,N_4717);
nand U6268 (N_6268,N_5145,N_4346);
nand U6269 (N_6269,N_5331,N_3967);
nand U6270 (N_6270,N_5206,N_5458);
and U6271 (N_6271,N_3748,N_3197);
and U6272 (N_6272,N_5152,N_3047);
nand U6273 (N_6273,N_5388,N_5399);
nor U6274 (N_6274,N_5124,N_5601);
or U6275 (N_6275,N_4754,N_5378);
xor U6276 (N_6276,N_4057,N_4921);
xnor U6277 (N_6277,N_4192,N_3747);
and U6278 (N_6278,N_5189,N_3015);
nor U6279 (N_6279,N_5231,N_3340);
xor U6280 (N_6280,N_5286,N_3762);
xnor U6281 (N_6281,N_3324,N_3832);
or U6282 (N_6282,N_5266,N_3302);
xnor U6283 (N_6283,N_3397,N_5000);
or U6284 (N_6284,N_4414,N_5907);
xnor U6285 (N_6285,N_4528,N_5533);
nor U6286 (N_6286,N_4541,N_3224);
xor U6287 (N_6287,N_4418,N_3261);
or U6288 (N_6288,N_4100,N_4763);
xor U6289 (N_6289,N_4877,N_4193);
xor U6290 (N_6290,N_3977,N_3636);
or U6291 (N_6291,N_5087,N_4318);
nor U6292 (N_6292,N_5474,N_4415);
and U6293 (N_6293,N_5539,N_3972);
or U6294 (N_6294,N_5621,N_5695);
or U6295 (N_6295,N_4083,N_5452);
nand U6296 (N_6296,N_5169,N_4694);
nor U6297 (N_6297,N_4722,N_4913);
and U6298 (N_6298,N_5184,N_3546);
and U6299 (N_6299,N_4063,N_4143);
xor U6300 (N_6300,N_5949,N_5840);
and U6301 (N_6301,N_4388,N_3820);
and U6302 (N_6302,N_4906,N_3474);
or U6303 (N_6303,N_3212,N_4796);
nor U6304 (N_6304,N_3804,N_3205);
nor U6305 (N_6305,N_3653,N_3814);
xnor U6306 (N_6306,N_4559,N_3218);
nor U6307 (N_6307,N_3477,N_3862);
or U6308 (N_6308,N_4145,N_3530);
nand U6309 (N_6309,N_4219,N_3149);
nand U6310 (N_6310,N_3885,N_4305);
nor U6311 (N_6311,N_4023,N_3979);
and U6312 (N_6312,N_5822,N_3464);
or U6313 (N_6313,N_4814,N_3973);
nand U6314 (N_6314,N_5439,N_3863);
or U6315 (N_6315,N_4080,N_3706);
or U6316 (N_6316,N_3027,N_4691);
or U6317 (N_6317,N_5218,N_4139);
xor U6318 (N_6318,N_5142,N_3560);
or U6319 (N_6319,N_5150,N_3045);
and U6320 (N_6320,N_3306,N_3110);
and U6321 (N_6321,N_3565,N_5304);
xnor U6322 (N_6322,N_3514,N_5225);
xnor U6323 (N_6323,N_4924,N_4172);
nand U6324 (N_6324,N_5251,N_5553);
nor U6325 (N_6325,N_5165,N_4330);
nand U6326 (N_6326,N_5376,N_4859);
nand U6327 (N_6327,N_5525,N_3626);
xor U6328 (N_6328,N_5357,N_5854);
nand U6329 (N_6329,N_5187,N_4958);
nand U6330 (N_6330,N_5511,N_3049);
or U6331 (N_6331,N_4433,N_3881);
nand U6332 (N_6332,N_3720,N_5214);
xor U6333 (N_6333,N_5503,N_5855);
nand U6334 (N_6334,N_4761,N_4512);
xor U6335 (N_6335,N_5687,N_3018);
or U6336 (N_6336,N_3736,N_5197);
xor U6337 (N_6337,N_5172,N_5252);
nand U6338 (N_6338,N_4177,N_5831);
xor U6339 (N_6339,N_5319,N_5422);
or U6340 (N_6340,N_4573,N_3982);
xnor U6341 (N_6341,N_5634,N_4222);
and U6342 (N_6342,N_4521,N_4634);
or U6343 (N_6343,N_3351,N_3040);
and U6344 (N_6344,N_3864,N_4199);
nand U6345 (N_6345,N_4891,N_3095);
and U6346 (N_6346,N_4534,N_5035);
nor U6347 (N_6347,N_4503,N_4938);
and U6348 (N_6348,N_4283,N_3752);
nor U6349 (N_6349,N_3461,N_3041);
xnor U6350 (N_6350,N_4068,N_5633);
xnor U6351 (N_6351,N_5008,N_4708);
and U6352 (N_6352,N_3895,N_4725);
or U6353 (N_6353,N_5488,N_5879);
nor U6354 (N_6354,N_5434,N_3154);
or U6355 (N_6355,N_3489,N_3337);
xor U6356 (N_6356,N_4742,N_3528);
xnor U6357 (N_6357,N_4348,N_5698);
xnor U6358 (N_6358,N_4976,N_4269);
and U6359 (N_6359,N_5158,N_3525);
xnor U6360 (N_6360,N_4853,N_4576);
xnor U6361 (N_6361,N_3960,N_5765);
xor U6362 (N_6362,N_5028,N_3800);
xnor U6363 (N_6363,N_5261,N_4397);
nand U6364 (N_6364,N_4558,N_3932);
nor U6365 (N_6365,N_5791,N_3770);
xnor U6366 (N_6366,N_4052,N_5925);
and U6367 (N_6367,N_3480,N_3558);
nor U6368 (N_6368,N_3939,N_5805);
or U6369 (N_6369,N_5190,N_4411);
nor U6370 (N_6370,N_3083,N_5204);
nor U6371 (N_6371,N_5199,N_4134);
or U6372 (N_6372,N_3874,N_5179);
nand U6373 (N_6373,N_4875,N_5077);
or U6374 (N_6374,N_5504,N_4735);
and U6375 (N_6375,N_3655,N_4601);
or U6376 (N_6376,N_4127,N_5056);
xor U6377 (N_6377,N_3750,N_5619);
xnor U6378 (N_6378,N_4533,N_4349);
and U6379 (N_6379,N_4161,N_4215);
nand U6380 (N_6380,N_3312,N_4463);
nand U6381 (N_6381,N_4306,N_4692);
and U6382 (N_6382,N_3066,N_5957);
and U6383 (N_6383,N_5089,N_4592);
and U6384 (N_6384,N_4266,N_3139);
nand U6385 (N_6385,N_4902,N_3054);
or U6386 (N_6386,N_5829,N_4148);
nor U6387 (N_6387,N_4311,N_4756);
and U6388 (N_6388,N_5893,N_4646);
and U6389 (N_6389,N_4322,N_4097);
nor U6390 (N_6390,N_5706,N_4846);
nor U6391 (N_6391,N_5409,N_5856);
nand U6392 (N_6392,N_3647,N_5546);
nand U6393 (N_6393,N_3082,N_5555);
nand U6394 (N_6394,N_3986,N_4223);
or U6395 (N_6395,N_4774,N_5371);
nand U6396 (N_6396,N_4965,N_3782);
or U6397 (N_6397,N_4899,N_5826);
and U6398 (N_6398,N_4497,N_5144);
nor U6399 (N_6399,N_4197,N_3778);
xnor U6400 (N_6400,N_4041,N_4442);
nor U6401 (N_6401,N_3755,N_3232);
nand U6402 (N_6402,N_3852,N_3585);
and U6403 (N_6403,N_3896,N_3724);
nand U6404 (N_6404,N_4581,N_3783);
xor U6405 (N_6405,N_5006,N_3215);
and U6406 (N_6406,N_3785,N_3633);
nand U6407 (N_6407,N_4935,N_4126);
and U6408 (N_6408,N_5374,N_4082);
xor U6409 (N_6409,N_5353,N_3768);
or U6410 (N_6410,N_3055,N_4813);
nand U6411 (N_6411,N_3429,N_5430);
and U6412 (N_6412,N_4970,N_5202);
nand U6413 (N_6413,N_4225,N_5005);
nor U6414 (N_6414,N_4547,N_3309);
and U6415 (N_6415,N_4849,N_5291);
nor U6416 (N_6416,N_3440,N_3754);
xor U6417 (N_6417,N_3233,N_5804);
nand U6418 (N_6418,N_5808,N_3230);
and U6419 (N_6419,N_3134,N_4994);
nand U6420 (N_6420,N_4252,N_5998);
nor U6421 (N_6421,N_4802,N_3247);
and U6422 (N_6422,N_3665,N_4762);
and U6423 (N_6423,N_3561,N_3072);
xnor U6424 (N_6424,N_4567,N_3532);
xnor U6425 (N_6425,N_3642,N_4308);
nor U6426 (N_6426,N_5872,N_4183);
nand U6427 (N_6427,N_3776,N_3473);
nor U6428 (N_6428,N_3927,N_5531);
nand U6429 (N_6429,N_4526,N_4404);
nand U6430 (N_6430,N_3572,N_3162);
nand U6431 (N_6431,N_3923,N_5548);
nand U6432 (N_6432,N_3206,N_4471);
and U6433 (N_6433,N_5904,N_4937);
and U6434 (N_6434,N_3446,N_3657);
xnor U6435 (N_6435,N_5026,N_4336);
and U6436 (N_6436,N_5497,N_4830);
xnor U6437 (N_6437,N_4816,N_3448);
and U6438 (N_6438,N_4298,N_5885);
nor U6439 (N_6439,N_4971,N_5061);
xor U6440 (N_6440,N_4498,N_5567);
nand U6441 (N_6441,N_3515,N_3221);
nand U6442 (N_6442,N_5764,N_3742);
nand U6443 (N_6443,N_5358,N_4981);
nor U6444 (N_6444,N_3059,N_4553);
or U6445 (N_6445,N_5824,N_5088);
xnor U6446 (N_6446,N_4538,N_3848);
nor U6447 (N_6447,N_5956,N_4954);
or U6448 (N_6448,N_4811,N_3316);
nand U6449 (N_6449,N_5079,N_3305);
nand U6450 (N_6450,N_4189,N_4539);
or U6451 (N_6451,N_5369,N_4554);
and U6452 (N_6452,N_3615,N_5836);
nand U6453 (N_6453,N_3502,N_5380);
and U6454 (N_6454,N_3985,N_4365);
nand U6455 (N_6455,N_4382,N_5735);
and U6456 (N_6456,N_5106,N_3690);
xor U6457 (N_6457,N_4504,N_5180);
and U6458 (N_6458,N_4568,N_4555);
or U6459 (N_6459,N_3840,N_3283);
nand U6460 (N_6460,N_4755,N_4927);
nor U6461 (N_6461,N_5253,N_3181);
or U6462 (N_6462,N_3638,N_5807);
nand U6463 (N_6463,N_4778,N_5941);
nand U6464 (N_6464,N_4757,N_5848);
nand U6465 (N_6465,N_5708,N_3837);
nand U6466 (N_6466,N_4460,N_3961);
nor U6467 (N_6467,N_4372,N_3611);
nor U6468 (N_6468,N_3931,N_5721);
or U6469 (N_6469,N_4825,N_4453);
nand U6470 (N_6470,N_5103,N_5921);
nor U6471 (N_6471,N_3944,N_3017);
or U6472 (N_6472,N_5166,N_5924);
xor U6473 (N_6473,N_5862,N_5060);
nor U6474 (N_6474,N_4940,N_5321);
xor U6475 (N_6475,N_5109,N_3523);
nand U6476 (N_6476,N_5160,N_5212);
xnor U6477 (N_6477,N_3402,N_3285);
and U6478 (N_6478,N_3465,N_5171);
nand U6479 (N_6479,N_4983,N_5043);
and U6480 (N_6480,N_5012,N_4900);
nor U6481 (N_6481,N_5193,N_5932);
xnor U6482 (N_6482,N_4276,N_4030);
or U6483 (N_6483,N_3375,N_3879);
or U6484 (N_6484,N_4394,N_5581);
nor U6485 (N_6485,N_5072,N_3012);
nand U6486 (N_6486,N_5161,N_4345);
and U6487 (N_6487,N_5234,N_3118);
nand U6488 (N_6488,N_5230,N_3595);
xnor U6489 (N_6489,N_4099,N_5700);
or U6490 (N_6490,N_4584,N_4956);
and U6491 (N_6491,N_3603,N_3699);
nand U6492 (N_6492,N_4812,N_4255);
nand U6493 (N_6493,N_5814,N_5502);
nand U6494 (N_6494,N_3812,N_4572);
or U6495 (N_6495,N_3042,N_5526);
and U6496 (N_6496,N_3411,N_4468);
nor U6497 (N_6497,N_5711,N_5159);
nor U6498 (N_6498,N_5527,N_5250);
xor U6499 (N_6499,N_3703,N_5310);
nor U6500 (N_6500,N_3201,N_4751);
nand U6501 (N_6501,N_4977,N_5945);
xor U6502 (N_6502,N_5799,N_3486);
nor U6503 (N_6503,N_5627,N_4310);
or U6504 (N_6504,N_5011,N_3681);
nand U6505 (N_6505,N_5997,N_4947);
nand U6506 (N_6506,N_4144,N_3567);
or U6507 (N_6507,N_4661,N_4141);
nor U6508 (N_6508,N_4797,N_5479);
and U6509 (N_6509,N_5537,N_3563);
and U6510 (N_6510,N_5864,N_3592);
or U6511 (N_6511,N_4107,N_5739);
or U6512 (N_6512,N_4704,N_3943);
xor U6513 (N_6513,N_3254,N_5303);
xor U6514 (N_6514,N_4695,N_4951);
or U6515 (N_6515,N_4364,N_3591);
xor U6516 (N_6516,N_3286,N_3000);
or U6517 (N_6517,N_5147,N_5002);
nor U6518 (N_6518,N_3409,N_5775);
and U6519 (N_6519,N_4764,N_5457);
nor U6520 (N_6520,N_5749,N_5887);
and U6521 (N_6521,N_3124,N_5701);
xor U6522 (N_6522,N_3543,N_3484);
or U6523 (N_6523,N_5080,N_3436);
nor U6524 (N_6524,N_3942,N_5522);
or U6525 (N_6525,N_4805,N_4419);
or U6526 (N_6526,N_5618,N_3359);
and U6527 (N_6527,N_4114,N_5936);
nand U6528 (N_6528,N_4633,N_3071);
nand U6529 (N_6529,N_4616,N_5530);
xor U6530 (N_6530,N_4031,N_5612);
and U6531 (N_6531,N_3976,N_5404);
nand U6532 (N_6532,N_5285,N_5606);
or U6533 (N_6533,N_5665,N_5348);
nand U6534 (N_6534,N_5615,N_5713);
xnor U6535 (N_6535,N_3136,N_5312);
nand U6536 (N_6536,N_5724,N_4745);
or U6537 (N_6537,N_5645,N_4485);
nand U6538 (N_6538,N_3046,N_3279);
or U6539 (N_6539,N_4896,N_4012);
xnor U6540 (N_6540,N_3918,N_4179);
nand U6541 (N_6541,N_3790,N_5138);
xnor U6542 (N_6542,N_4317,N_3651);
nor U6543 (N_6543,N_4719,N_4147);
and U6544 (N_6544,N_4758,N_5120);
nor U6545 (N_6545,N_4968,N_4799);
and U6546 (N_6546,N_4294,N_5365);
nand U6547 (N_6547,N_4518,N_5257);
xnor U6548 (N_6548,N_5975,N_5123);
nand U6549 (N_6549,N_3841,N_4187);
nand U6550 (N_6550,N_3873,N_5937);
nor U6551 (N_6551,N_4015,N_3771);
and U6552 (N_6552,N_4537,N_5447);
or U6553 (N_6553,N_4649,N_5918);
nand U6554 (N_6554,N_4780,N_5334);
nand U6555 (N_6555,N_5385,N_3069);
nand U6556 (N_6556,N_3103,N_5258);
nand U6557 (N_6557,N_3344,N_5988);
or U6558 (N_6558,N_4056,N_5865);
xnor U6559 (N_6559,N_4565,N_5487);
nor U6560 (N_6560,N_5569,N_3088);
xnor U6561 (N_6561,N_4879,N_4721);
xnor U6562 (N_6562,N_5305,N_3507);
or U6563 (N_6563,N_4782,N_5467);
nor U6564 (N_6564,N_5528,N_5599);
xnor U6565 (N_6565,N_5796,N_4595);
nand U6566 (N_6566,N_3512,N_4746);
or U6567 (N_6567,N_5586,N_3859);
and U6568 (N_6568,N_3079,N_4919);
and U6569 (N_6569,N_3001,N_5350);
or U6570 (N_6570,N_5678,N_5483);
and U6571 (N_6571,N_5425,N_4514);
and U6572 (N_6572,N_4714,N_5338);
nand U6573 (N_6573,N_5859,N_3521);
nor U6574 (N_6574,N_3301,N_3794);
or U6575 (N_6575,N_5373,N_3234);
or U6576 (N_6576,N_3019,N_4055);
and U6577 (N_6577,N_4438,N_5045);
nor U6578 (N_6578,N_4658,N_4486);
nor U6579 (N_6579,N_4446,N_5830);
xor U6580 (N_6580,N_3524,N_4284);
and U6581 (N_6581,N_4459,N_4233);
nand U6582 (N_6582,N_5978,N_5228);
nor U6583 (N_6583,N_5100,N_5164);
xor U6584 (N_6584,N_5493,N_5656);
nand U6585 (N_6585,N_4855,N_5170);
xor U6586 (N_6586,N_3151,N_4772);
xnor U6587 (N_6587,N_4332,N_5955);
xor U6588 (N_6588,N_4403,N_3555);
nand U6589 (N_6589,N_5648,N_4184);
and U6590 (N_6590,N_5630,N_3352);
and U6591 (N_6591,N_3255,N_4300);
or U6592 (N_6592,N_5344,N_4335);
nand U6593 (N_6593,N_5954,N_3672);
or U6594 (N_6594,N_5816,N_4495);
and U6595 (N_6595,N_3276,N_3260);
nand U6596 (N_6596,N_3304,N_5959);
nand U6597 (N_6597,N_5289,N_4798);
nand U6598 (N_6598,N_5475,N_3917);
xor U6599 (N_6599,N_3496,N_5916);
xnor U6600 (N_6600,N_4787,N_4016);
nor U6601 (N_6601,N_5647,N_4864);
nor U6602 (N_6602,N_4091,N_3211);
or U6603 (N_6603,N_3519,N_5613);
or U6604 (N_6604,N_3689,N_5354);
xor U6605 (N_6605,N_3529,N_3696);
nor U6606 (N_6606,N_3999,N_3715);
nor U6607 (N_6607,N_5162,N_5992);
nor U6608 (N_6608,N_3606,N_4808);
or U6609 (N_6609,N_4218,N_3198);
xor U6610 (N_6610,N_4273,N_4637);
nor U6611 (N_6611,N_5083,N_5969);
or U6612 (N_6612,N_4065,N_4651);
xor U6613 (N_6613,N_5501,N_4054);
and U6614 (N_6614,N_4371,N_3908);
and U6615 (N_6615,N_5262,N_4153);
nand U6616 (N_6616,N_3163,N_3273);
and U6617 (N_6617,N_5101,N_4216);
xnor U6618 (N_6618,N_5833,N_4806);
or U6619 (N_6619,N_4845,N_5758);
or U6620 (N_6620,N_4944,N_5460);
xor U6621 (N_6621,N_5543,N_4783);
and U6622 (N_6622,N_4061,N_4380);
nor U6623 (N_6623,N_4759,N_5363);
xor U6624 (N_6624,N_3143,N_3719);
or U6625 (N_6625,N_5549,N_3004);
and U6626 (N_6626,N_4683,N_3975);
nand U6627 (N_6627,N_5745,N_4070);
or U6628 (N_6628,N_5336,N_3679);
and U6629 (N_6629,N_5133,N_4480);
or U6630 (N_6630,N_5911,N_3434);
or U6631 (N_6631,N_5260,N_5464);
nand U6632 (N_6632,N_3907,N_4654);
nor U6633 (N_6633,N_4801,N_3122);
or U6634 (N_6634,N_4821,N_5018);
or U6635 (N_6635,N_5069,N_5326);
or U6636 (N_6636,N_3246,N_4039);
xnor U6637 (N_6637,N_5662,N_4051);
and U6638 (N_6638,N_4174,N_5943);
xor U6639 (N_6639,N_4355,N_3760);
nand U6640 (N_6640,N_3331,N_5020);
xnor U6641 (N_6641,N_4632,N_5991);
and U6642 (N_6642,N_4264,N_3030);
nand U6643 (N_6643,N_5308,N_5424);
xnor U6644 (N_6644,N_4086,N_4873);
xor U6645 (N_6645,N_3648,N_3635);
and U6646 (N_6646,N_5970,N_3376);
or U6647 (N_6647,N_4726,N_4237);
xnor U6648 (N_6648,N_4465,N_5140);
nand U6649 (N_6649,N_4379,N_5951);
nor U6650 (N_6650,N_4930,N_5010);
nor U6651 (N_6651,N_3725,N_5436);
or U6652 (N_6652,N_4049,N_3311);
nor U6653 (N_6653,N_4053,N_5227);
or U6654 (N_6654,N_5757,N_5747);
and U6655 (N_6655,N_3333,N_5316);
and U6656 (N_6656,N_5236,N_4591);
nand U6657 (N_6657,N_5743,N_3843);
xnor U6658 (N_6658,N_3065,N_4164);
and U6659 (N_6659,N_3637,N_4525);
nand U6660 (N_6660,N_4790,N_3691);
xor U6661 (N_6661,N_3887,N_5640);
nor U6662 (N_6662,N_4437,N_4128);
xor U6663 (N_6663,N_3940,N_3420);
or U6664 (N_6664,N_3810,N_3544);
or U6665 (N_6665,N_5426,N_4088);
or U6666 (N_6666,N_4933,N_5428);
nand U6667 (N_6667,N_4020,N_4509);
and U6668 (N_6668,N_5707,N_4399);
nor U6669 (N_6669,N_4925,N_4072);
nand U6670 (N_6670,N_5223,N_3856);
nor U6671 (N_6671,N_5558,N_3475);
nor U6672 (N_6672,N_5492,N_4354);
nor U6673 (N_6673,N_5347,N_3210);
or U6674 (N_6674,N_5671,N_5947);
xor U6675 (N_6675,N_5961,N_4232);
nand U6676 (N_6676,N_3580,N_5768);
nor U6677 (N_6677,N_3965,N_5741);
and U6678 (N_6678,N_4653,N_5752);
nand U6679 (N_6679,N_5269,N_5681);
nand U6680 (N_6680,N_3192,N_5355);
and U6681 (N_6681,N_4749,N_4234);
xnor U6682 (N_6682,N_5476,N_4398);
or U6683 (N_6683,N_5896,N_3138);
nor U6684 (N_6684,N_5986,N_4892);
and U6685 (N_6685,N_5134,N_3861);
and U6686 (N_6686,N_5054,N_3108);
and U6687 (N_6687,N_4113,N_3101);
nand U6688 (N_6688,N_5067,N_4777);
nor U6689 (N_6689,N_5632,N_5210);
nand U6690 (N_6690,N_5342,N_4048);
xnor U6691 (N_6691,N_3500,N_4730);
or U6692 (N_6692,N_3751,N_4106);
xor U6693 (N_6693,N_5867,N_5001);
nor U6694 (N_6694,N_3237,N_5753);
xor U6695 (N_6695,N_5096,N_4250);
nand U6696 (N_6696,N_3844,N_4878);
xor U6697 (N_6697,N_4304,N_3554);
nand U6698 (N_6698,N_5435,N_3036);
or U6699 (N_6699,N_5676,N_3094);
nand U6700 (N_6700,N_5438,N_5287);
or U6701 (N_6701,N_4123,N_5341);
nor U6702 (N_6702,N_3729,N_4928);
xor U6703 (N_6703,N_4093,N_4502);
xnor U6704 (N_6704,N_3245,N_4562);
or U6705 (N_6705,N_3834,N_5311);
nor U6706 (N_6706,N_4895,N_3338);
nand U6707 (N_6707,N_4996,N_5073);
nand U6708 (N_6708,N_3450,N_4548);
or U6709 (N_6709,N_4923,N_5301);
and U6710 (N_6710,N_3202,N_3632);
nand U6711 (N_6711,N_3363,N_5825);
xnor U6712 (N_6712,N_5176,N_4407);
nor U6713 (N_6713,N_4458,N_4917);
nand U6714 (N_6714,N_3610,N_4190);
nor U6715 (N_6715,N_4168,N_3387);
nand U6716 (N_6716,N_5652,N_4285);
or U6717 (N_6717,N_4328,N_5472);
nand U6718 (N_6718,N_3912,N_4211);
and U6719 (N_6719,N_4914,N_3614);
nand U6720 (N_6720,N_4085,N_4668);
nand U6721 (N_6721,N_4142,N_4718);
nor U6722 (N_6722,N_3380,N_4867);
nand U6723 (N_6723,N_4657,N_5697);
xor U6724 (N_6724,N_3292,N_4026);
nand U6725 (N_6725,N_4157,N_3296);
nand U6726 (N_6726,N_5093,N_3265);
or U6727 (N_6727,N_5877,N_5579);
nor U6728 (N_6728,N_3732,N_4244);
nor U6729 (N_6729,N_4915,N_4208);
and U6730 (N_6730,N_3214,N_3437);
nand U6731 (N_6731,N_3288,N_3817);
nand U6732 (N_6732,N_5841,N_4138);
and U6733 (N_6733,N_4140,N_5512);
and U6734 (N_6734,N_3169,N_4478);
and U6735 (N_6735,N_5256,N_5463);
nand U6736 (N_6736,N_4000,N_3188);
xnor U6737 (N_6737,N_3971,N_4076);
or U6738 (N_6738,N_3731,N_5847);
nand U6739 (N_6739,N_5897,N_4844);
nand U6740 (N_6740,N_4564,N_3893);
and U6741 (N_6741,N_5737,N_3325);
nor U6742 (N_6742,N_3601,N_5155);
or U6743 (N_6743,N_5726,N_5415);
and U6744 (N_6744,N_5570,N_5653);
and U6745 (N_6745,N_4227,N_5518);
or U6746 (N_6746,N_5248,N_3662);
nand U6747 (N_6747,N_5772,N_5769);
xor U6748 (N_6748,N_3677,N_4952);
nor U6749 (N_6749,N_3661,N_5299);
nor U6750 (N_6750,N_5677,N_5370);
xor U6751 (N_6751,N_4837,N_3877);
and U6752 (N_6752,N_3796,N_4282);
nor U6753 (N_6753,N_3372,N_3207);
nand U6754 (N_6754,N_5748,N_3195);
and U6755 (N_6755,N_5015,N_4771);
nor U6756 (N_6756,N_4420,N_5114);
nor U6757 (N_6757,N_3135,N_5317);
nor U6758 (N_6758,N_5964,N_5944);
or U6759 (N_6759,N_4618,N_3968);
nand U6760 (N_6760,N_5397,N_5084);
and U6761 (N_6761,N_3701,N_4287);
nor U6762 (N_6762,N_4496,N_5884);
and U6763 (N_6763,N_3913,N_4425);
and U6764 (N_6764,N_3505,N_5030);
and U6765 (N_6765,N_4280,N_4299);
nand U6766 (N_6766,N_4448,N_4773);
and U6767 (N_6767,N_5027,N_4492);
nand U6768 (N_6768,N_4549,N_3443);
xor U6769 (N_6769,N_3217,N_4779);
xnor U6770 (N_6770,N_3327,N_3415);
nand U6771 (N_6771,N_3184,N_4550);
and U6772 (N_6772,N_5952,N_4327);
or U6773 (N_6773,N_3759,N_4430);
nand U6774 (N_6774,N_3686,N_3328);
nor U6775 (N_6775,N_5722,N_4467);
nand U6776 (N_6776,N_3899,N_5869);
nor U6777 (N_6777,N_5053,N_5489);
nor U6778 (N_6778,N_5890,N_3935);
and U6779 (N_6779,N_3793,N_4551);
or U6780 (N_6780,N_4307,N_5607);
and U6781 (N_6781,N_3964,N_5423);
or U6782 (N_6782,N_5702,N_3761);
nor U6783 (N_6783,N_3022,N_4047);
nand U6784 (N_6784,N_4011,N_3044);
nand U6785 (N_6785,N_3321,N_5245);
or U6786 (N_6786,N_4456,N_5314);
xnor U6787 (N_6787,N_3307,N_4290);
and U6788 (N_6788,N_5478,N_5953);
xor U6789 (N_6789,N_3621,N_5294);
and U6790 (N_6790,N_3870,N_5448);
or U6791 (N_6791,N_5860,N_4439);
nand U6792 (N_6792,N_4422,N_5521);
and U6793 (N_6793,N_5575,N_4043);
xor U6794 (N_6794,N_3952,N_5064);
nand U6795 (N_6795,N_4402,N_3370);
xor U6796 (N_6796,N_4421,N_4619);
nor U6797 (N_6797,N_3707,N_3062);
nor U6798 (N_6798,N_3710,N_4625);
and U6799 (N_6799,N_3428,N_5693);
and U6800 (N_6800,N_4687,N_5573);
xor U6801 (N_6801,N_3427,N_4715);
and U6802 (N_6802,N_3479,N_3444);
and U6803 (N_6803,N_3491,N_4441);
or U6804 (N_6804,N_4271,N_3349);
and U6805 (N_6805,N_4881,N_3120);
and U6806 (N_6806,N_5554,N_5905);
and U6807 (N_6807,N_3538,N_5441);
nor U6808 (N_6808,N_3339,N_3469);
and U6809 (N_6809,N_4314,N_3430);
and U6810 (N_6810,N_3688,N_3244);
nand U6811 (N_6811,N_5861,N_5624);
or U6812 (N_6812,N_5429,N_4401);
xnor U6813 (N_6813,N_3791,N_4137);
and U6814 (N_6814,N_5198,N_5933);
xor U6815 (N_6815,N_3787,N_4369);
xnor U6816 (N_6816,N_3673,N_3739);
xor U6817 (N_6817,N_5818,N_4652);
or U6818 (N_6818,N_3953,N_5128);
or U6819 (N_6819,N_5629,N_4133);
nor U6820 (N_6820,N_3277,N_5696);
or U6821 (N_6821,N_4243,N_4929);
nor U6822 (N_6822,N_5908,N_5987);
xnor U6823 (N_6823,N_5788,N_4540);
nand U6824 (N_6824,N_4205,N_3357);
xor U6825 (N_6825,N_4556,N_3061);
nand U6826 (N_6826,N_5995,N_4667);
and U6827 (N_6827,N_3694,N_3227);
or U6828 (N_6828,N_4586,N_3291);
and U6829 (N_6829,N_3412,N_4836);
nor U6830 (N_6830,N_4876,N_3299);
and U6831 (N_6831,N_4752,N_3925);
or U6832 (N_6832,N_5126,N_4443);
nor U6833 (N_6833,N_5174,N_4810);
and U6834 (N_6834,N_3941,N_3107);
or U6835 (N_6835,N_5139,N_3057);
and U6836 (N_6836,N_4959,N_4961);
xor U6837 (N_6837,N_4874,N_5242);
or U6838 (N_6838,N_5534,N_5200);
xor U6839 (N_6839,N_5491,N_5972);
nor U6840 (N_6840,N_4111,N_5738);
nor U6841 (N_6841,N_5473,N_3494);
xnor U6842 (N_6842,N_4033,N_5582);
xor U6843 (N_6843,N_5496,N_3204);
nor U6844 (N_6844,N_5545,N_4800);
or U6845 (N_6845,N_3757,N_5105);
xor U6846 (N_6846,N_5744,N_4647);
nor U6847 (N_6847,N_4566,N_4988);
nor U6848 (N_6848,N_5345,N_4112);
and U6849 (N_6849,N_3105,N_4405);
xor U6850 (N_6850,N_3650,N_5520);
and U6851 (N_6851,N_3399,N_5853);
nor U6852 (N_6852,N_4426,N_3270);
nand U6853 (N_6853,N_3080,N_4457);
and U6854 (N_6854,N_3488,N_3605);
and U6855 (N_6855,N_3506,N_3594);
nor U6856 (N_6856,N_4338,N_4681);
xnor U6857 (N_6857,N_3125,N_4098);
and U6858 (N_6858,N_4720,N_5213);
nor U6859 (N_6859,N_4807,N_4775);
nand U6860 (N_6860,N_4315,N_5948);
xor U6861 (N_6861,N_4669,N_4630);
nand U6862 (N_6862,N_3559,N_4804);
nor U6863 (N_6863,N_4666,N_3462);
or U6864 (N_6864,N_3826,N_5742);
and U6865 (N_6865,N_3730,N_5812);
nor U6866 (N_6866,N_4435,N_3298);
nand U6867 (N_6867,N_5416,N_4684);
and U6868 (N_6868,N_4991,N_5517);
or U6869 (N_6869,N_4545,N_4170);
or U6870 (N_6870,N_3216,N_3294);
or U6871 (N_6871,N_4670,N_4854);
or U6872 (N_6872,N_5119,N_4375);
or U6873 (N_6873,N_4440,N_4036);
xor U6874 (N_6874,N_5297,N_5584);
nor U6875 (N_6875,N_5927,N_5052);
nor U6876 (N_6876,N_3463,N_3996);
or U6877 (N_6877,N_5714,N_4066);
nand U6878 (N_6878,N_3540,N_3187);
nand U6879 (N_6879,N_5580,N_5313);
or U6880 (N_6880,N_5092,N_5023);
or U6881 (N_6881,N_5974,N_3994);
and U6882 (N_6882,N_5746,N_5309);
and U6883 (N_6883,N_5787,N_5217);
and U6884 (N_6884,N_5219,N_3741);
nor U6885 (N_6885,N_5293,N_5411);
nand U6886 (N_6886,N_5111,N_5224);
or U6887 (N_6887,N_4152,N_4351);
nor U6888 (N_6888,N_5340,N_4990);
and U6889 (N_6889,N_3974,N_4905);
or U6890 (N_6890,N_5017,N_5188);
nand U6891 (N_6891,N_5505,N_5038);
or U6892 (N_6892,N_4636,N_3106);
and U6893 (N_6893,N_3622,N_5292);
xnor U6894 (N_6894,N_5229,N_5249);
and U6895 (N_6895,N_5211,N_3343);
nor U6896 (N_6896,N_5153,N_4362);
and U6897 (N_6897,N_3847,N_5903);
and U6898 (N_6898,N_5587,N_4588);
and U6899 (N_6899,N_5465,N_4482);
xnor U6900 (N_6900,N_5789,N_5792);
nor U6901 (N_6901,N_3727,N_4609);
or U6902 (N_6902,N_4155,N_5794);
xnor U6903 (N_6903,N_3310,N_4185);
nor U6904 (N_6904,N_3391,N_5614);
nand U6905 (N_6905,N_3743,N_3278);
and U6906 (N_6906,N_4081,N_3031);
and U6907 (N_6907,N_3683,N_5412);
nand U6908 (N_6908,N_4476,N_3590);
and U6909 (N_6909,N_5041,N_3009);
nor U6910 (N_6910,N_3389,N_5122);
or U6911 (N_6911,N_3394,N_3393);
nand U6912 (N_6912,N_3350,N_4973);
xnor U6913 (N_6913,N_3625,N_3226);
xnor U6914 (N_6914,N_3858,N_5222);
xnor U6915 (N_6915,N_4331,N_5149);
nand U6916 (N_6916,N_4251,N_3460);
and U6917 (N_6917,N_5075,N_3499);
nor U6918 (N_6918,N_5923,N_5300);
nor U6919 (N_6919,N_4519,N_4059);
xnor U6920 (N_6920,N_3644,N_5729);
and U6921 (N_6921,N_5608,N_5898);
or U6922 (N_6922,N_5928,N_4792);
nor U6923 (N_6923,N_4481,N_5330);
nor U6924 (N_6924,N_4136,N_3161);
or U6925 (N_6925,N_3792,N_3578);
nor U6926 (N_6926,N_5909,N_5719);
xnor U6927 (N_6927,N_3697,N_3158);
nor U6928 (N_6928,N_4383,N_4817);
nand U6929 (N_6929,N_3984,N_4373);
or U6930 (N_6930,N_5715,N_5185);
nor U6931 (N_6931,N_4835,N_3067);
xor U6932 (N_6932,N_3250,N_5994);
nand U6933 (N_6933,N_5650,N_5216);
nand U6934 (N_6934,N_3365,N_3086);
nand U6935 (N_6935,N_3239,N_5129);
nand U6936 (N_6936,N_5036,N_5683);
nor U6937 (N_6937,N_4396,N_3556);
nor U6938 (N_6938,N_5264,N_4524);
and U6939 (N_6939,N_3962,N_3607);
xor U6940 (N_6940,N_3846,N_3587);
nor U6941 (N_6941,N_4788,N_3811);
nor U6942 (N_6942,N_5894,N_5498);
nor U6943 (N_6943,N_5835,N_3764);
xor U6944 (N_6944,N_3269,N_4866);
or U6945 (N_6945,N_3780,N_5754);
nor U6946 (N_6946,N_3813,N_5971);
xnor U6947 (N_6947,N_3449,N_4275);
nor U6948 (N_6948,N_3588,N_5636);
nand U6949 (N_6949,N_3634,N_3916);
or U6950 (N_6950,N_3329,N_3076);
nor U6951 (N_6951,N_4013,N_3869);
xor U6952 (N_6952,N_5277,N_4918);
and U6953 (N_6953,N_4979,N_5914);
nor U6954 (N_6954,N_3268,N_4214);
xor U6955 (N_6955,N_4472,N_4527);
xor U6956 (N_6956,N_5468,N_4461);
nand U6957 (N_6957,N_4992,N_5778);
nand U6958 (N_6958,N_5776,N_3586);
or U6959 (N_6959,N_3684,N_4173);
nand U6960 (N_6960,N_4062,N_3152);
or U6961 (N_6961,N_4014,N_4596);
nand U6962 (N_6962,N_4323,N_4209);
nor U6963 (N_6963,N_3378,N_5443);
nand U6964 (N_6964,N_3367,N_5996);
or U6965 (N_6965,N_3495,N_4999);
nand U6966 (N_6966,N_4374,N_5362);
nand U6967 (N_6967,N_3133,N_4987);
nand U6968 (N_6968,N_5459,N_5007);
xnor U6969 (N_6969,N_3987,N_3833);
nor U6970 (N_6970,N_4203,N_4544);
and U6971 (N_6971,N_4103,N_3451);
or U6972 (N_6972,N_3177,N_3492);
or U6973 (N_6973,N_3081,N_4660);
nand U6974 (N_6974,N_3716,N_3483);
and U6975 (N_6975,N_3680,N_3617);
nor U6976 (N_6976,N_4196,N_4213);
nand U6977 (N_6977,N_5050,N_5598);
nand U6978 (N_6978,N_5902,N_3348);
or U6979 (N_6979,N_5104,N_5843);
nor U6980 (N_6980,N_3613,N_4733);
xnor U6981 (N_6981,N_4117,N_3920);
and U6982 (N_6982,N_5849,N_5366);
or U6983 (N_6983,N_4985,N_4641);
nand U6984 (N_6984,N_5761,N_4611);
nor U6985 (N_6985,N_4993,N_3970);
nand U6986 (N_6986,N_5332,N_5226);
nor U6987 (N_6987,N_4297,N_5692);
xor U6988 (N_6988,N_4698,N_5577);
nor U6989 (N_6989,N_4579,N_4819);
and U6990 (N_6990,N_4293,N_5795);
nand U6991 (N_6991,N_5931,N_5070);
or U6992 (N_6992,N_4962,N_4326);
or U6993 (N_6993,N_3956,N_4281);
or U6994 (N_6994,N_5667,N_5906);
and U6995 (N_6995,N_3236,N_5343);
xor U6996 (N_6996,N_5542,N_3534);
and U6997 (N_6997,N_3335,N_3884);
xor U6998 (N_6998,N_3208,N_5767);
and U6999 (N_6999,N_3539,N_3078);
xor U7000 (N_7000,N_5417,N_4069);
nand U7001 (N_7001,N_4980,N_3064);
xor U7002 (N_7002,N_5732,N_3775);
and U7003 (N_7003,N_3385,N_5643);
nand U7004 (N_7004,N_3640,N_4176);
xor U7005 (N_7005,N_3830,N_5414);
nor U7006 (N_7006,N_5797,N_5817);
xnor U7007 (N_7007,N_4295,N_5272);
or U7008 (N_7008,N_4408,N_5194);
and U7009 (N_7009,N_5116,N_4608);
nand U7010 (N_7010,N_3374,N_5819);
xnor U7011 (N_7011,N_5798,N_4358);
or U7012 (N_7012,N_4017,N_3517);
or U7013 (N_7013,N_4042,N_4249);
nor U7014 (N_7014,N_3395,N_4857);
nand U7015 (N_7015,N_3043,N_3165);
nand U7016 (N_7016,N_4500,N_3457);
nand U7017 (N_7017,N_5983,N_5029);
or U7018 (N_7018,N_3039,N_4766);
and U7019 (N_7019,N_4391,N_4470);
xor U7020 (N_7020,N_3914,N_3898);
xnor U7021 (N_7021,N_5440,N_3038);
and U7022 (N_7022,N_4631,N_3510);
and U7023 (N_7023,N_5510,N_4978);
nor U7024 (N_7024,N_4413,N_5790);
xor U7025 (N_7025,N_3346,N_4809);
nand U7026 (N_7026,N_5263,N_3034);
or U7027 (N_7027,N_5960,N_4531);
nand U7028 (N_7028,N_5090,N_4247);
and U7029 (N_7029,N_5280,N_3726);
or U7030 (N_7030,N_4887,N_3416);
xor U7031 (N_7031,N_3545,N_4046);
nor U7032 (N_7032,N_5989,N_5568);
or U7033 (N_7033,N_5756,N_3023);
nor U7034 (N_7034,N_5209,N_3392);
xor U7035 (N_7035,N_4998,N_3093);
nor U7036 (N_7036,N_3772,N_4747);
xnor U7037 (N_7037,N_4838,N_4911);
nand U7038 (N_7038,N_4945,N_3289);
or U7039 (N_7039,N_4180,N_3388);
or U7040 (N_7040,N_3248,N_4748);
xnor U7041 (N_7041,N_4605,N_3373);
xnor U7042 (N_7042,N_3315,N_4032);
nor U7043 (N_7043,N_3431,N_5382);
nor U7044 (N_7044,N_3949,N_5922);
nand U7045 (N_7045,N_4922,N_4986);
nor U7046 (N_7046,N_3978,N_5320);
nand U7047 (N_7047,N_4910,N_4449);
and U7048 (N_7048,N_3735,N_5963);
and U7049 (N_7049,N_3317,N_4230);
or U7050 (N_7050,N_3281,N_5540);
nand U7051 (N_7051,N_4546,N_3362);
or U7052 (N_7052,N_3035,N_4680);
or U7053 (N_7053,N_3142,N_5268);
or U7054 (N_7054,N_5950,N_5725);
nand U7055 (N_7055,N_3569,N_5594);
and U7056 (N_7056,N_4863,N_3478);
nand U7057 (N_7057,N_3200,N_5965);
or U7058 (N_7058,N_3835,N_5051);
or U7059 (N_7059,N_5076,N_5127);
nor U7060 (N_7060,N_4593,N_3878);
nor U7061 (N_7061,N_4974,N_3853);
nor U7062 (N_7062,N_3945,N_3901);
xor U7063 (N_7063,N_3379,N_4826);
and U7064 (N_7064,N_4455,N_3342);
and U7065 (N_7065,N_4368,N_4466);
nor U7066 (N_7066,N_4580,N_4431);
nor U7067 (N_7067,N_3002,N_3763);
or U7068 (N_7068,N_4587,N_5039);
nand U7069 (N_7069,N_3493,N_5889);
or U7070 (N_7070,N_4445,N_3903);
or U7071 (N_7071,N_4067,N_5565);
or U7072 (N_7072,N_4736,N_4261);
nor U7073 (N_7073,N_4325,N_4385);
xnor U7074 (N_7074,N_5717,N_5337);
nand U7075 (N_7075,N_4732,N_5421);
and U7076 (N_7076,N_4303,N_3551);
and U7077 (N_7077,N_5661,N_4622);
or U7078 (N_7078,N_3598,N_5660);
or U7079 (N_7079,N_4301,N_5649);
xor U7080 (N_7080,N_3891,N_4109);
or U7081 (N_7081,N_3173,N_5281);
and U7082 (N_7082,N_5396,N_4344);
or U7083 (N_7083,N_4904,N_5939);
nor U7084 (N_7084,N_5863,N_5156);
xor U7085 (N_7085,N_5410,N_3777);
and U7086 (N_7086,N_5302,N_3320);
or U7087 (N_7087,N_5850,N_3802);
nor U7088 (N_7088,N_5485,N_3511);
xnor U7089 (N_7089,N_5282,N_5393);
xnor U7090 (N_7090,N_5177,N_4972);
nand U7091 (N_7091,N_5857,N_4119);
nand U7092 (N_7092,N_3384,N_3405);
xnor U7093 (N_7093,N_3410,N_3382);
and U7094 (N_7094,N_3111,N_3981);
and U7095 (N_7095,N_4664,N_5058);
xnor U7096 (N_7096,N_5625,N_4869);
xnor U7097 (N_7097,N_4003,N_4508);
nand U7098 (N_7098,N_3630,N_3557);
or U7099 (N_7099,N_5059,N_5631);
nand U7100 (N_7100,N_4129,N_4220);
and U7101 (N_7101,N_5882,N_5779);
or U7102 (N_7102,N_5442,N_4104);
or U7103 (N_7103,N_3020,N_3520);
nor U7104 (N_7104,N_5576,N_3406);
and U7105 (N_7105,N_3766,N_4228);
nand U7106 (N_7106,N_5685,N_5731);
nor U7107 (N_7107,N_4861,N_4908);
or U7108 (N_7108,N_4387,N_3185);
and U7109 (N_7109,N_4931,N_3084);
nand U7110 (N_7110,N_3364,N_4427);
and U7111 (N_7111,N_5298,N_3799);
xor U7112 (N_7112,N_4130,N_5451);
xor U7113 (N_7113,N_4711,N_3737);
and U7114 (N_7114,N_4523,N_5684);
xor U7115 (N_7115,N_5886,N_3816);
and U7116 (N_7116,N_5668,N_5408);
and U7117 (N_7117,N_3381,N_4542);
and U7118 (N_7118,N_5157,N_5322);
xor U7119 (N_7119,N_3179,N_3109);
nor U7120 (N_7120,N_3998,N_3455);
nor U7121 (N_7121,N_5163,N_3537);
and U7122 (N_7122,N_4578,N_5515);
nand U7123 (N_7123,N_5394,N_3178);
nor U7124 (N_7124,N_5547,N_4964);
nor U7125 (N_7125,N_3641,N_5318);
nand U7126 (N_7126,N_3553,N_5387);
xor U7127 (N_7127,N_5400,N_3421);
or U7128 (N_7128,N_3746,N_3781);
xnor U7129 (N_7129,N_4833,N_3749);
nand U7130 (N_7130,N_4392,N_4409);
and U7131 (N_7131,N_5604,N_5295);
nand U7132 (N_7132,N_4563,N_3922);
nor U7133 (N_7133,N_4201,N_4131);
and U7134 (N_7134,N_3176,N_5689);
nor U7135 (N_7135,N_5324,N_4253);
and U7136 (N_7136,N_3414,N_4454);
and U7137 (N_7137,N_5445,N_4574);
and U7138 (N_7138,N_3113,N_4484);
nor U7139 (N_7139,N_5513,N_5405);
nor U7140 (N_7140,N_5196,N_5564);
and U7141 (N_7141,N_5620,N_4840);
nor U7142 (N_7142,N_5391,N_5360);
and U7143 (N_7143,N_3314,N_3326);
xor U7144 (N_7144,N_4267,N_3839);
or U7145 (N_7145,N_5888,N_4886);
and U7146 (N_7146,N_4115,N_4635);
nand U7147 (N_7147,N_4160,N_4377);
and U7148 (N_7148,N_3032,N_3228);
nor U7149 (N_7149,N_5871,N_4090);
xnor U7150 (N_7150,N_4175,N_4102);
nand U7151 (N_7151,N_3924,N_3003);
and U7152 (N_7152,N_3769,N_5081);
and U7153 (N_7153,N_5274,N_5838);
nor U7154 (N_7154,N_3575,N_4737);
or U7155 (N_7155,N_4926,N_4889);
and U7156 (N_7156,N_5777,N_4221);
xor U7157 (N_7157,N_4606,N_4505);
nor U7158 (N_7158,N_4851,N_3077);
xnor U7159 (N_7159,N_5881,N_4570);
or U7160 (N_7160,N_5019,N_4880);
nor U7161 (N_7161,N_4451,N_5589);
nand U7162 (N_7162,N_5004,N_3182);
nor U7163 (N_7163,N_3773,N_3552);
xnor U7164 (N_7164,N_5191,N_4288);
nand U7165 (N_7165,N_3240,N_3983);
xnor U7166 (N_7166,N_3784,N_4898);
nor U7167 (N_7167,N_5506,N_5827);
and U7168 (N_7168,N_4146,N_3253);
nor U7169 (N_7169,N_3203,N_5384);
nand U7170 (N_7170,N_4010,N_3168);
xnor U7171 (N_7171,N_3838,N_5110);
xnor U7172 (N_7172,N_3016,N_3472);
nor U7173 (N_7173,N_4444,N_4200);
nand U7174 (N_7174,N_3503,N_3259);
xnor U7175 (N_7175,N_4028,N_5178);
nand U7176 (N_7176,N_3718,N_5203);
nand U7177 (N_7177,N_5694,N_4473);
or U7178 (N_7178,N_3021,N_4108);
or U7179 (N_7179,N_3008,N_4024);
nand U7180 (N_7180,N_4035,N_4367);
or U7181 (N_7181,N_5709,N_4206);
nor U7182 (N_7182,N_5801,N_3670);
or U7183 (N_7183,N_5031,N_4920);
nand U7184 (N_7184,N_3006,N_3074);
nand U7185 (N_7185,N_4822,N_3167);
or U7186 (N_7186,N_5875,N_4333);
nand U7187 (N_7187,N_3602,N_4939);
nor U7188 (N_7188,N_3308,N_5398);
xor U7189 (N_7189,N_3371,N_3708);
and U7190 (N_7190,N_3526,N_4820);
xor U7191 (N_7191,N_5688,N_4795);
nand U7192 (N_7192,N_4696,N_4352);
and U7193 (N_7193,N_4610,N_4510);
nor U7194 (N_7194,N_3274,N_3654);
or U7195 (N_7195,N_3146,N_3950);
nand U7196 (N_7196,N_4073,N_5495);
and U7197 (N_7197,N_5682,N_5003);
nor U7198 (N_7198,N_4313,N_5431);
or U7199 (N_7199,N_3827,N_4417);
or U7200 (N_7200,N_5524,N_5655);
xor U7201 (N_7201,N_4888,N_5600);
nand U7202 (N_7202,N_3687,N_3937);
nand U7203 (N_7203,N_3490,N_5406);
or U7204 (N_7204,N_5895,N_3115);
nand U7205 (N_7205,N_5834,N_3656);
xor U7206 (N_7206,N_3789,N_5873);
or U7207 (N_7207,N_5507,N_5238);
or U7208 (N_7208,N_5962,N_4744);
nor U7209 (N_7209,N_3722,N_3262);
or U7210 (N_7210,N_3948,N_3148);
nor U7211 (N_7211,N_5874,N_4543);
and U7212 (N_7212,N_4614,N_4620);
nor U7213 (N_7213,N_3159,N_3290);
and U7214 (N_7214,N_5727,N_3303);
or U7215 (N_7215,N_5810,N_5552);
or U7216 (N_7216,N_3888,N_3052);
and U7217 (N_7217,N_5085,N_4894);
xor U7218 (N_7218,N_3435,N_4842);
nor U7219 (N_7219,N_5934,N_4089);
or U7220 (N_7220,N_3928,N_5082);
or U7221 (N_7221,N_5014,N_3533);
nor U7222 (N_7222,N_4607,N_3130);
xnor U7223 (N_7223,N_4884,N_3225);
nand U7224 (N_7224,N_5832,N_4162);
or U7225 (N_7225,N_3865,N_4723);
or U7226 (N_7226,N_5390,N_3645);
and U7227 (N_7227,N_4491,N_5013);
and U7228 (N_7228,N_4279,N_4872);
or U7229 (N_7229,N_3599,N_3566);
nand U7230 (N_7230,N_4124,N_4395);
or U7231 (N_7231,N_3969,N_5136);
or U7232 (N_7232,N_4390,N_3132);
nor U7233 (N_7233,N_4909,N_4410);
or U7234 (N_7234,N_4946,N_3438);
or U7235 (N_7235,N_4416,N_5639);
or U7236 (N_7236,N_3092,N_3263);
or U7237 (N_7237,N_4769,N_3779);
or U7238 (N_7238,N_4699,N_4789);
and U7239 (N_7239,N_4716,N_4277);
or U7240 (N_7240,N_3549,N_4957);
nand U7241 (N_7241,N_4474,N_3693);
nand U7242 (N_7242,N_5168,N_5022);
or U7243 (N_7243,N_5009,N_3906);
nand U7244 (N_7244,N_5484,N_3801);
and U7245 (N_7245,N_5806,N_3171);
nor U7246 (N_7246,N_4839,N_5762);
and U7247 (N_7247,N_5578,N_4029);
nor U7248 (N_7248,N_5113,N_5803);
and U7249 (N_7249,N_5561,N_3235);
xnor U7250 (N_7250,N_3129,N_5699);
and U7251 (N_7251,N_5704,N_5551);
and U7252 (N_7252,N_3467,N_5940);
nand U7253 (N_7253,N_4569,N_4257);
or U7254 (N_7254,N_5239,N_3946);
nand U7255 (N_7255,N_4613,N_4560);
nand U7256 (N_7256,N_4475,N_5935);
nor U7257 (N_7257,N_4685,N_4376);
xnor U7258 (N_7258,N_3267,N_3347);
xnor U7259 (N_7259,N_4501,N_4638);
and U7260 (N_7260,N_4675,N_3089);
nand U7261 (N_7261,N_5271,N_5915);
or U7262 (N_7262,N_3993,N_3767);
xor U7263 (N_7263,N_5167,N_3995);
xnor U7264 (N_7264,N_3282,N_5710);
or U7265 (N_7265,N_3190,N_4423);
xor U7266 (N_7266,N_5215,N_3121);
and U7267 (N_7267,N_5815,N_4022);
or U7268 (N_7268,N_4246,N_3700);
nand U7269 (N_7269,N_5866,N_3623);
or U7270 (N_7270,N_3481,N_4434);
nor U7271 (N_7271,N_5115,N_4357);
nand U7272 (N_7272,N_5389,N_4677);
nor U7273 (N_7273,N_4021,N_5065);
nor U7274 (N_7274,N_4248,N_3851);
nand U7275 (N_7275,N_4071,N_3574);
or U7276 (N_7276,N_5664,N_5500);
nor U7277 (N_7277,N_3476,N_4258);
xnor U7278 (N_7278,N_3936,N_5240);
nor U7279 (N_7279,N_3734,N_5919);
and U7280 (N_7280,N_4623,N_3786);
nor U7281 (N_7281,N_5235,N_4370);
xnor U7282 (N_7282,N_4154,N_3193);
nand U7283 (N_7283,N_4150,N_5723);
nand U7284 (N_7284,N_3498,N_3014);
nor U7285 (N_7285,N_4713,N_4561);
nor U7286 (N_7286,N_3243,N_4265);
nand U7287 (N_7287,N_3275,N_4340);
and U7288 (N_7288,N_3541,N_3550);
nand U7289 (N_7289,N_5146,N_5288);
and U7290 (N_7290,N_4254,N_5759);
nor U7291 (N_7291,N_3698,N_4381);
nor U7292 (N_7292,N_5712,N_5062);
and U7293 (N_7293,N_5183,N_3933);
nor U7294 (N_7294,N_3028,N_4642);
nor U7295 (N_7295,N_3604,N_5851);
xor U7296 (N_7296,N_5063,N_5143);
or U7297 (N_7297,N_5733,N_5760);
xnor U7298 (N_7298,N_3026,N_3855);
nor U7299 (N_7299,N_5670,N_3582);
and U7300 (N_7300,N_5691,N_3063);
and U7301 (N_7301,N_3468,N_5454);
or U7302 (N_7302,N_3991,N_3620);
and U7303 (N_7303,N_5686,N_5703);
xnor U7304 (N_7304,N_3513,N_5046);
nor U7305 (N_7305,N_3570,N_5346);
nor U7306 (N_7306,N_5845,N_4738);
xnor U7307 (N_7307,N_5208,N_4903);
xnor U7308 (N_7308,N_3404,N_3300);
or U7309 (N_7309,N_4832,N_3818);
and U7310 (N_7310,N_3921,N_4487);
xnor U7311 (N_7311,N_5899,N_4734);
nor U7312 (N_7312,N_5783,N_5766);
and U7313 (N_7313,N_4612,N_3471);
and U7314 (N_7314,N_5728,N_4393);
or U7315 (N_7315,N_4347,N_3867);
and U7316 (N_7316,N_5446,N_3815);
xnor U7317 (N_7317,N_3929,N_3522);
nor U7318 (N_7318,N_5750,N_4198);
or U7319 (N_7319,N_4767,N_3536);
nand U7320 (N_7320,N_4557,N_3774);
nand U7321 (N_7321,N_4224,N_5720);
nor U7322 (N_7322,N_4865,N_4105);
or U7323 (N_7323,N_4648,N_5680);
and U7324 (N_7324,N_4740,N_3669);
or U7325 (N_7325,N_5246,N_3619);
xor U7326 (N_7326,N_4429,N_3037);
nor U7327 (N_7327,N_3988,N_5610);
nand U7328 (N_7328,N_5466,N_5220);
nand U7329 (N_7329,N_3114,N_5057);
nor U7330 (N_7330,N_3487,N_5135);
nor U7331 (N_7331,N_4337,N_5244);
and U7332 (N_7332,N_5883,N_4975);
nor U7333 (N_7333,N_4768,N_5690);
xor U7334 (N_7334,N_5034,N_4760);
or U7335 (N_7335,N_5279,N_4226);
xor U7336 (N_7336,N_5679,N_5181);
xor U7337 (N_7337,N_4477,N_4750);
xnor U7338 (N_7338,N_4594,N_4672);
nand U7339 (N_7339,N_4727,N_3175);
xor U7340 (N_7340,N_5486,N_3628);
nand U7341 (N_7341,N_4329,N_4188);
nor U7342 (N_7342,N_4893,N_5529);
and U7343 (N_7343,N_3459,N_5450);
xnor U7344 (N_7344,N_4599,N_4121);
nor U7345 (N_7345,N_3345,N_4270);
xor U7346 (N_7346,N_4210,N_5107);
nor U7347 (N_7347,N_4950,N_4132);
and U7348 (N_7348,N_5979,N_5118);
nor U7349 (N_7349,N_5339,N_4710);
nand U7350 (N_7350,N_3860,N_5461);
nand U7351 (N_7351,N_4943,N_3548);
and U7352 (N_7352,N_4002,N_5641);
and U7353 (N_7353,N_3229,N_5427);
nor U7354 (N_7354,N_3882,N_3959);
nand U7355 (N_7355,N_3930,N_5432);
xnor U7356 (N_7356,N_3646,N_3627);
and U7357 (N_7357,N_3186,N_4803);
xnor U7358 (N_7358,N_3219,N_3390);
nand U7359 (N_7359,N_4673,N_4360);
nand U7360 (N_7360,N_4663,N_5912);
nand U7361 (N_7361,N_4552,N_5585);
or U7362 (N_7362,N_4643,N_4700);
and U7363 (N_7363,N_3117,N_4110);
nand U7364 (N_7364,N_4585,N_4361);
and U7365 (N_7365,N_4516,N_5659);
nor U7366 (N_7366,N_5628,N_3150);
nor U7367 (N_7367,N_3360,N_4078);
nor U7368 (N_7368,N_4731,N_5852);
nor U7369 (N_7369,N_4125,N_3191);
and U7370 (N_7370,N_5616,N_5868);
nor U7371 (N_7371,N_3432,N_4897);
and U7372 (N_7372,N_3692,N_5602);
nand U7373 (N_7373,N_5968,N_3989);
xor U7374 (N_7374,N_5574,N_4489);
and U7375 (N_7375,N_4953,N_3883);
xnor U7376 (N_7376,N_3671,N_4513);
xor U7377 (N_7377,N_4499,N_3439);
nand U7378 (N_7378,N_5420,N_4202);
nand U7379 (N_7379,N_5278,N_3649);
or U7380 (N_7380,N_5091,N_4707);
xor U7381 (N_7381,N_5993,N_3144);
and U7382 (N_7382,N_5375,N_5254);
or U7383 (N_7383,N_5821,N_3712);
nor U7384 (N_7384,N_4621,N_3318);
or U7385 (N_7385,N_5195,N_4058);
and U7386 (N_7386,N_3482,N_3714);
or U7387 (N_7387,N_4522,N_3183);
nor U7388 (N_7388,N_3900,N_3222);
and U7389 (N_7389,N_3579,N_4004);
and U7390 (N_7390,N_4074,N_4743);
nand U7391 (N_7391,N_4948,N_3568);
and U7392 (N_7392,N_3358,N_3624);
nor U7393 (N_7393,N_3958,N_5654);
and U7394 (N_7394,N_5383,N_4942);
nor U7395 (N_7395,N_3417,N_3821);
or U7396 (N_7396,N_4469,N_3220);
xnor U7397 (N_7397,N_5800,N_5102);
nor U7398 (N_7398,N_4583,N_3424);
or U7399 (N_7399,N_5837,N_3990);
nor U7400 (N_7400,N_4274,N_4791);
or U7401 (N_7401,N_4629,N_5437);
or U7402 (N_7402,N_3934,N_4339);
nor U7403 (N_7403,N_5049,N_4882);
and U7404 (N_7404,N_3915,N_4818);
nand U7405 (N_7405,N_4907,N_4464);
or U7406 (N_7406,N_3831,N_3926);
or U7407 (N_7407,N_3280,N_3196);
nor U7408 (N_7408,N_3258,N_5541);
or U7409 (N_7409,N_3119,N_4794);
nor U7410 (N_7410,N_5802,N_3319);
xnor U7411 (N_7411,N_3600,N_3905);
and U7412 (N_7412,N_3033,N_5367);
and U7413 (N_7413,N_5516,N_4969);
or U7414 (N_7414,N_3876,N_3819);
nand U7415 (N_7415,N_4116,N_5844);
or U7416 (N_7416,N_5596,N_4007);
and U7417 (N_7417,N_3297,N_3140);
xor U7418 (N_7418,N_5132,N_4995);
nor U7419 (N_7419,N_3854,N_4815);
or U7420 (N_7420,N_5644,N_4064);
nor U7421 (N_7421,N_4490,N_5477);
and U7422 (N_7422,N_4356,N_3542);
xor U7423 (N_7423,N_5333,N_4483);
or U7424 (N_7424,N_3209,N_3470);
and U7425 (N_7425,N_5232,N_4982);
or U7426 (N_7426,N_5755,N_5536);
and U7427 (N_7427,N_4384,N_3753);
nor U7428 (N_7428,N_4785,N_5666);
nor U7429 (N_7429,N_3053,N_3189);
xnor U7430 (N_7430,N_5716,N_3126);
nor U7431 (N_7431,N_4050,N_5591);
nor U7432 (N_7432,N_5328,N_3199);
nor U7433 (N_7433,N_5785,N_4092);
and U7434 (N_7434,N_4676,N_5763);
nor U7435 (N_7435,N_3058,N_4122);
nand U7436 (N_7436,N_5566,N_3745);
xor U7437 (N_7437,N_4245,N_3447);
xnor U7438 (N_7438,N_5283,N_5386);
or U7439 (N_7439,N_4452,N_5839);
nand U7440 (N_7440,N_3547,N_4045);
nand U7441 (N_7441,N_4639,N_5538);
nand U7442 (N_7442,N_5917,N_4037);
nand U7443 (N_7443,N_4963,N_4488);
and U7444 (N_7444,N_3807,N_4515);
nor U7445 (N_7445,N_3419,N_3527);
nand U7446 (N_7446,N_4741,N_5736);
xor U7447 (N_7447,N_4343,N_4571);
xnor U7448 (N_7448,N_5392,N_5086);
xnor U7449 (N_7449,N_5605,N_5509);
nand U7450 (N_7450,N_5449,N_5024);
and U7451 (N_7451,N_3803,N_5980);
xor U7452 (N_7452,N_5981,N_4679);
or U7453 (N_7453,N_4165,N_5130);
and U7454 (N_7454,N_3068,N_3341);
xor U7455 (N_7455,N_3400,N_4242);
or U7456 (N_7456,N_5207,N_4603);
or U7457 (N_7457,N_5544,N_4135);
nand U7458 (N_7458,N_5243,N_4118);
nand U7459 (N_7459,N_4786,N_4169);
and U7460 (N_7460,N_3466,N_4236);
or U7461 (N_7461,N_3584,N_3024);
nand U7462 (N_7462,N_5275,N_3147);
nand U7463 (N_7463,N_4532,N_5663);
nand U7464 (N_7464,N_5967,N_5718);
nand U7465 (N_7465,N_3386,N_4312);
nand U7466 (N_7466,N_5154,N_5910);
nor U7467 (N_7467,N_4615,N_3085);
nand U7468 (N_7468,N_4597,N_5097);
and U7469 (N_7469,N_3947,N_5611);
nand U7470 (N_7470,N_4665,N_5771);
xnor U7471 (N_7471,N_4644,N_5047);
and U7472 (N_7472,N_3355,N_4858);
nand U7473 (N_7473,N_4044,N_3366);
nand U7474 (N_7474,N_4671,N_4342);
xor U7475 (N_7475,N_3875,N_5068);
xor U7476 (N_7476,N_5284,N_5926);
xor U7477 (N_7477,N_5651,N_5078);
xor U7478 (N_7478,N_5455,N_5784);
nor U7479 (N_7479,N_5044,N_4589);
and U7480 (N_7480,N_3508,N_3581);
and U7481 (N_7481,N_5255,N_5192);
nor U7482 (N_7482,N_4966,N_3612);
nor U7483 (N_7483,N_5306,N_3702);
nor U7484 (N_7484,N_4706,N_5098);
and U7485 (N_7485,N_3573,N_5562);
nor U7486 (N_7486,N_4120,N_5148);
or U7487 (N_7487,N_4529,N_3966);
or U7488 (N_7488,N_3456,N_3194);
or U7489 (N_7489,N_4686,N_5482);
nand U7490 (N_7490,N_4241,N_3007);
xor U7491 (N_7491,N_3100,N_4038);
nor U7492 (N_7492,N_4598,N_3413);
or U7493 (N_7493,N_4272,N_5588);
and U7494 (N_7494,N_5705,N_5021);
nor U7495 (N_7495,N_4207,N_5982);
nand U7496 (N_7496,N_4829,N_5112);
and U7497 (N_7497,N_3075,N_4841);
nor U7498 (N_7498,N_5774,N_4167);
nor U7499 (N_7499,N_5913,N_4479);
nor U7500 (N_7500,N_3548,N_5211);
and U7501 (N_7501,N_4196,N_4334);
xor U7502 (N_7502,N_3999,N_5994);
or U7503 (N_7503,N_3910,N_4299);
or U7504 (N_7504,N_5547,N_5176);
nor U7505 (N_7505,N_5531,N_4431);
nand U7506 (N_7506,N_3518,N_4717);
nor U7507 (N_7507,N_3903,N_3484);
and U7508 (N_7508,N_5477,N_4160);
nor U7509 (N_7509,N_3078,N_4975);
and U7510 (N_7510,N_5813,N_5339);
nor U7511 (N_7511,N_4762,N_4361);
xnor U7512 (N_7512,N_3125,N_5223);
or U7513 (N_7513,N_4269,N_3286);
xor U7514 (N_7514,N_5555,N_4654);
xor U7515 (N_7515,N_3625,N_4545);
xor U7516 (N_7516,N_3992,N_4867);
or U7517 (N_7517,N_4932,N_4651);
nand U7518 (N_7518,N_5979,N_3249);
and U7519 (N_7519,N_3530,N_4679);
xor U7520 (N_7520,N_4687,N_5112);
xor U7521 (N_7521,N_5774,N_5197);
xnor U7522 (N_7522,N_3810,N_3901);
xnor U7523 (N_7523,N_4592,N_4643);
nor U7524 (N_7524,N_3804,N_4741);
and U7525 (N_7525,N_3171,N_5095);
xnor U7526 (N_7526,N_3228,N_5546);
xnor U7527 (N_7527,N_4858,N_4933);
nand U7528 (N_7528,N_4203,N_3621);
and U7529 (N_7529,N_5191,N_3163);
xnor U7530 (N_7530,N_4157,N_4521);
and U7531 (N_7531,N_3971,N_4394);
xor U7532 (N_7532,N_4614,N_5583);
nor U7533 (N_7533,N_5235,N_3669);
nor U7534 (N_7534,N_5425,N_3631);
or U7535 (N_7535,N_4286,N_4391);
nor U7536 (N_7536,N_5528,N_4410);
nor U7537 (N_7537,N_4106,N_5525);
nand U7538 (N_7538,N_5556,N_3182);
nor U7539 (N_7539,N_3722,N_3415);
nor U7540 (N_7540,N_3241,N_4642);
and U7541 (N_7541,N_5319,N_3032);
nor U7542 (N_7542,N_5593,N_4198);
xor U7543 (N_7543,N_4391,N_4021);
xnor U7544 (N_7544,N_3445,N_5111);
nand U7545 (N_7545,N_3184,N_4401);
nand U7546 (N_7546,N_3658,N_3198);
and U7547 (N_7547,N_3233,N_5404);
xnor U7548 (N_7548,N_4756,N_3455);
or U7549 (N_7549,N_5820,N_4341);
xnor U7550 (N_7550,N_3371,N_3049);
nand U7551 (N_7551,N_4941,N_4547);
or U7552 (N_7552,N_3172,N_4759);
nand U7553 (N_7553,N_5829,N_5005);
or U7554 (N_7554,N_5803,N_4938);
nor U7555 (N_7555,N_4634,N_5624);
nand U7556 (N_7556,N_5238,N_5434);
nor U7557 (N_7557,N_4314,N_4845);
and U7558 (N_7558,N_4934,N_4503);
xnor U7559 (N_7559,N_4837,N_3368);
xnor U7560 (N_7560,N_4463,N_4216);
nor U7561 (N_7561,N_5903,N_3766);
nand U7562 (N_7562,N_3556,N_4496);
or U7563 (N_7563,N_5448,N_3778);
or U7564 (N_7564,N_5365,N_5678);
nand U7565 (N_7565,N_5168,N_3110);
xnor U7566 (N_7566,N_5991,N_4068);
nand U7567 (N_7567,N_3149,N_5741);
nor U7568 (N_7568,N_4023,N_4322);
or U7569 (N_7569,N_5608,N_4151);
or U7570 (N_7570,N_3396,N_5912);
nor U7571 (N_7571,N_5443,N_3458);
nand U7572 (N_7572,N_3294,N_4437);
and U7573 (N_7573,N_3144,N_3164);
xor U7574 (N_7574,N_5098,N_3582);
or U7575 (N_7575,N_5567,N_4096);
or U7576 (N_7576,N_5902,N_5204);
xor U7577 (N_7577,N_4769,N_5142);
nand U7578 (N_7578,N_3620,N_5592);
nor U7579 (N_7579,N_5057,N_3345);
nor U7580 (N_7580,N_4166,N_3186);
nand U7581 (N_7581,N_4527,N_3721);
nand U7582 (N_7582,N_3985,N_5053);
nand U7583 (N_7583,N_4853,N_4749);
xnor U7584 (N_7584,N_3549,N_5483);
and U7585 (N_7585,N_4318,N_3806);
or U7586 (N_7586,N_3349,N_4240);
or U7587 (N_7587,N_3417,N_3676);
nand U7588 (N_7588,N_3989,N_5448);
nand U7589 (N_7589,N_4392,N_4611);
and U7590 (N_7590,N_5894,N_5841);
nand U7591 (N_7591,N_5948,N_4372);
xor U7592 (N_7592,N_5800,N_4987);
nor U7593 (N_7593,N_3129,N_3967);
nand U7594 (N_7594,N_5161,N_4821);
and U7595 (N_7595,N_5277,N_5489);
and U7596 (N_7596,N_5495,N_4033);
nand U7597 (N_7597,N_4398,N_5868);
nand U7598 (N_7598,N_5055,N_3910);
nand U7599 (N_7599,N_4707,N_4353);
xor U7600 (N_7600,N_4168,N_4505);
xnor U7601 (N_7601,N_4665,N_4344);
nor U7602 (N_7602,N_3971,N_4624);
and U7603 (N_7603,N_3791,N_4671);
and U7604 (N_7604,N_5430,N_3105);
nand U7605 (N_7605,N_3604,N_4493);
xor U7606 (N_7606,N_5156,N_4444);
nor U7607 (N_7607,N_3078,N_3522);
nor U7608 (N_7608,N_5045,N_4516);
and U7609 (N_7609,N_3835,N_4631);
or U7610 (N_7610,N_3851,N_5396);
and U7611 (N_7611,N_4947,N_4382);
nand U7612 (N_7612,N_5549,N_5430);
and U7613 (N_7613,N_4611,N_4936);
xor U7614 (N_7614,N_5205,N_4868);
nand U7615 (N_7615,N_5804,N_3744);
or U7616 (N_7616,N_4614,N_3324);
nand U7617 (N_7617,N_3170,N_3272);
or U7618 (N_7618,N_3322,N_4470);
nand U7619 (N_7619,N_4101,N_5335);
and U7620 (N_7620,N_4902,N_5664);
nor U7621 (N_7621,N_5597,N_3742);
nor U7622 (N_7622,N_5084,N_5123);
xnor U7623 (N_7623,N_5775,N_4214);
nand U7624 (N_7624,N_5240,N_5444);
or U7625 (N_7625,N_5467,N_4614);
nor U7626 (N_7626,N_5618,N_4318);
nor U7627 (N_7627,N_3920,N_3602);
xor U7628 (N_7628,N_3878,N_3356);
and U7629 (N_7629,N_4273,N_4716);
and U7630 (N_7630,N_3441,N_5108);
and U7631 (N_7631,N_3861,N_5474);
or U7632 (N_7632,N_4273,N_4147);
and U7633 (N_7633,N_5905,N_5275);
nand U7634 (N_7634,N_5854,N_4663);
or U7635 (N_7635,N_3973,N_3438);
nand U7636 (N_7636,N_5602,N_4525);
or U7637 (N_7637,N_4718,N_3532);
xnor U7638 (N_7638,N_5157,N_4166);
or U7639 (N_7639,N_3033,N_3109);
and U7640 (N_7640,N_4634,N_3334);
or U7641 (N_7641,N_5384,N_3297);
or U7642 (N_7642,N_3749,N_5594);
or U7643 (N_7643,N_3812,N_3082);
nor U7644 (N_7644,N_4393,N_4364);
nor U7645 (N_7645,N_4981,N_5667);
nor U7646 (N_7646,N_5300,N_5274);
or U7647 (N_7647,N_4195,N_5793);
and U7648 (N_7648,N_4025,N_4908);
or U7649 (N_7649,N_5534,N_5443);
and U7650 (N_7650,N_4830,N_5439);
nor U7651 (N_7651,N_3918,N_3584);
or U7652 (N_7652,N_4703,N_5866);
or U7653 (N_7653,N_3967,N_5152);
xnor U7654 (N_7654,N_3372,N_4013);
nor U7655 (N_7655,N_4188,N_3441);
or U7656 (N_7656,N_3344,N_5939);
nor U7657 (N_7657,N_3394,N_4272);
and U7658 (N_7658,N_3875,N_5005);
nand U7659 (N_7659,N_5106,N_3627);
and U7660 (N_7660,N_5465,N_4848);
nand U7661 (N_7661,N_3201,N_4277);
or U7662 (N_7662,N_3994,N_4728);
nor U7663 (N_7663,N_4239,N_5040);
xor U7664 (N_7664,N_5582,N_3678);
or U7665 (N_7665,N_3578,N_3234);
xnor U7666 (N_7666,N_3227,N_5041);
nor U7667 (N_7667,N_5719,N_3374);
or U7668 (N_7668,N_4868,N_4411);
or U7669 (N_7669,N_4707,N_4218);
and U7670 (N_7670,N_4049,N_5489);
or U7671 (N_7671,N_4288,N_4197);
nor U7672 (N_7672,N_3900,N_3476);
and U7673 (N_7673,N_3158,N_3323);
or U7674 (N_7674,N_5911,N_4260);
and U7675 (N_7675,N_3215,N_5438);
nand U7676 (N_7676,N_4395,N_4081);
and U7677 (N_7677,N_5085,N_4090);
xnor U7678 (N_7678,N_4598,N_4863);
or U7679 (N_7679,N_5626,N_4748);
nand U7680 (N_7680,N_4321,N_4867);
or U7681 (N_7681,N_3714,N_3992);
xnor U7682 (N_7682,N_5491,N_3406);
and U7683 (N_7683,N_5026,N_4316);
or U7684 (N_7684,N_5033,N_5167);
xor U7685 (N_7685,N_4187,N_4587);
and U7686 (N_7686,N_4260,N_5611);
nand U7687 (N_7687,N_5174,N_3884);
nand U7688 (N_7688,N_5935,N_4003);
and U7689 (N_7689,N_4185,N_5037);
or U7690 (N_7690,N_5089,N_5397);
xnor U7691 (N_7691,N_5691,N_3597);
or U7692 (N_7692,N_4470,N_3196);
nor U7693 (N_7693,N_3280,N_3367);
nand U7694 (N_7694,N_4900,N_4774);
nand U7695 (N_7695,N_5311,N_4794);
xor U7696 (N_7696,N_3108,N_3271);
nor U7697 (N_7697,N_5063,N_3209);
nand U7698 (N_7698,N_3863,N_4122);
nand U7699 (N_7699,N_4723,N_5326);
xor U7700 (N_7700,N_3785,N_4791);
nor U7701 (N_7701,N_4151,N_4136);
xnor U7702 (N_7702,N_5757,N_4598);
xor U7703 (N_7703,N_5740,N_4343);
and U7704 (N_7704,N_4978,N_5778);
nand U7705 (N_7705,N_3486,N_3265);
nand U7706 (N_7706,N_3564,N_4088);
nand U7707 (N_7707,N_3719,N_3706);
and U7708 (N_7708,N_3495,N_4153);
nand U7709 (N_7709,N_5500,N_3410);
xor U7710 (N_7710,N_5540,N_4756);
nor U7711 (N_7711,N_3894,N_5214);
nand U7712 (N_7712,N_3521,N_3031);
and U7713 (N_7713,N_4046,N_4896);
and U7714 (N_7714,N_4122,N_3927);
or U7715 (N_7715,N_4399,N_4267);
or U7716 (N_7716,N_3990,N_5032);
xor U7717 (N_7717,N_4917,N_3826);
nor U7718 (N_7718,N_5583,N_5195);
xor U7719 (N_7719,N_4695,N_5715);
and U7720 (N_7720,N_3468,N_4873);
xor U7721 (N_7721,N_4434,N_3283);
nor U7722 (N_7722,N_3857,N_3837);
or U7723 (N_7723,N_5843,N_4814);
and U7724 (N_7724,N_4548,N_4745);
and U7725 (N_7725,N_4674,N_4687);
or U7726 (N_7726,N_4531,N_5329);
or U7727 (N_7727,N_4349,N_5767);
nand U7728 (N_7728,N_4318,N_5527);
or U7729 (N_7729,N_5361,N_4744);
and U7730 (N_7730,N_3649,N_5279);
or U7731 (N_7731,N_5636,N_4605);
or U7732 (N_7732,N_4062,N_3562);
xor U7733 (N_7733,N_3670,N_4067);
and U7734 (N_7734,N_5132,N_4856);
and U7735 (N_7735,N_5432,N_5118);
or U7736 (N_7736,N_3087,N_4612);
nor U7737 (N_7737,N_4395,N_4806);
and U7738 (N_7738,N_5861,N_4121);
and U7739 (N_7739,N_4500,N_3906);
xor U7740 (N_7740,N_5316,N_4102);
xor U7741 (N_7741,N_4096,N_3727);
nand U7742 (N_7742,N_5857,N_5684);
nor U7743 (N_7743,N_4531,N_3927);
xor U7744 (N_7744,N_3893,N_5268);
nor U7745 (N_7745,N_3570,N_4879);
nor U7746 (N_7746,N_5914,N_5047);
nand U7747 (N_7747,N_4037,N_5021);
or U7748 (N_7748,N_5994,N_3506);
and U7749 (N_7749,N_3563,N_5538);
or U7750 (N_7750,N_4544,N_5169);
xor U7751 (N_7751,N_4925,N_3252);
and U7752 (N_7752,N_4500,N_5706);
and U7753 (N_7753,N_4567,N_4291);
xnor U7754 (N_7754,N_5257,N_5992);
xor U7755 (N_7755,N_3899,N_3497);
and U7756 (N_7756,N_5714,N_5987);
or U7757 (N_7757,N_5456,N_4117);
or U7758 (N_7758,N_4576,N_4037);
nor U7759 (N_7759,N_5769,N_3558);
xor U7760 (N_7760,N_4725,N_5312);
nand U7761 (N_7761,N_3550,N_3164);
nand U7762 (N_7762,N_5085,N_4948);
nor U7763 (N_7763,N_3020,N_3936);
xor U7764 (N_7764,N_4581,N_5950);
or U7765 (N_7765,N_4050,N_3871);
and U7766 (N_7766,N_4836,N_5969);
nor U7767 (N_7767,N_5515,N_5665);
nor U7768 (N_7768,N_3356,N_3367);
xor U7769 (N_7769,N_3629,N_4281);
nor U7770 (N_7770,N_5606,N_5363);
or U7771 (N_7771,N_4399,N_4305);
nor U7772 (N_7772,N_4131,N_4241);
nor U7773 (N_7773,N_3129,N_4041);
xnor U7774 (N_7774,N_3516,N_5543);
nand U7775 (N_7775,N_4388,N_5422);
nand U7776 (N_7776,N_3407,N_3518);
nor U7777 (N_7777,N_5107,N_3027);
or U7778 (N_7778,N_5647,N_4938);
nor U7779 (N_7779,N_3185,N_4797);
nand U7780 (N_7780,N_4273,N_3478);
and U7781 (N_7781,N_5885,N_5813);
xor U7782 (N_7782,N_5761,N_3011);
or U7783 (N_7783,N_5360,N_5358);
and U7784 (N_7784,N_5731,N_3194);
nor U7785 (N_7785,N_5791,N_3528);
nand U7786 (N_7786,N_4986,N_5686);
nor U7787 (N_7787,N_3941,N_4399);
xor U7788 (N_7788,N_3612,N_4245);
xor U7789 (N_7789,N_3566,N_3268);
nor U7790 (N_7790,N_4687,N_5741);
or U7791 (N_7791,N_3063,N_4955);
and U7792 (N_7792,N_3755,N_5726);
or U7793 (N_7793,N_4276,N_5651);
or U7794 (N_7794,N_5316,N_5746);
nand U7795 (N_7795,N_5557,N_5983);
xnor U7796 (N_7796,N_4911,N_5307);
nand U7797 (N_7797,N_3914,N_5327);
nor U7798 (N_7798,N_5361,N_4400);
xnor U7799 (N_7799,N_3528,N_5951);
and U7800 (N_7800,N_5462,N_4669);
nor U7801 (N_7801,N_5163,N_3430);
and U7802 (N_7802,N_3156,N_4317);
nand U7803 (N_7803,N_4622,N_4882);
and U7804 (N_7804,N_4740,N_5773);
and U7805 (N_7805,N_4423,N_4462);
nor U7806 (N_7806,N_4497,N_5053);
xor U7807 (N_7807,N_4951,N_5812);
xor U7808 (N_7808,N_4879,N_4745);
xor U7809 (N_7809,N_5949,N_3242);
or U7810 (N_7810,N_4288,N_5020);
or U7811 (N_7811,N_3211,N_3790);
nor U7812 (N_7812,N_3913,N_5077);
and U7813 (N_7813,N_3367,N_5706);
nor U7814 (N_7814,N_5654,N_3972);
and U7815 (N_7815,N_3851,N_5232);
nor U7816 (N_7816,N_3573,N_5600);
xor U7817 (N_7817,N_3960,N_4109);
or U7818 (N_7818,N_4014,N_4683);
nand U7819 (N_7819,N_5697,N_3452);
nor U7820 (N_7820,N_5461,N_3140);
xnor U7821 (N_7821,N_3941,N_3521);
nor U7822 (N_7822,N_4605,N_4608);
or U7823 (N_7823,N_5576,N_4406);
nor U7824 (N_7824,N_4976,N_3263);
or U7825 (N_7825,N_5923,N_3346);
and U7826 (N_7826,N_3982,N_4464);
and U7827 (N_7827,N_4119,N_5330);
and U7828 (N_7828,N_4441,N_3309);
nand U7829 (N_7829,N_5559,N_4497);
nor U7830 (N_7830,N_3779,N_3412);
and U7831 (N_7831,N_4265,N_3208);
nand U7832 (N_7832,N_4367,N_4186);
nor U7833 (N_7833,N_3477,N_3319);
and U7834 (N_7834,N_5284,N_4050);
xor U7835 (N_7835,N_5146,N_3861);
nor U7836 (N_7836,N_4714,N_5644);
nand U7837 (N_7837,N_3098,N_3286);
nand U7838 (N_7838,N_5143,N_4568);
or U7839 (N_7839,N_3090,N_3384);
and U7840 (N_7840,N_4672,N_5441);
nand U7841 (N_7841,N_4070,N_5395);
nor U7842 (N_7842,N_3638,N_4004);
xor U7843 (N_7843,N_3590,N_5065);
nor U7844 (N_7844,N_4863,N_4740);
nand U7845 (N_7845,N_5577,N_3384);
xor U7846 (N_7846,N_4581,N_5399);
xnor U7847 (N_7847,N_3476,N_3866);
nor U7848 (N_7848,N_4162,N_5398);
xor U7849 (N_7849,N_3467,N_3393);
and U7850 (N_7850,N_4524,N_4789);
and U7851 (N_7851,N_3659,N_4908);
and U7852 (N_7852,N_5368,N_4745);
xor U7853 (N_7853,N_3093,N_4721);
nor U7854 (N_7854,N_4896,N_3034);
and U7855 (N_7855,N_4387,N_4274);
nand U7856 (N_7856,N_3401,N_5916);
nor U7857 (N_7857,N_4583,N_4545);
and U7858 (N_7858,N_4570,N_5198);
or U7859 (N_7859,N_4818,N_5840);
or U7860 (N_7860,N_4040,N_3987);
xor U7861 (N_7861,N_4107,N_3960);
xor U7862 (N_7862,N_5208,N_3904);
xnor U7863 (N_7863,N_3480,N_5678);
nand U7864 (N_7864,N_4765,N_5400);
nand U7865 (N_7865,N_3562,N_5202);
nand U7866 (N_7866,N_4268,N_3676);
nor U7867 (N_7867,N_5661,N_4268);
or U7868 (N_7868,N_4033,N_4528);
or U7869 (N_7869,N_5156,N_5635);
xnor U7870 (N_7870,N_5250,N_4776);
nand U7871 (N_7871,N_3129,N_5991);
nand U7872 (N_7872,N_3763,N_3605);
or U7873 (N_7873,N_4991,N_5816);
nand U7874 (N_7874,N_4023,N_3080);
or U7875 (N_7875,N_5452,N_5622);
nand U7876 (N_7876,N_3281,N_5541);
nand U7877 (N_7877,N_5405,N_5602);
and U7878 (N_7878,N_5027,N_4185);
nand U7879 (N_7879,N_3075,N_5657);
and U7880 (N_7880,N_4574,N_4453);
or U7881 (N_7881,N_5025,N_4496);
nand U7882 (N_7882,N_5473,N_5369);
xnor U7883 (N_7883,N_3218,N_4053);
or U7884 (N_7884,N_5675,N_5340);
xnor U7885 (N_7885,N_5114,N_5737);
xor U7886 (N_7886,N_5388,N_4857);
xnor U7887 (N_7887,N_3194,N_4962);
nand U7888 (N_7888,N_4356,N_5863);
nor U7889 (N_7889,N_3619,N_5077);
nand U7890 (N_7890,N_3744,N_5965);
nand U7891 (N_7891,N_3803,N_5670);
or U7892 (N_7892,N_4362,N_4266);
or U7893 (N_7893,N_5205,N_3847);
xnor U7894 (N_7894,N_5585,N_3750);
nand U7895 (N_7895,N_4948,N_4536);
xor U7896 (N_7896,N_5574,N_5977);
nand U7897 (N_7897,N_5505,N_3946);
xnor U7898 (N_7898,N_4332,N_4581);
nand U7899 (N_7899,N_4794,N_3092);
nor U7900 (N_7900,N_5128,N_5647);
nand U7901 (N_7901,N_5324,N_5388);
nor U7902 (N_7902,N_4516,N_3763);
nand U7903 (N_7903,N_4663,N_3514);
xnor U7904 (N_7904,N_4214,N_4453);
nor U7905 (N_7905,N_3063,N_4759);
nand U7906 (N_7906,N_3747,N_5497);
or U7907 (N_7907,N_4495,N_4510);
and U7908 (N_7908,N_5633,N_3535);
xnor U7909 (N_7909,N_5034,N_5646);
and U7910 (N_7910,N_5741,N_4983);
nand U7911 (N_7911,N_3344,N_4759);
xor U7912 (N_7912,N_4428,N_5218);
and U7913 (N_7913,N_4597,N_5130);
nand U7914 (N_7914,N_4935,N_3982);
xor U7915 (N_7915,N_5598,N_3019);
and U7916 (N_7916,N_5058,N_3859);
and U7917 (N_7917,N_5444,N_3514);
nand U7918 (N_7918,N_5484,N_3083);
and U7919 (N_7919,N_3553,N_4050);
nand U7920 (N_7920,N_5677,N_4491);
or U7921 (N_7921,N_3292,N_4337);
or U7922 (N_7922,N_4067,N_5043);
xor U7923 (N_7923,N_3991,N_3453);
nand U7924 (N_7924,N_3941,N_5189);
or U7925 (N_7925,N_3328,N_5649);
nor U7926 (N_7926,N_3797,N_5936);
nor U7927 (N_7927,N_3229,N_4423);
xor U7928 (N_7928,N_5634,N_3129);
xor U7929 (N_7929,N_4232,N_3618);
nand U7930 (N_7930,N_4113,N_3017);
nor U7931 (N_7931,N_3858,N_3526);
xnor U7932 (N_7932,N_3604,N_5294);
nand U7933 (N_7933,N_4587,N_5249);
nand U7934 (N_7934,N_4889,N_3725);
or U7935 (N_7935,N_5509,N_3261);
xor U7936 (N_7936,N_4483,N_5758);
nor U7937 (N_7937,N_4094,N_5804);
xnor U7938 (N_7938,N_4627,N_3679);
or U7939 (N_7939,N_4677,N_3845);
nor U7940 (N_7940,N_3909,N_4266);
and U7941 (N_7941,N_5157,N_3670);
nor U7942 (N_7942,N_5235,N_3545);
or U7943 (N_7943,N_4322,N_3722);
nand U7944 (N_7944,N_3416,N_4340);
nor U7945 (N_7945,N_3275,N_4364);
xor U7946 (N_7946,N_3806,N_4084);
nor U7947 (N_7947,N_3592,N_5985);
nand U7948 (N_7948,N_3204,N_5629);
and U7949 (N_7949,N_5525,N_3658);
nor U7950 (N_7950,N_5792,N_3069);
xnor U7951 (N_7951,N_4297,N_4516);
xor U7952 (N_7952,N_4459,N_3116);
nand U7953 (N_7953,N_4864,N_5578);
and U7954 (N_7954,N_5052,N_4168);
nand U7955 (N_7955,N_4848,N_5224);
and U7956 (N_7956,N_5812,N_3106);
xnor U7957 (N_7957,N_4868,N_4687);
and U7958 (N_7958,N_5505,N_4046);
nor U7959 (N_7959,N_3669,N_3861);
and U7960 (N_7960,N_5647,N_3484);
nor U7961 (N_7961,N_4717,N_5262);
or U7962 (N_7962,N_5158,N_4941);
xor U7963 (N_7963,N_4944,N_3415);
nand U7964 (N_7964,N_3011,N_3017);
or U7965 (N_7965,N_3561,N_3220);
xnor U7966 (N_7966,N_4856,N_5253);
or U7967 (N_7967,N_5896,N_3921);
xor U7968 (N_7968,N_3705,N_4263);
nor U7969 (N_7969,N_3860,N_5436);
and U7970 (N_7970,N_5512,N_5200);
and U7971 (N_7971,N_3790,N_3217);
xor U7972 (N_7972,N_5718,N_5543);
and U7973 (N_7973,N_5757,N_5700);
xnor U7974 (N_7974,N_4433,N_3958);
nand U7975 (N_7975,N_5829,N_3311);
or U7976 (N_7976,N_4045,N_3463);
xnor U7977 (N_7977,N_5603,N_5077);
and U7978 (N_7978,N_4903,N_5820);
or U7979 (N_7979,N_3460,N_3090);
nand U7980 (N_7980,N_3059,N_5206);
or U7981 (N_7981,N_3169,N_3415);
and U7982 (N_7982,N_3316,N_4065);
nand U7983 (N_7983,N_5312,N_5164);
and U7984 (N_7984,N_5201,N_5724);
xor U7985 (N_7985,N_5380,N_5720);
nor U7986 (N_7986,N_3560,N_4295);
or U7987 (N_7987,N_4136,N_3787);
and U7988 (N_7988,N_5294,N_5581);
or U7989 (N_7989,N_3537,N_3229);
and U7990 (N_7990,N_5914,N_4303);
nor U7991 (N_7991,N_4733,N_3427);
xnor U7992 (N_7992,N_5863,N_5133);
nor U7993 (N_7993,N_4096,N_3071);
nor U7994 (N_7994,N_5457,N_3690);
nand U7995 (N_7995,N_3802,N_5841);
and U7996 (N_7996,N_5784,N_4995);
and U7997 (N_7997,N_3468,N_4813);
xnor U7998 (N_7998,N_5814,N_4688);
nand U7999 (N_7999,N_4931,N_5155);
and U8000 (N_8000,N_4205,N_5707);
nand U8001 (N_8001,N_4644,N_3122);
xnor U8002 (N_8002,N_5213,N_4996);
and U8003 (N_8003,N_5618,N_5501);
nand U8004 (N_8004,N_3431,N_3649);
nand U8005 (N_8005,N_3005,N_3666);
xnor U8006 (N_8006,N_3593,N_5967);
xnor U8007 (N_8007,N_3151,N_4454);
nand U8008 (N_8008,N_5106,N_4817);
nand U8009 (N_8009,N_5413,N_4564);
and U8010 (N_8010,N_3471,N_5490);
nor U8011 (N_8011,N_4874,N_4018);
nor U8012 (N_8012,N_3429,N_4474);
and U8013 (N_8013,N_4596,N_4165);
xor U8014 (N_8014,N_4455,N_4368);
and U8015 (N_8015,N_3252,N_5897);
or U8016 (N_8016,N_4482,N_3010);
and U8017 (N_8017,N_5741,N_5931);
nor U8018 (N_8018,N_4137,N_4986);
nand U8019 (N_8019,N_5937,N_5632);
nor U8020 (N_8020,N_4391,N_4059);
or U8021 (N_8021,N_4710,N_3738);
xnor U8022 (N_8022,N_3752,N_3309);
nand U8023 (N_8023,N_4380,N_3171);
nand U8024 (N_8024,N_3777,N_4701);
nand U8025 (N_8025,N_4186,N_4114);
and U8026 (N_8026,N_3890,N_3028);
xor U8027 (N_8027,N_4868,N_3700);
xor U8028 (N_8028,N_4157,N_3092);
nand U8029 (N_8029,N_4810,N_5371);
or U8030 (N_8030,N_3612,N_3021);
nor U8031 (N_8031,N_3783,N_4262);
nand U8032 (N_8032,N_5062,N_5377);
and U8033 (N_8033,N_5456,N_4489);
xnor U8034 (N_8034,N_5375,N_3768);
xnor U8035 (N_8035,N_4576,N_3795);
xnor U8036 (N_8036,N_3746,N_3315);
nand U8037 (N_8037,N_4265,N_4726);
nor U8038 (N_8038,N_4541,N_5825);
and U8039 (N_8039,N_4131,N_5666);
nand U8040 (N_8040,N_3297,N_3970);
xor U8041 (N_8041,N_4163,N_5768);
nand U8042 (N_8042,N_3128,N_4013);
or U8043 (N_8043,N_3184,N_4620);
or U8044 (N_8044,N_4256,N_5961);
nand U8045 (N_8045,N_3107,N_4701);
nand U8046 (N_8046,N_3898,N_3461);
and U8047 (N_8047,N_5408,N_4229);
nand U8048 (N_8048,N_5183,N_5447);
xnor U8049 (N_8049,N_4174,N_5797);
or U8050 (N_8050,N_3898,N_5972);
xor U8051 (N_8051,N_3424,N_5377);
xor U8052 (N_8052,N_4043,N_5601);
and U8053 (N_8053,N_4041,N_3537);
and U8054 (N_8054,N_5956,N_5495);
nand U8055 (N_8055,N_5264,N_3896);
and U8056 (N_8056,N_3867,N_4268);
nand U8057 (N_8057,N_5495,N_4334);
nand U8058 (N_8058,N_5657,N_4682);
or U8059 (N_8059,N_5463,N_4880);
xor U8060 (N_8060,N_5149,N_4418);
nor U8061 (N_8061,N_4496,N_3353);
nor U8062 (N_8062,N_5210,N_5657);
nand U8063 (N_8063,N_5721,N_5117);
and U8064 (N_8064,N_5399,N_3116);
and U8065 (N_8065,N_4296,N_3486);
nand U8066 (N_8066,N_5725,N_3478);
nor U8067 (N_8067,N_5220,N_3895);
or U8068 (N_8068,N_4681,N_4130);
nand U8069 (N_8069,N_4387,N_5304);
and U8070 (N_8070,N_4904,N_4738);
nand U8071 (N_8071,N_5539,N_4600);
nand U8072 (N_8072,N_4409,N_4222);
nor U8073 (N_8073,N_5805,N_5363);
nor U8074 (N_8074,N_4643,N_5786);
nor U8075 (N_8075,N_5715,N_3205);
or U8076 (N_8076,N_4158,N_4599);
nor U8077 (N_8077,N_4371,N_4564);
xnor U8078 (N_8078,N_5712,N_4550);
nand U8079 (N_8079,N_4524,N_5191);
or U8080 (N_8080,N_4802,N_4591);
nand U8081 (N_8081,N_3102,N_3658);
and U8082 (N_8082,N_5360,N_4567);
xnor U8083 (N_8083,N_5564,N_3009);
or U8084 (N_8084,N_5341,N_5445);
nand U8085 (N_8085,N_5254,N_4432);
nand U8086 (N_8086,N_5475,N_3650);
or U8087 (N_8087,N_3730,N_4779);
and U8088 (N_8088,N_3496,N_4666);
or U8089 (N_8089,N_3565,N_3210);
nand U8090 (N_8090,N_5757,N_4600);
xnor U8091 (N_8091,N_5960,N_3139);
or U8092 (N_8092,N_4305,N_5442);
nor U8093 (N_8093,N_5465,N_4628);
nand U8094 (N_8094,N_3576,N_5482);
xor U8095 (N_8095,N_5362,N_5069);
or U8096 (N_8096,N_5850,N_3022);
or U8097 (N_8097,N_4401,N_3959);
or U8098 (N_8098,N_3148,N_5294);
or U8099 (N_8099,N_3897,N_5032);
nor U8100 (N_8100,N_3115,N_3298);
nor U8101 (N_8101,N_4256,N_3939);
nand U8102 (N_8102,N_4935,N_5084);
or U8103 (N_8103,N_5522,N_4621);
or U8104 (N_8104,N_4590,N_4427);
xnor U8105 (N_8105,N_5466,N_3973);
or U8106 (N_8106,N_4762,N_4080);
nor U8107 (N_8107,N_3973,N_3974);
xor U8108 (N_8108,N_5533,N_5347);
xnor U8109 (N_8109,N_3584,N_5642);
xnor U8110 (N_8110,N_4848,N_4599);
or U8111 (N_8111,N_4043,N_5677);
nor U8112 (N_8112,N_4435,N_5078);
or U8113 (N_8113,N_5064,N_5386);
and U8114 (N_8114,N_4469,N_5536);
nor U8115 (N_8115,N_5811,N_5081);
xor U8116 (N_8116,N_5466,N_3808);
xor U8117 (N_8117,N_4970,N_5506);
nand U8118 (N_8118,N_4425,N_4504);
nand U8119 (N_8119,N_4389,N_3990);
xnor U8120 (N_8120,N_5518,N_5423);
and U8121 (N_8121,N_5263,N_4917);
nor U8122 (N_8122,N_5730,N_3771);
nor U8123 (N_8123,N_3714,N_5038);
xnor U8124 (N_8124,N_3495,N_5675);
or U8125 (N_8125,N_3762,N_5779);
or U8126 (N_8126,N_4196,N_5417);
nor U8127 (N_8127,N_5817,N_3202);
nand U8128 (N_8128,N_5121,N_3715);
nand U8129 (N_8129,N_3870,N_4494);
or U8130 (N_8130,N_5994,N_4773);
and U8131 (N_8131,N_3313,N_4975);
nor U8132 (N_8132,N_5411,N_3611);
nor U8133 (N_8133,N_5398,N_4324);
nand U8134 (N_8134,N_4078,N_3439);
nand U8135 (N_8135,N_4438,N_5163);
nand U8136 (N_8136,N_4844,N_3086);
nand U8137 (N_8137,N_4254,N_4631);
xor U8138 (N_8138,N_3536,N_5787);
nor U8139 (N_8139,N_4306,N_4871);
nand U8140 (N_8140,N_5379,N_5417);
or U8141 (N_8141,N_3727,N_5909);
or U8142 (N_8142,N_4366,N_5327);
or U8143 (N_8143,N_4372,N_4793);
xnor U8144 (N_8144,N_4450,N_4761);
and U8145 (N_8145,N_3497,N_3595);
or U8146 (N_8146,N_5208,N_5514);
nand U8147 (N_8147,N_5898,N_3544);
or U8148 (N_8148,N_3198,N_4771);
nand U8149 (N_8149,N_5520,N_4223);
nand U8150 (N_8150,N_4136,N_5008);
xor U8151 (N_8151,N_3052,N_3320);
or U8152 (N_8152,N_5586,N_5746);
and U8153 (N_8153,N_3189,N_3533);
nor U8154 (N_8154,N_3394,N_3651);
nand U8155 (N_8155,N_4874,N_3280);
nor U8156 (N_8156,N_5815,N_3109);
or U8157 (N_8157,N_3112,N_5311);
and U8158 (N_8158,N_3801,N_5025);
xnor U8159 (N_8159,N_5924,N_5132);
nor U8160 (N_8160,N_4245,N_5360);
and U8161 (N_8161,N_4743,N_4611);
nand U8162 (N_8162,N_4502,N_3810);
and U8163 (N_8163,N_3395,N_4968);
xor U8164 (N_8164,N_5048,N_4849);
nor U8165 (N_8165,N_5439,N_4319);
xnor U8166 (N_8166,N_4041,N_5345);
or U8167 (N_8167,N_3181,N_3903);
and U8168 (N_8168,N_5892,N_4637);
and U8169 (N_8169,N_4488,N_4911);
nand U8170 (N_8170,N_3427,N_4002);
or U8171 (N_8171,N_5221,N_5114);
and U8172 (N_8172,N_3275,N_4568);
or U8173 (N_8173,N_4431,N_4684);
xor U8174 (N_8174,N_3277,N_5024);
nor U8175 (N_8175,N_3695,N_3111);
nor U8176 (N_8176,N_3712,N_3099);
and U8177 (N_8177,N_4974,N_3148);
xor U8178 (N_8178,N_4010,N_3450);
xor U8179 (N_8179,N_4765,N_4352);
nand U8180 (N_8180,N_3986,N_3462);
nor U8181 (N_8181,N_5361,N_3073);
nand U8182 (N_8182,N_4614,N_5311);
and U8183 (N_8183,N_5345,N_3766);
or U8184 (N_8184,N_4547,N_5152);
nand U8185 (N_8185,N_4422,N_3616);
nor U8186 (N_8186,N_5048,N_3302);
or U8187 (N_8187,N_5128,N_5769);
or U8188 (N_8188,N_3741,N_3831);
and U8189 (N_8189,N_3138,N_5201);
and U8190 (N_8190,N_4907,N_5423);
nor U8191 (N_8191,N_4134,N_5815);
or U8192 (N_8192,N_5799,N_3839);
and U8193 (N_8193,N_4547,N_5847);
or U8194 (N_8194,N_4332,N_5316);
and U8195 (N_8195,N_3564,N_5611);
and U8196 (N_8196,N_4024,N_3680);
xnor U8197 (N_8197,N_5057,N_5583);
nor U8198 (N_8198,N_5348,N_3342);
nand U8199 (N_8199,N_3454,N_3461);
xor U8200 (N_8200,N_5975,N_5599);
xor U8201 (N_8201,N_3190,N_3573);
and U8202 (N_8202,N_4942,N_3948);
xor U8203 (N_8203,N_3035,N_3713);
nand U8204 (N_8204,N_4471,N_3554);
nand U8205 (N_8205,N_4220,N_3090);
nor U8206 (N_8206,N_3050,N_4877);
nand U8207 (N_8207,N_5456,N_5457);
and U8208 (N_8208,N_3022,N_3922);
or U8209 (N_8209,N_5732,N_4127);
or U8210 (N_8210,N_3444,N_5906);
nand U8211 (N_8211,N_5416,N_5932);
nand U8212 (N_8212,N_4598,N_3751);
nand U8213 (N_8213,N_5696,N_4132);
nand U8214 (N_8214,N_5243,N_3898);
or U8215 (N_8215,N_4053,N_3821);
nor U8216 (N_8216,N_4996,N_4547);
nand U8217 (N_8217,N_3219,N_4032);
nor U8218 (N_8218,N_5070,N_5962);
xor U8219 (N_8219,N_4779,N_3259);
or U8220 (N_8220,N_3728,N_4370);
nor U8221 (N_8221,N_5941,N_3116);
nand U8222 (N_8222,N_4422,N_5989);
and U8223 (N_8223,N_3828,N_5737);
xnor U8224 (N_8224,N_4853,N_3775);
xor U8225 (N_8225,N_5862,N_3526);
nor U8226 (N_8226,N_5319,N_4901);
xnor U8227 (N_8227,N_5427,N_5039);
xor U8228 (N_8228,N_5580,N_4579);
and U8229 (N_8229,N_5881,N_3988);
xnor U8230 (N_8230,N_3045,N_3307);
or U8231 (N_8231,N_4659,N_4309);
and U8232 (N_8232,N_3782,N_3663);
and U8233 (N_8233,N_4217,N_3324);
xnor U8234 (N_8234,N_5937,N_4647);
nor U8235 (N_8235,N_3041,N_3888);
or U8236 (N_8236,N_5939,N_3687);
nand U8237 (N_8237,N_4487,N_4375);
or U8238 (N_8238,N_4041,N_3219);
or U8239 (N_8239,N_4036,N_4225);
xnor U8240 (N_8240,N_4161,N_3539);
nor U8241 (N_8241,N_3261,N_4363);
or U8242 (N_8242,N_5703,N_4719);
xnor U8243 (N_8243,N_5104,N_4603);
and U8244 (N_8244,N_5967,N_4596);
nand U8245 (N_8245,N_5037,N_4585);
nand U8246 (N_8246,N_4436,N_5894);
or U8247 (N_8247,N_5155,N_4824);
nor U8248 (N_8248,N_3602,N_5576);
nand U8249 (N_8249,N_5473,N_3203);
nor U8250 (N_8250,N_3773,N_3747);
and U8251 (N_8251,N_3824,N_3698);
or U8252 (N_8252,N_5759,N_3870);
nand U8253 (N_8253,N_4812,N_5190);
nor U8254 (N_8254,N_3053,N_3221);
nor U8255 (N_8255,N_3251,N_3016);
xor U8256 (N_8256,N_5797,N_3331);
nand U8257 (N_8257,N_4068,N_4175);
and U8258 (N_8258,N_5947,N_3464);
or U8259 (N_8259,N_5719,N_4293);
xnor U8260 (N_8260,N_4733,N_4865);
xnor U8261 (N_8261,N_3347,N_5714);
and U8262 (N_8262,N_3209,N_5534);
nand U8263 (N_8263,N_3014,N_5054);
or U8264 (N_8264,N_4486,N_4236);
nand U8265 (N_8265,N_3067,N_3951);
nor U8266 (N_8266,N_4496,N_5919);
and U8267 (N_8267,N_5625,N_4938);
or U8268 (N_8268,N_4215,N_3829);
or U8269 (N_8269,N_4670,N_3562);
xnor U8270 (N_8270,N_4022,N_4395);
and U8271 (N_8271,N_4702,N_4794);
nor U8272 (N_8272,N_3637,N_5507);
and U8273 (N_8273,N_3559,N_5002);
xnor U8274 (N_8274,N_3995,N_4428);
and U8275 (N_8275,N_5851,N_5862);
and U8276 (N_8276,N_3931,N_3497);
and U8277 (N_8277,N_5809,N_4968);
nand U8278 (N_8278,N_5894,N_4158);
or U8279 (N_8279,N_3588,N_3177);
and U8280 (N_8280,N_4922,N_5921);
or U8281 (N_8281,N_4647,N_5855);
nor U8282 (N_8282,N_5344,N_5938);
nand U8283 (N_8283,N_3590,N_3485);
nand U8284 (N_8284,N_4516,N_4992);
xnor U8285 (N_8285,N_3239,N_3446);
nand U8286 (N_8286,N_3511,N_3473);
and U8287 (N_8287,N_4446,N_4143);
and U8288 (N_8288,N_5624,N_5854);
or U8289 (N_8289,N_5583,N_4115);
xor U8290 (N_8290,N_5600,N_3077);
xnor U8291 (N_8291,N_5419,N_4545);
or U8292 (N_8292,N_4514,N_3137);
nand U8293 (N_8293,N_3267,N_5177);
xor U8294 (N_8294,N_5627,N_3428);
nand U8295 (N_8295,N_4315,N_4932);
nand U8296 (N_8296,N_5501,N_5004);
xnor U8297 (N_8297,N_4047,N_4344);
nor U8298 (N_8298,N_5277,N_5358);
and U8299 (N_8299,N_3347,N_5908);
nor U8300 (N_8300,N_4595,N_5797);
nand U8301 (N_8301,N_5279,N_4242);
nand U8302 (N_8302,N_5955,N_4599);
or U8303 (N_8303,N_4140,N_5600);
nand U8304 (N_8304,N_5098,N_3126);
nor U8305 (N_8305,N_3123,N_4065);
and U8306 (N_8306,N_5961,N_5294);
and U8307 (N_8307,N_3387,N_4575);
or U8308 (N_8308,N_5580,N_5246);
or U8309 (N_8309,N_3191,N_4481);
nor U8310 (N_8310,N_4504,N_3210);
and U8311 (N_8311,N_3248,N_5689);
or U8312 (N_8312,N_4851,N_3982);
nand U8313 (N_8313,N_4866,N_3903);
or U8314 (N_8314,N_3034,N_4033);
xor U8315 (N_8315,N_4704,N_4226);
or U8316 (N_8316,N_5444,N_4867);
or U8317 (N_8317,N_5383,N_5005);
and U8318 (N_8318,N_3803,N_4484);
and U8319 (N_8319,N_3417,N_4524);
and U8320 (N_8320,N_4213,N_4086);
nand U8321 (N_8321,N_5009,N_3849);
or U8322 (N_8322,N_5690,N_4024);
and U8323 (N_8323,N_5629,N_3706);
xor U8324 (N_8324,N_5162,N_5781);
or U8325 (N_8325,N_3924,N_3206);
xor U8326 (N_8326,N_5630,N_5606);
or U8327 (N_8327,N_5197,N_5764);
nand U8328 (N_8328,N_3255,N_5763);
nand U8329 (N_8329,N_3403,N_3681);
or U8330 (N_8330,N_3914,N_5280);
nor U8331 (N_8331,N_4537,N_3342);
and U8332 (N_8332,N_5514,N_5199);
nand U8333 (N_8333,N_5748,N_5730);
xor U8334 (N_8334,N_5356,N_5665);
nand U8335 (N_8335,N_4447,N_4417);
xnor U8336 (N_8336,N_5046,N_5007);
or U8337 (N_8337,N_4864,N_5791);
or U8338 (N_8338,N_4994,N_3946);
nand U8339 (N_8339,N_4447,N_3202);
xor U8340 (N_8340,N_4808,N_5277);
and U8341 (N_8341,N_4523,N_4587);
and U8342 (N_8342,N_3898,N_5601);
and U8343 (N_8343,N_3106,N_3087);
xor U8344 (N_8344,N_3822,N_4622);
nor U8345 (N_8345,N_4512,N_3572);
and U8346 (N_8346,N_5268,N_4299);
xnor U8347 (N_8347,N_4213,N_3707);
nor U8348 (N_8348,N_4079,N_3005);
nor U8349 (N_8349,N_4766,N_5759);
nand U8350 (N_8350,N_5538,N_4145);
and U8351 (N_8351,N_3723,N_4651);
nand U8352 (N_8352,N_5677,N_3823);
nand U8353 (N_8353,N_3182,N_4908);
xnor U8354 (N_8354,N_4382,N_4426);
and U8355 (N_8355,N_5240,N_4899);
nor U8356 (N_8356,N_3192,N_5851);
xnor U8357 (N_8357,N_5374,N_4687);
xor U8358 (N_8358,N_3982,N_5818);
and U8359 (N_8359,N_3204,N_4465);
and U8360 (N_8360,N_3129,N_4109);
or U8361 (N_8361,N_3922,N_5601);
nand U8362 (N_8362,N_3041,N_3944);
and U8363 (N_8363,N_3672,N_3509);
and U8364 (N_8364,N_3235,N_5810);
nand U8365 (N_8365,N_4922,N_5649);
nand U8366 (N_8366,N_3498,N_3947);
nor U8367 (N_8367,N_5715,N_5138);
xor U8368 (N_8368,N_4779,N_3385);
nor U8369 (N_8369,N_5973,N_5119);
nand U8370 (N_8370,N_3339,N_4170);
and U8371 (N_8371,N_5675,N_3614);
nor U8372 (N_8372,N_4918,N_4183);
nand U8373 (N_8373,N_4158,N_4811);
and U8374 (N_8374,N_3080,N_3609);
and U8375 (N_8375,N_3611,N_4721);
nand U8376 (N_8376,N_4939,N_5990);
or U8377 (N_8377,N_3135,N_3961);
nor U8378 (N_8378,N_4862,N_3426);
nor U8379 (N_8379,N_3800,N_3555);
nand U8380 (N_8380,N_3432,N_3577);
nor U8381 (N_8381,N_4122,N_5111);
nand U8382 (N_8382,N_3225,N_4939);
xor U8383 (N_8383,N_3399,N_5472);
xnor U8384 (N_8384,N_3179,N_5581);
xnor U8385 (N_8385,N_5502,N_4219);
or U8386 (N_8386,N_5176,N_5419);
xnor U8387 (N_8387,N_3598,N_3090);
nand U8388 (N_8388,N_3061,N_4255);
and U8389 (N_8389,N_5619,N_3520);
or U8390 (N_8390,N_5242,N_3340);
and U8391 (N_8391,N_5548,N_5849);
xor U8392 (N_8392,N_4393,N_4218);
xnor U8393 (N_8393,N_4826,N_3643);
nand U8394 (N_8394,N_5641,N_4427);
nand U8395 (N_8395,N_5517,N_5943);
nand U8396 (N_8396,N_5844,N_4335);
and U8397 (N_8397,N_3813,N_3950);
nand U8398 (N_8398,N_4785,N_5316);
nor U8399 (N_8399,N_3095,N_4861);
xnor U8400 (N_8400,N_4711,N_4723);
and U8401 (N_8401,N_4151,N_4421);
nor U8402 (N_8402,N_4746,N_5301);
and U8403 (N_8403,N_5818,N_5696);
or U8404 (N_8404,N_4496,N_4925);
xnor U8405 (N_8405,N_5798,N_3855);
nor U8406 (N_8406,N_4287,N_4296);
and U8407 (N_8407,N_3215,N_4276);
nand U8408 (N_8408,N_3378,N_3230);
nand U8409 (N_8409,N_3813,N_5377);
xnor U8410 (N_8410,N_5048,N_4099);
xor U8411 (N_8411,N_4972,N_4305);
nand U8412 (N_8412,N_5983,N_4566);
nand U8413 (N_8413,N_4317,N_3318);
or U8414 (N_8414,N_5133,N_5506);
xor U8415 (N_8415,N_5174,N_3013);
and U8416 (N_8416,N_3356,N_4219);
nor U8417 (N_8417,N_3541,N_5863);
nor U8418 (N_8418,N_5332,N_3988);
nor U8419 (N_8419,N_3310,N_4928);
xor U8420 (N_8420,N_3869,N_3131);
nor U8421 (N_8421,N_5343,N_5498);
nand U8422 (N_8422,N_3770,N_3208);
xor U8423 (N_8423,N_5013,N_3491);
nand U8424 (N_8424,N_3150,N_4003);
and U8425 (N_8425,N_4357,N_5470);
or U8426 (N_8426,N_4171,N_5181);
xor U8427 (N_8427,N_3052,N_4325);
xnor U8428 (N_8428,N_3038,N_3430);
or U8429 (N_8429,N_5206,N_3900);
xor U8430 (N_8430,N_5684,N_3634);
and U8431 (N_8431,N_3724,N_5868);
or U8432 (N_8432,N_3241,N_5793);
xnor U8433 (N_8433,N_4404,N_4240);
nand U8434 (N_8434,N_5739,N_3784);
or U8435 (N_8435,N_4021,N_3605);
xor U8436 (N_8436,N_5390,N_4703);
nor U8437 (N_8437,N_4198,N_5511);
nand U8438 (N_8438,N_3407,N_4565);
nand U8439 (N_8439,N_3745,N_5149);
xnor U8440 (N_8440,N_5707,N_3950);
and U8441 (N_8441,N_3894,N_3615);
and U8442 (N_8442,N_3320,N_5624);
nor U8443 (N_8443,N_5806,N_4675);
xor U8444 (N_8444,N_4528,N_3069);
nand U8445 (N_8445,N_4735,N_3718);
and U8446 (N_8446,N_4504,N_4874);
and U8447 (N_8447,N_4975,N_4297);
nor U8448 (N_8448,N_4543,N_5498);
and U8449 (N_8449,N_3661,N_3053);
nor U8450 (N_8450,N_3107,N_4885);
nand U8451 (N_8451,N_3767,N_5508);
and U8452 (N_8452,N_4545,N_3616);
nor U8453 (N_8453,N_3913,N_3786);
or U8454 (N_8454,N_4606,N_3021);
xor U8455 (N_8455,N_3989,N_5748);
xnor U8456 (N_8456,N_5650,N_4528);
and U8457 (N_8457,N_3561,N_3091);
xnor U8458 (N_8458,N_3819,N_5705);
nor U8459 (N_8459,N_4748,N_3567);
and U8460 (N_8460,N_4174,N_4052);
nor U8461 (N_8461,N_4978,N_4069);
nor U8462 (N_8462,N_5434,N_3878);
nor U8463 (N_8463,N_5395,N_5756);
nor U8464 (N_8464,N_3615,N_3163);
or U8465 (N_8465,N_3190,N_3682);
nand U8466 (N_8466,N_3286,N_5920);
xor U8467 (N_8467,N_3386,N_4096);
nand U8468 (N_8468,N_4018,N_4396);
nor U8469 (N_8469,N_3984,N_3841);
nand U8470 (N_8470,N_5590,N_3976);
and U8471 (N_8471,N_4615,N_3277);
or U8472 (N_8472,N_4699,N_3170);
nor U8473 (N_8473,N_4639,N_3121);
nor U8474 (N_8474,N_5629,N_3237);
or U8475 (N_8475,N_5063,N_4066);
nand U8476 (N_8476,N_3124,N_4572);
and U8477 (N_8477,N_4468,N_3968);
nand U8478 (N_8478,N_5157,N_4666);
nand U8479 (N_8479,N_4418,N_3444);
and U8480 (N_8480,N_5106,N_3899);
nand U8481 (N_8481,N_4097,N_5552);
nor U8482 (N_8482,N_5851,N_4913);
nor U8483 (N_8483,N_5806,N_3498);
nand U8484 (N_8484,N_4340,N_4866);
xor U8485 (N_8485,N_5823,N_5461);
nand U8486 (N_8486,N_4894,N_3060);
or U8487 (N_8487,N_4323,N_4986);
nand U8488 (N_8488,N_4972,N_4491);
and U8489 (N_8489,N_5086,N_3622);
and U8490 (N_8490,N_3540,N_5261);
xor U8491 (N_8491,N_4072,N_4798);
nand U8492 (N_8492,N_4631,N_5665);
and U8493 (N_8493,N_3880,N_4582);
nor U8494 (N_8494,N_4603,N_5322);
nand U8495 (N_8495,N_3886,N_5775);
and U8496 (N_8496,N_5273,N_5582);
xnor U8497 (N_8497,N_5842,N_4847);
nand U8498 (N_8498,N_4109,N_4247);
xor U8499 (N_8499,N_5951,N_4889);
and U8500 (N_8500,N_5165,N_3210);
or U8501 (N_8501,N_4396,N_4887);
nand U8502 (N_8502,N_3415,N_5796);
xor U8503 (N_8503,N_5686,N_3351);
or U8504 (N_8504,N_4008,N_4782);
or U8505 (N_8505,N_5025,N_5321);
nor U8506 (N_8506,N_5659,N_3138);
nor U8507 (N_8507,N_5839,N_5816);
xnor U8508 (N_8508,N_5281,N_4494);
nand U8509 (N_8509,N_3965,N_3902);
and U8510 (N_8510,N_3350,N_3846);
xor U8511 (N_8511,N_3776,N_5682);
xnor U8512 (N_8512,N_4352,N_3095);
or U8513 (N_8513,N_5011,N_5528);
nor U8514 (N_8514,N_3447,N_5482);
nor U8515 (N_8515,N_3195,N_5230);
and U8516 (N_8516,N_5117,N_3204);
and U8517 (N_8517,N_4856,N_4904);
or U8518 (N_8518,N_5251,N_5790);
and U8519 (N_8519,N_5464,N_3357);
or U8520 (N_8520,N_3395,N_5657);
or U8521 (N_8521,N_5405,N_4374);
xor U8522 (N_8522,N_5463,N_3698);
and U8523 (N_8523,N_5837,N_3533);
and U8524 (N_8524,N_5782,N_5039);
or U8525 (N_8525,N_5651,N_3182);
and U8526 (N_8526,N_4847,N_3554);
nand U8527 (N_8527,N_4067,N_4737);
nor U8528 (N_8528,N_5183,N_5025);
and U8529 (N_8529,N_5819,N_5109);
or U8530 (N_8530,N_3175,N_4456);
nand U8531 (N_8531,N_3055,N_5667);
or U8532 (N_8532,N_5384,N_4962);
xnor U8533 (N_8533,N_5664,N_4642);
nor U8534 (N_8534,N_4496,N_4339);
nand U8535 (N_8535,N_5207,N_4221);
and U8536 (N_8536,N_3731,N_4564);
xnor U8537 (N_8537,N_3729,N_3395);
xnor U8538 (N_8538,N_5411,N_4549);
or U8539 (N_8539,N_5159,N_4905);
nor U8540 (N_8540,N_5366,N_3429);
xor U8541 (N_8541,N_4651,N_4996);
and U8542 (N_8542,N_4096,N_5556);
xor U8543 (N_8543,N_3109,N_3696);
nand U8544 (N_8544,N_5987,N_4692);
nand U8545 (N_8545,N_5018,N_4608);
nor U8546 (N_8546,N_4478,N_5517);
or U8547 (N_8547,N_5830,N_4589);
nand U8548 (N_8548,N_4317,N_3465);
and U8549 (N_8549,N_4489,N_5643);
nor U8550 (N_8550,N_4239,N_3772);
or U8551 (N_8551,N_3032,N_3238);
nor U8552 (N_8552,N_3780,N_3300);
or U8553 (N_8553,N_5030,N_5390);
or U8554 (N_8554,N_5607,N_5903);
and U8555 (N_8555,N_4238,N_3709);
and U8556 (N_8556,N_5839,N_5536);
nor U8557 (N_8557,N_4190,N_3051);
or U8558 (N_8558,N_4329,N_5644);
nand U8559 (N_8559,N_3675,N_3550);
or U8560 (N_8560,N_3743,N_5886);
and U8561 (N_8561,N_5543,N_4408);
or U8562 (N_8562,N_4436,N_3445);
xor U8563 (N_8563,N_5726,N_5013);
nand U8564 (N_8564,N_3234,N_3620);
xor U8565 (N_8565,N_4352,N_3379);
or U8566 (N_8566,N_4280,N_3265);
nor U8567 (N_8567,N_4608,N_4303);
xnor U8568 (N_8568,N_5079,N_3689);
nor U8569 (N_8569,N_3099,N_3543);
and U8570 (N_8570,N_5173,N_3011);
or U8571 (N_8571,N_3926,N_3355);
xnor U8572 (N_8572,N_5335,N_3122);
or U8573 (N_8573,N_5804,N_5391);
or U8574 (N_8574,N_5662,N_5703);
nor U8575 (N_8575,N_3340,N_5265);
or U8576 (N_8576,N_5791,N_3193);
or U8577 (N_8577,N_3560,N_5060);
nand U8578 (N_8578,N_4709,N_5841);
nand U8579 (N_8579,N_5474,N_5788);
nor U8580 (N_8580,N_3624,N_3295);
and U8581 (N_8581,N_4680,N_3324);
nand U8582 (N_8582,N_4713,N_3022);
nand U8583 (N_8583,N_5371,N_4821);
or U8584 (N_8584,N_4677,N_3596);
xnor U8585 (N_8585,N_3526,N_4047);
or U8586 (N_8586,N_3575,N_5499);
nor U8587 (N_8587,N_5750,N_4464);
nand U8588 (N_8588,N_5397,N_5894);
nand U8589 (N_8589,N_3011,N_5331);
and U8590 (N_8590,N_5305,N_3206);
and U8591 (N_8591,N_3499,N_4706);
xor U8592 (N_8592,N_4946,N_3411);
nand U8593 (N_8593,N_5316,N_3609);
or U8594 (N_8594,N_4881,N_4068);
nor U8595 (N_8595,N_4950,N_3893);
nor U8596 (N_8596,N_5017,N_4129);
xor U8597 (N_8597,N_3650,N_3599);
nor U8598 (N_8598,N_5514,N_5866);
nor U8599 (N_8599,N_5022,N_4186);
nand U8600 (N_8600,N_3644,N_4086);
or U8601 (N_8601,N_5700,N_5655);
nand U8602 (N_8602,N_5139,N_5107);
xor U8603 (N_8603,N_5731,N_4004);
and U8604 (N_8604,N_4839,N_4962);
or U8605 (N_8605,N_4016,N_5072);
and U8606 (N_8606,N_5814,N_4362);
xnor U8607 (N_8607,N_5164,N_3722);
and U8608 (N_8608,N_4466,N_4198);
nand U8609 (N_8609,N_4859,N_3285);
and U8610 (N_8610,N_4242,N_4644);
or U8611 (N_8611,N_5335,N_4757);
and U8612 (N_8612,N_5048,N_5356);
nor U8613 (N_8613,N_4520,N_4094);
xor U8614 (N_8614,N_4070,N_5160);
or U8615 (N_8615,N_3408,N_5793);
xor U8616 (N_8616,N_3636,N_4153);
or U8617 (N_8617,N_5375,N_4544);
and U8618 (N_8618,N_5446,N_5673);
and U8619 (N_8619,N_5347,N_3235);
nor U8620 (N_8620,N_4732,N_3145);
and U8621 (N_8621,N_3003,N_3462);
and U8622 (N_8622,N_3686,N_5991);
nand U8623 (N_8623,N_4947,N_4425);
nand U8624 (N_8624,N_3274,N_5037);
or U8625 (N_8625,N_5348,N_5812);
or U8626 (N_8626,N_5339,N_3386);
or U8627 (N_8627,N_3478,N_4113);
nor U8628 (N_8628,N_3854,N_4209);
and U8629 (N_8629,N_4326,N_3041);
or U8630 (N_8630,N_5705,N_5471);
or U8631 (N_8631,N_3878,N_4989);
xnor U8632 (N_8632,N_4947,N_3567);
nand U8633 (N_8633,N_4631,N_3634);
and U8634 (N_8634,N_4963,N_3655);
nor U8635 (N_8635,N_3876,N_5983);
nand U8636 (N_8636,N_4069,N_4384);
and U8637 (N_8637,N_5866,N_4524);
or U8638 (N_8638,N_5813,N_4136);
and U8639 (N_8639,N_3866,N_3180);
nand U8640 (N_8640,N_3840,N_5938);
nor U8641 (N_8641,N_3137,N_5406);
nor U8642 (N_8642,N_3380,N_4503);
nand U8643 (N_8643,N_5064,N_4095);
nor U8644 (N_8644,N_5260,N_5569);
nor U8645 (N_8645,N_3572,N_5638);
xor U8646 (N_8646,N_5020,N_3449);
xnor U8647 (N_8647,N_5759,N_3503);
nor U8648 (N_8648,N_5856,N_5098);
xor U8649 (N_8649,N_4255,N_4068);
xor U8650 (N_8650,N_5103,N_4490);
nand U8651 (N_8651,N_4668,N_3532);
nor U8652 (N_8652,N_3901,N_4054);
nand U8653 (N_8653,N_4087,N_3653);
nand U8654 (N_8654,N_3521,N_4672);
nor U8655 (N_8655,N_3812,N_5173);
nor U8656 (N_8656,N_4059,N_3241);
and U8657 (N_8657,N_3520,N_4110);
or U8658 (N_8658,N_3135,N_4915);
and U8659 (N_8659,N_3990,N_4643);
or U8660 (N_8660,N_5586,N_3856);
xnor U8661 (N_8661,N_5490,N_4427);
and U8662 (N_8662,N_5752,N_4704);
or U8663 (N_8663,N_3318,N_5419);
or U8664 (N_8664,N_4142,N_4786);
nor U8665 (N_8665,N_3290,N_3144);
and U8666 (N_8666,N_5704,N_3577);
or U8667 (N_8667,N_3601,N_3087);
nor U8668 (N_8668,N_5880,N_5227);
or U8669 (N_8669,N_5479,N_3765);
nand U8670 (N_8670,N_3609,N_5069);
nor U8671 (N_8671,N_3993,N_5693);
nand U8672 (N_8672,N_5650,N_3209);
and U8673 (N_8673,N_3687,N_4038);
nand U8674 (N_8674,N_5929,N_4961);
xnor U8675 (N_8675,N_4649,N_4458);
nand U8676 (N_8676,N_3974,N_4984);
xor U8677 (N_8677,N_4260,N_5226);
or U8678 (N_8678,N_3337,N_3956);
or U8679 (N_8679,N_3117,N_3965);
xnor U8680 (N_8680,N_3913,N_3623);
or U8681 (N_8681,N_4924,N_3704);
nor U8682 (N_8682,N_4343,N_3014);
and U8683 (N_8683,N_4102,N_5228);
and U8684 (N_8684,N_5114,N_4656);
and U8685 (N_8685,N_5640,N_3390);
nand U8686 (N_8686,N_4818,N_5399);
nand U8687 (N_8687,N_5381,N_3252);
nand U8688 (N_8688,N_4703,N_5611);
xor U8689 (N_8689,N_4023,N_5903);
and U8690 (N_8690,N_3460,N_4756);
and U8691 (N_8691,N_5490,N_4143);
nand U8692 (N_8692,N_5163,N_4913);
nand U8693 (N_8693,N_4730,N_5141);
and U8694 (N_8694,N_4516,N_3510);
or U8695 (N_8695,N_5445,N_5549);
or U8696 (N_8696,N_4838,N_5292);
or U8697 (N_8697,N_5019,N_3526);
nand U8698 (N_8698,N_4380,N_4548);
xnor U8699 (N_8699,N_4063,N_5126);
or U8700 (N_8700,N_4668,N_5707);
and U8701 (N_8701,N_4902,N_5226);
or U8702 (N_8702,N_4695,N_3497);
nor U8703 (N_8703,N_5802,N_4961);
nand U8704 (N_8704,N_4821,N_3141);
and U8705 (N_8705,N_3968,N_5744);
nor U8706 (N_8706,N_3872,N_4866);
xnor U8707 (N_8707,N_5060,N_4513);
nand U8708 (N_8708,N_4208,N_5069);
and U8709 (N_8709,N_5705,N_4517);
and U8710 (N_8710,N_5181,N_3517);
nand U8711 (N_8711,N_4760,N_4723);
nand U8712 (N_8712,N_4513,N_3380);
or U8713 (N_8713,N_3970,N_3383);
nand U8714 (N_8714,N_4214,N_5254);
and U8715 (N_8715,N_5382,N_5320);
nor U8716 (N_8716,N_3203,N_4692);
xnor U8717 (N_8717,N_3895,N_3781);
and U8718 (N_8718,N_3763,N_5935);
nor U8719 (N_8719,N_3311,N_3540);
nor U8720 (N_8720,N_3810,N_3683);
xor U8721 (N_8721,N_3267,N_4118);
nor U8722 (N_8722,N_5614,N_5733);
and U8723 (N_8723,N_3200,N_3638);
and U8724 (N_8724,N_3322,N_5933);
xor U8725 (N_8725,N_5263,N_5815);
xor U8726 (N_8726,N_5239,N_5306);
nor U8727 (N_8727,N_5348,N_3433);
and U8728 (N_8728,N_4736,N_3063);
and U8729 (N_8729,N_4413,N_3564);
and U8730 (N_8730,N_5247,N_4619);
or U8731 (N_8731,N_3440,N_4836);
xor U8732 (N_8732,N_5627,N_3879);
and U8733 (N_8733,N_5569,N_3925);
xnor U8734 (N_8734,N_4793,N_5653);
or U8735 (N_8735,N_4031,N_5513);
or U8736 (N_8736,N_5099,N_4024);
nand U8737 (N_8737,N_3779,N_3417);
or U8738 (N_8738,N_4637,N_4641);
nand U8739 (N_8739,N_4478,N_3072);
and U8740 (N_8740,N_4642,N_5378);
or U8741 (N_8741,N_3063,N_4582);
nor U8742 (N_8742,N_3568,N_5836);
xor U8743 (N_8743,N_3385,N_4283);
and U8744 (N_8744,N_5553,N_3323);
and U8745 (N_8745,N_4723,N_5936);
nand U8746 (N_8746,N_4707,N_3695);
or U8747 (N_8747,N_4724,N_4678);
and U8748 (N_8748,N_4927,N_3880);
nor U8749 (N_8749,N_4434,N_4207);
xor U8750 (N_8750,N_4156,N_4043);
nand U8751 (N_8751,N_4567,N_5162);
and U8752 (N_8752,N_5335,N_3045);
or U8753 (N_8753,N_3119,N_4258);
xnor U8754 (N_8754,N_4217,N_4156);
and U8755 (N_8755,N_3761,N_3832);
nor U8756 (N_8756,N_4947,N_5752);
nand U8757 (N_8757,N_4866,N_5827);
nand U8758 (N_8758,N_5306,N_3926);
nor U8759 (N_8759,N_4483,N_3874);
and U8760 (N_8760,N_4116,N_5555);
xor U8761 (N_8761,N_3425,N_3629);
or U8762 (N_8762,N_4472,N_3140);
and U8763 (N_8763,N_5847,N_4533);
and U8764 (N_8764,N_3992,N_3071);
and U8765 (N_8765,N_4205,N_5303);
nor U8766 (N_8766,N_3690,N_5753);
or U8767 (N_8767,N_3676,N_5720);
nor U8768 (N_8768,N_5842,N_5097);
nor U8769 (N_8769,N_4161,N_5023);
and U8770 (N_8770,N_5402,N_5111);
and U8771 (N_8771,N_4221,N_3914);
or U8772 (N_8772,N_3663,N_4977);
and U8773 (N_8773,N_5568,N_5110);
or U8774 (N_8774,N_3827,N_5808);
nand U8775 (N_8775,N_5261,N_5579);
nand U8776 (N_8776,N_5531,N_4546);
and U8777 (N_8777,N_4170,N_4101);
xnor U8778 (N_8778,N_3860,N_5144);
and U8779 (N_8779,N_4406,N_3766);
nand U8780 (N_8780,N_5856,N_4018);
or U8781 (N_8781,N_3170,N_4661);
nand U8782 (N_8782,N_4940,N_3284);
nand U8783 (N_8783,N_3711,N_4851);
nand U8784 (N_8784,N_3125,N_5533);
xnor U8785 (N_8785,N_4666,N_3605);
xnor U8786 (N_8786,N_4147,N_5437);
nand U8787 (N_8787,N_5041,N_4884);
nand U8788 (N_8788,N_3688,N_3611);
xor U8789 (N_8789,N_5869,N_5827);
nand U8790 (N_8790,N_4110,N_3799);
and U8791 (N_8791,N_4596,N_3033);
or U8792 (N_8792,N_3641,N_5170);
or U8793 (N_8793,N_3169,N_3667);
and U8794 (N_8794,N_3997,N_3296);
xnor U8795 (N_8795,N_4589,N_5608);
or U8796 (N_8796,N_5142,N_5691);
or U8797 (N_8797,N_5384,N_5029);
nor U8798 (N_8798,N_3252,N_3879);
nand U8799 (N_8799,N_4009,N_3800);
nand U8800 (N_8800,N_5253,N_3815);
or U8801 (N_8801,N_3190,N_5202);
nand U8802 (N_8802,N_5954,N_3291);
and U8803 (N_8803,N_3717,N_4271);
nand U8804 (N_8804,N_5501,N_4614);
and U8805 (N_8805,N_5505,N_3968);
nand U8806 (N_8806,N_4876,N_4655);
xnor U8807 (N_8807,N_3590,N_3689);
xnor U8808 (N_8808,N_5960,N_5636);
and U8809 (N_8809,N_4530,N_5015);
xnor U8810 (N_8810,N_4801,N_4365);
or U8811 (N_8811,N_3266,N_5945);
and U8812 (N_8812,N_5505,N_4996);
xnor U8813 (N_8813,N_5899,N_5201);
and U8814 (N_8814,N_4868,N_4376);
nand U8815 (N_8815,N_4778,N_5066);
nor U8816 (N_8816,N_5363,N_4892);
nand U8817 (N_8817,N_3835,N_5724);
xor U8818 (N_8818,N_4061,N_4681);
and U8819 (N_8819,N_4516,N_4956);
or U8820 (N_8820,N_5042,N_3775);
xor U8821 (N_8821,N_4468,N_3722);
nor U8822 (N_8822,N_3815,N_4858);
and U8823 (N_8823,N_3933,N_4721);
and U8824 (N_8824,N_5331,N_5132);
or U8825 (N_8825,N_3943,N_4536);
or U8826 (N_8826,N_3062,N_3346);
xor U8827 (N_8827,N_3569,N_3041);
nor U8828 (N_8828,N_5085,N_3731);
or U8829 (N_8829,N_4482,N_3339);
nand U8830 (N_8830,N_4213,N_5164);
xnor U8831 (N_8831,N_3419,N_3215);
nor U8832 (N_8832,N_3801,N_5689);
nor U8833 (N_8833,N_4589,N_4339);
nor U8834 (N_8834,N_3237,N_3319);
nor U8835 (N_8835,N_4892,N_4182);
nor U8836 (N_8836,N_3885,N_3298);
nor U8837 (N_8837,N_5185,N_4289);
nor U8838 (N_8838,N_5201,N_4240);
or U8839 (N_8839,N_4264,N_4083);
nand U8840 (N_8840,N_5815,N_4358);
xnor U8841 (N_8841,N_3428,N_5721);
and U8842 (N_8842,N_5401,N_5365);
or U8843 (N_8843,N_5989,N_5004);
and U8844 (N_8844,N_3717,N_5598);
nor U8845 (N_8845,N_3736,N_5642);
nor U8846 (N_8846,N_5694,N_5525);
or U8847 (N_8847,N_3375,N_3582);
xor U8848 (N_8848,N_3955,N_3061);
xnor U8849 (N_8849,N_5107,N_4458);
xnor U8850 (N_8850,N_3175,N_3331);
or U8851 (N_8851,N_3064,N_5804);
and U8852 (N_8852,N_4929,N_3611);
xor U8853 (N_8853,N_5740,N_4373);
nand U8854 (N_8854,N_3087,N_3757);
nand U8855 (N_8855,N_4473,N_4356);
or U8856 (N_8856,N_3010,N_5467);
or U8857 (N_8857,N_4216,N_5481);
and U8858 (N_8858,N_4529,N_3423);
and U8859 (N_8859,N_3188,N_4088);
and U8860 (N_8860,N_5646,N_5121);
and U8861 (N_8861,N_3338,N_5866);
nor U8862 (N_8862,N_5465,N_3480);
and U8863 (N_8863,N_3641,N_3659);
nand U8864 (N_8864,N_4319,N_4701);
xnor U8865 (N_8865,N_4975,N_5070);
nand U8866 (N_8866,N_4548,N_3305);
or U8867 (N_8867,N_4924,N_3400);
and U8868 (N_8868,N_5492,N_3957);
or U8869 (N_8869,N_5401,N_3294);
or U8870 (N_8870,N_3689,N_5033);
or U8871 (N_8871,N_5953,N_4857);
and U8872 (N_8872,N_3765,N_4749);
xor U8873 (N_8873,N_3680,N_5895);
nand U8874 (N_8874,N_5352,N_3740);
nor U8875 (N_8875,N_4555,N_5134);
and U8876 (N_8876,N_5920,N_5712);
and U8877 (N_8877,N_3052,N_5635);
and U8878 (N_8878,N_5769,N_3138);
nor U8879 (N_8879,N_4298,N_4013);
nand U8880 (N_8880,N_4481,N_3126);
and U8881 (N_8881,N_5653,N_5524);
and U8882 (N_8882,N_5632,N_3168);
and U8883 (N_8883,N_3620,N_5099);
and U8884 (N_8884,N_5127,N_4193);
or U8885 (N_8885,N_3187,N_5974);
and U8886 (N_8886,N_4055,N_5623);
nor U8887 (N_8887,N_4237,N_4386);
nor U8888 (N_8888,N_5259,N_5998);
nor U8889 (N_8889,N_5203,N_4691);
nor U8890 (N_8890,N_4004,N_4097);
or U8891 (N_8891,N_3873,N_4104);
xnor U8892 (N_8892,N_5246,N_3105);
nand U8893 (N_8893,N_4926,N_4037);
nand U8894 (N_8894,N_4363,N_4841);
nor U8895 (N_8895,N_4225,N_3474);
nor U8896 (N_8896,N_3499,N_4543);
and U8897 (N_8897,N_4684,N_3976);
or U8898 (N_8898,N_4334,N_3144);
nand U8899 (N_8899,N_3302,N_3889);
nor U8900 (N_8900,N_4260,N_4479);
nor U8901 (N_8901,N_5536,N_4087);
nand U8902 (N_8902,N_3790,N_5381);
nand U8903 (N_8903,N_4440,N_3160);
xnor U8904 (N_8904,N_5220,N_3106);
and U8905 (N_8905,N_5342,N_5830);
and U8906 (N_8906,N_5200,N_5020);
nor U8907 (N_8907,N_3717,N_4148);
and U8908 (N_8908,N_4140,N_3473);
nand U8909 (N_8909,N_3857,N_3237);
and U8910 (N_8910,N_4905,N_3110);
nand U8911 (N_8911,N_4814,N_5090);
nand U8912 (N_8912,N_4644,N_3601);
and U8913 (N_8913,N_3024,N_5113);
or U8914 (N_8914,N_3548,N_3703);
nor U8915 (N_8915,N_5319,N_3668);
or U8916 (N_8916,N_4909,N_5313);
or U8917 (N_8917,N_5035,N_3759);
or U8918 (N_8918,N_3737,N_4597);
nor U8919 (N_8919,N_4916,N_5038);
and U8920 (N_8920,N_5196,N_4849);
or U8921 (N_8921,N_3107,N_4904);
xnor U8922 (N_8922,N_3014,N_5661);
xor U8923 (N_8923,N_5887,N_4888);
xnor U8924 (N_8924,N_4516,N_5108);
nor U8925 (N_8925,N_3728,N_3401);
or U8926 (N_8926,N_4089,N_4330);
or U8927 (N_8927,N_5407,N_4775);
nand U8928 (N_8928,N_5099,N_5602);
or U8929 (N_8929,N_4211,N_5484);
and U8930 (N_8930,N_5405,N_3430);
and U8931 (N_8931,N_3933,N_4853);
nor U8932 (N_8932,N_5932,N_5044);
nor U8933 (N_8933,N_3515,N_4374);
nor U8934 (N_8934,N_5508,N_5100);
nor U8935 (N_8935,N_4057,N_3698);
and U8936 (N_8936,N_5210,N_3087);
nand U8937 (N_8937,N_3973,N_4196);
nand U8938 (N_8938,N_5838,N_4110);
nand U8939 (N_8939,N_3161,N_5313);
or U8940 (N_8940,N_5087,N_4378);
nor U8941 (N_8941,N_5823,N_4273);
and U8942 (N_8942,N_5208,N_5651);
nor U8943 (N_8943,N_3136,N_5957);
xnor U8944 (N_8944,N_4572,N_5954);
or U8945 (N_8945,N_3560,N_3527);
nor U8946 (N_8946,N_5069,N_5746);
nand U8947 (N_8947,N_3195,N_3380);
nand U8948 (N_8948,N_5012,N_3890);
nand U8949 (N_8949,N_5831,N_5569);
nand U8950 (N_8950,N_4934,N_3595);
and U8951 (N_8951,N_3847,N_3348);
xor U8952 (N_8952,N_4059,N_3840);
nand U8953 (N_8953,N_4833,N_4486);
xnor U8954 (N_8954,N_4517,N_5883);
xnor U8955 (N_8955,N_5872,N_3881);
or U8956 (N_8956,N_5261,N_4230);
nand U8957 (N_8957,N_5934,N_5817);
and U8958 (N_8958,N_4817,N_3470);
nor U8959 (N_8959,N_4453,N_4173);
and U8960 (N_8960,N_5173,N_5210);
nor U8961 (N_8961,N_3453,N_3365);
and U8962 (N_8962,N_3446,N_5821);
nand U8963 (N_8963,N_5953,N_4050);
or U8964 (N_8964,N_3680,N_4663);
nor U8965 (N_8965,N_5475,N_4438);
nand U8966 (N_8966,N_3070,N_3986);
nand U8967 (N_8967,N_5083,N_4401);
xnor U8968 (N_8968,N_5243,N_5088);
or U8969 (N_8969,N_3749,N_5427);
and U8970 (N_8970,N_5868,N_3810);
nor U8971 (N_8971,N_5072,N_4416);
nand U8972 (N_8972,N_3064,N_4095);
nor U8973 (N_8973,N_4635,N_4357);
nand U8974 (N_8974,N_4865,N_5031);
or U8975 (N_8975,N_3195,N_3052);
nand U8976 (N_8976,N_3743,N_5008);
and U8977 (N_8977,N_4205,N_4486);
xor U8978 (N_8978,N_5035,N_4182);
xnor U8979 (N_8979,N_3554,N_3349);
and U8980 (N_8980,N_4032,N_4015);
xor U8981 (N_8981,N_5296,N_4280);
nand U8982 (N_8982,N_4903,N_3152);
nand U8983 (N_8983,N_5795,N_5192);
nor U8984 (N_8984,N_3152,N_5809);
nor U8985 (N_8985,N_3604,N_3121);
or U8986 (N_8986,N_4532,N_3666);
or U8987 (N_8987,N_4231,N_5079);
xnor U8988 (N_8988,N_4499,N_5037);
and U8989 (N_8989,N_5807,N_5121);
nor U8990 (N_8990,N_4406,N_4883);
nor U8991 (N_8991,N_4053,N_3976);
nand U8992 (N_8992,N_5131,N_5511);
xor U8993 (N_8993,N_4634,N_4247);
xnor U8994 (N_8994,N_3541,N_4269);
or U8995 (N_8995,N_3550,N_4442);
xnor U8996 (N_8996,N_4400,N_4687);
nand U8997 (N_8997,N_5492,N_3300);
or U8998 (N_8998,N_4489,N_4778);
or U8999 (N_8999,N_3628,N_3318);
nand U9000 (N_9000,N_8267,N_7191);
nor U9001 (N_9001,N_7667,N_6275);
or U9002 (N_9002,N_7578,N_7937);
xnor U9003 (N_9003,N_8755,N_8505);
or U9004 (N_9004,N_6126,N_8557);
xor U9005 (N_9005,N_8279,N_8462);
nor U9006 (N_9006,N_6884,N_7832);
or U9007 (N_9007,N_8926,N_7278);
xnor U9008 (N_9008,N_8789,N_6585);
or U9009 (N_9009,N_7375,N_7285);
or U9010 (N_9010,N_8753,N_7416);
nand U9011 (N_9011,N_8830,N_8009);
xor U9012 (N_9012,N_8216,N_6639);
xor U9013 (N_9013,N_6453,N_6533);
nor U9014 (N_9014,N_7779,N_6317);
xor U9015 (N_9015,N_7855,N_7603);
xnor U9016 (N_9016,N_7351,N_6158);
or U9017 (N_9017,N_8787,N_7188);
nor U9018 (N_9018,N_6672,N_8726);
nand U9019 (N_9019,N_8620,N_7004);
xor U9020 (N_9020,N_6113,N_7982);
and U9021 (N_9021,N_7055,N_8366);
nor U9022 (N_9022,N_8409,N_8183);
nand U9023 (N_9023,N_6490,N_7861);
and U9024 (N_9024,N_8232,N_6274);
nand U9025 (N_9025,N_7638,N_8011);
or U9026 (N_9026,N_8206,N_8786);
nor U9027 (N_9027,N_7296,N_6277);
or U9028 (N_9028,N_7294,N_8800);
or U9029 (N_9029,N_6579,N_8284);
nor U9030 (N_9030,N_6219,N_8698);
or U9031 (N_9031,N_6504,N_6100);
and U9032 (N_9032,N_8508,N_7678);
nor U9033 (N_9033,N_7321,N_7629);
nor U9034 (N_9034,N_7595,N_7984);
nand U9035 (N_9035,N_6048,N_7061);
xnor U9036 (N_9036,N_8594,N_6228);
and U9037 (N_9037,N_8548,N_6649);
and U9038 (N_9038,N_7017,N_7802);
or U9039 (N_9039,N_6843,N_7356);
nand U9040 (N_9040,N_6471,N_7269);
nand U9041 (N_9041,N_6499,N_7340);
or U9042 (N_9042,N_6399,N_8130);
xnor U9043 (N_9043,N_7640,N_7027);
nor U9044 (N_9044,N_8427,N_6208);
nand U9045 (N_9045,N_7085,N_6822);
xor U9046 (N_9046,N_8129,N_7838);
nand U9047 (N_9047,N_7227,N_7486);
and U9048 (N_9048,N_6663,N_6510);
and U9049 (N_9049,N_7087,N_7734);
nor U9050 (N_9050,N_8408,N_8715);
nand U9051 (N_9051,N_8320,N_6160);
xor U9052 (N_9052,N_8621,N_6409);
or U9053 (N_9053,N_6134,N_7525);
xnor U9054 (N_9054,N_8092,N_8720);
xnor U9055 (N_9055,N_8870,N_8920);
and U9056 (N_9056,N_8510,N_8116);
nand U9057 (N_9057,N_8939,N_6526);
and U9058 (N_9058,N_7012,N_6738);
or U9059 (N_9059,N_8649,N_7418);
nand U9060 (N_9060,N_8230,N_8072);
and U9061 (N_9061,N_7909,N_7325);
nor U9062 (N_9062,N_7063,N_8218);
and U9063 (N_9063,N_7409,N_7954);
and U9064 (N_9064,N_8874,N_7005);
and U9065 (N_9065,N_6241,N_8217);
and U9066 (N_9066,N_8541,N_8815);
or U9067 (N_9067,N_6169,N_8764);
nor U9068 (N_9068,N_6632,N_6748);
or U9069 (N_9069,N_8795,N_6683);
xnor U9070 (N_9070,N_7350,N_8781);
or U9071 (N_9071,N_6175,N_6335);
nand U9072 (N_9072,N_8039,N_6302);
nor U9073 (N_9073,N_6911,N_6763);
or U9074 (N_9074,N_6596,N_8543);
nand U9075 (N_9075,N_6790,N_6122);
nand U9076 (N_9076,N_7167,N_6456);
nor U9077 (N_9077,N_7470,N_8724);
or U9078 (N_9078,N_7495,N_6703);
and U9079 (N_9079,N_6569,N_7746);
xnor U9080 (N_9080,N_8937,N_7732);
nor U9081 (N_9081,N_6700,N_7198);
or U9082 (N_9082,N_8438,N_7283);
and U9083 (N_9083,N_7704,N_8604);
or U9084 (N_9084,N_6411,N_8154);
xnor U9085 (N_9085,N_7083,N_8925);
or U9086 (N_9086,N_7711,N_6272);
xnor U9087 (N_9087,N_7592,N_7308);
and U9088 (N_9088,N_8455,N_8606);
or U9089 (N_9089,N_8812,N_8576);
and U9090 (N_9090,N_6873,N_8322);
nor U9091 (N_9091,N_8746,N_7482);
and U9092 (N_9092,N_6167,N_8856);
nor U9093 (N_9093,N_6052,N_6657);
or U9094 (N_9094,N_6008,N_8282);
xor U9095 (N_9095,N_8226,N_7385);
xnor U9096 (N_9096,N_8674,N_8212);
or U9097 (N_9097,N_6245,N_6749);
or U9098 (N_9098,N_7302,N_8325);
nand U9099 (N_9099,N_6772,N_7933);
or U9100 (N_9100,N_8632,N_6170);
or U9101 (N_9101,N_7096,N_7155);
and U9102 (N_9102,N_6146,N_8763);
xnor U9103 (N_9103,N_6566,N_8450);
nor U9104 (N_9104,N_7100,N_8445);
nand U9105 (N_9105,N_7123,N_8440);
nor U9106 (N_9106,N_7290,N_6321);
and U9107 (N_9107,N_6328,N_7488);
nor U9108 (N_9108,N_6732,N_8535);
nand U9109 (N_9109,N_7652,N_7972);
and U9110 (N_9110,N_7122,N_8103);
xnor U9111 (N_9111,N_6652,N_6375);
nor U9112 (N_9112,N_6037,N_7837);
nor U9113 (N_9113,N_8090,N_8121);
and U9114 (N_9114,N_7970,N_7111);
and U9115 (N_9115,N_8064,N_8690);
xor U9116 (N_9116,N_6725,N_8495);
or U9117 (N_9117,N_6083,N_7701);
xor U9118 (N_9118,N_8754,N_6412);
nand U9119 (N_9119,N_6868,N_7723);
nand U9120 (N_9120,N_7360,N_8909);
and U9121 (N_9121,N_7673,N_6580);
or U9122 (N_9122,N_7508,N_7580);
nor U9123 (N_9123,N_6060,N_6252);
and U9124 (N_9124,N_7435,N_8101);
and U9125 (N_9125,N_8118,N_8189);
xor U9126 (N_9126,N_6007,N_7824);
and U9127 (N_9127,N_6091,N_8307);
xnor U9128 (N_9128,N_8741,N_6929);
and U9129 (N_9129,N_7995,N_7774);
and U9130 (N_9130,N_7963,N_6559);
nor U9131 (N_9131,N_7020,N_7880);
nor U9132 (N_9132,N_8935,N_8014);
nor U9133 (N_9133,N_7266,N_7778);
nor U9134 (N_9134,N_7414,N_6390);
xor U9135 (N_9135,N_8147,N_8528);
xor U9136 (N_9136,N_8058,N_8210);
nor U9137 (N_9137,N_7519,N_7811);
nand U9138 (N_9138,N_8310,N_7310);
or U9139 (N_9139,N_8953,N_8088);
xor U9140 (N_9140,N_6305,N_7843);
or U9141 (N_9141,N_6650,N_6680);
nor U9142 (N_9142,N_6855,N_6201);
nor U9143 (N_9143,N_6183,N_6262);
nand U9144 (N_9144,N_7057,N_8613);
nand U9145 (N_9145,N_6155,N_7788);
nand U9146 (N_9146,N_8948,N_8544);
and U9147 (N_9147,N_8791,N_6668);
or U9148 (N_9148,N_7393,N_6845);
and U9149 (N_9149,N_7270,N_6147);
and U9150 (N_9150,N_8280,N_8405);
and U9151 (N_9151,N_6898,N_7165);
and U9152 (N_9152,N_6070,N_8418);
xnor U9153 (N_9153,N_6200,N_6303);
or U9154 (N_9154,N_6666,N_8084);
nand U9155 (N_9155,N_8105,N_7234);
or U9156 (N_9156,N_7612,N_6917);
and U9157 (N_9157,N_7383,N_6629);
xor U9158 (N_9158,N_6300,N_8941);
or U9159 (N_9159,N_8384,N_6432);
nor U9160 (N_9160,N_6350,N_7815);
nand U9161 (N_9161,N_7530,N_8809);
xnor U9162 (N_9162,N_8394,N_6662);
nand U9163 (N_9163,N_7468,N_8509);
and U9164 (N_9164,N_6475,N_6689);
nand U9165 (N_9165,N_7339,N_6821);
xor U9166 (N_9166,N_8037,N_8917);
and U9167 (N_9167,N_7960,N_8298);
nand U9168 (N_9168,N_6963,N_8444);
nand U9169 (N_9169,N_7413,N_6835);
nor U9170 (N_9170,N_6435,N_7421);
nor U9171 (N_9171,N_7658,N_8404);
or U9172 (N_9172,N_7107,N_7765);
and U9173 (N_9173,N_8711,N_6485);
xor U9174 (N_9174,N_7244,N_8550);
or U9175 (N_9175,N_6742,N_7596);
nor U9176 (N_9176,N_6227,N_8890);
nor U9177 (N_9177,N_7943,N_7881);
nand U9178 (N_9178,N_7259,N_6178);
nand U9179 (N_9179,N_6442,N_6144);
or U9180 (N_9180,N_7196,N_6391);
nand U9181 (N_9181,N_7023,N_8814);
xnor U9182 (N_9182,N_6810,N_8411);
xor U9183 (N_9183,N_8157,N_6258);
xor U9184 (N_9184,N_8646,N_6473);
nand U9185 (N_9185,N_8400,N_7391);
nor U9186 (N_9186,N_8113,N_6907);
or U9187 (N_9187,N_8179,N_6500);
nand U9188 (N_9188,N_7523,N_8045);
or U9189 (N_9189,N_6577,N_7280);
and U9190 (N_9190,N_6451,N_8916);
xnor U9191 (N_9191,N_7030,N_8422);
and U9192 (N_9192,N_7573,N_8251);
nand U9193 (N_9193,N_8231,N_8554);
nor U9194 (N_9194,N_7535,N_8790);
or U9195 (N_9195,N_8610,N_7128);
or U9196 (N_9196,N_6679,N_7715);
xor U9197 (N_9197,N_8355,N_6189);
nand U9198 (N_9198,N_8352,N_6468);
or U9199 (N_9199,N_6004,N_8608);
nand U9200 (N_9200,N_6910,N_6329);
nand U9201 (N_9201,N_7211,N_8175);
and U9202 (N_9202,N_7910,N_6033);
or U9203 (N_9203,N_6362,N_6728);
nor U9204 (N_9204,N_6179,N_6108);
or U9205 (N_9205,N_6168,N_7352);
xnor U9206 (N_9206,N_8016,N_7999);
or U9207 (N_9207,N_6531,N_6247);
nand U9208 (N_9208,N_6610,N_8335);
xnor U9209 (N_9209,N_6229,N_7170);
or U9210 (N_9210,N_7867,N_8759);
nor U9211 (N_9211,N_8693,N_7941);
nand U9212 (N_9212,N_8696,N_6349);
nor U9213 (N_9213,N_6202,N_8382);
and U9214 (N_9214,N_6207,N_7237);
nor U9215 (N_9215,N_7642,N_6752);
and U9216 (N_9216,N_8719,N_8141);
and U9217 (N_9217,N_8197,N_6781);
and U9218 (N_9218,N_7844,N_7347);
nand U9219 (N_9219,N_7448,N_7721);
nor U9220 (N_9220,N_8027,N_6393);
and U9221 (N_9221,N_8370,N_8805);
or U9222 (N_9222,N_7923,N_6906);
nand U9223 (N_9223,N_6421,N_6308);
or U9224 (N_9224,N_7876,N_7314);
xnor U9225 (N_9225,N_8365,N_6664);
xnor U9226 (N_9226,N_8599,N_8070);
or U9227 (N_9227,N_6159,N_7572);
and U9228 (N_9228,N_8131,N_7141);
and U9229 (N_9229,N_8447,N_8254);
xor U9230 (N_9230,N_7719,N_8562);
xnor U9231 (N_9231,N_8299,N_6494);
or U9232 (N_9232,N_8975,N_6978);
or U9233 (N_9233,N_8880,N_6373);
or U9234 (N_9234,N_7359,N_6086);
and U9235 (N_9235,N_8982,N_8669);
nor U9236 (N_9236,N_7420,N_6537);
xor U9237 (N_9237,N_8428,N_7432);
xnor U9238 (N_9238,N_8264,N_6894);
nand U9239 (N_9239,N_8517,N_8415);
and U9240 (N_9240,N_6582,N_6149);
nand U9241 (N_9241,N_7341,N_8785);
nand U9242 (N_9242,N_7307,N_6745);
and U9243 (N_9243,N_8395,N_8466);
and U9244 (N_9244,N_8356,N_7805);
or U9245 (N_9245,N_6065,N_8188);
or U9246 (N_9246,N_7126,N_7461);
or U9247 (N_9247,N_8593,N_6676);
xnor U9248 (N_9248,N_7473,N_6787);
nor U9249 (N_9249,N_8653,N_7865);
nor U9250 (N_9250,N_8957,N_7755);
xnor U9251 (N_9251,N_6476,N_6866);
or U9252 (N_9252,N_7725,N_6394);
nor U9253 (N_9253,N_6470,N_8624);
or U9254 (N_9254,N_8293,N_7478);
or U9255 (N_9255,N_8792,N_7134);
or U9256 (N_9256,N_7870,N_6392);
nand U9257 (N_9257,N_7474,N_8677);
and U9258 (N_9258,N_8031,N_7836);
xnor U9259 (N_9259,N_6982,N_6459);
nor U9260 (N_9260,N_6353,N_8729);
nor U9261 (N_9261,N_6243,N_8924);
and U9262 (N_9262,N_8184,N_8161);
and U9263 (N_9263,N_8582,N_6304);
and U9264 (N_9264,N_7090,N_8500);
nor U9265 (N_9265,N_6560,N_7953);
nand U9266 (N_9266,N_7009,N_8895);
xnor U9267 (N_9267,N_6628,N_6248);
nand U9268 (N_9268,N_8623,N_6572);
or U9269 (N_9269,N_6831,N_6933);
or U9270 (N_9270,N_7145,N_7271);
nor U9271 (N_9271,N_6647,N_8087);
or U9272 (N_9272,N_6828,N_7444);
nand U9273 (N_9273,N_8364,N_8017);
nor U9274 (N_9274,N_6592,N_8659);
or U9275 (N_9275,N_8170,N_8727);
nand U9276 (N_9276,N_8196,N_7586);
xnor U9277 (N_9277,N_8859,N_7037);
xor U9278 (N_9278,N_6612,N_6968);
nor U9279 (N_9279,N_6590,N_8964);
xor U9280 (N_9280,N_6646,N_8174);
or U9281 (N_9281,N_8481,N_8581);
or U9282 (N_9282,N_6705,N_8884);
nor U9283 (N_9283,N_6055,N_7641);
or U9284 (N_9284,N_8507,N_7967);
or U9285 (N_9285,N_6151,N_6690);
nor U9286 (N_9286,N_8200,N_7274);
nand U9287 (N_9287,N_6836,N_7785);
xor U9288 (N_9288,N_6753,N_6889);
nor U9289 (N_9289,N_7769,N_7924);
and U9290 (N_9290,N_6547,N_7276);
nor U9291 (N_9291,N_7557,N_8695);
nor U9292 (N_9292,N_6961,N_7829);
nor U9293 (N_9293,N_6669,N_7847);
nor U9294 (N_9294,N_8896,N_8263);
and U9295 (N_9295,N_8052,N_6237);
nor U9296 (N_9296,N_8579,N_8342);
or U9297 (N_9297,N_7770,N_8272);
nand U9298 (N_9298,N_8756,N_8803);
and U9299 (N_9299,N_8533,N_8337);
and U9300 (N_9300,N_8849,N_7029);
or U9301 (N_9301,N_6452,N_6403);
nor U9302 (N_9302,N_6895,N_6408);
and U9303 (N_9303,N_7898,N_7944);
xnor U9304 (N_9304,N_7514,N_6789);
xnor U9305 (N_9305,N_6257,N_6769);
or U9306 (N_9306,N_8449,N_8819);
nor U9307 (N_9307,N_7007,N_6900);
nand U9308 (N_9308,N_7616,N_7354);
nand U9309 (N_9309,N_6722,N_7506);
xor U9310 (N_9310,N_8373,N_8585);
or U9311 (N_9311,N_7043,N_7192);
or U9312 (N_9312,N_8420,N_7707);
xnor U9313 (N_9313,N_7254,N_8845);
nand U9314 (N_9314,N_8910,N_7477);
nand U9315 (N_9315,N_7694,N_8357);
nand U9316 (N_9316,N_7498,N_6901);
nand U9317 (N_9317,N_7938,N_6838);
or U9318 (N_9318,N_8228,N_8246);
nand U9319 (N_9319,N_6486,N_7058);
xnor U9320 (N_9320,N_8708,N_8467);
and U9321 (N_9321,N_6278,N_8234);
and U9322 (N_9322,N_8810,N_6865);
nand U9323 (N_9323,N_6716,N_6182);
or U9324 (N_9324,N_8032,N_8306);
xor U9325 (N_9325,N_6434,N_8497);
and U9326 (N_9326,N_8514,N_6054);
or U9327 (N_9327,N_7273,N_8164);
nor U9328 (N_9328,N_6603,N_7659);
nand U9329 (N_9329,N_8911,N_6484);
xor U9330 (N_9330,N_7547,N_8458);
nor U9331 (N_9331,N_8801,N_8402);
or U9332 (N_9332,N_6503,N_7367);
or U9333 (N_9333,N_7753,N_6892);
and U9334 (N_9334,N_8124,N_6024);
nor U9335 (N_9335,N_7232,N_6595);
xor U9336 (N_9336,N_7239,N_6334);
xnor U9337 (N_9337,N_6636,N_6808);
and U9338 (N_9338,N_7405,N_7670);
nand U9339 (N_9339,N_8704,N_8343);
xor U9340 (N_9340,N_7781,N_7284);
or U9341 (N_9341,N_7159,N_7842);
and U9342 (N_9342,N_6957,N_7998);
nor U9343 (N_9343,N_6852,N_7233);
and U9344 (N_9344,N_6496,N_7577);
and U9345 (N_9345,N_6110,N_8861);
or U9346 (N_9346,N_8275,N_7873);
nor U9347 (N_9347,N_8662,N_7863);
nand U9348 (N_9348,N_8133,N_7289);
and U9349 (N_9349,N_8046,N_6851);
nand U9350 (N_9350,N_7761,N_6544);
xor U9351 (N_9351,N_8679,N_6265);
nor U9352 (N_9352,N_6326,N_6543);
nand U9353 (N_9353,N_7118,N_7460);
and U9354 (N_9354,N_7248,N_8048);
xor U9355 (N_9355,N_8705,N_8877);
nor U9356 (N_9356,N_6023,N_6564);
nand U9357 (N_9357,N_8793,N_6932);
or U9358 (N_9358,N_7471,N_6163);
nand U9359 (N_9359,N_6527,N_6800);
nand U9360 (N_9360,N_7653,N_7793);
or U9361 (N_9361,N_7241,N_6859);
nor U9362 (N_9362,N_8634,N_6803);
or U9363 (N_9363,N_7113,N_7666);
xor U9364 (N_9364,N_8778,N_7258);
or U9365 (N_9365,N_6574,N_7373);
nand U9366 (N_9366,N_7336,N_8540);
nand U9367 (N_9367,N_8999,N_8607);
nand U9368 (N_9368,N_8112,N_7971);
or U9369 (N_9369,N_8765,N_8327);
or U9370 (N_9370,N_7546,N_7148);
and U9371 (N_9371,N_7487,N_8914);
nor U9372 (N_9372,N_6990,N_8068);
nand U9373 (N_9373,N_6358,N_7539);
or U9374 (N_9374,N_6436,N_7651);
nor U9375 (N_9375,N_6594,N_7019);
or U9376 (N_9376,N_7509,N_8127);
or U9377 (N_9377,N_8635,N_7455);
xor U9378 (N_9378,N_6867,N_6491);
xnor U9379 (N_9379,N_8168,N_7160);
xnor U9380 (N_9380,N_8779,N_6637);
xor U9381 (N_9381,N_7630,N_7220);
xnor U9382 (N_9382,N_8177,N_7047);
nand U9383 (N_9383,N_8903,N_6254);
nor U9384 (N_9384,N_8598,N_8201);
or U9385 (N_9385,N_7689,N_6264);
nand U9386 (N_9386,N_8551,N_6809);
nand U9387 (N_9387,N_7099,N_6427);
or U9388 (N_9388,N_7064,N_6114);
nor U9389 (N_9389,N_6715,N_7550);
nand U9390 (N_9390,N_6726,N_8005);
nand U9391 (N_9391,N_7194,N_7883);
nand U9392 (N_9392,N_6864,N_7527);
or U9393 (N_9393,N_6215,N_7635);
and U9394 (N_9394,N_8843,N_6806);
and U9395 (N_9395,N_7091,N_6986);
nor U9396 (N_9396,N_8923,N_8813);
or U9397 (N_9397,N_8056,N_6717);
nor U9398 (N_9398,N_7363,N_7562);
or U9399 (N_9399,N_8030,N_8996);
and U9400 (N_9400,N_8181,N_8530);
nor U9401 (N_9401,N_7402,N_8691);
nand U9402 (N_9402,N_8612,N_6407);
xnor U9403 (N_9403,N_8430,N_8371);
nand U9404 (N_9404,N_8463,N_7025);
or U9405 (N_9405,N_6554,N_7764);
xnor U9406 (N_9406,N_6947,N_7442);
and U9407 (N_9407,N_7928,N_8997);
nor U9408 (N_9408,N_7252,N_6665);
nor U9409 (N_9409,N_6764,N_8149);
nand U9410 (N_9410,N_6627,N_6509);
nor U9411 (N_9411,N_7889,N_6641);
or U9412 (N_9412,N_6562,N_6697);
or U9413 (N_9413,N_6567,N_8292);
and U9414 (N_9414,N_8943,N_6840);
nor U9415 (N_9415,N_7623,N_6222);
or U9416 (N_9416,N_6481,N_8361);
nand U9417 (N_9417,N_7001,N_6401);
nand U9418 (N_9418,N_8252,N_7959);
nor U9419 (N_9419,N_6903,N_8380);
or U9420 (N_9420,N_7922,N_7784);
nor U9421 (N_9421,N_6991,N_7812);
or U9422 (N_9422,N_8678,N_8652);
nor U9423 (N_9423,N_6285,N_7911);
and U9424 (N_9424,N_7210,N_7655);
and U9425 (N_9425,N_8000,N_8140);
and U9426 (N_9426,N_8297,N_6972);
xnor U9427 (N_9427,N_7245,N_8762);
xnor U9428 (N_9428,N_6288,N_8584);
nand U9429 (N_9429,N_6369,N_7696);
xor U9430 (N_9430,N_7268,N_7318);
and U9431 (N_9431,N_7767,N_6619);
and U9432 (N_9432,N_7445,N_6042);
and U9433 (N_9433,N_8477,N_7965);
and U9434 (N_9434,N_8879,N_8436);
xnor U9435 (N_9435,N_8419,N_6330);
nand U9436 (N_9436,N_7300,N_8243);
xor U9437 (N_9437,N_7263,N_7319);
nand U9438 (N_9438,N_7900,N_7361);
xor U9439 (N_9439,N_7879,N_8172);
xor U9440 (N_9440,N_6681,N_8050);
and U9441 (N_9441,N_6995,N_7071);
nand U9442 (N_9442,N_8132,N_8296);
nor U9443 (N_9443,N_6755,N_7895);
nand U9444 (N_9444,N_8207,N_8213);
and U9445 (N_9445,N_7695,N_7317);
nor U9446 (N_9446,N_6458,N_7443);
nand U9447 (N_9447,N_6255,N_6143);
or U9448 (N_9448,N_8004,N_8714);
or U9449 (N_9449,N_8564,N_6234);
xnor U9450 (N_9450,N_8622,N_7993);
and U9451 (N_9451,N_7371,N_8578);
nand U9452 (N_9452,N_6363,N_6936);
or U9453 (N_9453,N_6754,N_8358);
xor U9454 (N_9454,N_7479,N_7627);
or U9455 (N_9455,N_8558,N_6919);
or U9456 (N_9456,N_6534,N_8381);
and U9457 (N_9457,N_6487,N_6332);
nor U9458 (N_9458,N_7874,N_7989);
xnor U9459 (N_9459,N_8303,N_7127);
or U9460 (N_9460,N_7932,N_7262);
xor U9461 (N_9461,N_6480,N_8474);
nor U9462 (N_9462,N_7181,N_6224);
or U9463 (N_9463,N_6736,N_7758);
and U9464 (N_9464,N_7125,N_8223);
and U9465 (N_9465,N_8142,N_8651);
nor U9466 (N_9466,N_8918,N_6983);
and U9467 (N_9467,N_7594,N_7968);
nand U9468 (N_9468,N_6863,N_7979);
and U9469 (N_9469,N_7554,N_8503);
nor U9470 (N_9470,N_7489,N_6677);
and U9471 (N_9471,N_6940,N_8618);
and U9472 (N_9472,N_7894,N_8725);
or U9473 (N_9473,N_8748,N_7353);
and U9474 (N_9474,N_7890,N_6857);
and U9475 (N_9475,N_7175,N_8976);
and U9476 (N_9476,N_6814,N_6309);
xnor U9477 (N_9477,N_7287,N_7888);
and U9478 (N_9478,N_7992,N_8962);
xor U9479 (N_9479,N_8194,N_7311);
xnor U9480 (N_9480,N_8826,N_7337);
nand U9481 (N_9481,N_8836,N_6012);
nand U9482 (N_9482,N_8966,N_8950);
xor U9483 (N_9483,N_7948,N_8109);
or U9484 (N_9484,N_8960,N_8097);
xor U9485 (N_9485,N_8848,N_8972);
nand U9486 (N_9486,N_6626,N_7102);
or U9487 (N_9487,N_7093,N_7808);
nand U9488 (N_9488,N_8348,N_6552);
nor U9489 (N_9489,N_6172,N_6871);
xor U9490 (N_9490,N_7295,N_8323);
nand U9491 (N_9491,N_8774,N_8947);
and U9492 (N_9492,N_6320,N_6276);
xor U9493 (N_9493,N_7583,N_7293);
nand U9494 (N_9494,N_6775,N_6960);
nand U9495 (N_9495,N_7345,N_6440);
xnor U9496 (N_9496,N_6085,N_8930);
or U9497 (N_9497,N_8592,N_8702);
or U9498 (N_9498,N_7885,N_8012);
nor U9499 (N_9499,N_8270,N_7332);
and U9500 (N_9500,N_8432,N_6331);
and U9501 (N_9501,N_8833,N_8434);
and U9502 (N_9502,N_7201,N_7738);
nand U9503 (N_9503,N_6315,N_6997);
nand U9504 (N_9504,N_7522,N_7281);
xor U9505 (N_9505,N_7384,N_6779);
nor U9506 (N_9506,N_6294,N_8736);
or U9507 (N_9507,N_7497,N_6128);
xnor U9508 (N_9508,N_8522,N_7313);
xor U9509 (N_9509,N_7124,N_7576);
nand U9510 (N_9510,N_8688,N_6181);
nand U9511 (N_9511,N_8008,N_8208);
xor U9512 (N_9512,N_8028,N_6951);
and U9513 (N_9513,N_8406,N_8491);
or U9514 (N_9514,N_6020,N_7282);
and U9515 (N_9515,N_7400,N_7112);
or U9516 (N_9516,N_8931,N_7597);
or U9517 (N_9517,N_8616,N_8998);
xor U9518 (N_9518,N_7077,N_8586);
and U9519 (N_9519,N_6102,N_8399);
and U9520 (N_9520,N_8531,N_7291);
or U9521 (N_9521,N_7224,N_8086);
nand U9522 (N_9522,N_6774,N_6364);
xor U9523 (N_9523,N_7925,N_6206);
or U9524 (N_9524,N_7657,N_7412);
and U9525 (N_9525,N_7173,N_8077);
nor U9526 (N_9526,N_8734,N_8227);
xnor U9527 (N_9527,N_7830,N_8229);
nand U9528 (N_9528,N_6106,N_8818);
or U9529 (N_9529,N_8002,N_7875);
and U9530 (N_9530,N_8363,N_6782);
nor U9531 (N_9531,N_7026,N_6777);
nor U9532 (N_9532,N_7505,N_7260);
nor U9533 (N_9533,N_7121,N_6720);
or U9534 (N_9534,N_8098,N_8166);
and U9535 (N_9535,N_7864,N_7563);
xor U9536 (N_9536,N_8831,N_6946);
xor U9537 (N_9537,N_6778,N_7054);
nand U9538 (N_9538,N_6162,N_8331);
xnor U9539 (N_9539,N_6077,N_7759);
nor U9540 (N_9540,N_8967,N_7411);
xnor U9541 (N_9541,N_7048,N_8628);
xnor U9542 (N_9542,N_8281,N_8534);
xor U9543 (N_9543,N_7078,N_8431);
nand U9544 (N_9544,N_7074,N_6702);
nand U9545 (N_9545,N_7022,N_7073);
nand U9546 (N_9546,N_8311,N_7364);
and U9547 (N_9547,N_8772,N_6058);
xor U9548 (N_9548,N_7344,N_8283);
or U9549 (N_9549,N_6123,N_6545);
nand U9550 (N_9550,N_8882,N_6727);
and U9551 (N_9551,N_8044,N_6949);
xor U9552 (N_9552,N_8013,N_6075);
nand U9553 (N_9553,N_8955,N_8609);
nor U9554 (N_9554,N_8523,N_8317);
or U9555 (N_9555,N_8460,N_7771);
and U9556 (N_9556,N_6188,N_6423);
nor U9557 (N_9557,N_8784,N_7240);
nand U9558 (N_9558,N_7499,N_7534);
and U9559 (N_9559,N_6850,N_6140);
xor U9560 (N_9560,N_8214,N_7831);
and U9561 (N_9561,N_7382,N_6519);
nor U9562 (N_9562,N_8588,N_8487);
or U9563 (N_9563,N_6830,N_8858);
xor U9564 (N_9564,N_7335,N_8965);
nand U9565 (N_9565,N_7731,N_7069);
xnor U9566 (N_9566,N_8205,N_7430);
and U9567 (N_9567,N_6578,N_7555);
nand U9568 (N_9568,N_8421,N_7951);
nor U9569 (N_9569,N_6575,N_7153);
xnor U9570 (N_9570,N_6418,N_7171);
nor U9571 (N_9571,N_6266,N_6097);
xor U9572 (N_9572,N_7604,N_7397);
nand U9573 (N_9573,N_7206,N_7164);
xnor U9574 (N_9574,N_8872,N_8590);
or U9575 (N_9575,N_8290,N_8316);
xor U9576 (N_9576,N_7915,N_6542);
or U9577 (N_9577,N_8825,N_7343);
nand U9578 (N_9578,N_8658,N_6081);
xor U9579 (N_9579,N_7510,N_6263);
nor U9580 (N_9580,N_6682,N_6489);
and U9581 (N_9581,N_6756,N_8457);
xor U9582 (N_9582,N_6121,N_7135);
nor U9583 (N_9583,N_6483,N_7439);
and U9584 (N_9584,N_8577,N_8318);
nor U9585 (N_9585,N_6221,N_6952);
nand U9586 (N_9586,N_7656,N_6801);
nand U9587 (N_9587,N_8692,N_6209);
nor U9588 (N_9588,N_6751,N_7469);
or U9589 (N_9589,N_8111,N_7726);
or U9590 (N_9590,N_7685,N_7699);
nand U9591 (N_9591,N_8766,N_8739);
nor U9592 (N_9592,N_7620,N_8666);
or U9593 (N_9593,N_6540,N_6620);
nand U9594 (N_9594,N_8685,N_6909);
nand U9595 (N_9595,N_6372,N_8171);
nor U9596 (N_9596,N_6029,N_7503);
and U9597 (N_9597,N_6584,N_7480);
xor U9598 (N_9598,N_8993,N_8398);
nand U9599 (N_9599,N_7092,N_6343);
or U9600 (N_9600,N_7417,N_8767);
or U9601 (N_9601,N_6671,N_8108);
or U9602 (N_9602,N_6290,N_7028);
nor U9603 (N_9603,N_7182,N_6239);
or U9604 (N_9604,N_8878,N_6057);
nand U9605 (N_9605,N_7401,N_8153);
or U9606 (N_9606,N_6888,N_7306);
and U9607 (N_9607,N_8821,N_6558);
nand U9608 (N_9608,N_6444,N_7905);
xor U9609 (N_9609,N_7365,N_8047);
xor U9610 (N_9610,N_7143,N_8126);
nand U9611 (N_9611,N_6402,N_7654);
or U9612 (N_9612,N_7301,N_7710);
nor U9613 (N_9613,N_8580,N_8940);
nor U9614 (N_9614,N_8407,N_7187);
xor U9615 (N_9615,N_6109,N_7613);
nor U9616 (N_9616,N_6886,N_8029);
and U9617 (N_9617,N_6735,N_6299);
nand U9618 (N_9618,N_7109,N_6338);
and U9619 (N_9619,N_8003,N_7016);
nor U9620 (N_9620,N_6015,N_6478);
xnor U9621 (N_9621,N_7637,N_7045);
xnor U9622 (N_9622,N_7377,N_7209);
and U9623 (N_9623,N_7833,N_8829);
xnor U9624 (N_9624,N_7609,N_7940);
nor U9625 (N_9625,N_7800,N_6638);
xor U9626 (N_9626,N_7856,N_7702);
nand U9627 (N_9627,N_7436,N_7406);
xor U9628 (N_9628,N_8069,N_6931);
xnor U9629 (N_9629,N_7366,N_8783);
and U9630 (N_9630,N_8682,N_6529);
xor U9631 (N_9631,N_6443,N_8392);
xor U9632 (N_9632,N_7893,N_8922);
nor U9633 (N_9633,N_7010,N_6858);
xor U9634 (N_9634,N_7762,N_8148);
and U9635 (N_9635,N_6994,N_6236);
nor U9636 (N_9636,N_7231,N_6005);
nor U9637 (N_9637,N_6462,N_6516);
or U9638 (N_9638,N_6670,N_8209);
and U9639 (N_9639,N_6635,N_8680);
xnor U9640 (N_9640,N_6107,N_8117);
and U9641 (N_9641,N_8139,N_6938);
nand U9642 (N_9642,N_7098,N_7229);
or U9643 (N_9643,N_7398,N_8631);
nor U9644 (N_9644,N_7185,N_6977);
nor U9645 (N_9645,N_8393,N_8513);
nor U9646 (N_9646,N_8876,N_7803);
and U9647 (N_9647,N_6116,N_8868);
nand U9648 (N_9648,N_6969,N_7942);
nand U9649 (N_9649,N_6425,N_6367);
and U9650 (N_9650,N_8549,N_8555);
or U9651 (N_9651,N_8315,N_7821);
xor U9652 (N_9652,N_7661,N_8828);
or U9653 (N_9653,N_7679,N_6718);
xor U9654 (N_9654,N_8459,N_8639);
nor U9655 (N_9655,N_7177,N_8396);
nor U9656 (N_9656,N_6479,N_8341);
nand U9657 (N_9657,N_6724,N_7903);
nand U9658 (N_9658,N_6071,N_7230);
nand U9659 (N_9659,N_6044,N_7139);
and U9660 (N_9660,N_6536,N_6565);
or U9661 (N_9661,N_6142,N_8847);
or U9662 (N_9662,N_6347,N_7649);
nand U9663 (N_9663,N_7541,N_8871);
nor U9664 (N_9664,N_7749,N_7977);
or U9665 (N_9665,N_6104,N_8574);
xnor U9666 (N_9666,N_7008,N_6400);
nor U9667 (N_9667,N_6950,N_8151);
xnor U9668 (N_9668,N_8388,N_7590);
and U9669 (N_9669,N_8022,N_8067);
nor U9670 (N_9670,N_8253,N_8591);
nor U9671 (N_9671,N_7740,N_7067);
and U9672 (N_9672,N_7687,N_6419);
nand U9673 (N_9673,N_6796,N_8260);
nand U9674 (N_9674,N_6497,N_7491);
nand U9675 (N_9675,N_6238,N_6153);
nor U9676 (N_9676,N_6406,N_6607);
xor U9677 (N_9677,N_8992,N_7034);
xor U9678 (N_9678,N_8285,N_7481);
nor U9679 (N_9679,N_8464,N_8096);
nand U9680 (N_9680,N_6477,N_8596);
and U9681 (N_9681,N_8561,N_6599);
nor U9682 (N_9682,N_7434,N_6230);
or U9683 (N_9683,N_8978,N_6156);
nand U9684 (N_9684,N_7780,N_8961);
nor U9685 (N_9685,N_6883,N_8169);
nor U9686 (N_9686,N_6319,N_8934);
nor U9687 (N_9687,N_6093,N_7607);
and U9688 (N_9688,N_7264,N_6766);
or U9689 (N_9689,N_7835,N_6342);
nand U9690 (N_9690,N_6825,N_7265);
and U9691 (N_9691,N_7570,N_6598);
or U9692 (N_9692,N_6848,N_7097);
nor U9693 (N_9693,N_6498,N_8660);
xnor U9694 (N_9694,N_7906,N_7044);
and U9695 (N_9695,N_6244,N_8482);
nand U9696 (N_9696,N_6040,N_6853);
and U9697 (N_9697,N_6090,N_8990);
and U9698 (N_9698,N_6062,N_6719);
nand U9699 (N_9699,N_8636,N_6913);
nand U9700 (N_9700,N_6211,N_8817);
nand U9701 (N_9701,N_6785,N_6758);
and U9702 (N_9702,N_8289,N_7381);
or U9703 (N_9703,N_8330,N_6341);
nor U9704 (N_9704,N_6881,N_7329);
xnor U9705 (N_9705,N_6133,N_8273);
nor U9706 (N_9706,N_8360,N_8959);
nor U9707 (N_9707,N_8269,N_6253);
and U9708 (N_9708,N_6035,N_8423);
xor U9709 (N_9709,N_8390,N_7682);
and U9710 (N_9710,N_6381,N_8456);
nor U9711 (N_9711,N_7598,N_8255);
nand U9712 (N_9712,N_6279,N_8123);
and U9713 (N_9713,N_8894,N_7154);
nand U9714 (N_9714,N_6360,N_8426);
and U9715 (N_9715,N_8686,N_6914);
or U9716 (N_9716,N_8107,N_6387);
nor U9717 (N_9717,N_6989,N_8887);
nand U9718 (N_9718,N_6430,N_7859);
or U9719 (N_9719,N_8650,N_8379);
nor U9720 (N_9720,N_8471,N_8838);
nand U9721 (N_9721,N_6291,N_7452);
xnor U9722 (N_9722,N_7303,N_6000);
xnor U9723 (N_9723,N_8024,N_8664);
and U9724 (N_9724,N_6195,N_6522);
nor U9725 (N_9725,N_6112,N_7011);
and U9726 (N_9726,N_8465,N_8338);
nand U9727 (N_9727,N_8042,N_6025);
nand U9728 (N_9728,N_6450,N_8899);
and U9729 (N_9729,N_8912,N_6355);
nor U9730 (N_9730,N_8043,N_8951);
and U9731 (N_9731,N_7647,N_7466);
xnor U9732 (N_9732,N_8150,N_7200);
xnor U9733 (N_9733,N_8747,N_7212);
and U9734 (N_9734,N_7564,N_6095);
and U9735 (N_9735,N_6084,N_7179);
and U9736 (N_9736,N_7253,N_7327);
nand U9737 (N_9737,N_7138,N_7978);
xor U9738 (N_9738,N_6625,N_8626);
nor U9739 (N_9739,N_6414,N_7372);
xor U9740 (N_9740,N_7939,N_8256);
nor U9741 (N_9741,N_8259,N_8737);
and U9742 (N_9742,N_8511,N_6927);
and U9743 (N_9743,N_6313,N_8344);
and U9744 (N_9744,N_6833,N_7787);
nor U9745 (N_9745,N_6570,N_6210);
nor U9746 (N_9746,N_7545,N_7917);
and U9747 (N_9747,N_6388,N_7305);
nand U9748 (N_9748,N_7574,N_8744);
nor U9749 (N_9749,N_8671,N_7002);
xor U9750 (N_9750,N_6597,N_6365);
nor U9751 (N_9751,N_7997,N_6617);
or U9752 (N_9752,N_7877,N_6424);
and U9753 (N_9753,N_7088,N_6505);
nand U9754 (N_9754,N_6921,N_6078);
or U9755 (N_9755,N_6872,N_6270);
xnor U9756 (N_9756,N_8470,N_8240);
nand U9757 (N_9757,N_8385,N_6038);
nor U9758 (N_9758,N_8268,N_6640);
nand U9759 (N_9759,N_6767,N_6684);
nand U9760 (N_9760,N_8672,N_7003);
nand U9761 (N_9761,N_8145,N_8262);
xnor U9762 (N_9762,N_7672,N_8271);
nand U9763 (N_9763,N_6213,N_8901);
and U9764 (N_9764,N_7814,N_6073);
xor U9765 (N_9765,N_6539,N_7315);
and U9766 (N_9766,N_8743,N_8742);
and U9767 (N_9767,N_7458,N_6017);
or U9768 (N_9768,N_8502,N_8376);
or U9769 (N_9769,N_8771,N_6696);
and U9770 (N_9770,N_8573,N_8553);
and U9771 (N_9771,N_8835,N_7823);
or U9772 (N_9772,N_7674,N_7288);
nor U9773 (N_9773,N_7095,N_7976);
and U9774 (N_9774,N_8367,N_7644);
or U9775 (N_9775,N_7848,N_7860);
or U9776 (N_9776,N_7101,N_6386);
or U9777 (N_9777,N_6098,N_7463);
and U9778 (N_9778,N_8656,N_7698);
xnor U9779 (N_9779,N_6021,N_8443);
nand U9780 (N_9780,N_6966,N_7907);
or U9781 (N_9781,N_6431,N_8572);
nand U9782 (N_9782,N_8191,N_8475);
and U9783 (N_9783,N_6733,N_6079);
and U9784 (N_9784,N_7724,N_8203);
nand U9785 (N_9785,N_8973,N_6807);
xor U9786 (N_9786,N_8345,N_8424);
xor U9787 (N_9787,N_8673,N_6551);
nor U9788 (N_9788,N_7718,N_8294);
or U9789 (N_9789,N_7358,N_7650);
or U9790 (N_9790,N_7946,N_6549);
and U9791 (N_9791,N_7075,N_8770);
or U9792 (N_9792,N_8350,N_6069);
nor U9793 (N_9793,N_8391,N_7228);
xnor U9794 (N_9794,N_6281,N_8034);
nor U9795 (N_9795,N_8035,N_6973);
and U9796 (N_9796,N_8319,N_7399);
nand U9797 (N_9797,N_8053,N_7449);
or U9798 (N_9798,N_6583,N_7548);
or U9799 (N_9799,N_8198,N_8723);
nor U9800 (N_9800,N_8286,N_7465);
nand U9801 (N_9801,N_6943,N_8820);
or U9802 (N_9802,N_8377,N_7691);
nand U9803 (N_9803,N_7429,N_6944);
or U9804 (N_9804,N_8738,N_7810);
xnor U9805 (N_9805,N_6644,N_6856);
xnor U9806 (N_9806,N_7215,N_7660);
xnor U9807 (N_9807,N_6261,N_8907);
or U9808 (N_9808,N_6521,N_6651);
nor U9809 (N_9809,N_6067,N_8694);
xnor U9810 (N_9810,N_7105,N_6377);
and U9811 (N_9811,N_7426,N_7713);
nand U9812 (N_9812,N_6908,N_6765);
nand U9813 (N_9813,N_8332,N_7735);
or U9814 (N_9814,N_7207,N_7585);
xnor U9815 (N_9815,N_7544,N_7056);
nand U9816 (N_9816,N_8560,N_8942);
nand U9817 (N_9817,N_8125,N_8881);
or U9818 (N_9818,N_7080,N_8933);
xor U9819 (N_9819,N_6292,N_8796);
nand U9820 (N_9820,N_7018,N_7919);
nor U9821 (N_9821,N_6231,N_7850);
nand U9822 (N_9822,N_7728,N_7868);
and U9823 (N_9823,N_6197,N_7727);
xnor U9824 (N_9824,N_6061,N_7816);
and U9825 (N_9825,N_6370,N_6242);
or U9826 (N_9826,N_7106,N_8862);
nor U9827 (N_9827,N_6618,N_7549);
xor U9828 (N_9828,N_7257,N_6926);
or U9829 (N_9829,N_6357,N_6082);
or U9830 (N_9830,N_8655,N_7568);
xor U9831 (N_9831,N_7887,N_7684);
and U9832 (N_9832,N_6849,N_7899);
and U9833 (N_9833,N_8701,N_6988);
xnor U9834 (N_9834,N_8033,N_8485);
nor U9835 (N_9835,N_7783,N_8258);
or U9836 (N_9836,N_7869,N_8242);
xor U9837 (N_9837,N_8851,N_7186);
nor U9838 (N_9838,N_7914,N_6366);
nand U9839 (N_9839,N_6511,N_8403);
xnor U9840 (N_9840,N_6389,N_7451);
or U9841 (N_9841,N_8389,N_7150);
and U9842 (N_9842,N_7743,N_7957);
nor U9843 (N_9843,N_6563,N_7741);
nor U9844 (N_9844,N_6026,N_8472);
xnor U9845 (N_9845,N_7346,N_6837);
nor U9846 (N_9846,N_7849,N_8414);
or U9847 (N_9847,N_8799,N_6220);
and U9848 (N_9848,N_8100,N_8102);
nand U9849 (N_9849,N_8834,N_8369);
or U9850 (N_9850,N_6693,N_6216);
nor U9851 (N_9851,N_7947,N_6622);
nand U9852 (N_9852,N_6930,N_7736);
xnor U9853 (N_9853,N_7553,N_6383);
nand U9854 (N_9854,N_8644,N_7828);
nor U9855 (N_9855,N_7261,N_7798);
xor U9856 (N_9856,N_7916,N_7021);
or U9857 (N_9857,N_7089,N_7060);
nor U9858 (N_9858,N_8324,N_6240);
and U9859 (N_9859,N_7062,N_6187);
xor U9860 (N_9860,N_8699,N_7324);
nor U9861 (N_9861,N_7326,N_6232);
nand U9862 (N_9862,N_6191,N_7015);
xor U9863 (N_9863,N_6792,N_7243);
nor U9864 (N_9864,N_8927,N_7389);
xnor U9865 (N_9865,N_6379,N_7593);
xnor U9866 (N_9866,N_7540,N_6455);
xnor U9867 (N_9867,N_6437,N_7333);
or U9868 (N_9868,N_8115,N_7066);
or U9869 (N_9869,N_8633,N_8015);
nor U9870 (N_9870,N_7913,N_7161);
nor U9871 (N_9871,N_7292,N_8136);
nor U9872 (N_9872,N_6712,N_6979);
or U9873 (N_9873,N_6148,N_7985);
or U9874 (N_9874,N_6447,N_8120);
and U9875 (N_9875,N_8094,N_8897);
and U9876 (N_9876,N_7676,N_6854);
nor U9877 (N_9877,N_6905,N_6643);
nor U9878 (N_9878,N_6860,N_6713);
nor U9879 (N_9879,N_8062,N_7567);
or U9880 (N_9880,N_7453,N_6096);
nor U9881 (N_9881,N_8915,N_8026);
nand U9882 (N_9882,N_8518,N_8867);
nor U9883 (N_9883,N_8823,N_8645);
xnor U9884 (N_9884,N_7817,N_6034);
nor U9885 (N_9885,N_6747,N_8906);
nor U9886 (N_9886,N_8970,N_8236);
nor U9887 (N_9887,N_8248,N_8413);
and U9888 (N_9888,N_7433,N_8241);
or U9889 (N_9889,N_8832,N_6322);
nor U9890 (N_9890,N_7934,N_7834);
or U9891 (N_9891,N_7450,N_6124);
nor U9892 (N_9892,N_8448,N_8842);
xnor U9893 (N_9893,N_6730,N_7739);
nand U9894 (N_9894,N_7663,N_6834);
xnor U9895 (N_9895,N_7927,N_6019);
and U9896 (N_9896,N_7404,N_7608);
nand U9897 (N_9897,N_6556,N_6659);
nor U9898 (N_9898,N_8625,N_6346);
nand U9899 (N_9899,N_8244,N_6958);
nor U9900 (N_9900,N_7199,N_8041);
nor U9901 (N_9901,N_6129,N_6161);
xor U9902 (N_9902,N_8854,N_6862);
nor U9903 (N_9903,N_6251,N_8665);
or U9904 (N_9904,N_8333,N_6698);
or U9905 (N_9905,N_8190,N_6955);
or U9906 (N_9906,N_7511,N_6658);
or U9907 (N_9907,N_8728,N_6154);
and U9908 (N_9908,N_6474,N_7446);
nor U9909 (N_9909,N_7987,N_7994);
or U9910 (N_9910,N_6939,N_6874);
xor U9911 (N_9911,N_6987,N_6928);
nand U9912 (N_9912,N_8049,N_8222);
nand U9913 (N_9913,N_8936,N_7267);
or U9914 (N_9914,N_8204,N_6398);
nand U9915 (N_9915,N_7866,N_7110);
xnor U9916 (N_9916,N_6352,N_8308);
and U9917 (N_9917,N_8302,N_6541);
xor U9918 (N_9918,N_7675,N_6199);
or U9919 (N_9919,N_8353,N_6368);
nand U9920 (N_9920,N_7348,N_6041);
xor U9921 (N_9921,N_7852,N_7589);
nor U9922 (N_9922,N_8055,N_8159);
nor U9923 (N_9923,N_6535,N_6514);
and U9924 (N_9924,N_6333,N_7516);
or U9925 (N_9925,N_7584,N_6959);
nand U9926 (N_9926,N_7826,N_6439);
and U9927 (N_9927,N_7751,N_6815);
xnor U9928 (N_9928,N_8716,N_6694);
xnor U9929 (N_9929,N_7304,N_8776);
or U9930 (N_9930,N_8314,N_7149);
xor U9931 (N_9931,N_7789,N_8944);
and U9932 (N_9932,N_8888,N_8615);
and U9933 (N_9933,N_6385,N_6176);
nand U9934 (N_9934,N_6887,N_7775);
nor U9935 (N_9935,N_8630,N_7208);
nand U9936 (N_9936,N_6118,N_8104);
nand U9937 (N_9937,N_6538,N_8277);
nor U9938 (N_9938,N_7380,N_7447);
nor U9939 (N_9939,N_8850,N_7152);
or U9940 (N_9940,N_6066,N_6267);
or U9941 (N_9941,N_6791,N_7983);
and U9942 (N_9942,N_6214,N_6573);
nand U9943 (N_9943,N_6941,N_6190);
nand U9944 (N_9944,N_6426,N_8493);
and U9945 (N_9945,N_6965,N_6131);
nor U9946 (N_9946,N_8496,N_6212);
and U9947 (N_9947,N_8900,N_6691);
or U9948 (N_9948,N_8983,N_7222);
xnor U9949 (N_9949,N_6817,N_7423);
xnor U9950 (N_9950,N_6286,N_7065);
and U9951 (N_9951,N_6378,N_7431);
nand U9952 (N_9952,N_8484,N_6177);
nor U9953 (N_9953,N_8155,N_6137);
xor U9954 (N_9954,N_6166,N_7981);
or U9955 (N_9955,N_6396,N_8889);
nand U9956 (N_9956,N_7582,N_6998);
nor U9957 (N_9957,N_8902,N_6454);
xor U9958 (N_9958,N_8860,N_7032);
xor U9959 (N_9959,N_6818,N_7791);
xor U9960 (N_9960,N_7528,N_6298);
nand U9961 (N_9961,N_6512,N_7617);
and U9962 (N_9962,N_6374,N_7892);
or U9963 (N_9963,N_6217,N_6508);
or U9964 (N_9964,N_6336,N_6816);
and U9965 (N_9965,N_6688,N_6686);
xnor U9966 (N_9966,N_7496,N_6203);
and U9967 (N_9967,N_7744,N_8010);
nand U9968 (N_9968,N_7162,N_6912);
or U9969 (N_9969,N_8760,N_8751);
nand U9970 (N_9970,N_7051,N_7205);
or U9971 (N_9971,N_6985,N_7130);
xor U9972 (N_9972,N_6283,N_6729);
or U9973 (N_9973,N_7140,N_7757);
nor U9974 (N_9974,N_6761,N_7700);
nand U9975 (N_9975,N_6192,N_6310);
nand U9976 (N_9976,N_7403,N_8225);
xor U9977 (N_9977,N_8733,N_8641);
and U9978 (N_9978,N_7040,N_8780);
xor U9979 (N_9979,N_7708,N_6465);
nor U9980 (N_9980,N_7249,N_7116);
and U9981 (N_9981,N_6589,N_6323);
nor U9982 (N_9982,N_6287,N_6706);
nor U9983 (N_9983,N_8946,N_8684);
and U9984 (N_9984,N_7216,N_8468);
xor U9985 (N_9985,N_7441,N_7219);
and U9986 (N_9986,N_6550,N_7664);
nand U9987 (N_9987,N_8547,N_7878);
xor U9988 (N_9988,N_7822,N_7566);
and U9989 (N_9989,N_7921,N_7277);
nor U9990 (N_9990,N_6546,N_8865);
nand U9991 (N_9991,N_8804,N_8757);
or U9992 (N_9992,N_7218,N_6942);
or U9993 (N_9993,N_8707,N_6878);
and U9994 (N_9994,N_6861,N_6870);
and U9995 (N_9995,N_7622,N_6593);
nor U9996 (N_9996,N_7677,N_7157);
or U9997 (N_9997,N_7163,N_8354);
nor U9998 (N_9998,N_6904,N_7729);
or U9999 (N_9999,N_8773,N_6893);
or U10000 (N_10000,N_7046,N_8515);
nor U10001 (N_10001,N_7472,N_7370);
and U10002 (N_10002,N_8637,N_8898);
nor U10003 (N_10003,N_7683,N_8984);
nor U10004 (N_10004,N_7636,N_7813);
xor U10005 (N_10005,N_8313,N_7587);
nor U10006 (N_10006,N_8486,N_6036);
nand U10007 (N_10007,N_6687,N_8782);
nand U10008 (N_10008,N_6841,N_7766);
nand U10009 (N_10009,N_7945,N_7133);
xnor U10010 (N_10010,N_6711,N_7223);
nand U10011 (N_10011,N_7697,N_7991);
xnor U10012 (N_10012,N_7084,N_7388);
nand U10013 (N_10013,N_7646,N_7882);
or U10014 (N_10014,N_8007,N_7610);
and U10015 (N_10015,N_8687,N_8506);
or U10016 (N_10016,N_8654,N_7825);
and U10017 (N_10017,N_6415,N_7858);
or U10018 (N_10018,N_7777,N_7119);
xor U10019 (N_10019,N_6506,N_8563);
and U10020 (N_10020,N_6513,N_6502);
xnor U10021 (N_10021,N_6920,N_7396);
nand U10022 (N_10022,N_7144,N_6410);
nand U10023 (N_10023,N_6734,N_7936);
nand U10024 (N_10024,N_7872,N_7794);
nand U10025 (N_10025,N_7013,N_7120);
xor U10026 (N_10026,N_7485,N_7795);
and U10027 (N_10027,N_7591,N_6371);
and U10028 (N_10028,N_8480,N_6648);
nor U10029 (N_10029,N_7014,N_6351);
nand U10030 (N_10030,N_7376,N_6273);
xor U10031 (N_10031,N_6250,N_6050);
xnor U10032 (N_10032,N_6417,N_7132);
nand U10033 (N_10033,N_6045,N_7425);
nand U10034 (N_10034,N_8237,N_7896);
nor U10035 (N_10035,N_8274,N_7320);
nand U10036 (N_10036,N_6954,N_8891);
or U10037 (N_10037,N_6581,N_6088);
nand U10038 (N_10038,N_7217,N_6068);
and U10039 (N_10039,N_7368,N_8073);
or U10040 (N_10040,N_8492,N_6517);
nand U10041 (N_10041,N_6046,N_8095);
xnor U10042 (N_10042,N_6441,N_7845);
and U10043 (N_10043,N_6846,N_6249);
nor U10044 (N_10044,N_7786,N_7804);
and U10045 (N_10045,N_8186,N_7394);
and U10046 (N_10046,N_6268,N_7961);
or U10047 (N_10047,N_8156,N_8956);
and U10048 (N_10048,N_7039,N_8619);
xor U10049 (N_10049,N_6359,N_8559);
and U10050 (N_10050,N_7602,N_8883);
xnor U10051 (N_10051,N_6576,N_8709);
nor U10052 (N_10052,N_8529,N_6135);
nor U10053 (N_10053,N_7853,N_6030);
xor U10054 (N_10054,N_8079,N_7297);
and U10055 (N_10055,N_6013,N_6557);
nand U10056 (N_10056,N_6771,N_7773);
or U10057 (N_10057,N_8336,N_6653);
xor U10058 (N_10058,N_8383,N_6520);
or U10059 (N_10059,N_7419,N_6880);
nand U10060 (N_10060,N_8036,N_8401);
nand U10061 (N_10061,N_7131,N_8587);
xor U10062 (N_10062,N_8019,N_8605);
or U10063 (N_10063,N_6548,N_7569);
nand U10064 (N_10064,N_8106,N_8378);
nand U10065 (N_10065,N_6695,N_6674);
and U10066 (N_10066,N_7524,N_7330);
nand U10067 (N_10067,N_6602,N_8339);
nand U10068 (N_10068,N_6631,N_8346);
xnor U10069 (N_10069,N_6145,N_6404);
nor U10070 (N_10070,N_8642,N_6993);
nand U10071 (N_10071,N_7668,N_7632);
nor U10072 (N_10072,N_8839,N_6185);
nand U10073 (N_10073,N_8768,N_6006);
and U10074 (N_10074,N_7819,N_8362);
nand U10075 (N_10075,N_7551,N_7286);
or U10076 (N_10076,N_7599,N_8532);
and U10077 (N_10077,N_7962,N_8220);
or U10078 (N_10078,N_7606,N_7279);
nand U10079 (N_10079,N_7665,N_7841);
xnor U10080 (N_10080,N_8417,N_7357);
nand U10081 (N_10081,N_6460,N_7639);
or U10082 (N_10082,N_7038,N_7108);
xor U10083 (N_10083,N_6194,N_6555);
or U10084 (N_10084,N_7645,N_8501);
and U10085 (N_10085,N_8952,N_6469);
and U10086 (N_10086,N_6031,N_7955);
and U10087 (N_10087,N_6125,N_7952);
and U10088 (N_10088,N_6847,N_7275);
and U10089 (N_10089,N_7717,N_6339);
and U10090 (N_10090,N_8721,N_8717);
and U10091 (N_10091,N_7986,N_6119);
xor U10092 (N_10092,N_7756,N_8276);
and U10093 (N_10093,N_8938,N_6890);
or U10094 (N_10094,N_7328,N_7747);
or U10095 (N_10095,N_6773,N_7619);
or U10096 (N_10096,N_6740,N_8309);
nand U10097 (N_10097,N_7560,N_7183);
nor U10098 (N_10098,N_7626,N_8893);
nor U10099 (N_10099,N_6235,N_7312);
nand U10100 (N_10100,N_6770,N_6981);
xor U10101 (N_10101,N_6260,N_8869);
xor U10102 (N_10102,N_7851,N_7969);
nand U10103 (N_10103,N_7839,N_8538);
nand U10104 (N_10104,N_6937,N_7387);
nor U10105 (N_10105,N_7031,N_8556);
and U10106 (N_10106,N_7601,N_7628);
nor U10107 (N_10107,N_6976,N_8128);
and U10108 (N_10108,N_7552,N_8152);
nand U10109 (N_10109,N_7529,N_6047);
nand U10110 (N_10110,N_6002,N_7531);
and U10111 (N_10111,N_6667,N_6996);
nor U10112 (N_10112,N_7820,N_8446);
xor U10113 (N_10113,N_8885,N_8059);
nor U10114 (N_10114,N_8473,N_8706);
nor U10115 (N_10115,N_6604,N_6325);
nand U10116 (N_10116,N_7147,N_6072);
or U10117 (N_10117,N_8065,N_6380);
nand U10118 (N_10118,N_8647,N_7671);
xor U10119 (N_10119,N_6011,N_8568);
or U10120 (N_10120,N_8986,N_6885);
nor U10121 (N_10121,N_6587,N_8080);
and U10122 (N_10122,N_6553,N_7754);
and U10123 (N_10123,N_6032,N_8178);
xor U10124 (N_10124,N_7309,N_8278);
and U10125 (N_10125,N_8777,N_7166);
or U10126 (N_10126,N_8397,N_6495);
and U10127 (N_10127,N_8775,N_6488);
xnor U10128 (N_10128,N_7854,N_7349);
nand U10129 (N_10129,N_7492,N_7256);
and U10130 (N_10130,N_7760,N_6223);
xnor U10131 (N_10131,N_8575,N_6157);
and U10132 (N_10132,N_8387,N_6956);
xor U10133 (N_10133,N_7818,N_6971);
nor U10134 (N_10134,N_7512,N_7035);
xor U10135 (N_10135,N_6438,N_7369);
or U10136 (N_10136,N_7581,N_6634);
and U10137 (N_10137,N_8020,N_8857);
nor U10138 (N_10138,N_8974,N_6924);
and U10139 (N_10139,N_8144,N_6186);
xor U10140 (N_10140,N_6842,N_7467);
xnor U10141 (N_10141,N_8076,N_7203);
nand U10142 (N_10142,N_8730,N_7518);
and U10143 (N_10143,N_6624,N_6289);
xnor U10144 (N_10144,N_8469,N_8963);
or U10145 (N_10145,N_8182,N_7807);
xnor U10146 (N_10146,N_8689,N_7190);
xnor U10147 (N_10147,N_8295,N_7709);
and U10148 (N_10148,N_6492,N_6844);
nand U10149 (N_10149,N_8841,N_6601);
and U10150 (N_10150,N_7536,N_6945);
and U10151 (N_10151,N_7681,N_6312);
or U10152 (N_10152,N_6141,N_7104);
or U10153 (N_10153,N_7950,N_6524);
and U10154 (N_10154,N_8452,N_6405);
and U10155 (N_10155,N_6152,N_6571);
xor U10156 (N_10156,N_7053,N_6992);
and U10157 (N_10157,N_7964,N_8710);
or U10158 (N_10158,N_6923,N_8083);
nand U10159 (N_10159,N_7172,N_8981);
nand U10160 (N_10160,N_7115,N_7558);
nor U10161 (N_10161,N_6092,N_8638);
nor U10162 (N_10162,N_6780,N_7776);
nand U10163 (N_10163,N_6089,N_8057);
or U10164 (N_10164,N_7513,N_7507);
or U10165 (N_10165,N_7966,N_7680);
nor U10166 (N_10166,N_6616,N_6269);
nand U10167 (N_10167,N_8994,N_6180);
nor U10168 (N_10168,N_7904,N_6819);
or U10169 (N_10169,N_6614,N_7797);
xor U10170 (N_10170,N_7614,N_7716);
or U10171 (N_10171,N_6826,N_6675);
xor U10172 (N_10172,N_8536,N_6737);
xnor U10173 (N_10173,N_7862,N_8504);
nor U10174 (N_10174,N_8091,N_8712);
or U10175 (N_10175,N_6130,N_7809);
xnor U10176 (N_10176,N_7605,N_7571);
and U10177 (N_10177,N_7720,N_8866);
xor U10178 (N_10178,N_6964,N_7440);
nand U10179 (N_10179,N_7996,N_6709);
and U10180 (N_10180,N_7768,N_8827);
nand U10181 (N_10181,N_7006,N_6039);
nand U10182 (N_10182,N_6701,N_7213);
xor U10183 (N_10183,N_8304,N_8904);
nand U10184 (N_10184,N_7926,N_6916);
and U10185 (N_10185,N_6482,N_6297);
nand U10186 (N_10186,N_6739,N_6043);
xnor U10187 (N_10187,N_8989,N_6811);
and U10188 (N_10188,N_7225,N_7438);
and U10189 (N_10189,N_8571,N_7517);
xor U10190 (N_10190,N_7322,N_6493);
or U10191 (N_10191,N_7990,N_6467);
or U10192 (N_10192,N_6376,N_8442);
or U10193 (N_10193,N_8162,N_6799);
or U10194 (N_10194,N_8066,N_8266);
and U10195 (N_10195,N_6416,N_7195);
and U10196 (N_10196,N_6306,N_6915);
or U10197 (N_10197,N_8250,N_6466);
nor U10198 (N_10198,N_7180,N_8134);
nor U10199 (N_10199,N_8119,N_8215);
and U10200 (N_10200,N_7792,N_8811);
or U10201 (N_10201,N_6970,N_8600);
and U10202 (N_10202,N_6829,N_6301);
nand U10203 (N_10203,N_7931,N_7156);
nand U10204 (N_10204,N_6101,N_7730);
nand U10205 (N_10205,N_8185,N_6953);
nand U10206 (N_10206,N_7079,N_7956);
nor U10207 (N_10207,N_8224,N_6962);
nand U10208 (N_10208,N_7221,N_7958);
and U10209 (N_10209,N_8873,N_8195);
and U10210 (N_10210,N_7493,N_6561);
nor U10211 (N_10211,N_6507,N_7395);
xnor U10212 (N_10212,N_7094,N_6115);
or U10213 (N_10213,N_6080,N_6661);
xnor U10214 (N_10214,N_8601,N_8545);
nand U10215 (N_10215,N_8488,N_7634);
nand U10216 (N_10216,N_8525,N_7247);
nor U10217 (N_10217,N_7575,N_6824);
or U10218 (N_10218,N_8921,N_6731);
xnor U10219 (N_10219,N_7714,N_6525);
nor U10220 (N_10220,N_8969,N_6586);
xnor U10221 (N_10221,N_6139,N_6397);
nor U10222 (N_10222,N_8221,N_7533);
and U10223 (N_10223,N_7168,N_6395);
nand U10224 (N_10224,N_6746,N_8257);
nor U10225 (N_10225,N_6173,N_7214);
nand U10226 (N_10226,N_7520,N_8193);
nor U10227 (N_10227,N_6103,N_8454);
xnor U10228 (N_10228,N_8245,N_6523);
xor U10229 (N_10229,N_7891,N_8932);
nand U10230 (N_10230,N_6461,N_8750);
nor U10231 (N_10231,N_7763,N_8569);
nor U10232 (N_10232,N_7024,N_8054);
nor U10233 (N_10233,N_7272,N_6063);
or U10234 (N_10234,N_8368,N_7386);
and U10235 (N_10235,N_8949,N_7980);
nor U10236 (N_10236,N_7142,N_6463);
nor U10237 (N_10237,N_8441,N_8863);
nand U10238 (N_10238,N_8629,N_7801);
or U10239 (N_10239,N_7722,N_6820);
xor U10240 (N_10240,N_6879,N_6999);
nand U10241 (N_10241,N_7542,N_8566);
xnor U10242 (N_10242,N_7137,N_7129);
nor U10243 (N_10243,N_6642,N_7235);
or U10244 (N_10244,N_7151,N_8082);
and U10245 (N_10245,N_8852,N_7042);
nand U10246 (N_10246,N_7501,N_8071);
nor U10247 (N_10247,N_6699,N_6016);
xor U10248 (N_10248,N_6823,N_7476);
and U10249 (N_10249,N_8657,N_6656);
nand U10250 (N_10250,N_7427,N_8697);
nor U10251 (N_10251,N_7158,N_7334);
or U10252 (N_10252,N_6171,N_7454);
and U10253 (N_10253,N_8160,N_7464);
nor U10254 (N_10254,N_7688,N_6613);
nor U10255 (N_10255,N_6218,N_8051);
xor U10256 (N_10256,N_6935,N_8060);
nand U10257 (N_10257,N_8542,N_8524);
xor U10258 (N_10258,N_6010,N_8300);
or U10259 (N_10259,N_6361,N_8138);
and U10260 (N_10260,N_8093,N_8021);
or U10261 (N_10261,N_6605,N_8971);
or U10262 (N_10262,N_8602,N_6198);
nand U10263 (N_10263,N_8565,N_6164);
nand U10264 (N_10264,N_7176,N_6271);
xor U10265 (N_10265,N_7242,N_7897);
nand U10266 (N_10266,N_8476,N_8412);
nand U10267 (N_10267,N_6049,N_8165);
nand U10268 (N_10268,N_6018,N_6532);
nand U10269 (N_10269,N_6784,N_8995);
nand U10270 (N_10270,N_7631,N_8199);
xor U10271 (N_10271,N_6318,N_7250);
nand U10272 (N_10272,N_8163,N_8461);
xor U10273 (N_10273,N_7238,N_6316);
nand U10274 (N_10274,N_7745,N_6295);
nor U10275 (N_10275,N_7407,N_7686);
and U10276 (N_10276,N_7886,N_8552);
xor U10277 (N_10277,N_8681,N_8211);
and U10278 (N_10278,N_6882,N_7502);
xnor U10279 (N_10279,N_6788,N_6138);
nand U10280 (N_10280,N_8864,N_7041);
and U10281 (N_10281,N_6022,N_7615);
or U10282 (N_10282,N_6588,N_7082);
nor U10283 (N_10283,N_7076,N_7255);
and U10284 (N_10284,N_8570,N_7342);
nand U10285 (N_10285,N_6591,N_8479);
or U10286 (N_10286,N_6307,N_7362);
nand U10287 (N_10287,N_7459,N_7579);
xnor U10288 (N_10288,N_6786,N_7975);
nor U10289 (N_10289,N_7052,N_8372);
nor U10290 (N_10290,N_8627,N_8291);
xnor U10291 (N_10291,N_6621,N_6233);
xor U10292 (N_10292,N_6918,N_7000);
xnor U10293 (N_10293,N_7236,N_7556);
xnor U10294 (N_10294,N_6382,N_7070);
nand U10295 (N_10295,N_7705,N_6196);
and U10296 (N_10296,N_8816,N_7901);
nand U10297 (N_10297,N_6259,N_6707);
nand U10298 (N_10298,N_7457,N_7920);
and U10299 (N_10299,N_6282,N_7424);
nand U10300 (N_10300,N_6660,N_8892);
and U10301 (N_10301,N_8837,N_8261);
nor U10302 (N_10302,N_7068,N_7500);
nand U10303 (N_10303,N_8512,N_6608);
or U10304 (N_10304,N_7483,N_8913);
xor U10305 (N_10305,N_7174,N_8075);
xnor U10306 (N_10306,N_7189,N_6762);
nand U10307 (N_10307,N_8807,N_7561);
nor U10308 (N_10308,N_7538,N_6053);
nor U10309 (N_10309,N_8919,N_8676);
or U10310 (N_10310,N_8954,N_7840);
or U10311 (N_10311,N_6226,N_6059);
nand U10312 (N_10312,N_6225,N_6869);
nor U10313 (N_10313,N_6654,N_8265);
or U10314 (N_10314,N_6710,N_6446);
nand U10315 (N_10315,N_7410,N_7532);
and U10316 (N_10316,N_8374,N_6064);
nor U10317 (N_10317,N_7537,N_7437);
nor U10318 (N_10318,N_8180,N_8478);
nor U10319 (N_10319,N_8794,N_6356);
and U10320 (N_10320,N_6980,N_6615);
or U10321 (N_10321,N_6087,N_8875);
nor U10322 (N_10322,N_7490,N_7565);
and U10323 (N_10323,N_8425,N_6014);
and U10324 (N_10324,N_6714,N_8661);
or U10325 (N_10325,N_8439,N_6136);
nand U10326 (N_10326,N_8640,N_7415);
or U10327 (N_10327,N_8985,N_6794);
xor U10328 (N_10328,N_6280,N_6464);
or U10329 (N_10329,N_8758,N_7884);
nor U10330 (N_10330,N_7930,N_8074);
nand U10331 (N_10331,N_8683,N_6827);
nand U10332 (N_10332,N_8375,N_8173);
or U10333 (N_10333,N_8713,N_6630);
xor U10334 (N_10334,N_8063,N_7588);
and U10335 (N_10335,N_8788,N_6327);
and U10336 (N_10336,N_6284,N_6759);
xnor U10337 (N_10337,N_6678,N_8192);
nand U10338 (N_10338,N_6673,N_8908);
nor U10339 (N_10339,N_8749,N_8520);
nand U10340 (N_10340,N_8061,N_7918);
or U10341 (N_10341,N_7251,N_7624);
nor U10342 (N_10342,N_7988,N_6472);
and U10343 (N_10343,N_6984,N_7456);
and U10344 (N_10344,N_7559,N_7706);
and U10345 (N_10345,N_6704,N_7871);
or U10346 (N_10346,N_7912,N_8167);
nand U10347 (N_10347,N_6150,N_6422);
nand U10348 (N_10348,N_7846,N_8135);
and U10349 (N_10349,N_6655,N_8038);
nand U10350 (N_10350,N_6802,N_6925);
xnor U10351 (N_10351,N_8078,N_8340);
xor U10352 (N_10352,N_8740,N_8451);
or U10353 (N_10353,N_7712,N_6027);
and U10354 (N_10354,N_8980,N_7693);
nand U10355 (N_10355,N_7462,N_7935);
and U10356 (N_10356,N_8176,N_6813);
nor U10357 (N_10357,N_7204,N_8483);
xor U10358 (N_10358,N_7036,N_6967);
nor U10359 (N_10359,N_6344,N_7737);
or U10360 (N_10360,N_6606,N_7072);
xnor U10361 (N_10361,N_8840,N_6120);
xor U10362 (N_10362,N_8928,N_8735);
xnor U10363 (N_10363,N_6832,N_6293);
nand U10364 (N_10364,N_6922,N_6685);
or U10365 (N_10365,N_8539,N_7600);
xnor U10366 (N_10366,N_6623,N_8855);
and U10367 (N_10367,N_8001,N_6743);
xnor U10368 (N_10368,N_7662,N_7908);
or U10369 (N_10369,N_7428,N_6515);
and U10370 (N_10370,N_7526,N_8703);
xnor U10371 (N_10371,N_6433,N_8187);
and U10372 (N_10372,N_8595,N_7742);
nand U10373 (N_10373,N_7331,N_7648);
nor U10374 (N_10374,N_8435,N_8416);
nor U10375 (N_10375,N_7086,N_6094);
or U10376 (N_10376,N_8202,N_7974);
nand U10377 (N_10377,N_6256,N_7422);
and U10378 (N_10378,N_7703,N_8670);
and U10379 (N_10379,N_7902,N_8668);
nand U10380 (N_10380,N_6600,N_7475);
nand U10381 (N_10381,N_6812,N_6896);
and U10382 (N_10382,N_6165,N_7772);
nand U10383 (N_10383,N_8326,N_8968);
nor U10384 (N_10384,N_7625,N_7392);
nand U10385 (N_10385,N_6609,N_8301);
and U10386 (N_10386,N_8722,N_6184);
nor U10387 (N_10387,N_7103,N_6768);
xnor U10388 (N_10388,N_6324,N_8018);
and U10389 (N_10389,N_7146,N_6337);
nor U10390 (N_10390,N_8219,N_8494);
nand U10391 (N_10391,N_6384,N_6839);
and U10392 (N_10392,N_8305,N_8844);
and U10393 (N_10393,N_8769,N_6457);
and U10394 (N_10394,N_6692,N_6127);
or U10395 (N_10395,N_6723,N_7515);
nor U10396 (N_10396,N_6001,N_8349);
nor U10397 (N_10397,N_6296,N_6445);
and U10398 (N_10398,N_7543,N_8806);
nand U10399 (N_10399,N_8099,N_8603);
nor U10400 (N_10400,N_7750,N_8675);
and U10401 (N_10401,N_7226,N_7193);
nor U10402 (N_10402,N_7197,N_8802);
nand U10403 (N_10403,N_8614,N_7136);
and U10404 (N_10404,N_7379,N_7521);
and U10405 (N_10405,N_7618,N_6348);
nand U10406 (N_10406,N_6204,N_7390);
nand U10407 (N_10407,N_6744,N_6449);
or U10408 (N_10408,N_8546,N_7790);
xnor U10409 (N_10409,N_8745,N_8617);
xor U10410 (N_10410,N_7184,N_6875);
and U10411 (N_10411,N_8238,N_6448);
nor U10412 (N_10412,N_6051,N_8089);
and U10413 (N_10413,N_8433,N_8752);
and U10414 (N_10414,N_8359,N_6340);
nor U10415 (N_10415,N_8334,N_8700);
xor U10416 (N_10416,N_8122,N_6501);
nor U10417 (N_10417,N_7643,N_8081);
nor U10418 (N_10418,N_7782,N_6429);
xor U10419 (N_10419,N_6568,N_7690);
xnor U10420 (N_10420,N_8905,N_6174);
xor U10421 (N_10421,N_6902,N_8761);
nor U10422 (N_10422,N_6899,N_8006);
nor U10423 (N_10423,N_8429,N_8040);
xor U10424 (N_10424,N_7949,N_7796);
nor U10425 (N_10425,N_8137,N_6974);
nor U10426 (N_10426,N_8143,N_8643);
nor U10427 (N_10427,N_8498,N_8329);
nand U10428 (N_10428,N_6645,N_6948);
nand U10429 (N_10429,N_7246,N_8527);
and U10430 (N_10430,N_8114,N_8410);
nor U10431 (N_10431,N_8386,N_8589);
nor U10432 (N_10432,N_8732,N_7316);
nand U10433 (N_10433,N_7611,N_6099);
or U10434 (N_10434,N_7050,N_7633);
nand U10435 (N_10435,N_8797,N_6193);
nor U10436 (N_10436,N_6311,N_8453);
nor U10437 (N_10437,N_6132,N_6757);
nand U10438 (N_10438,N_8235,N_6776);
xnor U10439 (N_10439,N_6783,N_7323);
or U10440 (N_10440,N_7504,N_8521);
and U10441 (N_10441,N_8822,N_7081);
or U10442 (N_10442,N_7669,N_8023);
nand U10443 (N_10443,N_8886,N_8288);
nor U10444 (N_10444,N_6750,N_6891);
or U10445 (N_10445,N_7857,N_8597);
and U10446 (N_10446,N_8977,N_6633);
nor U10447 (N_10447,N_8945,N_8490);
nor U10448 (N_10448,N_6611,N_7169);
or U10449 (N_10449,N_7484,N_7973);
nand U10450 (N_10450,N_6074,N_7733);
xor U10451 (N_10451,N_7114,N_6798);
and U10452 (N_10452,N_8239,N_8312);
xnor U10453 (N_10453,N_6354,N_7494);
xor U10454 (N_10454,N_6876,N_7338);
nand U10455 (N_10455,N_8110,N_7374);
nand U10456 (N_10456,N_8979,N_8085);
and U10457 (N_10457,N_7752,N_7033);
or U10458 (N_10458,N_6028,N_8731);
and U10459 (N_10459,N_8846,N_7049);
nand U10460 (N_10460,N_8321,N_8991);
and U10461 (N_10461,N_6117,N_7806);
xor U10462 (N_10462,N_8025,N_6804);
nand U10463 (N_10463,N_6314,N_6076);
or U10464 (N_10464,N_6795,N_8146);
nand U10465 (N_10465,N_8611,N_6721);
or U10466 (N_10466,N_8489,N_7378);
nor U10467 (N_10467,N_7827,N_7692);
xor U10468 (N_10468,N_8437,N_8249);
nand U10469 (N_10469,N_6934,N_7799);
or U10470 (N_10470,N_8663,N_8988);
and U10471 (N_10471,N_6528,N_7299);
and U10472 (N_10472,N_7748,N_6741);
nand U10473 (N_10473,N_6205,N_6003);
and U10474 (N_10474,N_6793,N_6345);
and U10475 (N_10475,N_6428,N_8667);
xor U10476 (N_10476,N_8247,N_8287);
nand U10477 (N_10477,N_6797,N_8567);
xor U10478 (N_10478,N_6518,N_6975);
nand U10479 (N_10479,N_6877,N_8347);
xnor U10480 (N_10480,N_6413,N_7355);
or U10481 (N_10481,N_6530,N_6246);
nand U10482 (N_10482,N_8516,N_7298);
nor U10483 (N_10483,N_7621,N_8233);
nand U10484 (N_10484,N_6805,N_8853);
nor U10485 (N_10485,N_8519,N_6708);
xnor U10486 (N_10486,N_6897,N_8718);
or U10487 (N_10487,N_6111,N_8499);
xor U10488 (N_10488,N_8987,N_8929);
xnor U10489 (N_10489,N_6760,N_8158);
nand U10490 (N_10490,N_7059,N_8328);
nor U10491 (N_10491,N_6105,N_7178);
or U10492 (N_10492,N_6009,N_8351);
and U10493 (N_10493,N_7929,N_8808);
xnor U10494 (N_10494,N_7202,N_6420);
or U10495 (N_10495,N_7408,N_8583);
or U10496 (N_10496,N_6056,N_8824);
and U10497 (N_10497,N_8958,N_8798);
nor U10498 (N_10498,N_8648,N_8526);
and U10499 (N_10499,N_7117,N_8537);
or U10500 (N_10500,N_6851,N_6257);
xor U10501 (N_10501,N_7877,N_8412);
or U10502 (N_10502,N_6120,N_6856);
nand U10503 (N_10503,N_8722,N_7732);
and U10504 (N_10504,N_6329,N_6663);
or U10505 (N_10505,N_7061,N_6231);
xnor U10506 (N_10506,N_8679,N_8933);
xor U10507 (N_10507,N_6554,N_8373);
or U10508 (N_10508,N_8274,N_7616);
nand U10509 (N_10509,N_6803,N_7344);
nor U10510 (N_10510,N_8707,N_7727);
xnor U10511 (N_10511,N_6206,N_7004);
xor U10512 (N_10512,N_7253,N_6730);
xnor U10513 (N_10513,N_7779,N_6369);
nand U10514 (N_10514,N_7023,N_8344);
nor U10515 (N_10515,N_7841,N_8809);
xnor U10516 (N_10516,N_7724,N_6680);
and U10517 (N_10517,N_6795,N_8752);
nor U10518 (N_10518,N_8022,N_8191);
nor U10519 (N_10519,N_7138,N_6336);
xnor U10520 (N_10520,N_6687,N_8627);
nand U10521 (N_10521,N_8170,N_6060);
nand U10522 (N_10522,N_8228,N_8713);
nand U10523 (N_10523,N_7736,N_7846);
and U10524 (N_10524,N_7699,N_8507);
or U10525 (N_10525,N_7994,N_6698);
and U10526 (N_10526,N_8228,N_6637);
nor U10527 (N_10527,N_6654,N_7258);
or U10528 (N_10528,N_7203,N_6114);
and U10529 (N_10529,N_8814,N_8554);
xnor U10530 (N_10530,N_7205,N_7790);
and U10531 (N_10531,N_7193,N_6938);
and U10532 (N_10532,N_7191,N_8962);
nor U10533 (N_10533,N_7283,N_6721);
and U10534 (N_10534,N_7795,N_7506);
and U10535 (N_10535,N_8002,N_8032);
nor U10536 (N_10536,N_6599,N_7168);
and U10537 (N_10537,N_6076,N_8730);
or U10538 (N_10538,N_7432,N_8576);
and U10539 (N_10539,N_8396,N_7665);
and U10540 (N_10540,N_7193,N_7430);
and U10541 (N_10541,N_6732,N_7533);
nand U10542 (N_10542,N_7874,N_8784);
nor U10543 (N_10543,N_8207,N_6756);
xor U10544 (N_10544,N_7924,N_7816);
or U10545 (N_10545,N_7285,N_7221);
nor U10546 (N_10546,N_7177,N_8637);
nor U10547 (N_10547,N_7354,N_7289);
xnor U10548 (N_10548,N_7192,N_7939);
and U10549 (N_10549,N_8778,N_8214);
nand U10550 (N_10550,N_6084,N_6718);
nor U10551 (N_10551,N_8235,N_8023);
nor U10552 (N_10552,N_8524,N_8014);
or U10553 (N_10553,N_7186,N_6513);
xor U10554 (N_10554,N_7387,N_8557);
and U10555 (N_10555,N_7960,N_7590);
nand U10556 (N_10556,N_7424,N_7388);
or U10557 (N_10557,N_8630,N_7706);
nand U10558 (N_10558,N_7009,N_6403);
and U10559 (N_10559,N_7515,N_6001);
and U10560 (N_10560,N_7293,N_7131);
nand U10561 (N_10561,N_7172,N_6515);
and U10562 (N_10562,N_6328,N_8361);
and U10563 (N_10563,N_7584,N_6153);
or U10564 (N_10564,N_6672,N_6354);
or U10565 (N_10565,N_8832,N_8421);
nand U10566 (N_10566,N_8418,N_8628);
nand U10567 (N_10567,N_7676,N_8627);
and U10568 (N_10568,N_8033,N_8849);
or U10569 (N_10569,N_7828,N_7152);
nand U10570 (N_10570,N_8244,N_6203);
nor U10571 (N_10571,N_7165,N_7081);
nand U10572 (N_10572,N_6477,N_7157);
or U10573 (N_10573,N_6363,N_6758);
nand U10574 (N_10574,N_7589,N_8574);
or U10575 (N_10575,N_8586,N_6751);
nor U10576 (N_10576,N_6016,N_6940);
xor U10577 (N_10577,N_7777,N_8671);
nor U10578 (N_10578,N_8617,N_7119);
and U10579 (N_10579,N_7536,N_8904);
or U10580 (N_10580,N_8422,N_8676);
or U10581 (N_10581,N_6648,N_7183);
and U10582 (N_10582,N_7185,N_7484);
and U10583 (N_10583,N_7139,N_6311);
xnor U10584 (N_10584,N_7366,N_6542);
and U10585 (N_10585,N_6525,N_6228);
xnor U10586 (N_10586,N_8104,N_6601);
xor U10587 (N_10587,N_6976,N_6364);
xor U10588 (N_10588,N_7675,N_6128);
xor U10589 (N_10589,N_7961,N_8290);
or U10590 (N_10590,N_7030,N_8060);
nand U10591 (N_10591,N_6606,N_6254);
or U10592 (N_10592,N_8081,N_7327);
and U10593 (N_10593,N_7080,N_6667);
xnor U10594 (N_10594,N_6989,N_8959);
and U10595 (N_10595,N_6179,N_7292);
nand U10596 (N_10596,N_7762,N_8844);
nor U10597 (N_10597,N_6082,N_6330);
nor U10598 (N_10598,N_6368,N_8134);
and U10599 (N_10599,N_6003,N_7536);
and U10600 (N_10600,N_8955,N_7629);
or U10601 (N_10601,N_6089,N_6349);
xor U10602 (N_10602,N_7401,N_8125);
nor U10603 (N_10603,N_8417,N_8445);
nor U10604 (N_10604,N_8188,N_6633);
and U10605 (N_10605,N_6620,N_8700);
nor U10606 (N_10606,N_8808,N_8699);
and U10607 (N_10607,N_7721,N_8500);
nor U10608 (N_10608,N_6414,N_8234);
and U10609 (N_10609,N_6996,N_6717);
nand U10610 (N_10610,N_6309,N_8317);
nand U10611 (N_10611,N_8276,N_7664);
xor U10612 (N_10612,N_7682,N_8911);
and U10613 (N_10613,N_8896,N_7556);
or U10614 (N_10614,N_7313,N_8489);
nor U10615 (N_10615,N_7495,N_6791);
or U10616 (N_10616,N_6931,N_8234);
xor U10617 (N_10617,N_8927,N_8196);
xnor U10618 (N_10618,N_7339,N_7014);
nand U10619 (N_10619,N_8515,N_6502);
nor U10620 (N_10620,N_7154,N_6551);
xor U10621 (N_10621,N_8077,N_7023);
or U10622 (N_10622,N_8519,N_7842);
nand U10623 (N_10623,N_6616,N_8330);
nand U10624 (N_10624,N_6939,N_8904);
and U10625 (N_10625,N_6839,N_6088);
nand U10626 (N_10626,N_6144,N_7484);
or U10627 (N_10627,N_8804,N_6096);
nand U10628 (N_10628,N_8524,N_7987);
nor U10629 (N_10629,N_7187,N_7288);
nand U10630 (N_10630,N_6520,N_8616);
xor U10631 (N_10631,N_8133,N_6218);
or U10632 (N_10632,N_6433,N_6707);
nand U10633 (N_10633,N_7859,N_7170);
and U10634 (N_10634,N_7990,N_8880);
xnor U10635 (N_10635,N_8241,N_6415);
nor U10636 (N_10636,N_8535,N_6966);
or U10637 (N_10637,N_6281,N_8757);
nor U10638 (N_10638,N_7343,N_8930);
and U10639 (N_10639,N_8128,N_8552);
or U10640 (N_10640,N_6946,N_7035);
xnor U10641 (N_10641,N_6249,N_6243);
and U10642 (N_10642,N_6098,N_7906);
or U10643 (N_10643,N_7651,N_6760);
nor U10644 (N_10644,N_7302,N_8377);
nor U10645 (N_10645,N_7240,N_8899);
and U10646 (N_10646,N_8019,N_8853);
nand U10647 (N_10647,N_8579,N_7556);
or U10648 (N_10648,N_7681,N_8136);
nor U10649 (N_10649,N_6541,N_6380);
or U10650 (N_10650,N_6227,N_7420);
nor U10651 (N_10651,N_8992,N_6876);
xor U10652 (N_10652,N_8098,N_7050);
nand U10653 (N_10653,N_7739,N_8109);
or U10654 (N_10654,N_8564,N_8485);
and U10655 (N_10655,N_6727,N_7276);
nand U10656 (N_10656,N_7855,N_7046);
and U10657 (N_10657,N_8483,N_7126);
xor U10658 (N_10658,N_6236,N_7336);
nand U10659 (N_10659,N_7980,N_7967);
nand U10660 (N_10660,N_6453,N_8330);
and U10661 (N_10661,N_7192,N_8036);
nand U10662 (N_10662,N_6646,N_7300);
or U10663 (N_10663,N_6169,N_6671);
xor U10664 (N_10664,N_8111,N_7551);
xnor U10665 (N_10665,N_8924,N_7418);
or U10666 (N_10666,N_6386,N_7443);
and U10667 (N_10667,N_8810,N_6291);
nand U10668 (N_10668,N_8966,N_6037);
and U10669 (N_10669,N_6119,N_7173);
or U10670 (N_10670,N_6535,N_6450);
and U10671 (N_10671,N_7295,N_6024);
and U10672 (N_10672,N_7372,N_6094);
and U10673 (N_10673,N_7796,N_8183);
xnor U10674 (N_10674,N_7238,N_6177);
or U10675 (N_10675,N_7794,N_7319);
and U10676 (N_10676,N_8169,N_8059);
nand U10677 (N_10677,N_8342,N_8131);
nor U10678 (N_10678,N_7457,N_6661);
or U10679 (N_10679,N_6770,N_7811);
nor U10680 (N_10680,N_7571,N_7616);
nor U10681 (N_10681,N_8899,N_7341);
nand U10682 (N_10682,N_8268,N_8127);
or U10683 (N_10683,N_6335,N_7439);
and U10684 (N_10684,N_7726,N_7014);
nor U10685 (N_10685,N_8463,N_7774);
and U10686 (N_10686,N_7398,N_8993);
xnor U10687 (N_10687,N_7524,N_7618);
and U10688 (N_10688,N_8680,N_7944);
xnor U10689 (N_10689,N_7984,N_7242);
nand U10690 (N_10690,N_8770,N_8071);
nand U10691 (N_10691,N_8163,N_7097);
and U10692 (N_10692,N_7979,N_7576);
nor U10693 (N_10693,N_6766,N_8098);
or U10694 (N_10694,N_7965,N_7381);
xor U10695 (N_10695,N_7147,N_6035);
nand U10696 (N_10696,N_6142,N_8207);
nand U10697 (N_10697,N_8444,N_8717);
or U10698 (N_10698,N_7020,N_6594);
or U10699 (N_10699,N_6876,N_7828);
nor U10700 (N_10700,N_6809,N_7560);
xnor U10701 (N_10701,N_6149,N_6394);
or U10702 (N_10702,N_8447,N_8277);
xnor U10703 (N_10703,N_8649,N_8817);
nand U10704 (N_10704,N_8177,N_7226);
and U10705 (N_10705,N_7135,N_8976);
or U10706 (N_10706,N_7992,N_6609);
or U10707 (N_10707,N_6156,N_8184);
and U10708 (N_10708,N_8458,N_6525);
nor U10709 (N_10709,N_8556,N_8677);
xor U10710 (N_10710,N_7738,N_6745);
xnor U10711 (N_10711,N_6589,N_7201);
nor U10712 (N_10712,N_8981,N_6694);
nand U10713 (N_10713,N_7084,N_8383);
nand U10714 (N_10714,N_8818,N_6221);
or U10715 (N_10715,N_7648,N_7880);
or U10716 (N_10716,N_7202,N_7168);
nand U10717 (N_10717,N_8999,N_7042);
xnor U10718 (N_10718,N_8846,N_6911);
xnor U10719 (N_10719,N_6715,N_8475);
xor U10720 (N_10720,N_8465,N_6065);
and U10721 (N_10721,N_8022,N_7806);
nand U10722 (N_10722,N_8205,N_7200);
nor U10723 (N_10723,N_7785,N_6450);
and U10724 (N_10724,N_7174,N_7206);
xnor U10725 (N_10725,N_8979,N_7173);
and U10726 (N_10726,N_8802,N_8554);
nor U10727 (N_10727,N_6329,N_8958);
nor U10728 (N_10728,N_6312,N_7259);
nor U10729 (N_10729,N_6755,N_7902);
xor U10730 (N_10730,N_8509,N_7170);
or U10731 (N_10731,N_8592,N_7860);
nand U10732 (N_10732,N_6026,N_8123);
nor U10733 (N_10733,N_7641,N_8809);
xor U10734 (N_10734,N_7250,N_7985);
or U10735 (N_10735,N_7295,N_8647);
and U10736 (N_10736,N_8875,N_6334);
and U10737 (N_10737,N_8835,N_6397);
nand U10738 (N_10738,N_8569,N_7328);
or U10739 (N_10739,N_8637,N_8140);
or U10740 (N_10740,N_7982,N_6521);
or U10741 (N_10741,N_8217,N_8008);
nand U10742 (N_10742,N_8609,N_7772);
nand U10743 (N_10743,N_7975,N_6894);
xor U10744 (N_10744,N_7106,N_6326);
nor U10745 (N_10745,N_8097,N_8593);
nor U10746 (N_10746,N_6859,N_8459);
and U10747 (N_10747,N_7976,N_7664);
and U10748 (N_10748,N_7464,N_8187);
nor U10749 (N_10749,N_8637,N_8679);
xnor U10750 (N_10750,N_6799,N_7161);
nor U10751 (N_10751,N_8620,N_8165);
and U10752 (N_10752,N_6655,N_7338);
xnor U10753 (N_10753,N_6172,N_7119);
nand U10754 (N_10754,N_7849,N_7831);
or U10755 (N_10755,N_8508,N_8890);
xnor U10756 (N_10756,N_8333,N_8055);
xor U10757 (N_10757,N_7037,N_8061);
xor U10758 (N_10758,N_7900,N_8454);
and U10759 (N_10759,N_7984,N_8342);
or U10760 (N_10760,N_8005,N_6441);
nand U10761 (N_10761,N_6935,N_8520);
nor U10762 (N_10762,N_6548,N_7372);
or U10763 (N_10763,N_8902,N_8288);
nor U10764 (N_10764,N_7185,N_8999);
xnor U10765 (N_10765,N_7638,N_7964);
nor U10766 (N_10766,N_6546,N_8562);
nand U10767 (N_10767,N_7240,N_7231);
nor U10768 (N_10768,N_7763,N_7297);
xnor U10769 (N_10769,N_6351,N_8335);
xnor U10770 (N_10770,N_8001,N_7184);
or U10771 (N_10771,N_6309,N_6396);
xor U10772 (N_10772,N_7640,N_7325);
and U10773 (N_10773,N_8650,N_8769);
nand U10774 (N_10774,N_8217,N_8873);
nand U10775 (N_10775,N_8916,N_6556);
nand U10776 (N_10776,N_7076,N_6833);
nor U10777 (N_10777,N_6835,N_6862);
nor U10778 (N_10778,N_8262,N_6639);
xnor U10779 (N_10779,N_7075,N_8816);
and U10780 (N_10780,N_6659,N_7424);
nor U10781 (N_10781,N_7021,N_6394);
and U10782 (N_10782,N_6442,N_6403);
or U10783 (N_10783,N_7719,N_8288);
or U10784 (N_10784,N_6347,N_7826);
nand U10785 (N_10785,N_8232,N_6622);
nor U10786 (N_10786,N_7205,N_6390);
xnor U10787 (N_10787,N_7112,N_7626);
and U10788 (N_10788,N_7716,N_7326);
and U10789 (N_10789,N_6387,N_7319);
xor U10790 (N_10790,N_7463,N_8553);
xnor U10791 (N_10791,N_7066,N_8823);
xor U10792 (N_10792,N_7277,N_6902);
nand U10793 (N_10793,N_8618,N_7056);
xor U10794 (N_10794,N_8046,N_6081);
nor U10795 (N_10795,N_7539,N_8489);
nand U10796 (N_10796,N_6233,N_7934);
xnor U10797 (N_10797,N_7321,N_7256);
or U10798 (N_10798,N_7552,N_8053);
nor U10799 (N_10799,N_8302,N_8585);
nand U10800 (N_10800,N_7043,N_7720);
and U10801 (N_10801,N_6996,N_8257);
or U10802 (N_10802,N_7505,N_7371);
or U10803 (N_10803,N_6363,N_6541);
nor U10804 (N_10804,N_7286,N_8457);
and U10805 (N_10805,N_6244,N_7470);
and U10806 (N_10806,N_8636,N_6910);
nor U10807 (N_10807,N_6120,N_8075);
nor U10808 (N_10808,N_6841,N_8283);
nor U10809 (N_10809,N_7303,N_8250);
nand U10810 (N_10810,N_6315,N_8348);
xor U10811 (N_10811,N_7476,N_6782);
nand U10812 (N_10812,N_7424,N_8313);
or U10813 (N_10813,N_8862,N_8126);
and U10814 (N_10814,N_6660,N_7881);
and U10815 (N_10815,N_7683,N_7404);
or U10816 (N_10816,N_8616,N_7941);
nand U10817 (N_10817,N_6705,N_7514);
and U10818 (N_10818,N_6588,N_7429);
or U10819 (N_10819,N_6900,N_6158);
and U10820 (N_10820,N_7751,N_7305);
or U10821 (N_10821,N_6576,N_7220);
xnor U10822 (N_10822,N_7792,N_6010);
nand U10823 (N_10823,N_6058,N_6184);
or U10824 (N_10824,N_8039,N_7639);
xor U10825 (N_10825,N_7058,N_7772);
nor U10826 (N_10826,N_6933,N_7298);
or U10827 (N_10827,N_7474,N_8957);
and U10828 (N_10828,N_6346,N_8903);
and U10829 (N_10829,N_6937,N_7417);
or U10830 (N_10830,N_7751,N_8162);
and U10831 (N_10831,N_8483,N_7564);
xor U10832 (N_10832,N_7081,N_7875);
and U10833 (N_10833,N_7626,N_8951);
and U10834 (N_10834,N_6395,N_8504);
or U10835 (N_10835,N_8892,N_7404);
xnor U10836 (N_10836,N_7967,N_7209);
and U10837 (N_10837,N_8719,N_6357);
or U10838 (N_10838,N_6838,N_8580);
and U10839 (N_10839,N_6952,N_6181);
nand U10840 (N_10840,N_6089,N_6859);
and U10841 (N_10841,N_8663,N_8915);
nand U10842 (N_10842,N_8118,N_7033);
xnor U10843 (N_10843,N_7202,N_8113);
nand U10844 (N_10844,N_6074,N_6335);
and U10845 (N_10845,N_7029,N_8384);
and U10846 (N_10846,N_7505,N_7664);
or U10847 (N_10847,N_7968,N_8551);
nor U10848 (N_10848,N_7774,N_6548);
xnor U10849 (N_10849,N_6331,N_8470);
and U10850 (N_10850,N_7905,N_7681);
xor U10851 (N_10851,N_8651,N_8993);
nand U10852 (N_10852,N_6772,N_7255);
nor U10853 (N_10853,N_7485,N_7536);
nor U10854 (N_10854,N_8984,N_6147);
nor U10855 (N_10855,N_7473,N_7236);
nand U10856 (N_10856,N_7115,N_7386);
nor U10857 (N_10857,N_8907,N_8936);
nor U10858 (N_10858,N_6489,N_7070);
nor U10859 (N_10859,N_7693,N_7106);
or U10860 (N_10860,N_7198,N_8982);
nor U10861 (N_10861,N_7424,N_6720);
nor U10862 (N_10862,N_6145,N_6535);
and U10863 (N_10863,N_6108,N_6889);
nor U10864 (N_10864,N_7976,N_6803);
or U10865 (N_10865,N_6356,N_8579);
or U10866 (N_10866,N_7978,N_6796);
nand U10867 (N_10867,N_6599,N_6578);
and U10868 (N_10868,N_6910,N_7442);
nand U10869 (N_10869,N_6229,N_6874);
nor U10870 (N_10870,N_8595,N_8719);
nor U10871 (N_10871,N_8092,N_8275);
nor U10872 (N_10872,N_7253,N_7230);
or U10873 (N_10873,N_7028,N_7728);
or U10874 (N_10874,N_6181,N_7906);
and U10875 (N_10875,N_7094,N_8279);
nor U10876 (N_10876,N_7158,N_6965);
and U10877 (N_10877,N_7223,N_7402);
or U10878 (N_10878,N_6935,N_6440);
and U10879 (N_10879,N_6794,N_8858);
nand U10880 (N_10880,N_8568,N_7629);
or U10881 (N_10881,N_6516,N_7952);
xnor U10882 (N_10882,N_8251,N_8958);
or U10883 (N_10883,N_7259,N_8286);
nor U10884 (N_10884,N_8262,N_8575);
nand U10885 (N_10885,N_7910,N_6360);
nand U10886 (N_10886,N_8888,N_8170);
nand U10887 (N_10887,N_7244,N_6256);
nand U10888 (N_10888,N_8689,N_8674);
xor U10889 (N_10889,N_7553,N_8731);
or U10890 (N_10890,N_8088,N_8579);
or U10891 (N_10891,N_7091,N_8573);
nor U10892 (N_10892,N_6948,N_8496);
nor U10893 (N_10893,N_6273,N_6553);
nand U10894 (N_10894,N_8222,N_7889);
xnor U10895 (N_10895,N_8909,N_7319);
and U10896 (N_10896,N_8676,N_6129);
and U10897 (N_10897,N_8123,N_8599);
or U10898 (N_10898,N_8988,N_7859);
nand U10899 (N_10899,N_7844,N_7036);
nand U10900 (N_10900,N_8009,N_8724);
xor U10901 (N_10901,N_8195,N_6283);
and U10902 (N_10902,N_6644,N_8322);
nor U10903 (N_10903,N_7307,N_8886);
xnor U10904 (N_10904,N_7649,N_8358);
or U10905 (N_10905,N_6287,N_8529);
nand U10906 (N_10906,N_8243,N_6520);
or U10907 (N_10907,N_8437,N_8420);
nor U10908 (N_10908,N_8206,N_8654);
nand U10909 (N_10909,N_8665,N_8935);
xnor U10910 (N_10910,N_7210,N_7311);
nand U10911 (N_10911,N_7142,N_8904);
nand U10912 (N_10912,N_8695,N_8107);
or U10913 (N_10913,N_7189,N_7701);
xnor U10914 (N_10914,N_7273,N_6412);
nor U10915 (N_10915,N_7175,N_8253);
and U10916 (N_10916,N_8220,N_8160);
xor U10917 (N_10917,N_8950,N_7015);
nor U10918 (N_10918,N_6559,N_6188);
and U10919 (N_10919,N_8433,N_6964);
and U10920 (N_10920,N_6526,N_7854);
or U10921 (N_10921,N_6654,N_6876);
or U10922 (N_10922,N_7285,N_6403);
nand U10923 (N_10923,N_6522,N_7764);
nor U10924 (N_10924,N_6807,N_6870);
xor U10925 (N_10925,N_7916,N_7462);
nand U10926 (N_10926,N_6232,N_7766);
xor U10927 (N_10927,N_6149,N_7140);
nand U10928 (N_10928,N_6670,N_7676);
xor U10929 (N_10929,N_6637,N_8826);
nand U10930 (N_10930,N_6433,N_6051);
and U10931 (N_10931,N_8605,N_8263);
nor U10932 (N_10932,N_8895,N_8821);
and U10933 (N_10933,N_7671,N_8924);
and U10934 (N_10934,N_6054,N_6660);
nand U10935 (N_10935,N_8289,N_8537);
and U10936 (N_10936,N_6706,N_7324);
or U10937 (N_10937,N_7558,N_6904);
nor U10938 (N_10938,N_6528,N_6620);
xor U10939 (N_10939,N_8084,N_8845);
xnor U10940 (N_10940,N_6494,N_6762);
and U10941 (N_10941,N_8766,N_8158);
nand U10942 (N_10942,N_6297,N_8021);
nor U10943 (N_10943,N_8379,N_7220);
xor U10944 (N_10944,N_6014,N_7316);
or U10945 (N_10945,N_7707,N_8931);
and U10946 (N_10946,N_8686,N_8892);
xor U10947 (N_10947,N_8460,N_7753);
and U10948 (N_10948,N_6227,N_8517);
and U10949 (N_10949,N_7323,N_8367);
nand U10950 (N_10950,N_8782,N_6359);
xnor U10951 (N_10951,N_7810,N_6129);
nand U10952 (N_10952,N_8581,N_7284);
xnor U10953 (N_10953,N_8337,N_6014);
xnor U10954 (N_10954,N_8578,N_7511);
xor U10955 (N_10955,N_6449,N_7053);
and U10956 (N_10956,N_8153,N_7933);
and U10957 (N_10957,N_8364,N_6292);
nand U10958 (N_10958,N_6584,N_8165);
xor U10959 (N_10959,N_6975,N_6591);
nor U10960 (N_10960,N_7086,N_6809);
nand U10961 (N_10961,N_8940,N_6503);
or U10962 (N_10962,N_6676,N_6127);
or U10963 (N_10963,N_7755,N_7198);
xnor U10964 (N_10964,N_8834,N_8657);
xor U10965 (N_10965,N_8956,N_8079);
xnor U10966 (N_10966,N_6173,N_7079);
xnor U10967 (N_10967,N_8081,N_8993);
nand U10968 (N_10968,N_6415,N_8894);
xnor U10969 (N_10969,N_7526,N_6141);
and U10970 (N_10970,N_6663,N_6531);
xnor U10971 (N_10971,N_7902,N_8580);
nand U10972 (N_10972,N_6151,N_8203);
nand U10973 (N_10973,N_8785,N_6789);
nor U10974 (N_10974,N_6840,N_8706);
xnor U10975 (N_10975,N_8350,N_8718);
nand U10976 (N_10976,N_7362,N_6215);
nor U10977 (N_10977,N_6411,N_7449);
or U10978 (N_10978,N_7859,N_7638);
and U10979 (N_10979,N_7322,N_8755);
xor U10980 (N_10980,N_7333,N_6306);
nand U10981 (N_10981,N_7080,N_8180);
or U10982 (N_10982,N_6462,N_6992);
and U10983 (N_10983,N_8285,N_6516);
xnor U10984 (N_10984,N_7263,N_8772);
xor U10985 (N_10985,N_7766,N_8385);
xor U10986 (N_10986,N_8448,N_8995);
nor U10987 (N_10987,N_8657,N_6566);
nand U10988 (N_10988,N_6284,N_8680);
and U10989 (N_10989,N_8803,N_6590);
or U10990 (N_10990,N_7460,N_7187);
nand U10991 (N_10991,N_8961,N_6353);
nor U10992 (N_10992,N_7296,N_6163);
xor U10993 (N_10993,N_6277,N_6679);
nand U10994 (N_10994,N_7786,N_8074);
nand U10995 (N_10995,N_7176,N_6627);
or U10996 (N_10996,N_6907,N_6611);
or U10997 (N_10997,N_7696,N_8377);
and U10998 (N_10998,N_7330,N_8656);
nor U10999 (N_10999,N_6793,N_7954);
xor U11000 (N_11000,N_6049,N_7993);
xnor U11001 (N_11001,N_7899,N_8612);
xnor U11002 (N_11002,N_6428,N_6940);
xor U11003 (N_11003,N_6526,N_6903);
nor U11004 (N_11004,N_6549,N_8414);
xnor U11005 (N_11005,N_6731,N_8687);
or U11006 (N_11006,N_7610,N_7353);
xor U11007 (N_11007,N_6399,N_7744);
or U11008 (N_11008,N_7584,N_6718);
xnor U11009 (N_11009,N_7240,N_8126);
or U11010 (N_11010,N_8560,N_7933);
or U11011 (N_11011,N_7981,N_7647);
and U11012 (N_11012,N_6153,N_6331);
and U11013 (N_11013,N_6503,N_7153);
xnor U11014 (N_11014,N_8514,N_6790);
or U11015 (N_11015,N_8527,N_7723);
or U11016 (N_11016,N_6448,N_7130);
nand U11017 (N_11017,N_7612,N_7094);
xor U11018 (N_11018,N_6580,N_7537);
and U11019 (N_11019,N_6568,N_7560);
xor U11020 (N_11020,N_7655,N_8721);
nand U11021 (N_11021,N_7099,N_8758);
nor U11022 (N_11022,N_6903,N_7515);
nand U11023 (N_11023,N_8787,N_6501);
nor U11024 (N_11024,N_6224,N_6766);
nor U11025 (N_11025,N_6365,N_6273);
or U11026 (N_11026,N_7194,N_7169);
nor U11027 (N_11027,N_7878,N_6452);
and U11028 (N_11028,N_6491,N_7022);
or U11029 (N_11029,N_6922,N_7422);
or U11030 (N_11030,N_7287,N_6490);
xnor U11031 (N_11031,N_7323,N_6973);
nor U11032 (N_11032,N_6957,N_8009);
or U11033 (N_11033,N_6238,N_6450);
nor U11034 (N_11034,N_7299,N_7689);
nand U11035 (N_11035,N_8107,N_7281);
nor U11036 (N_11036,N_7521,N_8075);
nand U11037 (N_11037,N_8325,N_6988);
nand U11038 (N_11038,N_7895,N_7548);
nor U11039 (N_11039,N_8781,N_6138);
nor U11040 (N_11040,N_6772,N_6391);
xor U11041 (N_11041,N_7809,N_8965);
and U11042 (N_11042,N_7592,N_6860);
xor U11043 (N_11043,N_6108,N_8227);
or U11044 (N_11044,N_8081,N_7620);
nand U11045 (N_11045,N_8900,N_7040);
nor U11046 (N_11046,N_7021,N_8656);
nand U11047 (N_11047,N_7109,N_8519);
nor U11048 (N_11048,N_8869,N_7501);
nand U11049 (N_11049,N_6231,N_7152);
xnor U11050 (N_11050,N_7011,N_8748);
nor U11051 (N_11051,N_7235,N_8946);
and U11052 (N_11052,N_7669,N_6167);
xor U11053 (N_11053,N_8131,N_6780);
nand U11054 (N_11054,N_8481,N_6992);
and U11055 (N_11055,N_8234,N_6840);
xor U11056 (N_11056,N_7915,N_6505);
and U11057 (N_11057,N_7102,N_7717);
xor U11058 (N_11058,N_8268,N_6871);
nand U11059 (N_11059,N_6345,N_7649);
nor U11060 (N_11060,N_6316,N_8705);
and U11061 (N_11061,N_7560,N_7467);
nor U11062 (N_11062,N_6196,N_6610);
and U11063 (N_11063,N_8699,N_8562);
nor U11064 (N_11064,N_8549,N_6606);
xor U11065 (N_11065,N_6907,N_7433);
or U11066 (N_11066,N_6757,N_7284);
nand U11067 (N_11067,N_8513,N_8014);
and U11068 (N_11068,N_7603,N_7688);
xnor U11069 (N_11069,N_7450,N_6550);
nor U11070 (N_11070,N_7704,N_7020);
xnor U11071 (N_11071,N_6812,N_7626);
nand U11072 (N_11072,N_6207,N_8561);
or U11073 (N_11073,N_6828,N_8080);
nor U11074 (N_11074,N_6339,N_6219);
nand U11075 (N_11075,N_8353,N_7865);
and U11076 (N_11076,N_8215,N_7239);
xor U11077 (N_11077,N_6057,N_8515);
nor U11078 (N_11078,N_7891,N_8758);
nor U11079 (N_11079,N_6449,N_8642);
and U11080 (N_11080,N_6781,N_6885);
nand U11081 (N_11081,N_7573,N_7729);
and U11082 (N_11082,N_7899,N_8263);
xor U11083 (N_11083,N_8256,N_8612);
nand U11084 (N_11084,N_8699,N_8277);
nor U11085 (N_11085,N_7673,N_6362);
or U11086 (N_11086,N_6898,N_6542);
xnor U11087 (N_11087,N_8886,N_7490);
or U11088 (N_11088,N_6936,N_8296);
and U11089 (N_11089,N_7772,N_8658);
nand U11090 (N_11090,N_7890,N_7030);
nor U11091 (N_11091,N_8037,N_6894);
or U11092 (N_11092,N_7820,N_7156);
nand U11093 (N_11093,N_8024,N_7813);
and U11094 (N_11094,N_7450,N_8841);
or U11095 (N_11095,N_6419,N_6855);
nand U11096 (N_11096,N_6731,N_6313);
nor U11097 (N_11097,N_6377,N_6182);
nor U11098 (N_11098,N_6523,N_8991);
or U11099 (N_11099,N_7994,N_7419);
xor U11100 (N_11100,N_7336,N_6549);
and U11101 (N_11101,N_6669,N_8233);
xor U11102 (N_11102,N_6409,N_8599);
or U11103 (N_11103,N_7575,N_7780);
nor U11104 (N_11104,N_7215,N_6701);
or U11105 (N_11105,N_6499,N_6364);
and U11106 (N_11106,N_8344,N_8353);
nor U11107 (N_11107,N_8424,N_6948);
or U11108 (N_11108,N_6326,N_8986);
xor U11109 (N_11109,N_8873,N_8554);
and U11110 (N_11110,N_6768,N_6635);
xnor U11111 (N_11111,N_8870,N_7670);
nand U11112 (N_11112,N_8168,N_8216);
and U11113 (N_11113,N_7664,N_8765);
or U11114 (N_11114,N_6149,N_8566);
and U11115 (N_11115,N_6585,N_6401);
xor U11116 (N_11116,N_8479,N_8569);
and U11117 (N_11117,N_8883,N_8314);
or U11118 (N_11118,N_7318,N_8304);
xnor U11119 (N_11119,N_7175,N_8480);
and U11120 (N_11120,N_6907,N_7027);
nand U11121 (N_11121,N_6009,N_6178);
and U11122 (N_11122,N_6717,N_6725);
nor U11123 (N_11123,N_6299,N_8064);
or U11124 (N_11124,N_7035,N_8931);
nor U11125 (N_11125,N_6374,N_6208);
nor U11126 (N_11126,N_6465,N_8439);
nor U11127 (N_11127,N_8644,N_7817);
or U11128 (N_11128,N_7309,N_8345);
nor U11129 (N_11129,N_6064,N_8542);
nor U11130 (N_11130,N_6525,N_8939);
nor U11131 (N_11131,N_6175,N_8834);
nor U11132 (N_11132,N_7149,N_8556);
nand U11133 (N_11133,N_7105,N_6614);
nand U11134 (N_11134,N_7287,N_7670);
nor U11135 (N_11135,N_8952,N_7777);
and U11136 (N_11136,N_8016,N_7769);
and U11137 (N_11137,N_6014,N_7184);
xor U11138 (N_11138,N_7425,N_7936);
xor U11139 (N_11139,N_8690,N_8378);
or U11140 (N_11140,N_8035,N_6937);
and U11141 (N_11141,N_6663,N_7111);
nand U11142 (N_11142,N_6418,N_8233);
nand U11143 (N_11143,N_6809,N_7977);
nand U11144 (N_11144,N_8431,N_7008);
xnor U11145 (N_11145,N_8208,N_8571);
nor U11146 (N_11146,N_6056,N_6975);
nor U11147 (N_11147,N_7016,N_8381);
and U11148 (N_11148,N_7798,N_6613);
nand U11149 (N_11149,N_8151,N_7468);
and U11150 (N_11150,N_7632,N_7728);
nor U11151 (N_11151,N_6351,N_8104);
or U11152 (N_11152,N_6691,N_6809);
or U11153 (N_11153,N_7700,N_7835);
and U11154 (N_11154,N_7033,N_8060);
and U11155 (N_11155,N_8757,N_8861);
or U11156 (N_11156,N_6237,N_7193);
nor U11157 (N_11157,N_8082,N_8108);
nor U11158 (N_11158,N_8210,N_7045);
nor U11159 (N_11159,N_7791,N_6559);
xor U11160 (N_11160,N_6795,N_7488);
and U11161 (N_11161,N_6548,N_7462);
or U11162 (N_11162,N_8910,N_7806);
nor U11163 (N_11163,N_6393,N_6026);
xor U11164 (N_11164,N_6561,N_8741);
nand U11165 (N_11165,N_6154,N_7527);
nor U11166 (N_11166,N_6849,N_8819);
xnor U11167 (N_11167,N_8730,N_7307);
and U11168 (N_11168,N_8007,N_6624);
nand U11169 (N_11169,N_6421,N_7861);
nand U11170 (N_11170,N_7478,N_8233);
nand U11171 (N_11171,N_6258,N_7332);
and U11172 (N_11172,N_6071,N_7345);
or U11173 (N_11173,N_8774,N_7316);
nor U11174 (N_11174,N_8996,N_6250);
xor U11175 (N_11175,N_6729,N_8954);
and U11176 (N_11176,N_8580,N_8431);
xor U11177 (N_11177,N_6253,N_6456);
xor U11178 (N_11178,N_6020,N_7355);
nor U11179 (N_11179,N_8145,N_6077);
nand U11180 (N_11180,N_6229,N_8574);
and U11181 (N_11181,N_8850,N_6300);
xor U11182 (N_11182,N_8531,N_8037);
nand U11183 (N_11183,N_7880,N_6545);
and U11184 (N_11184,N_7083,N_8110);
nor U11185 (N_11185,N_8075,N_8326);
xor U11186 (N_11186,N_6809,N_7604);
nor U11187 (N_11187,N_8995,N_6161);
nand U11188 (N_11188,N_8561,N_8960);
or U11189 (N_11189,N_6403,N_8511);
or U11190 (N_11190,N_6423,N_7864);
nand U11191 (N_11191,N_7877,N_6008);
or U11192 (N_11192,N_7986,N_8572);
nand U11193 (N_11193,N_6696,N_6119);
or U11194 (N_11194,N_6469,N_6068);
or U11195 (N_11195,N_7039,N_6459);
xnor U11196 (N_11196,N_7230,N_6777);
and U11197 (N_11197,N_6728,N_8948);
xnor U11198 (N_11198,N_6816,N_8859);
and U11199 (N_11199,N_7021,N_7601);
nor U11200 (N_11200,N_8927,N_8655);
and U11201 (N_11201,N_8071,N_6586);
xnor U11202 (N_11202,N_8387,N_7187);
or U11203 (N_11203,N_6908,N_8410);
nor U11204 (N_11204,N_6697,N_8001);
nand U11205 (N_11205,N_7589,N_7443);
and U11206 (N_11206,N_8596,N_8990);
and U11207 (N_11207,N_7731,N_6194);
nor U11208 (N_11208,N_7667,N_7072);
and U11209 (N_11209,N_8749,N_7197);
nand U11210 (N_11210,N_6901,N_6584);
and U11211 (N_11211,N_8000,N_7870);
xor U11212 (N_11212,N_6527,N_7799);
nor U11213 (N_11213,N_6626,N_8906);
xnor U11214 (N_11214,N_7815,N_8462);
and U11215 (N_11215,N_7154,N_8969);
nand U11216 (N_11216,N_7585,N_6372);
or U11217 (N_11217,N_8107,N_7018);
nand U11218 (N_11218,N_7768,N_8155);
and U11219 (N_11219,N_7619,N_7707);
nor U11220 (N_11220,N_7781,N_8577);
and U11221 (N_11221,N_8351,N_7690);
xnor U11222 (N_11222,N_7940,N_8632);
xor U11223 (N_11223,N_7915,N_8763);
xor U11224 (N_11224,N_7837,N_8765);
xor U11225 (N_11225,N_7204,N_7762);
or U11226 (N_11226,N_8940,N_7569);
xnor U11227 (N_11227,N_6657,N_6223);
or U11228 (N_11228,N_6862,N_7991);
nand U11229 (N_11229,N_6691,N_8939);
or U11230 (N_11230,N_8773,N_6721);
nand U11231 (N_11231,N_7153,N_8439);
xnor U11232 (N_11232,N_8376,N_6990);
and U11233 (N_11233,N_6121,N_6066);
nor U11234 (N_11234,N_6252,N_7328);
or U11235 (N_11235,N_8316,N_6930);
or U11236 (N_11236,N_6495,N_8529);
and U11237 (N_11237,N_7517,N_8972);
or U11238 (N_11238,N_8746,N_8722);
xnor U11239 (N_11239,N_8111,N_6066);
and U11240 (N_11240,N_7791,N_8035);
xor U11241 (N_11241,N_7568,N_8334);
or U11242 (N_11242,N_6262,N_6258);
and U11243 (N_11243,N_7728,N_8038);
or U11244 (N_11244,N_7424,N_7833);
xnor U11245 (N_11245,N_7975,N_6514);
and U11246 (N_11246,N_6848,N_8877);
xor U11247 (N_11247,N_7369,N_7446);
and U11248 (N_11248,N_7312,N_7151);
nor U11249 (N_11249,N_7008,N_7472);
or U11250 (N_11250,N_7890,N_6246);
nor U11251 (N_11251,N_6679,N_8311);
xnor U11252 (N_11252,N_8453,N_6455);
nand U11253 (N_11253,N_8965,N_6946);
xor U11254 (N_11254,N_7341,N_6382);
xor U11255 (N_11255,N_7471,N_8139);
or U11256 (N_11256,N_6157,N_7416);
nand U11257 (N_11257,N_8905,N_6597);
and U11258 (N_11258,N_6913,N_6495);
xnor U11259 (N_11259,N_6723,N_6000);
nor U11260 (N_11260,N_7992,N_8150);
nor U11261 (N_11261,N_7263,N_8288);
or U11262 (N_11262,N_8492,N_8886);
and U11263 (N_11263,N_6706,N_8622);
and U11264 (N_11264,N_6293,N_6934);
and U11265 (N_11265,N_7767,N_7540);
nand U11266 (N_11266,N_8209,N_8018);
and U11267 (N_11267,N_8668,N_8009);
nor U11268 (N_11268,N_7775,N_6748);
nand U11269 (N_11269,N_7639,N_8105);
and U11270 (N_11270,N_7657,N_8795);
or U11271 (N_11271,N_7861,N_7754);
nand U11272 (N_11272,N_8287,N_6730);
or U11273 (N_11273,N_6717,N_6221);
nand U11274 (N_11274,N_7417,N_8987);
xnor U11275 (N_11275,N_6900,N_7031);
nand U11276 (N_11276,N_7861,N_7660);
nor U11277 (N_11277,N_7640,N_6355);
nor U11278 (N_11278,N_7788,N_6857);
and U11279 (N_11279,N_8780,N_6753);
or U11280 (N_11280,N_8440,N_8683);
nand U11281 (N_11281,N_6923,N_6180);
nand U11282 (N_11282,N_6541,N_8337);
and U11283 (N_11283,N_6322,N_6554);
and U11284 (N_11284,N_6401,N_6042);
and U11285 (N_11285,N_6358,N_7328);
and U11286 (N_11286,N_7192,N_6948);
xnor U11287 (N_11287,N_6296,N_7089);
nor U11288 (N_11288,N_6246,N_7786);
and U11289 (N_11289,N_8189,N_6336);
or U11290 (N_11290,N_7759,N_7738);
or U11291 (N_11291,N_8876,N_6860);
and U11292 (N_11292,N_7344,N_8433);
nand U11293 (N_11293,N_8851,N_7175);
and U11294 (N_11294,N_8829,N_8768);
nand U11295 (N_11295,N_6785,N_7969);
or U11296 (N_11296,N_8135,N_7497);
and U11297 (N_11297,N_8521,N_8701);
nand U11298 (N_11298,N_6245,N_7408);
and U11299 (N_11299,N_7399,N_6149);
nor U11300 (N_11300,N_7979,N_8231);
and U11301 (N_11301,N_7989,N_6636);
and U11302 (N_11302,N_6137,N_7447);
xor U11303 (N_11303,N_8292,N_8573);
nand U11304 (N_11304,N_6370,N_6747);
or U11305 (N_11305,N_6002,N_7208);
and U11306 (N_11306,N_6980,N_6826);
and U11307 (N_11307,N_8143,N_7187);
or U11308 (N_11308,N_6481,N_7609);
xor U11309 (N_11309,N_7974,N_8286);
xnor U11310 (N_11310,N_7199,N_8308);
nor U11311 (N_11311,N_8264,N_7687);
nor U11312 (N_11312,N_8456,N_8065);
and U11313 (N_11313,N_8340,N_6046);
nor U11314 (N_11314,N_7008,N_7405);
and U11315 (N_11315,N_8145,N_7627);
xnor U11316 (N_11316,N_7879,N_6737);
nand U11317 (N_11317,N_7791,N_8160);
or U11318 (N_11318,N_8583,N_6166);
xor U11319 (N_11319,N_6302,N_6307);
nor U11320 (N_11320,N_6028,N_6995);
xnor U11321 (N_11321,N_6653,N_6594);
nand U11322 (N_11322,N_8652,N_6659);
nor U11323 (N_11323,N_6828,N_8933);
and U11324 (N_11324,N_6362,N_6025);
nor U11325 (N_11325,N_8053,N_7930);
xnor U11326 (N_11326,N_8087,N_7146);
nor U11327 (N_11327,N_8323,N_8262);
nor U11328 (N_11328,N_7674,N_7121);
nand U11329 (N_11329,N_8939,N_6052);
and U11330 (N_11330,N_7392,N_7987);
and U11331 (N_11331,N_8163,N_7954);
xnor U11332 (N_11332,N_7091,N_6041);
nand U11333 (N_11333,N_8690,N_8666);
xnor U11334 (N_11334,N_6386,N_8186);
and U11335 (N_11335,N_6784,N_7868);
nand U11336 (N_11336,N_8365,N_6299);
and U11337 (N_11337,N_7183,N_8056);
nand U11338 (N_11338,N_6667,N_8143);
and U11339 (N_11339,N_6868,N_8575);
and U11340 (N_11340,N_7960,N_8293);
xnor U11341 (N_11341,N_6164,N_6769);
and U11342 (N_11342,N_6819,N_7124);
nor U11343 (N_11343,N_8737,N_8849);
nor U11344 (N_11344,N_7323,N_7888);
nor U11345 (N_11345,N_8490,N_6707);
nand U11346 (N_11346,N_6660,N_8248);
and U11347 (N_11347,N_6393,N_8548);
and U11348 (N_11348,N_7461,N_8253);
nand U11349 (N_11349,N_6372,N_6007);
nor U11350 (N_11350,N_6113,N_7429);
nor U11351 (N_11351,N_7730,N_6940);
or U11352 (N_11352,N_8091,N_8160);
nor U11353 (N_11353,N_8711,N_8241);
or U11354 (N_11354,N_7807,N_6755);
xnor U11355 (N_11355,N_6588,N_6932);
xnor U11356 (N_11356,N_6278,N_7770);
and U11357 (N_11357,N_7585,N_7998);
nor U11358 (N_11358,N_8009,N_8194);
nor U11359 (N_11359,N_8594,N_8206);
xnor U11360 (N_11360,N_8919,N_8684);
nand U11361 (N_11361,N_7992,N_6142);
nor U11362 (N_11362,N_6575,N_8421);
or U11363 (N_11363,N_6292,N_7838);
or U11364 (N_11364,N_6451,N_6404);
nor U11365 (N_11365,N_8411,N_7225);
and U11366 (N_11366,N_7349,N_7888);
or U11367 (N_11367,N_7605,N_8619);
or U11368 (N_11368,N_6375,N_6167);
nand U11369 (N_11369,N_8624,N_7497);
and U11370 (N_11370,N_7037,N_8367);
and U11371 (N_11371,N_7925,N_7473);
or U11372 (N_11372,N_7914,N_6816);
xnor U11373 (N_11373,N_7447,N_7537);
xnor U11374 (N_11374,N_7298,N_8322);
and U11375 (N_11375,N_8071,N_7211);
nand U11376 (N_11376,N_6785,N_6364);
and U11377 (N_11377,N_8594,N_6681);
nand U11378 (N_11378,N_8624,N_8712);
xor U11379 (N_11379,N_7454,N_8558);
nor U11380 (N_11380,N_7699,N_7768);
and U11381 (N_11381,N_7348,N_8959);
xor U11382 (N_11382,N_8737,N_8607);
xnor U11383 (N_11383,N_7677,N_7057);
nor U11384 (N_11384,N_6993,N_6497);
xor U11385 (N_11385,N_6536,N_7749);
xor U11386 (N_11386,N_8682,N_7139);
xnor U11387 (N_11387,N_8669,N_6479);
nor U11388 (N_11388,N_8515,N_8865);
or U11389 (N_11389,N_6270,N_7824);
and U11390 (N_11390,N_6297,N_8053);
nor U11391 (N_11391,N_7185,N_7960);
nand U11392 (N_11392,N_7493,N_8970);
xor U11393 (N_11393,N_6646,N_6883);
nor U11394 (N_11394,N_6763,N_7756);
xor U11395 (N_11395,N_7574,N_8740);
nand U11396 (N_11396,N_7088,N_6907);
and U11397 (N_11397,N_6808,N_8758);
nor U11398 (N_11398,N_8922,N_7251);
xor U11399 (N_11399,N_7061,N_7279);
nand U11400 (N_11400,N_8551,N_7732);
or U11401 (N_11401,N_6161,N_7049);
nand U11402 (N_11402,N_8356,N_8091);
xor U11403 (N_11403,N_6325,N_8204);
or U11404 (N_11404,N_7061,N_8332);
and U11405 (N_11405,N_8693,N_7893);
xnor U11406 (N_11406,N_8117,N_6421);
and U11407 (N_11407,N_7664,N_7831);
and U11408 (N_11408,N_6291,N_8156);
and U11409 (N_11409,N_6699,N_7886);
nand U11410 (N_11410,N_7476,N_7539);
or U11411 (N_11411,N_6134,N_8241);
or U11412 (N_11412,N_8060,N_6726);
xnor U11413 (N_11413,N_6482,N_7939);
nor U11414 (N_11414,N_7746,N_6088);
xnor U11415 (N_11415,N_6474,N_7144);
or U11416 (N_11416,N_7158,N_6339);
or U11417 (N_11417,N_8452,N_6509);
or U11418 (N_11418,N_7855,N_8713);
nor U11419 (N_11419,N_8291,N_6184);
and U11420 (N_11420,N_7771,N_6427);
nand U11421 (N_11421,N_7610,N_7570);
or U11422 (N_11422,N_6717,N_8395);
xor U11423 (N_11423,N_8201,N_6939);
or U11424 (N_11424,N_7601,N_7927);
and U11425 (N_11425,N_7916,N_6912);
and U11426 (N_11426,N_8915,N_8082);
and U11427 (N_11427,N_7650,N_6593);
nor U11428 (N_11428,N_7613,N_8490);
and U11429 (N_11429,N_7471,N_8854);
or U11430 (N_11430,N_8105,N_8385);
nand U11431 (N_11431,N_6760,N_7133);
nor U11432 (N_11432,N_8105,N_8168);
or U11433 (N_11433,N_6111,N_7456);
or U11434 (N_11434,N_7527,N_7032);
or U11435 (N_11435,N_6706,N_8065);
xnor U11436 (N_11436,N_8262,N_6464);
or U11437 (N_11437,N_7650,N_6301);
or U11438 (N_11438,N_7195,N_8617);
nand U11439 (N_11439,N_7971,N_6764);
and U11440 (N_11440,N_8531,N_6960);
nor U11441 (N_11441,N_6475,N_8690);
nand U11442 (N_11442,N_8499,N_6529);
nand U11443 (N_11443,N_7794,N_6911);
xor U11444 (N_11444,N_8510,N_8814);
nor U11445 (N_11445,N_7499,N_8236);
or U11446 (N_11446,N_8054,N_8335);
and U11447 (N_11447,N_6901,N_7053);
or U11448 (N_11448,N_8240,N_6216);
nand U11449 (N_11449,N_7583,N_8598);
or U11450 (N_11450,N_8995,N_6187);
and U11451 (N_11451,N_6622,N_8801);
nor U11452 (N_11452,N_7322,N_8107);
xnor U11453 (N_11453,N_7599,N_7479);
nand U11454 (N_11454,N_8267,N_8291);
and U11455 (N_11455,N_7194,N_6843);
nand U11456 (N_11456,N_7200,N_6465);
xor U11457 (N_11457,N_7437,N_6209);
or U11458 (N_11458,N_6660,N_6831);
nand U11459 (N_11459,N_6312,N_6201);
nand U11460 (N_11460,N_7319,N_7093);
xnor U11461 (N_11461,N_8336,N_7213);
or U11462 (N_11462,N_6024,N_8768);
nand U11463 (N_11463,N_7106,N_8557);
xnor U11464 (N_11464,N_8180,N_7558);
xnor U11465 (N_11465,N_7763,N_8415);
nand U11466 (N_11466,N_6297,N_8935);
and U11467 (N_11467,N_7648,N_6397);
nor U11468 (N_11468,N_6118,N_6137);
nand U11469 (N_11469,N_7470,N_6910);
nand U11470 (N_11470,N_8124,N_7162);
nand U11471 (N_11471,N_6562,N_8471);
nand U11472 (N_11472,N_7583,N_6669);
nand U11473 (N_11473,N_6312,N_7633);
and U11474 (N_11474,N_7511,N_6985);
or U11475 (N_11475,N_6999,N_6048);
nor U11476 (N_11476,N_7513,N_8605);
or U11477 (N_11477,N_6930,N_7600);
or U11478 (N_11478,N_7813,N_6340);
xnor U11479 (N_11479,N_6466,N_7738);
and U11480 (N_11480,N_7203,N_8054);
nor U11481 (N_11481,N_7118,N_6526);
or U11482 (N_11482,N_7273,N_6291);
or U11483 (N_11483,N_8506,N_7685);
and U11484 (N_11484,N_7517,N_6332);
and U11485 (N_11485,N_6102,N_8302);
nor U11486 (N_11486,N_8997,N_7856);
xnor U11487 (N_11487,N_7627,N_8022);
xnor U11488 (N_11488,N_6957,N_6126);
nor U11489 (N_11489,N_7772,N_6202);
and U11490 (N_11490,N_8145,N_8355);
nand U11491 (N_11491,N_6431,N_6043);
nand U11492 (N_11492,N_7116,N_7410);
nor U11493 (N_11493,N_7290,N_6384);
and U11494 (N_11494,N_8684,N_6734);
nand U11495 (N_11495,N_6061,N_7168);
or U11496 (N_11496,N_6197,N_6884);
nor U11497 (N_11497,N_6383,N_6837);
xnor U11498 (N_11498,N_8341,N_8955);
xor U11499 (N_11499,N_7040,N_8776);
nand U11500 (N_11500,N_6417,N_8203);
and U11501 (N_11501,N_8244,N_6829);
nand U11502 (N_11502,N_6086,N_8804);
xor U11503 (N_11503,N_8299,N_8933);
nor U11504 (N_11504,N_6260,N_7405);
and U11505 (N_11505,N_6989,N_6717);
and U11506 (N_11506,N_6298,N_6659);
nor U11507 (N_11507,N_6616,N_8878);
xor U11508 (N_11508,N_8596,N_6174);
or U11509 (N_11509,N_6944,N_8177);
or U11510 (N_11510,N_7705,N_6274);
nand U11511 (N_11511,N_7730,N_6236);
and U11512 (N_11512,N_8380,N_8887);
nor U11513 (N_11513,N_8755,N_6536);
or U11514 (N_11514,N_8738,N_8485);
nand U11515 (N_11515,N_6401,N_8779);
xor U11516 (N_11516,N_7032,N_8775);
nor U11517 (N_11517,N_6959,N_6722);
or U11518 (N_11518,N_8960,N_7199);
and U11519 (N_11519,N_6513,N_7341);
xnor U11520 (N_11520,N_6016,N_8174);
or U11521 (N_11521,N_8054,N_7721);
and U11522 (N_11522,N_6588,N_6805);
or U11523 (N_11523,N_7101,N_6956);
nor U11524 (N_11524,N_6251,N_6632);
xor U11525 (N_11525,N_6474,N_6282);
nor U11526 (N_11526,N_6444,N_8602);
nor U11527 (N_11527,N_7834,N_7303);
nand U11528 (N_11528,N_6590,N_7208);
or U11529 (N_11529,N_8414,N_7730);
and U11530 (N_11530,N_8910,N_8111);
xnor U11531 (N_11531,N_6039,N_8698);
nor U11532 (N_11532,N_8103,N_7306);
or U11533 (N_11533,N_6320,N_7854);
and U11534 (N_11534,N_7482,N_6463);
nor U11535 (N_11535,N_8665,N_7651);
xnor U11536 (N_11536,N_7133,N_8874);
nand U11537 (N_11537,N_8354,N_7696);
nor U11538 (N_11538,N_8793,N_6572);
nor U11539 (N_11539,N_6280,N_8684);
and U11540 (N_11540,N_6785,N_6307);
nand U11541 (N_11541,N_8779,N_8986);
and U11542 (N_11542,N_7457,N_6106);
xnor U11543 (N_11543,N_8758,N_6824);
xor U11544 (N_11544,N_6587,N_6227);
and U11545 (N_11545,N_8525,N_8752);
nand U11546 (N_11546,N_8945,N_6838);
nand U11547 (N_11547,N_7319,N_7540);
nor U11548 (N_11548,N_6162,N_6561);
or U11549 (N_11549,N_7897,N_7113);
xor U11550 (N_11550,N_6932,N_6162);
nand U11551 (N_11551,N_6228,N_8877);
and U11552 (N_11552,N_6315,N_8963);
nor U11553 (N_11553,N_8432,N_6280);
xnor U11554 (N_11554,N_7475,N_7485);
nand U11555 (N_11555,N_7353,N_7221);
or U11556 (N_11556,N_7114,N_7633);
or U11557 (N_11557,N_6135,N_8818);
and U11558 (N_11558,N_8398,N_8896);
nand U11559 (N_11559,N_8055,N_6059);
and U11560 (N_11560,N_6545,N_7163);
nor U11561 (N_11561,N_7370,N_6530);
xor U11562 (N_11562,N_7696,N_6649);
xor U11563 (N_11563,N_7968,N_6538);
nand U11564 (N_11564,N_7650,N_8497);
xor U11565 (N_11565,N_7093,N_6987);
nor U11566 (N_11566,N_6786,N_8319);
nor U11567 (N_11567,N_6611,N_6365);
nand U11568 (N_11568,N_6028,N_8916);
xor U11569 (N_11569,N_6592,N_8169);
and U11570 (N_11570,N_6579,N_6225);
nand U11571 (N_11571,N_6577,N_7847);
nor U11572 (N_11572,N_6043,N_8281);
nand U11573 (N_11573,N_7166,N_6683);
xnor U11574 (N_11574,N_8240,N_8698);
xor U11575 (N_11575,N_7783,N_8651);
and U11576 (N_11576,N_8979,N_6612);
xnor U11577 (N_11577,N_8684,N_6744);
xnor U11578 (N_11578,N_6054,N_6076);
or U11579 (N_11579,N_7058,N_8551);
nand U11580 (N_11580,N_7032,N_8306);
nand U11581 (N_11581,N_7604,N_7934);
and U11582 (N_11582,N_8471,N_6669);
or U11583 (N_11583,N_7299,N_6083);
xor U11584 (N_11584,N_7138,N_6071);
or U11585 (N_11585,N_8150,N_8336);
nand U11586 (N_11586,N_6683,N_6129);
nor U11587 (N_11587,N_8687,N_8407);
nand U11588 (N_11588,N_8198,N_7884);
nor U11589 (N_11589,N_7890,N_8670);
or U11590 (N_11590,N_8629,N_6729);
xor U11591 (N_11591,N_6732,N_6494);
nand U11592 (N_11592,N_8862,N_6098);
nor U11593 (N_11593,N_8668,N_7218);
nor U11594 (N_11594,N_6852,N_7434);
or U11595 (N_11595,N_7234,N_7372);
nand U11596 (N_11596,N_7559,N_8783);
nor U11597 (N_11597,N_6169,N_7772);
xnor U11598 (N_11598,N_6359,N_6838);
xor U11599 (N_11599,N_6251,N_7810);
xor U11600 (N_11600,N_7614,N_8008);
nor U11601 (N_11601,N_8892,N_7889);
nor U11602 (N_11602,N_6187,N_6086);
or U11603 (N_11603,N_7716,N_8013);
nand U11604 (N_11604,N_8588,N_6541);
nand U11605 (N_11605,N_7993,N_6356);
or U11606 (N_11606,N_7562,N_8470);
nand U11607 (N_11607,N_7140,N_6772);
xnor U11608 (N_11608,N_7440,N_6942);
nand U11609 (N_11609,N_6629,N_6635);
nand U11610 (N_11610,N_7423,N_8429);
nor U11611 (N_11611,N_6384,N_6675);
and U11612 (N_11612,N_6012,N_8117);
nor U11613 (N_11613,N_6627,N_7684);
nor U11614 (N_11614,N_8052,N_6056);
or U11615 (N_11615,N_6451,N_8745);
nor U11616 (N_11616,N_6469,N_6197);
nand U11617 (N_11617,N_7211,N_7816);
and U11618 (N_11618,N_6050,N_6967);
or U11619 (N_11619,N_8956,N_6331);
nand U11620 (N_11620,N_7896,N_8793);
xnor U11621 (N_11621,N_6286,N_6277);
nor U11622 (N_11622,N_8327,N_8546);
nand U11623 (N_11623,N_6397,N_6180);
and U11624 (N_11624,N_6864,N_8717);
xor U11625 (N_11625,N_8433,N_8468);
nand U11626 (N_11626,N_6795,N_8189);
nor U11627 (N_11627,N_7243,N_6276);
or U11628 (N_11628,N_8432,N_7696);
or U11629 (N_11629,N_7651,N_8449);
nor U11630 (N_11630,N_8115,N_6236);
xnor U11631 (N_11631,N_6247,N_7330);
nor U11632 (N_11632,N_6147,N_8616);
nor U11633 (N_11633,N_6872,N_6512);
nand U11634 (N_11634,N_7603,N_8326);
nor U11635 (N_11635,N_8423,N_6420);
nor U11636 (N_11636,N_8938,N_8520);
xor U11637 (N_11637,N_6142,N_7899);
nand U11638 (N_11638,N_8190,N_7367);
xnor U11639 (N_11639,N_7364,N_8932);
xnor U11640 (N_11640,N_8700,N_7156);
nand U11641 (N_11641,N_8252,N_8650);
nor U11642 (N_11642,N_7601,N_6059);
xnor U11643 (N_11643,N_8759,N_7556);
xnor U11644 (N_11644,N_7998,N_8761);
or U11645 (N_11645,N_6204,N_6863);
and U11646 (N_11646,N_6671,N_6321);
and U11647 (N_11647,N_8848,N_6188);
and U11648 (N_11648,N_8718,N_7305);
or U11649 (N_11649,N_7176,N_6042);
nand U11650 (N_11650,N_8319,N_8047);
xnor U11651 (N_11651,N_6056,N_7259);
or U11652 (N_11652,N_8956,N_8535);
nor U11653 (N_11653,N_7047,N_7095);
nor U11654 (N_11654,N_6764,N_6338);
xor U11655 (N_11655,N_7503,N_6193);
or U11656 (N_11656,N_6765,N_6451);
or U11657 (N_11657,N_7223,N_8045);
nor U11658 (N_11658,N_8435,N_8832);
nor U11659 (N_11659,N_6410,N_8164);
nand U11660 (N_11660,N_8312,N_8206);
xor U11661 (N_11661,N_7868,N_7528);
and U11662 (N_11662,N_6540,N_8671);
nor U11663 (N_11663,N_7289,N_6379);
nor U11664 (N_11664,N_8317,N_6972);
nand U11665 (N_11665,N_7092,N_6356);
nor U11666 (N_11666,N_7889,N_8248);
and U11667 (N_11667,N_7906,N_7391);
or U11668 (N_11668,N_6272,N_7843);
nor U11669 (N_11669,N_6471,N_8068);
nand U11670 (N_11670,N_6772,N_6285);
or U11671 (N_11671,N_6578,N_7795);
xnor U11672 (N_11672,N_7478,N_6206);
or U11673 (N_11673,N_7740,N_6458);
or U11674 (N_11674,N_7903,N_7567);
nand U11675 (N_11675,N_7794,N_7593);
or U11676 (N_11676,N_7157,N_8250);
nor U11677 (N_11677,N_7604,N_6460);
nor U11678 (N_11678,N_8193,N_7412);
and U11679 (N_11679,N_8910,N_7354);
nand U11680 (N_11680,N_7836,N_6399);
nor U11681 (N_11681,N_6559,N_7312);
nor U11682 (N_11682,N_6212,N_6980);
xor U11683 (N_11683,N_8470,N_7380);
or U11684 (N_11684,N_8842,N_7040);
and U11685 (N_11685,N_6714,N_6698);
nor U11686 (N_11686,N_7021,N_6748);
and U11687 (N_11687,N_8970,N_7223);
or U11688 (N_11688,N_7667,N_6979);
xor U11689 (N_11689,N_6327,N_7973);
nor U11690 (N_11690,N_8176,N_7275);
xnor U11691 (N_11691,N_8182,N_6696);
xor U11692 (N_11692,N_7529,N_7632);
xor U11693 (N_11693,N_8760,N_8965);
or U11694 (N_11694,N_7825,N_7832);
or U11695 (N_11695,N_7531,N_6675);
or U11696 (N_11696,N_7160,N_8282);
nor U11697 (N_11697,N_6150,N_6823);
nor U11698 (N_11698,N_6035,N_7383);
nand U11699 (N_11699,N_8934,N_6848);
and U11700 (N_11700,N_7421,N_6957);
and U11701 (N_11701,N_7039,N_7669);
nor U11702 (N_11702,N_8625,N_8127);
or U11703 (N_11703,N_7682,N_8082);
xnor U11704 (N_11704,N_6245,N_7604);
or U11705 (N_11705,N_6170,N_7423);
and U11706 (N_11706,N_7413,N_6398);
or U11707 (N_11707,N_7135,N_8209);
xnor U11708 (N_11708,N_8839,N_7757);
xnor U11709 (N_11709,N_7022,N_6576);
nand U11710 (N_11710,N_8313,N_7461);
or U11711 (N_11711,N_8136,N_8119);
nor U11712 (N_11712,N_6783,N_6409);
and U11713 (N_11713,N_7378,N_8613);
xor U11714 (N_11714,N_7637,N_6277);
xor U11715 (N_11715,N_7408,N_6077);
or U11716 (N_11716,N_8372,N_6218);
nor U11717 (N_11717,N_8933,N_6814);
nand U11718 (N_11718,N_7693,N_7553);
and U11719 (N_11719,N_7685,N_6601);
nor U11720 (N_11720,N_7319,N_7099);
or U11721 (N_11721,N_7992,N_7450);
nand U11722 (N_11722,N_6273,N_8085);
and U11723 (N_11723,N_8261,N_8356);
xnor U11724 (N_11724,N_6762,N_6649);
nand U11725 (N_11725,N_6266,N_8233);
xor U11726 (N_11726,N_6285,N_7575);
and U11727 (N_11727,N_6106,N_6473);
or U11728 (N_11728,N_7916,N_7854);
xor U11729 (N_11729,N_7154,N_6012);
nand U11730 (N_11730,N_8172,N_6073);
and U11731 (N_11731,N_6086,N_8222);
nor U11732 (N_11732,N_7381,N_7539);
or U11733 (N_11733,N_7837,N_6809);
and U11734 (N_11734,N_6785,N_8869);
xor U11735 (N_11735,N_8205,N_6228);
xor U11736 (N_11736,N_6993,N_7497);
and U11737 (N_11737,N_7980,N_6489);
xnor U11738 (N_11738,N_8770,N_8080);
and U11739 (N_11739,N_8165,N_6982);
xor U11740 (N_11740,N_8399,N_7432);
xor U11741 (N_11741,N_8214,N_7601);
nor U11742 (N_11742,N_6375,N_8202);
and U11743 (N_11743,N_7775,N_7758);
and U11744 (N_11744,N_6201,N_7084);
or U11745 (N_11745,N_6581,N_8869);
nor U11746 (N_11746,N_8531,N_7094);
nor U11747 (N_11747,N_7721,N_8980);
and U11748 (N_11748,N_7087,N_6252);
and U11749 (N_11749,N_8023,N_7437);
or U11750 (N_11750,N_6745,N_8531);
xor U11751 (N_11751,N_6214,N_8330);
or U11752 (N_11752,N_6273,N_7325);
and U11753 (N_11753,N_6914,N_7073);
or U11754 (N_11754,N_6576,N_7504);
nor U11755 (N_11755,N_6929,N_8361);
or U11756 (N_11756,N_7953,N_7652);
xor U11757 (N_11757,N_6219,N_8096);
nand U11758 (N_11758,N_8690,N_7966);
and U11759 (N_11759,N_7793,N_7399);
nand U11760 (N_11760,N_7324,N_7606);
or U11761 (N_11761,N_7535,N_8470);
nand U11762 (N_11762,N_8897,N_8618);
nand U11763 (N_11763,N_8602,N_6436);
xor U11764 (N_11764,N_8948,N_8532);
nor U11765 (N_11765,N_7925,N_7569);
and U11766 (N_11766,N_6068,N_6278);
xnor U11767 (N_11767,N_7324,N_6458);
nand U11768 (N_11768,N_7264,N_7803);
and U11769 (N_11769,N_8041,N_6130);
nor U11770 (N_11770,N_8693,N_7547);
nor U11771 (N_11771,N_8402,N_8969);
nor U11772 (N_11772,N_8859,N_6171);
or U11773 (N_11773,N_8881,N_8098);
and U11774 (N_11774,N_6906,N_7242);
and U11775 (N_11775,N_7327,N_6095);
or U11776 (N_11776,N_8097,N_6400);
or U11777 (N_11777,N_7258,N_8537);
xor U11778 (N_11778,N_8529,N_7437);
nor U11779 (N_11779,N_8581,N_6429);
nand U11780 (N_11780,N_6279,N_7300);
xnor U11781 (N_11781,N_8534,N_8892);
or U11782 (N_11782,N_8460,N_8598);
nor U11783 (N_11783,N_6260,N_8283);
xor U11784 (N_11784,N_7178,N_6330);
nor U11785 (N_11785,N_6990,N_6848);
and U11786 (N_11786,N_8679,N_6680);
nor U11787 (N_11787,N_7747,N_6536);
nor U11788 (N_11788,N_6772,N_7438);
or U11789 (N_11789,N_7505,N_6826);
nor U11790 (N_11790,N_8333,N_8781);
nand U11791 (N_11791,N_7667,N_6966);
nor U11792 (N_11792,N_6361,N_8379);
and U11793 (N_11793,N_6856,N_8054);
and U11794 (N_11794,N_6323,N_7894);
or U11795 (N_11795,N_7415,N_8844);
nor U11796 (N_11796,N_8209,N_7810);
nand U11797 (N_11797,N_8248,N_8730);
nand U11798 (N_11798,N_6439,N_7756);
nor U11799 (N_11799,N_6850,N_6993);
and U11800 (N_11800,N_6383,N_6403);
nand U11801 (N_11801,N_7570,N_8418);
and U11802 (N_11802,N_8065,N_7543);
xor U11803 (N_11803,N_6061,N_8593);
or U11804 (N_11804,N_7496,N_7328);
xor U11805 (N_11805,N_6731,N_8156);
nor U11806 (N_11806,N_8883,N_6767);
or U11807 (N_11807,N_8365,N_7879);
or U11808 (N_11808,N_7205,N_7324);
xnor U11809 (N_11809,N_7465,N_8723);
and U11810 (N_11810,N_6823,N_7377);
or U11811 (N_11811,N_6278,N_8241);
and U11812 (N_11812,N_8347,N_8115);
and U11813 (N_11813,N_6629,N_7716);
xnor U11814 (N_11814,N_6979,N_8104);
or U11815 (N_11815,N_8868,N_8909);
and U11816 (N_11816,N_8647,N_6589);
nor U11817 (N_11817,N_8548,N_7112);
or U11818 (N_11818,N_8304,N_7941);
xnor U11819 (N_11819,N_8925,N_6976);
and U11820 (N_11820,N_7971,N_7767);
or U11821 (N_11821,N_6145,N_7093);
or U11822 (N_11822,N_8195,N_8124);
nand U11823 (N_11823,N_8666,N_8993);
or U11824 (N_11824,N_6969,N_8759);
xor U11825 (N_11825,N_7076,N_7817);
xnor U11826 (N_11826,N_8407,N_8343);
xor U11827 (N_11827,N_7566,N_7317);
and U11828 (N_11828,N_7446,N_6306);
nor U11829 (N_11829,N_7799,N_7285);
or U11830 (N_11830,N_7815,N_6131);
nor U11831 (N_11831,N_7831,N_6482);
xor U11832 (N_11832,N_8251,N_7388);
nor U11833 (N_11833,N_7851,N_7387);
and U11834 (N_11834,N_6460,N_7832);
and U11835 (N_11835,N_8387,N_8307);
or U11836 (N_11836,N_6224,N_6893);
nand U11837 (N_11837,N_8358,N_7398);
nand U11838 (N_11838,N_7260,N_7756);
xnor U11839 (N_11839,N_7845,N_8851);
or U11840 (N_11840,N_7700,N_6182);
xnor U11841 (N_11841,N_6802,N_8381);
nor U11842 (N_11842,N_6974,N_6249);
xnor U11843 (N_11843,N_6553,N_6253);
nor U11844 (N_11844,N_7636,N_8344);
xor U11845 (N_11845,N_7646,N_7434);
nor U11846 (N_11846,N_8092,N_7425);
xnor U11847 (N_11847,N_7447,N_6042);
or U11848 (N_11848,N_8702,N_8874);
xor U11849 (N_11849,N_6386,N_6214);
nor U11850 (N_11850,N_6852,N_6644);
and U11851 (N_11851,N_8820,N_7341);
xor U11852 (N_11852,N_8552,N_6837);
xnor U11853 (N_11853,N_8965,N_6782);
nor U11854 (N_11854,N_6142,N_7735);
xor U11855 (N_11855,N_8054,N_7350);
or U11856 (N_11856,N_6484,N_8872);
and U11857 (N_11857,N_7649,N_7982);
nor U11858 (N_11858,N_7591,N_8972);
and U11859 (N_11859,N_7436,N_6356);
nor U11860 (N_11860,N_7175,N_8877);
and U11861 (N_11861,N_7411,N_7145);
and U11862 (N_11862,N_8882,N_8552);
and U11863 (N_11863,N_7448,N_6715);
xnor U11864 (N_11864,N_6305,N_6015);
and U11865 (N_11865,N_6539,N_8864);
and U11866 (N_11866,N_6881,N_6782);
xnor U11867 (N_11867,N_8976,N_8383);
nand U11868 (N_11868,N_6866,N_8080);
and U11869 (N_11869,N_7221,N_6488);
nand U11870 (N_11870,N_8258,N_6369);
nor U11871 (N_11871,N_8455,N_6269);
xor U11872 (N_11872,N_7939,N_7166);
xnor U11873 (N_11873,N_8218,N_8978);
and U11874 (N_11874,N_7344,N_8507);
xor U11875 (N_11875,N_6390,N_7665);
nand U11876 (N_11876,N_7853,N_6336);
and U11877 (N_11877,N_6996,N_7915);
xnor U11878 (N_11878,N_6222,N_8373);
nor U11879 (N_11879,N_7559,N_7202);
nand U11880 (N_11880,N_8049,N_8733);
nand U11881 (N_11881,N_7465,N_6212);
and U11882 (N_11882,N_6521,N_8217);
or U11883 (N_11883,N_8300,N_7192);
or U11884 (N_11884,N_6953,N_7303);
or U11885 (N_11885,N_8172,N_8699);
and U11886 (N_11886,N_7160,N_8008);
or U11887 (N_11887,N_8463,N_8705);
xor U11888 (N_11888,N_8484,N_6768);
nor U11889 (N_11889,N_8421,N_6386);
or U11890 (N_11890,N_7689,N_6109);
xor U11891 (N_11891,N_8483,N_6488);
or U11892 (N_11892,N_7967,N_7158);
and U11893 (N_11893,N_7075,N_7445);
nor U11894 (N_11894,N_6079,N_6023);
and U11895 (N_11895,N_8234,N_8087);
nor U11896 (N_11896,N_7218,N_7442);
xor U11897 (N_11897,N_7238,N_8884);
nand U11898 (N_11898,N_6638,N_6031);
xnor U11899 (N_11899,N_8123,N_6872);
and U11900 (N_11900,N_8634,N_6708);
or U11901 (N_11901,N_6539,N_6148);
nand U11902 (N_11902,N_7486,N_7617);
and U11903 (N_11903,N_8732,N_8306);
xor U11904 (N_11904,N_7123,N_8960);
xnor U11905 (N_11905,N_7840,N_8393);
nand U11906 (N_11906,N_6158,N_7882);
or U11907 (N_11907,N_7664,N_6503);
and U11908 (N_11908,N_7524,N_8240);
nor U11909 (N_11909,N_6260,N_8453);
and U11910 (N_11910,N_7310,N_6590);
nand U11911 (N_11911,N_7994,N_6844);
or U11912 (N_11912,N_7608,N_7170);
xor U11913 (N_11913,N_8786,N_6693);
or U11914 (N_11914,N_7996,N_6510);
or U11915 (N_11915,N_7973,N_7043);
nand U11916 (N_11916,N_6901,N_8992);
and U11917 (N_11917,N_8580,N_8343);
nor U11918 (N_11918,N_6057,N_7097);
nor U11919 (N_11919,N_6627,N_8615);
and U11920 (N_11920,N_6841,N_7437);
xnor U11921 (N_11921,N_6456,N_6526);
nor U11922 (N_11922,N_6733,N_6806);
nand U11923 (N_11923,N_7832,N_8490);
nor U11924 (N_11924,N_7026,N_8846);
nand U11925 (N_11925,N_7747,N_7499);
xor U11926 (N_11926,N_6195,N_8278);
and U11927 (N_11927,N_7893,N_6465);
or U11928 (N_11928,N_6006,N_7349);
nand U11929 (N_11929,N_6784,N_7610);
nor U11930 (N_11930,N_7709,N_8941);
nor U11931 (N_11931,N_6247,N_7366);
nand U11932 (N_11932,N_8274,N_7324);
nand U11933 (N_11933,N_7323,N_8702);
or U11934 (N_11934,N_8352,N_7357);
or U11935 (N_11935,N_7118,N_7007);
and U11936 (N_11936,N_6315,N_7463);
nand U11937 (N_11937,N_8240,N_8336);
xor U11938 (N_11938,N_8632,N_7657);
nor U11939 (N_11939,N_7895,N_6871);
nand U11940 (N_11940,N_8695,N_8065);
nand U11941 (N_11941,N_7210,N_8951);
nor U11942 (N_11942,N_7853,N_7030);
or U11943 (N_11943,N_7836,N_7148);
and U11944 (N_11944,N_6507,N_7446);
and U11945 (N_11945,N_7205,N_7477);
xnor U11946 (N_11946,N_8796,N_8524);
or U11947 (N_11947,N_7512,N_8049);
nand U11948 (N_11948,N_6417,N_7040);
or U11949 (N_11949,N_7824,N_7045);
xnor U11950 (N_11950,N_8677,N_7817);
or U11951 (N_11951,N_8208,N_7135);
or U11952 (N_11952,N_8873,N_7875);
nand U11953 (N_11953,N_6750,N_6820);
and U11954 (N_11954,N_8675,N_6168);
or U11955 (N_11955,N_8042,N_7116);
or U11956 (N_11956,N_7028,N_7849);
or U11957 (N_11957,N_8358,N_6614);
or U11958 (N_11958,N_6222,N_8310);
or U11959 (N_11959,N_8925,N_7139);
nand U11960 (N_11960,N_7933,N_7052);
nand U11961 (N_11961,N_7616,N_6761);
or U11962 (N_11962,N_6570,N_7536);
or U11963 (N_11963,N_7270,N_7140);
xor U11964 (N_11964,N_8589,N_6117);
xnor U11965 (N_11965,N_7375,N_8928);
nor U11966 (N_11966,N_8567,N_6484);
nor U11967 (N_11967,N_7208,N_7842);
nand U11968 (N_11968,N_8176,N_7542);
nor U11969 (N_11969,N_6678,N_8797);
and U11970 (N_11970,N_6461,N_6611);
and U11971 (N_11971,N_6834,N_7246);
or U11972 (N_11972,N_8425,N_7102);
nor U11973 (N_11973,N_8247,N_8463);
xor U11974 (N_11974,N_7279,N_8929);
nor U11975 (N_11975,N_6673,N_6684);
or U11976 (N_11976,N_7058,N_6466);
and U11977 (N_11977,N_6017,N_8641);
xor U11978 (N_11978,N_7802,N_6269);
and U11979 (N_11979,N_6459,N_6299);
or U11980 (N_11980,N_8010,N_8367);
and U11981 (N_11981,N_6417,N_8436);
nor U11982 (N_11982,N_7093,N_8894);
nand U11983 (N_11983,N_8382,N_7353);
nor U11984 (N_11984,N_7882,N_7452);
and U11985 (N_11985,N_6283,N_8956);
and U11986 (N_11986,N_6938,N_7391);
or U11987 (N_11987,N_8830,N_6463);
and U11988 (N_11988,N_6805,N_6194);
or U11989 (N_11989,N_8086,N_7252);
nand U11990 (N_11990,N_7140,N_6005);
xnor U11991 (N_11991,N_6193,N_7214);
and U11992 (N_11992,N_7212,N_7226);
nand U11993 (N_11993,N_6269,N_6146);
xor U11994 (N_11994,N_8408,N_8770);
nor U11995 (N_11995,N_8513,N_8493);
nor U11996 (N_11996,N_6613,N_7584);
xnor U11997 (N_11997,N_6087,N_7886);
nand U11998 (N_11998,N_8430,N_7922);
and U11999 (N_11999,N_8906,N_6828);
nor U12000 (N_12000,N_10805,N_10158);
xor U12001 (N_12001,N_9198,N_10584);
xor U12002 (N_12002,N_10346,N_9313);
or U12003 (N_12003,N_10445,N_11249);
or U12004 (N_12004,N_11035,N_11996);
and U12005 (N_12005,N_10570,N_10798);
xnor U12006 (N_12006,N_11207,N_11937);
and U12007 (N_12007,N_9137,N_10088);
and U12008 (N_12008,N_11679,N_10603);
and U12009 (N_12009,N_11517,N_10030);
nand U12010 (N_12010,N_11390,N_10174);
nor U12011 (N_12011,N_9207,N_11787);
nor U12012 (N_12012,N_9893,N_9534);
or U12013 (N_12013,N_9699,N_10077);
and U12014 (N_12014,N_9077,N_10604);
and U12015 (N_12015,N_9242,N_11220);
xnor U12016 (N_12016,N_10500,N_10385);
or U12017 (N_12017,N_10457,N_11840);
xor U12018 (N_12018,N_10530,N_10964);
xor U12019 (N_12019,N_10770,N_9188);
or U12020 (N_12020,N_10315,N_9233);
xnor U12021 (N_12021,N_11545,N_10237);
xnor U12022 (N_12022,N_9468,N_11537);
xnor U12023 (N_12023,N_9049,N_9870);
xnor U12024 (N_12024,N_9656,N_11610);
or U12025 (N_12025,N_10840,N_11083);
nand U12026 (N_12026,N_10723,N_11757);
xor U12027 (N_12027,N_10637,N_9814);
and U12028 (N_12028,N_9598,N_10134);
and U12029 (N_12029,N_9709,N_9469);
or U12030 (N_12030,N_10187,N_10109);
xnor U12031 (N_12031,N_9585,N_10156);
xnor U12032 (N_12032,N_11123,N_11255);
xnor U12033 (N_12033,N_11033,N_11809);
xor U12034 (N_12034,N_10463,N_11741);
nor U12035 (N_12035,N_11010,N_10976);
and U12036 (N_12036,N_11524,N_9296);
or U12037 (N_12037,N_9248,N_11192);
nand U12038 (N_12038,N_11142,N_9748);
or U12039 (N_12039,N_10998,N_10915);
or U12040 (N_12040,N_10355,N_11089);
xor U12041 (N_12041,N_9453,N_11362);
and U12042 (N_12042,N_11122,N_10135);
and U12043 (N_12043,N_10873,N_10348);
or U12044 (N_12044,N_11539,N_11723);
xor U12045 (N_12045,N_9231,N_9519);
nor U12046 (N_12046,N_10794,N_9247);
and U12047 (N_12047,N_9079,N_9877);
or U12048 (N_12048,N_11344,N_11898);
nor U12049 (N_12049,N_9727,N_10185);
nand U12050 (N_12050,N_11931,N_10248);
nor U12051 (N_12051,N_11989,N_11146);
or U12052 (N_12052,N_10425,N_10953);
and U12053 (N_12053,N_11941,N_10903);
xnor U12054 (N_12054,N_9511,N_11737);
nand U12055 (N_12055,N_10528,N_11124);
xor U12056 (N_12056,N_11072,N_9367);
nand U12057 (N_12057,N_9048,N_9029);
nor U12058 (N_12058,N_9266,N_11775);
and U12059 (N_12059,N_11167,N_10594);
xor U12060 (N_12060,N_10215,N_10577);
nor U12061 (N_12061,N_11606,N_11644);
xor U12062 (N_12062,N_11502,N_9543);
nor U12063 (N_12063,N_11882,N_10945);
and U12064 (N_12064,N_9662,N_9928);
nor U12065 (N_12065,N_10299,N_11237);
xor U12066 (N_12066,N_9508,N_11654);
nand U12067 (N_12067,N_10947,N_11385);
nand U12068 (N_12068,N_9769,N_11994);
nand U12069 (N_12069,N_9629,N_11183);
xnor U12070 (N_12070,N_11997,N_11678);
nor U12071 (N_12071,N_10833,N_10443);
nand U12072 (N_12072,N_9552,N_11351);
or U12073 (N_12073,N_11149,N_9818);
nor U12074 (N_12074,N_10183,N_9963);
nor U12075 (N_12075,N_10890,N_10830);
or U12076 (N_12076,N_9887,N_9310);
xnor U12077 (N_12077,N_11155,N_9240);
nor U12078 (N_12078,N_9906,N_9745);
xnor U12079 (N_12079,N_11844,N_10095);
nor U12080 (N_12080,N_9985,N_9530);
or U12081 (N_12081,N_9341,N_10051);
nor U12082 (N_12082,N_11747,N_9251);
nor U12083 (N_12083,N_9895,N_9679);
xor U12084 (N_12084,N_9702,N_11190);
and U12085 (N_12085,N_9631,N_10949);
or U12086 (N_12086,N_9352,N_9064);
xor U12087 (N_12087,N_11012,N_10785);
and U12088 (N_12088,N_11962,N_11990);
nand U12089 (N_12089,N_9236,N_11592);
nand U12090 (N_12090,N_9326,N_9124);
nor U12091 (N_12091,N_10234,N_11193);
nor U12092 (N_12092,N_9066,N_10005);
or U12093 (N_12093,N_11267,N_10857);
nand U12094 (N_12094,N_10126,N_9862);
nor U12095 (N_12095,N_9471,N_11055);
xnor U12096 (N_12096,N_11661,N_11949);
nand U12097 (N_12097,N_11622,N_10452);
and U12098 (N_12098,N_11693,N_11415);
xor U12099 (N_12099,N_11566,N_9861);
nor U12100 (N_12100,N_9210,N_10628);
nor U12101 (N_12101,N_10569,N_9217);
and U12102 (N_12102,N_10467,N_9558);
xnor U12103 (N_12103,N_9704,N_10605);
nor U12104 (N_12104,N_10148,N_11743);
or U12105 (N_12105,N_11384,N_10480);
nand U12106 (N_12106,N_10968,N_11579);
nand U12107 (N_12107,N_10193,N_9355);
xnor U12108 (N_12108,N_11536,N_9403);
and U12109 (N_12109,N_9966,N_9324);
and U12110 (N_12110,N_11369,N_9271);
nand U12111 (N_12111,N_11272,N_9160);
and U12112 (N_12112,N_11871,N_10329);
nor U12113 (N_12113,N_11530,N_10450);
nor U12114 (N_12114,N_10195,N_11806);
and U12115 (N_12115,N_11712,N_10004);
nand U12116 (N_12116,N_11869,N_9421);
or U12117 (N_12117,N_9990,N_9641);
xor U12118 (N_12118,N_9993,N_9987);
or U12119 (N_12119,N_10626,N_10598);
nand U12120 (N_12120,N_9696,N_11458);
xnor U12121 (N_12121,N_9839,N_11292);
xnor U12122 (N_12122,N_11805,N_11600);
nand U12123 (N_12123,N_11366,N_10880);
xnor U12124 (N_12124,N_10506,N_11211);
nor U12125 (N_12125,N_11224,N_11578);
or U12126 (N_12126,N_11746,N_11084);
nand U12127 (N_12127,N_9388,N_10521);
and U12128 (N_12128,N_10102,N_9920);
nand U12129 (N_12129,N_10847,N_9434);
nand U12130 (N_12130,N_10176,N_10260);
and U12131 (N_12131,N_10474,N_11497);
or U12132 (N_12132,N_9106,N_10013);
xor U12133 (N_12133,N_9135,N_11336);
and U12134 (N_12134,N_9357,N_11554);
and U12135 (N_12135,N_10323,N_11480);
nand U12136 (N_12136,N_10571,N_9295);
and U12137 (N_12137,N_9884,N_11498);
and U12138 (N_12138,N_11375,N_11819);
and U12139 (N_12139,N_11413,N_10032);
nor U12140 (N_12140,N_10600,N_10842);
nand U12141 (N_12141,N_10057,N_9622);
and U12142 (N_12142,N_9400,N_11347);
nand U12143 (N_12143,N_9022,N_11280);
nor U12144 (N_12144,N_9601,N_9956);
xor U12145 (N_12145,N_9875,N_9196);
nand U12146 (N_12146,N_9512,N_10455);
nor U12147 (N_12147,N_10067,N_9849);
and U12148 (N_12148,N_10305,N_10575);
and U12149 (N_12149,N_10122,N_11241);
and U12150 (N_12150,N_10550,N_10314);
and U12151 (N_12151,N_9268,N_9105);
or U12152 (N_12152,N_10327,N_10713);
and U12153 (N_12153,N_10536,N_9476);
nor U12154 (N_12154,N_9611,N_11125);
xnor U12155 (N_12155,N_9460,N_11427);
and U12156 (N_12156,N_11619,N_9683);
nand U12157 (N_12157,N_10415,N_11097);
nor U12158 (N_12158,N_9724,N_10357);
or U12159 (N_12159,N_11234,N_10317);
xnor U12160 (N_12160,N_10461,N_11635);
xnor U12161 (N_12161,N_11748,N_10621);
and U12162 (N_12162,N_10410,N_9024);
nand U12163 (N_12163,N_9654,N_10416);
nor U12164 (N_12164,N_11236,N_10812);
nand U12165 (N_12165,N_11812,N_9908);
and U12166 (N_12166,N_11031,N_11409);
nand U12167 (N_12167,N_9626,N_11297);
nand U12168 (N_12168,N_10336,N_9871);
nand U12169 (N_12169,N_11238,N_11643);
xnor U12170 (N_12170,N_11034,N_11667);
xor U12171 (N_12171,N_11750,N_9499);
and U12172 (N_12172,N_10276,N_9058);
or U12173 (N_12173,N_9931,N_10912);
and U12174 (N_12174,N_11309,N_9382);
nor U12175 (N_12175,N_9362,N_11404);
nor U12176 (N_12176,N_10779,N_11675);
nand U12177 (N_12177,N_11228,N_10140);
or U12178 (N_12178,N_10369,N_11328);
nor U12179 (N_12179,N_9316,N_11656);
nor U12180 (N_12180,N_9873,N_11910);
or U12181 (N_12181,N_10251,N_9789);
nand U12182 (N_12182,N_10732,N_10063);
and U12183 (N_12183,N_10627,N_9441);
nand U12184 (N_12184,N_9114,N_10647);
nand U12185 (N_12185,N_11153,N_9506);
xnor U12186 (N_12186,N_10339,N_11572);
and U12187 (N_12187,N_11810,N_11259);
nor U12188 (N_12188,N_9510,N_11186);
nor U12189 (N_12189,N_11711,N_9312);
and U12190 (N_12190,N_10921,N_10618);
and U12191 (N_12191,N_9718,N_10432);
xor U12192 (N_12192,N_11360,N_10611);
and U12193 (N_12193,N_11551,N_9147);
or U12194 (N_12194,N_10046,N_11864);
nand U12195 (N_12195,N_10108,N_10780);
or U12196 (N_12196,N_11525,N_10422);
nor U12197 (N_12197,N_9821,N_10472);
xnor U12198 (N_12198,N_10381,N_10629);
and U12199 (N_12199,N_9098,N_10619);
nor U12200 (N_12200,N_9811,N_9951);
or U12201 (N_12201,N_11363,N_9334);
and U12202 (N_12202,N_11916,N_10007);
nor U12203 (N_12203,N_9776,N_11611);
nand U12204 (N_12204,N_11768,N_9785);
nand U12205 (N_12205,N_9384,N_9161);
xor U12206 (N_12206,N_10935,N_11065);
nand U12207 (N_12207,N_10166,N_10045);
or U12208 (N_12208,N_11042,N_10331);
nor U12209 (N_12209,N_9596,N_11802);
nor U12210 (N_12210,N_11002,N_10849);
nor U12211 (N_12211,N_11728,N_10518);
nand U12212 (N_12212,N_11274,N_10661);
xor U12213 (N_12213,N_11912,N_11529);
and U12214 (N_12214,N_10539,N_9712);
xor U12215 (N_12215,N_11117,N_9673);
or U12216 (N_12216,N_9097,N_10739);
nor U12217 (N_12217,N_11063,N_11121);
xnor U12218 (N_12218,N_11273,N_9151);
xnor U12219 (N_12219,N_10612,N_9376);
xnor U12220 (N_12220,N_10981,N_10652);
and U12221 (N_12221,N_9689,N_9803);
nor U12222 (N_12222,N_9164,N_10275);
nor U12223 (N_12223,N_10241,N_10649);
xor U12224 (N_12224,N_9809,N_9968);
xnor U12225 (N_12225,N_9529,N_10560);
nor U12226 (N_12226,N_10219,N_9491);
nor U12227 (N_12227,N_9387,N_11247);
or U12228 (N_12228,N_11185,N_10145);
or U12229 (N_12229,N_11815,N_9256);
xnor U12230 (N_12230,N_10803,N_10267);
xnor U12231 (N_12231,N_10820,N_10200);
xor U12232 (N_12232,N_10939,N_11485);
or U12233 (N_12233,N_9459,N_9182);
and U12234 (N_12234,N_10100,N_9381);
xnor U12235 (N_12235,N_10653,N_9193);
and U12236 (N_12236,N_10103,N_10292);
nor U12237 (N_12237,N_10910,N_11509);
xor U12238 (N_12238,N_11513,N_11858);
xnor U12239 (N_12239,N_9886,N_9758);
and U12240 (N_12240,N_9498,N_10716);
xor U12241 (N_12241,N_11209,N_11000);
nor U12242 (N_12242,N_11357,N_11172);
nand U12243 (N_12243,N_9719,N_9041);
xor U12244 (N_12244,N_10634,N_9916);
and U12245 (N_12245,N_10035,N_11648);
xor U12246 (N_12246,N_9068,N_11219);
or U12247 (N_12247,N_10679,N_9995);
xor U12248 (N_12248,N_9345,N_11928);
xnor U12249 (N_12249,N_9455,N_9044);
nand U12250 (N_12250,N_10875,N_10549);
and U12251 (N_12251,N_10966,N_10610);
or U12252 (N_12252,N_11900,N_11573);
nand U12253 (N_12253,N_10105,N_10919);
nand U12254 (N_12254,N_9806,N_9778);
xnor U12255 (N_12255,N_9915,N_9447);
and U12256 (N_12256,N_9343,N_10497);
and U12257 (N_12257,N_10459,N_11521);
or U12258 (N_12258,N_9674,N_11461);
nand U12259 (N_12259,N_9396,N_9675);
nor U12260 (N_12260,N_10245,N_9548);
and U12261 (N_12261,N_11804,N_11132);
and U12262 (N_12262,N_11977,N_9320);
nor U12263 (N_12263,N_10133,N_9292);
xnor U12264 (N_12264,N_10831,N_11531);
or U12265 (N_12265,N_10316,N_11637);
or U12266 (N_12266,N_10520,N_10017);
and U12267 (N_12267,N_10635,N_9408);
and U12268 (N_12268,N_11792,N_10021);
xor U12269 (N_12269,N_10169,N_11368);
or U12270 (N_12270,N_11535,N_11841);
xnor U12271 (N_12271,N_11173,N_10059);
nor U12272 (N_12272,N_11716,N_9687);
xnor U12273 (N_12273,N_11543,N_9813);
nand U12274 (N_12274,N_9201,N_10392);
nand U12275 (N_12275,N_10042,N_10913);
nor U12276 (N_12276,N_11188,N_11473);
nor U12277 (N_12277,N_11602,N_11086);
nand U12278 (N_12278,N_9043,N_11668);
and U12279 (N_12279,N_11423,N_9574);
nand U12280 (N_12280,N_9903,N_10147);
nand U12281 (N_12281,N_9448,N_9964);
nor U12282 (N_12282,N_11260,N_10162);
xor U12283 (N_12283,N_10202,N_11329);
nand U12284 (N_12284,N_9439,N_11103);
and U12285 (N_12285,N_9697,N_9998);
nor U12286 (N_12286,N_9853,N_9083);
or U12287 (N_12287,N_11090,N_10424);
nand U12288 (N_12288,N_10591,N_9040);
nor U12289 (N_12289,N_10428,N_10413);
and U12290 (N_12290,N_10850,N_11338);
xnor U12291 (N_12291,N_10426,N_11909);
nor U12292 (N_12292,N_9805,N_9136);
or U12293 (N_12293,N_10361,N_9593);
nor U12294 (N_12294,N_10124,N_10885);
nand U12295 (N_12295,N_9801,N_9435);
nor U12296 (N_12296,N_11432,N_10483);
nor U12297 (N_12297,N_11682,N_9793);
xnor U12298 (N_12298,N_10640,N_9836);
xnor U12299 (N_12299,N_11947,N_9649);
xor U12300 (N_12300,N_11331,N_9405);
nor U12301 (N_12301,N_9138,N_10561);
nand U12302 (N_12302,N_10883,N_10396);
nor U12303 (N_12303,N_9905,N_11282);
nor U12304 (N_12304,N_11951,N_9166);
nand U12305 (N_12305,N_9738,N_9544);
nand U12306 (N_12306,N_10685,N_9226);
nor U12307 (N_12307,N_9630,N_9402);
or U12308 (N_12308,N_9346,N_11963);
nor U12309 (N_12309,N_11288,N_11923);
and U12310 (N_12310,N_9186,N_9669);
nand U12311 (N_12311,N_9464,N_11814);
or U12312 (N_12312,N_9329,N_9094);
nor U12313 (N_12313,N_11612,N_10283);
or U12314 (N_12314,N_10554,N_9483);
xnor U12315 (N_12315,N_9713,N_9907);
and U12316 (N_12316,N_10658,N_10181);
xnor U12317 (N_12317,N_11345,N_10250);
nand U12318 (N_12318,N_11742,N_11891);
nor U12319 (N_12319,N_9777,N_9122);
and U12320 (N_12320,N_10670,N_9981);
xor U12321 (N_12321,N_10468,N_11367);
nand U12322 (N_12322,N_10651,N_11283);
nand U12323 (N_12323,N_9281,N_11713);
xor U12324 (N_12324,N_10983,N_10889);
nor U12325 (N_12325,N_10789,N_9866);
nor U12326 (N_12326,N_11129,N_9314);
xnor U12327 (N_12327,N_9034,N_11040);
or U12328 (N_12328,N_9411,N_11957);
or U12329 (N_12329,N_11647,N_11137);
or U12330 (N_12330,N_9187,N_10226);
and U12331 (N_12331,N_10839,N_11334);
xnor U12332 (N_12332,N_9695,N_9501);
nand U12333 (N_12333,N_9762,N_10697);
or U12334 (N_12334,N_9072,N_9723);
nand U12335 (N_12335,N_9315,N_11587);
xor U12336 (N_12336,N_9131,N_11616);
nand U12337 (N_12337,N_9734,N_11901);
nand U12338 (N_12338,N_10249,N_9797);
or U12339 (N_12339,N_11917,N_10695);
nand U12340 (N_12340,N_9834,N_10863);
xnor U12341 (N_12341,N_10282,N_11223);
nor U12342 (N_12342,N_11455,N_11009);
xnor U12343 (N_12343,N_10993,N_10279);
or U12344 (N_12344,N_11570,N_10496);
nand U12345 (N_12345,N_9235,N_9211);
nand U12346 (N_12346,N_9133,N_11683);
nand U12347 (N_12347,N_11196,N_9204);
nor U12348 (N_12348,N_9017,N_10878);
or U12349 (N_12349,N_10982,N_10344);
nand U12350 (N_12350,N_10137,N_9795);
and U12351 (N_12351,N_10777,N_11617);
and U12352 (N_12352,N_11976,N_10493);
or U12353 (N_12353,N_9358,N_10099);
nand U12354 (N_12354,N_11721,N_11333);
or U12355 (N_12355,N_11230,N_11403);
or U12356 (N_12356,N_10535,N_11310);
xor U12357 (N_12357,N_9747,N_9191);
nand U12358 (N_12358,N_9978,N_9130);
and U12359 (N_12359,N_11460,N_9577);
nand U12360 (N_12360,N_10892,N_9994);
nor U12361 (N_12361,N_10907,N_11674);
nor U12362 (N_12362,N_11968,N_9688);
nor U12363 (N_12363,N_9898,N_10213);
xnor U12364 (N_12364,N_9567,N_9791);
or U12365 (N_12365,N_11965,N_11440);
xor U12366 (N_12366,N_11704,N_10920);
xor U12367 (N_12367,N_9216,N_10866);
nor U12368 (N_12368,N_10720,N_10934);
xor U12369 (N_12369,N_9370,N_10268);
or U12370 (N_12370,N_11684,N_11689);
or U12371 (N_12371,N_9527,N_11753);
nor U12372 (N_12372,N_10583,N_10741);
nor U12373 (N_12373,N_10714,N_10039);
or U12374 (N_12374,N_11411,N_11522);
and U12375 (N_12375,N_11439,N_11181);
and U12376 (N_12376,N_9609,N_9684);
nand U12377 (N_12377,N_10265,N_10227);
nor U12378 (N_12378,N_9472,N_11029);
nor U12379 (N_12379,N_9178,N_10548);
xor U12380 (N_12380,N_9588,N_11975);
or U12381 (N_12381,N_9430,N_11846);
and U12382 (N_12382,N_9897,N_10079);
or U12383 (N_12383,N_9982,N_11350);
and U12384 (N_12384,N_9282,N_9804);
xor U12385 (N_12385,N_9890,N_9466);
nand U12386 (N_12386,N_11527,N_9115);
nand U12387 (N_12387,N_10688,N_9280);
and U12388 (N_12388,N_11377,N_10269);
nand U12389 (N_12389,N_11549,N_11852);
and U12390 (N_12390,N_10198,N_11599);
or U12391 (N_12391,N_9715,N_9375);
nor U12392 (N_12392,N_10358,N_10264);
xnor U12393 (N_12393,N_11897,N_10318);
nand U12394 (N_12394,N_10752,N_10871);
nor U12395 (N_12395,N_10936,N_10904);
and U12396 (N_12396,N_11469,N_11519);
and U12397 (N_12397,N_11795,N_11094);
nand U12398 (N_12398,N_10545,N_9613);
nand U12399 (N_12399,N_11257,N_11091);
xor U12400 (N_12400,N_11569,N_11099);
and U12401 (N_12401,N_9194,N_11346);
xnor U12402 (N_12402,N_11774,N_11457);
nor U12403 (N_12403,N_11293,N_11623);
nand U12404 (N_12404,N_11349,N_11722);
xnor U12405 (N_12405,N_9359,N_11066);
nand U12406 (N_12406,N_11225,N_10877);
nand U12407 (N_12407,N_11553,N_10748);
nand U12408 (N_12408,N_10655,N_11200);
nand U12409 (N_12409,N_9788,N_11163);
and U12410 (N_12410,N_10371,N_10350);
xor U12411 (N_12411,N_11176,N_11179);
xnor U12412 (N_12412,N_10131,N_11630);
or U12413 (N_12413,N_11791,N_9433);
nor U12414 (N_12414,N_11051,N_9220);
nor U12415 (N_12415,N_10220,N_11087);
or U12416 (N_12416,N_11286,N_11402);
nand U12417 (N_12417,N_11581,N_10683);
and U12418 (N_12418,N_10524,N_9970);
nand U12419 (N_12419,N_11836,N_9290);
and U12420 (N_12420,N_10448,N_9063);
nor U12421 (N_12421,N_9011,N_10471);
or U12422 (N_12422,N_11902,N_11811);
and U12423 (N_12423,N_10252,N_9227);
nor U12424 (N_12424,N_11317,N_9002);
nor U12425 (N_12425,N_10663,N_10146);
and U12426 (N_12426,N_9270,N_10356);
and U12427 (N_12427,N_10261,N_9183);
nand U12428 (N_12428,N_11184,N_11300);
or U12429 (N_12429,N_9423,N_11490);
or U12430 (N_12430,N_11491,N_11863);
or U12431 (N_12431,N_11904,N_9333);
nor U12432 (N_12432,N_9680,N_10730);
nand U12433 (N_12433,N_11203,N_9865);
xnor U12434 (N_12434,N_11391,N_11355);
nor U12435 (N_12435,N_9417,N_9550);
or U12436 (N_12436,N_11641,N_11755);
or U12437 (N_12437,N_11006,N_11662);
nand U12438 (N_12438,N_10091,N_10078);
nor U12439 (N_12439,N_10565,N_10048);
nand U12440 (N_12440,N_10313,N_9933);
nor U12441 (N_12441,N_10853,N_11294);
xor U12442 (N_12442,N_11178,N_9031);
or U12443 (N_12443,N_9286,N_9635);
xnor U12444 (N_12444,N_10387,N_10433);
xnor U12445 (N_12445,N_11613,N_10121);
nor U12446 (N_12446,N_11061,N_10094);
xor U12447 (N_12447,N_9379,N_10544);
or U12448 (N_12448,N_9992,N_10946);
nand U12449 (N_12449,N_9323,N_11974);
and U12450 (N_12450,N_11538,N_11725);
xnor U12451 (N_12451,N_9036,N_11835);
nor U12452 (N_12452,N_10581,N_11004);
and U12453 (N_12453,N_11435,N_10072);
or U12454 (N_12454,N_9073,N_10563);
nand U12455 (N_12455,N_11177,N_9639);
and U12456 (N_12456,N_10893,N_11405);
xor U12457 (N_12457,N_9515,N_10613);
nand U12458 (N_12458,N_9910,N_10796);
xor U12459 (N_12459,N_9482,N_9497);
nor U12460 (N_12460,N_11943,N_11915);
nor U12461 (N_12461,N_10572,N_11905);
and U12462 (N_12462,N_10222,N_10816);
or U12463 (N_12463,N_9856,N_11053);
or U12464 (N_12464,N_11306,N_10191);
or U12465 (N_12465,N_9504,N_10645);
or U12466 (N_12466,N_10111,N_11598);
nor U12467 (N_12467,N_10793,N_11341);
and U12468 (N_12468,N_11546,N_11966);
xor U12469 (N_12469,N_9395,N_10308);
and U12470 (N_12470,N_9152,N_10991);
xor U12471 (N_12471,N_11204,N_9035);
or U12472 (N_12472,N_10391,N_11107);
xor U12473 (N_12473,N_9962,N_11467);
xnor U12474 (N_12474,N_10351,N_9787);
and U12475 (N_12475,N_11821,N_9168);
nor U12476 (N_12476,N_10182,N_10044);
nor U12477 (N_12477,N_9901,N_10025);
nor U12478 (N_12478,N_11295,N_9786);
and U12479 (N_12479,N_11304,N_10884);
and U12480 (N_12480,N_11954,N_10441);
xor U12481 (N_12481,N_10876,N_10733);
nor U12482 (N_12482,N_11567,N_10322);
and U12483 (N_12483,N_9580,N_9001);
and U12484 (N_12484,N_9822,N_9607);
nor U12485 (N_12485,N_10574,N_11050);
nand U12486 (N_12486,N_10475,N_10582);
and U12487 (N_12487,N_9616,N_9067);
xor U12488 (N_12488,N_11454,N_9944);
or U12489 (N_12489,N_10874,N_11466);
or U12490 (N_12490,N_9302,N_10034);
and U12491 (N_12491,N_10916,N_10207);
nor U12492 (N_12492,N_10050,N_9941);
and U12493 (N_12493,N_9935,N_9949);
and U12494 (N_12494,N_11762,N_11770);
xnor U12495 (N_12495,N_10901,N_9700);
nand U12496 (N_12496,N_11143,N_11270);
nor U12497 (N_12497,N_10484,N_11421);
or U12498 (N_12498,N_10469,N_10098);
nor U12499 (N_12499,N_9012,N_9560);
and U12500 (N_12500,N_11585,N_11922);
nand U12501 (N_12501,N_11269,N_11380);
and U12502 (N_12502,N_9756,N_10588);
nor U12503 (N_12503,N_11197,N_11240);
or U12504 (N_12504,N_10974,N_10186);
xnor U12505 (N_12505,N_9249,N_9045);
nor U12506 (N_12506,N_9707,N_11324);
xnor U12507 (N_12507,N_9535,N_9042);
xnor U12508 (N_12508,N_9652,N_9061);
or U12509 (N_12509,N_9647,N_9409);
nand U12510 (N_12510,N_10066,N_10810);
and U12511 (N_12511,N_9934,N_9470);
or U12512 (N_12512,N_9663,N_11649);
xnor U12513 (N_12513,N_11032,N_11729);
nand U12514 (N_12514,N_11154,N_11511);
nand U12515 (N_12515,N_11879,N_11991);
or U12516 (N_12516,N_10214,N_9410);
nor U12517 (N_12517,N_10390,N_9595);
or U12518 (N_12518,N_11348,N_11972);
nor U12519 (N_12519,N_9306,N_11505);
xnor U12520 (N_12520,N_11321,N_11077);
nor U12521 (N_12521,N_9109,N_9911);
or U12522 (N_12522,N_11894,N_9516);
or U12523 (N_12523,N_10644,N_10881);
xor U12524 (N_12524,N_9751,N_9028);
xor U12525 (N_12525,N_10896,N_10337);
nand U12526 (N_12526,N_9380,N_11314);
or U12527 (N_12527,N_9112,N_10141);
nor U12528 (N_12528,N_10080,N_11052);
xor U12529 (N_12529,N_9243,N_11636);
nand U12530 (N_12530,N_11515,N_10144);
or U12531 (N_12531,N_10675,N_10819);
or U12532 (N_12532,N_10206,N_10236);
and U12533 (N_12533,N_10625,N_9859);
nand U12534 (N_12534,N_10427,N_11964);
nand U12535 (N_12535,N_11779,N_9693);
nand U12536 (N_12536,N_10404,N_11938);
nand U12537 (N_12537,N_9730,N_10931);
xnor U12538 (N_12538,N_9522,N_11206);
xnor U12539 (N_12539,N_9015,N_9819);
xnor U12540 (N_12540,N_10401,N_11896);
and U12541 (N_12541,N_9092,N_11591);
xnor U12542 (N_12542,N_9729,N_11239);
and U12543 (N_12543,N_9880,N_10960);
nand U12544 (N_12544,N_10096,N_10012);
xor U12545 (N_12545,N_10143,N_10076);
nor U12546 (N_12546,N_9838,N_9495);
or U12547 (N_12547,N_10822,N_10786);
and U12548 (N_12548,N_11832,N_10989);
nand U12549 (N_12549,N_10373,N_10037);
nor U12550 (N_12550,N_10825,N_9304);
nand U12551 (N_12551,N_11870,N_10386);
and U12552 (N_12552,N_11232,N_10473);
and U12553 (N_12553,N_11803,N_10809);
xor U12554 (N_12554,N_9568,N_11484);
nand U12555 (N_12555,N_9579,N_11424);
or U12556 (N_12556,N_9761,N_9869);
and U12557 (N_12557,N_9200,N_10221);
nand U12558 (N_12558,N_10362,N_10055);
nand U12559 (N_12559,N_10879,N_11494);
nand U12560 (N_12560,N_11281,N_10498);
nand U12561 (N_12561,N_10589,N_11120);
nor U12562 (N_12562,N_9848,N_9953);
and U12563 (N_12563,N_10152,N_10409);
xnor U12564 (N_12564,N_10542,N_10854);
nand U12565 (N_12565,N_11855,N_11574);
xnor U12566 (N_12566,N_10160,N_10586);
or U12567 (N_12567,N_10027,N_11766);
or U12568 (N_12568,N_10054,N_10590);
xor U12569 (N_12569,N_11769,N_11939);
nor U12570 (N_12570,N_11215,N_11182);
or U12571 (N_12571,N_11101,N_11699);
and U12572 (N_12572,N_11265,N_9958);
xor U12573 (N_12573,N_10389,N_10895);
or U12574 (N_12574,N_10928,N_10902);
xnor U12575 (N_12575,N_10699,N_10418);
xnor U12576 (N_12576,N_9288,N_11463);
xnor U12577 (N_12577,N_9815,N_9961);
nand U12578 (N_12578,N_10746,N_10278);
or U12579 (N_12579,N_9300,N_11337);
or U12580 (N_12580,N_9705,N_11924);
nand U12581 (N_12581,N_10755,N_11231);
nand U12582 (N_12582,N_10795,N_11807);
or U12583 (N_12583,N_10087,N_10963);
or U12584 (N_12584,N_9157,N_11374);
xnor U12585 (N_12585,N_11315,N_9845);
nor U12586 (N_12586,N_10325,N_9406);
and U12587 (N_12587,N_10421,N_11881);
nor U12588 (N_12588,N_11595,N_10811);
or U12589 (N_12589,N_10580,N_10927);
xor U12590 (N_12590,N_11828,N_10343);
xor U12591 (N_12591,N_11731,N_9454);
xor U12592 (N_12592,N_9142,N_9878);
xor U12593 (N_12593,N_9372,N_10808);
nand U12594 (N_12594,N_11942,N_11724);
nor U12595 (N_12595,N_9425,N_11156);
or U12596 (N_12596,N_9254,N_11320);
or U12597 (N_12597,N_10082,N_11046);
xnor U12598 (N_12598,N_10925,N_10821);
xor U12599 (N_12599,N_10616,N_10737);
xnor U12600 (N_12600,N_9181,N_10400);
and U12601 (N_12601,N_10402,N_11441);
nor U12602 (N_12602,N_10273,N_11642);
and U12603 (N_12603,N_9189,N_9540);
nand U12604 (N_12604,N_9190,N_11562);
and U12605 (N_12605,N_11703,N_9457);
xor U12606 (N_12606,N_11174,N_11495);
or U12607 (N_12607,N_9752,N_10224);
or U12608 (N_12608,N_11734,N_10489);
or U12609 (N_12609,N_11788,N_10994);
or U12610 (N_12610,N_9619,N_9018);
nand U12611 (N_12611,N_10287,N_9443);
or U12612 (N_12612,N_11376,N_10481);
nand U12613 (N_12613,N_10701,N_9426);
nor U12614 (N_12614,N_9781,N_10036);
nand U12615 (N_12615,N_9285,N_11605);
or U12616 (N_12616,N_9605,N_9846);
nand U12617 (N_12617,N_9807,N_10607);
and U12618 (N_12618,N_9037,N_11064);
nand U12619 (N_12619,N_11885,N_9000);
nand U12620 (N_12620,N_9490,N_9864);
and U12621 (N_12621,N_11685,N_9823);
or U12622 (N_12622,N_9977,N_11168);
nor U12623 (N_12623,N_10556,N_9252);
xor U12624 (N_12624,N_9549,N_9746);
nand U12625 (N_12625,N_11056,N_9692);
and U12626 (N_12626,N_9420,N_10073);
and U12627 (N_12627,N_9563,N_10513);
or U12628 (N_12628,N_10157,N_11967);
nand U12629 (N_12629,N_10440,N_9371);
xor U12630 (N_12630,N_11911,N_10068);
xnor U12631 (N_12631,N_9123,N_10952);
or U12632 (N_12632,N_11372,N_10687);
or U12633 (N_12633,N_11959,N_11701);
and U12634 (N_12634,N_10957,N_11507);
and U12635 (N_12635,N_9657,N_10462);
and U12636 (N_12636,N_9798,N_11170);
and U12637 (N_12637,N_10255,N_10302);
or U12638 (N_12638,N_9404,N_9835);
or U12639 (N_12639,N_10769,N_10664);
nor U12640 (N_12640,N_9642,N_9971);
and U12641 (N_12641,N_10439,N_10700);
nand U12642 (N_12642,N_11389,N_11354);
nand U12643 (N_12643,N_10987,N_11359);
nor U12644 (N_12644,N_9110,N_11078);
and U12645 (N_12645,N_11710,N_9531);
or U12646 (N_12646,N_10024,N_11246);
xnor U12647 (N_12647,N_10019,N_11226);
nor U12648 (N_12648,N_11732,N_11071);
nor U12649 (N_12649,N_11092,N_10001);
nor U12650 (N_12650,N_9591,N_9922);
and U12651 (N_12651,N_10745,N_10861);
nand U12652 (N_12652,N_11597,N_11115);
and U12653 (N_12653,N_11586,N_9368);
nand U12654 (N_12654,N_10764,N_10304);
xor U12655 (N_12655,N_11829,N_11845);
nor U12656 (N_12656,N_10110,N_10965);
and U12657 (N_12657,N_9986,N_10646);
nand U12658 (N_12658,N_9069,N_10394);
and U12659 (N_12659,N_11601,N_10064);
nand U12660 (N_12660,N_10016,N_10667);
xnor U12661 (N_12661,N_10406,N_11459);
or U12662 (N_12662,N_9445,N_10593);
and U12663 (N_12663,N_11518,N_10725);
xor U12664 (N_12664,N_10058,N_11817);
and U12665 (N_12665,N_9957,N_11822);
or U12666 (N_12666,N_11145,N_9437);
or U12667 (N_12667,N_10277,N_9494);
nor U12668 (N_12668,N_11007,N_11555);
or U12669 (N_12669,N_11892,N_10692);
or U12670 (N_12670,N_10060,N_10799);
xor U12671 (N_12671,N_9610,N_11751);
and U12672 (N_12672,N_10801,N_10774);
nor U12673 (N_12673,N_10383,N_11969);
nor U12674 (N_12674,N_9121,N_11978);
xnor U12675 (N_12675,N_11568,N_9289);
nor U12676 (N_12676,N_9974,N_10074);
nor U12677 (N_12677,N_9309,N_9339);
and U12678 (N_12678,N_10508,N_10938);
xnor U12679 (N_12679,N_10754,N_11625);
or U12680 (N_12680,N_9363,N_9456);
or U12681 (N_12681,N_10197,N_9891);
and U12682 (N_12682,N_11532,N_11018);
or U12683 (N_12683,N_9754,N_11694);
nor U12684 (N_12684,N_11212,N_11417);
xor U12685 (N_12685,N_11030,N_10223);
nand U12686 (N_12686,N_9914,N_10852);
nor U12687 (N_12687,N_11199,N_10188);
xor U12688 (N_12688,N_11982,N_10740);
or U12689 (N_12689,N_11198,N_10334);
or U12690 (N_12690,N_11629,N_10204);
nand U12691 (N_12691,N_9489,N_10086);
nand U12692 (N_12692,N_9881,N_10326);
nor U12693 (N_12693,N_11658,N_11652);
and U12694 (N_12694,N_9946,N_9139);
nor U12695 (N_12695,N_11727,N_11127);
xnor U12696 (N_12696,N_10306,N_10324);
nand U12697 (N_12697,N_9478,N_10636);
or U12698 (N_12698,N_11038,N_11284);
nor U12699 (N_12699,N_9507,N_9284);
and U12700 (N_12700,N_9269,N_10753);
nand U12701 (N_12701,N_9074,N_9274);
nand U12702 (N_12702,N_9257,N_9768);
or U12703 (N_12703,N_9374,N_9213);
xor U12704 (N_12704,N_11104,N_10681);
and U12705 (N_12705,N_11243,N_11278);
xnor U12706 (N_12706,N_11878,N_9082);
or U12707 (N_12707,N_9060,N_11883);
xnor U12708 (N_12708,N_10824,N_11202);
nand U12709 (N_12709,N_9180,N_11058);
xor U12710 (N_12710,N_9344,N_10835);
nand U12711 (N_12711,N_10837,N_11489);
nand U12712 (N_12712,N_10167,N_11510);
nand U12713 (N_12713,N_9894,N_10052);
and U12714 (N_12714,N_11434,N_9602);
nor U12715 (N_12715,N_10407,N_10487);
and U12716 (N_12716,N_11074,N_9892);
nand U12717 (N_12717,N_10458,N_11446);
nand U12718 (N_12718,N_11893,N_9857);
or U12719 (N_12719,N_11399,N_11082);
nor U12720 (N_12720,N_9241,N_11062);
nand U12721 (N_12721,N_9575,N_9486);
nor U12722 (N_12722,N_10378,N_10829);
nor U12723 (N_12723,N_11877,N_10205);
xnor U12724 (N_12724,N_10116,N_9004);
and U12725 (N_12725,N_10708,N_9008);
nand U12726 (N_12726,N_10639,N_9509);
nor U12727 (N_12727,N_11765,N_11169);
or U12728 (N_12728,N_11659,N_10368);
or U12729 (N_12729,N_11119,N_10296);
xor U12730 (N_12730,N_10376,N_10807);
xnor U12731 (N_12731,N_9634,N_11945);
nand U12732 (N_12732,N_11820,N_9348);
nand U12733 (N_12733,N_9937,N_11958);
or U12734 (N_12734,N_10882,N_11425);
and U12735 (N_12735,N_9156,N_11794);
and U12736 (N_12736,N_10791,N_9192);
nand U12737 (N_12737,N_11396,N_11998);
nand U12738 (N_12738,N_9904,N_11847);
and U12739 (N_12739,N_9129,N_10388);
nand U12740 (N_12740,N_10941,N_9199);
and U12741 (N_12741,N_10408,N_10380);
xor U12742 (N_12742,N_11735,N_9927);
and U12743 (N_12743,N_10944,N_11971);
nor U12744 (N_12744,N_11733,N_9996);
nor U12745 (N_12745,N_10958,N_11256);
or U12746 (N_12746,N_11452,N_11839);
and U12747 (N_12747,N_11447,N_9093);
nand U12748 (N_12748,N_9655,N_11070);
xnor U12749 (N_12749,N_11857,N_10429);
nor U12750 (N_12750,N_9973,N_11730);
and U12751 (N_12751,N_9475,N_11849);
xor U12752 (N_12752,N_11024,N_10107);
or U12753 (N_12753,N_10682,N_9056);
or U12754 (N_12754,N_9872,N_9770);
and U12755 (N_12755,N_10235,N_11843);
xnor U12756 (N_12756,N_10806,N_10620);
nor U12757 (N_12757,N_10161,N_11868);
xor U12758 (N_12758,N_9477,N_11895);
or U12759 (N_12759,N_11992,N_11934);
xor U12760 (N_12760,N_11157,N_9913);
and U12761 (N_12761,N_10826,N_10231);
nor U12762 (N_12762,N_10838,N_10239);
or U12763 (N_12763,N_9615,N_10727);
xor U12764 (N_12764,N_11873,N_9013);
xnor U12765 (N_12765,N_10022,N_11690);
and U12766 (N_12766,N_10781,N_10229);
nand U12767 (N_12767,N_11301,N_11416);
or U12768 (N_12768,N_9338,N_10000);
nor U12769 (N_12769,N_9997,N_10547);
and U12770 (N_12770,N_9900,N_10320);
and U12771 (N_12771,N_11688,N_9677);
xnor U12772 (N_12772,N_10546,N_10671);
and U12773 (N_12773,N_10196,N_10367);
and U12774 (N_12774,N_9812,N_11340);
and U12775 (N_12775,N_10155,N_11474);
nand U12776 (N_12776,N_9947,N_10674);
nand U12777 (N_12777,N_11165,N_9925);
and U12778 (N_12778,N_10555,N_9141);
or U12779 (N_12779,N_9422,N_10527);
xnor U12780 (N_12780,N_11113,N_11218);
nand U12781 (N_12781,N_11589,N_10735);
nor U12782 (N_12782,N_11624,N_10728);
nand U12783 (N_12783,N_11047,N_9263);
xor U12784 (N_12784,N_9592,N_9007);
nor U12785 (N_12785,N_11229,N_10668);
nand U12786 (N_12786,N_11488,N_9438);
xor U12787 (N_12787,N_9373,N_9038);
and U12788 (N_12788,N_10606,N_9331);
nand U12789 (N_12789,N_9101,N_9972);
nor U12790 (N_12790,N_9945,N_9319);
nor U12791 (N_12791,N_11720,N_9023);
nand U12792 (N_12792,N_10541,N_11604);
and U12793 (N_12793,N_11838,N_11638);
xor U12794 (N_12794,N_9179,N_10848);
and U12795 (N_12795,N_9062,N_11462);
nand U12796 (N_12796,N_11187,N_11342);
or U12797 (N_12797,N_10743,N_10760);
and U12798 (N_12798,N_11477,N_9144);
nand U12799 (N_12799,N_11726,N_11523);
or U12800 (N_12800,N_9393,N_9860);
nand U12801 (N_12801,N_11686,N_10417);
xor U12802 (N_12802,N_9735,N_11487);
nor U12803 (N_12803,N_11936,N_9808);
nand U12804 (N_12804,N_10023,N_9095);
nand U12805 (N_12805,N_9162,N_11714);
or U12806 (N_12806,N_10482,N_11548);
nand U12807 (N_12807,N_11540,N_11194);
nor U12808 (N_12808,N_9128,N_9843);
nor U12809 (N_12809,N_10525,N_11771);
nand U12810 (N_12810,N_10684,N_10776);
nor U12811 (N_12811,N_10130,N_11316);
and U12812 (N_12812,N_10552,N_9583);
and U12813 (N_12813,N_10395,N_10056);
nand U12814 (N_12814,N_10006,N_10721);
xnor U12815 (N_12815,N_9463,N_11607);
xnor U12816 (N_12816,N_11650,N_9514);
and U12817 (N_12817,N_11105,N_10749);
nand U12818 (N_12818,N_10514,N_10932);
nand U12819 (N_12819,N_10717,N_9706);
or U12820 (N_12820,N_11013,N_11961);
or U12821 (N_12821,N_10194,N_9676);
xor U12822 (N_12822,N_11680,N_11995);
or U12823 (N_12823,N_11479,N_11783);
nor U12824 (N_12824,N_9195,N_10192);
nor U12825 (N_12825,N_10511,N_10163);
and U12826 (N_12826,N_9354,N_10379);
nor U12827 (N_12827,N_9882,N_11634);
nor U12828 (N_12828,N_9722,N_10382);
and U12829 (N_12829,N_10002,N_9759);
xor U12830 (N_12830,N_9664,N_11470);
and U12831 (N_12831,N_11615,N_9571);
nand U12832 (N_12832,N_11571,N_9969);
nor U12833 (N_12833,N_9644,N_11528);
xor U12834 (N_12834,N_11420,N_10531);
and U12835 (N_12835,N_10800,N_11110);
nand U12836 (N_12836,N_11290,N_9020);
and U12837 (N_12837,N_10272,N_11276);
or U12838 (N_12838,N_9276,N_11575);
or U12839 (N_12839,N_11118,N_10284);
and U12840 (N_12840,N_11296,N_10942);
nand U12841 (N_12841,N_11332,N_11456);
xnor U12842 (N_12842,N_9492,N_10009);
nor U12843 (N_12843,N_11854,N_9461);
and U12844 (N_12844,N_10123,N_9939);
xnor U12845 (N_12845,N_11664,N_9148);
nor U12846 (N_12846,N_11214,N_9087);
xor U12847 (N_12847,N_9234,N_9650);
xor U12848 (N_12848,N_11430,N_11271);
xnor U12849 (N_12849,N_9620,N_11287);
nor U12850 (N_12850,N_9720,N_9980);
nor U12851 (N_12851,N_10978,N_9377);
xnor U12852 (N_12852,N_9790,N_11790);
nand U12853 (N_12853,N_10650,N_10827);
xor U12854 (N_12854,N_9317,N_9526);
nor U12855 (N_12855,N_10085,N_9203);
and U12856 (N_12856,N_10813,N_10783);
or U12857 (N_12857,N_9833,N_9976);
nand U12858 (N_12858,N_10595,N_10859);
nand U12859 (N_12859,N_9902,N_10669);
nand U12860 (N_12860,N_10689,N_11789);
nand U12861 (N_12861,N_11210,N_10996);
and U12862 (N_12862,N_10844,N_9078);
nor U12863 (N_12863,N_10632,N_9581);
and U12864 (N_12864,N_11026,N_11017);
nor U12865 (N_12865,N_9154,N_9016);
nor U12866 (N_12866,N_9599,N_9167);
xnor U12867 (N_12867,N_11899,N_10293);
and U12868 (N_12868,N_9107,N_11401);
xnor U12869 (N_12869,N_10118,N_9888);
nor U12870 (N_12870,N_9416,N_11503);
xnor U12871 (N_12871,N_11383,N_10430);
nand U12872 (N_12872,N_10984,N_10986);
nor U12873 (N_12873,N_10217,N_11867);
xnor U12874 (N_12874,N_10494,N_11983);
nor U12875 (N_12875,N_9215,N_9661);
and U12876 (N_12876,N_9794,N_9019);
and U12877 (N_12877,N_11011,N_9999);
xor U12878 (N_12878,N_11558,N_10985);
or U12879 (N_12879,N_10972,N_11657);
xnor U12880 (N_12880,N_10784,N_9555);
nand U12881 (N_12881,N_11275,N_9989);
nor U12882 (N_12882,N_10767,N_10660);
or U12883 (N_12883,N_10295,N_9694);
or U12884 (N_12884,N_10184,N_11312);
xor U12885 (N_12885,N_9369,N_11217);
or U12886 (N_12886,N_11862,N_10576);
nor U12887 (N_12887,N_10254,N_9983);
nor U12888 (N_12888,N_9926,N_9918);
nand U12889 (N_12889,N_10310,N_10125);
and U12890 (N_12890,N_11164,N_10353);
or U12891 (N_12891,N_10540,N_10041);
or U12892 (N_12892,N_10112,N_9899);
and U12893 (N_12893,N_10698,N_11673);
or U12894 (N_12894,N_11874,N_10359);
nand U12895 (N_12895,N_9955,N_11472);
or U12896 (N_12896,N_11526,N_10106);
xor U12897 (N_12897,N_10579,N_9632);
and U12898 (N_12898,N_10909,N_9033);
nand U12899 (N_12899,N_11813,N_10132);
nor U12900 (N_12900,N_11946,N_10887);
xor U12901 (N_12901,N_11079,N_10666);
or U12902 (N_12902,N_10142,N_10648);
or U12903 (N_12903,N_9909,N_10690);
xnor U12904 (N_12904,N_10171,N_9450);
and U12905 (N_12905,N_10499,N_11189);
or U12906 (N_12906,N_10762,N_11319);
nor U12907 (N_12907,N_10341,N_11364);
or U12908 (N_12908,N_11075,N_9767);
xor U12909 (N_12909,N_11067,N_9701);
or U12910 (N_12910,N_11918,N_11665);
or U12911 (N_12911,N_11772,N_9452);
and U12912 (N_12912,N_11250,N_9005);
or U12913 (N_12913,N_9943,N_11003);
or U12914 (N_12914,N_10300,N_11593);
nand U12915 (N_12915,N_9744,N_11422);
or U12916 (N_12916,N_11496,N_11326);
nor U12917 (N_12917,N_11028,N_9327);
or U12918 (N_12918,N_9424,N_11609);
nor U12919 (N_12919,N_9842,N_11005);
nand U12920 (N_12920,N_11436,N_11706);
nor U12921 (N_12921,N_9604,N_9481);
or U12922 (N_12922,N_9342,N_9025);
nor U12923 (N_12923,N_11764,N_9879);
or U12924 (N_12924,N_10309,N_11195);
or U12925 (N_12925,N_10456,N_11036);
xor U12926 (N_12926,N_11833,N_9799);
and U12927 (N_12927,N_10377,N_10139);
xor U12928 (N_12928,N_9134,N_11039);
and U12929 (N_12929,N_10507,N_9867);
nand U12930 (N_12930,N_9883,N_9783);
and U12931 (N_12931,N_11520,N_9255);
and U12932 (N_12932,N_10436,N_9929);
or U12933 (N_12933,N_11653,N_11512);
xor U12934 (N_12934,N_11707,N_10990);
or U12935 (N_12935,N_9774,N_10271);
nor U12936 (N_12936,N_9086,N_10018);
and U12937 (N_12937,N_10558,N_9561);
nand U12938 (N_12938,N_10501,N_11620);
or U12939 (N_12939,N_10707,N_9009);
and U12940 (N_12940,N_9952,N_9975);
nand U12941 (N_12941,N_11140,N_11596);
nor U12942 (N_12942,N_9779,N_11266);
nor U12943 (N_12943,N_9244,N_10676);
and U12944 (N_12944,N_9480,N_9565);
or U12945 (N_12945,N_9089,N_10075);
and U12946 (N_12946,N_9868,N_10973);
nand U12947 (N_12947,N_9827,N_9698);
or U12948 (N_12948,N_10364,N_9513);
nor U12949 (N_12949,N_9102,N_11785);
and U12950 (N_12950,N_9643,N_10170);
nand U12951 (N_12951,N_11191,N_9502);
nand U12952 (N_12952,N_11471,N_9832);
or U12953 (N_12953,N_11476,N_10374);
and U12954 (N_12954,N_11356,N_11180);
or U12955 (N_12955,N_10891,N_9923);
nand U12956 (N_12956,N_9260,N_11428);
and U12957 (N_12957,N_11482,N_10177);
and U12958 (N_12958,N_10868,N_10775);
xor U12959 (N_12959,N_9361,N_11944);
nor U12960 (N_12960,N_11888,N_10138);
xnor U12961 (N_12961,N_11371,N_11818);
and U12962 (N_12962,N_10930,N_11861);
and U12963 (N_12963,N_10967,N_10656);
nor U12964 (N_12964,N_9717,N_10899);
and U12965 (N_12965,N_10773,N_11128);
nor U12966 (N_12966,N_10948,N_10961);
nand U12967 (N_12967,N_9587,N_10867);
or U12968 (N_12968,N_10977,N_11095);
xor U12969 (N_12969,N_10083,N_11277);
and U12970 (N_12970,N_9820,N_10734);
or U12971 (N_12971,N_11580,N_11025);
nand U12972 (N_12972,N_11744,N_10212);
nor U12973 (N_12973,N_10686,N_9442);
xor U12974 (N_12974,N_9299,N_10992);
xnor U12975 (N_12975,N_10843,N_10330);
nand U12976 (N_12976,N_9524,N_9760);
or U12977 (N_12977,N_9645,N_9311);
nor U12978 (N_12978,N_9640,N_9127);
xor U12979 (N_12979,N_9398,N_10706);
xnor U12980 (N_12980,N_9542,N_9633);
nand U12981 (N_12981,N_9399,N_9125);
or U12982 (N_12982,N_9841,N_10845);
xnor U12983 (N_12983,N_10431,N_10538);
and U12984 (N_12984,N_10172,N_11865);
or U12985 (N_12985,N_10465,N_9126);
or U12986 (N_12986,N_11760,N_11144);
and U12987 (N_12987,N_10031,N_11859);
nor U12988 (N_12988,N_9030,N_10384);
xnor U12989 (N_12989,N_10641,N_9763);
nand U12990 (N_12990,N_11561,N_11449);
nor U12991 (N_12991,N_11325,N_9938);
or U12992 (N_12992,N_11175,N_11999);
or U12993 (N_12993,N_9537,N_9749);
nand U12994 (N_12994,N_9851,N_10179);
xor U12995 (N_12995,N_11698,N_11608);
xnor U12996 (N_12996,N_9740,N_11171);
and U12997 (N_12997,N_10503,N_11577);
and U12998 (N_12998,N_10092,N_10956);
or U12999 (N_12999,N_10747,N_11020);
or U13000 (N_13000,N_10335,N_10495);
and U13001 (N_13001,N_10592,N_11588);
nor U13002 (N_13002,N_11279,N_9026);
xnor U13003 (N_13003,N_10672,N_9027);
xor U13004 (N_13004,N_10712,N_9681);
and U13005 (N_13005,N_9394,N_9764);
nand U13006 (N_13006,N_11148,N_11508);
or U13007 (N_13007,N_10090,N_10997);
nor U13008 (N_13008,N_11692,N_10657);
and U13009 (N_13009,N_9737,N_11465);
and U13010 (N_13010,N_10566,N_11394);
nand U13011 (N_13011,N_9113,N_9356);
or U13012 (N_13012,N_10372,N_10815);
and U13013 (N_13013,N_9010,N_11386);
xor U13014 (N_13014,N_11663,N_11438);
and U13015 (N_13015,N_11687,N_9597);
xor U13016 (N_13016,N_10120,N_11138);
nand U13017 (N_13017,N_10526,N_9850);
or U13018 (N_13018,N_9143,N_10307);
nand U13019 (N_13019,N_10460,N_9149);
xor U13020 (N_13020,N_11926,N_10084);
nor U13021 (N_13021,N_9293,N_10559);
and U13022 (N_13022,N_9383,N_9924);
and U13023 (N_13023,N_9250,N_9446);
and U13024 (N_13024,N_9685,N_9172);
nor U13025 (N_13025,N_10638,N_9775);
nor U13026 (N_13026,N_10529,N_10765);
nor U13027 (N_13027,N_10534,N_10093);
nand U13028 (N_13028,N_9817,N_10442);
nand U13029 (N_13029,N_11780,N_9991);
or U13030 (N_13030,N_9415,N_9553);
xnor U13031 (N_13031,N_11514,N_10505);
nand U13032 (N_13032,N_9503,N_10438);
nor U13033 (N_13033,N_11773,N_10557);
or U13034 (N_13034,N_11311,N_11986);
or U13035 (N_13035,N_9229,N_9385);
xnor U13036 (N_13036,N_10319,N_11059);
nor U13037 (N_13037,N_9521,N_10454);
and U13038 (N_13038,N_11373,N_9784);
and U13039 (N_13039,N_10128,N_11853);
xor U13040 (N_13040,N_11880,N_10119);
nand U13041 (N_13041,N_9921,N_9021);
nand U13042 (N_13042,N_11264,N_10015);
nor U13043 (N_13043,N_11776,N_10397);
and U13044 (N_13044,N_10218,N_10726);
nand U13045 (N_13045,N_11700,N_9726);
and U13046 (N_13046,N_11443,N_10136);
and U13047 (N_13047,N_9091,N_10010);
and U13048 (N_13048,N_11057,N_9390);
xor U13049 (N_13049,N_9538,N_10828);
and U13050 (N_13050,N_9528,N_10768);
nor U13051 (N_13051,N_10778,N_11956);
nor U13052 (N_13052,N_9624,N_10924);
nand U13053 (N_13053,N_11318,N_11227);
and U13054 (N_13054,N_10097,N_9336);
xor U13055 (N_13055,N_10238,N_10246);
nor U13056 (N_13056,N_9085,N_11253);
nand U13057 (N_13057,N_10347,N_11875);
nand U13058 (N_13058,N_10115,N_9006);
nor U13059 (N_13059,N_10772,N_9594);
nor U13060 (N_13060,N_11378,N_11213);
or U13061 (N_13061,N_9660,N_10312);
nand U13062 (N_13062,N_10230,N_10297);
nand U13063 (N_13063,N_11626,N_11023);
and U13064 (N_13064,N_10342,N_10349);
or U13065 (N_13065,N_10301,N_11044);
or U13066 (N_13066,N_10345,N_10553);
nor U13067 (N_13067,N_11929,N_9627);
xnor U13068 (N_13068,N_9366,N_10865);
nand U13069 (N_13069,N_10366,N_11481);
or U13070 (N_13070,N_11135,N_9721);
or U13071 (N_13071,N_9096,N_9119);
or U13072 (N_13072,N_10788,N_11948);
or U13073 (N_13073,N_9351,N_9444);
xnor U13074 (N_13074,N_10771,N_9628);
xor U13075 (N_13075,N_10864,N_10333);
nor U13076 (N_13076,N_9237,N_10043);
or U13077 (N_13077,N_10937,N_9071);
or U13078 (N_13078,N_11906,N_10398);
nand U13079 (N_13079,N_10164,N_10321);
xnor U13080 (N_13080,N_9230,N_10189);
nor U13081 (N_13081,N_11633,N_9582);
nand U13082 (N_13082,N_10485,N_11955);
or U13083 (N_13083,N_11330,N_10933);
and U13084 (N_13084,N_10906,N_9451);
nor U13085 (N_13085,N_9711,N_9075);
nor U13086 (N_13086,N_9988,N_11981);
nand U13087 (N_13087,N_11913,N_10841);
xnor U13088 (N_13088,N_11953,N_9279);
and U13089 (N_13089,N_9118,N_11979);
nand U13090 (N_13090,N_9294,N_10370);
and U13091 (N_13091,N_10894,N_11302);
and U13092 (N_13092,N_11393,N_10405);
nand U13093 (N_13093,N_10970,N_9150);
nand U13094 (N_13094,N_9099,N_9340);
nand U13095 (N_13095,N_11761,N_9668);
nand U13096 (N_13096,N_10855,N_9484);
xor U13097 (N_13097,N_11932,N_9335);
xor U13098 (N_13098,N_9111,N_9401);
xnor U13099 (N_13099,N_9232,N_9831);
or U13100 (N_13100,N_11940,N_10451);
xor U13101 (N_13101,N_11993,N_9612);
or U13102 (N_13102,N_10522,N_9275);
xnor U13103 (N_13103,N_9225,N_9330);
nand U13104 (N_13104,N_11920,N_11506);
nor U13105 (N_13105,N_9397,N_10190);
xor U13106 (N_13106,N_10173,N_9431);
xnor U13107 (N_13107,N_10943,N_9816);
nand U13108 (N_13108,N_11358,N_10599);
xnor U13109 (N_13109,N_9419,N_10763);
and U13110 (N_13110,N_10423,N_10490);
and U13111 (N_13111,N_10270,N_11299);
and U13112 (N_13112,N_10061,N_10003);
or U13113 (N_13113,N_11834,N_11001);
and U13114 (N_13114,N_10199,N_11400);
nand U13115 (N_13115,N_9569,N_10026);
and U13116 (N_13116,N_11823,N_10165);
xor U13117 (N_13117,N_11759,N_11102);
and U13118 (N_13118,N_11486,N_9636);
or U13119 (N_13119,N_9950,N_11876);
and U13120 (N_13120,N_11824,N_11927);
xor U13121 (N_13121,N_9896,N_10149);
xor U13122 (N_13122,N_11100,N_10914);
xnor U13123 (N_13123,N_10340,N_9039);
or U13124 (N_13124,N_9780,N_10757);
nor U13125 (N_13125,N_11019,N_10729);
and U13126 (N_13126,N_9589,N_9608);
and U13127 (N_13127,N_10259,N_10817);
xnor U13128 (N_13128,N_11109,N_10444);
nor U13129 (N_13129,N_10832,N_9557);
nand U13130 (N_13130,N_11670,N_9059);
and U13131 (N_13131,N_9523,N_11984);
and U13132 (N_13132,N_11914,N_11793);
nand U13133 (N_13133,N_11559,N_11049);
nand U13134 (N_13134,N_11408,N_10908);
nand U13135 (N_13135,N_10694,N_9638);
and U13136 (N_13136,N_9559,N_11639);
nand U13137 (N_13137,N_11980,N_10719);
xor U13138 (N_13138,N_9474,N_11327);
xor U13139 (N_13139,N_10047,N_10659);
xnor U13140 (N_13140,N_10578,N_10089);
or U13141 (N_13141,N_9826,N_11671);
xor U13142 (N_13142,N_11889,N_11045);
and U13143 (N_13143,N_9584,N_11261);
nor U13144 (N_13144,N_9536,N_11504);
nor U13145 (N_13145,N_10399,N_11763);
and U13146 (N_13146,N_10028,N_11808);
or U13147 (N_13147,N_9603,N_9670);
nand U13148 (N_13148,N_10523,N_10168);
nor U13149 (N_13149,N_10782,N_9796);
nor U13150 (N_13150,N_10065,N_9427);
or U13151 (N_13151,N_11672,N_10117);
nand U13152 (N_13152,N_10691,N_9145);
nor U13153 (N_13153,N_10285,N_10615);
xnor U13154 (N_13154,N_11669,N_9184);
and U13155 (N_13155,N_9245,N_10851);
xnor U13156 (N_13156,N_10298,N_10623);
and U13157 (N_13157,N_9573,N_9625);
xor U13158 (N_13158,N_10216,N_9303);
or U13159 (N_13159,N_9500,N_11907);
and U13160 (N_13160,N_11106,N_9267);
and U13161 (N_13161,N_9473,N_10274);
nor U13162 (N_13162,N_9440,N_9076);
nor U13163 (N_13163,N_11767,N_11096);
nand U13164 (N_13164,N_9708,N_9349);
and U13165 (N_13165,N_11475,N_9214);
xnor U13166 (N_13166,N_9479,N_9755);
nor U13167 (N_13167,N_10564,N_10897);
or U13168 (N_13168,N_10014,N_9488);
and U13169 (N_13169,N_9052,N_10923);
and U13170 (N_13170,N_11631,N_10738);
xnor U13171 (N_13171,N_11800,N_10477);
and U13172 (N_13172,N_10792,N_11921);
xnor U13173 (N_13173,N_11925,N_10872);
xor U13174 (N_13174,N_9228,N_9487);
nor U13175 (N_13175,N_11492,N_9297);
or U13176 (N_13176,N_9810,N_11533);
nand U13177 (N_13177,N_10180,N_10233);
and U13178 (N_13178,N_11392,N_9710);
xnor U13179 (N_13179,N_10332,N_10492);
nor U13180 (N_13180,N_11233,N_11738);
nand U13181 (N_13181,N_11884,N_9854);
nand U13182 (N_13182,N_9090,N_11493);
xor U13183 (N_13183,N_11242,N_11313);
or U13184 (N_13184,N_10127,N_11516);
and U13185 (N_13185,N_9919,N_11108);
nand U13186 (N_13186,N_9505,N_10678);
and U13187 (N_13187,N_11717,N_11453);
nand U13188 (N_13188,N_9350,N_10113);
and U13189 (N_13189,N_11041,N_9175);
and U13190 (N_13190,N_9825,N_10758);
and U13191 (N_13191,N_11258,N_11483);
nor U13192 (N_13192,N_11152,N_9678);
and U13193 (N_13193,N_9837,N_11445);
nor U13194 (N_13194,N_9047,N_10999);
xor U13195 (N_13195,N_11429,N_9562);
and U13196 (N_13196,N_11621,N_10532);
xor U13197 (N_13197,N_10263,N_10512);
and U13198 (N_13198,N_11379,N_11850);
nand U13199 (N_13199,N_11398,N_10926);
nand U13200 (N_13200,N_11335,N_11043);
xor U13201 (N_13201,N_11660,N_11388);
xor U13202 (N_13202,N_10519,N_11666);
or U13203 (N_13203,N_11848,N_10435);
and U13204 (N_13204,N_11085,N_11708);
and U13205 (N_13205,N_11715,N_10446);
nor U13206 (N_13206,N_9750,N_9176);
and U13207 (N_13207,N_9948,N_10225);
nand U13208 (N_13208,N_10568,N_10587);
and U13209 (N_13209,N_9782,N_10466);
xor U13210 (N_13210,N_9772,N_9205);
and U13211 (N_13211,N_9648,N_10922);
xor U13212 (N_13212,N_10724,N_11291);
or U13213 (N_13213,N_9003,N_10918);
nor U13214 (N_13214,N_10543,N_9449);
and U13215 (N_13215,N_9353,N_9493);
nor U13216 (N_13216,N_11651,N_11412);
and U13217 (N_13217,N_11361,N_10642);
xor U13218 (N_13218,N_9858,N_9800);
xnor U13219 (N_13219,N_9170,N_9462);
nor U13220 (N_13220,N_11134,N_9307);
nor U13221 (N_13221,N_9053,N_9876);
nor U13222 (N_13222,N_10567,N_11081);
xnor U13223 (N_13223,N_9753,N_9889);
nand U13224 (N_13224,N_10414,N_9533);
nor U13225 (N_13225,N_11205,N_10403);
xor U13226 (N_13226,N_11251,N_10159);
xnor U13227 (N_13227,N_10693,N_10969);
nor U13228 (N_13228,N_9546,N_10262);
nor U13229 (N_13229,N_11444,N_10447);
or U13230 (N_13230,N_10354,N_9539);
or U13231 (N_13231,N_11614,N_10209);
nor U13232 (N_13232,N_9741,N_10643);
and U13233 (N_13233,N_10870,N_10955);
or U13234 (N_13234,N_11161,N_10823);
xor U13235 (N_13235,N_10988,N_10858);
nand U13236 (N_13236,N_10258,N_9525);
or U13237 (N_13237,N_11448,N_10232);
and U13238 (N_13238,N_11150,N_11758);
nor U13239 (N_13239,N_9088,N_10029);
and U13240 (N_13240,N_9467,N_9332);
nor U13241 (N_13241,N_9174,N_11037);
nor U13242 (N_13242,N_11796,N_9050);
or U13243 (N_13243,N_11244,N_11126);
or U13244 (N_13244,N_9155,N_10602);
or U13245 (N_13245,N_11068,N_9912);
nor U13246 (N_13246,N_11702,N_11705);
and U13247 (N_13247,N_9570,N_9614);
and U13248 (N_13248,N_11139,N_11908);
or U13249 (N_13249,N_9218,N_9246);
xor U13250 (N_13250,N_10962,N_11322);
and U13251 (N_13251,N_10736,N_10940);
nor U13252 (N_13252,N_9100,N_10488);
or U13253 (N_13253,N_9163,N_10208);
nand U13254 (N_13254,N_11560,N_10040);
or U13255 (N_13255,N_9967,N_11116);
nand U13256 (N_13256,N_11131,N_10081);
nand U13257 (N_13257,N_9465,N_11825);
or U13258 (N_13258,N_11407,N_11098);
or U13259 (N_13259,N_10761,N_11534);
nand U13260 (N_13260,N_10288,N_11339);
and U13261 (N_13261,N_9221,N_9517);
and U13262 (N_13262,N_10975,N_11887);
or U13263 (N_13263,N_10585,N_10280);
or U13264 (N_13264,N_10718,N_11695);
nor U13265 (N_13265,N_11627,N_9265);
xor U13266 (N_13266,N_10617,N_11151);
xnor U13267 (N_13267,N_11221,N_10751);
or U13268 (N_13268,N_10951,N_11797);
nand U13269 (N_13269,N_10633,N_9407);
nor U13270 (N_13270,N_11387,N_9960);
xnor U13271 (N_13271,N_11111,N_10363);
nor U13272 (N_13272,N_11831,N_9646);
and U13273 (N_13273,N_10954,N_9686);
or U13274 (N_13274,N_10479,N_11784);
nor U13275 (N_13275,N_9283,N_11960);
and U13276 (N_13276,N_9665,N_11499);
nor U13277 (N_13277,N_10228,N_9739);
and U13278 (N_13278,N_11216,N_9032);
nand U13279 (N_13279,N_10011,N_10038);
or U13280 (N_13280,N_9223,N_10818);
and U13281 (N_13281,N_9253,N_11696);
nor U13282 (N_13282,N_9140,N_11093);
nor U13283 (N_13283,N_11451,N_11557);
nand U13284 (N_13284,N_9829,N_9733);
nand U13285 (N_13285,N_10412,N_11433);
or U13286 (N_13286,N_10478,N_10759);
and U13287 (N_13287,N_9855,N_11718);
xnor U13288 (N_13288,N_9932,N_9606);
and U13289 (N_13289,N_9566,N_11014);
nor U13290 (N_13290,N_10766,N_10750);
nand U13291 (N_13291,N_11048,N_10597);
or U13292 (N_13292,N_11777,N_9173);
xor U13293 (N_13293,N_9618,N_9054);
nand U13294 (N_13294,N_11736,N_9365);
nor U13295 (N_13295,N_10129,N_9743);
nand U13296 (N_13296,N_9291,N_9863);
and U13297 (N_13297,N_11343,N_10114);
or U13298 (N_13298,N_10434,N_9378);
nor U13299 (N_13299,N_11406,N_9572);
nor U13300 (N_13300,N_10294,N_9659);
xor U13301 (N_13301,N_11298,N_9278);
nand U13302 (N_13302,N_10151,N_9328);
nand U13303 (N_13303,N_11681,N_11381);
and U13304 (N_13304,N_10790,N_9412);
xor U13305 (N_13305,N_11147,N_9885);
and U13306 (N_13306,N_10601,N_11827);
nand U13307 (N_13307,N_9224,N_11080);
nor U13308 (N_13308,N_9413,N_11054);
nand U13309 (N_13309,N_10290,N_10680);
or U13310 (N_13310,N_11166,N_9672);
nand U13311 (N_13311,N_9547,N_11872);
xor U13312 (N_13312,N_10328,N_10240);
nand U13313 (N_13313,N_11450,N_9824);
nor U13314 (N_13314,N_11632,N_10950);
and U13315 (N_13315,N_11603,N_11564);
or U13316 (N_13316,N_11919,N_11655);
and U13317 (N_13317,N_10502,N_9551);
nor U13318 (N_13318,N_9954,N_10797);
xor U13319 (N_13319,N_9070,N_9432);
or U13320 (N_13320,N_11756,N_10929);
nor U13321 (N_13321,N_9337,N_9386);
or U13322 (N_13322,N_10846,N_9308);
xnor U13323 (N_13323,N_11930,N_10662);
xor U13324 (N_13324,N_9259,N_9428);
xnor U13325 (N_13325,N_9666,N_11565);
or U13326 (N_13326,N_9057,N_9171);
and U13327 (N_13327,N_11752,N_10311);
xnor U13328 (N_13328,N_10257,N_11985);
and U13329 (N_13329,N_10630,N_9418);
or U13330 (N_13330,N_9959,N_11782);
nor U13331 (N_13331,N_11382,N_9728);
or U13332 (N_13332,N_10281,N_9765);
xnor U13333 (N_13333,N_11303,N_10201);
and U13334 (N_13334,N_11158,N_9732);
or U13335 (N_13335,N_10437,N_11252);
xor U13336 (N_13336,N_10420,N_11952);
or U13337 (N_13337,N_9238,N_9046);
nor U13338 (N_13338,N_10886,N_10979);
xnor U13339 (N_13339,N_9084,N_9014);
nor U13340 (N_13340,N_10836,N_9258);
or U13341 (N_13341,N_11201,N_11544);
nand U13342 (N_13342,N_9691,N_10869);
nand U13343 (N_13343,N_9158,N_10071);
nor U13344 (N_13344,N_10453,N_11159);
or U13345 (N_13345,N_10709,N_9600);
xnor U13346 (N_13346,N_10702,N_9940);
or U13347 (N_13347,N_9364,N_10289);
nand U13348 (N_13348,N_11365,N_10352);
xor U13349 (N_13349,N_11245,N_9219);
nand U13350 (N_13350,N_10393,N_11826);
or U13351 (N_13351,N_11130,N_11323);
nand U13352 (N_13352,N_10609,N_11060);
and U13353 (N_13353,N_11798,N_9532);
nor U13354 (N_13354,N_11268,N_10562);
nor U13355 (N_13355,N_10101,N_10980);
and U13356 (N_13356,N_9065,N_11719);
nand U13357 (N_13357,N_10178,N_11162);
and U13358 (N_13358,N_9436,N_11370);
xor U13359 (N_13359,N_10971,N_10710);
xor U13360 (N_13360,N_11970,N_11008);
and U13361 (N_13361,N_10756,N_11988);
xnor U13362 (N_13362,N_10705,N_10742);
xor U13363 (N_13363,N_9653,N_11816);
or U13364 (N_13364,N_9874,N_11676);
xnor U13365 (N_13365,N_10631,N_11307);
and U13366 (N_13366,N_9773,N_10665);
or U13367 (N_13367,N_11073,N_10787);
xor U13368 (N_13368,N_9736,N_11749);
and U13369 (N_13369,N_9771,N_9429);
xor U13370 (N_13370,N_11133,N_11289);
or U13371 (N_13371,N_11552,N_11866);
and U13372 (N_13372,N_11419,N_11903);
and U13373 (N_13373,N_9578,N_9518);
or U13374 (N_13374,N_9458,N_11628);
xnor U13375 (N_13375,N_11136,N_9496);
xor U13376 (N_13376,N_9725,N_9930);
xor U13377 (N_13377,N_11584,N_9623);
nor U13378 (N_13378,N_10624,N_10256);
nor U13379 (N_13379,N_11254,N_9212);
and U13380 (N_13380,N_9576,N_11464);
nand U13381 (N_13381,N_9347,N_11677);
nand U13382 (N_13382,N_9301,N_10696);
nand U13383 (N_13383,N_10247,N_10470);
nand U13384 (N_13384,N_10243,N_11740);
nand U13385 (N_13385,N_10203,N_11352);
xnor U13386 (N_13386,N_9830,N_11478);
and U13387 (N_13387,N_10898,N_9159);
xor U13388 (N_13388,N_10905,N_11500);
xor U13389 (N_13389,N_10677,N_11468);
nand U13390 (N_13390,N_11541,N_11697);
xor U13391 (N_13391,N_11563,N_10515);
nor U13392 (N_13392,N_11262,N_9586);
or U13393 (N_13393,N_11935,N_9847);
nand U13394 (N_13394,N_11112,N_10419);
xor U13395 (N_13395,N_11645,N_9360);
and U13396 (N_13396,N_10533,N_9261);
nor U13397 (N_13397,N_11305,N_10210);
nand U13398 (N_13398,N_9556,N_11933);
xor U13399 (N_13399,N_9051,N_9671);
xnor U13400 (N_13400,N_10242,N_9208);
or U13401 (N_13401,N_9120,N_11395);
nand U13402 (N_13402,N_11501,N_11576);
and U13403 (N_13403,N_9658,N_11778);
nand U13404 (N_13404,N_9104,N_10411);
nand U13405 (N_13405,N_10153,N_11801);
and U13406 (N_13406,N_9132,N_11842);
or U13407 (N_13407,N_9541,N_9392);
or U13408 (N_13408,N_10303,N_9197);
xnor U13409 (N_13409,N_11582,N_9165);
nor U13410 (N_13410,N_10517,N_9979);
nor U13411 (N_13411,N_9262,N_10375);
nor U13412 (N_13412,N_9298,N_9554);
nor U13413 (N_13413,N_11016,N_11431);
nor U13414 (N_13414,N_9742,N_10150);
nor U13415 (N_13415,N_9984,N_11973);
or U13416 (N_13416,N_10911,N_9485);
nand U13417 (N_13417,N_11781,N_10715);
nand U13418 (N_13418,N_10722,N_10491);
xnor U13419 (N_13419,N_9108,N_10069);
and U13420 (N_13420,N_10900,N_11426);
nand U13421 (N_13421,N_11076,N_9277);
xor U13422 (N_13422,N_10509,N_9177);
nor U13423 (N_13423,N_11583,N_9209);
xnor U13424 (N_13424,N_9682,N_9222);
or U13425 (N_13425,N_10804,N_9844);
and U13426 (N_13426,N_9802,N_10286);
and U13427 (N_13427,N_10654,N_9264);
or U13428 (N_13428,N_10573,N_11208);
or U13429 (N_13429,N_10862,N_11739);
nor U13430 (N_13430,N_11830,N_9690);
nor U13431 (N_13431,N_9617,N_11640);
nand U13432 (N_13432,N_11542,N_10291);
or U13433 (N_13433,N_11285,N_9055);
nor U13434 (N_13434,N_11799,N_9936);
xor U13435 (N_13435,N_11837,N_11856);
or U13436 (N_13436,N_11950,N_10814);
and U13437 (N_13437,N_11987,N_9828);
and U13438 (N_13438,N_10033,N_10253);
nor U13439 (N_13439,N_10020,N_10608);
xor U13440 (N_13440,N_9325,N_9080);
nand U13441 (N_13441,N_11235,N_11308);
and U13442 (N_13442,N_11550,N_11418);
or U13443 (N_13443,N_11088,N_11263);
xor U13444 (N_13444,N_10802,N_11027);
and U13445 (N_13445,N_10244,N_11691);
or U13446 (N_13446,N_11709,N_11397);
nand U13447 (N_13447,N_10486,N_10008);
and U13448 (N_13448,N_11222,N_10049);
nor U13449 (N_13449,N_9169,N_10834);
xor U13450 (N_13450,N_9146,N_9414);
nand U13451 (N_13451,N_11069,N_9637);
and U13452 (N_13452,N_9206,N_9766);
and U13453 (N_13453,N_11437,N_9716);
and U13454 (N_13454,N_9318,N_10622);
and U13455 (N_13455,N_11646,N_10104);
nand U13456 (N_13456,N_10464,N_10856);
nor U13457 (N_13457,N_9391,N_9520);
or U13458 (N_13458,N_11248,N_9714);
xor U13459 (N_13459,N_11141,N_11160);
nand U13460 (N_13460,N_9153,N_9942);
nand U13461 (N_13461,N_10365,N_9116);
and U13462 (N_13462,N_11021,N_10596);
and U13463 (N_13463,N_10504,N_11590);
and U13464 (N_13464,N_10860,N_10211);
nor U13465 (N_13465,N_9564,N_9322);
and U13466 (N_13466,N_10476,N_11860);
nand U13467 (N_13467,N_9185,N_10703);
and U13468 (N_13468,N_11114,N_9731);
and U13469 (N_13469,N_10888,N_11353);
and U13470 (N_13470,N_9321,N_9917);
xor U13471 (N_13471,N_10744,N_11410);
or U13472 (N_13472,N_9305,N_11754);
or U13473 (N_13473,N_10731,N_11618);
and U13474 (N_13474,N_11786,N_11015);
and U13475 (N_13475,N_9287,N_11414);
xor U13476 (N_13476,N_9239,N_9389);
and U13477 (N_13477,N_11594,N_10510);
and U13478 (N_13478,N_11886,N_11442);
xnor U13479 (N_13479,N_10053,N_9852);
nand U13480 (N_13480,N_10175,N_10516);
nand U13481 (N_13481,N_9117,N_10062);
xor U13482 (N_13482,N_11851,N_10995);
nor U13483 (N_13483,N_10959,N_11745);
xor U13484 (N_13484,N_9103,N_11890);
xor U13485 (N_13485,N_9272,N_9621);
nor U13486 (N_13486,N_10704,N_9792);
xnor U13487 (N_13487,N_9651,N_9667);
nor U13488 (N_13488,N_10614,N_9081);
or U13489 (N_13489,N_10070,N_10338);
nor U13490 (N_13490,N_9703,N_11022);
nand U13491 (N_13491,N_9545,N_10551);
xnor U13492 (N_13492,N_10917,N_9273);
or U13493 (N_13493,N_11556,N_10673);
nor U13494 (N_13494,N_10537,N_10711);
and U13495 (N_13495,N_9202,N_9965);
xor U13496 (N_13496,N_9840,N_10266);
and U13497 (N_13497,N_11547,N_9590);
nor U13498 (N_13498,N_9757,N_10449);
or U13499 (N_13499,N_10360,N_10154);
nor U13500 (N_13500,N_11074,N_11064);
or U13501 (N_13501,N_11756,N_10010);
xor U13502 (N_13502,N_9239,N_10767);
nor U13503 (N_13503,N_11175,N_10279);
nor U13504 (N_13504,N_9813,N_10662);
or U13505 (N_13505,N_10770,N_11861);
and U13506 (N_13506,N_10360,N_9746);
or U13507 (N_13507,N_11910,N_11803);
or U13508 (N_13508,N_10779,N_10566);
nand U13509 (N_13509,N_9089,N_11169);
or U13510 (N_13510,N_10603,N_9351);
xor U13511 (N_13511,N_11485,N_10708);
and U13512 (N_13512,N_11050,N_10557);
and U13513 (N_13513,N_11134,N_11710);
or U13514 (N_13514,N_10320,N_9073);
or U13515 (N_13515,N_11712,N_10290);
xor U13516 (N_13516,N_11914,N_10936);
nor U13517 (N_13517,N_10737,N_11515);
nor U13518 (N_13518,N_10617,N_11431);
nand U13519 (N_13519,N_10968,N_10533);
nand U13520 (N_13520,N_9860,N_11560);
nand U13521 (N_13521,N_11811,N_10664);
and U13522 (N_13522,N_11214,N_11977);
nor U13523 (N_13523,N_9875,N_10542);
or U13524 (N_13524,N_10618,N_11516);
nor U13525 (N_13525,N_11732,N_9960);
nand U13526 (N_13526,N_11516,N_11097);
nand U13527 (N_13527,N_10982,N_9615);
nand U13528 (N_13528,N_10382,N_10965);
nor U13529 (N_13529,N_9239,N_11149);
and U13530 (N_13530,N_10182,N_9703);
nand U13531 (N_13531,N_11947,N_10624);
xnor U13532 (N_13532,N_11262,N_11851);
nor U13533 (N_13533,N_9811,N_11014);
nand U13534 (N_13534,N_10960,N_10710);
nand U13535 (N_13535,N_9526,N_10138);
nand U13536 (N_13536,N_11224,N_9797);
nand U13537 (N_13537,N_9081,N_10016);
and U13538 (N_13538,N_9644,N_11494);
or U13539 (N_13539,N_9697,N_11084);
nor U13540 (N_13540,N_9541,N_9637);
and U13541 (N_13541,N_9543,N_10131);
and U13542 (N_13542,N_11598,N_10113);
nor U13543 (N_13543,N_10957,N_9858);
nand U13544 (N_13544,N_11890,N_11732);
nor U13545 (N_13545,N_9715,N_10722);
xnor U13546 (N_13546,N_10890,N_9540);
and U13547 (N_13547,N_10913,N_11070);
nand U13548 (N_13548,N_10964,N_10628);
and U13549 (N_13549,N_10631,N_10455);
nor U13550 (N_13550,N_11026,N_11515);
nand U13551 (N_13551,N_11748,N_10098);
and U13552 (N_13552,N_11226,N_9139);
and U13553 (N_13553,N_11272,N_11640);
or U13554 (N_13554,N_9726,N_10377);
and U13555 (N_13555,N_9887,N_11456);
nor U13556 (N_13556,N_10998,N_11708);
and U13557 (N_13557,N_11791,N_10738);
xor U13558 (N_13558,N_11536,N_11525);
nor U13559 (N_13559,N_9689,N_9450);
nor U13560 (N_13560,N_11119,N_11541);
and U13561 (N_13561,N_10531,N_9634);
nor U13562 (N_13562,N_9832,N_10973);
and U13563 (N_13563,N_11534,N_11321);
xnor U13564 (N_13564,N_9697,N_11012);
xnor U13565 (N_13565,N_9445,N_11764);
xnor U13566 (N_13566,N_11910,N_10285);
nor U13567 (N_13567,N_10483,N_10285);
xor U13568 (N_13568,N_9162,N_10137);
nor U13569 (N_13569,N_11947,N_9357);
xnor U13570 (N_13570,N_10542,N_10446);
or U13571 (N_13571,N_9914,N_10686);
nor U13572 (N_13572,N_11552,N_11718);
and U13573 (N_13573,N_11729,N_11045);
nand U13574 (N_13574,N_11410,N_11664);
and U13575 (N_13575,N_9162,N_9059);
and U13576 (N_13576,N_10445,N_10731);
or U13577 (N_13577,N_9475,N_9091);
xnor U13578 (N_13578,N_10657,N_11158);
nor U13579 (N_13579,N_9557,N_11472);
nand U13580 (N_13580,N_11086,N_10421);
nor U13581 (N_13581,N_9570,N_9932);
and U13582 (N_13582,N_10174,N_10789);
nand U13583 (N_13583,N_9595,N_10771);
and U13584 (N_13584,N_11152,N_9874);
nor U13585 (N_13585,N_10387,N_10019);
xnor U13586 (N_13586,N_11950,N_10700);
nand U13587 (N_13587,N_10808,N_11206);
and U13588 (N_13588,N_9678,N_10569);
nor U13589 (N_13589,N_11027,N_10559);
xor U13590 (N_13590,N_10329,N_10525);
or U13591 (N_13591,N_10251,N_10532);
and U13592 (N_13592,N_11133,N_10776);
or U13593 (N_13593,N_11108,N_11413);
and U13594 (N_13594,N_11591,N_10402);
nand U13595 (N_13595,N_9243,N_10633);
nand U13596 (N_13596,N_10011,N_9873);
and U13597 (N_13597,N_11642,N_11804);
nand U13598 (N_13598,N_11658,N_9208);
or U13599 (N_13599,N_9316,N_11170);
xor U13600 (N_13600,N_10651,N_10182);
or U13601 (N_13601,N_9222,N_11685);
and U13602 (N_13602,N_10165,N_11339);
nand U13603 (N_13603,N_9844,N_9103);
or U13604 (N_13604,N_10044,N_11547);
nand U13605 (N_13605,N_10090,N_11778);
and U13606 (N_13606,N_9735,N_11816);
or U13607 (N_13607,N_9684,N_10789);
or U13608 (N_13608,N_11645,N_9411);
nor U13609 (N_13609,N_11856,N_11525);
and U13610 (N_13610,N_9852,N_10083);
and U13611 (N_13611,N_9138,N_11296);
xnor U13612 (N_13612,N_10801,N_10426);
or U13613 (N_13613,N_10721,N_10191);
and U13614 (N_13614,N_10411,N_9039);
nor U13615 (N_13615,N_10575,N_9777);
nor U13616 (N_13616,N_9426,N_11207);
nand U13617 (N_13617,N_9458,N_9647);
and U13618 (N_13618,N_10677,N_10378);
xnor U13619 (N_13619,N_9648,N_10237);
xor U13620 (N_13620,N_10592,N_9261);
and U13621 (N_13621,N_10406,N_9726);
xnor U13622 (N_13622,N_10799,N_10628);
nand U13623 (N_13623,N_10940,N_9616);
or U13624 (N_13624,N_11660,N_10715);
nor U13625 (N_13625,N_9403,N_11995);
or U13626 (N_13626,N_9603,N_11053);
and U13627 (N_13627,N_9353,N_10326);
and U13628 (N_13628,N_10080,N_10168);
nand U13629 (N_13629,N_10825,N_9463);
nor U13630 (N_13630,N_9650,N_10430);
nor U13631 (N_13631,N_11459,N_11321);
nor U13632 (N_13632,N_9149,N_11444);
or U13633 (N_13633,N_11842,N_10167);
nand U13634 (N_13634,N_11451,N_11943);
nand U13635 (N_13635,N_10426,N_9463);
nor U13636 (N_13636,N_9981,N_10145);
and U13637 (N_13637,N_11408,N_11560);
nor U13638 (N_13638,N_9941,N_10550);
or U13639 (N_13639,N_9682,N_11702);
nor U13640 (N_13640,N_9049,N_9529);
or U13641 (N_13641,N_11330,N_9091);
nand U13642 (N_13642,N_11799,N_9531);
or U13643 (N_13643,N_9284,N_9779);
nor U13644 (N_13644,N_10649,N_11519);
or U13645 (N_13645,N_11699,N_10515);
xor U13646 (N_13646,N_11633,N_10209);
nor U13647 (N_13647,N_9442,N_9351);
and U13648 (N_13648,N_9192,N_9890);
nor U13649 (N_13649,N_11525,N_10621);
and U13650 (N_13650,N_9352,N_9274);
and U13651 (N_13651,N_9722,N_9784);
and U13652 (N_13652,N_9934,N_9089);
and U13653 (N_13653,N_10228,N_11092);
xor U13654 (N_13654,N_10094,N_10462);
and U13655 (N_13655,N_11719,N_10926);
nor U13656 (N_13656,N_11515,N_10912);
or U13657 (N_13657,N_11706,N_10262);
nand U13658 (N_13658,N_10624,N_10519);
xnor U13659 (N_13659,N_10317,N_10855);
and U13660 (N_13660,N_9368,N_9164);
xor U13661 (N_13661,N_11039,N_11726);
and U13662 (N_13662,N_9396,N_11448);
xor U13663 (N_13663,N_10014,N_9272);
or U13664 (N_13664,N_10743,N_11688);
or U13665 (N_13665,N_11765,N_11130);
xnor U13666 (N_13666,N_11551,N_9777);
and U13667 (N_13667,N_10086,N_11057);
and U13668 (N_13668,N_11003,N_10124);
or U13669 (N_13669,N_9608,N_9059);
nand U13670 (N_13670,N_9811,N_11556);
and U13671 (N_13671,N_9220,N_11501);
or U13672 (N_13672,N_11399,N_10699);
nand U13673 (N_13673,N_9157,N_11296);
xor U13674 (N_13674,N_10305,N_10315);
xnor U13675 (N_13675,N_10206,N_11566);
xnor U13676 (N_13676,N_9507,N_11900);
nor U13677 (N_13677,N_10874,N_9442);
and U13678 (N_13678,N_9985,N_11242);
xnor U13679 (N_13679,N_10636,N_9560);
or U13680 (N_13680,N_11900,N_10132);
xnor U13681 (N_13681,N_9299,N_10370);
xnor U13682 (N_13682,N_10891,N_11715);
and U13683 (N_13683,N_9628,N_11294);
and U13684 (N_13684,N_10997,N_9318);
nand U13685 (N_13685,N_9916,N_9898);
or U13686 (N_13686,N_11597,N_10395);
nand U13687 (N_13687,N_11879,N_10991);
nand U13688 (N_13688,N_9024,N_10646);
and U13689 (N_13689,N_11666,N_11430);
nor U13690 (N_13690,N_11000,N_11819);
or U13691 (N_13691,N_10603,N_10980);
nor U13692 (N_13692,N_9546,N_11704);
and U13693 (N_13693,N_11658,N_9867);
xnor U13694 (N_13694,N_11887,N_11505);
nor U13695 (N_13695,N_11959,N_9441);
nor U13696 (N_13696,N_11948,N_9537);
xnor U13697 (N_13697,N_10090,N_10372);
xor U13698 (N_13698,N_11615,N_11301);
nand U13699 (N_13699,N_11210,N_11707);
and U13700 (N_13700,N_11445,N_10121);
and U13701 (N_13701,N_9877,N_9284);
nor U13702 (N_13702,N_11453,N_10074);
and U13703 (N_13703,N_11067,N_10922);
nand U13704 (N_13704,N_10401,N_11054);
xnor U13705 (N_13705,N_10580,N_11216);
nand U13706 (N_13706,N_9058,N_11781);
nand U13707 (N_13707,N_9557,N_9847);
nor U13708 (N_13708,N_10356,N_11765);
nand U13709 (N_13709,N_11204,N_9132);
xnor U13710 (N_13710,N_9880,N_11173);
or U13711 (N_13711,N_9307,N_11439);
or U13712 (N_13712,N_11366,N_10608);
or U13713 (N_13713,N_9114,N_11604);
or U13714 (N_13714,N_11626,N_9578);
nor U13715 (N_13715,N_10585,N_10810);
xor U13716 (N_13716,N_10129,N_11299);
or U13717 (N_13717,N_9265,N_10371);
xor U13718 (N_13718,N_11638,N_9313);
xnor U13719 (N_13719,N_11450,N_9096);
or U13720 (N_13720,N_11602,N_11271);
nor U13721 (N_13721,N_11739,N_9971);
or U13722 (N_13722,N_9703,N_10758);
xnor U13723 (N_13723,N_10996,N_9369);
xor U13724 (N_13724,N_9652,N_9745);
nand U13725 (N_13725,N_10805,N_9476);
xnor U13726 (N_13726,N_10511,N_9230);
nor U13727 (N_13727,N_10164,N_10058);
or U13728 (N_13728,N_9219,N_10002);
or U13729 (N_13729,N_10739,N_11546);
xor U13730 (N_13730,N_9336,N_9687);
or U13731 (N_13731,N_11964,N_11360);
and U13732 (N_13732,N_9827,N_9009);
xnor U13733 (N_13733,N_11774,N_11725);
xor U13734 (N_13734,N_10997,N_11285);
nor U13735 (N_13735,N_10468,N_10969);
and U13736 (N_13736,N_9413,N_9730);
and U13737 (N_13737,N_11858,N_10402);
or U13738 (N_13738,N_9995,N_11337);
nand U13739 (N_13739,N_9554,N_10284);
or U13740 (N_13740,N_9812,N_9135);
xnor U13741 (N_13741,N_11985,N_10118);
xor U13742 (N_13742,N_9064,N_9093);
or U13743 (N_13743,N_10722,N_11325);
xnor U13744 (N_13744,N_10621,N_9149);
xor U13745 (N_13745,N_9014,N_11614);
nand U13746 (N_13746,N_9595,N_9437);
nor U13747 (N_13747,N_9980,N_9049);
nor U13748 (N_13748,N_10856,N_10711);
and U13749 (N_13749,N_11437,N_9123);
and U13750 (N_13750,N_11762,N_9958);
xnor U13751 (N_13751,N_9817,N_10082);
or U13752 (N_13752,N_9696,N_11190);
nand U13753 (N_13753,N_10443,N_9157);
or U13754 (N_13754,N_9247,N_9282);
and U13755 (N_13755,N_9145,N_10395);
nand U13756 (N_13756,N_10309,N_9643);
nor U13757 (N_13757,N_11079,N_9895);
or U13758 (N_13758,N_9606,N_10094);
or U13759 (N_13759,N_11897,N_10164);
nor U13760 (N_13760,N_10035,N_9676);
nor U13761 (N_13761,N_11254,N_11189);
nor U13762 (N_13762,N_11882,N_10568);
nand U13763 (N_13763,N_9463,N_10654);
or U13764 (N_13764,N_9699,N_11944);
and U13765 (N_13765,N_9786,N_10885);
nor U13766 (N_13766,N_11083,N_10549);
nor U13767 (N_13767,N_9518,N_11561);
or U13768 (N_13768,N_10212,N_9880);
and U13769 (N_13769,N_9942,N_9303);
xnor U13770 (N_13770,N_9923,N_11457);
or U13771 (N_13771,N_10399,N_9625);
nor U13772 (N_13772,N_11857,N_11532);
xor U13773 (N_13773,N_9809,N_11060);
nand U13774 (N_13774,N_9616,N_9309);
nor U13775 (N_13775,N_9185,N_10998);
or U13776 (N_13776,N_9086,N_9710);
or U13777 (N_13777,N_9313,N_11075);
or U13778 (N_13778,N_9649,N_9786);
and U13779 (N_13779,N_9464,N_11351);
and U13780 (N_13780,N_10770,N_11149);
nand U13781 (N_13781,N_9512,N_10639);
nor U13782 (N_13782,N_9899,N_11015);
and U13783 (N_13783,N_11408,N_11378);
xnor U13784 (N_13784,N_9851,N_10812);
or U13785 (N_13785,N_9900,N_11259);
xnor U13786 (N_13786,N_9721,N_10146);
or U13787 (N_13787,N_11245,N_11132);
or U13788 (N_13788,N_10080,N_10980);
xor U13789 (N_13789,N_11059,N_9388);
and U13790 (N_13790,N_10652,N_10459);
xnor U13791 (N_13791,N_9350,N_11727);
nor U13792 (N_13792,N_11288,N_10227);
or U13793 (N_13793,N_11378,N_10055);
and U13794 (N_13794,N_10566,N_11243);
or U13795 (N_13795,N_10388,N_11676);
or U13796 (N_13796,N_9016,N_11843);
and U13797 (N_13797,N_9023,N_9205);
nor U13798 (N_13798,N_9161,N_9721);
or U13799 (N_13799,N_11950,N_11021);
and U13800 (N_13800,N_10061,N_10694);
xor U13801 (N_13801,N_9720,N_10241);
and U13802 (N_13802,N_9058,N_11954);
nor U13803 (N_13803,N_9757,N_9941);
xor U13804 (N_13804,N_11202,N_10195);
nand U13805 (N_13805,N_10768,N_9560);
nor U13806 (N_13806,N_11599,N_9904);
xor U13807 (N_13807,N_9208,N_10686);
or U13808 (N_13808,N_10905,N_10779);
nand U13809 (N_13809,N_10625,N_9270);
nor U13810 (N_13810,N_10114,N_10348);
and U13811 (N_13811,N_11645,N_10918);
and U13812 (N_13812,N_10927,N_11812);
xor U13813 (N_13813,N_11530,N_10348);
nand U13814 (N_13814,N_11351,N_10830);
or U13815 (N_13815,N_10314,N_9535);
or U13816 (N_13816,N_10637,N_9598);
and U13817 (N_13817,N_10891,N_11890);
and U13818 (N_13818,N_10514,N_10452);
nand U13819 (N_13819,N_10657,N_9453);
nor U13820 (N_13820,N_9729,N_9602);
xor U13821 (N_13821,N_9832,N_10283);
nor U13822 (N_13822,N_11275,N_10636);
nand U13823 (N_13823,N_10447,N_10605);
nor U13824 (N_13824,N_10094,N_9944);
nand U13825 (N_13825,N_9619,N_9632);
nor U13826 (N_13826,N_11050,N_9899);
nand U13827 (N_13827,N_11771,N_11355);
xnor U13828 (N_13828,N_11269,N_11154);
nor U13829 (N_13829,N_10503,N_11047);
or U13830 (N_13830,N_9166,N_9064);
nand U13831 (N_13831,N_9412,N_10188);
and U13832 (N_13832,N_10108,N_11535);
xnor U13833 (N_13833,N_10247,N_11343);
and U13834 (N_13834,N_11741,N_11497);
nand U13835 (N_13835,N_10702,N_10325);
and U13836 (N_13836,N_10622,N_11625);
xor U13837 (N_13837,N_10434,N_11587);
and U13838 (N_13838,N_11273,N_10493);
nor U13839 (N_13839,N_10530,N_10049);
nand U13840 (N_13840,N_11684,N_9369);
and U13841 (N_13841,N_11280,N_9342);
xnor U13842 (N_13842,N_9097,N_9325);
nand U13843 (N_13843,N_9500,N_9895);
xor U13844 (N_13844,N_11333,N_10065);
nand U13845 (N_13845,N_9134,N_10341);
xor U13846 (N_13846,N_10289,N_11802);
and U13847 (N_13847,N_9100,N_9299);
nand U13848 (N_13848,N_10804,N_10080);
xnor U13849 (N_13849,N_11914,N_10012);
nand U13850 (N_13850,N_10969,N_9809);
nand U13851 (N_13851,N_10540,N_10760);
and U13852 (N_13852,N_10509,N_11711);
or U13853 (N_13853,N_10790,N_9934);
xnor U13854 (N_13854,N_9085,N_11138);
and U13855 (N_13855,N_10577,N_9152);
and U13856 (N_13856,N_11675,N_11045);
or U13857 (N_13857,N_11605,N_11519);
nand U13858 (N_13858,N_10936,N_11075);
nor U13859 (N_13859,N_11873,N_11350);
and U13860 (N_13860,N_11838,N_9156);
nor U13861 (N_13861,N_10749,N_11590);
or U13862 (N_13862,N_9729,N_11218);
or U13863 (N_13863,N_9078,N_10448);
nor U13864 (N_13864,N_9940,N_9825);
and U13865 (N_13865,N_9406,N_11565);
nand U13866 (N_13866,N_11964,N_11526);
xnor U13867 (N_13867,N_9592,N_11536);
and U13868 (N_13868,N_10189,N_11720);
or U13869 (N_13869,N_9623,N_9124);
and U13870 (N_13870,N_10395,N_9777);
nand U13871 (N_13871,N_10211,N_11216);
nor U13872 (N_13872,N_9239,N_11078);
or U13873 (N_13873,N_11011,N_10804);
or U13874 (N_13874,N_10310,N_9151);
nor U13875 (N_13875,N_9721,N_11455);
nor U13876 (N_13876,N_9367,N_9425);
or U13877 (N_13877,N_11029,N_9303);
nand U13878 (N_13878,N_10111,N_10998);
xnor U13879 (N_13879,N_9651,N_9199);
xnor U13880 (N_13880,N_11705,N_11413);
nand U13881 (N_13881,N_9385,N_11885);
or U13882 (N_13882,N_11361,N_10045);
and U13883 (N_13883,N_9779,N_9453);
nor U13884 (N_13884,N_10759,N_9877);
xor U13885 (N_13885,N_9808,N_11811);
nand U13886 (N_13886,N_9127,N_10453);
xnor U13887 (N_13887,N_9049,N_9892);
or U13888 (N_13888,N_10729,N_11898);
nor U13889 (N_13889,N_9326,N_9493);
and U13890 (N_13890,N_9184,N_11211);
or U13891 (N_13891,N_10855,N_11155);
and U13892 (N_13892,N_10653,N_11431);
xor U13893 (N_13893,N_10127,N_11187);
and U13894 (N_13894,N_10877,N_10139);
xor U13895 (N_13895,N_9988,N_10657);
nand U13896 (N_13896,N_10643,N_9904);
nand U13897 (N_13897,N_11292,N_9884);
xnor U13898 (N_13898,N_11572,N_9934);
nand U13899 (N_13899,N_10086,N_11503);
or U13900 (N_13900,N_10242,N_10416);
xor U13901 (N_13901,N_10843,N_9638);
xor U13902 (N_13902,N_9242,N_9595);
nand U13903 (N_13903,N_9381,N_9840);
nand U13904 (N_13904,N_10754,N_10379);
and U13905 (N_13905,N_11964,N_9695);
or U13906 (N_13906,N_10670,N_11998);
nor U13907 (N_13907,N_10164,N_10439);
nand U13908 (N_13908,N_9710,N_9333);
and U13909 (N_13909,N_9858,N_10642);
and U13910 (N_13910,N_9603,N_11754);
xnor U13911 (N_13911,N_11179,N_10094);
xor U13912 (N_13912,N_10030,N_10063);
and U13913 (N_13913,N_11909,N_9133);
nand U13914 (N_13914,N_10685,N_9708);
xnor U13915 (N_13915,N_9666,N_11355);
nand U13916 (N_13916,N_11695,N_9932);
nor U13917 (N_13917,N_9049,N_10449);
or U13918 (N_13918,N_10294,N_11515);
and U13919 (N_13919,N_9896,N_9041);
xor U13920 (N_13920,N_9373,N_10054);
xor U13921 (N_13921,N_10853,N_11312);
xnor U13922 (N_13922,N_11467,N_11936);
or U13923 (N_13923,N_9647,N_10646);
xnor U13924 (N_13924,N_11950,N_10734);
xor U13925 (N_13925,N_9078,N_10161);
nor U13926 (N_13926,N_10665,N_11996);
nand U13927 (N_13927,N_11401,N_9040);
xor U13928 (N_13928,N_9408,N_9922);
and U13929 (N_13929,N_10214,N_9707);
and U13930 (N_13930,N_11855,N_10772);
xnor U13931 (N_13931,N_9268,N_9093);
or U13932 (N_13932,N_11162,N_9839);
nand U13933 (N_13933,N_9685,N_11702);
or U13934 (N_13934,N_10421,N_10121);
xnor U13935 (N_13935,N_11786,N_10381);
nand U13936 (N_13936,N_9019,N_9755);
xnor U13937 (N_13937,N_10009,N_10203);
nor U13938 (N_13938,N_9548,N_11013);
or U13939 (N_13939,N_10743,N_11143);
and U13940 (N_13940,N_11483,N_10719);
and U13941 (N_13941,N_9865,N_9870);
and U13942 (N_13942,N_11690,N_9010);
or U13943 (N_13943,N_10227,N_11058);
nor U13944 (N_13944,N_11941,N_9531);
nand U13945 (N_13945,N_9055,N_9635);
nor U13946 (N_13946,N_10763,N_11344);
or U13947 (N_13947,N_10616,N_11868);
or U13948 (N_13948,N_11104,N_9996);
xnor U13949 (N_13949,N_10605,N_10190);
nand U13950 (N_13950,N_11241,N_10970);
or U13951 (N_13951,N_9817,N_11067);
xor U13952 (N_13952,N_11075,N_9299);
or U13953 (N_13953,N_10246,N_10337);
or U13954 (N_13954,N_9897,N_11469);
xor U13955 (N_13955,N_11772,N_10384);
nor U13956 (N_13956,N_9764,N_10624);
nand U13957 (N_13957,N_10355,N_10779);
and U13958 (N_13958,N_9489,N_9554);
nand U13959 (N_13959,N_11613,N_11923);
xnor U13960 (N_13960,N_11288,N_9197);
xor U13961 (N_13961,N_9964,N_10770);
xnor U13962 (N_13962,N_10048,N_10472);
xor U13963 (N_13963,N_10562,N_11470);
nand U13964 (N_13964,N_11187,N_11181);
and U13965 (N_13965,N_9098,N_10795);
and U13966 (N_13966,N_9693,N_9786);
nor U13967 (N_13967,N_11096,N_9583);
or U13968 (N_13968,N_10433,N_9896);
xor U13969 (N_13969,N_10554,N_11592);
and U13970 (N_13970,N_10717,N_11155);
xor U13971 (N_13971,N_9040,N_10887);
xnor U13972 (N_13972,N_10665,N_11220);
nor U13973 (N_13973,N_11132,N_11571);
nand U13974 (N_13974,N_10661,N_10246);
and U13975 (N_13975,N_10008,N_11401);
nor U13976 (N_13976,N_11579,N_10839);
nand U13977 (N_13977,N_9421,N_11003);
nand U13978 (N_13978,N_11202,N_11653);
or U13979 (N_13979,N_10981,N_10893);
and U13980 (N_13980,N_9161,N_10674);
or U13981 (N_13981,N_11140,N_11448);
and U13982 (N_13982,N_11000,N_9978);
and U13983 (N_13983,N_11610,N_10394);
and U13984 (N_13984,N_11422,N_10894);
xor U13985 (N_13985,N_11574,N_9968);
and U13986 (N_13986,N_11947,N_10850);
or U13987 (N_13987,N_9517,N_10037);
nand U13988 (N_13988,N_10081,N_11463);
or U13989 (N_13989,N_10218,N_10550);
or U13990 (N_13990,N_10631,N_9634);
and U13991 (N_13991,N_11311,N_9409);
nand U13992 (N_13992,N_11005,N_10231);
and U13993 (N_13993,N_10518,N_9931);
and U13994 (N_13994,N_11577,N_11609);
nor U13995 (N_13995,N_11110,N_9955);
or U13996 (N_13996,N_11760,N_10863);
nor U13997 (N_13997,N_10768,N_9652);
or U13998 (N_13998,N_10388,N_9105);
or U13999 (N_13999,N_9632,N_11264);
and U14000 (N_14000,N_11421,N_11260);
or U14001 (N_14001,N_11917,N_11695);
xor U14002 (N_14002,N_10651,N_11759);
and U14003 (N_14003,N_10994,N_11786);
nand U14004 (N_14004,N_9250,N_10840);
or U14005 (N_14005,N_9278,N_9464);
nand U14006 (N_14006,N_9001,N_11409);
or U14007 (N_14007,N_11067,N_11151);
xor U14008 (N_14008,N_9429,N_11025);
xor U14009 (N_14009,N_10850,N_9724);
nor U14010 (N_14010,N_11555,N_11995);
nor U14011 (N_14011,N_10541,N_10223);
and U14012 (N_14012,N_10855,N_9514);
xor U14013 (N_14013,N_11933,N_10120);
xnor U14014 (N_14014,N_10839,N_10002);
nand U14015 (N_14015,N_11668,N_11399);
or U14016 (N_14016,N_11598,N_10520);
nand U14017 (N_14017,N_9011,N_9876);
xor U14018 (N_14018,N_11920,N_9981);
nor U14019 (N_14019,N_9437,N_11599);
nor U14020 (N_14020,N_11013,N_10099);
xor U14021 (N_14021,N_11420,N_10972);
nor U14022 (N_14022,N_9353,N_9052);
xnor U14023 (N_14023,N_11775,N_9927);
nand U14024 (N_14024,N_11327,N_10806);
and U14025 (N_14025,N_9615,N_9304);
or U14026 (N_14026,N_11688,N_11443);
and U14027 (N_14027,N_10243,N_11079);
and U14028 (N_14028,N_9993,N_10960);
nand U14029 (N_14029,N_9982,N_9724);
or U14030 (N_14030,N_9509,N_11717);
xor U14031 (N_14031,N_10240,N_9487);
xor U14032 (N_14032,N_10055,N_9875);
and U14033 (N_14033,N_9982,N_11499);
nand U14034 (N_14034,N_10610,N_11607);
nor U14035 (N_14035,N_9666,N_10463);
xor U14036 (N_14036,N_10513,N_10475);
or U14037 (N_14037,N_10735,N_11871);
nor U14038 (N_14038,N_9032,N_11953);
nor U14039 (N_14039,N_9773,N_10375);
and U14040 (N_14040,N_9014,N_9356);
and U14041 (N_14041,N_11900,N_9323);
xor U14042 (N_14042,N_11037,N_10954);
and U14043 (N_14043,N_9491,N_11954);
or U14044 (N_14044,N_9179,N_11951);
nand U14045 (N_14045,N_9207,N_11912);
or U14046 (N_14046,N_10369,N_10026);
nand U14047 (N_14047,N_11806,N_11661);
nor U14048 (N_14048,N_9273,N_9604);
nand U14049 (N_14049,N_11219,N_10761);
or U14050 (N_14050,N_9560,N_9420);
nor U14051 (N_14051,N_10754,N_9107);
and U14052 (N_14052,N_10296,N_10601);
xor U14053 (N_14053,N_11106,N_10363);
nor U14054 (N_14054,N_10259,N_9650);
or U14055 (N_14055,N_11585,N_10827);
or U14056 (N_14056,N_9282,N_10473);
nor U14057 (N_14057,N_10205,N_11524);
nand U14058 (N_14058,N_11437,N_10685);
or U14059 (N_14059,N_11695,N_10710);
and U14060 (N_14060,N_11141,N_9115);
nand U14061 (N_14061,N_10891,N_10527);
xor U14062 (N_14062,N_9815,N_9760);
xor U14063 (N_14063,N_9116,N_9390);
and U14064 (N_14064,N_11451,N_9253);
xor U14065 (N_14065,N_10017,N_9371);
xor U14066 (N_14066,N_9883,N_10740);
nand U14067 (N_14067,N_11386,N_10133);
or U14068 (N_14068,N_11909,N_9386);
and U14069 (N_14069,N_9518,N_10399);
nand U14070 (N_14070,N_10311,N_10560);
or U14071 (N_14071,N_11381,N_10701);
nor U14072 (N_14072,N_9499,N_9768);
or U14073 (N_14073,N_10262,N_11977);
or U14074 (N_14074,N_10412,N_11340);
xor U14075 (N_14075,N_10579,N_11805);
or U14076 (N_14076,N_10021,N_11092);
nor U14077 (N_14077,N_9639,N_11262);
or U14078 (N_14078,N_10913,N_9967);
or U14079 (N_14079,N_11550,N_11716);
xnor U14080 (N_14080,N_9922,N_11461);
and U14081 (N_14081,N_10621,N_9895);
nor U14082 (N_14082,N_10754,N_10012);
and U14083 (N_14083,N_9969,N_11008);
or U14084 (N_14084,N_9030,N_10669);
xor U14085 (N_14085,N_11876,N_10553);
and U14086 (N_14086,N_11930,N_10834);
xor U14087 (N_14087,N_9969,N_10850);
xnor U14088 (N_14088,N_11979,N_9428);
xor U14089 (N_14089,N_9021,N_9093);
nand U14090 (N_14090,N_10641,N_10636);
nand U14091 (N_14091,N_9826,N_11347);
xor U14092 (N_14092,N_10802,N_9914);
nand U14093 (N_14093,N_10066,N_10627);
xor U14094 (N_14094,N_11983,N_11666);
xnor U14095 (N_14095,N_9284,N_11263);
and U14096 (N_14096,N_10623,N_10523);
nand U14097 (N_14097,N_11857,N_10158);
and U14098 (N_14098,N_11209,N_11599);
or U14099 (N_14099,N_11444,N_10502);
nor U14100 (N_14100,N_11276,N_9606);
nand U14101 (N_14101,N_11286,N_10700);
nand U14102 (N_14102,N_9873,N_11693);
nand U14103 (N_14103,N_9381,N_10493);
xnor U14104 (N_14104,N_10241,N_9522);
xor U14105 (N_14105,N_11469,N_10382);
nand U14106 (N_14106,N_10957,N_10087);
xor U14107 (N_14107,N_10846,N_10397);
xnor U14108 (N_14108,N_11716,N_9573);
and U14109 (N_14109,N_11292,N_10437);
nor U14110 (N_14110,N_10936,N_9320);
nor U14111 (N_14111,N_9322,N_10554);
nand U14112 (N_14112,N_10163,N_9461);
or U14113 (N_14113,N_10704,N_9040);
xnor U14114 (N_14114,N_11622,N_10117);
xnor U14115 (N_14115,N_9351,N_11343);
xnor U14116 (N_14116,N_11678,N_11727);
xnor U14117 (N_14117,N_11275,N_9577);
nor U14118 (N_14118,N_11290,N_10281);
nand U14119 (N_14119,N_10620,N_9345);
and U14120 (N_14120,N_9821,N_10744);
nor U14121 (N_14121,N_10029,N_10529);
and U14122 (N_14122,N_9286,N_11229);
xnor U14123 (N_14123,N_9044,N_10243);
and U14124 (N_14124,N_9942,N_10019);
nand U14125 (N_14125,N_11155,N_10291);
xor U14126 (N_14126,N_11395,N_11547);
xnor U14127 (N_14127,N_10737,N_11778);
nor U14128 (N_14128,N_11107,N_10056);
nor U14129 (N_14129,N_10291,N_11410);
nor U14130 (N_14130,N_11001,N_10272);
or U14131 (N_14131,N_9474,N_9863);
nor U14132 (N_14132,N_11590,N_9059);
xor U14133 (N_14133,N_9768,N_9806);
xor U14134 (N_14134,N_9485,N_10854);
and U14135 (N_14135,N_11059,N_11108);
and U14136 (N_14136,N_9337,N_11393);
nor U14137 (N_14137,N_10214,N_11507);
nor U14138 (N_14138,N_10017,N_9055);
and U14139 (N_14139,N_10133,N_9254);
xor U14140 (N_14140,N_9391,N_11813);
nand U14141 (N_14141,N_9479,N_9182);
and U14142 (N_14142,N_10339,N_9964);
nand U14143 (N_14143,N_9584,N_11006);
xnor U14144 (N_14144,N_11314,N_10449);
nor U14145 (N_14145,N_9069,N_10986);
or U14146 (N_14146,N_10255,N_10392);
or U14147 (N_14147,N_11189,N_9418);
or U14148 (N_14148,N_10066,N_10769);
xor U14149 (N_14149,N_9568,N_10280);
nand U14150 (N_14150,N_11342,N_10565);
nand U14151 (N_14151,N_10181,N_11959);
nand U14152 (N_14152,N_11186,N_9455);
or U14153 (N_14153,N_11459,N_11728);
nor U14154 (N_14154,N_11349,N_11718);
nand U14155 (N_14155,N_9932,N_9961);
or U14156 (N_14156,N_11038,N_11451);
or U14157 (N_14157,N_11235,N_11840);
nor U14158 (N_14158,N_9202,N_10619);
and U14159 (N_14159,N_10340,N_11041);
or U14160 (N_14160,N_9216,N_11466);
xor U14161 (N_14161,N_11922,N_10459);
nand U14162 (N_14162,N_9237,N_11168);
or U14163 (N_14163,N_9162,N_11167);
xnor U14164 (N_14164,N_11922,N_9068);
nor U14165 (N_14165,N_11245,N_9354);
or U14166 (N_14166,N_9940,N_11359);
and U14167 (N_14167,N_10882,N_9968);
or U14168 (N_14168,N_9681,N_9490);
and U14169 (N_14169,N_9455,N_10900);
or U14170 (N_14170,N_11178,N_9267);
xnor U14171 (N_14171,N_9772,N_11036);
and U14172 (N_14172,N_11172,N_9450);
nor U14173 (N_14173,N_10282,N_9978);
nor U14174 (N_14174,N_10547,N_9066);
or U14175 (N_14175,N_9451,N_11532);
nor U14176 (N_14176,N_10042,N_9044);
or U14177 (N_14177,N_10313,N_11007);
and U14178 (N_14178,N_9613,N_11123);
nor U14179 (N_14179,N_11354,N_9131);
or U14180 (N_14180,N_10539,N_9625);
or U14181 (N_14181,N_10456,N_10410);
nor U14182 (N_14182,N_11495,N_9821);
or U14183 (N_14183,N_9810,N_10233);
and U14184 (N_14184,N_11761,N_10428);
nand U14185 (N_14185,N_11022,N_10119);
nand U14186 (N_14186,N_10906,N_11677);
xnor U14187 (N_14187,N_10734,N_9390);
and U14188 (N_14188,N_10672,N_10906);
nor U14189 (N_14189,N_9796,N_9454);
nand U14190 (N_14190,N_9049,N_10640);
or U14191 (N_14191,N_9851,N_10848);
or U14192 (N_14192,N_9249,N_10295);
nor U14193 (N_14193,N_10654,N_10197);
or U14194 (N_14194,N_11772,N_9851);
and U14195 (N_14195,N_9265,N_10303);
and U14196 (N_14196,N_10314,N_11504);
or U14197 (N_14197,N_11821,N_10112);
xnor U14198 (N_14198,N_9494,N_9777);
nor U14199 (N_14199,N_11552,N_9981);
and U14200 (N_14200,N_11051,N_11072);
nand U14201 (N_14201,N_11075,N_9698);
or U14202 (N_14202,N_11773,N_9790);
nor U14203 (N_14203,N_10733,N_11776);
nor U14204 (N_14204,N_9407,N_9982);
and U14205 (N_14205,N_10143,N_11094);
or U14206 (N_14206,N_10950,N_11890);
xor U14207 (N_14207,N_11054,N_10046);
nand U14208 (N_14208,N_11584,N_11517);
nor U14209 (N_14209,N_11067,N_11213);
nand U14210 (N_14210,N_9847,N_11224);
xor U14211 (N_14211,N_9149,N_11182);
xnor U14212 (N_14212,N_9080,N_10800);
nand U14213 (N_14213,N_9129,N_9495);
nor U14214 (N_14214,N_9078,N_10683);
xnor U14215 (N_14215,N_10699,N_10863);
and U14216 (N_14216,N_10257,N_9698);
nor U14217 (N_14217,N_10583,N_9910);
nor U14218 (N_14218,N_11578,N_9294);
xnor U14219 (N_14219,N_9298,N_10031);
nand U14220 (N_14220,N_9451,N_9168);
nor U14221 (N_14221,N_9238,N_10029);
nand U14222 (N_14222,N_9379,N_9606);
nor U14223 (N_14223,N_9139,N_11054);
and U14224 (N_14224,N_9926,N_10385);
nand U14225 (N_14225,N_9316,N_9169);
and U14226 (N_14226,N_9758,N_11600);
or U14227 (N_14227,N_10237,N_9389);
or U14228 (N_14228,N_9410,N_11853);
xnor U14229 (N_14229,N_9076,N_10763);
nor U14230 (N_14230,N_10111,N_10304);
nand U14231 (N_14231,N_11975,N_10828);
nor U14232 (N_14232,N_10028,N_10948);
xnor U14233 (N_14233,N_11326,N_10355);
nor U14234 (N_14234,N_11102,N_10826);
nand U14235 (N_14235,N_11538,N_9671);
nor U14236 (N_14236,N_9885,N_10212);
and U14237 (N_14237,N_11782,N_10399);
xor U14238 (N_14238,N_9041,N_10839);
and U14239 (N_14239,N_10539,N_11651);
nor U14240 (N_14240,N_10521,N_9476);
and U14241 (N_14241,N_11680,N_9716);
or U14242 (N_14242,N_9167,N_9753);
nand U14243 (N_14243,N_9159,N_10352);
nand U14244 (N_14244,N_9503,N_10127);
and U14245 (N_14245,N_10328,N_11739);
xnor U14246 (N_14246,N_9953,N_11612);
and U14247 (N_14247,N_11672,N_11908);
nor U14248 (N_14248,N_10090,N_9646);
and U14249 (N_14249,N_10291,N_11863);
xnor U14250 (N_14250,N_11793,N_11362);
xor U14251 (N_14251,N_10044,N_11643);
xor U14252 (N_14252,N_11279,N_9954);
or U14253 (N_14253,N_9784,N_11698);
nor U14254 (N_14254,N_11702,N_9634);
nand U14255 (N_14255,N_11427,N_11738);
nor U14256 (N_14256,N_9052,N_10657);
xor U14257 (N_14257,N_10911,N_9487);
or U14258 (N_14258,N_10110,N_10494);
and U14259 (N_14259,N_11534,N_10923);
nor U14260 (N_14260,N_9170,N_10367);
nor U14261 (N_14261,N_9856,N_10482);
nand U14262 (N_14262,N_10865,N_9466);
or U14263 (N_14263,N_9820,N_11720);
xor U14264 (N_14264,N_10239,N_11691);
xor U14265 (N_14265,N_10873,N_9466);
or U14266 (N_14266,N_10870,N_9541);
xor U14267 (N_14267,N_9455,N_11682);
and U14268 (N_14268,N_11066,N_10965);
nor U14269 (N_14269,N_10190,N_11902);
or U14270 (N_14270,N_10207,N_11264);
and U14271 (N_14271,N_11082,N_10490);
nor U14272 (N_14272,N_10644,N_11914);
or U14273 (N_14273,N_9698,N_11895);
xnor U14274 (N_14274,N_10265,N_9460);
nand U14275 (N_14275,N_11922,N_9081);
nor U14276 (N_14276,N_9277,N_10115);
nand U14277 (N_14277,N_9137,N_10973);
and U14278 (N_14278,N_9051,N_10375);
xor U14279 (N_14279,N_11421,N_10447);
xor U14280 (N_14280,N_11814,N_11073);
and U14281 (N_14281,N_11453,N_9014);
or U14282 (N_14282,N_10317,N_9295);
or U14283 (N_14283,N_9982,N_9123);
nor U14284 (N_14284,N_11685,N_11176);
nor U14285 (N_14285,N_11382,N_11225);
and U14286 (N_14286,N_11892,N_9414);
and U14287 (N_14287,N_9128,N_9225);
nand U14288 (N_14288,N_9166,N_10579);
nor U14289 (N_14289,N_10986,N_10703);
and U14290 (N_14290,N_10764,N_11959);
nor U14291 (N_14291,N_11506,N_11588);
xor U14292 (N_14292,N_11763,N_10200);
or U14293 (N_14293,N_10368,N_9681);
and U14294 (N_14294,N_9803,N_9237);
xnor U14295 (N_14295,N_10588,N_11570);
or U14296 (N_14296,N_9084,N_11212);
xnor U14297 (N_14297,N_9581,N_11558);
xnor U14298 (N_14298,N_9408,N_9229);
nor U14299 (N_14299,N_9582,N_10506);
xnor U14300 (N_14300,N_11322,N_9565);
nand U14301 (N_14301,N_9646,N_9330);
xnor U14302 (N_14302,N_11599,N_9610);
and U14303 (N_14303,N_10955,N_9386);
nor U14304 (N_14304,N_9619,N_10281);
xor U14305 (N_14305,N_10258,N_10254);
and U14306 (N_14306,N_9873,N_11115);
nor U14307 (N_14307,N_11248,N_11997);
and U14308 (N_14308,N_9929,N_10288);
or U14309 (N_14309,N_9153,N_11955);
nand U14310 (N_14310,N_9206,N_11695);
nor U14311 (N_14311,N_10913,N_10948);
or U14312 (N_14312,N_10136,N_9689);
or U14313 (N_14313,N_11699,N_11860);
xor U14314 (N_14314,N_10090,N_10297);
or U14315 (N_14315,N_9254,N_9991);
nand U14316 (N_14316,N_10344,N_11847);
xnor U14317 (N_14317,N_9028,N_10785);
nor U14318 (N_14318,N_9160,N_10460);
xnor U14319 (N_14319,N_11161,N_11681);
xnor U14320 (N_14320,N_11071,N_11349);
nand U14321 (N_14321,N_11669,N_9993);
xnor U14322 (N_14322,N_11744,N_9410);
xor U14323 (N_14323,N_9219,N_9404);
xor U14324 (N_14324,N_11044,N_11742);
xnor U14325 (N_14325,N_11815,N_10925);
nand U14326 (N_14326,N_10702,N_11369);
nor U14327 (N_14327,N_11068,N_10943);
nand U14328 (N_14328,N_11619,N_9630);
nor U14329 (N_14329,N_10687,N_10317);
and U14330 (N_14330,N_9709,N_10114);
nor U14331 (N_14331,N_9725,N_9666);
xnor U14332 (N_14332,N_10622,N_10093);
nand U14333 (N_14333,N_9240,N_9648);
xnor U14334 (N_14334,N_11318,N_9564);
nand U14335 (N_14335,N_9337,N_9302);
nor U14336 (N_14336,N_11375,N_10247);
xor U14337 (N_14337,N_10504,N_10487);
nand U14338 (N_14338,N_10994,N_10950);
nand U14339 (N_14339,N_9170,N_11940);
nand U14340 (N_14340,N_11029,N_9299);
xnor U14341 (N_14341,N_9336,N_10999);
xor U14342 (N_14342,N_11734,N_10401);
or U14343 (N_14343,N_9600,N_10455);
nand U14344 (N_14344,N_9749,N_9318);
and U14345 (N_14345,N_9126,N_9704);
nor U14346 (N_14346,N_10696,N_9998);
nand U14347 (N_14347,N_11271,N_9191);
and U14348 (N_14348,N_11573,N_10250);
and U14349 (N_14349,N_9120,N_10728);
xnor U14350 (N_14350,N_10702,N_11756);
or U14351 (N_14351,N_11108,N_9816);
nor U14352 (N_14352,N_9867,N_10717);
nand U14353 (N_14353,N_11860,N_10666);
xor U14354 (N_14354,N_10253,N_11831);
or U14355 (N_14355,N_10939,N_9742);
and U14356 (N_14356,N_10410,N_10577);
nor U14357 (N_14357,N_9071,N_11309);
nand U14358 (N_14358,N_11995,N_11975);
or U14359 (N_14359,N_9382,N_11724);
xnor U14360 (N_14360,N_11859,N_10516);
nand U14361 (N_14361,N_9030,N_9802);
nor U14362 (N_14362,N_10745,N_9260);
xnor U14363 (N_14363,N_10312,N_9611);
xor U14364 (N_14364,N_10662,N_10379);
and U14365 (N_14365,N_9598,N_9409);
or U14366 (N_14366,N_9745,N_9293);
nor U14367 (N_14367,N_11205,N_9873);
nand U14368 (N_14368,N_10354,N_9007);
nor U14369 (N_14369,N_10491,N_11171);
nor U14370 (N_14370,N_11549,N_11892);
or U14371 (N_14371,N_11449,N_11224);
and U14372 (N_14372,N_9847,N_9532);
nor U14373 (N_14373,N_10566,N_10255);
and U14374 (N_14374,N_10582,N_10480);
nor U14375 (N_14375,N_11191,N_9107);
xor U14376 (N_14376,N_11097,N_10184);
and U14377 (N_14377,N_10548,N_9839);
nor U14378 (N_14378,N_11649,N_11806);
or U14379 (N_14379,N_9511,N_11865);
or U14380 (N_14380,N_10647,N_11124);
and U14381 (N_14381,N_10598,N_9287);
nand U14382 (N_14382,N_9978,N_9434);
nor U14383 (N_14383,N_11691,N_9978);
and U14384 (N_14384,N_11813,N_11025);
nor U14385 (N_14385,N_11672,N_9921);
nor U14386 (N_14386,N_9376,N_9369);
xor U14387 (N_14387,N_10417,N_10219);
nand U14388 (N_14388,N_9326,N_11135);
nor U14389 (N_14389,N_11791,N_11463);
or U14390 (N_14390,N_11950,N_9199);
nor U14391 (N_14391,N_10935,N_9355);
nand U14392 (N_14392,N_10899,N_9073);
xor U14393 (N_14393,N_9328,N_11095);
nor U14394 (N_14394,N_11601,N_10399);
xnor U14395 (N_14395,N_9971,N_11376);
nand U14396 (N_14396,N_10475,N_11667);
and U14397 (N_14397,N_9898,N_11220);
nor U14398 (N_14398,N_11155,N_9828);
nor U14399 (N_14399,N_9737,N_10870);
nor U14400 (N_14400,N_11889,N_10878);
or U14401 (N_14401,N_11160,N_9722);
nor U14402 (N_14402,N_10914,N_10720);
nor U14403 (N_14403,N_11238,N_11897);
nand U14404 (N_14404,N_11656,N_11436);
and U14405 (N_14405,N_9764,N_9691);
nand U14406 (N_14406,N_9672,N_9912);
xnor U14407 (N_14407,N_10411,N_9497);
nand U14408 (N_14408,N_10755,N_10056);
nor U14409 (N_14409,N_11667,N_10353);
nand U14410 (N_14410,N_10429,N_10091);
nor U14411 (N_14411,N_10381,N_10771);
nand U14412 (N_14412,N_10978,N_11235);
nand U14413 (N_14413,N_11393,N_11180);
and U14414 (N_14414,N_11067,N_11477);
nor U14415 (N_14415,N_10635,N_10168);
or U14416 (N_14416,N_11878,N_9098);
or U14417 (N_14417,N_9362,N_11369);
xnor U14418 (N_14418,N_9494,N_9630);
nor U14419 (N_14419,N_10866,N_10519);
xor U14420 (N_14420,N_9735,N_10975);
nand U14421 (N_14421,N_11964,N_11472);
nand U14422 (N_14422,N_11005,N_11382);
nand U14423 (N_14423,N_11063,N_11300);
xnor U14424 (N_14424,N_10116,N_10884);
nand U14425 (N_14425,N_10407,N_10604);
and U14426 (N_14426,N_11581,N_11325);
nor U14427 (N_14427,N_9940,N_10559);
or U14428 (N_14428,N_9735,N_10483);
xnor U14429 (N_14429,N_11867,N_10604);
and U14430 (N_14430,N_10707,N_11742);
nand U14431 (N_14431,N_11463,N_10998);
nand U14432 (N_14432,N_11844,N_9001);
nand U14433 (N_14433,N_11562,N_9409);
and U14434 (N_14434,N_9820,N_10251);
and U14435 (N_14435,N_10802,N_10448);
nor U14436 (N_14436,N_9292,N_11845);
xnor U14437 (N_14437,N_11627,N_9227);
nor U14438 (N_14438,N_11472,N_10081);
xnor U14439 (N_14439,N_10468,N_9852);
or U14440 (N_14440,N_11408,N_11128);
nand U14441 (N_14441,N_10056,N_9437);
or U14442 (N_14442,N_9316,N_10728);
and U14443 (N_14443,N_11396,N_9256);
nor U14444 (N_14444,N_10830,N_11141);
xnor U14445 (N_14445,N_10778,N_9246);
nand U14446 (N_14446,N_11835,N_10234);
nand U14447 (N_14447,N_10342,N_10425);
and U14448 (N_14448,N_10685,N_11552);
or U14449 (N_14449,N_11137,N_11828);
or U14450 (N_14450,N_10906,N_9410);
nor U14451 (N_14451,N_9359,N_10735);
or U14452 (N_14452,N_11414,N_9497);
xnor U14453 (N_14453,N_10112,N_11234);
nand U14454 (N_14454,N_9234,N_10775);
nand U14455 (N_14455,N_10810,N_9641);
nand U14456 (N_14456,N_11226,N_9917);
or U14457 (N_14457,N_9995,N_9746);
or U14458 (N_14458,N_9365,N_9893);
nor U14459 (N_14459,N_9746,N_11660);
xor U14460 (N_14460,N_9348,N_10346);
xnor U14461 (N_14461,N_10161,N_10646);
and U14462 (N_14462,N_10048,N_10303);
and U14463 (N_14463,N_10983,N_9883);
xor U14464 (N_14464,N_9737,N_10682);
nor U14465 (N_14465,N_9447,N_10753);
or U14466 (N_14466,N_9913,N_10308);
or U14467 (N_14467,N_9777,N_9582);
nand U14468 (N_14468,N_9821,N_9977);
xor U14469 (N_14469,N_11277,N_9322);
nand U14470 (N_14470,N_10704,N_10640);
and U14471 (N_14471,N_10570,N_11772);
and U14472 (N_14472,N_10390,N_11612);
nand U14473 (N_14473,N_11305,N_10308);
xor U14474 (N_14474,N_11543,N_10245);
nand U14475 (N_14475,N_10850,N_9683);
nand U14476 (N_14476,N_11756,N_9581);
nand U14477 (N_14477,N_9155,N_11871);
or U14478 (N_14478,N_9865,N_9226);
or U14479 (N_14479,N_11190,N_10431);
nand U14480 (N_14480,N_11836,N_11639);
and U14481 (N_14481,N_10573,N_11724);
and U14482 (N_14482,N_11185,N_9268);
or U14483 (N_14483,N_10610,N_11451);
or U14484 (N_14484,N_11060,N_10810);
nand U14485 (N_14485,N_11833,N_11953);
and U14486 (N_14486,N_11048,N_9849);
nor U14487 (N_14487,N_11582,N_11461);
nor U14488 (N_14488,N_9677,N_10637);
nor U14489 (N_14489,N_10853,N_9653);
nor U14490 (N_14490,N_10238,N_10777);
and U14491 (N_14491,N_9780,N_9897);
and U14492 (N_14492,N_9878,N_10365);
nand U14493 (N_14493,N_9534,N_11397);
nand U14494 (N_14494,N_10919,N_11366);
or U14495 (N_14495,N_10202,N_11267);
nor U14496 (N_14496,N_11055,N_9725);
nand U14497 (N_14497,N_9073,N_10307);
nor U14498 (N_14498,N_11494,N_10693);
and U14499 (N_14499,N_10822,N_9505);
or U14500 (N_14500,N_9422,N_10541);
nand U14501 (N_14501,N_11555,N_9898);
nand U14502 (N_14502,N_11839,N_9087);
xor U14503 (N_14503,N_11901,N_10367);
or U14504 (N_14504,N_11787,N_11470);
and U14505 (N_14505,N_10671,N_9822);
and U14506 (N_14506,N_9720,N_10639);
or U14507 (N_14507,N_10533,N_9403);
or U14508 (N_14508,N_9494,N_11562);
nand U14509 (N_14509,N_9906,N_9215);
nand U14510 (N_14510,N_9177,N_10373);
nor U14511 (N_14511,N_9555,N_10557);
and U14512 (N_14512,N_10064,N_10801);
and U14513 (N_14513,N_10723,N_9768);
nand U14514 (N_14514,N_9617,N_10876);
xnor U14515 (N_14515,N_10291,N_10210);
and U14516 (N_14516,N_10387,N_9429);
and U14517 (N_14517,N_11573,N_10279);
or U14518 (N_14518,N_11726,N_10259);
nor U14519 (N_14519,N_10669,N_11613);
xnor U14520 (N_14520,N_9426,N_10850);
and U14521 (N_14521,N_11330,N_10319);
nor U14522 (N_14522,N_11085,N_10641);
and U14523 (N_14523,N_9228,N_11367);
nand U14524 (N_14524,N_9612,N_10192);
or U14525 (N_14525,N_10482,N_10654);
xnor U14526 (N_14526,N_11454,N_10090);
nand U14527 (N_14527,N_11200,N_10117);
and U14528 (N_14528,N_11254,N_9854);
nor U14529 (N_14529,N_11002,N_9627);
and U14530 (N_14530,N_10369,N_10497);
and U14531 (N_14531,N_10005,N_11807);
nand U14532 (N_14532,N_11316,N_9116);
nand U14533 (N_14533,N_10822,N_11505);
nor U14534 (N_14534,N_11906,N_11475);
or U14535 (N_14535,N_10904,N_11314);
nand U14536 (N_14536,N_10937,N_10283);
nor U14537 (N_14537,N_10393,N_10317);
or U14538 (N_14538,N_11619,N_9010);
nand U14539 (N_14539,N_10691,N_11828);
or U14540 (N_14540,N_10981,N_10056);
xnor U14541 (N_14541,N_9409,N_9837);
nand U14542 (N_14542,N_10175,N_10405);
xor U14543 (N_14543,N_10770,N_10142);
xor U14544 (N_14544,N_11978,N_9315);
nand U14545 (N_14545,N_9395,N_11516);
or U14546 (N_14546,N_10192,N_9000);
xnor U14547 (N_14547,N_11278,N_10033);
nor U14548 (N_14548,N_10953,N_11944);
nor U14549 (N_14549,N_10832,N_9503);
and U14550 (N_14550,N_9807,N_10319);
nand U14551 (N_14551,N_9740,N_10824);
nor U14552 (N_14552,N_9317,N_9203);
nor U14553 (N_14553,N_10427,N_10955);
nand U14554 (N_14554,N_11548,N_11364);
nor U14555 (N_14555,N_9359,N_11822);
xor U14556 (N_14556,N_10232,N_9976);
or U14557 (N_14557,N_11813,N_9256);
xor U14558 (N_14558,N_10806,N_10855);
or U14559 (N_14559,N_11401,N_11496);
or U14560 (N_14560,N_10817,N_9203);
nor U14561 (N_14561,N_11630,N_9533);
xor U14562 (N_14562,N_11705,N_10681);
nand U14563 (N_14563,N_10700,N_9149);
nor U14564 (N_14564,N_10637,N_10332);
xor U14565 (N_14565,N_10366,N_11576);
xor U14566 (N_14566,N_9482,N_9415);
nor U14567 (N_14567,N_11911,N_11506);
xnor U14568 (N_14568,N_10842,N_11553);
xor U14569 (N_14569,N_10819,N_11248);
or U14570 (N_14570,N_9832,N_9072);
xor U14571 (N_14571,N_11710,N_10297);
or U14572 (N_14572,N_10292,N_9558);
and U14573 (N_14573,N_10813,N_9408);
or U14574 (N_14574,N_11729,N_9665);
nand U14575 (N_14575,N_10829,N_11548);
or U14576 (N_14576,N_10934,N_9135);
xnor U14577 (N_14577,N_9680,N_9789);
xnor U14578 (N_14578,N_10017,N_11146);
and U14579 (N_14579,N_9768,N_10379);
xor U14580 (N_14580,N_11388,N_11491);
or U14581 (N_14581,N_9217,N_10623);
nand U14582 (N_14582,N_9155,N_10232);
nand U14583 (N_14583,N_11973,N_11141);
nand U14584 (N_14584,N_10702,N_10984);
nor U14585 (N_14585,N_10054,N_10612);
and U14586 (N_14586,N_11917,N_10798);
nand U14587 (N_14587,N_9988,N_11537);
nor U14588 (N_14588,N_11596,N_10544);
xnor U14589 (N_14589,N_9219,N_10528);
xnor U14590 (N_14590,N_11267,N_10224);
or U14591 (N_14591,N_10295,N_10102);
or U14592 (N_14592,N_9163,N_9920);
nor U14593 (N_14593,N_10132,N_9835);
nor U14594 (N_14594,N_11814,N_11967);
or U14595 (N_14595,N_11678,N_9827);
or U14596 (N_14596,N_10887,N_9002);
and U14597 (N_14597,N_9488,N_9603);
nor U14598 (N_14598,N_10853,N_10966);
xor U14599 (N_14599,N_11342,N_9734);
and U14600 (N_14600,N_10885,N_9768);
nor U14601 (N_14601,N_10841,N_9924);
xor U14602 (N_14602,N_10322,N_11306);
xnor U14603 (N_14603,N_9095,N_10956);
and U14604 (N_14604,N_9157,N_10798);
xor U14605 (N_14605,N_9029,N_9761);
xor U14606 (N_14606,N_11040,N_11757);
and U14607 (N_14607,N_11494,N_9546);
xnor U14608 (N_14608,N_10594,N_9528);
or U14609 (N_14609,N_11589,N_9970);
xnor U14610 (N_14610,N_11395,N_10140);
xor U14611 (N_14611,N_9185,N_9956);
and U14612 (N_14612,N_11344,N_10401);
and U14613 (N_14613,N_11448,N_9920);
and U14614 (N_14614,N_9514,N_9088);
xor U14615 (N_14615,N_11685,N_9830);
or U14616 (N_14616,N_10989,N_10442);
nand U14617 (N_14617,N_9105,N_10295);
nor U14618 (N_14618,N_9306,N_11948);
or U14619 (N_14619,N_9778,N_10702);
nor U14620 (N_14620,N_11628,N_10891);
nand U14621 (N_14621,N_10767,N_10645);
or U14622 (N_14622,N_10320,N_11007);
or U14623 (N_14623,N_11767,N_10013);
nand U14624 (N_14624,N_11955,N_11226);
nor U14625 (N_14625,N_11139,N_10683);
nor U14626 (N_14626,N_11702,N_11718);
nor U14627 (N_14627,N_11295,N_10944);
nor U14628 (N_14628,N_9182,N_10837);
and U14629 (N_14629,N_10576,N_11779);
and U14630 (N_14630,N_9177,N_10555);
nor U14631 (N_14631,N_9012,N_9623);
xnor U14632 (N_14632,N_9457,N_10415);
xnor U14633 (N_14633,N_11320,N_10121);
nand U14634 (N_14634,N_9810,N_9011);
xor U14635 (N_14635,N_9220,N_10971);
or U14636 (N_14636,N_9330,N_10746);
nor U14637 (N_14637,N_10147,N_10911);
nand U14638 (N_14638,N_9568,N_9085);
xor U14639 (N_14639,N_11723,N_9964);
and U14640 (N_14640,N_11608,N_11116);
and U14641 (N_14641,N_9537,N_9398);
xor U14642 (N_14642,N_9930,N_9673);
nor U14643 (N_14643,N_9848,N_10965);
nor U14644 (N_14644,N_9204,N_11044);
nand U14645 (N_14645,N_10797,N_9228);
or U14646 (N_14646,N_9117,N_10135);
and U14647 (N_14647,N_11923,N_10576);
nand U14648 (N_14648,N_11809,N_10067);
nand U14649 (N_14649,N_10239,N_9447);
nor U14650 (N_14650,N_9303,N_9827);
nand U14651 (N_14651,N_9113,N_9036);
nor U14652 (N_14652,N_10152,N_10656);
or U14653 (N_14653,N_11522,N_10598);
or U14654 (N_14654,N_11358,N_9800);
nor U14655 (N_14655,N_11973,N_11474);
and U14656 (N_14656,N_10763,N_9707);
or U14657 (N_14657,N_9245,N_10705);
or U14658 (N_14658,N_9808,N_10713);
nor U14659 (N_14659,N_11661,N_9016);
nand U14660 (N_14660,N_11456,N_10020);
or U14661 (N_14661,N_11338,N_10083);
and U14662 (N_14662,N_10681,N_10410);
and U14663 (N_14663,N_10431,N_10365);
nand U14664 (N_14664,N_11716,N_11589);
and U14665 (N_14665,N_11245,N_9346);
or U14666 (N_14666,N_11613,N_11419);
xnor U14667 (N_14667,N_11299,N_9164);
xor U14668 (N_14668,N_9824,N_11345);
or U14669 (N_14669,N_11600,N_10705);
nand U14670 (N_14670,N_11284,N_11544);
or U14671 (N_14671,N_9071,N_10379);
nand U14672 (N_14672,N_10365,N_11263);
nand U14673 (N_14673,N_9985,N_10384);
nand U14674 (N_14674,N_11981,N_11716);
nand U14675 (N_14675,N_9506,N_9857);
and U14676 (N_14676,N_11569,N_11053);
xnor U14677 (N_14677,N_10812,N_9085);
xnor U14678 (N_14678,N_10722,N_9658);
nand U14679 (N_14679,N_9551,N_11697);
and U14680 (N_14680,N_9049,N_10493);
nand U14681 (N_14681,N_11922,N_10075);
and U14682 (N_14682,N_10227,N_10970);
nand U14683 (N_14683,N_10031,N_11311);
and U14684 (N_14684,N_9739,N_11840);
nand U14685 (N_14685,N_11879,N_11102);
xnor U14686 (N_14686,N_10356,N_9961);
nor U14687 (N_14687,N_10434,N_10606);
or U14688 (N_14688,N_11533,N_9369);
xor U14689 (N_14689,N_11456,N_10803);
nand U14690 (N_14690,N_9058,N_9445);
nor U14691 (N_14691,N_10439,N_11711);
xnor U14692 (N_14692,N_10056,N_10628);
xor U14693 (N_14693,N_9858,N_10246);
and U14694 (N_14694,N_9409,N_10149);
nor U14695 (N_14695,N_10629,N_11847);
and U14696 (N_14696,N_9926,N_11121);
nor U14697 (N_14697,N_9171,N_9573);
xnor U14698 (N_14698,N_11085,N_11404);
nand U14699 (N_14699,N_9758,N_10414);
or U14700 (N_14700,N_11988,N_9985);
and U14701 (N_14701,N_9826,N_10757);
and U14702 (N_14702,N_11200,N_9780);
or U14703 (N_14703,N_10383,N_11867);
nand U14704 (N_14704,N_11337,N_10401);
and U14705 (N_14705,N_11426,N_10920);
or U14706 (N_14706,N_9526,N_11007);
nor U14707 (N_14707,N_11231,N_10196);
nand U14708 (N_14708,N_11106,N_10349);
nand U14709 (N_14709,N_9053,N_9926);
nor U14710 (N_14710,N_11045,N_10876);
and U14711 (N_14711,N_11839,N_11553);
or U14712 (N_14712,N_10809,N_11012);
and U14713 (N_14713,N_10518,N_10242);
or U14714 (N_14714,N_10005,N_9286);
nor U14715 (N_14715,N_9737,N_11898);
nor U14716 (N_14716,N_11236,N_10462);
or U14717 (N_14717,N_9081,N_10951);
and U14718 (N_14718,N_10213,N_11552);
nor U14719 (N_14719,N_9088,N_9338);
nand U14720 (N_14720,N_10774,N_9613);
or U14721 (N_14721,N_10502,N_11735);
xor U14722 (N_14722,N_11452,N_9135);
and U14723 (N_14723,N_10933,N_9788);
nand U14724 (N_14724,N_11305,N_11927);
or U14725 (N_14725,N_9337,N_11317);
or U14726 (N_14726,N_11770,N_10136);
xnor U14727 (N_14727,N_10676,N_10637);
and U14728 (N_14728,N_11314,N_9629);
or U14729 (N_14729,N_9891,N_10120);
nand U14730 (N_14730,N_11106,N_11742);
nor U14731 (N_14731,N_10271,N_10592);
or U14732 (N_14732,N_10101,N_10137);
and U14733 (N_14733,N_9909,N_10847);
and U14734 (N_14734,N_9851,N_11230);
or U14735 (N_14735,N_10756,N_9900);
nand U14736 (N_14736,N_11967,N_10226);
or U14737 (N_14737,N_10652,N_9000);
and U14738 (N_14738,N_10650,N_10781);
xor U14739 (N_14739,N_11918,N_9128);
nor U14740 (N_14740,N_11394,N_10757);
or U14741 (N_14741,N_11290,N_10689);
xor U14742 (N_14742,N_9797,N_11799);
nand U14743 (N_14743,N_9202,N_11913);
xor U14744 (N_14744,N_10390,N_10192);
or U14745 (N_14745,N_9209,N_10925);
xnor U14746 (N_14746,N_9105,N_10629);
and U14747 (N_14747,N_11239,N_10937);
and U14748 (N_14748,N_11256,N_9697);
nand U14749 (N_14749,N_10654,N_10149);
and U14750 (N_14750,N_10131,N_10847);
or U14751 (N_14751,N_10161,N_9503);
nand U14752 (N_14752,N_11122,N_10965);
nand U14753 (N_14753,N_11462,N_9605);
or U14754 (N_14754,N_11908,N_9301);
nor U14755 (N_14755,N_9851,N_11687);
or U14756 (N_14756,N_11090,N_11951);
xor U14757 (N_14757,N_10693,N_10578);
xnor U14758 (N_14758,N_9361,N_10832);
xor U14759 (N_14759,N_11490,N_11796);
nand U14760 (N_14760,N_10664,N_10624);
nor U14761 (N_14761,N_11392,N_11481);
xnor U14762 (N_14762,N_9644,N_11579);
nor U14763 (N_14763,N_9875,N_11292);
and U14764 (N_14764,N_9058,N_9251);
xor U14765 (N_14765,N_11175,N_9882);
or U14766 (N_14766,N_11888,N_11286);
or U14767 (N_14767,N_10106,N_10032);
nand U14768 (N_14768,N_11145,N_10572);
or U14769 (N_14769,N_9799,N_9542);
and U14770 (N_14770,N_11039,N_11930);
and U14771 (N_14771,N_11733,N_10911);
nand U14772 (N_14772,N_10038,N_10431);
or U14773 (N_14773,N_9795,N_11147);
xor U14774 (N_14774,N_10031,N_10104);
or U14775 (N_14775,N_10929,N_9543);
nand U14776 (N_14776,N_9577,N_9410);
or U14777 (N_14777,N_11017,N_10258);
or U14778 (N_14778,N_9221,N_11133);
nor U14779 (N_14779,N_11441,N_9182);
nand U14780 (N_14780,N_9677,N_10448);
nor U14781 (N_14781,N_11178,N_10036);
or U14782 (N_14782,N_10864,N_10852);
xnor U14783 (N_14783,N_9800,N_10697);
and U14784 (N_14784,N_9292,N_11783);
nand U14785 (N_14785,N_10034,N_9450);
nor U14786 (N_14786,N_10043,N_11511);
and U14787 (N_14787,N_10463,N_10202);
xnor U14788 (N_14788,N_11370,N_10868);
or U14789 (N_14789,N_9742,N_11005);
and U14790 (N_14790,N_10835,N_9379);
xor U14791 (N_14791,N_9330,N_10947);
or U14792 (N_14792,N_9831,N_10973);
xor U14793 (N_14793,N_11961,N_10051);
nor U14794 (N_14794,N_9115,N_11881);
or U14795 (N_14795,N_11202,N_11522);
xor U14796 (N_14796,N_10121,N_10445);
nor U14797 (N_14797,N_11381,N_11746);
or U14798 (N_14798,N_9007,N_10053);
and U14799 (N_14799,N_10465,N_11129);
and U14800 (N_14800,N_11557,N_11683);
xnor U14801 (N_14801,N_9354,N_10170);
nand U14802 (N_14802,N_11241,N_11805);
xnor U14803 (N_14803,N_10221,N_10845);
or U14804 (N_14804,N_9779,N_10815);
xnor U14805 (N_14805,N_11377,N_9577);
xor U14806 (N_14806,N_11204,N_10966);
or U14807 (N_14807,N_11572,N_9235);
nand U14808 (N_14808,N_11521,N_9024);
nand U14809 (N_14809,N_10140,N_11131);
nor U14810 (N_14810,N_11339,N_9990);
or U14811 (N_14811,N_10350,N_11115);
and U14812 (N_14812,N_11781,N_11733);
nand U14813 (N_14813,N_10734,N_11250);
xor U14814 (N_14814,N_10759,N_10260);
nor U14815 (N_14815,N_9783,N_10844);
and U14816 (N_14816,N_11546,N_9791);
or U14817 (N_14817,N_10453,N_10749);
or U14818 (N_14818,N_9093,N_11430);
or U14819 (N_14819,N_9725,N_9999);
or U14820 (N_14820,N_11292,N_9498);
nor U14821 (N_14821,N_10488,N_9870);
or U14822 (N_14822,N_10229,N_9061);
or U14823 (N_14823,N_10138,N_10356);
nand U14824 (N_14824,N_10443,N_10560);
and U14825 (N_14825,N_11373,N_10854);
and U14826 (N_14826,N_10773,N_10912);
xnor U14827 (N_14827,N_9866,N_9071);
xor U14828 (N_14828,N_11922,N_11588);
or U14829 (N_14829,N_9058,N_9588);
or U14830 (N_14830,N_10639,N_11043);
and U14831 (N_14831,N_10734,N_9414);
nand U14832 (N_14832,N_10428,N_9906);
xnor U14833 (N_14833,N_10417,N_9117);
xor U14834 (N_14834,N_9559,N_9957);
or U14835 (N_14835,N_10449,N_11771);
xnor U14836 (N_14836,N_11680,N_11911);
nor U14837 (N_14837,N_10064,N_11604);
nor U14838 (N_14838,N_10626,N_9934);
and U14839 (N_14839,N_10557,N_9334);
xnor U14840 (N_14840,N_10321,N_10650);
xnor U14841 (N_14841,N_11024,N_11949);
nand U14842 (N_14842,N_11083,N_11774);
nand U14843 (N_14843,N_10794,N_11532);
nand U14844 (N_14844,N_9551,N_9048);
or U14845 (N_14845,N_10976,N_10248);
nand U14846 (N_14846,N_9243,N_10230);
xnor U14847 (N_14847,N_9170,N_10000);
xor U14848 (N_14848,N_10534,N_9473);
nand U14849 (N_14849,N_11854,N_11092);
nor U14850 (N_14850,N_11715,N_11925);
nand U14851 (N_14851,N_11985,N_9476);
nor U14852 (N_14852,N_10072,N_9262);
nor U14853 (N_14853,N_9461,N_11432);
xor U14854 (N_14854,N_9084,N_10278);
nor U14855 (N_14855,N_10383,N_10629);
nand U14856 (N_14856,N_10783,N_10929);
xor U14857 (N_14857,N_11579,N_9692);
nor U14858 (N_14858,N_11775,N_11784);
nand U14859 (N_14859,N_10555,N_9465);
nor U14860 (N_14860,N_10859,N_11292);
xnor U14861 (N_14861,N_11538,N_11330);
or U14862 (N_14862,N_11251,N_10611);
and U14863 (N_14863,N_11546,N_10658);
or U14864 (N_14864,N_11496,N_10758);
or U14865 (N_14865,N_11699,N_10285);
nor U14866 (N_14866,N_11450,N_9026);
xor U14867 (N_14867,N_11582,N_10712);
nor U14868 (N_14868,N_10078,N_11214);
and U14869 (N_14869,N_9993,N_9877);
and U14870 (N_14870,N_11006,N_9030);
xor U14871 (N_14871,N_9198,N_9068);
nand U14872 (N_14872,N_10230,N_10843);
xor U14873 (N_14873,N_10557,N_10773);
and U14874 (N_14874,N_9276,N_9508);
or U14875 (N_14875,N_10201,N_11249);
nand U14876 (N_14876,N_10652,N_10003);
nor U14877 (N_14877,N_11920,N_11766);
and U14878 (N_14878,N_11048,N_9135);
xor U14879 (N_14879,N_11490,N_10188);
nor U14880 (N_14880,N_11730,N_11070);
nand U14881 (N_14881,N_11857,N_11301);
nand U14882 (N_14882,N_9354,N_9085);
or U14883 (N_14883,N_11771,N_9676);
nand U14884 (N_14884,N_9878,N_11111);
nand U14885 (N_14885,N_9693,N_11161);
nand U14886 (N_14886,N_11038,N_9567);
xor U14887 (N_14887,N_9798,N_9329);
nand U14888 (N_14888,N_9272,N_9923);
or U14889 (N_14889,N_10448,N_9398);
xnor U14890 (N_14890,N_11959,N_10961);
and U14891 (N_14891,N_9957,N_11697);
nor U14892 (N_14892,N_10744,N_11517);
xor U14893 (N_14893,N_9307,N_10888);
or U14894 (N_14894,N_10624,N_10225);
nand U14895 (N_14895,N_10573,N_11687);
and U14896 (N_14896,N_10959,N_11064);
or U14897 (N_14897,N_9647,N_10577);
nand U14898 (N_14898,N_11938,N_9024);
nor U14899 (N_14899,N_10091,N_10635);
nand U14900 (N_14900,N_10566,N_11981);
xnor U14901 (N_14901,N_9731,N_10331);
xor U14902 (N_14902,N_11229,N_9106);
nand U14903 (N_14903,N_9351,N_11144);
nand U14904 (N_14904,N_11329,N_10568);
or U14905 (N_14905,N_10214,N_10071);
or U14906 (N_14906,N_11075,N_10191);
nor U14907 (N_14907,N_9965,N_11291);
xor U14908 (N_14908,N_9574,N_10055);
nand U14909 (N_14909,N_10839,N_11577);
nand U14910 (N_14910,N_11210,N_9003);
nor U14911 (N_14911,N_9791,N_11317);
xnor U14912 (N_14912,N_9788,N_9401);
nand U14913 (N_14913,N_9435,N_10375);
nand U14914 (N_14914,N_9090,N_11585);
and U14915 (N_14915,N_11839,N_11948);
xor U14916 (N_14916,N_9948,N_9615);
and U14917 (N_14917,N_10219,N_9097);
nor U14918 (N_14918,N_10517,N_10974);
xnor U14919 (N_14919,N_11938,N_10473);
nand U14920 (N_14920,N_10903,N_10788);
and U14921 (N_14921,N_9068,N_10460);
or U14922 (N_14922,N_9389,N_10634);
or U14923 (N_14923,N_11304,N_10845);
and U14924 (N_14924,N_9684,N_11015);
nor U14925 (N_14925,N_9172,N_11896);
or U14926 (N_14926,N_9671,N_11906);
nand U14927 (N_14927,N_10961,N_11032);
and U14928 (N_14928,N_10208,N_10040);
and U14929 (N_14929,N_9642,N_10705);
nor U14930 (N_14930,N_9268,N_10319);
xnor U14931 (N_14931,N_10328,N_11548);
nand U14932 (N_14932,N_10471,N_10331);
xnor U14933 (N_14933,N_11380,N_10984);
nand U14934 (N_14934,N_9707,N_11483);
and U14935 (N_14935,N_9859,N_9076);
nand U14936 (N_14936,N_10834,N_10447);
and U14937 (N_14937,N_9203,N_9806);
and U14938 (N_14938,N_11534,N_9604);
nor U14939 (N_14939,N_10832,N_9727);
xnor U14940 (N_14940,N_10020,N_11108);
nand U14941 (N_14941,N_9814,N_10366);
or U14942 (N_14942,N_11597,N_9290);
and U14943 (N_14943,N_9355,N_9965);
or U14944 (N_14944,N_10308,N_9396);
or U14945 (N_14945,N_10266,N_11528);
nor U14946 (N_14946,N_11628,N_10629);
nor U14947 (N_14947,N_11714,N_11169);
xnor U14948 (N_14948,N_9972,N_11340);
nand U14949 (N_14949,N_9937,N_11601);
or U14950 (N_14950,N_9027,N_9407);
and U14951 (N_14951,N_10466,N_11528);
and U14952 (N_14952,N_10320,N_10165);
nand U14953 (N_14953,N_11807,N_11296);
xnor U14954 (N_14954,N_9287,N_10825);
xor U14955 (N_14955,N_10684,N_9183);
nand U14956 (N_14956,N_11000,N_9095);
xor U14957 (N_14957,N_9649,N_10736);
and U14958 (N_14958,N_11494,N_9980);
nand U14959 (N_14959,N_11019,N_11983);
and U14960 (N_14960,N_10274,N_11607);
or U14961 (N_14961,N_10950,N_9415);
nand U14962 (N_14962,N_11548,N_10782);
xor U14963 (N_14963,N_10603,N_9866);
nand U14964 (N_14964,N_9351,N_11643);
nor U14965 (N_14965,N_10876,N_11583);
nand U14966 (N_14966,N_10596,N_11296);
nor U14967 (N_14967,N_10325,N_9373);
nand U14968 (N_14968,N_11025,N_9056);
nor U14969 (N_14969,N_10382,N_11168);
xnor U14970 (N_14970,N_11159,N_9315);
and U14971 (N_14971,N_11539,N_11261);
or U14972 (N_14972,N_10232,N_10658);
nand U14973 (N_14973,N_11995,N_11561);
nand U14974 (N_14974,N_11569,N_11654);
xnor U14975 (N_14975,N_11837,N_10280);
xor U14976 (N_14976,N_11916,N_9289);
or U14977 (N_14977,N_11390,N_11815);
or U14978 (N_14978,N_9182,N_11479);
or U14979 (N_14979,N_10092,N_11949);
nand U14980 (N_14980,N_10681,N_11027);
nor U14981 (N_14981,N_10368,N_11165);
and U14982 (N_14982,N_11111,N_11538);
nor U14983 (N_14983,N_9400,N_11122);
xor U14984 (N_14984,N_10863,N_10790);
xor U14985 (N_14985,N_10145,N_10272);
nor U14986 (N_14986,N_11284,N_10560);
or U14987 (N_14987,N_11290,N_10672);
xor U14988 (N_14988,N_11585,N_10250);
or U14989 (N_14989,N_11290,N_11925);
and U14990 (N_14990,N_9713,N_10679);
xnor U14991 (N_14991,N_9528,N_10011);
xor U14992 (N_14992,N_10508,N_10593);
xnor U14993 (N_14993,N_9796,N_9741);
or U14994 (N_14994,N_10236,N_10889);
and U14995 (N_14995,N_10923,N_10474);
xor U14996 (N_14996,N_9587,N_9173);
or U14997 (N_14997,N_9206,N_11720);
xor U14998 (N_14998,N_10368,N_11549);
or U14999 (N_14999,N_10912,N_11035);
and UO_0 (O_0,N_12217,N_13137);
xor UO_1 (O_1,N_12630,N_13806);
or UO_2 (O_2,N_14966,N_13290);
and UO_3 (O_3,N_14564,N_14175);
xor UO_4 (O_4,N_13065,N_13502);
and UO_5 (O_5,N_12895,N_13033);
nor UO_6 (O_6,N_14565,N_13061);
and UO_7 (O_7,N_12522,N_13251);
nand UO_8 (O_8,N_12908,N_12806);
nor UO_9 (O_9,N_13490,N_14082);
and UO_10 (O_10,N_13935,N_14752);
and UO_11 (O_11,N_12305,N_12225);
xnor UO_12 (O_12,N_14091,N_13788);
or UO_13 (O_13,N_14078,N_13712);
nor UO_14 (O_14,N_13909,N_14346);
xnor UO_15 (O_15,N_14363,N_14669);
nor UO_16 (O_16,N_12770,N_13482);
and UO_17 (O_17,N_14526,N_12061);
and UO_18 (O_18,N_14786,N_13441);
or UO_19 (O_19,N_14248,N_12173);
nor UO_20 (O_20,N_13354,N_12257);
nor UO_21 (O_21,N_12476,N_14465);
xnor UO_22 (O_22,N_12366,N_12104);
xor UO_23 (O_23,N_13440,N_14069);
xor UO_24 (O_24,N_14320,N_14850);
and UO_25 (O_25,N_14764,N_12315);
or UO_26 (O_26,N_12206,N_12262);
or UO_27 (O_27,N_12538,N_13685);
nor UO_28 (O_28,N_12736,N_14234);
and UO_29 (O_29,N_13604,N_13116);
xnor UO_30 (O_30,N_12775,N_12319);
xnor UO_31 (O_31,N_13901,N_12480);
and UO_32 (O_32,N_14798,N_13207);
and UO_33 (O_33,N_13467,N_13107);
or UO_34 (O_34,N_14173,N_13631);
nor UO_35 (O_35,N_14802,N_14781);
xor UO_36 (O_36,N_14751,N_13818);
nand UO_37 (O_37,N_13808,N_14704);
nand UO_38 (O_38,N_14235,N_13851);
and UO_39 (O_39,N_14260,N_13573);
or UO_40 (O_40,N_13980,N_12232);
xor UO_41 (O_41,N_14128,N_13224);
or UO_42 (O_42,N_14711,N_13105);
nand UO_43 (O_43,N_13549,N_12561);
nand UO_44 (O_44,N_14858,N_13465);
nor UO_45 (O_45,N_12082,N_12479);
and UO_46 (O_46,N_12750,N_14596);
nor UO_47 (O_47,N_13991,N_13182);
or UO_48 (O_48,N_13123,N_13929);
and UO_49 (O_49,N_13617,N_14396);
and UO_50 (O_50,N_13072,N_14199);
nand UO_51 (O_51,N_12326,N_13134);
nand UO_52 (O_52,N_14827,N_12610);
nor UO_53 (O_53,N_14093,N_13443);
nor UO_54 (O_54,N_13176,N_13825);
nor UO_55 (O_55,N_12518,N_12752);
and UO_56 (O_56,N_14575,N_13492);
nor UO_57 (O_57,N_12245,N_13816);
or UO_58 (O_58,N_13800,N_13704);
xor UO_59 (O_59,N_14950,N_12352);
xor UO_60 (O_60,N_13879,N_12025);
xor UO_61 (O_61,N_13585,N_14621);
xor UO_62 (O_62,N_12491,N_14723);
and UO_63 (O_63,N_12397,N_13041);
nor UO_64 (O_64,N_12608,N_12194);
nor UO_65 (O_65,N_14187,N_14815);
or UO_66 (O_66,N_12556,N_12488);
or UO_67 (O_67,N_14369,N_14989);
or UO_68 (O_68,N_12696,N_14608);
and UO_69 (O_69,N_13097,N_13200);
and UO_70 (O_70,N_12048,N_14887);
and UO_71 (O_71,N_12815,N_13472);
xor UO_72 (O_72,N_14624,N_12286);
nand UO_73 (O_73,N_14742,N_12125);
nor UO_74 (O_74,N_12606,N_13510);
nand UO_75 (O_75,N_12541,N_13646);
nand UO_76 (O_76,N_12673,N_14415);
xnor UO_77 (O_77,N_14634,N_14744);
nor UO_78 (O_78,N_13367,N_13821);
xor UO_79 (O_79,N_13498,N_12519);
or UO_80 (O_80,N_14698,N_14637);
xor UO_81 (O_81,N_13770,N_12951);
or UO_82 (O_82,N_13075,N_13926);
and UO_83 (O_83,N_14072,N_12439);
nor UO_84 (O_84,N_12228,N_12391);
or UO_85 (O_85,N_13272,N_12495);
nor UO_86 (O_86,N_13986,N_12502);
nand UO_87 (O_87,N_12337,N_12621);
and UO_88 (O_88,N_13539,N_13691);
or UO_89 (O_89,N_14216,N_13512);
nor UO_90 (O_90,N_12080,N_12791);
xnor UO_91 (O_91,N_14108,N_14374);
and UO_92 (O_92,N_14405,N_12186);
nand UO_93 (O_93,N_13168,N_14993);
and UO_94 (O_94,N_12669,N_13535);
and UO_95 (O_95,N_12230,N_13634);
and UO_96 (O_96,N_13130,N_13974);
nand UO_97 (O_97,N_13811,N_12546);
nor UO_98 (O_98,N_12364,N_13464);
or UO_99 (O_99,N_13608,N_12441);
and UO_100 (O_100,N_13112,N_14452);
xnor UO_101 (O_101,N_14653,N_12953);
nand UO_102 (O_102,N_13532,N_13504);
xor UO_103 (O_103,N_13639,N_14677);
and UO_104 (O_104,N_14506,N_13673);
nand UO_105 (O_105,N_13771,N_12345);
nand UO_106 (O_106,N_14172,N_14541);
or UO_107 (O_107,N_13835,N_12301);
xor UO_108 (O_108,N_13192,N_14717);
nand UO_109 (O_109,N_13841,N_13454);
nor UO_110 (O_110,N_13344,N_14514);
nand UO_111 (O_111,N_14103,N_12701);
and UO_112 (O_112,N_12901,N_14951);
or UO_113 (O_113,N_12427,N_12341);
and UO_114 (O_114,N_14807,N_14992);
nand UO_115 (O_115,N_12207,N_14042);
nor UO_116 (O_116,N_13784,N_14762);
or UO_117 (O_117,N_12818,N_13892);
xor UO_118 (O_118,N_12498,N_13042);
nand UO_119 (O_119,N_14979,N_13180);
nor UO_120 (O_120,N_12725,N_13270);
and UO_121 (O_121,N_14052,N_13777);
or UO_122 (O_122,N_12184,N_14694);
xor UO_123 (O_123,N_13320,N_12654);
nand UO_124 (O_124,N_13775,N_14083);
nand UO_125 (O_125,N_12849,N_13106);
nand UO_126 (O_126,N_12607,N_14144);
or UO_127 (O_127,N_12848,N_14530);
and UO_128 (O_128,N_14321,N_12963);
nor UO_129 (O_129,N_14371,N_13473);
nor UO_130 (O_130,N_12619,N_14382);
nand UO_131 (O_131,N_12764,N_13908);
and UO_132 (O_132,N_14423,N_13526);
nor UO_133 (O_133,N_13247,N_14229);
nor UO_134 (O_134,N_12302,N_13726);
or UO_135 (O_135,N_13150,N_13032);
or UO_136 (O_136,N_12615,N_14462);
xor UO_137 (O_137,N_12066,N_13566);
and UO_138 (O_138,N_13397,N_13419);
nand UO_139 (O_139,N_14376,N_14599);
nor UO_140 (O_140,N_13206,N_12042);
or UO_141 (O_141,N_12322,N_14963);
nor UO_142 (O_142,N_12817,N_12943);
nor UO_143 (O_143,N_13491,N_14714);
nor UO_144 (O_144,N_13735,N_12112);
nand UO_145 (O_145,N_12907,N_12704);
nand UO_146 (O_146,N_12841,N_14336);
nor UO_147 (O_147,N_13853,N_12708);
or UO_148 (O_148,N_14882,N_13556);
or UO_149 (O_149,N_14293,N_14839);
or UO_150 (O_150,N_13794,N_12292);
or UO_151 (O_151,N_14194,N_12832);
nand UO_152 (O_152,N_14112,N_13342);
xor UO_153 (O_153,N_13462,N_13244);
or UO_154 (O_154,N_12497,N_13546);
or UO_155 (O_155,N_14883,N_13776);
xor UO_156 (O_156,N_12827,N_12467);
nand UO_157 (O_157,N_12967,N_14058);
or UO_158 (O_158,N_14618,N_14748);
nand UO_159 (O_159,N_14613,N_12244);
and UO_160 (O_160,N_13749,N_13972);
and UO_161 (O_161,N_14094,N_14038);
xor UO_162 (O_162,N_14425,N_12779);
or UO_163 (O_163,N_14603,N_12418);
nand UO_164 (O_164,N_13621,N_13311);
nor UO_165 (O_165,N_14349,N_13830);
xnor UO_166 (O_166,N_12380,N_12012);
nand UO_167 (O_167,N_14885,N_12079);
nor UO_168 (O_168,N_14693,N_13804);
nand UO_169 (O_169,N_12393,N_14005);
xor UO_170 (O_170,N_14829,N_13678);
xor UO_171 (O_171,N_13162,N_13839);
xor UO_172 (O_172,N_12989,N_14746);
xor UO_173 (O_173,N_12800,N_14870);
or UO_174 (O_174,N_12904,N_14952);
or UO_175 (O_175,N_12124,N_14844);
xor UO_176 (O_176,N_12512,N_13852);
or UO_177 (O_177,N_14645,N_13667);
xor UO_178 (O_178,N_13336,N_14967);
nor UO_179 (O_179,N_12471,N_14962);
xnor UO_180 (O_180,N_14011,N_12369);
nand UO_181 (O_181,N_14939,N_12636);
or UO_182 (O_182,N_12202,N_12898);
xor UO_183 (O_183,N_14857,N_13897);
nor UO_184 (O_184,N_14337,N_13188);
nor UO_185 (O_185,N_14938,N_14877);
or UO_186 (O_186,N_13923,N_14820);
or UO_187 (O_187,N_12043,N_14237);
and UO_188 (O_188,N_12870,N_14045);
or UO_189 (O_189,N_13423,N_14995);
nor UO_190 (O_190,N_13199,N_14214);
and UO_191 (O_191,N_13226,N_13717);
xnor UO_192 (O_192,N_12069,N_13907);
nor UO_193 (O_193,N_13672,N_13094);
nor UO_194 (O_194,N_13683,N_13073);
and UO_195 (O_195,N_13418,N_12600);
nand UO_196 (O_196,N_12576,N_14410);
xor UO_197 (O_197,N_13316,N_13999);
nor UO_198 (O_198,N_12761,N_12405);
or UO_199 (O_199,N_14206,N_12068);
xor UO_200 (O_200,N_13607,N_12277);
and UO_201 (O_201,N_13475,N_12390);
nand UO_202 (O_202,N_12762,N_14907);
nand UO_203 (O_203,N_13092,N_13402);
nand UO_204 (O_204,N_12182,N_14500);
or UO_205 (O_205,N_13362,N_14016);
xnor UO_206 (O_206,N_12067,N_14513);
nor UO_207 (O_207,N_14957,N_14115);
and UO_208 (O_208,N_13417,N_13594);
xnor UO_209 (O_209,N_14988,N_12490);
and UO_210 (O_210,N_13146,N_14310);
and UO_211 (O_211,N_13438,N_14440);
nor UO_212 (O_212,N_12647,N_13896);
nor UO_213 (O_213,N_14118,N_13763);
nor UO_214 (O_214,N_12516,N_12887);
xnor UO_215 (O_215,N_14441,N_12771);
nand UO_216 (O_216,N_14239,N_14292);
nand UO_217 (O_217,N_12440,N_14166);
or UO_218 (O_218,N_12598,N_14426);
nand UO_219 (O_219,N_13317,N_13355);
nand UO_220 (O_220,N_12039,N_13343);
nand UO_221 (O_221,N_12313,N_13487);
nand UO_222 (O_222,N_12999,N_12937);
xor UO_223 (O_223,N_13541,N_12246);
nand UO_224 (O_224,N_12002,N_13627);
nand UO_225 (O_225,N_13846,N_14546);
and UO_226 (O_226,N_14648,N_14322);
nand UO_227 (O_227,N_12683,N_12871);
and UO_228 (O_228,N_14906,N_12671);
nand UO_229 (O_229,N_14153,N_12551);
nand UO_230 (O_230,N_14889,N_14975);
and UO_231 (O_231,N_14960,N_12339);
nand UO_232 (O_232,N_14976,N_12719);
and UO_233 (O_233,N_14490,N_14431);
and UO_234 (O_234,N_13714,N_12765);
and UO_235 (O_235,N_13826,N_12991);
and UO_236 (O_236,N_14602,N_13345);
and UO_237 (O_237,N_13086,N_13111);
nand UO_238 (O_238,N_13327,N_14463);
nand UO_239 (O_239,N_12142,N_14804);
xor UO_240 (O_240,N_14845,N_14605);
nor UO_241 (O_241,N_13005,N_13881);
and UO_242 (O_242,N_14587,N_12709);
or UO_243 (O_243,N_14551,N_13817);
nand UO_244 (O_244,N_14826,N_14550);
or UO_245 (O_245,N_12836,N_13420);
xnor UO_246 (O_246,N_13873,N_14201);
or UO_247 (O_247,N_12422,N_13956);
nand UO_248 (O_248,N_14945,N_13283);
and UO_249 (O_249,N_12521,N_12674);
xor UO_250 (O_250,N_14417,N_14429);
and UO_251 (O_251,N_13891,N_12306);
and UO_252 (O_252,N_12013,N_12811);
xnor UO_253 (O_253,N_12562,N_13983);
or UO_254 (O_254,N_13118,N_12549);
nand UO_255 (O_255,N_12289,N_13968);
and UO_256 (O_256,N_14317,N_14935);
nand UO_257 (O_257,N_14604,N_13476);
and UO_258 (O_258,N_13214,N_13758);
or UO_259 (O_259,N_12094,N_14066);
nand UO_260 (O_260,N_14563,N_14033);
nor UO_261 (O_261,N_12947,N_13383);
xnor UO_262 (O_262,N_14443,N_13941);
or UO_263 (O_263,N_14539,N_12592);
and UO_264 (O_264,N_14942,N_13700);
or UO_265 (O_265,N_14508,N_13727);
nand UO_266 (O_266,N_14155,N_14584);
nor UO_267 (O_267,N_13738,N_14932);
nand UO_268 (O_268,N_14198,N_12411);
or UO_269 (O_269,N_13082,N_12846);
nand UO_270 (O_270,N_14344,N_13411);
and UO_271 (O_271,N_14049,N_12987);
and UO_272 (O_272,N_12156,N_13364);
xnor UO_273 (O_273,N_12220,N_13016);
xnor UO_274 (O_274,N_14903,N_13857);
and UO_275 (O_275,N_13630,N_14543);
xor UO_276 (O_276,N_14763,N_13981);
nor UO_277 (O_277,N_12119,N_13401);
nor UO_278 (O_278,N_13416,N_13074);
xnor UO_279 (O_279,N_12948,N_13715);
xnor UO_280 (O_280,N_12567,N_14837);
or UO_281 (O_281,N_12945,N_12501);
or UO_282 (O_282,N_14135,N_13866);
nand UO_283 (O_283,N_14361,N_13480);
nand UO_284 (O_284,N_13921,N_14895);
and UO_285 (O_285,N_12523,N_14614);
and UO_286 (O_286,N_13944,N_13024);
or UO_287 (O_287,N_13071,N_14771);
nand UO_288 (O_288,N_13733,N_13632);
nand UO_289 (O_289,N_13893,N_13305);
xor UO_290 (O_290,N_12477,N_14666);
nand UO_291 (O_291,N_13414,N_13643);
nand UO_292 (O_292,N_13792,N_14394);
nor UO_293 (O_293,N_13867,N_14330);
and UO_294 (O_294,N_12392,N_14088);
or UO_295 (O_295,N_14619,N_13133);
nor UO_296 (O_296,N_13553,N_14690);
xor UO_297 (O_297,N_12912,N_13596);
xnor UO_298 (O_298,N_14811,N_12539);
and UO_299 (O_299,N_14727,N_13756);
or UO_300 (O_300,N_12348,N_12197);
or UO_301 (O_301,N_12215,N_13185);
xor UO_302 (O_302,N_14097,N_12545);
or UO_303 (O_303,N_14222,N_14110);
or UO_304 (O_304,N_12457,N_12766);
or UO_305 (O_305,N_14672,N_12687);
nor UO_306 (O_306,N_14721,N_13790);
xor UO_307 (O_307,N_14847,N_13959);
nand UO_308 (O_308,N_14209,N_12312);
or UO_309 (O_309,N_12446,N_14912);
xor UO_310 (O_310,N_14085,N_12227);
or UO_311 (O_311,N_12755,N_13789);
nor UO_312 (O_312,N_13842,N_12417);
nand UO_313 (O_313,N_14842,N_14456);
and UO_314 (O_314,N_13064,N_13212);
xor UO_315 (O_315,N_13521,N_14778);
xor UO_316 (O_316,N_14611,N_13698);
xnor UO_317 (O_317,N_12645,N_14079);
nor UO_318 (O_318,N_12604,N_12639);
and UO_319 (O_319,N_13151,N_12022);
nor UO_320 (O_320,N_13237,N_14205);
nor UO_321 (O_321,N_14174,N_12127);
and UO_322 (O_322,N_14986,N_13095);
xor UO_323 (O_323,N_14731,N_12078);
xnor UO_324 (O_324,N_13989,N_13353);
and UO_325 (O_325,N_14557,N_13201);
nor UO_326 (O_326,N_13755,N_14638);
nand UO_327 (O_327,N_14768,N_13163);
and UO_328 (O_328,N_13127,N_14354);
nand UO_329 (O_329,N_13970,N_14958);
nand UO_330 (O_330,N_12075,N_12782);
nand UO_331 (O_331,N_12367,N_13936);
nor UO_332 (O_332,N_13950,N_14105);
xor UO_333 (O_333,N_13805,N_14338);
or UO_334 (O_334,N_14294,N_14535);
or UO_335 (O_335,N_12087,N_12796);
and UO_336 (O_336,N_12862,N_12327);
and UO_337 (O_337,N_12885,N_14809);
or UO_338 (O_338,N_12040,N_14560);
or UO_339 (O_339,N_14300,N_14961);
nand UO_340 (O_340,N_12627,N_14032);
nor UO_341 (O_341,N_12726,N_12196);
and UO_342 (O_342,N_13572,N_14039);
or UO_343 (O_343,N_14077,N_14245);
nor UO_344 (O_344,N_13753,N_13450);
xor UO_345 (O_345,N_13508,N_14503);
and UO_346 (O_346,N_12651,N_12279);
nor UO_347 (O_347,N_13910,N_12083);
or UO_348 (O_348,N_13413,N_12992);
nand UO_349 (O_349,N_13388,N_12475);
nor UO_350 (O_350,N_14424,N_12425);
and UO_351 (O_351,N_13503,N_13149);
nand UO_352 (O_352,N_13298,N_13705);
nand UO_353 (O_353,N_12748,N_14994);
nor UO_354 (O_354,N_12926,N_14190);
nand UO_355 (O_355,N_14460,N_12866);
xor UO_356 (O_356,N_14578,N_13276);
nor UO_357 (O_357,N_13445,N_14674);
and UO_358 (O_358,N_13593,N_12136);
xor UO_359 (O_359,N_12860,N_14348);
nand UO_360 (O_360,N_12029,N_13459);
xnor UO_361 (O_361,N_13113,N_13729);
nand UO_362 (O_362,N_14197,N_12448);
xnor UO_363 (O_363,N_12178,N_14092);
xor UO_364 (O_364,N_12915,N_14387);
and UO_365 (O_365,N_13716,N_13040);
nand UO_366 (O_366,N_12413,N_12208);
or UO_367 (O_367,N_12238,N_13122);
xnor UO_368 (O_368,N_13523,N_13096);
and UO_369 (O_369,N_12805,N_13170);
nand UO_370 (O_370,N_12065,N_12387);
nor UO_371 (O_371,N_12930,N_13529);
nor UO_372 (O_372,N_14521,N_14357);
and UO_373 (O_373,N_13091,N_12020);
xor UO_374 (O_374,N_12381,N_13507);
xor UO_375 (O_375,N_12646,N_13942);
or UO_376 (O_376,N_12675,N_13554);
or UO_377 (O_377,N_12580,N_14356);
nand UO_378 (O_378,N_14664,N_13937);
nand UO_379 (O_379,N_14444,N_14267);
or UO_380 (O_380,N_14304,N_13385);
xnor UO_381 (O_381,N_12459,N_14326);
and UO_382 (O_382,N_13571,N_14136);
nand UO_383 (O_383,N_13590,N_13348);
nor UO_384 (O_384,N_13550,N_12874);
xnor UO_385 (O_385,N_14832,N_14592);
xnor UO_386 (O_386,N_13056,N_13222);
nand UO_387 (O_387,N_12176,N_14678);
and UO_388 (O_388,N_14707,N_12095);
nor UO_389 (O_389,N_12064,N_14902);
or UO_390 (O_390,N_13931,N_13679);
or UO_391 (O_391,N_14428,N_12308);
nor UO_392 (O_392,N_13802,N_12685);
nor UO_393 (O_393,N_12650,N_13647);
xor UO_394 (O_394,N_13747,N_12853);
nor UO_395 (O_395,N_14439,N_14397);
nand UO_396 (O_396,N_13325,N_12557);
xor UO_397 (O_397,N_12754,N_14099);
xor UO_398 (O_398,N_13292,N_13813);
nor UO_399 (O_399,N_12211,N_14623);
nor UO_400 (O_400,N_13680,N_12702);
or UO_401 (O_401,N_14914,N_13469);
and UO_402 (O_402,N_13803,N_12378);
nand UO_403 (O_403,N_12118,N_12547);
and UO_404 (O_404,N_14341,N_12834);
xor UO_405 (O_405,N_14133,N_12404);
nor UO_406 (O_406,N_12310,N_12278);
nand UO_407 (O_407,N_12192,N_12788);
nand UO_408 (O_408,N_13053,N_13474);
xor UO_409 (O_409,N_13511,N_12251);
and UO_410 (O_410,N_13046,N_14864);
and UO_411 (O_411,N_12642,N_13169);
xnor UO_412 (O_412,N_13245,N_12810);
nand UO_413 (O_413,N_13990,N_12216);
or UO_414 (O_414,N_14542,N_12993);
or UO_415 (O_415,N_13648,N_12285);
or UO_416 (O_416,N_12299,N_13628);
xor UO_417 (O_417,N_12548,N_14067);
xor UO_418 (O_418,N_13204,N_13155);
or UO_419 (O_419,N_13856,N_14185);
xnor UO_420 (O_420,N_12955,N_14745);
and UO_421 (O_421,N_14287,N_12062);
xnor UO_422 (O_422,N_12485,N_12699);
or UO_423 (O_423,N_13036,N_14026);
or UO_424 (O_424,N_13779,N_12504);
xnor UO_425 (O_425,N_14335,N_13448);
xor UO_426 (O_426,N_14920,N_12213);
nand UO_427 (O_427,N_14037,N_14483);
and UO_428 (O_428,N_12662,N_12377);
nor UO_429 (O_429,N_12151,N_14132);
or UO_430 (O_430,N_13934,N_12656);
nand UO_431 (O_431,N_14379,N_13368);
nand UO_432 (O_432,N_13256,N_12949);
nor UO_433 (O_433,N_14461,N_12535);
and UO_434 (O_434,N_14703,N_12964);
or UO_435 (O_435,N_14388,N_13057);
nor UO_436 (O_436,N_14656,N_14090);
or UO_437 (O_437,N_14270,N_14775);
nor UO_438 (O_438,N_14880,N_12737);
xor UO_439 (O_439,N_12786,N_14089);
nand UO_440 (O_440,N_14481,N_14586);
nor UO_441 (O_441,N_14800,N_13253);
nor UO_442 (O_442,N_14226,N_14000);
nor UO_443 (O_443,N_14457,N_14876);
xor UO_444 (O_444,N_13961,N_14616);
xor UO_445 (O_445,N_12714,N_13565);
and UO_446 (O_446,N_13542,N_14878);
nand UO_447 (O_447,N_14485,N_14195);
xnor UO_448 (O_448,N_13318,N_14980);
nor UO_449 (O_449,N_13693,N_12093);
xor UO_450 (O_450,N_13898,N_12812);
or UO_451 (O_451,N_13277,N_14271);
xor UO_452 (O_452,N_14242,N_12825);
nand UO_453 (O_453,N_12711,N_12307);
nand UO_454 (O_454,N_14401,N_13663);
nor UO_455 (O_455,N_12593,N_13220);
nand UO_456 (O_456,N_13778,N_12747);
and UO_457 (O_457,N_12481,N_12931);
and UO_458 (O_458,N_12236,N_14353);
or UO_459 (O_459,N_12720,N_12638);
xor UO_460 (O_460,N_13267,N_14590);
and UO_461 (O_461,N_14908,N_12988);
nand UO_462 (O_462,N_14724,N_13548);
xnor UO_463 (O_463,N_14430,N_14087);
nor UO_464 (O_464,N_14534,N_12981);
nor UO_465 (O_465,N_13489,N_14302);
and UO_466 (O_466,N_13004,N_14400);
xnor UO_467 (O_467,N_12373,N_13587);
xor UO_468 (O_468,N_13555,N_14340);
nor UO_469 (O_469,N_14726,N_12362);
and UO_470 (O_470,N_13447,N_13421);
xnor UO_471 (O_471,N_14795,N_12970);
xor UO_472 (O_472,N_12879,N_14411);
nand UO_473 (O_473,N_12936,N_14488);
and UO_474 (O_474,N_13025,N_12044);
and UO_475 (O_475,N_12962,N_14170);
xnor UO_476 (O_476,N_13386,N_12034);
and UO_477 (O_477,N_13102,N_14881);
or UO_478 (O_478,N_13589,N_13302);
nor UO_479 (O_479,N_12632,N_14265);
or UO_480 (O_480,N_12582,N_12275);
and UO_481 (O_481,N_14259,N_12325);
or UO_482 (O_482,N_12614,N_14025);
or UO_483 (O_483,N_14009,N_14657);
nor UO_484 (O_484,N_12098,N_13156);
xnor UO_485 (O_485,N_12900,N_14846);
xnor UO_486 (O_486,N_13746,N_12590);
nand UO_487 (O_487,N_12330,N_14367);
xnor UO_488 (O_488,N_13457,N_13831);
xor UO_489 (O_489,N_12554,N_13139);
nand UO_490 (O_490,N_12445,N_14047);
xnor UO_491 (O_491,N_14263,N_14893);
and UO_492 (O_492,N_14368,N_12396);
or UO_493 (O_493,N_14455,N_12426);
or UO_494 (O_494,N_12976,N_13173);
nor UO_495 (O_495,N_12792,N_12728);
and UO_496 (O_496,N_12803,N_12563);
nand UO_497 (O_497,N_14249,N_12016);
nand UO_498 (O_498,N_14305,N_14327);
or UO_499 (O_499,N_14673,N_12528);
or UO_500 (O_500,N_14733,N_14710);
or UO_501 (O_501,N_12667,N_12316);
or UO_502 (O_502,N_14470,N_13141);
or UO_503 (O_503,N_12804,N_14498);
xor UO_504 (O_504,N_13221,N_12778);
and UO_505 (O_505,N_12137,N_13126);
or UO_506 (O_506,N_13062,N_13391);
xor UO_507 (O_507,N_14567,N_13496);
xor UO_508 (O_508,N_12643,N_12526);
xor UO_509 (O_509,N_12819,N_13424);
nor UO_510 (O_510,N_13306,N_14757);
or UO_511 (O_511,N_13819,N_14559);
or UO_512 (O_512,N_14897,N_13987);
and UO_513 (O_513,N_12284,N_12121);
and UO_514 (O_514,N_14389,N_12478);
and UO_515 (O_515,N_14275,N_12768);
xor UO_516 (O_516,N_13171,N_13791);
and UO_517 (O_517,N_13906,N_14124);
nor UO_518 (O_518,N_12729,N_12536);
or UO_519 (O_519,N_12049,N_13389);
xnor UO_520 (O_520,N_13000,N_14484);
or UO_521 (O_521,N_13164,N_14773);
or UO_522 (O_522,N_14477,N_14900);
nor UO_523 (O_523,N_12969,N_13799);
and UO_524 (O_524,N_14591,N_14171);
nand UO_525 (O_525,N_12384,N_14048);
nand UO_526 (O_526,N_14816,N_13377);
nand UO_527 (O_527,N_13449,N_14636);
nor UO_528 (O_528,N_13925,N_12823);
xor UO_529 (O_529,N_12550,N_13323);
or UO_530 (O_530,N_12665,N_12581);
nor UO_531 (O_531,N_13861,N_13677);
nor UO_532 (O_532,N_13297,N_13708);
nor UO_533 (O_533,N_12344,N_13904);
or UO_534 (O_534,N_12116,N_14595);
and UO_535 (O_535,N_12270,N_14081);
and UO_536 (O_536,N_14738,N_12054);
nor UO_537 (O_537,N_12296,N_13455);
nand UO_538 (O_538,N_13570,N_13279);
nand UO_539 (O_539,N_13958,N_12058);
xnor UO_540 (O_540,N_13858,N_12437);
nand UO_541 (O_541,N_14879,N_13750);
xor UO_542 (O_542,N_12126,N_14814);
or UO_543 (O_543,N_14244,N_12865);
nand UO_544 (O_544,N_12631,N_14134);
nor UO_545 (O_545,N_13131,N_14675);
or UO_546 (O_546,N_13359,N_14972);
xor UO_547 (O_547,N_14019,N_12613);
and UO_548 (O_548,N_14251,N_13668);
and UO_549 (O_549,N_14871,N_12293);
and UO_550 (O_550,N_12543,N_14101);
and UO_551 (O_551,N_13870,N_13381);
nand UO_552 (O_552,N_14020,N_12376);
xor UO_553 (O_553,N_12980,N_13128);
or UO_554 (O_554,N_14898,N_12648);
or UO_555 (O_555,N_12894,N_12532);
xor UO_556 (O_556,N_12724,N_13850);
and UO_557 (O_557,N_13954,N_13458);
and UO_558 (O_558,N_12171,N_12787);
nor UO_559 (O_559,N_13871,N_14494);
nor UO_560 (O_560,N_12096,N_12052);
and UO_561 (O_561,N_12454,N_12273);
xor UO_562 (O_562,N_12605,N_14347);
nor UO_563 (O_563,N_14610,N_12386);
nor UO_564 (O_564,N_13132,N_12406);
nand UO_565 (O_565,N_12240,N_12430);
xor UO_566 (O_566,N_12431,N_13373);
nand UO_567 (O_567,N_13766,N_14568);
or UO_568 (O_568,N_12160,N_13578);
and UO_569 (O_569,N_14224,N_14630);
nor UO_570 (O_570,N_12453,N_13829);
nand UO_571 (O_571,N_14495,N_13658);
nand UO_572 (O_572,N_13055,N_14257);
and UO_573 (O_573,N_14433,N_12594);
xnor UO_574 (O_574,N_14262,N_14824);
xor UO_575 (O_575,N_13543,N_13860);
xor UO_576 (O_576,N_13798,N_12146);
xnor UO_577 (O_577,N_13828,N_13254);
or UO_578 (O_578,N_13930,N_14179);
nand UO_579 (O_579,N_12715,N_13051);
xor UO_580 (O_580,N_13390,N_14803);
or UO_581 (O_581,N_14531,N_14414);
nand UO_582 (O_582,N_14776,N_13545);
nand UO_583 (O_583,N_13938,N_14609);
nor UO_584 (O_584,N_14947,N_13560);
and UO_585 (O_585,N_13271,N_14035);
nor UO_586 (O_586,N_12814,N_14713);
xor UO_587 (O_587,N_14186,N_12328);
nor UO_588 (O_588,N_14312,N_13669);
nand UO_589 (O_589,N_12670,N_12482);
nand UO_590 (O_590,N_12655,N_13725);
nand UO_591 (O_591,N_13395,N_12017);
nor UO_592 (O_592,N_13718,N_14031);
xnor UO_593 (O_593,N_14700,N_14973);
nand UO_594 (O_594,N_12351,N_12982);
nand UO_595 (O_595,N_13899,N_14866);
nor UO_596 (O_596,N_12868,N_13837);
and UO_597 (O_597,N_13997,N_13161);
and UO_598 (O_598,N_12959,N_14003);
nor UO_599 (O_599,N_13157,N_12132);
nand UO_600 (O_600,N_12388,N_13697);
nor UO_601 (O_601,N_14113,N_14873);
nand UO_602 (O_602,N_13186,N_14734);
or UO_603 (O_603,N_14372,N_12047);
nor UO_604 (O_604,N_13595,N_14632);
xnor UO_605 (O_605,N_14398,N_12070);
nand UO_606 (O_606,N_14918,N_13326);
xor UO_607 (O_607,N_12802,N_13882);
xnor UO_608 (O_608,N_14665,N_13069);
nor UO_609 (O_609,N_13361,N_13845);
and UO_610 (O_610,N_13258,N_12617);
or UO_611 (O_611,N_14215,N_12789);
nor UO_612 (O_612,N_12767,N_13274);
and UO_613 (O_613,N_12060,N_13399);
xnor UO_614 (O_614,N_13265,N_12465);
nand UO_615 (O_615,N_12785,N_13217);
nor UO_616 (O_616,N_14626,N_14892);
nor UO_617 (O_617,N_13228,N_12584);
or UO_618 (O_618,N_12731,N_13234);
and UO_619 (O_619,N_12688,N_14949);
xor UO_620 (O_620,N_14987,N_12231);
and UO_621 (O_621,N_14570,N_13313);
or UO_622 (O_622,N_14100,N_13872);
xor UO_623 (O_623,N_14663,N_14296);
nor UO_624 (O_624,N_14549,N_12722);
xor UO_625 (O_625,N_13081,N_14909);
and UO_626 (O_626,N_12534,N_14188);
and UO_627 (O_627,N_14221,N_13088);
nand UO_628 (O_628,N_13190,N_12294);
nand UO_629 (O_629,N_12644,N_13752);
nand UO_630 (O_630,N_13347,N_14766);
xnor UO_631 (O_631,N_14562,N_12822);
nor UO_632 (O_632,N_14279,N_13178);
and UO_633 (O_633,N_13034,N_14712);
xnor UO_634 (O_634,N_13408,N_12474);
or UO_635 (O_635,N_13012,N_13994);
and UO_636 (O_636,N_14243,N_14030);
nor UO_637 (O_637,N_14306,N_12681);
xor UO_638 (O_638,N_13396,N_12371);
nor UO_639 (O_639,N_14552,N_12875);
xor UO_640 (O_640,N_14152,N_13108);
xor UO_641 (O_641,N_12914,N_14601);
and UO_642 (O_642,N_14588,N_12429);
nor UO_643 (O_643,N_13849,N_12952);
and UO_644 (O_644,N_13376,N_14841);
and UO_645 (O_645,N_14965,N_14915);
or UO_646 (O_646,N_13461,N_14278);
or UO_647 (O_647,N_12346,N_12260);
nand UO_648 (O_648,N_13078,N_13285);
nor UO_649 (O_649,N_12902,N_13241);
or UO_650 (O_650,N_14323,N_12110);
xor UO_651 (O_651,N_14059,N_14480);
and UO_652 (O_652,N_12705,N_14288);
xnor UO_653 (O_653,N_13027,N_12304);
or UO_654 (O_654,N_13619,N_14849);
nor UO_655 (O_655,N_13079,N_14266);
nand UO_656 (O_656,N_13339,N_14612);
xnor UO_657 (O_657,N_12283,N_13610);
nand UO_658 (O_658,N_12589,N_13887);
nor UO_659 (O_659,N_13730,N_12324);
xnor UO_660 (O_660,N_13497,N_13524);
xor UO_661 (O_661,N_12837,N_12544);
nand UO_662 (O_662,N_13706,N_12091);
nor UO_663 (O_663,N_12579,N_12727);
nand UO_664 (O_664,N_12011,N_13470);
nand UO_665 (O_665,N_13223,N_12157);
xnor UO_666 (O_666,N_13728,N_14708);
xor UO_667 (O_667,N_14068,N_13885);
nor UO_668 (O_668,N_14982,N_12668);
nand UO_669 (O_669,N_12869,N_13175);
and UO_670 (O_670,N_13742,N_12383);
or UO_671 (O_671,N_14686,N_13029);
nor UO_672 (O_672,N_14659,N_14553);
or UO_673 (O_673,N_13193,N_14150);
nand UO_674 (O_674,N_14997,N_12150);
or UO_675 (O_675,N_13483,N_14217);
and UO_676 (O_676,N_12004,N_14886);
nand UO_677 (O_677,N_14002,N_12412);
or UO_678 (O_678,N_13694,N_13745);
and UO_679 (O_679,N_14996,N_12596);
and UO_680 (O_680,N_13559,N_14487);
and UO_681 (O_681,N_12218,N_12891);
xor UO_682 (O_682,N_13015,N_14577);
xnor UO_683 (O_683,N_14974,N_12198);
or UO_684 (O_684,N_14790,N_13488);
nand UO_685 (O_685,N_14473,N_13196);
and UO_686 (O_686,N_14268,N_12399);
nand UO_687 (O_687,N_13760,N_14719);
xnor UO_688 (O_688,N_12928,N_12564);
xor UO_689 (O_689,N_14308,N_13992);
and UO_690 (O_690,N_13696,N_14313);
and UO_691 (O_691,N_14865,N_12692);
nand UO_692 (O_692,N_13823,N_12718);
xor UO_693 (O_693,N_13300,N_13003);
and UO_694 (O_694,N_13093,N_12249);
or UO_695 (O_695,N_13054,N_13181);
xor UO_696 (O_696,N_13815,N_13142);
or UO_697 (O_697,N_14735,N_12055);
and UO_698 (O_698,N_12571,N_13946);
nor UO_699 (O_699,N_12253,N_14192);
and UO_700 (O_700,N_14040,N_14840);
and UO_701 (O_701,N_13843,N_14923);
or UO_702 (O_702,N_13591,N_12698);
xor UO_703 (O_703,N_12633,N_14797);
nor UO_704 (O_704,N_14593,N_12695);
and UO_705 (O_705,N_13605,N_13350);
or UO_706 (O_706,N_13965,N_13514);
or UO_707 (O_707,N_13583,N_13446);
nor UO_708 (O_708,N_12629,N_13664);
xnor UO_709 (O_709,N_12977,N_13439);
nand UO_710 (O_710,N_14084,N_13859);
and UO_711 (O_711,N_12063,N_14819);
nand UO_712 (O_712,N_14165,N_14053);
or UO_713 (O_713,N_14756,N_13531);
nand UO_714 (O_714,N_14023,N_14073);
and UO_715 (O_715,N_12555,N_12155);
or UO_716 (O_716,N_13198,N_14916);
nand UO_717 (O_717,N_14223,N_13324);
xnor UO_718 (O_718,N_13426,N_12998);
nand UO_719 (O_719,N_14576,N_12201);
nor UO_720 (O_720,N_13356,N_14143);
nand UO_721 (O_721,N_13932,N_13037);
or UO_722 (O_722,N_13219,N_12824);
and UO_723 (O_723,N_13257,N_13795);
nand UO_724 (O_724,N_12408,N_14569);
nand UO_725 (O_725,N_14228,N_13289);
nand UO_726 (O_726,N_12033,N_13264);
nand UO_727 (O_727,N_12857,N_13335);
and UO_728 (O_728,N_13520,N_12784);
or UO_729 (O_729,N_13121,N_13374);
or UO_730 (O_730,N_12569,N_13814);
nand UO_731 (O_731,N_13824,N_12336);
xor UO_732 (O_732,N_12780,N_13509);
or UO_733 (O_733,N_14661,N_12925);
nand UO_734 (O_734,N_13235,N_14301);
or UO_735 (O_735,N_12858,N_13623);
or UO_736 (O_736,N_12831,N_14339);
and UO_737 (O_737,N_12795,N_14922);
nor UO_738 (O_738,N_12682,N_14863);
nor UO_739 (O_739,N_12145,N_12774);
or UO_740 (O_740,N_13655,N_14830);
nand UO_741 (O_741,N_13603,N_13043);
nand UO_742 (O_742,N_13048,N_13500);
or UO_743 (O_743,N_12966,N_13626);
xor UO_744 (O_744,N_12434,N_14747);
and UO_745 (O_745,N_14730,N_14767);
xnor UO_746 (O_746,N_13144,N_12753);
nand UO_747 (O_747,N_13280,N_12420);
and UO_748 (O_748,N_14761,N_12983);
nor UO_749 (O_749,N_12239,N_13636);
nand UO_750 (O_750,N_14706,N_13864);
and UO_751 (O_751,N_13400,N_13996);
and UO_752 (O_752,N_13369,N_14720);
nor UO_753 (O_753,N_13659,N_13435);
or UO_754 (O_754,N_13466,N_12241);
xor UO_755 (O_755,N_14001,N_14753);
and UO_756 (O_756,N_12347,N_12520);
or UO_757 (O_757,N_13499,N_14823);
nor UO_758 (O_758,N_14311,N_13291);
xnor UO_759 (O_759,N_14419,N_12212);
nand UO_760 (O_760,N_14558,N_14475);
xor UO_761 (O_761,N_13516,N_12469);
nand UO_762 (O_762,N_12965,N_13844);
or UO_763 (O_763,N_14822,N_14458);
or UO_764 (O_764,N_13721,N_14022);
nand UO_765 (O_765,N_12880,N_14759);
nand UO_766 (O_766,N_14545,N_12009);
and UO_767 (O_767,N_14365,N_12961);
nand UO_768 (O_768,N_12599,N_12525);
nor UO_769 (O_769,N_13903,N_14254);
xor UO_770 (O_770,N_13743,N_12677);
nand UO_771 (O_771,N_13939,N_12053);
or UO_772 (O_772,N_13259,N_12140);
nor UO_773 (O_773,N_14163,N_13880);
and UO_774 (O_774,N_13273,N_14036);
nand UO_775 (O_775,N_13661,N_14635);
or UO_776 (O_776,N_12205,N_12282);
and UO_777 (O_777,N_14137,N_14782);
or UO_778 (O_778,N_12143,N_12507);
and UO_779 (O_779,N_13309,N_13645);
or UO_780 (O_780,N_13662,N_14732);
or UO_781 (O_781,N_14012,N_13767);
nand UO_782 (O_782,N_12932,N_13427);
xnor UO_783 (O_783,N_12172,N_12923);
xor UO_784 (O_784,N_13331,N_13660);
and UO_785 (O_785,N_12783,N_13505);
nand UO_786 (O_786,N_12773,N_14496);
xnor UO_787 (O_787,N_14784,N_13371);
nor UO_788 (O_788,N_12442,N_14373);
nand UO_789 (O_789,N_14924,N_13649);
nand UO_790 (O_790,N_14060,N_13208);
nand UO_791 (O_791,N_12842,N_13674);
nor UO_792 (O_792,N_14459,N_14981);
nand UO_793 (O_793,N_12838,N_13203);
xor UO_794 (O_794,N_14141,N_13050);
nor UO_795 (O_795,N_13184,N_12100);
xor UO_796 (O_796,N_12174,N_14158);
or UO_797 (O_797,N_12735,N_12073);
or UO_798 (O_798,N_14872,N_13098);
nor UO_799 (O_799,N_13409,N_13366);
and UO_800 (O_800,N_12128,N_12801);
xor UO_801 (O_801,N_14617,N_14261);
or UO_802 (O_802,N_12200,N_12006);
nor UO_803 (O_803,N_14471,N_14176);
xor UO_804 (O_804,N_14582,N_14250);
and UO_805 (O_805,N_14796,N_13995);
or UO_806 (O_806,N_13314,N_12007);
nor UO_807 (O_807,N_12037,N_12487);
nor UO_808 (O_808,N_13787,N_13653);
nand UO_809 (O_809,N_12298,N_14901);
nor UO_810 (O_810,N_12153,N_14606);
nor UO_811 (O_811,N_13616,N_12790);
or UO_812 (O_812,N_13681,N_12807);
and UO_813 (O_813,N_14937,N_13322);
or UO_814 (O_814,N_12845,N_13544);
or UO_815 (O_815,N_13977,N_12559);
and UO_816 (O_816,N_13557,N_13847);
nand UO_817 (O_817,N_12944,N_12092);
nor UO_818 (O_818,N_12379,N_13310);
or UO_819 (O_819,N_12106,N_12933);
nand UO_820 (O_820,N_12152,N_13754);
xnor UO_821 (O_821,N_12913,N_13741);
nand UO_822 (O_822,N_12109,N_13363);
nand UO_823 (O_823,N_13701,N_12015);
and UO_824 (O_824,N_12335,N_13940);
xnor UO_825 (O_825,N_14788,N_14189);
nor UO_826 (O_826,N_14855,N_13820);
or UO_827 (O_827,N_13515,N_12553);
nor UO_828 (O_828,N_12759,N_13099);
or UO_829 (O_829,N_14467,N_14524);
or UO_830 (O_830,N_14679,N_12637);
xnor UO_831 (O_831,N_13387,N_14671);
xor UO_832 (O_832,N_12129,N_14933);
xor UO_833 (O_833,N_13567,N_13993);
and UO_834 (O_834,N_13268,N_13912);
and UO_835 (O_835,N_12700,N_13969);
and UO_836 (O_836,N_12628,N_14643);
xor UO_837 (O_837,N_12586,N_14572);
or UO_838 (O_838,N_12123,N_14104);
nor UO_839 (O_839,N_13666,N_14868);
nand UO_840 (O_840,N_12649,N_13782);
nor UO_841 (O_841,N_12266,N_13020);
nand UO_842 (O_842,N_12694,N_13284);
nand UO_843 (O_843,N_14875,N_13900);
and UO_844 (O_844,N_12323,N_12023);
xnor UO_845 (O_845,N_14780,N_12461);
and UO_846 (O_846,N_12575,N_14754);
and UO_847 (O_847,N_13877,N_12623);
nor UO_848 (O_848,N_13246,N_13478);
xnor UO_849 (O_849,N_14787,N_13460);
and UO_850 (O_850,N_14725,N_13442);
or UO_851 (O_851,N_13809,N_14366);
and UO_852 (O_852,N_14114,N_14940);
nand UO_853 (O_853,N_12300,N_14130);
nor UO_854 (O_854,N_12888,N_14765);
and UO_855 (O_855,N_14157,N_12881);
nand UO_856 (O_856,N_12269,N_14164);
or UO_857 (O_857,N_12585,N_14109);
or UO_858 (O_858,N_14127,N_12686);
nand UO_859 (O_859,N_12626,N_14504);
xor UO_860 (O_860,N_12946,N_12835);
and UO_861 (O_861,N_14051,N_14984);
or UO_862 (O_862,N_14303,N_12187);
or UO_863 (O_863,N_13564,N_14013);
nand UO_864 (O_864,N_13179,N_13174);
xnor UO_865 (O_865,N_12222,N_13709);
and UO_866 (O_866,N_13719,N_13773);
or UO_867 (O_867,N_12972,N_14739);
nor UO_868 (O_868,N_12443,N_12188);
nor UO_869 (O_869,N_14131,N_14427);
nand UO_870 (O_870,N_14537,N_13836);
or UO_871 (O_871,N_13109,N_13519);
or UO_872 (O_872,N_13644,N_12338);
and UO_873 (O_873,N_12181,N_13260);
nor UO_874 (O_874,N_12618,N_12954);
or UO_875 (O_875,N_14755,N_14095);
or UO_876 (O_876,N_13021,N_12463);
or UO_877 (O_877,N_14086,N_12342);
xnor UO_878 (O_878,N_13740,N_13493);
and UO_879 (O_879,N_13576,N_14696);
nand UO_880 (O_880,N_12855,N_13618);
or UO_881 (O_881,N_13656,N_12861);
nor UO_882 (O_882,N_13334,N_12428);
xnor UO_883 (O_883,N_13953,N_14284);
xnor UO_884 (O_884,N_14056,N_14283);
xor UO_885 (O_885,N_12573,N_13902);
and UO_886 (O_886,N_14160,N_13011);
nand UO_887 (O_887,N_12107,N_12102);
or UO_888 (O_888,N_12248,N_13444);
nor UO_889 (O_889,N_14421,N_13269);
nor UO_890 (O_890,N_14370,N_12777);
and UO_891 (O_891,N_14896,N_12115);
and UO_892 (O_892,N_13068,N_13229);
nand UO_893 (O_893,N_12272,N_14533);
nand UO_894 (O_894,N_12158,N_13671);
and UO_895 (O_895,N_14453,N_12533);
xor UO_896 (O_896,N_14193,N_14805);
or UO_897 (O_897,N_14377,N_13100);
xnor UO_898 (O_898,N_14662,N_13286);
nor UO_899 (O_899,N_14548,N_14395);
nand UO_900 (O_900,N_13586,N_12542);
xor UO_901 (O_901,N_14835,N_13278);
nand UO_902 (O_902,N_13905,N_13597);
nor UO_903 (O_903,N_12863,N_12237);
or UO_904 (O_904,N_14126,N_13834);
nand UO_905 (O_905,N_12927,N_12167);
nor UO_906 (O_906,N_12361,N_13379);
and UO_907 (O_907,N_14502,N_14948);
nor UO_908 (O_908,N_14977,N_13945);
nand UO_909 (O_909,N_13315,N_12072);
or UO_910 (O_910,N_14869,N_14378);
xnor UO_911 (O_911,N_12986,N_13955);
or UO_912 (O_912,N_14971,N_14622);
or UO_913 (O_913,N_12739,N_13120);
nor UO_914 (O_914,N_13927,N_13875);
nand UO_915 (O_915,N_14107,N_12893);
or UO_916 (O_916,N_12721,N_12370);
xnor UO_917 (O_917,N_14269,N_13437);
nand UO_918 (O_918,N_13622,N_12566);
nor UO_919 (O_919,N_14070,N_12135);
nor UO_920 (O_920,N_13422,N_13477);
and UO_921 (O_921,N_13598,N_14862);
xnor UO_922 (O_922,N_13452,N_13686);
nand UO_923 (O_923,N_12941,N_13002);
and UO_924 (O_924,N_12994,N_14934);
xor UO_925 (O_925,N_12130,N_14154);
xor UO_926 (O_926,N_12968,N_14911);
nand UO_927 (O_927,N_14978,N_13191);
xnor UO_928 (O_928,N_14350,N_12852);
nor UO_929 (O_929,N_13884,N_14813);
and UO_930 (O_930,N_14196,N_14538);
nand UO_931 (O_931,N_13988,N_13352);
and UO_932 (O_932,N_13687,N_12297);
nand UO_933 (O_933,N_12280,N_14325);
xor UO_934 (O_934,N_13392,N_14364);
or UO_935 (O_935,N_14282,N_13287);
or UO_936 (O_936,N_14540,N_12214);
xor UO_937 (O_937,N_14769,N_13205);
and UO_938 (O_938,N_12359,N_14298);
or UO_939 (O_939,N_12653,N_12938);
and UO_940 (O_940,N_14178,N_13998);
xor UO_941 (O_941,N_13479,N_14921);
nand UO_942 (O_942,N_14817,N_12274);
or UO_943 (O_943,N_14953,N_12864);
nor UO_944 (O_944,N_13640,N_14793);
and UO_945 (O_945,N_13865,N_13957);
nand UO_946 (O_946,N_14928,N_14281);
nor UO_947 (O_947,N_13985,N_14054);
and UO_948 (O_948,N_14930,N_14512);
and UO_949 (O_949,N_14063,N_13690);
nand UO_950 (O_950,N_12473,N_12084);
xor UO_951 (O_951,N_12077,N_12210);
nor UO_952 (O_952,N_14585,N_14437);
and UO_953 (O_953,N_14080,N_12353);
xnor UO_954 (O_954,N_14203,N_13759);
nand UO_955 (O_955,N_12496,N_12509);
and UO_956 (O_956,N_12407,N_13890);
nand UO_957 (O_957,N_13232,N_12233);
nor UO_958 (O_958,N_13962,N_13761);
or UO_959 (O_959,N_12436,N_12652);
or UO_960 (O_960,N_13964,N_12247);
and UO_961 (O_961,N_12971,N_14667);
and UO_962 (O_962,N_13255,N_12910);
nor UO_963 (O_963,N_13568,N_14655);
nor UO_964 (O_964,N_13136,N_13372);
nand UO_965 (O_965,N_12224,N_13215);
and UO_966 (O_966,N_14231,N_12609);
and UO_967 (O_967,N_13341,N_13463);
or UO_968 (O_968,N_12493,N_14843);
nor UO_969 (O_969,N_13966,N_14681);
xnor UO_970 (O_970,N_13774,N_12354);
xor UO_971 (O_971,N_14277,N_13888);
and UO_972 (O_972,N_14151,N_12424);
and UO_973 (O_973,N_13360,N_14381);
nor UO_974 (O_974,N_12658,N_13840);
and UO_975 (O_975,N_14116,N_12840);
nor UO_976 (O_976,N_13183,N_13584);
or UO_977 (O_977,N_13913,N_14985);
nand UO_978 (O_978,N_13551,N_13243);
xor UO_979 (O_979,N_14329,N_12134);
nor UO_980 (O_980,N_12956,N_14161);
and UO_981 (O_981,N_12742,N_14718);
and UO_982 (O_982,N_12678,N_12693);
and UO_983 (O_983,N_14676,N_13960);
nor UO_984 (O_984,N_14685,N_14836);
or UO_985 (O_985,N_13495,N_14516);
xor UO_986 (O_986,N_13080,N_14383);
and UO_987 (O_987,N_12769,N_13534);
and UO_988 (O_988,N_12265,N_13398);
nor UO_989 (O_989,N_13087,N_13262);
nand UO_990 (O_990,N_13615,N_13506);
and UO_991 (O_991,N_14891,N_14812);
xnor UO_992 (O_992,N_12760,N_13160);
nand UO_993 (O_993,N_14749,N_12508);
and UO_994 (O_994,N_13434,N_13633);
and UO_995 (O_995,N_14055,N_13009);
nor UO_996 (O_996,N_14515,N_14065);
or UO_997 (O_997,N_12175,N_14917);
and UO_998 (O_998,N_12089,N_12045);
or UO_999 (O_999,N_13785,N_12934);
xor UO_1000 (O_1000,N_12886,N_13528);
nor UO_1001 (O_1001,N_12138,N_14519);
nor UO_1002 (O_1002,N_13707,N_12611);
xnor UO_1003 (O_1003,N_12416,N_14331);
nand UO_1004 (O_1004,N_14695,N_12612);
nand UO_1005 (O_1005,N_12464,N_14253);
and UO_1006 (O_1006,N_12026,N_13303);
or UO_1007 (O_1007,N_12400,N_13713);
and UO_1008 (O_1008,N_14380,N_14652);
xor UO_1009 (O_1009,N_14600,N_14017);
or UO_1010 (O_1010,N_14699,N_12659);
xor UO_1011 (O_1011,N_12531,N_14125);
xnor UO_1012 (O_1012,N_12375,N_12027);
xnor UO_1013 (O_1013,N_14213,N_12529);
and UO_1014 (O_1014,N_14280,N_13436);
nand UO_1015 (O_1015,N_14999,N_14008);
nor UO_1016 (O_1016,N_13143,N_14208);
or UO_1017 (O_1017,N_12031,N_14505);
nor UO_1018 (O_1018,N_12148,N_13060);
and UO_1019 (O_1019,N_14448,N_14027);
or UO_1020 (O_1020,N_13307,N_12349);
or UO_1021 (O_1021,N_13606,N_14123);
and UO_1022 (O_1022,N_12716,N_13430);
or UO_1023 (O_1023,N_12758,N_14273);
nor UO_1024 (O_1024,N_13047,N_13167);
nor UO_1025 (O_1025,N_13281,N_12568);
xor UO_1026 (O_1026,N_13744,N_13035);
xnor UO_1027 (O_1027,N_13240,N_13675);
nor UO_1028 (O_1028,N_14062,N_12622);
xnor UO_1029 (O_1029,N_13135,N_12833);
nor UO_1030 (O_1030,N_12514,N_14299);
nand UO_1031 (O_1031,N_14651,N_14716);
nor UO_1032 (O_1032,N_13365,N_14384);
xnor UO_1033 (O_1033,N_14256,N_13827);
nand UO_1034 (O_1034,N_13582,N_12259);
xnor UO_1035 (O_1035,N_12290,N_14220);
nor UO_1036 (O_1036,N_13296,N_12395);
nand UO_1037 (O_1037,N_14159,N_13971);
or UO_1038 (O_1038,N_12839,N_12450);
xnor UO_1039 (O_1039,N_14491,N_14991);
or UO_1040 (O_1040,N_12821,N_14351);
or UO_1041 (O_1041,N_13066,N_12117);
and UO_1042 (O_1042,N_13807,N_14233);
nand UO_1043 (O_1043,N_12672,N_13230);
xnor UO_1044 (O_1044,N_14509,N_12746);
nor UO_1045 (O_1045,N_12940,N_14970);
and UO_1046 (O_1046,N_14451,N_12661);
nor UO_1047 (O_1047,N_14391,N_12603);
and UO_1048 (O_1048,N_13076,N_13045);
and UO_1049 (O_1049,N_14291,N_14644);
nor UO_1050 (O_1050,N_12360,N_12101);
nand UO_1051 (O_1051,N_14806,N_13148);
or UO_1052 (O_1052,N_13358,N_12041);
nand UO_1053 (O_1053,N_12703,N_13911);
nor UO_1054 (O_1054,N_12235,N_12793);
nor UO_1055 (O_1055,N_14450,N_13346);
or UO_1056 (O_1056,N_12808,N_12267);
nor UO_1057 (O_1057,N_12334,N_12851);
nor UO_1058 (O_1058,N_13299,N_12419);
nor UO_1059 (O_1059,N_14167,N_14884);
xor UO_1060 (O_1060,N_14860,N_12899);
nand UO_1061 (O_1061,N_12415,N_14598);
nor UO_1062 (O_1062,N_14004,N_12403);
xor UO_1063 (O_1063,N_12854,N_13732);
nor UO_1064 (O_1064,N_14854,N_12243);
xnor UO_1065 (O_1065,N_14607,N_14386);
or UO_1066 (O_1066,N_14010,N_13211);
xor UO_1067 (O_1067,N_14511,N_12595);
nand UO_1068 (O_1068,N_13720,N_12358);
xnor UO_1069 (O_1069,N_12957,N_12221);
or UO_1070 (O_1070,N_12572,N_12882);
and UO_1071 (O_1071,N_13797,N_13129);
or UO_1072 (O_1072,N_14525,N_12019);
or UO_1073 (O_1073,N_12975,N_14041);
nor UO_1074 (O_1074,N_14145,N_14434);
and UO_1075 (O_1075,N_12922,N_14639);
and UO_1076 (O_1076,N_12484,N_14779);
or UO_1077 (O_1077,N_12877,N_13922);
xnor UO_1078 (O_1078,N_14286,N_13158);
xor UO_1079 (O_1079,N_12872,N_14407);
nor UO_1080 (O_1080,N_13848,N_12276);
xor UO_1081 (O_1081,N_13085,N_12483);
nand UO_1082 (O_1082,N_13008,N_14392);
or UO_1083 (O_1083,N_13119,N_14583);
nor UO_1084 (O_1084,N_13115,N_13031);
and UO_1085 (O_1085,N_13394,N_14833);
xnor UO_1086 (O_1086,N_14236,N_14191);
nor UO_1087 (O_1087,N_14246,N_14760);
and UO_1088 (O_1088,N_12984,N_13793);
or UO_1089 (O_1089,N_12892,N_14472);
nor UO_1090 (O_1090,N_12185,N_13338);
xnor UO_1091 (O_1091,N_13165,N_14925);
xnor UO_1092 (O_1092,N_13635,N_13577);
nand UO_1093 (O_1093,N_14204,N_12890);
xnor UO_1094 (O_1094,N_13152,N_13052);
xnor UO_1095 (O_1095,N_13563,N_13433);
xor UO_1096 (O_1096,N_12859,N_14285);
or UO_1097 (O_1097,N_13486,N_14919);
nor UO_1098 (O_1098,N_13261,N_14046);
nor UO_1099 (O_1099,N_14510,N_14018);
or UO_1100 (O_1100,N_12500,N_13780);
xnor UO_1101 (O_1101,N_14740,N_12867);
xnor UO_1102 (O_1102,N_13916,N_14589);
nand UO_1103 (O_1103,N_14856,N_14687);
or UO_1104 (O_1104,N_14647,N_14573);
nor UO_1105 (O_1105,N_14728,N_12878);
and UO_1106 (O_1106,N_14561,N_14913);
nor UO_1107 (O_1107,N_13609,N_13862);
nand UO_1108 (O_1108,N_13304,N_12565);
nor UO_1109 (O_1109,N_13832,N_14969);
xnor UO_1110 (O_1110,N_12183,N_12616);
nand UO_1111 (O_1111,N_14682,N_12432);
and UO_1112 (O_1112,N_13406,N_12577);
and UO_1113 (O_1113,N_13569,N_12466);
nor UO_1114 (O_1114,N_13948,N_13468);
xor UO_1115 (O_1115,N_13657,N_12382);
or UO_1116 (O_1116,N_13006,N_12730);
and UO_1117 (O_1117,N_13189,N_12876);
nor UO_1118 (O_1118,N_14422,N_13293);
and UO_1119 (O_1119,N_12641,N_14852);
nand UO_1120 (O_1120,N_14006,N_12350);
nand UO_1121 (O_1121,N_12515,N_13404);
nand UO_1122 (O_1122,N_14149,N_12271);
nor UO_1123 (O_1123,N_14684,N_12690);
or UO_1124 (O_1124,N_12924,N_12578);
and UO_1125 (O_1125,N_12657,N_13889);
and UO_1126 (O_1126,N_14736,N_12664);
nand UO_1127 (O_1127,N_13676,N_12410);
xor UO_1128 (O_1128,N_13731,N_12000);
nand UO_1129 (O_1129,N_12919,N_14894);
xnor UO_1130 (O_1130,N_12261,N_14121);
or UO_1131 (O_1131,N_14594,N_14772);
xnor UO_1132 (O_1132,N_14697,N_12252);
nor UO_1133 (O_1133,N_13382,N_13522);
xor UO_1134 (O_1134,N_14043,N_12433);
and UO_1135 (O_1135,N_12906,N_12710);
or UO_1136 (O_1136,N_14096,N_13838);
xnor UO_1137 (O_1137,N_13924,N_13751);
xnor UO_1138 (O_1138,N_13692,N_14777);
or UO_1139 (O_1139,N_14021,N_14183);
xnor UO_1140 (O_1140,N_13340,N_13917);
or UO_1141 (O_1141,N_12081,N_14034);
or UO_1142 (O_1142,N_13007,N_13238);
and UO_1143 (O_1143,N_14409,N_14435);
and UO_1144 (O_1144,N_12939,N_12035);
and UO_1145 (O_1145,N_14574,N_13145);
nand UO_1146 (O_1146,N_13682,N_12295);
or UO_1147 (O_1147,N_13883,N_13063);
or UO_1148 (O_1148,N_14098,N_12113);
xor UO_1149 (O_1149,N_13059,N_12435);
and UO_1150 (O_1150,N_13308,N_12050);
xnor UO_1151 (O_1151,N_14834,N_12303);
nor UO_1152 (O_1152,N_12159,N_12097);
nand UO_1153 (O_1153,N_14014,N_14177);
nand UO_1154 (O_1154,N_14486,N_12255);
or UO_1155 (O_1155,N_14057,N_14701);
or UO_1156 (O_1156,N_12401,N_14328);
xor UO_1157 (O_1157,N_14828,N_14818);
nand UO_1158 (O_1158,N_13432,N_12311);
nor UO_1159 (O_1159,N_12133,N_12847);
and UO_1160 (O_1160,N_13579,N_13453);
xor UO_1161 (O_1161,N_12883,N_12799);
and UO_1162 (O_1162,N_13518,N_12909);
nand UO_1163 (O_1163,N_14615,N_12903);
nand UO_1164 (O_1164,N_13976,N_12763);
or UO_1165 (O_1165,N_12776,N_13781);
or UO_1166 (O_1166,N_14355,N_14990);
nor UO_1167 (O_1167,N_13947,N_12154);
nor UO_1168 (O_1168,N_12513,N_12340);
xnor UO_1169 (O_1169,N_14142,N_13928);
and UO_1170 (O_1170,N_14492,N_14770);
and UO_1171 (O_1171,N_12288,N_12828);
or UO_1172 (O_1172,N_12139,N_14532);
xnor UO_1173 (O_1173,N_13117,N_12660);
nand UO_1174 (O_1174,N_13249,N_14359);
and UO_1175 (O_1175,N_14420,N_13979);
or UO_1176 (O_1176,N_14529,N_12229);
and UO_1177 (O_1177,N_12918,N_13768);
nor UO_1178 (O_1178,N_12505,N_13652);
and UO_1179 (O_1179,N_13762,N_14028);
or UO_1180 (O_1180,N_12712,N_12193);
or UO_1181 (O_1181,N_14210,N_14670);
and UO_1182 (O_1182,N_14941,N_14633);
xnor UO_1183 (O_1183,N_13147,N_12144);
or UO_1184 (O_1184,N_14362,N_13517);
nand UO_1185 (O_1185,N_13537,N_14792);
and UO_1186 (O_1186,N_12844,N_12409);
and UO_1187 (O_1187,N_13018,N_12447);
xnor UO_1188 (O_1188,N_13822,N_13915);
nor UO_1189 (O_1189,N_13588,N_12663);
xnor UO_1190 (O_1190,N_13471,N_14111);
nor UO_1191 (O_1191,N_12389,N_13410);
or UO_1192 (O_1192,N_13026,N_12057);
xor UO_1193 (O_1193,N_14274,N_12996);
xnor UO_1194 (O_1194,N_12640,N_14861);
nand UO_1195 (O_1195,N_13485,N_14936);
or UO_1196 (O_1196,N_12195,N_12997);
nor UO_1197 (O_1197,N_12460,N_12489);
nor UO_1198 (O_1198,N_13125,N_14408);
and UO_1199 (O_1199,N_12451,N_13527);
and UO_1200 (O_1200,N_12517,N_14789);
nand UO_1201 (O_1201,N_13975,N_12506);
xor UO_1202 (O_1202,N_12756,N_14225);
xnor UO_1203 (O_1203,N_14029,N_12333);
and UO_1204 (O_1204,N_14649,N_13044);
xnor UO_1205 (O_1205,N_13187,N_14264);
or UO_1206 (O_1206,N_12741,N_13070);
and UO_1207 (O_1207,N_12088,N_13154);
nor UO_1208 (O_1208,N_13614,N_12830);
xnor UO_1209 (O_1209,N_12929,N_13650);
nor UO_1210 (O_1210,N_13248,N_13878);
or UO_1211 (O_1211,N_12189,N_14432);
and UO_1212 (O_1212,N_13978,N_13202);
xnor UO_1213 (O_1213,N_12028,N_14518);
nor UO_1214 (O_1214,N_14182,N_13077);
nand UO_1215 (O_1215,N_12958,N_12226);
nand UO_1216 (O_1216,N_13177,N_14227);
nor UO_1217 (O_1217,N_13695,N_14295);
nor UO_1218 (O_1218,N_12979,N_14848);
xor UO_1219 (O_1219,N_13084,N_14743);
and UO_1220 (O_1220,N_12751,N_14482);
nand UO_1221 (O_1221,N_12164,N_14076);
and UO_1222 (O_1222,N_14831,N_14162);
nor UO_1223 (O_1223,N_14750,N_14680);
and UO_1224 (O_1224,N_12263,N_14929);
xor UO_1225 (O_1225,N_14688,N_13919);
or UO_1226 (O_1226,N_14927,N_14252);
nand UO_1227 (O_1227,N_14705,N_12470);
nor UO_1228 (O_1228,N_13233,N_13038);
nor UO_1229 (O_1229,N_14702,N_12527);
xnor UO_1230 (O_1230,N_13197,N_13868);
nand UO_1231 (O_1231,N_14715,N_14071);
or UO_1232 (O_1232,N_12601,N_14808);
xnor UO_1233 (O_1233,N_14345,N_12365);
nand UO_1234 (O_1234,N_14314,N_12331);
nor UO_1235 (O_1235,N_12798,N_12264);
nand UO_1236 (O_1236,N_12374,N_14956);
xnor UO_1237 (O_1237,N_12170,N_13384);
or UO_1238 (O_1238,N_13967,N_12394);
nor UO_1239 (O_1239,N_12950,N_12850);
or UO_1240 (O_1240,N_12510,N_12291);
nand UO_1241 (O_1241,N_14683,N_12177);
or UO_1242 (O_1242,N_12597,N_12826);
nand UO_1243 (O_1243,N_13602,N_13333);
and UO_1244 (O_1244,N_13195,N_13451);
and UO_1245 (O_1245,N_12494,N_12530);
nor UO_1246 (O_1246,N_12676,N_13481);
nand UO_1247 (O_1247,N_14140,N_12190);
nor UO_1248 (O_1248,N_12363,N_14825);
xor UO_1249 (O_1249,N_12456,N_14899);
xor UO_1250 (O_1250,N_13943,N_12717);
or UO_1251 (O_1251,N_12018,N_12960);
or UO_1252 (O_1252,N_14689,N_14289);
or UO_1253 (O_1253,N_12749,N_13159);
or UO_1254 (O_1254,N_12438,N_14015);
nand UO_1255 (O_1255,N_12974,N_13854);
nor UO_1256 (O_1256,N_12809,N_12014);
nor UO_1257 (O_1257,N_12161,N_12743);
nand UO_1258 (O_1258,N_13547,N_13227);
and UO_1259 (O_1259,N_13266,N_14968);
xor UO_1260 (O_1260,N_13375,N_14910);
and UO_1261 (O_1261,N_14641,N_13017);
nand UO_1262 (O_1262,N_14853,N_12732);
nor UO_1263 (O_1263,N_12794,N_14859);
and UO_1264 (O_1264,N_13039,N_13378);
and UO_1265 (O_1265,N_13330,N_12314);
nand UO_1266 (O_1266,N_12332,N_12587);
nand UO_1267 (O_1267,N_12772,N_14741);
xnor UO_1268 (O_1268,N_13963,N_14138);
nor UO_1269 (O_1269,N_14597,N_12356);
nand UO_1270 (O_1270,N_13010,N_14413);
nor UO_1271 (O_1271,N_13724,N_12843);
or UO_1272 (O_1272,N_12917,N_13022);
nor UO_1273 (O_1273,N_14230,N_12090);
xor UO_1274 (O_1274,N_13982,N_12281);
and UO_1275 (O_1275,N_12149,N_14147);
nor UO_1276 (O_1276,N_12038,N_14169);
nand UO_1277 (O_1277,N_14867,N_12978);
or UO_1278 (O_1278,N_13231,N_12588);
or UO_1279 (O_1279,N_13561,N_14061);
xor UO_1280 (O_1280,N_14122,N_13090);
xnor UO_1281 (O_1281,N_12560,N_14983);
and UO_1282 (O_1282,N_14442,N_14501);
and UO_1283 (O_1283,N_13252,N_13737);
and UO_1284 (O_1284,N_14729,N_14075);
xnor UO_1285 (O_1285,N_12503,N_14660);
xor UO_1286 (O_1286,N_12321,N_12010);
and UO_1287 (O_1287,N_12468,N_14232);
or UO_1288 (O_1288,N_14691,N_12738);
and UO_1289 (O_1289,N_14402,N_12723);
nand UO_1290 (O_1290,N_14658,N_14579);
and UO_1291 (O_1291,N_14904,N_12414);
xnor UO_1292 (O_1292,N_12234,N_14580);
or UO_1293 (O_1293,N_13013,N_12896);
nor UO_1294 (O_1294,N_14555,N_13772);
or UO_1295 (O_1295,N_12103,N_13918);
and UO_1296 (O_1296,N_14418,N_14466);
or UO_1297 (O_1297,N_12085,N_14307);
nand UO_1298 (O_1298,N_12329,N_13739);
and UO_1299 (O_1299,N_12003,N_13600);
nor UO_1300 (O_1300,N_12105,N_14181);
or UO_1301 (O_1301,N_13213,N_14785);
nor UO_1302 (O_1302,N_13431,N_14794);
or UO_1303 (O_1303,N_12385,N_13484);
or UO_1304 (O_1304,N_12036,N_12030);
nand UO_1305 (O_1305,N_14499,N_12147);
xnor UO_1306 (O_1306,N_14959,N_12813);
nor UO_1307 (O_1307,N_12122,N_12733);
nand UO_1308 (O_1308,N_14219,N_12625);
xnor UO_1309 (O_1309,N_13530,N_14044);
xnor UO_1310 (O_1310,N_14464,N_12162);
nand UO_1311 (O_1311,N_14955,N_14758);
nor UO_1312 (O_1312,N_12570,N_13319);
and UO_1313 (O_1313,N_14316,N_14385);
or UO_1314 (O_1314,N_14120,N_12713);
or UO_1315 (O_1315,N_13140,N_12462);
xnor UO_1316 (O_1316,N_12199,N_13914);
xor UO_1317 (O_1317,N_12706,N_13172);
nor UO_1318 (O_1318,N_13236,N_12889);
or UO_1319 (O_1319,N_13670,N_13769);
nor UO_1320 (O_1320,N_12697,N_14964);
and UO_1321 (O_1321,N_13796,N_14324);
xor UO_1322 (O_1322,N_12008,N_14581);
or UO_1323 (O_1323,N_14631,N_12309);
and UO_1324 (O_1324,N_13089,N_13722);
nand UO_1325 (O_1325,N_12111,N_14620);
xnor UO_1326 (O_1326,N_13637,N_13592);
xnor UO_1327 (O_1327,N_13321,N_12492);
xnor UO_1328 (O_1328,N_13023,N_13103);
and UO_1329 (O_1329,N_13642,N_12141);
and UO_1330 (O_1330,N_13581,N_14692);
nand UO_1331 (O_1331,N_13801,N_13357);
nor UO_1332 (O_1332,N_14783,N_14168);
and UO_1333 (O_1333,N_12287,N_14489);
and UO_1334 (O_1334,N_14438,N_14628);
or UO_1335 (O_1335,N_12120,N_13104);
xor UO_1336 (O_1336,N_12032,N_13629);
xor UO_1337 (O_1337,N_12056,N_14468);
xor UO_1338 (O_1338,N_13886,N_13863);
xor UO_1339 (O_1339,N_12935,N_14469);
or UO_1340 (O_1340,N_13599,N_13638);
nor UO_1341 (O_1341,N_14050,N_12166);
nor UO_1342 (O_1342,N_12691,N_13393);
xor UO_1343 (O_1343,N_13562,N_13312);
or UO_1344 (O_1344,N_14791,N_13351);
nand UO_1345 (O_1345,N_14318,N_14493);
and UO_1346 (O_1346,N_14905,N_13014);
xnor UO_1347 (O_1347,N_12707,N_14454);
and UO_1348 (O_1348,N_12734,N_12829);
nand UO_1349 (O_1349,N_12320,N_12223);
nor UO_1350 (O_1350,N_12921,N_12511);
xor UO_1351 (O_1351,N_13058,N_13282);
nand UO_1352 (O_1352,N_14211,N_13263);
xor UO_1353 (O_1353,N_12071,N_14352);
and UO_1354 (O_1354,N_13250,N_13428);
or UO_1355 (O_1355,N_12990,N_14255);
or UO_1356 (O_1356,N_14343,N_14556);
nor UO_1357 (O_1357,N_12180,N_12051);
or UO_1358 (O_1358,N_14358,N_14478);
nor UO_1359 (O_1359,N_13783,N_14416);
and UO_1360 (O_1360,N_12458,N_12856);
and UO_1361 (O_1361,N_13574,N_12916);
and UO_1362 (O_1362,N_14943,N_13651);
xnor UO_1363 (O_1363,N_13575,N_14946);
xnor UO_1364 (O_1364,N_14156,N_13580);
nand UO_1365 (O_1365,N_13920,N_12099);
xor UO_1366 (O_1366,N_12421,N_14646);
nor UO_1367 (O_1367,N_12357,N_14207);
or UO_1368 (O_1368,N_13124,N_12203);
and UO_1369 (O_1369,N_13407,N_14139);
nand UO_1370 (O_1370,N_13855,N_12634);
and UO_1371 (O_1371,N_13030,N_14200);
or UO_1372 (O_1372,N_12250,N_13153);
nand UO_1373 (O_1373,N_13684,N_14944);
xor UO_1374 (O_1374,N_14319,N_12021);
nor UO_1375 (O_1375,N_12635,N_14024);
nand UO_1376 (O_1376,N_13723,N_14332);
nor UO_1377 (O_1377,N_14315,N_13525);
and UO_1378 (O_1378,N_14799,N_13625);
and UO_1379 (O_1379,N_14522,N_13601);
and UO_1380 (O_1380,N_13702,N_14117);
or UO_1381 (O_1381,N_13703,N_14709);
xor UO_1382 (O_1382,N_14479,N_12499);
and UO_1383 (O_1383,N_13765,N_14375);
nand UO_1384 (O_1384,N_13869,N_14119);
xnor UO_1385 (O_1385,N_13067,N_14403);
xnor UO_1386 (O_1386,N_13501,N_12973);
and UO_1387 (O_1387,N_13403,N_14390);
nor UO_1388 (O_1388,N_13349,N_12191);
xor UO_1389 (O_1389,N_13328,N_14737);
nor UO_1390 (O_1390,N_13612,N_14497);
nor UO_1391 (O_1391,N_12355,N_14449);
xnor UO_1392 (O_1392,N_14954,N_13558);
and UO_1393 (O_1393,N_12537,N_14218);
or UO_1394 (O_1394,N_13405,N_13654);
and UO_1395 (O_1395,N_12995,N_13415);
nand UO_1396 (O_1396,N_13225,N_14334);
or UO_1397 (O_1397,N_14544,N_13239);
nand UO_1398 (O_1398,N_12318,N_12540);
and UO_1399 (O_1399,N_12209,N_14007);
xor UO_1400 (O_1400,N_14931,N_13242);
and UO_1401 (O_1401,N_12343,N_13028);
or UO_1402 (O_1402,N_13540,N_12108);
xnor UO_1403 (O_1403,N_12884,N_14309);
nor UO_1404 (O_1404,N_12985,N_12591);
xnor UO_1405 (O_1405,N_13275,N_12179);
or UO_1406 (O_1406,N_14446,N_12059);
nor UO_1407 (O_1407,N_13332,N_12486);
and UO_1408 (O_1408,N_14810,N_12873);
xor UO_1409 (O_1409,N_13949,N_14148);
nor UO_1410 (O_1410,N_12256,N_13736);
nor UO_1411 (O_1411,N_14625,N_14447);
or UO_1412 (O_1412,N_12583,N_13786);
or UO_1413 (O_1413,N_12204,N_14445);
nand UO_1414 (O_1414,N_14890,N_14272);
nand UO_1415 (O_1415,N_14436,N_13689);
or UO_1416 (O_1416,N_14238,N_13699);
or UO_1417 (O_1417,N_12781,N_13114);
nor UO_1418 (O_1418,N_13138,N_13665);
xnor UO_1419 (O_1419,N_12679,N_14517);
nor UO_1420 (O_1420,N_13536,N_14406);
nand UO_1421 (O_1421,N_13895,N_12423);
or UO_1422 (O_1422,N_14722,N_14668);
and UO_1423 (O_1423,N_12816,N_14627);
and UO_1424 (O_1424,N_12368,N_14297);
nand UO_1425 (O_1425,N_12317,N_12574);
xor UO_1426 (O_1426,N_13110,N_13295);
nor UO_1427 (O_1427,N_13083,N_12258);
or UO_1428 (O_1428,N_12444,N_12684);
and UO_1429 (O_1429,N_14240,N_12757);
or UO_1430 (O_1430,N_13711,N_13513);
xor UO_1431 (O_1431,N_13337,N_12165);
xnor UO_1432 (O_1432,N_13218,N_12740);
nand UO_1433 (O_1433,N_13611,N_13210);
and UO_1434 (O_1434,N_14106,N_13641);
nor UO_1435 (O_1435,N_13209,N_14520);
xnor UO_1436 (O_1436,N_12689,N_12602);
nand UO_1437 (O_1437,N_14838,N_12820);
xnor UO_1438 (O_1438,N_13216,N_12242);
or UO_1439 (O_1439,N_13101,N_13425);
nand UO_1440 (O_1440,N_12911,N_13710);
nor UO_1441 (O_1441,N_14642,N_13613);
nor UO_1442 (O_1442,N_13380,N_14528);
xnor UO_1443 (O_1443,N_12744,N_14874);
nand UO_1444 (O_1444,N_12372,N_13833);
nor UO_1445 (O_1445,N_14102,N_13294);
and UO_1446 (O_1446,N_14821,N_14566);
nor UO_1447 (O_1447,N_13874,N_13533);
nand UO_1448 (O_1448,N_14527,N_13984);
nor UO_1449 (O_1449,N_14412,N_14554);
nand UO_1450 (O_1450,N_14476,N_13494);
xor UO_1451 (O_1451,N_14801,N_14276);
and UO_1452 (O_1452,N_13620,N_13288);
xor UO_1453 (O_1453,N_12163,N_14571);
nor UO_1454 (O_1454,N_12524,N_13951);
nor UO_1455 (O_1455,N_12797,N_13456);
or UO_1456 (O_1456,N_14474,N_14074);
nor UO_1457 (O_1457,N_12001,N_14926);
or UO_1458 (O_1458,N_12620,N_12680);
nor UO_1459 (O_1459,N_14202,N_13973);
nor UO_1460 (O_1460,N_13734,N_14654);
nor UO_1461 (O_1461,N_13933,N_12005);
nand UO_1462 (O_1462,N_12745,N_12074);
nor UO_1463 (O_1463,N_13429,N_13764);
nand UO_1464 (O_1464,N_13876,N_12449);
nor UO_1465 (O_1465,N_13757,N_13688);
or UO_1466 (O_1466,N_12472,N_13166);
xnor UO_1467 (O_1467,N_13194,N_12169);
and UO_1468 (O_1468,N_13019,N_12114);
xnor UO_1469 (O_1469,N_13329,N_14180);
or UO_1470 (O_1470,N_14404,N_14536);
and UO_1471 (O_1471,N_14247,N_13624);
and UO_1472 (O_1472,N_12624,N_12046);
xnor UO_1473 (O_1473,N_12086,N_13001);
or UO_1474 (O_1474,N_14241,N_14888);
nor UO_1475 (O_1475,N_14507,N_14393);
nand UO_1476 (O_1476,N_13552,N_13049);
nand UO_1477 (O_1477,N_14360,N_13748);
and UO_1478 (O_1478,N_12268,N_12168);
nor UO_1479 (O_1479,N_14399,N_14851);
or UO_1480 (O_1480,N_12254,N_14064);
or UO_1481 (O_1481,N_14290,N_14212);
or UO_1482 (O_1482,N_12455,N_12024);
nor UO_1483 (O_1483,N_14523,N_14629);
or UO_1484 (O_1484,N_14998,N_13412);
nor UO_1485 (O_1485,N_12131,N_13810);
xor UO_1486 (O_1486,N_12905,N_13370);
xor UO_1487 (O_1487,N_14650,N_13301);
xor UO_1488 (O_1488,N_12558,N_12920);
and UO_1489 (O_1489,N_13538,N_14333);
or UO_1490 (O_1490,N_13894,N_14774);
and UO_1491 (O_1491,N_13812,N_13952);
xor UO_1492 (O_1492,N_12942,N_12398);
nand UO_1493 (O_1493,N_12219,N_14184);
nand UO_1494 (O_1494,N_14547,N_12076);
nand UO_1495 (O_1495,N_14640,N_14146);
and UO_1496 (O_1496,N_12402,N_12666);
xnor UO_1497 (O_1497,N_12452,N_14129);
nor UO_1498 (O_1498,N_14258,N_14342);
nor UO_1499 (O_1499,N_12552,N_12897);
xor UO_1500 (O_1500,N_12822,N_12238);
nor UO_1501 (O_1501,N_14568,N_14012);
xnor UO_1502 (O_1502,N_14094,N_13736);
nor UO_1503 (O_1503,N_12100,N_12579);
xor UO_1504 (O_1504,N_14969,N_13277);
nand UO_1505 (O_1505,N_13481,N_12808);
and UO_1506 (O_1506,N_14426,N_13837);
and UO_1507 (O_1507,N_12371,N_13831);
nor UO_1508 (O_1508,N_12148,N_13393);
nor UO_1509 (O_1509,N_12807,N_14356);
nor UO_1510 (O_1510,N_13726,N_12909);
nor UO_1511 (O_1511,N_12056,N_12271);
and UO_1512 (O_1512,N_12101,N_13620);
nor UO_1513 (O_1513,N_14602,N_14302);
or UO_1514 (O_1514,N_12547,N_12163);
nand UO_1515 (O_1515,N_14398,N_12503);
xnor UO_1516 (O_1516,N_13430,N_14155);
or UO_1517 (O_1517,N_14608,N_14932);
and UO_1518 (O_1518,N_13596,N_12099);
and UO_1519 (O_1519,N_13794,N_14173);
or UO_1520 (O_1520,N_14211,N_13492);
or UO_1521 (O_1521,N_13639,N_12010);
and UO_1522 (O_1522,N_14887,N_13981);
nand UO_1523 (O_1523,N_12259,N_13152);
and UO_1524 (O_1524,N_12578,N_14116);
nand UO_1525 (O_1525,N_12093,N_14010);
or UO_1526 (O_1526,N_13926,N_12597);
nor UO_1527 (O_1527,N_14458,N_14938);
and UO_1528 (O_1528,N_14655,N_13860);
or UO_1529 (O_1529,N_12170,N_13318);
nand UO_1530 (O_1530,N_13090,N_12309);
and UO_1531 (O_1531,N_12346,N_12044);
nand UO_1532 (O_1532,N_14734,N_12176);
xnor UO_1533 (O_1533,N_13380,N_14635);
xor UO_1534 (O_1534,N_14684,N_13513);
nand UO_1535 (O_1535,N_13457,N_12319);
or UO_1536 (O_1536,N_14692,N_14580);
and UO_1537 (O_1537,N_12505,N_12437);
and UO_1538 (O_1538,N_12982,N_13930);
and UO_1539 (O_1539,N_13860,N_13981);
xor UO_1540 (O_1540,N_12827,N_12599);
or UO_1541 (O_1541,N_13953,N_13651);
xnor UO_1542 (O_1542,N_12982,N_12637);
or UO_1543 (O_1543,N_13272,N_14580);
nand UO_1544 (O_1544,N_12153,N_14436);
or UO_1545 (O_1545,N_14827,N_13391);
or UO_1546 (O_1546,N_12311,N_14545);
nand UO_1547 (O_1547,N_13638,N_12683);
xnor UO_1548 (O_1548,N_12382,N_14268);
or UO_1549 (O_1549,N_14021,N_14979);
and UO_1550 (O_1550,N_13648,N_14543);
nor UO_1551 (O_1551,N_12990,N_13538);
nand UO_1552 (O_1552,N_12898,N_13666);
and UO_1553 (O_1553,N_14556,N_12650);
xor UO_1554 (O_1554,N_14396,N_13859);
and UO_1555 (O_1555,N_13151,N_13890);
xnor UO_1556 (O_1556,N_13391,N_13888);
or UO_1557 (O_1557,N_13659,N_14069);
nand UO_1558 (O_1558,N_12162,N_14160);
and UO_1559 (O_1559,N_13658,N_12145);
nand UO_1560 (O_1560,N_13606,N_12946);
or UO_1561 (O_1561,N_12865,N_13273);
nand UO_1562 (O_1562,N_14972,N_13288);
nand UO_1563 (O_1563,N_12861,N_13381);
nor UO_1564 (O_1564,N_12125,N_13523);
and UO_1565 (O_1565,N_14430,N_14798);
and UO_1566 (O_1566,N_14035,N_13742);
and UO_1567 (O_1567,N_14732,N_12082);
or UO_1568 (O_1568,N_14592,N_13093);
xor UO_1569 (O_1569,N_12390,N_12786);
xnor UO_1570 (O_1570,N_14353,N_12246);
and UO_1571 (O_1571,N_12440,N_13053);
xor UO_1572 (O_1572,N_14123,N_14383);
and UO_1573 (O_1573,N_12851,N_12762);
or UO_1574 (O_1574,N_12255,N_12535);
nand UO_1575 (O_1575,N_13428,N_12045);
and UO_1576 (O_1576,N_14656,N_14559);
nand UO_1577 (O_1577,N_13906,N_12460);
or UO_1578 (O_1578,N_13428,N_13758);
nand UO_1579 (O_1579,N_12033,N_12479);
or UO_1580 (O_1580,N_14744,N_13685);
nand UO_1581 (O_1581,N_14957,N_13641);
nand UO_1582 (O_1582,N_13263,N_14101);
xor UO_1583 (O_1583,N_13002,N_14022);
nand UO_1584 (O_1584,N_13723,N_12288);
nor UO_1585 (O_1585,N_12472,N_12188);
xnor UO_1586 (O_1586,N_12447,N_13100);
nand UO_1587 (O_1587,N_14114,N_12914);
or UO_1588 (O_1588,N_12677,N_12500);
nor UO_1589 (O_1589,N_13975,N_12031);
and UO_1590 (O_1590,N_14969,N_12965);
or UO_1591 (O_1591,N_13782,N_14373);
and UO_1592 (O_1592,N_13311,N_14994);
xnor UO_1593 (O_1593,N_12563,N_14477);
nor UO_1594 (O_1594,N_12757,N_13351);
xnor UO_1595 (O_1595,N_14758,N_13480);
nand UO_1596 (O_1596,N_14879,N_13339);
nand UO_1597 (O_1597,N_12049,N_14138);
nor UO_1598 (O_1598,N_13811,N_13275);
or UO_1599 (O_1599,N_13620,N_14425);
xnor UO_1600 (O_1600,N_14912,N_13725);
nand UO_1601 (O_1601,N_14712,N_13726);
or UO_1602 (O_1602,N_14702,N_14426);
and UO_1603 (O_1603,N_12176,N_13829);
or UO_1604 (O_1604,N_13166,N_14135);
xor UO_1605 (O_1605,N_13577,N_13514);
or UO_1606 (O_1606,N_12082,N_13716);
nor UO_1607 (O_1607,N_12414,N_13139);
nand UO_1608 (O_1608,N_14170,N_12897);
and UO_1609 (O_1609,N_13932,N_13971);
nand UO_1610 (O_1610,N_12476,N_14349);
xnor UO_1611 (O_1611,N_14341,N_12534);
or UO_1612 (O_1612,N_12241,N_14716);
xnor UO_1613 (O_1613,N_12970,N_14627);
or UO_1614 (O_1614,N_12081,N_14356);
nor UO_1615 (O_1615,N_12172,N_12824);
xor UO_1616 (O_1616,N_12030,N_14512);
nor UO_1617 (O_1617,N_14049,N_12338);
nand UO_1618 (O_1618,N_12890,N_12920);
xor UO_1619 (O_1619,N_12474,N_14613);
nor UO_1620 (O_1620,N_14513,N_14245);
nor UO_1621 (O_1621,N_12437,N_14440);
nor UO_1622 (O_1622,N_13277,N_13411);
nor UO_1623 (O_1623,N_14899,N_13207);
xor UO_1624 (O_1624,N_12713,N_12839);
nand UO_1625 (O_1625,N_13154,N_13524);
nor UO_1626 (O_1626,N_14085,N_14466);
and UO_1627 (O_1627,N_13412,N_13637);
and UO_1628 (O_1628,N_13586,N_14763);
nand UO_1629 (O_1629,N_13480,N_12201);
nand UO_1630 (O_1630,N_13754,N_13687);
nand UO_1631 (O_1631,N_13180,N_13529);
nor UO_1632 (O_1632,N_12498,N_12276);
nor UO_1633 (O_1633,N_13013,N_14999);
nand UO_1634 (O_1634,N_14798,N_13522);
xnor UO_1635 (O_1635,N_12425,N_12720);
nand UO_1636 (O_1636,N_12771,N_13720);
xnor UO_1637 (O_1637,N_12717,N_13916);
xnor UO_1638 (O_1638,N_13717,N_14147);
nand UO_1639 (O_1639,N_13501,N_14489);
or UO_1640 (O_1640,N_12470,N_13070);
nor UO_1641 (O_1641,N_14164,N_14143);
nand UO_1642 (O_1642,N_12177,N_12355);
or UO_1643 (O_1643,N_12796,N_13405);
xor UO_1644 (O_1644,N_14730,N_13085);
xor UO_1645 (O_1645,N_13359,N_12318);
xnor UO_1646 (O_1646,N_12130,N_13305);
or UO_1647 (O_1647,N_14574,N_12468);
xnor UO_1648 (O_1648,N_13653,N_12581);
nor UO_1649 (O_1649,N_14233,N_13236);
or UO_1650 (O_1650,N_14056,N_13608);
or UO_1651 (O_1651,N_12094,N_14764);
nor UO_1652 (O_1652,N_13447,N_14183);
xnor UO_1653 (O_1653,N_12955,N_13100);
nor UO_1654 (O_1654,N_14663,N_14657);
nor UO_1655 (O_1655,N_14495,N_12851);
xor UO_1656 (O_1656,N_14372,N_13785);
nand UO_1657 (O_1657,N_13298,N_12109);
xnor UO_1658 (O_1658,N_13275,N_12566);
nand UO_1659 (O_1659,N_12736,N_12468);
or UO_1660 (O_1660,N_12179,N_14370);
xor UO_1661 (O_1661,N_12404,N_13166);
xor UO_1662 (O_1662,N_12677,N_12512);
nand UO_1663 (O_1663,N_12059,N_14336);
or UO_1664 (O_1664,N_14086,N_14379);
xor UO_1665 (O_1665,N_14022,N_14539);
nand UO_1666 (O_1666,N_12496,N_13037);
or UO_1667 (O_1667,N_12926,N_13963);
nor UO_1668 (O_1668,N_12094,N_12555);
nand UO_1669 (O_1669,N_12131,N_14494);
or UO_1670 (O_1670,N_12226,N_13324);
xnor UO_1671 (O_1671,N_12273,N_14806);
and UO_1672 (O_1672,N_12437,N_13687);
or UO_1673 (O_1673,N_14689,N_12968);
xor UO_1674 (O_1674,N_13373,N_13999);
xnor UO_1675 (O_1675,N_13326,N_13765);
xor UO_1676 (O_1676,N_13844,N_13603);
xnor UO_1677 (O_1677,N_14499,N_14830);
nor UO_1678 (O_1678,N_12366,N_12617);
nand UO_1679 (O_1679,N_12111,N_14130);
and UO_1680 (O_1680,N_14700,N_13095);
nand UO_1681 (O_1681,N_12852,N_14692);
and UO_1682 (O_1682,N_12402,N_12798);
nor UO_1683 (O_1683,N_12069,N_12688);
or UO_1684 (O_1684,N_13193,N_13166);
or UO_1685 (O_1685,N_12739,N_12366);
xnor UO_1686 (O_1686,N_12956,N_12816);
nor UO_1687 (O_1687,N_12128,N_14548);
and UO_1688 (O_1688,N_12654,N_12586);
xnor UO_1689 (O_1689,N_12555,N_13644);
nand UO_1690 (O_1690,N_12102,N_14116);
and UO_1691 (O_1691,N_13398,N_13277);
nand UO_1692 (O_1692,N_12029,N_13044);
and UO_1693 (O_1693,N_14724,N_12582);
xnor UO_1694 (O_1694,N_12274,N_14997);
nor UO_1695 (O_1695,N_13284,N_14860);
xor UO_1696 (O_1696,N_12664,N_13123);
nor UO_1697 (O_1697,N_12666,N_13369);
or UO_1698 (O_1698,N_13228,N_12169);
nand UO_1699 (O_1699,N_12132,N_13381);
nand UO_1700 (O_1700,N_13542,N_12974);
or UO_1701 (O_1701,N_12966,N_12524);
xnor UO_1702 (O_1702,N_12976,N_12012);
and UO_1703 (O_1703,N_13168,N_14053);
nand UO_1704 (O_1704,N_14571,N_13930);
nor UO_1705 (O_1705,N_13461,N_14719);
nor UO_1706 (O_1706,N_14331,N_14189);
xor UO_1707 (O_1707,N_14946,N_12861);
or UO_1708 (O_1708,N_13187,N_12736);
xor UO_1709 (O_1709,N_13797,N_13595);
nor UO_1710 (O_1710,N_13882,N_12423);
and UO_1711 (O_1711,N_12090,N_14891);
and UO_1712 (O_1712,N_13960,N_12831);
nand UO_1713 (O_1713,N_13367,N_14649);
and UO_1714 (O_1714,N_12487,N_14673);
and UO_1715 (O_1715,N_13003,N_14825);
xnor UO_1716 (O_1716,N_13760,N_12560);
nor UO_1717 (O_1717,N_13406,N_12461);
xnor UO_1718 (O_1718,N_14843,N_14206);
or UO_1719 (O_1719,N_13416,N_14915);
and UO_1720 (O_1720,N_13832,N_14332);
xnor UO_1721 (O_1721,N_13118,N_13367);
or UO_1722 (O_1722,N_12482,N_13180);
or UO_1723 (O_1723,N_14384,N_13098);
or UO_1724 (O_1724,N_14439,N_12257);
nor UO_1725 (O_1725,N_14275,N_12909);
xor UO_1726 (O_1726,N_12373,N_13656);
nor UO_1727 (O_1727,N_12602,N_14080);
or UO_1728 (O_1728,N_14243,N_12571);
and UO_1729 (O_1729,N_14627,N_12458);
nor UO_1730 (O_1730,N_12137,N_13243);
or UO_1731 (O_1731,N_14708,N_14834);
nor UO_1732 (O_1732,N_14119,N_14808);
nor UO_1733 (O_1733,N_14685,N_14355);
nand UO_1734 (O_1734,N_13909,N_12128);
or UO_1735 (O_1735,N_13995,N_14839);
xor UO_1736 (O_1736,N_12634,N_13192);
xor UO_1737 (O_1737,N_13837,N_13681);
and UO_1738 (O_1738,N_12267,N_14168);
xor UO_1739 (O_1739,N_14421,N_12158);
nor UO_1740 (O_1740,N_12190,N_12584);
or UO_1741 (O_1741,N_14917,N_12964);
xor UO_1742 (O_1742,N_13951,N_13612);
nor UO_1743 (O_1743,N_13807,N_13450);
nor UO_1744 (O_1744,N_12784,N_14433);
or UO_1745 (O_1745,N_13989,N_14360);
nor UO_1746 (O_1746,N_13487,N_14968);
or UO_1747 (O_1747,N_13706,N_14077);
and UO_1748 (O_1748,N_14416,N_14956);
nor UO_1749 (O_1749,N_12426,N_12346);
and UO_1750 (O_1750,N_12632,N_13223);
and UO_1751 (O_1751,N_13602,N_13861);
nand UO_1752 (O_1752,N_14641,N_13731);
xnor UO_1753 (O_1753,N_13439,N_14777);
xor UO_1754 (O_1754,N_13145,N_14457);
and UO_1755 (O_1755,N_14562,N_12417);
and UO_1756 (O_1756,N_12795,N_12641);
and UO_1757 (O_1757,N_13229,N_12366);
xnor UO_1758 (O_1758,N_12773,N_14881);
xnor UO_1759 (O_1759,N_12525,N_14604);
nor UO_1760 (O_1760,N_13734,N_12222);
nand UO_1761 (O_1761,N_12970,N_13015);
nand UO_1762 (O_1762,N_12759,N_12494);
nor UO_1763 (O_1763,N_14594,N_12253);
nand UO_1764 (O_1764,N_13160,N_12089);
xor UO_1765 (O_1765,N_13516,N_13017);
nand UO_1766 (O_1766,N_14042,N_13874);
nand UO_1767 (O_1767,N_14727,N_12920);
nor UO_1768 (O_1768,N_14909,N_14505);
xnor UO_1769 (O_1769,N_12515,N_12610);
nand UO_1770 (O_1770,N_12364,N_12777);
or UO_1771 (O_1771,N_12722,N_13979);
nor UO_1772 (O_1772,N_14424,N_12094);
nor UO_1773 (O_1773,N_13213,N_12637);
and UO_1774 (O_1774,N_14695,N_12170);
nor UO_1775 (O_1775,N_14203,N_14106);
or UO_1776 (O_1776,N_14444,N_12828);
xor UO_1777 (O_1777,N_12879,N_13298);
xor UO_1778 (O_1778,N_13428,N_12109);
nor UO_1779 (O_1779,N_13566,N_14699);
nand UO_1780 (O_1780,N_12523,N_13089);
xor UO_1781 (O_1781,N_12596,N_13331);
nor UO_1782 (O_1782,N_14108,N_14176);
or UO_1783 (O_1783,N_14117,N_13333);
nand UO_1784 (O_1784,N_12365,N_12483);
nand UO_1785 (O_1785,N_13979,N_13323);
or UO_1786 (O_1786,N_13633,N_13227);
nor UO_1787 (O_1787,N_12637,N_14326);
nand UO_1788 (O_1788,N_13058,N_13123);
nor UO_1789 (O_1789,N_14055,N_13527);
and UO_1790 (O_1790,N_14235,N_13680);
nand UO_1791 (O_1791,N_12794,N_12992);
nand UO_1792 (O_1792,N_13622,N_14789);
and UO_1793 (O_1793,N_14199,N_12105);
or UO_1794 (O_1794,N_14999,N_13612);
xnor UO_1795 (O_1795,N_14966,N_13384);
nor UO_1796 (O_1796,N_14074,N_12558);
xor UO_1797 (O_1797,N_14313,N_14894);
nand UO_1798 (O_1798,N_12176,N_14543);
nor UO_1799 (O_1799,N_12530,N_13472);
and UO_1800 (O_1800,N_12337,N_13555);
and UO_1801 (O_1801,N_13578,N_13888);
or UO_1802 (O_1802,N_13803,N_13014);
and UO_1803 (O_1803,N_12203,N_13035);
or UO_1804 (O_1804,N_13850,N_13361);
or UO_1805 (O_1805,N_14029,N_12668);
xor UO_1806 (O_1806,N_14217,N_13284);
nor UO_1807 (O_1807,N_12230,N_13935);
xor UO_1808 (O_1808,N_13005,N_12815);
nand UO_1809 (O_1809,N_14465,N_12468);
nand UO_1810 (O_1810,N_13745,N_13227);
nor UO_1811 (O_1811,N_14473,N_14678);
or UO_1812 (O_1812,N_14116,N_14771);
or UO_1813 (O_1813,N_14917,N_14513);
and UO_1814 (O_1814,N_12354,N_14608);
nor UO_1815 (O_1815,N_12454,N_12051);
or UO_1816 (O_1816,N_13916,N_12287);
xnor UO_1817 (O_1817,N_13642,N_14508);
and UO_1818 (O_1818,N_12468,N_14036);
or UO_1819 (O_1819,N_12229,N_13241);
and UO_1820 (O_1820,N_14220,N_14884);
and UO_1821 (O_1821,N_13243,N_13015);
nand UO_1822 (O_1822,N_14541,N_12215);
nor UO_1823 (O_1823,N_14164,N_14331);
or UO_1824 (O_1824,N_12877,N_12188);
nor UO_1825 (O_1825,N_12164,N_12643);
or UO_1826 (O_1826,N_13194,N_12268);
or UO_1827 (O_1827,N_13877,N_12855);
nand UO_1828 (O_1828,N_14493,N_13895);
or UO_1829 (O_1829,N_13406,N_14379);
nand UO_1830 (O_1830,N_14599,N_14239);
nor UO_1831 (O_1831,N_14460,N_14420);
or UO_1832 (O_1832,N_14575,N_14937);
xor UO_1833 (O_1833,N_14484,N_14966);
nand UO_1834 (O_1834,N_13338,N_12504);
nor UO_1835 (O_1835,N_12092,N_14673);
and UO_1836 (O_1836,N_12250,N_14709);
nand UO_1837 (O_1837,N_13288,N_14861);
nand UO_1838 (O_1838,N_14958,N_12040);
and UO_1839 (O_1839,N_14924,N_13855);
nor UO_1840 (O_1840,N_14962,N_14622);
or UO_1841 (O_1841,N_13482,N_13050);
nor UO_1842 (O_1842,N_13441,N_13385);
and UO_1843 (O_1843,N_14189,N_13852);
nor UO_1844 (O_1844,N_14569,N_12394);
xor UO_1845 (O_1845,N_13148,N_14897);
and UO_1846 (O_1846,N_13164,N_14525);
xor UO_1847 (O_1847,N_12491,N_14787);
nor UO_1848 (O_1848,N_13609,N_12894);
or UO_1849 (O_1849,N_13002,N_14582);
xor UO_1850 (O_1850,N_14556,N_12585);
nand UO_1851 (O_1851,N_12811,N_13328);
nor UO_1852 (O_1852,N_14033,N_14011);
nand UO_1853 (O_1853,N_13876,N_13957);
or UO_1854 (O_1854,N_12046,N_14170);
nand UO_1855 (O_1855,N_12194,N_13088);
and UO_1856 (O_1856,N_14707,N_12013);
xnor UO_1857 (O_1857,N_14018,N_14802);
xnor UO_1858 (O_1858,N_12431,N_14890);
nand UO_1859 (O_1859,N_14022,N_13949);
nand UO_1860 (O_1860,N_12809,N_12204);
nor UO_1861 (O_1861,N_14763,N_12857);
xnor UO_1862 (O_1862,N_14907,N_13618);
xnor UO_1863 (O_1863,N_12045,N_12874);
or UO_1864 (O_1864,N_14738,N_13154);
nand UO_1865 (O_1865,N_13812,N_13594);
or UO_1866 (O_1866,N_14969,N_14138);
xnor UO_1867 (O_1867,N_13178,N_14292);
or UO_1868 (O_1868,N_12580,N_12694);
and UO_1869 (O_1869,N_13370,N_13491);
and UO_1870 (O_1870,N_12093,N_12328);
nand UO_1871 (O_1871,N_13397,N_12498);
xnor UO_1872 (O_1872,N_13358,N_12772);
nand UO_1873 (O_1873,N_13088,N_14583);
and UO_1874 (O_1874,N_13012,N_14133);
nand UO_1875 (O_1875,N_13309,N_14803);
nand UO_1876 (O_1876,N_13474,N_14795);
or UO_1877 (O_1877,N_13654,N_12943);
or UO_1878 (O_1878,N_13174,N_13534);
or UO_1879 (O_1879,N_14535,N_12052);
nand UO_1880 (O_1880,N_14929,N_14609);
and UO_1881 (O_1881,N_14989,N_13250);
nand UO_1882 (O_1882,N_14526,N_12709);
xor UO_1883 (O_1883,N_12264,N_14461);
and UO_1884 (O_1884,N_13418,N_13250);
nor UO_1885 (O_1885,N_13005,N_12976);
nand UO_1886 (O_1886,N_12349,N_12170);
nor UO_1887 (O_1887,N_13933,N_13375);
xnor UO_1888 (O_1888,N_14853,N_13413);
or UO_1889 (O_1889,N_14281,N_14193);
nand UO_1890 (O_1890,N_14744,N_13159);
nor UO_1891 (O_1891,N_13438,N_13295);
and UO_1892 (O_1892,N_12656,N_14335);
or UO_1893 (O_1893,N_12190,N_13455);
and UO_1894 (O_1894,N_14037,N_13103);
nor UO_1895 (O_1895,N_12182,N_13102);
xnor UO_1896 (O_1896,N_13321,N_12443);
or UO_1897 (O_1897,N_14764,N_14489);
nand UO_1898 (O_1898,N_12839,N_12925);
nand UO_1899 (O_1899,N_14151,N_13001);
nor UO_1900 (O_1900,N_12554,N_14345);
xnor UO_1901 (O_1901,N_14495,N_13779);
xnor UO_1902 (O_1902,N_14825,N_13457);
xor UO_1903 (O_1903,N_12292,N_14946);
nand UO_1904 (O_1904,N_14812,N_12054);
nor UO_1905 (O_1905,N_13568,N_13427);
or UO_1906 (O_1906,N_12320,N_13028);
nand UO_1907 (O_1907,N_13069,N_14065);
or UO_1908 (O_1908,N_14378,N_14799);
xor UO_1909 (O_1909,N_12933,N_12199);
xnor UO_1910 (O_1910,N_13702,N_13917);
nand UO_1911 (O_1911,N_13871,N_13289);
or UO_1912 (O_1912,N_14383,N_12634);
nor UO_1913 (O_1913,N_14220,N_12156);
nor UO_1914 (O_1914,N_14675,N_14337);
or UO_1915 (O_1915,N_13556,N_12909);
and UO_1916 (O_1916,N_14498,N_12911);
xnor UO_1917 (O_1917,N_13517,N_14215);
nor UO_1918 (O_1918,N_12302,N_13190);
or UO_1919 (O_1919,N_13120,N_12936);
nor UO_1920 (O_1920,N_14886,N_14221);
xnor UO_1921 (O_1921,N_14547,N_14520);
nor UO_1922 (O_1922,N_12517,N_14950);
xor UO_1923 (O_1923,N_13387,N_13104);
xor UO_1924 (O_1924,N_12242,N_13429);
xnor UO_1925 (O_1925,N_14258,N_13360);
nor UO_1926 (O_1926,N_12174,N_13622);
xor UO_1927 (O_1927,N_14925,N_12439);
xor UO_1928 (O_1928,N_12023,N_12767);
and UO_1929 (O_1929,N_14514,N_12951);
nor UO_1930 (O_1930,N_12643,N_13626);
or UO_1931 (O_1931,N_13768,N_13381);
and UO_1932 (O_1932,N_12151,N_12782);
xor UO_1933 (O_1933,N_13923,N_14115);
xor UO_1934 (O_1934,N_14338,N_12102);
and UO_1935 (O_1935,N_13575,N_14066);
nor UO_1936 (O_1936,N_14342,N_12297);
or UO_1937 (O_1937,N_12474,N_13819);
nor UO_1938 (O_1938,N_12809,N_12854);
or UO_1939 (O_1939,N_13766,N_12404);
and UO_1940 (O_1940,N_13361,N_14847);
and UO_1941 (O_1941,N_14535,N_14764);
xnor UO_1942 (O_1942,N_12043,N_13983);
and UO_1943 (O_1943,N_12257,N_12022);
and UO_1944 (O_1944,N_13346,N_13169);
nor UO_1945 (O_1945,N_12238,N_14076);
xor UO_1946 (O_1946,N_12463,N_12635);
and UO_1947 (O_1947,N_13683,N_12079);
and UO_1948 (O_1948,N_14682,N_14226);
nor UO_1949 (O_1949,N_12321,N_14821);
or UO_1950 (O_1950,N_14724,N_12390);
nand UO_1951 (O_1951,N_14725,N_12773);
nor UO_1952 (O_1952,N_14966,N_14013);
or UO_1953 (O_1953,N_13496,N_14966);
xor UO_1954 (O_1954,N_12533,N_13853);
and UO_1955 (O_1955,N_14364,N_12920);
or UO_1956 (O_1956,N_13225,N_14112);
or UO_1957 (O_1957,N_12322,N_13738);
or UO_1958 (O_1958,N_13815,N_12316);
or UO_1959 (O_1959,N_14265,N_13398);
nand UO_1960 (O_1960,N_14376,N_12938);
or UO_1961 (O_1961,N_14015,N_13485);
xnor UO_1962 (O_1962,N_14897,N_13517);
xnor UO_1963 (O_1963,N_12424,N_13031);
xor UO_1964 (O_1964,N_14017,N_13090);
nor UO_1965 (O_1965,N_12828,N_13916);
and UO_1966 (O_1966,N_14300,N_14539);
xnor UO_1967 (O_1967,N_14379,N_12073);
nand UO_1968 (O_1968,N_13163,N_12610);
or UO_1969 (O_1969,N_13431,N_14238);
xor UO_1970 (O_1970,N_14034,N_12341);
xnor UO_1971 (O_1971,N_14513,N_13980);
or UO_1972 (O_1972,N_13873,N_12650);
nand UO_1973 (O_1973,N_13637,N_12400);
nand UO_1974 (O_1974,N_14365,N_12907);
xnor UO_1975 (O_1975,N_13254,N_12877);
nand UO_1976 (O_1976,N_13991,N_13243);
nor UO_1977 (O_1977,N_12655,N_13430);
and UO_1978 (O_1978,N_14815,N_13137);
nand UO_1979 (O_1979,N_12762,N_14228);
and UO_1980 (O_1980,N_13578,N_12562);
or UO_1981 (O_1981,N_12695,N_13670);
xnor UO_1982 (O_1982,N_14752,N_12310);
nand UO_1983 (O_1983,N_14970,N_13045);
nor UO_1984 (O_1984,N_14497,N_14744);
xnor UO_1985 (O_1985,N_13627,N_13918);
nand UO_1986 (O_1986,N_13311,N_12839);
and UO_1987 (O_1987,N_13944,N_13454);
or UO_1988 (O_1988,N_13487,N_14050);
or UO_1989 (O_1989,N_13540,N_14977);
xor UO_1990 (O_1990,N_12576,N_14684);
nand UO_1991 (O_1991,N_13083,N_14465);
nor UO_1992 (O_1992,N_12349,N_14614);
nor UO_1993 (O_1993,N_12938,N_12468);
or UO_1994 (O_1994,N_13137,N_13260);
or UO_1995 (O_1995,N_12380,N_13058);
and UO_1996 (O_1996,N_14941,N_13333);
nand UO_1997 (O_1997,N_13152,N_12630);
nor UO_1998 (O_1998,N_12069,N_13755);
nor UO_1999 (O_1999,N_13142,N_14697);
endmodule