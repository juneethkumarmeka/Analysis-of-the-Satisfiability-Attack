module basic_2000_20000_2500_5_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1244,In_754);
and U1 (N_1,In_480,In_1804);
or U2 (N_2,In_923,In_517);
nor U3 (N_3,In_751,In_783);
nor U4 (N_4,In_1507,In_895);
nor U5 (N_5,In_494,In_507);
or U6 (N_6,In_1220,In_1834);
and U7 (N_7,In_1577,In_1955);
nand U8 (N_8,In_1491,In_270);
or U9 (N_9,In_1318,In_1166);
nor U10 (N_10,In_141,In_840);
nand U11 (N_11,In_631,In_20);
nand U12 (N_12,In_676,In_687);
nor U13 (N_13,In_1580,In_1432);
nor U14 (N_14,In_886,In_1987);
nand U15 (N_15,In_1143,In_168);
nor U16 (N_16,In_1963,In_1036);
nand U17 (N_17,In_881,In_487);
and U18 (N_18,In_1661,In_1392);
or U19 (N_19,In_818,In_1409);
nand U20 (N_20,In_1650,In_1422);
and U21 (N_21,In_336,In_1606);
nor U22 (N_22,In_1836,In_1099);
and U23 (N_23,In_1271,In_712);
nand U24 (N_24,In_597,In_256);
xor U25 (N_25,In_1717,In_1696);
nand U26 (N_26,In_994,In_1512);
and U27 (N_27,In_273,In_603);
and U28 (N_28,In_1935,In_607);
or U29 (N_29,In_1436,In_1574);
nor U30 (N_30,In_1904,In_972);
or U31 (N_31,In_866,In_1969);
or U32 (N_32,In_1229,In_1918);
nand U33 (N_33,In_1346,In_1452);
nand U34 (N_34,In_147,In_76);
or U35 (N_35,In_718,In_1303);
nor U36 (N_36,In_1594,In_1769);
nor U37 (N_37,In_1351,In_1479);
xnor U38 (N_38,In_1371,In_1757);
and U39 (N_39,In_1224,In_1015);
and U40 (N_40,In_700,In_56);
xnor U41 (N_41,In_1498,In_1389);
nand U42 (N_42,In_1533,In_945);
nand U43 (N_43,In_1,In_1932);
nand U44 (N_44,In_1334,In_239);
nand U45 (N_45,In_1078,In_1654);
and U46 (N_46,In_417,In_1849);
and U47 (N_47,In_341,In_1196);
nor U48 (N_48,In_1793,In_1352);
xnor U49 (N_49,In_442,In_102);
xor U50 (N_50,In_1828,In_1767);
nor U51 (N_51,In_1554,In_734);
nand U52 (N_52,In_218,In_1807);
or U53 (N_53,In_965,In_1130);
and U54 (N_54,In_1879,In_1892);
or U55 (N_55,In_842,In_544);
and U56 (N_56,In_422,In_1556);
nand U57 (N_57,In_1517,In_28);
nor U58 (N_58,In_1226,In_660);
nand U59 (N_59,In_784,In_41);
or U60 (N_60,In_755,In_777);
nor U61 (N_61,In_1230,In_1047);
xnor U62 (N_62,In_1476,In_1764);
nand U63 (N_63,In_1178,In_694);
nand U64 (N_64,In_1949,In_690);
nand U65 (N_65,In_1321,In_741);
or U66 (N_66,In_1617,In_1273);
or U67 (N_67,In_760,In_1845);
or U68 (N_68,In_430,In_1658);
and U69 (N_69,In_1189,In_1798);
nor U70 (N_70,In_397,In_987);
nand U71 (N_71,In_974,In_1296);
nor U72 (N_72,In_1778,In_95);
nor U73 (N_73,In_641,In_1900);
nor U74 (N_74,In_1823,In_816);
and U75 (N_75,In_1232,In_1140);
or U76 (N_76,In_101,In_546);
or U77 (N_77,In_1265,In_6);
nor U78 (N_78,In_497,In_1528);
or U79 (N_79,In_366,In_1298);
and U80 (N_80,In_1869,In_1282);
nand U81 (N_81,In_635,In_405);
nand U82 (N_82,In_1379,In_1890);
and U83 (N_83,In_390,In_1020);
or U84 (N_84,In_899,In_431);
or U85 (N_85,In_1384,In_1366);
and U86 (N_86,In_991,In_950);
nand U87 (N_87,In_1234,In_1284);
and U88 (N_88,In_1593,In_549);
nor U89 (N_89,In_1103,In_1876);
nand U90 (N_90,In_1250,In_1923);
nor U91 (N_91,In_268,In_1263);
nand U92 (N_92,In_815,In_992);
nor U93 (N_93,In_1309,In_1082);
nor U94 (N_94,In_304,In_155);
nor U95 (N_95,In_524,In_161);
xor U96 (N_96,In_902,In_1182);
xnor U97 (N_97,In_496,In_329);
and U98 (N_98,In_512,In_677);
nand U99 (N_99,In_1449,In_1427);
and U100 (N_100,In_1564,In_327);
and U101 (N_101,In_1456,In_1046);
or U102 (N_102,In_1655,In_684);
and U103 (N_103,In_1790,In_423);
nor U104 (N_104,In_583,In_1114);
or U105 (N_105,In_36,In_1733);
and U106 (N_106,In_1494,In_449);
and U107 (N_107,In_484,In_1687);
nor U108 (N_108,In_115,In_1348);
nand U109 (N_109,In_1252,In_1181);
xor U110 (N_110,In_547,In_1728);
or U111 (N_111,In_404,In_1602);
nand U112 (N_112,In_1508,In_1908);
and U113 (N_113,In_403,In_692);
nor U114 (N_114,In_1920,In_282);
or U115 (N_115,In_514,In_1947);
nand U116 (N_116,In_339,In_295);
or U117 (N_117,In_1221,In_666);
or U118 (N_118,In_858,In_1722);
and U119 (N_119,In_697,In_535);
nand U120 (N_120,In_503,In_1051);
nor U121 (N_121,In_1489,In_10);
and U122 (N_122,In_1727,In_340);
and U123 (N_123,In_444,In_811);
nand U124 (N_124,In_861,In_1780);
or U125 (N_125,In_675,In_1522);
and U126 (N_126,In_771,In_647);
xor U127 (N_127,In_817,In_427);
and U128 (N_128,In_800,In_707);
xor U129 (N_129,In_1608,In_1360);
xnor U130 (N_130,In_636,In_1510);
nor U131 (N_131,In_1450,In_1715);
nor U132 (N_132,In_1830,In_1172);
nand U133 (N_133,In_306,In_511);
or U134 (N_134,In_605,In_1610);
and U135 (N_135,In_1744,In_890);
or U136 (N_136,In_1647,In_468);
nor U137 (N_137,In_1419,In_633);
or U138 (N_138,In_960,In_1493);
nand U139 (N_139,In_1395,In_1964);
nor U140 (N_140,In_195,In_98);
or U141 (N_141,In_1812,In_1848);
or U142 (N_142,In_964,In_1049);
nand U143 (N_143,In_1913,In_222);
nand U144 (N_144,In_180,In_1803);
or U145 (N_145,In_352,In_1154);
nand U146 (N_146,In_399,In_714);
or U147 (N_147,In_587,In_164);
nand U148 (N_148,In_1177,In_111);
xor U149 (N_149,In_1705,In_383);
and U150 (N_150,In_542,In_22);
or U151 (N_151,In_778,In_1539);
and U152 (N_152,In_61,In_318);
xor U153 (N_153,In_826,In_148);
nand U154 (N_154,In_735,In_1745);
xor U155 (N_155,In_1292,In_223);
or U156 (N_156,In_903,In_1361);
and U157 (N_157,In_841,In_411);
nand U158 (N_158,In_1576,In_303);
nor U159 (N_159,In_129,In_1041);
or U160 (N_160,In_516,In_1219);
nor U161 (N_161,In_371,In_1458);
nor U162 (N_162,In_1482,In_710);
and U163 (N_163,In_130,In_1938);
or U164 (N_164,In_458,In_326);
or U165 (N_165,In_679,In_1560);
nor U166 (N_166,In_1865,In_49);
and U167 (N_167,In_1741,In_1754);
nor U168 (N_168,In_1989,In_259);
or U169 (N_169,In_1162,In_1894);
nand U170 (N_170,In_254,In_1697);
xnor U171 (N_171,In_642,In_1978);
nand U172 (N_172,In_1363,In_1994);
or U173 (N_173,In_1710,In_181);
or U174 (N_174,In_1365,In_884);
nor U175 (N_175,In_478,In_443);
nand U176 (N_176,In_725,In_1338);
xnor U177 (N_177,In_309,In_1990);
nand U178 (N_178,In_1446,In_17);
or U179 (N_179,In_913,In_1312);
and U180 (N_180,In_646,In_196);
nand U181 (N_181,In_1711,In_1626);
xor U182 (N_182,In_145,In_324);
and U183 (N_183,In_412,In_1055);
nor U184 (N_184,In_1797,In_1101);
nor U185 (N_185,In_823,In_1095);
and U186 (N_186,In_810,In_1683);
nor U187 (N_187,In_16,In_1972);
nand U188 (N_188,In_37,In_733);
nand U189 (N_189,In_1618,In_1277);
and U190 (N_190,In_765,In_809);
and U191 (N_191,In_271,In_183);
and U192 (N_192,In_1437,In_998);
and U193 (N_193,In_433,In_1299);
nor U194 (N_194,In_1042,In_525);
nand U195 (N_195,In_1153,In_1185);
or U196 (N_196,In_1811,In_864);
nor U197 (N_197,In_1521,In_1285);
nor U198 (N_198,In_272,In_590);
and U199 (N_199,In_1006,In_658);
or U200 (N_200,In_81,In_1061);
nand U201 (N_201,In_192,In_66);
nand U202 (N_202,In_1704,In_199);
nand U203 (N_203,In_1958,In_563);
nor U204 (N_204,In_1463,In_1835);
nor U205 (N_205,In_434,In_188);
and U206 (N_206,In_578,In_420);
nor U207 (N_207,In_1541,In_703);
or U208 (N_208,In_1833,In_1942);
or U209 (N_209,In_1414,In_1474);
nor U210 (N_210,In_9,In_1943);
nand U211 (N_211,In_1759,In_612);
nand U212 (N_212,In_1155,In_1753);
and U213 (N_213,In_565,In_1660);
nand U214 (N_214,In_638,In_1123);
xnor U215 (N_215,In_720,In_351);
or U216 (N_216,In_1550,In_1817);
nor U217 (N_217,In_797,In_1968);
and U218 (N_218,In_1806,In_21);
nor U219 (N_219,In_314,In_911);
nand U220 (N_220,In_182,In_1513);
xnor U221 (N_221,In_1581,In_1117);
nor U222 (N_222,In_796,In_1852);
or U223 (N_223,In_1345,In_1448);
or U224 (N_224,In_159,In_600);
nand U225 (N_225,In_246,In_806);
xnor U226 (N_226,In_1256,In_781);
nor U227 (N_227,In_360,In_387);
and U228 (N_228,In_280,In_202);
and U229 (N_229,In_743,In_523);
and U230 (N_230,In_618,In_951);
or U231 (N_231,In_232,In_678);
or U232 (N_232,In_723,In_576);
xor U233 (N_233,In_581,In_485);
and U234 (N_234,In_1597,In_1021);
xnor U235 (N_235,In_933,In_1930);
nand U236 (N_236,In_1552,In_162);
nor U237 (N_237,In_586,In_1975);
nand U238 (N_238,In_1686,In_1695);
and U239 (N_239,In_601,In_1547);
nor U240 (N_240,In_1623,In_1418);
nor U241 (N_241,In_439,In_997);
xor U242 (N_242,In_122,In_1354);
nor U243 (N_243,In_1628,In_1570);
xor U244 (N_244,In_1984,In_1022);
nand U245 (N_245,In_1281,In_1897);
and U246 (N_246,In_928,In_986);
or U247 (N_247,In_713,In_926);
nor U248 (N_248,In_455,In_1136);
or U249 (N_249,In_473,In_486);
or U250 (N_250,In_1846,In_51);
and U251 (N_251,In_1497,In_833);
or U252 (N_252,In_1538,In_1258);
xnor U253 (N_253,In_1108,In_406);
xnor U254 (N_254,In_200,In_1625);
nor U255 (N_255,In_1784,In_1748);
nand U256 (N_256,In_990,In_1065);
nand U257 (N_257,In_252,In_1619);
or U258 (N_258,In_1156,In_1163);
nor U259 (N_259,In_1680,In_839);
and U260 (N_260,In_745,In_1566);
nand U261 (N_261,In_1295,In_1239);
or U262 (N_262,In_1573,In_189);
nor U263 (N_263,In_165,In_1037);
xor U264 (N_264,In_1428,In_379);
nor U265 (N_265,In_1067,In_1643);
nand U266 (N_266,In_33,In_330);
nand U267 (N_267,In_1212,In_1358);
or U268 (N_268,In_668,In_1648);
and U269 (N_269,In_1819,In_1131);
nor U270 (N_270,In_1433,In_764);
xnor U271 (N_271,In_1287,In_1031);
nor U272 (N_272,In_622,In_263);
nor U273 (N_273,In_298,In_149);
and U274 (N_274,In_435,In_146);
or U275 (N_275,In_1763,In_1124);
xor U276 (N_276,In_1774,In_1884);
xor U277 (N_277,In_606,In_975);
and U278 (N_278,In_961,In_1758);
nor U279 (N_279,In_344,In_1575);
and U280 (N_280,In_1887,In_1330);
nor U281 (N_281,In_1813,In_1927);
nor U282 (N_282,In_1200,In_84);
and U283 (N_283,In_619,In_135);
and U284 (N_284,In_1035,In_1262);
nor U285 (N_285,In_758,In_110);
nor U286 (N_286,In_845,In_60);
nor U287 (N_287,In_1018,In_1116);
xor U288 (N_288,In_1486,In_1732);
and U289 (N_289,In_802,In_686);
xnor U290 (N_290,In_325,In_943);
or U291 (N_291,In_140,In_1504);
nor U292 (N_292,In_1701,In_644);
nand U293 (N_293,In_1126,In_955);
and U294 (N_294,In_892,In_1786);
nand U295 (N_295,In_898,In_410);
or U296 (N_296,In_551,In_1612);
and U297 (N_297,In_973,In_1261);
or U298 (N_298,In_785,In_812);
nor U299 (N_299,In_64,In_626);
or U300 (N_300,In_979,In_495);
and U301 (N_301,In_1291,In_1011);
and U302 (N_302,In_805,In_748);
nand U303 (N_303,In_1777,In_787);
or U304 (N_304,In_333,In_871);
and U305 (N_305,In_1926,In_1783);
xnor U306 (N_306,In_1090,In_334);
or U307 (N_307,In_1546,In_1922);
or U308 (N_308,In_332,In_493);
or U309 (N_309,In_1344,In_169);
nand U310 (N_310,In_1052,In_1138);
or U311 (N_311,In_1870,In_846);
nand U312 (N_312,In_1310,In_1272);
nand U313 (N_313,In_392,In_721);
nand U314 (N_314,In_885,In_851);
nor U315 (N_315,In_391,In_1132);
nor U316 (N_316,In_331,In_1158);
nor U317 (N_317,In_1615,In_1677);
nand U318 (N_318,In_464,In_1856);
nand U319 (N_319,In_873,In_85);
nand U320 (N_320,In_1454,In_1364);
nand U321 (N_321,In_1919,In_1151);
and U322 (N_322,In_1034,In_970);
or U323 (N_323,In_989,In_401);
or U324 (N_324,In_918,In_377);
and U325 (N_325,In_118,In_693);
or U326 (N_326,In_1639,In_996);
nor U327 (N_327,In_1825,In_627);
nand U328 (N_328,In_416,In_1341);
and U329 (N_329,In_1472,In_1703);
nor U330 (N_330,In_99,In_1864);
or U331 (N_331,In_780,In_1731);
nor U332 (N_332,In_133,In_1652);
xor U333 (N_333,In_1776,In_1614);
and U334 (N_334,In_215,In_388);
nor U335 (N_335,In_1954,In_167);
xor U336 (N_336,In_510,In_782);
nor U337 (N_337,In_1630,In_463);
and U338 (N_338,In_887,In_1141);
and U339 (N_339,In_216,In_1227);
or U340 (N_340,In_437,In_1698);
or U341 (N_341,In_505,In_79);
nand U342 (N_342,In_1622,In_592);
nand U343 (N_343,In_749,In_948);
nand U344 (N_344,In_1631,In_211);
and U345 (N_345,In_908,In_3);
nor U346 (N_346,In_185,In_18);
or U347 (N_347,In_501,In_204);
and U348 (N_348,In_2,In_29);
nor U349 (N_349,In_1316,In_1716);
nor U350 (N_350,In_1308,In_1981);
or U351 (N_351,In_1511,In_657);
and U352 (N_352,In_867,In_428);
xor U353 (N_353,In_355,In_1050);
and U354 (N_354,In_82,In_1578);
nor U355 (N_355,In_1276,In_156);
nor U356 (N_356,In_1359,In_1604);
nor U357 (N_357,In_214,In_207);
and U358 (N_358,In_154,In_289);
and U359 (N_359,In_850,In_1462);
nor U360 (N_360,In_1146,In_294);
nor U361 (N_361,In_1323,In_863);
or U362 (N_362,In_1700,In_367);
xnor U363 (N_363,In_1469,In_386);
and U364 (N_364,In_1007,In_1467);
and U365 (N_365,In_322,In_1266);
or U366 (N_366,In_52,In_844);
or U367 (N_367,In_264,In_1257);
and U368 (N_368,In_984,In_1195);
or U369 (N_369,In_1438,In_381);
nor U370 (N_370,In_1214,In_681);
nor U371 (N_371,In_490,In_767);
xnor U372 (N_372,In_1821,In_402);
and U373 (N_373,In_374,In_1233);
xnor U374 (N_374,In_1331,In_556);
nor U375 (N_375,In_1746,In_203);
nand U376 (N_376,In_70,In_1304);
and U377 (N_377,In_498,In_1339);
nand U378 (N_378,In_127,In_830);
and U379 (N_379,In_469,In_126);
nor U380 (N_380,In_1815,In_317);
and U381 (N_381,In_424,In_1125);
or U382 (N_382,In_398,In_461);
or U383 (N_383,In_571,In_1500);
xnor U384 (N_384,In_980,In_136);
nor U385 (N_385,In_1871,In_31);
and U386 (N_386,In_38,In_1673);
and U387 (N_387,In_1860,In_1336);
or U388 (N_388,In_1937,In_1142);
and U389 (N_389,In_529,In_930);
nand U390 (N_390,In_39,In_134);
xor U391 (N_391,In_302,In_1656);
nand U392 (N_392,In_1723,In_1267);
and U393 (N_393,In_1442,In_1157);
and U394 (N_394,In_1997,In_1740);
nor U395 (N_395,In_819,In_1079);
or U396 (N_396,In_457,In_157);
nor U397 (N_397,In_829,In_1053);
and U398 (N_398,In_373,In_615);
nor U399 (N_399,In_260,In_1164);
nor U400 (N_400,In_1264,In_1645);
or U401 (N_401,In_151,In_481);
nor U402 (N_402,In_836,In_569);
nand U403 (N_403,In_255,In_1071);
nand U404 (N_404,In_1374,In_176);
nand U405 (N_405,In_682,In_451);
nor U406 (N_406,In_1470,In_985);
or U407 (N_407,In_1858,In_1872);
and U408 (N_408,In_1888,In_1314);
or U409 (N_409,In_649,In_1816);
nand U410 (N_410,In_1399,In_1290);
and U411 (N_411,In_247,In_1995);
and U412 (N_412,In_691,In_1691);
and U413 (N_413,In_359,In_175);
or U414 (N_414,In_1902,In_491);
nand U415 (N_415,In_801,In_872);
and U416 (N_416,In_993,In_1324);
and U417 (N_417,In_319,In_875);
nor U418 (N_418,In_1464,In_265);
xor U419 (N_419,In_105,In_515);
and U420 (N_420,In_905,In_893);
or U421 (N_421,In_1487,In_1083);
or U422 (N_422,In_1558,In_1599);
or U423 (N_423,In_171,In_1337);
and U424 (N_424,In_1976,In_574);
and U425 (N_425,In_794,In_465);
nor U426 (N_426,In_227,In_1009);
and U427 (N_427,In_1326,In_747);
nor U428 (N_428,In_1796,In_1001);
and U429 (N_429,In_564,In_716);
nor U430 (N_430,In_883,In_1885);
nor U431 (N_431,In_874,In_798);
nor U432 (N_432,In_143,In_1135);
or U433 (N_433,In_593,In_1174);
or U434 (N_434,In_1880,In_1674);
xor U435 (N_435,In_629,In_768);
or U436 (N_436,In_1045,In_1147);
or U437 (N_437,In_937,In_1914);
nand U438 (N_438,In_1317,In_1620);
xor U439 (N_439,In_909,In_1057);
nor U440 (N_440,In_1663,In_672);
or U441 (N_441,In_349,In_1184);
and U442 (N_442,In_1043,In_1186);
nand U443 (N_443,In_1062,In_814);
or U444 (N_444,In_1729,In_346);
or U445 (N_445,In_936,In_1685);
or U446 (N_446,In_1038,In_552);
nand U447 (N_447,In_825,In_1853);
nor U448 (N_448,In_372,In_297);
nor U449 (N_449,In_369,In_1843);
nor U450 (N_450,In_910,In_897);
or U451 (N_451,In_774,In_438);
nor U452 (N_452,In_1420,In_1466);
xnor U453 (N_453,In_1781,In_1115);
and U454 (N_454,In_579,In_1012);
and U455 (N_455,In_1974,In_1353);
nand U456 (N_456,In_243,In_1385);
or U457 (N_457,In_804,In_532);
and U458 (N_458,In_361,In_1702);
and U459 (N_459,In_59,In_1523);
xor U460 (N_460,In_942,In_1693);
xnor U461 (N_461,In_1542,In_882);
and U462 (N_462,In_1225,In_621);
nor U463 (N_463,In_634,In_94);
nor U464 (N_464,In_394,In_1669);
and U465 (N_465,In_1313,In_561);
or U466 (N_466,In_1411,In_1553);
or U467 (N_467,In_1910,In_400);
and U468 (N_468,In_962,In_1190);
nor U469 (N_469,In_759,In_14);
nand U470 (N_470,In_1726,In_1983);
nor U471 (N_471,In_504,In_160);
and U472 (N_472,In_640,In_1100);
and U473 (N_473,In_924,In_762);
or U474 (N_474,In_944,In_981);
nor U475 (N_475,In_821,In_912);
nor U476 (N_476,In_1555,In_971);
or U477 (N_477,In_1952,In_611);
nor U478 (N_478,In_396,In_1059);
nor U479 (N_479,In_1004,In_1165);
nand U480 (N_480,In_1810,In_1953);
or U481 (N_481,In_1861,In_1412);
nand U482 (N_482,In_868,In_452);
nand U483 (N_483,In_1627,In_1960);
nor U484 (N_484,In_307,In_1621);
and U485 (N_485,In_522,In_1592);
xor U486 (N_486,In_1005,In_940);
and U487 (N_487,In_1237,In_1386);
or U488 (N_488,In_1213,In_1202);
nor U489 (N_489,In_1706,In_234);
xor U490 (N_490,In_958,In_445);
nor U491 (N_491,In_533,In_1761);
nand U492 (N_492,In_1516,In_753);
and U493 (N_493,In_376,In_286);
xor U494 (N_494,In_1249,In_876);
nand U495 (N_495,In_166,In_1073);
or U496 (N_496,In_89,In_1531);
or U497 (N_497,In_604,In_466);
nor U498 (N_498,In_88,In_109);
nand U499 (N_499,In_1788,In_1562);
and U500 (N_500,In_1127,In_1644);
nor U501 (N_501,In_91,In_1561);
xnor U502 (N_502,In_949,In_240);
or U503 (N_503,In_1120,In_1329);
nand U504 (N_504,In_1519,In_1525);
nand U505 (N_505,In_1439,In_673);
xor U506 (N_506,In_267,In_432);
xnor U507 (N_507,In_1077,In_1368);
or U508 (N_508,In_312,In_1598);
or U509 (N_509,In_1492,In_409);
nand U510 (N_510,In_1898,In_43);
xor U511 (N_511,In_173,In_1718);
and U512 (N_512,In_348,In_1657);
or U513 (N_513,In_775,In_1097);
and U514 (N_514,In_1205,In_299);
nand U515 (N_515,In_791,In_1133);
nor U516 (N_516,In_1294,In_1085);
or U517 (N_517,In_1283,In_828);
and U518 (N_518,In_711,In_1207);
or U519 (N_519,In_1875,In_11);
nand U520 (N_520,In_952,In_1445);
nand U521 (N_521,In_393,In_795);
nand U522 (N_522,In_1372,In_1795);
nand U523 (N_523,In_32,In_1391);
nor U524 (N_524,In_1300,In_1637);
and U525 (N_525,In_727,In_193);
and U526 (N_526,In_1571,In_648);
or U527 (N_527,In_462,In_1128);
nor U528 (N_528,In_705,In_1167);
nand U529 (N_529,In_1595,In_1026);
nand U530 (N_530,In_174,In_1370);
or U531 (N_531,In_1678,In_1030);
or U532 (N_532,In_1530,In_1569);
and U533 (N_533,In_1242,In_562);
nor U534 (N_534,In_1505,In_1883);
or U535 (N_535,In_1915,In_609);
nand U536 (N_536,In_1394,In_1600);
xnor U537 (N_537,In_1951,In_1443);
xor U538 (N_538,In_835,In_901);
nand U539 (N_539,In_356,In_116);
nand U540 (N_540,In_1000,In_1144);
and U541 (N_541,In_1407,In_378);
and U542 (N_542,In_1268,In_93);
or U543 (N_543,In_1682,In_667);
nand U544 (N_544,In_1425,In_1785);
and U545 (N_545,In_1089,In_1072);
or U546 (N_546,In_1199,In_257);
nand U547 (N_547,In_362,In_1613);
and U548 (N_548,In_878,In_281);
or U549 (N_549,In_655,In_722);
and U550 (N_550,In_1563,In_221);
nor U551 (N_551,In_100,In_338);
nor U552 (N_552,In_554,In_1098);
and U553 (N_553,In_1985,In_580);
xor U554 (N_554,In_1899,In_894);
nand U555 (N_555,In_55,In_112);
nand U556 (N_556,In_1223,In_1070);
and U557 (N_557,In_1286,In_1398);
or U558 (N_558,In_1565,In_843);
nand U559 (N_559,In_1624,In_235);
nand U560 (N_560,In_1387,In_1475);
and U561 (N_561,In_1966,In_1536);
nor U562 (N_562,In_739,In_1651);
and U563 (N_563,In_78,In_357);
nand U564 (N_564,In_521,In_588);
and U565 (N_565,In_228,In_12);
or U566 (N_566,In_855,In_217);
nor U567 (N_567,In_630,In_1794);
or U568 (N_568,In_1991,In_1148);
or U569 (N_569,In_1096,In_158);
or U570 (N_570,In_519,In_1434);
and U571 (N_571,In_669,In_287);
and U572 (N_572,In_71,In_1818);
and U573 (N_573,In_1724,In_1641);
or U574 (N_574,In_1518,In_832);
nand U575 (N_575,In_1549,In_1461);
nor U576 (N_576,In_717,In_1435);
nor U577 (N_577,In_1534,In_527);
nor U578 (N_578,In_1901,In_1842);
xor U579 (N_579,In_857,In_1211);
nand U580 (N_580,In_128,In_572);
or U581 (N_581,In_489,In_756);
nor U582 (N_582,In_1929,In_1023);
or U583 (N_583,In_956,In_1585);
or U584 (N_584,In_1931,In_1662);
and U585 (N_585,In_1054,In_1245);
nor U586 (N_586,In_1088,In_891);
and U587 (N_587,In_947,In_250);
or U588 (N_588,In_96,In_1340);
or U589 (N_589,In_1863,In_639);
xnor U590 (N_590,In_1405,In_375);
nor U591 (N_591,In_1274,In_1841);
nor U592 (N_592,In_1529,In_328);
nor U593 (N_593,In_380,In_799);
nand U594 (N_594,In_853,In_57);
nor U595 (N_595,In_1191,In_1509);
and U596 (N_596,In_1139,In_1404);
or U597 (N_597,In_1996,In_24);
nand U598 (N_598,In_142,In_1906);
or U599 (N_599,In_1532,In_1916);
nor U600 (N_600,In_1749,In_363);
nand U601 (N_601,In_1709,In_1771);
and U602 (N_602,In_1979,In_186);
or U603 (N_603,In_1122,In_907);
nand U604 (N_604,In_922,In_1909);
or U605 (N_605,In_929,In_40);
or U606 (N_606,In_1333,In_1862);
xor U607 (N_607,In_591,In_1940);
nor U608 (N_608,In_1679,In_1699);
nor U609 (N_609,In_1150,In_450);
and U610 (N_610,In_219,In_1765);
or U611 (N_611,In_198,In_358);
and U612 (N_612,In_1393,In_995);
nand U613 (N_613,In_368,In_1988);
nand U614 (N_614,In_932,In_896);
and U615 (N_615,In_1289,In_1567);
nand U616 (N_616,In_915,In_1243);
and U617 (N_617,In_624,In_460);
nand U618 (N_618,In_1998,In_471);
and U619 (N_619,In_1453,In_1993);
nor U620 (N_620,In_365,In_1801);
nand U621 (N_621,In_80,In_671);
nand U622 (N_622,In_1684,In_1217);
nand U623 (N_623,In_1659,In_1255);
nand U624 (N_624,In_125,In_1543);
and U625 (N_625,In_408,In_482);
and U626 (N_626,In_1583,In_608);
nand U627 (N_627,In_1839,In_766);
or U628 (N_628,In_770,In_120);
nor U629 (N_629,In_447,In_620);
nand U630 (N_630,In_1665,In_45);
nor U631 (N_631,In_610,In_1459);
nor U632 (N_632,In_685,In_1430);
and U633 (N_633,In_506,In_1579);
or U634 (N_634,In_205,In_1939);
xnor U635 (N_635,In_1676,In_83);
nand U636 (N_636,In_479,In_1965);
or U637 (N_637,In_27,In_1501);
and U638 (N_638,In_1447,In_350);
and U639 (N_639,In_72,In_637);
or U640 (N_640,In_172,In_170);
and U641 (N_641,In_582,In_1490);
or U642 (N_642,In_1840,In_1403);
and U643 (N_643,In_34,In_1629);
and U644 (N_644,In_1415,In_1113);
nand U645 (N_645,In_744,In_1714);
nor U646 (N_646,In_1649,In_233);
or U647 (N_647,In_518,In_335);
nand U648 (N_648,In_1209,In_1413);
nor U649 (N_649,In_1634,In_889);
nor U650 (N_650,In_650,In_1750);
or U651 (N_651,In_1889,In_702);
xor U652 (N_652,In_599,In_847);
nor U653 (N_653,In_595,In_1792);
or U654 (N_654,In_305,In_792);
and U655 (N_655,In_477,In_385);
nor U656 (N_656,In_1253,In_1928);
or U657 (N_657,In_114,In_1934);
xor U658 (N_658,In_803,In_750);
and U659 (N_659,In_1973,In_1933);
nand U660 (N_660,In_1121,In_585);
nor U661 (N_661,In_1247,In_1587);
nand U662 (N_662,In_1204,In_1048);
and U663 (N_663,In_1260,In_888);
and U664 (N_664,In_1917,In_773);
nand U665 (N_665,In_1468,In_1254);
nand U666 (N_666,In_1485,In_824);
nor U667 (N_667,In_87,In_1670);
and U668 (N_668,In_1768,In_862);
nor U669 (N_669,In_680,In_1877);
nor U670 (N_670,In_1607,In_738);
nor U671 (N_671,In_1376,In_1328);
or U672 (N_672,In_1950,In_1850);
nand U673 (N_673,In_1514,In_292);
nor U674 (N_674,In_1406,In_178);
nor U675 (N_675,In_1311,In_342);
and U676 (N_676,In_1441,In_917);
and U677 (N_677,In_1160,In_1401);
or U678 (N_678,In_119,In_904);
nand U679 (N_679,In_1847,In_197);
xor U680 (N_680,In_138,In_107);
and U681 (N_681,In_476,In_1236);
and U682 (N_682,In_1465,In_441);
nor U683 (N_683,In_277,In_179);
nor U684 (N_684,In_935,In_1106);
nand U685 (N_685,In_1327,In_959);
nor U686 (N_686,In_632,In_1367);
nor U687 (N_687,In_1664,In_26);
nand U688 (N_688,In_1332,In_1028);
and U689 (N_689,In_1946,In_67);
nor U690 (N_690,In_659,In_194);
xor U691 (N_691,In_1540,In_695);
or U692 (N_692,In_467,In_1609);
nor U693 (N_693,In_520,In_269);
nor U694 (N_694,In_1738,In_859);
nand U695 (N_695,In_488,In_837);
xnor U696 (N_696,In_849,In_536);
or U697 (N_697,In_1874,In_213);
nor U698 (N_698,In_1799,In_1349);
nand U699 (N_699,In_1911,In_1616);
or U700 (N_700,In_1484,In_1596);
or U701 (N_701,In_1343,In_1238);
nor U702 (N_702,In_1800,In_1248);
or U703 (N_703,In_1721,In_58);
and U704 (N_704,In_793,In_1945);
nor U705 (N_705,In_651,In_1168);
nand U706 (N_706,In_869,In_1739);
nor U707 (N_707,In_1279,In_251);
nor U708 (N_708,In_757,In_616);
nor U709 (N_709,In_1524,In_139);
nor U710 (N_710,In_425,In_541);
xnor U711 (N_711,In_1736,In_310);
nand U712 (N_712,In_1208,In_384);
and U713 (N_713,In_1590,In_1805);
and U714 (N_714,In_1455,In_1019);
or U715 (N_715,In_1636,In_709);
nor U716 (N_716,In_1956,In_1179);
nand U717 (N_717,In_472,In_1373);
nand U718 (N_718,In_1014,In_1112);
nand U719 (N_719,In_701,In_1109);
xnor U720 (N_720,In_1725,In_288);
nand U721 (N_721,In_1408,In_1719);
nand U722 (N_722,In_1218,In_245);
xnor U723 (N_723,In_1866,In_1058);
nor U724 (N_724,In_48,In_284);
nor U725 (N_725,In_1712,In_1826);
or U726 (N_726,In_1827,In_1690);
and U727 (N_727,In_1152,In_1878);
xnor U728 (N_728,In_1557,In_1369);
nor U729 (N_729,In_1791,In_283);
and U730 (N_730,In_1176,In_919);
xnor U731 (N_731,In_1222,In_1451);
or U732 (N_732,In_1180,In_628);
nor U733 (N_733,In_613,In_1388);
and U734 (N_734,In_407,In_236);
or U735 (N_735,In_249,In_276);
or U736 (N_736,In_1137,In_1457);
xor U737 (N_737,In_1377,In_1868);
xnor U738 (N_738,In_448,In_1751);
or U739 (N_739,In_1081,In_1259);
nor U740 (N_740,In_1269,In_1170);
or U741 (N_741,In_1881,In_1789);
and U742 (N_742,In_1779,In_1194);
and U743 (N_743,In_1822,In_1040);
nand U744 (N_744,In_459,In_726);
or U745 (N_745,In_1893,In_1895);
and U746 (N_746,In_1526,In_820);
and U747 (N_747,In_7,In_35);
and U748 (N_748,In_661,In_1424);
nand U749 (N_749,In_1322,In_301);
and U750 (N_750,In_1844,In_740);
xnor U751 (N_751,In_1149,In_291);
nor U752 (N_752,In_854,In_558);
nand U753 (N_753,In_526,In_1228);
xor U754 (N_754,In_1762,In_1896);
nand U755 (N_755,In_1235,In_1766);
nor U756 (N_756,In_1551,In_1572);
and U757 (N_757,In_1672,In_865);
and U758 (N_758,In_321,In_1192);
nor U759 (N_759,In_1173,In_1808);
or U760 (N_760,In_736,In_279);
xnor U761 (N_761,In_969,In_278);
nand U762 (N_762,In_1591,In_1110);
or U763 (N_763,In_123,In_1635);
nand U764 (N_764,In_545,In_454);
and U765 (N_765,In_210,In_106);
nor U766 (N_766,In_900,In_75);
nand U767 (N_767,In_584,In_1426);
nor U768 (N_768,In_209,In_772);
and U769 (N_769,In_1201,In_1350);
or U770 (N_770,In_1390,In_1925);
nand U771 (N_771,In_742,In_786);
nor U772 (N_772,In_1134,In_808);
and U773 (N_773,In_788,In_1601);
nor U774 (N_774,In_737,In_238);
nor U775 (N_775,In_870,In_665);
nand U776 (N_776,In_557,In_108);
or U777 (N_777,In_1431,In_1809);
nor U778 (N_778,In_860,In_1084);
nand U779 (N_779,In_1402,In_856);
xor U780 (N_780,In_662,In_1924);
or U781 (N_781,In_1473,In_1423);
nand U782 (N_782,In_594,In_1692);
nand U783 (N_783,In_1382,In_25);
or U784 (N_784,In_920,In_1075);
nand U785 (N_785,In_1066,In_1198);
or U786 (N_786,In_838,In_983);
and U787 (N_787,In_999,In_1488);
or U788 (N_788,In_1280,In_880);
nor U789 (N_789,In_231,In_44);
and U790 (N_790,In_1707,In_982);
or U791 (N_791,In_688,In_1986);
and U792 (N_792,In_1068,In_1495);
nand U793 (N_793,In_953,In_187);
and U794 (N_794,In_1017,In_1159);
and U795 (N_795,In_1111,In_1787);
nor U796 (N_796,In_77,In_931);
and U797 (N_797,In_719,In_954);
nor U798 (N_798,In_440,In_1477);
or U799 (N_799,In_1301,In_86);
and U800 (N_800,In_1824,In_1381);
and U801 (N_801,In_131,In_1851);
nand U802 (N_802,In_337,In_938);
and U803 (N_803,In_266,In_1060);
nand U804 (N_804,In_1747,In_274);
nor U805 (N_805,In_1912,In_1535);
and U806 (N_806,In_879,In_5);
and U807 (N_807,In_528,In_623);
nand U808 (N_808,In_1171,In_429);
or U809 (N_809,In_500,In_1380);
nand U810 (N_810,In_311,In_242);
or U811 (N_811,In_852,In_1905);
nand U812 (N_812,In_285,In_728);
nand U813 (N_813,In_674,In_939);
nand U814 (N_814,In_475,In_446);
or U815 (N_815,In_1044,In_1633);
nor U816 (N_816,In_1537,In_177);
nor U817 (N_817,In_23,In_789);
nor U818 (N_818,In_1814,In_508);
or U819 (N_819,In_1188,In_229);
nand U820 (N_820,In_752,In_1091);
and U821 (N_821,In_201,In_1873);
nand U822 (N_822,In_241,In_353);
or U823 (N_823,In_1356,In_1770);
or U824 (N_824,In_663,In_1175);
nor U825 (N_825,In_706,In_509);
and U826 (N_826,In_696,In_1187);
or U827 (N_827,In_1056,In_906);
or U828 (N_828,In_1992,In_1832);
or U829 (N_829,In_499,In_62);
and U830 (N_830,In_46,In_1362);
nand U831 (N_831,In_1008,In_1396);
nor U832 (N_832,In_963,In_1527);
nor U833 (N_833,In_413,In_1094);
xor U834 (N_834,In_656,In_0);
nor U835 (N_835,In_1193,In_1671);
nand U836 (N_836,In_921,In_73);
nor U837 (N_837,In_1586,In_968);
xor U838 (N_838,In_1891,In_1640);
nand U839 (N_839,In_934,In_225);
and U840 (N_840,In_90,In_244);
and U841 (N_841,In_290,In_1241);
nor U842 (N_842,In_614,In_577);
and U843 (N_843,In_1838,In_50);
nor U844 (N_844,In_65,In_502);
nor U845 (N_845,In_483,In_230);
or U846 (N_846,In_1320,In_596);
nor U847 (N_847,In_1667,In_1886);
or U848 (N_848,In_347,In_1589);
nand U849 (N_849,In_1632,In_54);
nand U850 (N_850,In_320,In_1355);
or U851 (N_851,In_208,In_1013);
nand U852 (N_852,In_1307,In_370);
and U853 (N_853,In_1270,In_976);
nor U854 (N_854,In_704,In_30);
nor U855 (N_855,In_1357,In_470);
and U856 (N_856,In_1967,In_113);
xnor U857 (N_857,In_1400,In_560);
and U858 (N_858,In_1802,In_988);
nand U859 (N_859,In_414,In_1638);
and U860 (N_860,In_1568,In_1039);
and U861 (N_861,In_8,In_831);
nor U862 (N_862,In_1416,In_121);
and U863 (N_863,In_296,In_97);
or U864 (N_864,In_1944,In_550);
or U865 (N_865,In_670,In_538);
nand U866 (N_866,In_1820,In_1756);
xor U867 (N_867,In_553,In_1027);
nand U868 (N_868,In_1002,In_1971);
xnor U869 (N_869,In_848,In_1755);
or U870 (N_870,In_47,In_1107);
nand U871 (N_871,In_1480,In_1582);
nor U872 (N_872,In_1735,In_813);
xnor U873 (N_873,In_689,In_1772);
or U874 (N_874,In_1024,In_539);
or U875 (N_875,In_1867,In_137);
or U876 (N_876,In_555,In_531);
nor U877 (N_877,In_1069,In_1941);
or U878 (N_878,In_602,In_300);
and U879 (N_879,In_1689,In_1483);
nand U880 (N_880,In_4,In_543);
nor U881 (N_881,In_275,In_1502);
or U882 (N_882,In_1742,In_1216);
and U883 (N_883,In_1713,In_1957);
nor U884 (N_884,In_653,In_153);
or U885 (N_885,In_568,In_237);
and U886 (N_886,In_1429,In_822);
or U887 (N_887,In_625,In_1417);
or U888 (N_888,In_315,In_1093);
and U889 (N_889,In_389,In_1496);
nand U890 (N_890,In_914,In_323);
nand U891 (N_891,In_776,In_1169);
nand U892 (N_892,In_1708,In_566);
nor U893 (N_893,In_1145,In_1297);
and U894 (N_894,In_645,In_967);
nand U895 (N_895,In_293,In_308);
nand U896 (N_896,In_977,In_1203);
or U897 (N_897,In_68,In_573);
nand U898 (N_898,In_652,In_1246);
nand U899 (N_899,In_916,In_1206);
nand U900 (N_900,In_1064,In_724);
xnor U901 (N_901,In_152,In_978);
nand U902 (N_902,In_1251,In_1666);
and U903 (N_903,In_1694,In_1503);
nand U904 (N_904,In_364,In_1325);
and U905 (N_905,In_1605,In_124);
and U906 (N_906,In_421,In_790);
nor U907 (N_907,In_53,In_1921);
and U908 (N_908,In_1980,In_453);
nor U909 (N_909,In_1829,In_1293);
nor U910 (N_910,In_1688,In_761);
nor U911 (N_911,In_1999,In_74);
nand U912 (N_912,In_1773,In_132);
nand U913 (N_913,In_1278,In_1653);
xor U914 (N_914,In_834,In_1016);
and U915 (N_915,In_382,In_1730);
nand U916 (N_916,In_418,In_575);
nand U917 (N_917,In_104,In_1319);
or U918 (N_918,In_570,In_1118);
nand U919 (N_919,In_212,In_827);
nand U920 (N_920,In_220,In_708);
nand U921 (N_921,In_1548,In_534);
and U922 (N_922,In_419,In_1010);
or U923 (N_923,In_492,In_1306);
nand U924 (N_924,In_262,In_732);
and U925 (N_925,In_1646,In_258);
and U926 (N_926,In_1275,In_1720);
nand U927 (N_927,In_1471,In_1086);
or U928 (N_928,In_1855,In_1305);
nor U929 (N_929,In_540,In_683);
nor U930 (N_930,In_1961,In_474);
nor U931 (N_931,In_1105,In_184);
or U932 (N_932,In_354,In_1857);
or U933 (N_933,In_1611,In_13);
nand U934 (N_934,In_1063,In_1197);
and U935 (N_935,In_1559,In_1315);
xor U936 (N_936,In_248,In_729);
or U937 (N_937,In_316,In_1087);
nand U938 (N_938,In_190,In_1003);
nor U939 (N_939,In_42,In_15);
or U940 (N_940,In_1347,In_1854);
and U941 (N_941,In_589,In_567);
or U942 (N_942,In_1231,In_1775);
nor U943 (N_943,In_769,In_1515);
and U944 (N_944,In_117,In_927);
nor U945 (N_945,In_1397,In_1642);
nand U946 (N_946,In_1378,In_1240);
and U947 (N_947,In_1210,In_1440);
or U948 (N_948,In_1410,In_1335);
nand U949 (N_949,In_1478,In_1161);
nand U950 (N_950,In_1903,In_1831);
or U951 (N_951,In_1288,In_163);
xnor U952 (N_952,In_1032,In_1129);
nand U953 (N_953,In_226,In_731);
nor U954 (N_954,In_1545,In_103);
xnor U955 (N_955,In_715,In_537);
or U956 (N_956,In_1948,In_1104);
nor U957 (N_957,In_261,In_1302);
nor U958 (N_958,In_957,In_1080);
nand U959 (N_959,In_191,In_925);
or U960 (N_960,In_1074,In_395);
xnor U961 (N_961,In_1460,In_1734);
nand U962 (N_962,In_1603,In_1215);
and U963 (N_963,In_763,In_746);
or U964 (N_964,In_1029,In_877);
nor U965 (N_965,In_1584,In_92);
nand U966 (N_966,In_1506,In_1375);
xor U967 (N_967,In_1481,In_1977);
nand U968 (N_968,In_1962,In_1444);
nand U969 (N_969,In_1752,In_1499);
and U970 (N_970,In_1025,In_807);
and U971 (N_971,In_946,In_1076);
xor U972 (N_972,In_426,In_1760);
nand U973 (N_973,In_617,In_1936);
nand U974 (N_974,In_1342,In_548);
xor U975 (N_975,In_69,In_456);
xnor U976 (N_976,In_1668,In_654);
nor U977 (N_977,In_345,In_1033);
xor U978 (N_978,In_643,In_1837);
and U979 (N_979,In_559,In_1681);
and U980 (N_980,In_436,In_343);
and U981 (N_981,In_1544,In_415);
and U982 (N_982,In_150,In_1421);
nand U983 (N_983,In_313,In_730);
or U984 (N_984,In_1588,In_1092);
nor U985 (N_985,In_1383,In_63);
or U986 (N_986,In_598,In_1782);
or U987 (N_987,In_513,In_941);
nand U988 (N_988,In_1737,In_1982);
or U989 (N_989,In_1907,In_530);
xor U990 (N_990,In_224,In_1102);
nand U991 (N_991,In_1970,In_664);
and U992 (N_992,In_1520,In_1119);
nand U993 (N_993,In_206,In_1859);
xnor U994 (N_994,In_1183,In_253);
nor U995 (N_995,In_966,In_779);
nor U996 (N_996,In_144,In_699);
or U997 (N_997,In_698,In_1743);
and U998 (N_998,In_1882,In_1959);
and U999 (N_999,In_1675,In_19);
nand U1000 (N_1000,In_1165,In_571);
and U1001 (N_1001,In_1907,In_1638);
nor U1002 (N_1002,In_1059,In_684);
and U1003 (N_1003,In_1479,In_1736);
xor U1004 (N_1004,In_931,In_1268);
and U1005 (N_1005,In_1884,In_829);
nand U1006 (N_1006,In_861,In_767);
nand U1007 (N_1007,In_552,In_1981);
and U1008 (N_1008,In_1019,In_672);
xnor U1009 (N_1009,In_1868,In_1391);
and U1010 (N_1010,In_1984,In_227);
and U1011 (N_1011,In_800,In_1269);
or U1012 (N_1012,In_1313,In_789);
xor U1013 (N_1013,In_887,In_1486);
and U1014 (N_1014,In_776,In_158);
or U1015 (N_1015,In_369,In_121);
or U1016 (N_1016,In_770,In_1999);
nand U1017 (N_1017,In_1705,In_1956);
nand U1018 (N_1018,In_1069,In_1153);
nor U1019 (N_1019,In_1419,In_1519);
or U1020 (N_1020,In_137,In_1813);
nand U1021 (N_1021,In_485,In_702);
and U1022 (N_1022,In_199,In_1744);
xnor U1023 (N_1023,In_438,In_1586);
nor U1024 (N_1024,In_1471,In_1772);
and U1025 (N_1025,In_1367,In_1713);
and U1026 (N_1026,In_1919,In_958);
nand U1027 (N_1027,In_655,In_643);
nand U1028 (N_1028,In_427,In_991);
nand U1029 (N_1029,In_1657,In_703);
nor U1030 (N_1030,In_1028,In_1636);
xor U1031 (N_1031,In_1986,In_1308);
nor U1032 (N_1032,In_406,In_71);
and U1033 (N_1033,In_1362,In_1379);
or U1034 (N_1034,In_1481,In_385);
or U1035 (N_1035,In_1721,In_1237);
nor U1036 (N_1036,In_1123,In_109);
or U1037 (N_1037,In_1975,In_998);
and U1038 (N_1038,In_961,In_3);
nand U1039 (N_1039,In_1411,In_292);
and U1040 (N_1040,In_977,In_429);
or U1041 (N_1041,In_597,In_1659);
xnor U1042 (N_1042,In_1126,In_890);
nor U1043 (N_1043,In_1511,In_668);
xor U1044 (N_1044,In_1630,In_941);
nor U1045 (N_1045,In_1201,In_478);
and U1046 (N_1046,In_683,In_879);
nand U1047 (N_1047,In_1760,In_1728);
and U1048 (N_1048,In_1569,In_376);
or U1049 (N_1049,In_1574,In_227);
or U1050 (N_1050,In_545,In_770);
nand U1051 (N_1051,In_80,In_1601);
nor U1052 (N_1052,In_1323,In_647);
nor U1053 (N_1053,In_1277,In_141);
or U1054 (N_1054,In_531,In_327);
and U1055 (N_1055,In_1142,In_1957);
nand U1056 (N_1056,In_1681,In_1224);
nor U1057 (N_1057,In_819,In_1409);
xor U1058 (N_1058,In_1635,In_121);
and U1059 (N_1059,In_1746,In_1205);
nand U1060 (N_1060,In_1187,In_1474);
and U1061 (N_1061,In_297,In_681);
and U1062 (N_1062,In_1245,In_465);
nor U1063 (N_1063,In_548,In_532);
or U1064 (N_1064,In_1083,In_888);
and U1065 (N_1065,In_462,In_562);
nor U1066 (N_1066,In_1757,In_1844);
or U1067 (N_1067,In_839,In_1302);
nand U1068 (N_1068,In_1321,In_1557);
nand U1069 (N_1069,In_1081,In_17);
or U1070 (N_1070,In_1446,In_745);
nand U1071 (N_1071,In_924,In_30);
and U1072 (N_1072,In_21,In_703);
nor U1073 (N_1073,In_1232,In_495);
or U1074 (N_1074,In_1878,In_127);
nand U1075 (N_1075,In_1760,In_1192);
nand U1076 (N_1076,In_748,In_1054);
or U1077 (N_1077,In_1269,In_1651);
nand U1078 (N_1078,In_1945,In_1241);
and U1079 (N_1079,In_1546,In_1126);
or U1080 (N_1080,In_324,In_587);
nor U1081 (N_1081,In_1384,In_159);
and U1082 (N_1082,In_553,In_121);
nor U1083 (N_1083,In_950,In_834);
and U1084 (N_1084,In_1389,In_272);
or U1085 (N_1085,In_788,In_1941);
and U1086 (N_1086,In_241,In_631);
nor U1087 (N_1087,In_327,In_1144);
or U1088 (N_1088,In_543,In_1772);
nor U1089 (N_1089,In_320,In_1565);
nand U1090 (N_1090,In_228,In_1309);
nor U1091 (N_1091,In_196,In_1344);
and U1092 (N_1092,In_1855,In_1019);
xor U1093 (N_1093,In_1345,In_551);
nor U1094 (N_1094,In_1570,In_965);
xor U1095 (N_1095,In_1080,In_1726);
and U1096 (N_1096,In_1948,In_336);
nor U1097 (N_1097,In_1910,In_1333);
or U1098 (N_1098,In_898,In_359);
and U1099 (N_1099,In_1333,In_1441);
or U1100 (N_1100,In_1808,In_1901);
and U1101 (N_1101,In_1902,In_591);
nor U1102 (N_1102,In_453,In_231);
xor U1103 (N_1103,In_854,In_374);
nand U1104 (N_1104,In_1732,In_1995);
or U1105 (N_1105,In_1571,In_1137);
nand U1106 (N_1106,In_510,In_1385);
or U1107 (N_1107,In_1586,In_1490);
or U1108 (N_1108,In_570,In_240);
or U1109 (N_1109,In_1256,In_119);
or U1110 (N_1110,In_87,In_1922);
nor U1111 (N_1111,In_652,In_1978);
or U1112 (N_1112,In_1978,In_746);
and U1113 (N_1113,In_1951,In_81);
and U1114 (N_1114,In_1880,In_134);
and U1115 (N_1115,In_1630,In_1293);
or U1116 (N_1116,In_1440,In_1511);
nand U1117 (N_1117,In_388,In_468);
and U1118 (N_1118,In_1626,In_185);
nor U1119 (N_1119,In_1847,In_257);
and U1120 (N_1120,In_1732,In_1027);
and U1121 (N_1121,In_73,In_1652);
or U1122 (N_1122,In_489,In_146);
nand U1123 (N_1123,In_852,In_380);
xor U1124 (N_1124,In_231,In_1493);
nand U1125 (N_1125,In_1103,In_344);
or U1126 (N_1126,In_1576,In_406);
or U1127 (N_1127,In_1307,In_841);
xnor U1128 (N_1128,In_1454,In_194);
or U1129 (N_1129,In_1735,In_848);
nand U1130 (N_1130,In_1996,In_1253);
and U1131 (N_1131,In_127,In_90);
xor U1132 (N_1132,In_1814,In_315);
xor U1133 (N_1133,In_1706,In_1281);
nor U1134 (N_1134,In_1474,In_1289);
nor U1135 (N_1135,In_109,In_763);
and U1136 (N_1136,In_973,In_1043);
nor U1137 (N_1137,In_394,In_428);
or U1138 (N_1138,In_644,In_820);
or U1139 (N_1139,In_1509,In_323);
xnor U1140 (N_1140,In_1066,In_1274);
or U1141 (N_1141,In_1553,In_1694);
or U1142 (N_1142,In_1496,In_797);
nor U1143 (N_1143,In_1689,In_490);
xor U1144 (N_1144,In_724,In_358);
nand U1145 (N_1145,In_728,In_1441);
and U1146 (N_1146,In_1734,In_831);
nor U1147 (N_1147,In_1536,In_1940);
xor U1148 (N_1148,In_135,In_1702);
and U1149 (N_1149,In_446,In_439);
or U1150 (N_1150,In_1640,In_356);
nand U1151 (N_1151,In_463,In_1678);
nor U1152 (N_1152,In_805,In_16);
nor U1153 (N_1153,In_1374,In_438);
and U1154 (N_1154,In_1709,In_911);
and U1155 (N_1155,In_90,In_1750);
and U1156 (N_1156,In_916,In_44);
and U1157 (N_1157,In_140,In_120);
or U1158 (N_1158,In_807,In_153);
and U1159 (N_1159,In_128,In_217);
or U1160 (N_1160,In_1089,In_74);
nand U1161 (N_1161,In_700,In_347);
and U1162 (N_1162,In_1105,In_383);
nand U1163 (N_1163,In_1513,In_701);
xor U1164 (N_1164,In_922,In_255);
or U1165 (N_1165,In_1694,In_685);
and U1166 (N_1166,In_1843,In_630);
xor U1167 (N_1167,In_589,In_1143);
nor U1168 (N_1168,In_1106,In_1934);
xnor U1169 (N_1169,In_1476,In_1426);
nand U1170 (N_1170,In_1339,In_757);
or U1171 (N_1171,In_1331,In_709);
or U1172 (N_1172,In_703,In_247);
xnor U1173 (N_1173,In_839,In_1947);
nand U1174 (N_1174,In_150,In_1677);
nand U1175 (N_1175,In_33,In_1152);
nand U1176 (N_1176,In_298,In_189);
nor U1177 (N_1177,In_1720,In_1938);
xor U1178 (N_1178,In_498,In_1396);
nor U1179 (N_1179,In_1460,In_1466);
or U1180 (N_1180,In_459,In_834);
nand U1181 (N_1181,In_1481,In_739);
nor U1182 (N_1182,In_1892,In_1937);
nor U1183 (N_1183,In_1169,In_1576);
or U1184 (N_1184,In_1171,In_1518);
nor U1185 (N_1185,In_792,In_1298);
and U1186 (N_1186,In_1979,In_1950);
or U1187 (N_1187,In_1453,In_1549);
or U1188 (N_1188,In_653,In_516);
nand U1189 (N_1189,In_1597,In_1427);
or U1190 (N_1190,In_1160,In_1226);
nor U1191 (N_1191,In_549,In_1380);
xor U1192 (N_1192,In_630,In_1750);
nand U1193 (N_1193,In_1902,In_539);
and U1194 (N_1194,In_881,In_757);
nand U1195 (N_1195,In_1467,In_1468);
nor U1196 (N_1196,In_939,In_1439);
nand U1197 (N_1197,In_315,In_55);
nand U1198 (N_1198,In_669,In_1909);
nand U1199 (N_1199,In_1390,In_593);
nor U1200 (N_1200,In_1010,In_677);
nor U1201 (N_1201,In_1832,In_1522);
or U1202 (N_1202,In_1589,In_180);
or U1203 (N_1203,In_583,In_1559);
nand U1204 (N_1204,In_1084,In_700);
nand U1205 (N_1205,In_1154,In_35);
nand U1206 (N_1206,In_1721,In_1048);
or U1207 (N_1207,In_1570,In_1554);
or U1208 (N_1208,In_1807,In_1374);
or U1209 (N_1209,In_520,In_1510);
and U1210 (N_1210,In_7,In_1490);
or U1211 (N_1211,In_1441,In_445);
nand U1212 (N_1212,In_53,In_1553);
or U1213 (N_1213,In_112,In_53);
nor U1214 (N_1214,In_936,In_1337);
and U1215 (N_1215,In_1231,In_44);
or U1216 (N_1216,In_124,In_1291);
or U1217 (N_1217,In_415,In_1534);
nor U1218 (N_1218,In_685,In_1412);
nand U1219 (N_1219,In_1623,In_743);
nand U1220 (N_1220,In_668,In_197);
xor U1221 (N_1221,In_951,In_441);
and U1222 (N_1222,In_1072,In_1944);
nand U1223 (N_1223,In_345,In_101);
xor U1224 (N_1224,In_856,In_670);
xor U1225 (N_1225,In_528,In_55);
nand U1226 (N_1226,In_890,In_142);
or U1227 (N_1227,In_1881,In_584);
nor U1228 (N_1228,In_1687,In_52);
and U1229 (N_1229,In_1166,In_90);
nand U1230 (N_1230,In_74,In_614);
nor U1231 (N_1231,In_1261,In_1065);
nor U1232 (N_1232,In_492,In_823);
nor U1233 (N_1233,In_538,In_1886);
and U1234 (N_1234,In_1683,In_1319);
and U1235 (N_1235,In_132,In_1585);
and U1236 (N_1236,In_10,In_130);
nor U1237 (N_1237,In_106,In_1358);
nand U1238 (N_1238,In_802,In_1569);
or U1239 (N_1239,In_690,In_1138);
nand U1240 (N_1240,In_200,In_1864);
xor U1241 (N_1241,In_1041,In_397);
or U1242 (N_1242,In_1353,In_1971);
nor U1243 (N_1243,In_389,In_1195);
and U1244 (N_1244,In_1445,In_699);
and U1245 (N_1245,In_1670,In_232);
nor U1246 (N_1246,In_1463,In_368);
and U1247 (N_1247,In_1495,In_673);
nor U1248 (N_1248,In_1475,In_1040);
and U1249 (N_1249,In_638,In_755);
or U1250 (N_1250,In_1481,In_193);
nand U1251 (N_1251,In_1467,In_1542);
nand U1252 (N_1252,In_1404,In_1703);
and U1253 (N_1253,In_1848,In_1160);
or U1254 (N_1254,In_465,In_1865);
and U1255 (N_1255,In_690,In_1634);
nor U1256 (N_1256,In_664,In_785);
xor U1257 (N_1257,In_243,In_19);
nor U1258 (N_1258,In_1038,In_1181);
nand U1259 (N_1259,In_708,In_77);
nor U1260 (N_1260,In_427,In_1777);
xor U1261 (N_1261,In_106,In_291);
or U1262 (N_1262,In_1968,In_121);
and U1263 (N_1263,In_47,In_1919);
nor U1264 (N_1264,In_1407,In_899);
or U1265 (N_1265,In_1138,In_11);
and U1266 (N_1266,In_987,In_1392);
or U1267 (N_1267,In_1639,In_162);
nand U1268 (N_1268,In_552,In_1725);
and U1269 (N_1269,In_295,In_1026);
or U1270 (N_1270,In_1890,In_401);
nand U1271 (N_1271,In_1325,In_478);
and U1272 (N_1272,In_1543,In_86);
xor U1273 (N_1273,In_1591,In_1087);
xnor U1274 (N_1274,In_1677,In_287);
nand U1275 (N_1275,In_1163,In_1782);
and U1276 (N_1276,In_1813,In_663);
or U1277 (N_1277,In_684,In_1629);
or U1278 (N_1278,In_71,In_1314);
and U1279 (N_1279,In_1776,In_292);
and U1280 (N_1280,In_1528,In_1461);
nor U1281 (N_1281,In_57,In_1911);
and U1282 (N_1282,In_934,In_1747);
nor U1283 (N_1283,In_1061,In_784);
nor U1284 (N_1284,In_592,In_71);
nor U1285 (N_1285,In_1502,In_356);
or U1286 (N_1286,In_826,In_9);
xnor U1287 (N_1287,In_912,In_1780);
and U1288 (N_1288,In_1497,In_187);
nand U1289 (N_1289,In_217,In_1453);
xnor U1290 (N_1290,In_974,In_28);
and U1291 (N_1291,In_261,In_906);
and U1292 (N_1292,In_237,In_94);
xor U1293 (N_1293,In_297,In_497);
nand U1294 (N_1294,In_982,In_1451);
and U1295 (N_1295,In_10,In_1165);
or U1296 (N_1296,In_416,In_486);
and U1297 (N_1297,In_1901,In_807);
and U1298 (N_1298,In_1039,In_33);
xnor U1299 (N_1299,In_1500,In_1540);
or U1300 (N_1300,In_235,In_1635);
nor U1301 (N_1301,In_1948,In_1875);
xor U1302 (N_1302,In_5,In_1174);
nand U1303 (N_1303,In_1169,In_1179);
and U1304 (N_1304,In_1369,In_1165);
and U1305 (N_1305,In_1460,In_1082);
or U1306 (N_1306,In_1141,In_901);
nand U1307 (N_1307,In_466,In_1872);
and U1308 (N_1308,In_227,In_1389);
or U1309 (N_1309,In_855,In_170);
nor U1310 (N_1310,In_1968,In_1112);
nand U1311 (N_1311,In_1326,In_1343);
nor U1312 (N_1312,In_924,In_213);
and U1313 (N_1313,In_1821,In_1281);
and U1314 (N_1314,In_402,In_333);
nor U1315 (N_1315,In_1657,In_701);
or U1316 (N_1316,In_1622,In_963);
or U1317 (N_1317,In_534,In_1010);
and U1318 (N_1318,In_1767,In_1248);
or U1319 (N_1319,In_1113,In_1566);
nor U1320 (N_1320,In_140,In_729);
and U1321 (N_1321,In_72,In_1817);
nor U1322 (N_1322,In_375,In_1572);
nor U1323 (N_1323,In_418,In_598);
nor U1324 (N_1324,In_1821,In_891);
or U1325 (N_1325,In_1053,In_175);
xor U1326 (N_1326,In_1583,In_1661);
nand U1327 (N_1327,In_652,In_1042);
xor U1328 (N_1328,In_1402,In_773);
or U1329 (N_1329,In_463,In_1742);
and U1330 (N_1330,In_958,In_1103);
and U1331 (N_1331,In_1513,In_993);
xor U1332 (N_1332,In_1683,In_1105);
nand U1333 (N_1333,In_1961,In_1820);
xnor U1334 (N_1334,In_482,In_1378);
nand U1335 (N_1335,In_980,In_752);
and U1336 (N_1336,In_353,In_765);
nand U1337 (N_1337,In_1967,In_1145);
nand U1338 (N_1338,In_743,In_605);
or U1339 (N_1339,In_1047,In_1445);
nor U1340 (N_1340,In_1818,In_82);
or U1341 (N_1341,In_1094,In_1640);
or U1342 (N_1342,In_281,In_299);
and U1343 (N_1343,In_853,In_511);
or U1344 (N_1344,In_1340,In_1119);
xor U1345 (N_1345,In_1,In_552);
xor U1346 (N_1346,In_883,In_977);
or U1347 (N_1347,In_359,In_1032);
nor U1348 (N_1348,In_795,In_1708);
xor U1349 (N_1349,In_518,In_1540);
nand U1350 (N_1350,In_697,In_1677);
nor U1351 (N_1351,In_664,In_8);
or U1352 (N_1352,In_1463,In_1622);
nand U1353 (N_1353,In_1617,In_131);
and U1354 (N_1354,In_1155,In_654);
nor U1355 (N_1355,In_166,In_1821);
nand U1356 (N_1356,In_1266,In_652);
or U1357 (N_1357,In_1179,In_879);
nor U1358 (N_1358,In_148,In_839);
or U1359 (N_1359,In_1438,In_541);
nand U1360 (N_1360,In_631,In_327);
xnor U1361 (N_1361,In_246,In_1649);
nand U1362 (N_1362,In_1435,In_1886);
and U1363 (N_1363,In_410,In_702);
or U1364 (N_1364,In_1485,In_953);
nand U1365 (N_1365,In_1526,In_1865);
nor U1366 (N_1366,In_1143,In_1569);
nand U1367 (N_1367,In_1349,In_663);
nor U1368 (N_1368,In_130,In_209);
or U1369 (N_1369,In_1759,In_1526);
nor U1370 (N_1370,In_1506,In_1518);
and U1371 (N_1371,In_1972,In_1859);
or U1372 (N_1372,In_1048,In_1929);
nor U1373 (N_1373,In_52,In_932);
and U1374 (N_1374,In_687,In_807);
or U1375 (N_1375,In_1267,In_1602);
nor U1376 (N_1376,In_217,In_1119);
nor U1377 (N_1377,In_1992,In_1304);
nor U1378 (N_1378,In_338,In_1694);
and U1379 (N_1379,In_430,In_1725);
nand U1380 (N_1380,In_1654,In_1120);
nand U1381 (N_1381,In_1567,In_1898);
or U1382 (N_1382,In_748,In_1583);
and U1383 (N_1383,In_8,In_542);
or U1384 (N_1384,In_825,In_1922);
or U1385 (N_1385,In_946,In_1998);
and U1386 (N_1386,In_550,In_1157);
and U1387 (N_1387,In_770,In_1285);
nor U1388 (N_1388,In_293,In_237);
or U1389 (N_1389,In_1052,In_261);
nand U1390 (N_1390,In_1862,In_1816);
xor U1391 (N_1391,In_1975,In_1939);
and U1392 (N_1392,In_1725,In_385);
and U1393 (N_1393,In_1854,In_724);
nand U1394 (N_1394,In_1744,In_1693);
or U1395 (N_1395,In_1518,In_1676);
nor U1396 (N_1396,In_1401,In_42);
nand U1397 (N_1397,In_1368,In_534);
xnor U1398 (N_1398,In_150,In_1542);
and U1399 (N_1399,In_74,In_851);
nor U1400 (N_1400,In_230,In_943);
xor U1401 (N_1401,In_1343,In_200);
or U1402 (N_1402,In_508,In_1063);
or U1403 (N_1403,In_1604,In_216);
xnor U1404 (N_1404,In_1019,In_843);
or U1405 (N_1405,In_1432,In_70);
or U1406 (N_1406,In_171,In_920);
nor U1407 (N_1407,In_994,In_1075);
nand U1408 (N_1408,In_1587,In_259);
and U1409 (N_1409,In_1857,In_818);
xor U1410 (N_1410,In_170,In_1238);
nand U1411 (N_1411,In_1646,In_1831);
nor U1412 (N_1412,In_1095,In_1960);
nand U1413 (N_1413,In_913,In_58);
nand U1414 (N_1414,In_1274,In_1525);
and U1415 (N_1415,In_1639,In_819);
and U1416 (N_1416,In_1634,In_1624);
nor U1417 (N_1417,In_1268,In_620);
or U1418 (N_1418,In_1612,In_774);
nor U1419 (N_1419,In_1128,In_1449);
or U1420 (N_1420,In_147,In_1152);
or U1421 (N_1421,In_891,In_1763);
nor U1422 (N_1422,In_712,In_92);
or U1423 (N_1423,In_103,In_1398);
nand U1424 (N_1424,In_340,In_164);
nand U1425 (N_1425,In_35,In_802);
nand U1426 (N_1426,In_1303,In_1865);
xor U1427 (N_1427,In_1972,In_727);
nand U1428 (N_1428,In_446,In_1788);
nor U1429 (N_1429,In_769,In_699);
nor U1430 (N_1430,In_313,In_1790);
and U1431 (N_1431,In_1019,In_148);
nand U1432 (N_1432,In_1567,In_1660);
nand U1433 (N_1433,In_1061,In_572);
or U1434 (N_1434,In_726,In_770);
and U1435 (N_1435,In_1841,In_829);
nor U1436 (N_1436,In_1486,In_1831);
and U1437 (N_1437,In_308,In_1337);
or U1438 (N_1438,In_1572,In_287);
nand U1439 (N_1439,In_1176,In_1682);
nand U1440 (N_1440,In_1828,In_1454);
or U1441 (N_1441,In_580,In_975);
and U1442 (N_1442,In_1270,In_1242);
and U1443 (N_1443,In_888,In_1637);
nand U1444 (N_1444,In_963,In_569);
or U1445 (N_1445,In_671,In_1344);
nor U1446 (N_1446,In_116,In_157);
nand U1447 (N_1447,In_40,In_1634);
and U1448 (N_1448,In_1055,In_793);
and U1449 (N_1449,In_606,In_33);
nand U1450 (N_1450,In_146,In_1302);
and U1451 (N_1451,In_1093,In_1897);
nand U1452 (N_1452,In_452,In_1746);
or U1453 (N_1453,In_1035,In_174);
xnor U1454 (N_1454,In_615,In_1621);
nor U1455 (N_1455,In_1622,In_170);
nand U1456 (N_1456,In_1149,In_1505);
xnor U1457 (N_1457,In_1598,In_1832);
xnor U1458 (N_1458,In_630,In_1456);
nor U1459 (N_1459,In_1400,In_242);
or U1460 (N_1460,In_171,In_1609);
or U1461 (N_1461,In_1547,In_1569);
or U1462 (N_1462,In_1798,In_1757);
and U1463 (N_1463,In_1396,In_1938);
or U1464 (N_1464,In_1995,In_1392);
nor U1465 (N_1465,In_1480,In_75);
nor U1466 (N_1466,In_963,In_203);
or U1467 (N_1467,In_1964,In_1748);
nand U1468 (N_1468,In_1774,In_1167);
nand U1469 (N_1469,In_264,In_1979);
nand U1470 (N_1470,In_787,In_1174);
and U1471 (N_1471,In_116,In_1641);
nor U1472 (N_1472,In_1318,In_652);
nand U1473 (N_1473,In_65,In_455);
xor U1474 (N_1474,In_85,In_914);
nor U1475 (N_1475,In_102,In_1146);
or U1476 (N_1476,In_400,In_1303);
nor U1477 (N_1477,In_1562,In_508);
and U1478 (N_1478,In_56,In_1866);
nor U1479 (N_1479,In_859,In_1712);
nand U1480 (N_1480,In_1294,In_933);
nand U1481 (N_1481,In_1826,In_886);
nor U1482 (N_1482,In_975,In_1766);
or U1483 (N_1483,In_1131,In_1628);
nor U1484 (N_1484,In_1095,In_843);
nor U1485 (N_1485,In_362,In_1897);
nand U1486 (N_1486,In_1806,In_1254);
and U1487 (N_1487,In_284,In_917);
and U1488 (N_1488,In_1820,In_53);
and U1489 (N_1489,In_1665,In_1704);
nand U1490 (N_1490,In_1870,In_1471);
and U1491 (N_1491,In_1257,In_225);
and U1492 (N_1492,In_1108,In_1394);
nand U1493 (N_1493,In_514,In_446);
nand U1494 (N_1494,In_1668,In_256);
and U1495 (N_1495,In_1176,In_745);
or U1496 (N_1496,In_928,In_910);
or U1497 (N_1497,In_1841,In_1280);
and U1498 (N_1498,In_1643,In_146);
nand U1499 (N_1499,In_222,In_1985);
nand U1500 (N_1500,In_1616,In_1077);
nand U1501 (N_1501,In_293,In_1529);
and U1502 (N_1502,In_1691,In_1278);
nor U1503 (N_1503,In_1699,In_1991);
or U1504 (N_1504,In_1895,In_432);
nor U1505 (N_1505,In_1917,In_570);
and U1506 (N_1506,In_205,In_1837);
nand U1507 (N_1507,In_965,In_743);
nand U1508 (N_1508,In_509,In_1518);
nor U1509 (N_1509,In_116,In_962);
and U1510 (N_1510,In_1567,In_1090);
xor U1511 (N_1511,In_1128,In_1751);
nor U1512 (N_1512,In_302,In_1181);
xnor U1513 (N_1513,In_863,In_1379);
or U1514 (N_1514,In_1458,In_1729);
or U1515 (N_1515,In_211,In_958);
or U1516 (N_1516,In_416,In_260);
nor U1517 (N_1517,In_910,In_1228);
nor U1518 (N_1518,In_151,In_1740);
or U1519 (N_1519,In_1,In_825);
nand U1520 (N_1520,In_1553,In_1672);
xor U1521 (N_1521,In_635,In_55);
xor U1522 (N_1522,In_1319,In_1444);
nand U1523 (N_1523,In_1810,In_1710);
xnor U1524 (N_1524,In_1153,In_1210);
or U1525 (N_1525,In_999,In_235);
nand U1526 (N_1526,In_482,In_1759);
nor U1527 (N_1527,In_818,In_1634);
nand U1528 (N_1528,In_400,In_1388);
nand U1529 (N_1529,In_1806,In_1352);
or U1530 (N_1530,In_1697,In_1700);
nand U1531 (N_1531,In_731,In_1803);
nor U1532 (N_1532,In_1401,In_1311);
nor U1533 (N_1533,In_1612,In_1972);
nor U1534 (N_1534,In_1875,In_402);
nand U1535 (N_1535,In_1737,In_1438);
nor U1536 (N_1536,In_968,In_1083);
xor U1537 (N_1537,In_1409,In_1859);
and U1538 (N_1538,In_252,In_266);
nor U1539 (N_1539,In_49,In_1061);
nor U1540 (N_1540,In_272,In_703);
nand U1541 (N_1541,In_195,In_230);
nand U1542 (N_1542,In_927,In_372);
nand U1543 (N_1543,In_42,In_1424);
nor U1544 (N_1544,In_990,In_1723);
and U1545 (N_1545,In_1163,In_658);
nor U1546 (N_1546,In_1312,In_570);
and U1547 (N_1547,In_1185,In_229);
nand U1548 (N_1548,In_525,In_225);
and U1549 (N_1549,In_1437,In_273);
nand U1550 (N_1550,In_1785,In_233);
nor U1551 (N_1551,In_657,In_775);
nor U1552 (N_1552,In_991,In_1861);
or U1553 (N_1553,In_662,In_755);
nand U1554 (N_1554,In_897,In_700);
or U1555 (N_1555,In_103,In_35);
and U1556 (N_1556,In_134,In_651);
nand U1557 (N_1557,In_1805,In_1782);
xnor U1558 (N_1558,In_1888,In_25);
nor U1559 (N_1559,In_1213,In_537);
or U1560 (N_1560,In_977,In_1961);
or U1561 (N_1561,In_1548,In_322);
nand U1562 (N_1562,In_1733,In_50);
nor U1563 (N_1563,In_456,In_1600);
and U1564 (N_1564,In_283,In_637);
nor U1565 (N_1565,In_607,In_1223);
nand U1566 (N_1566,In_1420,In_1594);
or U1567 (N_1567,In_1297,In_1863);
and U1568 (N_1568,In_1886,In_213);
nor U1569 (N_1569,In_710,In_371);
or U1570 (N_1570,In_110,In_781);
nand U1571 (N_1571,In_1395,In_535);
nand U1572 (N_1572,In_1668,In_144);
nand U1573 (N_1573,In_163,In_479);
xor U1574 (N_1574,In_759,In_1306);
and U1575 (N_1575,In_465,In_1175);
or U1576 (N_1576,In_712,In_442);
xor U1577 (N_1577,In_1767,In_1683);
or U1578 (N_1578,In_64,In_798);
or U1579 (N_1579,In_1136,In_1236);
nor U1580 (N_1580,In_1671,In_858);
and U1581 (N_1581,In_667,In_684);
or U1582 (N_1582,In_1489,In_1334);
and U1583 (N_1583,In_42,In_516);
xnor U1584 (N_1584,In_1096,In_1879);
and U1585 (N_1585,In_48,In_65);
or U1586 (N_1586,In_1819,In_1764);
nor U1587 (N_1587,In_1738,In_187);
nand U1588 (N_1588,In_1103,In_1207);
nand U1589 (N_1589,In_758,In_1413);
nor U1590 (N_1590,In_1465,In_1528);
or U1591 (N_1591,In_1399,In_1302);
and U1592 (N_1592,In_1058,In_24);
xor U1593 (N_1593,In_1277,In_11);
and U1594 (N_1594,In_261,In_983);
nor U1595 (N_1595,In_373,In_121);
nand U1596 (N_1596,In_756,In_1649);
nor U1597 (N_1597,In_643,In_707);
nor U1598 (N_1598,In_1194,In_658);
nor U1599 (N_1599,In_478,In_397);
nand U1600 (N_1600,In_1529,In_539);
and U1601 (N_1601,In_481,In_184);
or U1602 (N_1602,In_452,In_1016);
nor U1603 (N_1603,In_140,In_1838);
nand U1604 (N_1604,In_1959,In_1114);
nor U1605 (N_1605,In_978,In_1531);
or U1606 (N_1606,In_1344,In_581);
and U1607 (N_1607,In_1629,In_1014);
and U1608 (N_1608,In_940,In_428);
xor U1609 (N_1609,In_772,In_361);
nor U1610 (N_1610,In_1715,In_1126);
xor U1611 (N_1611,In_176,In_235);
nor U1612 (N_1612,In_737,In_584);
or U1613 (N_1613,In_1480,In_1304);
xor U1614 (N_1614,In_131,In_33);
or U1615 (N_1615,In_1512,In_909);
nor U1616 (N_1616,In_1746,In_1538);
or U1617 (N_1617,In_1988,In_1341);
nand U1618 (N_1618,In_1923,In_642);
nor U1619 (N_1619,In_1470,In_1433);
nor U1620 (N_1620,In_1262,In_1294);
nand U1621 (N_1621,In_1256,In_776);
and U1622 (N_1622,In_1690,In_1142);
nor U1623 (N_1623,In_490,In_344);
nand U1624 (N_1624,In_293,In_1568);
and U1625 (N_1625,In_1788,In_1322);
nand U1626 (N_1626,In_766,In_217);
nand U1627 (N_1627,In_1227,In_960);
and U1628 (N_1628,In_188,In_939);
and U1629 (N_1629,In_1154,In_381);
nand U1630 (N_1630,In_1150,In_1034);
or U1631 (N_1631,In_4,In_1008);
and U1632 (N_1632,In_1814,In_233);
and U1633 (N_1633,In_1237,In_952);
xor U1634 (N_1634,In_1512,In_49);
nand U1635 (N_1635,In_46,In_1310);
nor U1636 (N_1636,In_1624,In_178);
or U1637 (N_1637,In_1327,In_1913);
or U1638 (N_1638,In_293,In_306);
and U1639 (N_1639,In_1538,In_1411);
and U1640 (N_1640,In_1816,In_339);
nor U1641 (N_1641,In_1520,In_1993);
xnor U1642 (N_1642,In_1001,In_773);
nand U1643 (N_1643,In_1680,In_452);
or U1644 (N_1644,In_1083,In_1998);
nand U1645 (N_1645,In_1780,In_300);
and U1646 (N_1646,In_1084,In_1089);
or U1647 (N_1647,In_1300,In_1399);
and U1648 (N_1648,In_908,In_505);
nor U1649 (N_1649,In_1551,In_293);
xor U1650 (N_1650,In_377,In_705);
xnor U1651 (N_1651,In_110,In_1421);
xnor U1652 (N_1652,In_279,In_1924);
and U1653 (N_1653,In_1578,In_1265);
and U1654 (N_1654,In_1881,In_106);
and U1655 (N_1655,In_973,In_1864);
and U1656 (N_1656,In_362,In_258);
nor U1657 (N_1657,In_1103,In_1892);
nand U1658 (N_1658,In_1551,In_949);
nor U1659 (N_1659,In_519,In_509);
and U1660 (N_1660,In_1026,In_443);
nor U1661 (N_1661,In_1731,In_442);
and U1662 (N_1662,In_1814,In_852);
nand U1663 (N_1663,In_1659,In_640);
nor U1664 (N_1664,In_517,In_1223);
or U1665 (N_1665,In_1587,In_1569);
or U1666 (N_1666,In_1601,In_1850);
nand U1667 (N_1667,In_715,In_1953);
nand U1668 (N_1668,In_1450,In_893);
nor U1669 (N_1669,In_300,In_919);
nand U1670 (N_1670,In_19,In_418);
nand U1671 (N_1671,In_432,In_1758);
nor U1672 (N_1672,In_692,In_1612);
and U1673 (N_1673,In_1943,In_103);
xnor U1674 (N_1674,In_1386,In_1204);
nand U1675 (N_1675,In_940,In_80);
nor U1676 (N_1676,In_1151,In_598);
nand U1677 (N_1677,In_324,In_218);
nand U1678 (N_1678,In_1502,In_617);
nand U1679 (N_1679,In_858,In_624);
or U1680 (N_1680,In_23,In_546);
nand U1681 (N_1681,In_193,In_1944);
or U1682 (N_1682,In_1199,In_1448);
nor U1683 (N_1683,In_250,In_700);
nor U1684 (N_1684,In_1088,In_441);
nor U1685 (N_1685,In_779,In_1812);
nand U1686 (N_1686,In_821,In_1203);
and U1687 (N_1687,In_1988,In_785);
nor U1688 (N_1688,In_986,In_1179);
or U1689 (N_1689,In_1962,In_586);
xnor U1690 (N_1690,In_1735,In_69);
or U1691 (N_1691,In_1388,In_862);
nor U1692 (N_1692,In_1915,In_1548);
nor U1693 (N_1693,In_502,In_1183);
and U1694 (N_1694,In_1387,In_1083);
or U1695 (N_1695,In_1783,In_1083);
nand U1696 (N_1696,In_1968,In_385);
xor U1697 (N_1697,In_1250,In_15);
and U1698 (N_1698,In_382,In_1824);
nor U1699 (N_1699,In_1216,In_896);
xnor U1700 (N_1700,In_524,In_464);
or U1701 (N_1701,In_1224,In_469);
and U1702 (N_1702,In_1721,In_1936);
nor U1703 (N_1703,In_1182,In_1183);
or U1704 (N_1704,In_266,In_426);
xor U1705 (N_1705,In_362,In_174);
and U1706 (N_1706,In_13,In_1468);
nor U1707 (N_1707,In_1980,In_440);
nand U1708 (N_1708,In_1786,In_953);
nor U1709 (N_1709,In_1038,In_1415);
xor U1710 (N_1710,In_1609,In_649);
nor U1711 (N_1711,In_176,In_1621);
nand U1712 (N_1712,In_1353,In_589);
or U1713 (N_1713,In_517,In_25);
nor U1714 (N_1714,In_955,In_1448);
or U1715 (N_1715,In_465,In_1204);
or U1716 (N_1716,In_1920,In_1560);
xnor U1717 (N_1717,In_1618,In_599);
and U1718 (N_1718,In_1346,In_252);
nor U1719 (N_1719,In_616,In_1914);
and U1720 (N_1720,In_1231,In_937);
or U1721 (N_1721,In_535,In_855);
nand U1722 (N_1722,In_314,In_1955);
or U1723 (N_1723,In_960,In_1759);
nor U1724 (N_1724,In_1247,In_60);
nand U1725 (N_1725,In_1297,In_558);
or U1726 (N_1726,In_564,In_1141);
xor U1727 (N_1727,In_1345,In_1878);
or U1728 (N_1728,In_1730,In_1074);
xnor U1729 (N_1729,In_1277,In_1917);
nor U1730 (N_1730,In_1799,In_727);
nand U1731 (N_1731,In_286,In_1293);
and U1732 (N_1732,In_259,In_1347);
and U1733 (N_1733,In_366,In_1394);
xor U1734 (N_1734,In_1780,In_1959);
or U1735 (N_1735,In_544,In_135);
and U1736 (N_1736,In_817,In_1618);
nand U1737 (N_1737,In_237,In_1141);
nand U1738 (N_1738,In_1518,In_1603);
nor U1739 (N_1739,In_407,In_1042);
and U1740 (N_1740,In_916,In_1913);
and U1741 (N_1741,In_981,In_116);
nor U1742 (N_1742,In_614,In_242);
nor U1743 (N_1743,In_1468,In_650);
nor U1744 (N_1744,In_1099,In_1001);
nand U1745 (N_1745,In_288,In_63);
xor U1746 (N_1746,In_836,In_658);
or U1747 (N_1747,In_1617,In_1576);
or U1748 (N_1748,In_1971,In_1400);
nor U1749 (N_1749,In_343,In_400);
nand U1750 (N_1750,In_490,In_133);
nor U1751 (N_1751,In_1846,In_236);
and U1752 (N_1752,In_732,In_360);
nand U1753 (N_1753,In_1098,In_532);
nand U1754 (N_1754,In_1421,In_1952);
and U1755 (N_1755,In_370,In_1878);
and U1756 (N_1756,In_482,In_468);
or U1757 (N_1757,In_1814,In_1204);
nand U1758 (N_1758,In_118,In_1983);
nand U1759 (N_1759,In_1786,In_1634);
xnor U1760 (N_1760,In_283,In_201);
or U1761 (N_1761,In_1207,In_1209);
or U1762 (N_1762,In_435,In_937);
nand U1763 (N_1763,In_1552,In_1139);
nand U1764 (N_1764,In_1412,In_515);
and U1765 (N_1765,In_1101,In_797);
nand U1766 (N_1766,In_1178,In_508);
or U1767 (N_1767,In_68,In_463);
nor U1768 (N_1768,In_1867,In_1934);
and U1769 (N_1769,In_110,In_788);
nand U1770 (N_1770,In_1709,In_885);
or U1771 (N_1771,In_623,In_829);
and U1772 (N_1772,In_473,In_1629);
and U1773 (N_1773,In_518,In_879);
nand U1774 (N_1774,In_768,In_64);
nor U1775 (N_1775,In_1784,In_1280);
nand U1776 (N_1776,In_701,In_609);
nor U1777 (N_1777,In_1240,In_237);
nor U1778 (N_1778,In_218,In_1099);
nor U1779 (N_1779,In_1233,In_428);
nor U1780 (N_1780,In_788,In_1442);
nand U1781 (N_1781,In_898,In_883);
nand U1782 (N_1782,In_461,In_1115);
and U1783 (N_1783,In_1789,In_985);
or U1784 (N_1784,In_1290,In_981);
xor U1785 (N_1785,In_1250,In_1345);
and U1786 (N_1786,In_56,In_1609);
nand U1787 (N_1787,In_1297,In_1471);
nor U1788 (N_1788,In_989,In_1567);
and U1789 (N_1789,In_488,In_1779);
or U1790 (N_1790,In_891,In_529);
nand U1791 (N_1791,In_929,In_846);
and U1792 (N_1792,In_1208,In_803);
nand U1793 (N_1793,In_672,In_35);
or U1794 (N_1794,In_648,In_926);
nor U1795 (N_1795,In_1762,In_1171);
nand U1796 (N_1796,In_268,In_1342);
or U1797 (N_1797,In_1071,In_1318);
and U1798 (N_1798,In_923,In_1007);
nand U1799 (N_1799,In_1071,In_835);
and U1800 (N_1800,In_20,In_1412);
nand U1801 (N_1801,In_849,In_1881);
nor U1802 (N_1802,In_1728,In_880);
nand U1803 (N_1803,In_1391,In_636);
or U1804 (N_1804,In_962,In_584);
xor U1805 (N_1805,In_1989,In_1697);
nor U1806 (N_1806,In_493,In_240);
nor U1807 (N_1807,In_942,In_1524);
xnor U1808 (N_1808,In_1809,In_1593);
or U1809 (N_1809,In_1914,In_778);
nor U1810 (N_1810,In_978,In_124);
or U1811 (N_1811,In_949,In_1366);
or U1812 (N_1812,In_1395,In_1315);
and U1813 (N_1813,In_146,In_121);
and U1814 (N_1814,In_1344,In_848);
or U1815 (N_1815,In_1961,In_639);
and U1816 (N_1816,In_505,In_1780);
nor U1817 (N_1817,In_1338,In_1880);
xor U1818 (N_1818,In_1834,In_916);
nand U1819 (N_1819,In_1839,In_1452);
or U1820 (N_1820,In_1443,In_424);
or U1821 (N_1821,In_1759,In_335);
and U1822 (N_1822,In_902,In_242);
and U1823 (N_1823,In_745,In_800);
xnor U1824 (N_1824,In_369,In_1518);
nor U1825 (N_1825,In_215,In_526);
or U1826 (N_1826,In_1329,In_1130);
nor U1827 (N_1827,In_176,In_693);
nor U1828 (N_1828,In_560,In_1085);
or U1829 (N_1829,In_51,In_1689);
nand U1830 (N_1830,In_1277,In_1116);
and U1831 (N_1831,In_1870,In_28);
nor U1832 (N_1832,In_310,In_1372);
or U1833 (N_1833,In_523,In_1149);
or U1834 (N_1834,In_1153,In_525);
or U1835 (N_1835,In_806,In_963);
xnor U1836 (N_1836,In_690,In_1937);
nor U1837 (N_1837,In_310,In_1269);
or U1838 (N_1838,In_372,In_1313);
and U1839 (N_1839,In_358,In_943);
nand U1840 (N_1840,In_1100,In_860);
nor U1841 (N_1841,In_1999,In_803);
nor U1842 (N_1842,In_1968,In_515);
and U1843 (N_1843,In_1781,In_502);
nor U1844 (N_1844,In_606,In_331);
and U1845 (N_1845,In_1505,In_553);
nand U1846 (N_1846,In_926,In_251);
nor U1847 (N_1847,In_892,In_1256);
and U1848 (N_1848,In_1480,In_761);
nor U1849 (N_1849,In_1396,In_841);
nand U1850 (N_1850,In_1731,In_1593);
nor U1851 (N_1851,In_891,In_897);
xor U1852 (N_1852,In_219,In_239);
nor U1853 (N_1853,In_150,In_943);
and U1854 (N_1854,In_910,In_602);
nor U1855 (N_1855,In_850,In_1483);
nand U1856 (N_1856,In_1817,In_919);
nand U1857 (N_1857,In_762,In_1918);
nand U1858 (N_1858,In_119,In_713);
and U1859 (N_1859,In_24,In_1900);
or U1860 (N_1860,In_1234,In_962);
xor U1861 (N_1861,In_629,In_1853);
xnor U1862 (N_1862,In_1129,In_578);
and U1863 (N_1863,In_1106,In_1663);
and U1864 (N_1864,In_1716,In_1297);
or U1865 (N_1865,In_40,In_1990);
xor U1866 (N_1866,In_707,In_1611);
xnor U1867 (N_1867,In_1661,In_790);
nor U1868 (N_1868,In_1479,In_800);
or U1869 (N_1869,In_255,In_84);
nand U1870 (N_1870,In_1451,In_154);
or U1871 (N_1871,In_1555,In_617);
and U1872 (N_1872,In_1441,In_42);
nand U1873 (N_1873,In_101,In_1416);
or U1874 (N_1874,In_1061,In_547);
xor U1875 (N_1875,In_818,In_1722);
nor U1876 (N_1876,In_256,In_1224);
nand U1877 (N_1877,In_45,In_114);
nand U1878 (N_1878,In_894,In_1599);
or U1879 (N_1879,In_1693,In_1173);
nand U1880 (N_1880,In_1871,In_213);
and U1881 (N_1881,In_384,In_870);
or U1882 (N_1882,In_1202,In_1007);
xnor U1883 (N_1883,In_1560,In_1620);
nor U1884 (N_1884,In_1194,In_709);
and U1885 (N_1885,In_936,In_1410);
and U1886 (N_1886,In_738,In_1776);
nand U1887 (N_1887,In_1621,In_265);
nand U1888 (N_1888,In_1245,In_851);
and U1889 (N_1889,In_1126,In_1665);
xor U1890 (N_1890,In_1842,In_167);
or U1891 (N_1891,In_1790,In_1363);
nand U1892 (N_1892,In_392,In_978);
and U1893 (N_1893,In_533,In_1808);
nor U1894 (N_1894,In_1733,In_439);
nor U1895 (N_1895,In_958,In_1585);
and U1896 (N_1896,In_1152,In_517);
nand U1897 (N_1897,In_652,In_637);
nor U1898 (N_1898,In_1232,In_613);
xnor U1899 (N_1899,In_1042,In_400);
or U1900 (N_1900,In_1038,In_465);
xor U1901 (N_1901,In_1612,In_1181);
nand U1902 (N_1902,In_1461,In_1454);
or U1903 (N_1903,In_700,In_1874);
nand U1904 (N_1904,In_236,In_1755);
nor U1905 (N_1905,In_1547,In_1864);
nor U1906 (N_1906,In_1304,In_1178);
nor U1907 (N_1907,In_827,In_1281);
nor U1908 (N_1908,In_221,In_1871);
nand U1909 (N_1909,In_394,In_779);
or U1910 (N_1910,In_191,In_780);
xnor U1911 (N_1911,In_1920,In_1625);
and U1912 (N_1912,In_1743,In_1858);
or U1913 (N_1913,In_1575,In_717);
nor U1914 (N_1914,In_436,In_538);
nand U1915 (N_1915,In_918,In_213);
nor U1916 (N_1916,In_1461,In_85);
nand U1917 (N_1917,In_850,In_497);
nand U1918 (N_1918,In_1532,In_927);
and U1919 (N_1919,In_1230,In_1612);
or U1920 (N_1920,In_1334,In_1087);
nor U1921 (N_1921,In_718,In_1919);
nor U1922 (N_1922,In_340,In_803);
or U1923 (N_1923,In_37,In_159);
nor U1924 (N_1924,In_821,In_1261);
nand U1925 (N_1925,In_150,In_1134);
nor U1926 (N_1926,In_262,In_818);
nor U1927 (N_1927,In_351,In_1580);
or U1928 (N_1928,In_553,In_1984);
nand U1929 (N_1929,In_1720,In_1536);
and U1930 (N_1930,In_1412,In_42);
and U1931 (N_1931,In_1685,In_1352);
and U1932 (N_1932,In_679,In_123);
nand U1933 (N_1933,In_724,In_387);
nor U1934 (N_1934,In_557,In_597);
nor U1935 (N_1935,In_655,In_872);
and U1936 (N_1936,In_1886,In_1984);
nor U1937 (N_1937,In_1587,In_1886);
or U1938 (N_1938,In_1949,In_230);
nand U1939 (N_1939,In_116,In_820);
nor U1940 (N_1940,In_1986,In_1222);
and U1941 (N_1941,In_330,In_285);
nand U1942 (N_1942,In_1098,In_1909);
nor U1943 (N_1943,In_1475,In_1011);
nor U1944 (N_1944,In_1753,In_1750);
nand U1945 (N_1945,In_774,In_451);
and U1946 (N_1946,In_1265,In_1293);
or U1947 (N_1947,In_1586,In_1579);
xnor U1948 (N_1948,In_1929,In_1506);
or U1949 (N_1949,In_1773,In_1546);
nand U1950 (N_1950,In_161,In_1796);
nand U1951 (N_1951,In_169,In_603);
nand U1952 (N_1952,In_1367,In_1864);
nand U1953 (N_1953,In_1992,In_777);
or U1954 (N_1954,In_1851,In_1167);
and U1955 (N_1955,In_472,In_1553);
nand U1956 (N_1956,In_27,In_1529);
nand U1957 (N_1957,In_342,In_1343);
nand U1958 (N_1958,In_353,In_1711);
nor U1959 (N_1959,In_580,In_438);
nand U1960 (N_1960,In_512,In_100);
or U1961 (N_1961,In_1843,In_837);
or U1962 (N_1962,In_797,In_1504);
or U1963 (N_1963,In_1931,In_1105);
nand U1964 (N_1964,In_23,In_1104);
nand U1965 (N_1965,In_485,In_1566);
and U1966 (N_1966,In_1054,In_1604);
or U1967 (N_1967,In_902,In_325);
nor U1968 (N_1968,In_1325,In_1319);
nor U1969 (N_1969,In_172,In_418);
nand U1970 (N_1970,In_1139,In_1641);
xor U1971 (N_1971,In_792,In_1745);
or U1972 (N_1972,In_872,In_1132);
nand U1973 (N_1973,In_766,In_512);
or U1974 (N_1974,In_1992,In_646);
or U1975 (N_1975,In_1173,In_1074);
nand U1976 (N_1976,In_1987,In_1701);
nor U1977 (N_1977,In_31,In_1231);
and U1978 (N_1978,In_940,In_1606);
nor U1979 (N_1979,In_1297,In_1144);
or U1980 (N_1980,In_221,In_378);
and U1981 (N_1981,In_712,In_1535);
xor U1982 (N_1982,In_715,In_103);
nor U1983 (N_1983,In_1737,In_782);
and U1984 (N_1984,In_983,In_517);
and U1985 (N_1985,In_764,In_1612);
nand U1986 (N_1986,In_414,In_1193);
nand U1987 (N_1987,In_1578,In_1646);
xnor U1988 (N_1988,In_1294,In_394);
or U1989 (N_1989,In_746,In_1459);
and U1990 (N_1990,In_469,In_1113);
or U1991 (N_1991,In_1832,In_674);
or U1992 (N_1992,In_1341,In_638);
xnor U1993 (N_1993,In_1458,In_1531);
xor U1994 (N_1994,In_700,In_1445);
nor U1995 (N_1995,In_335,In_1545);
nor U1996 (N_1996,In_1202,In_1232);
nor U1997 (N_1997,In_1719,In_196);
or U1998 (N_1998,In_284,In_153);
or U1999 (N_1999,In_1464,In_1232);
xor U2000 (N_2000,In_1226,In_955);
nand U2001 (N_2001,In_767,In_456);
xor U2002 (N_2002,In_1883,In_93);
and U2003 (N_2003,In_246,In_1922);
or U2004 (N_2004,In_1315,In_752);
nand U2005 (N_2005,In_210,In_1161);
or U2006 (N_2006,In_343,In_780);
nor U2007 (N_2007,In_1839,In_1941);
nand U2008 (N_2008,In_1646,In_1002);
nor U2009 (N_2009,In_1019,In_276);
or U2010 (N_2010,In_1732,In_1613);
nor U2011 (N_2011,In_1971,In_577);
or U2012 (N_2012,In_1079,In_1180);
nor U2013 (N_2013,In_353,In_603);
nor U2014 (N_2014,In_1343,In_473);
nand U2015 (N_2015,In_1348,In_764);
nand U2016 (N_2016,In_1002,In_1407);
or U2017 (N_2017,In_823,In_1737);
nand U2018 (N_2018,In_129,In_542);
and U2019 (N_2019,In_323,In_1251);
or U2020 (N_2020,In_281,In_1931);
xnor U2021 (N_2021,In_688,In_1668);
nand U2022 (N_2022,In_1407,In_247);
xnor U2023 (N_2023,In_1300,In_1666);
and U2024 (N_2024,In_1508,In_691);
xor U2025 (N_2025,In_882,In_1650);
nand U2026 (N_2026,In_538,In_588);
xnor U2027 (N_2027,In_1207,In_1465);
or U2028 (N_2028,In_1007,In_142);
or U2029 (N_2029,In_302,In_1030);
nor U2030 (N_2030,In_707,In_836);
nor U2031 (N_2031,In_1682,In_799);
xor U2032 (N_2032,In_300,In_1708);
nor U2033 (N_2033,In_297,In_676);
or U2034 (N_2034,In_1116,In_1557);
nand U2035 (N_2035,In_1199,In_597);
or U2036 (N_2036,In_464,In_1072);
nand U2037 (N_2037,In_2,In_232);
nand U2038 (N_2038,In_253,In_231);
nor U2039 (N_2039,In_672,In_1379);
or U2040 (N_2040,In_1795,In_1816);
and U2041 (N_2041,In_1797,In_1324);
nor U2042 (N_2042,In_770,In_1332);
and U2043 (N_2043,In_1836,In_1879);
nand U2044 (N_2044,In_1456,In_781);
and U2045 (N_2045,In_1517,In_630);
or U2046 (N_2046,In_900,In_382);
xnor U2047 (N_2047,In_1439,In_229);
or U2048 (N_2048,In_621,In_77);
or U2049 (N_2049,In_253,In_1233);
or U2050 (N_2050,In_947,In_490);
or U2051 (N_2051,In_1162,In_516);
and U2052 (N_2052,In_953,In_1080);
and U2053 (N_2053,In_1787,In_1093);
nor U2054 (N_2054,In_1749,In_1139);
and U2055 (N_2055,In_1102,In_1135);
nor U2056 (N_2056,In_845,In_608);
nand U2057 (N_2057,In_947,In_323);
nand U2058 (N_2058,In_535,In_787);
and U2059 (N_2059,In_54,In_948);
nand U2060 (N_2060,In_1790,In_467);
or U2061 (N_2061,In_505,In_1065);
nor U2062 (N_2062,In_287,In_1338);
nand U2063 (N_2063,In_940,In_1535);
and U2064 (N_2064,In_1581,In_1269);
or U2065 (N_2065,In_1396,In_1607);
or U2066 (N_2066,In_715,In_1623);
or U2067 (N_2067,In_345,In_1512);
or U2068 (N_2068,In_1082,In_1176);
and U2069 (N_2069,In_90,In_135);
nor U2070 (N_2070,In_839,In_806);
nor U2071 (N_2071,In_1674,In_345);
nor U2072 (N_2072,In_1676,In_1892);
or U2073 (N_2073,In_86,In_1465);
nor U2074 (N_2074,In_1129,In_1712);
or U2075 (N_2075,In_994,In_1422);
xnor U2076 (N_2076,In_1599,In_795);
nand U2077 (N_2077,In_162,In_1289);
xor U2078 (N_2078,In_1342,In_713);
or U2079 (N_2079,In_1603,In_51);
or U2080 (N_2080,In_48,In_1313);
and U2081 (N_2081,In_237,In_97);
nor U2082 (N_2082,In_1773,In_1363);
nand U2083 (N_2083,In_1642,In_224);
xor U2084 (N_2084,In_293,In_1982);
xor U2085 (N_2085,In_1024,In_562);
and U2086 (N_2086,In_1768,In_630);
or U2087 (N_2087,In_945,In_1678);
and U2088 (N_2088,In_105,In_875);
nand U2089 (N_2089,In_1017,In_1755);
or U2090 (N_2090,In_360,In_709);
and U2091 (N_2091,In_971,In_1512);
or U2092 (N_2092,In_689,In_746);
or U2093 (N_2093,In_337,In_1881);
xnor U2094 (N_2094,In_1171,In_820);
and U2095 (N_2095,In_1860,In_1946);
nor U2096 (N_2096,In_388,In_401);
or U2097 (N_2097,In_609,In_311);
nor U2098 (N_2098,In_579,In_1913);
nor U2099 (N_2099,In_1795,In_1447);
and U2100 (N_2100,In_1913,In_479);
nand U2101 (N_2101,In_1565,In_913);
nor U2102 (N_2102,In_331,In_1364);
or U2103 (N_2103,In_398,In_21);
nor U2104 (N_2104,In_1657,In_1699);
or U2105 (N_2105,In_345,In_1107);
nand U2106 (N_2106,In_554,In_980);
nand U2107 (N_2107,In_1311,In_1960);
nor U2108 (N_2108,In_1548,In_1354);
xnor U2109 (N_2109,In_805,In_379);
nor U2110 (N_2110,In_1977,In_53);
and U2111 (N_2111,In_65,In_1998);
xor U2112 (N_2112,In_459,In_1367);
or U2113 (N_2113,In_453,In_486);
and U2114 (N_2114,In_319,In_388);
and U2115 (N_2115,In_1934,In_1166);
nor U2116 (N_2116,In_324,In_870);
nor U2117 (N_2117,In_1001,In_1506);
or U2118 (N_2118,In_1709,In_1344);
nand U2119 (N_2119,In_811,In_1421);
nor U2120 (N_2120,In_677,In_638);
nor U2121 (N_2121,In_1332,In_1483);
nor U2122 (N_2122,In_1403,In_1171);
or U2123 (N_2123,In_1230,In_1693);
nor U2124 (N_2124,In_1586,In_1006);
nor U2125 (N_2125,In_1493,In_1007);
and U2126 (N_2126,In_261,In_1839);
and U2127 (N_2127,In_12,In_1039);
and U2128 (N_2128,In_1363,In_745);
or U2129 (N_2129,In_1173,In_682);
nor U2130 (N_2130,In_1447,In_828);
or U2131 (N_2131,In_393,In_1043);
or U2132 (N_2132,In_630,In_34);
or U2133 (N_2133,In_692,In_938);
or U2134 (N_2134,In_1342,In_171);
nor U2135 (N_2135,In_723,In_747);
or U2136 (N_2136,In_240,In_1441);
nor U2137 (N_2137,In_1817,In_1308);
and U2138 (N_2138,In_628,In_1038);
xnor U2139 (N_2139,In_744,In_1799);
or U2140 (N_2140,In_92,In_881);
and U2141 (N_2141,In_1519,In_896);
xor U2142 (N_2142,In_1210,In_436);
or U2143 (N_2143,In_1432,In_1746);
xnor U2144 (N_2144,In_300,In_1930);
nor U2145 (N_2145,In_414,In_534);
or U2146 (N_2146,In_1059,In_1510);
nor U2147 (N_2147,In_9,In_1901);
and U2148 (N_2148,In_1215,In_1319);
nand U2149 (N_2149,In_120,In_1757);
xnor U2150 (N_2150,In_1761,In_504);
nand U2151 (N_2151,In_773,In_800);
xnor U2152 (N_2152,In_1424,In_1869);
or U2153 (N_2153,In_53,In_789);
nor U2154 (N_2154,In_426,In_1312);
and U2155 (N_2155,In_340,In_136);
xor U2156 (N_2156,In_1880,In_901);
or U2157 (N_2157,In_2,In_48);
nand U2158 (N_2158,In_1203,In_425);
and U2159 (N_2159,In_1882,In_623);
xor U2160 (N_2160,In_1279,In_602);
nor U2161 (N_2161,In_738,In_1030);
or U2162 (N_2162,In_428,In_815);
and U2163 (N_2163,In_1819,In_1365);
xnor U2164 (N_2164,In_1929,In_1133);
nand U2165 (N_2165,In_1155,In_964);
nand U2166 (N_2166,In_1286,In_1174);
and U2167 (N_2167,In_932,In_477);
nand U2168 (N_2168,In_1302,In_679);
and U2169 (N_2169,In_1949,In_1223);
xnor U2170 (N_2170,In_110,In_237);
nand U2171 (N_2171,In_30,In_493);
nor U2172 (N_2172,In_640,In_405);
nand U2173 (N_2173,In_709,In_1533);
nor U2174 (N_2174,In_3,In_1972);
nand U2175 (N_2175,In_1530,In_441);
nand U2176 (N_2176,In_1001,In_289);
and U2177 (N_2177,In_1908,In_800);
nand U2178 (N_2178,In_966,In_785);
or U2179 (N_2179,In_778,In_631);
or U2180 (N_2180,In_630,In_1336);
nor U2181 (N_2181,In_1648,In_145);
nand U2182 (N_2182,In_720,In_568);
nand U2183 (N_2183,In_1200,In_294);
nand U2184 (N_2184,In_500,In_27);
and U2185 (N_2185,In_188,In_1531);
nor U2186 (N_2186,In_666,In_1373);
or U2187 (N_2187,In_425,In_301);
nand U2188 (N_2188,In_1571,In_915);
nor U2189 (N_2189,In_1493,In_1692);
and U2190 (N_2190,In_594,In_258);
and U2191 (N_2191,In_1108,In_222);
or U2192 (N_2192,In_745,In_919);
and U2193 (N_2193,In_328,In_70);
and U2194 (N_2194,In_704,In_929);
nand U2195 (N_2195,In_1939,In_631);
nor U2196 (N_2196,In_538,In_249);
nand U2197 (N_2197,In_1517,In_207);
nand U2198 (N_2198,In_575,In_1167);
nand U2199 (N_2199,In_1873,In_753);
and U2200 (N_2200,In_1415,In_389);
nand U2201 (N_2201,In_571,In_1100);
or U2202 (N_2202,In_1730,In_1433);
nand U2203 (N_2203,In_390,In_681);
nand U2204 (N_2204,In_1137,In_322);
nand U2205 (N_2205,In_1412,In_9);
and U2206 (N_2206,In_1827,In_904);
nand U2207 (N_2207,In_1133,In_469);
nand U2208 (N_2208,In_1835,In_387);
and U2209 (N_2209,In_660,In_1344);
xor U2210 (N_2210,In_1895,In_796);
nor U2211 (N_2211,In_1015,In_544);
or U2212 (N_2212,In_314,In_1835);
and U2213 (N_2213,In_171,In_944);
nor U2214 (N_2214,In_18,In_1244);
nor U2215 (N_2215,In_1161,In_1550);
and U2216 (N_2216,In_447,In_929);
nor U2217 (N_2217,In_1018,In_580);
nand U2218 (N_2218,In_954,In_192);
and U2219 (N_2219,In_839,In_1710);
and U2220 (N_2220,In_1416,In_602);
nor U2221 (N_2221,In_1546,In_517);
or U2222 (N_2222,In_754,In_620);
nor U2223 (N_2223,In_1740,In_1403);
nand U2224 (N_2224,In_503,In_876);
and U2225 (N_2225,In_1511,In_587);
nor U2226 (N_2226,In_1540,In_315);
nand U2227 (N_2227,In_499,In_582);
or U2228 (N_2228,In_830,In_1723);
and U2229 (N_2229,In_354,In_904);
nor U2230 (N_2230,In_1103,In_1760);
nor U2231 (N_2231,In_1222,In_39);
nor U2232 (N_2232,In_885,In_1363);
nor U2233 (N_2233,In_731,In_606);
and U2234 (N_2234,In_397,In_1508);
xor U2235 (N_2235,In_1863,In_467);
or U2236 (N_2236,In_1529,In_1093);
and U2237 (N_2237,In_934,In_195);
and U2238 (N_2238,In_856,In_686);
nor U2239 (N_2239,In_182,In_919);
or U2240 (N_2240,In_195,In_1007);
nand U2241 (N_2241,In_289,In_205);
or U2242 (N_2242,In_577,In_89);
nand U2243 (N_2243,In_1675,In_1352);
nor U2244 (N_2244,In_581,In_1769);
or U2245 (N_2245,In_343,In_379);
or U2246 (N_2246,In_1704,In_1677);
nor U2247 (N_2247,In_1470,In_1391);
xnor U2248 (N_2248,In_1710,In_891);
or U2249 (N_2249,In_535,In_209);
nand U2250 (N_2250,In_556,In_1002);
nor U2251 (N_2251,In_1897,In_758);
and U2252 (N_2252,In_1988,In_414);
nand U2253 (N_2253,In_943,In_915);
nor U2254 (N_2254,In_440,In_1508);
and U2255 (N_2255,In_1519,In_1350);
nor U2256 (N_2256,In_117,In_1217);
nand U2257 (N_2257,In_167,In_188);
and U2258 (N_2258,In_1642,In_1508);
xor U2259 (N_2259,In_1049,In_1054);
and U2260 (N_2260,In_1398,In_1789);
nand U2261 (N_2261,In_1632,In_1039);
and U2262 (N_2262,In_1509,In_1059);
or U2263 (N_2263,In_1893,In_1053);
nor U2264 (N_2264,In_747,In_685);
and U2265 (N_2265,In_1974,In_818);
nor U2266 (N_2266,In_1534,In_191);
xor U2267 (N_2267,In_1080,In_1327);
xnor U2268 (N_2268,In_258,In_935);
nor U2269 (N_2269,In_939,In_501);
nand U2270 (N_2270,In_1552,In_430);
and U2271 (N_2271,In_1930,In_227);
nor U2272 (N_2272,In_873,In_966);
nor U2273 (N_2273,In_486,In_1505);
nand U2274 (N_2274,In_606,In_916);
and U2275 (N_2275,In_275,In_464);
and U2276 (N_2276,In_864,In_1880);
and U2277 (N_2277,In_455,In_1087);
and U2278 (N_2278,In_1761,In_773);
or U2279 (N_2279,In_1269,In_1798);
or U2280 (N_2280,In_995,In_236);
nand U2281 (N_2281,In_906,In_1443);
nor U2282 (N_2282,In_1634,In_1499);
nand U2283 (N_2283,In_1201,In_1705);
or U2284 (N_2284,In_1164,In_1004);
and U2285 (N_2285,In_1046,In_1332);
xnor U2286 (N_2286,In_1385,In_394);
or U2287 (N_2287,In_705,In_1840);
nor U2288 (N_2288,In_1088,In_743);
nor U2289 (N_2289,In_1485,In_440);
and U2290 (N_2290,In_823,In_1697);
nand U2291 (N_2291,In_1752,In_1432);
and U2292 (N_2292,In_325,In_524);
or U2293 (N_2293,In_1522,In_1128);
and U2294 (N_2294,In_1007,In_733);
nand U2295 (N_2295,In_260,In_267);
and U2296 (N_2296,In_56,In_409);
or U2297 (N_2297,In_899,In_1155);
or U2298 (N_2298,In_875,In_251);
nor U2299 (N_2299,In_634,In_343);
nand U2300 (N_2300,In_373,In_1386);
nor U2301 (N_2301,In_1607,In_449);
or U2302 (N_2302,In_33,In_334);
nor U2303 (N_2303,In_1812,In_501);
and U2304 (N_2304,In_1560,In_1497);
or U2305 (N_2305,In_1142,In_427);
and U2306 (N_2306,In_1016,In_367);
or U2307 (N_2307,In_76,In_985);
and U2308 (N_2308,In_637,In_1317);
or U2309 (N_2309,In_507,In_344);
and U2310 (N_2310,In_1497,In_731);
or U2311 (N_2311,In_1966,In_432);
nand U2312 (N_2312,In_1497,In_134);
and U2313 (N_2313,In_1545,In_1297);
nor U2314 (N_2314,In_939,In_998);
or U2315 (N_2315,In_301,In_143);
nand U2316 (N_2316,In_250,In_519);
nor U2317 (N_2317,In_1257,In_851);
and U2318 (N_2318,In_1909,In_1876);
and U2319 (N_2319,In_1540,In_1807);
and U2320 (N_2320,In_305,In_1022);
xnor U2321 (N_2321,In_182,In_284);
or U2322 (N_2322,In_646,In_1857);
or U2323 (N_2323,In_996,In_900);
nor U2324 (N_2324,In_526,In_323);
and U2325 (N_2325,In_1516,In_1966);
nand U2326 (N_2326,In_491,In_506);
xnor U2327 (N_2327,In_355,In_1809);
nand U2328 (N_2328,In_1195,In_1453);
nand U2329 (N_2329,In_1852,In_1567);
or U2330 (N_2330,In_124,In_543);
nor U2331 (N_2331,In_1969,In_275);
nor U2332 (N_2332,In_573,In_1231);
xnor U2333 (N_2333,In_833,In_830);
or U2334 (N_2334,In_847,In_1343);
and U2335 (N_2335,In_1237,In_1376);
nand U2336 (N_2336,In_1144,In_1993);
nor U2337 (N_2337,In_958,In_1283);
or U2338 (N_2338,In_1688,In_574);
nor U2339 (N_2339,In_672,In_918);
nor U2340 (N_2340,In_522,In_1517);
and U2341 (N_2341,In_858,In_1963);
or U2342 (N_2342,In_1685,In_872);
and U2343 (N_2343,In_1874,In_1601);
or U2344 (N_2344,In_1643,In_1011);
nor U2345 (N_2345,In_417,In_1707);
nand U2346 (N_2346,In_768,In_1422);
xnor U2347 (N_2347,In_243,In_652);
xor U2348 (N_2348,In_40,In_374);
nor U2349 (N_2349,In_425,In_1879);
nor U2350 (N_2350,In_119,In_1840);
nand U2351 (N_2351,In_1673,In_1324);
and U2352 (N_2352,In_367,In_1724);
and U2353 (N_2353,In_1731,In_1932);
and U2354 (N_2354,In_403,In_405);
and U2355 (N_2355,In_651,In_548);
and U2356 (N_2356,In_1215,In_1063);
or U2357 (N_2357,In_446,In_897);
nand U2358 (N_2358,In_1341,In_1709);
or U2359 (N_2359,In_619,In_1890);
nand U2360 (N_2360,In_395,In_1231);
or U2361 (N_2361,In_710,In_9);
nor U2362 (N_2362,In_762,In_457);
or U2363 (N_2363,In_139,In_1097);
and U2364 (N_2364,In_774,In_3);
and U2365 (N_2365,In_1597,In_684);
nand U2366 (N_2366,In_1151,In_716);
and U2367 (N_2367,In_1487,In_439);
and U2368 (N_2368,In_1087,In_1910);
nand U2369 (N_2369,In_1834,In_62);
nor U2370 (N_2370,In_1183,In_1379);
and U2371 (N_2371,In_1339,In_1220);
or U2372 (N_2372,In_864,In_1634);
nand U2373 (N_2373,In_858,In_391);
nand U2374 (N_2374,In_1868,In_1375);
and U2375 (N_2375,In_1165,In_1188);
nor U2376 (N_2376,In_1438,In_699);
and U2377 (N_2377,In_1709,In_1363);
and U2378 (N_2378,In_1228,In_79);
and U2379 (N_2379,In_1055,In_991);
nand U2380 (N_2380,In_715,In_1367);
or U2381 (N_2381,In_1544,In_843);
nand U2382 (N_2382,In_890,In_1396);
nor U2383 (N_2383,In_558,In_1534);
or U2384 (N_2384,In_537,In_870);
xor U2385 (N_2385,In_1037,In_1268);
or U2386 (N_2386,In_541,In_655);
or U2387 (N_2387,In_1047,In_1724);
and U2388 (N_2388,In_288,In_1068);
nand U2389 (N_2389,In_1266,In_849);
nor U2390 (N_2390,In_1923,In_235);
xnor U2391 (N_2391,In_1037,In_1397);
nand U2392 (N_2392,In_780,In_1113);
or U2393 (N_2393,In_1670,In_277);
nor U2394 (N_2394,In_23,In_888);
or U2395 (N_2395,In_1936,In_1679);
and U2396 (N_2396,In_1739,In_704);
nand U2397 (N_2397,In_312,In_513);
nand U2398 (N_2398,In_1316,In_1012);
nor U2399 (N_2399,In_198,In_1369);
nand U2400 (N_2400,In_1520,In_320);
nand U2401 (N_2401,In_1969,In_1041);
nor U2402 (N_2402,In_1625,In_1622);
and U2403 (N_2403,In_1229,In_833);
nor U2404 (N_2404,In_533,In_1516);
nand U2405 (N_2405,In_1275,In_1331);
xor U2406 (N_2406,In_68,In_633);
xor U2407 (N_2407,In_1826,In_173);
nor U2408 (N_2408,In_191,In_810);
nor U2409 (N_2409,In_264,In_1786);
nand U2410 (N_2410,In_118,In_1206);
nand U2411 (N_2411,In_532,In_1335);
or U2412 (N_2412,In_1112,In_1815);
or U2413 (N_2413,In_1261,In_183);
nor U2414 (N_2414,In_1262,In_1051);
and U2415 (N_2415,In_510,In_1034);
or U2416 (N_2416,In_1342,In_294);
and U2417 (N_2417,In_723,In_1698);
or U2418 (N_2418,In_1379,In_407);
and U2419 (N_2419,In_1542,In_1042);
nand U2420 (N_2420,In_1371,In_171);
xor U2421 (N_2421,In_1808,In_1673);
or U2422 (N_2422,In_658,In_1323);
nor U2423 (N_2423,In_385,In_298);
nor U2424 (N_2424,In_390,In_587);
nand U2425 (N_2425,In_1235,In_1446);
nor U2426 (N_2426,In_1502,In_414);
nand U2427 (N_2427,In_1649,In_538);
xor U2428 (N_2428,In_1198,In_1964);
xnor U2429 (N_2429,In_256,In_1164);
nand U2430 (N_2430,In_56,In_1298);
or U2431 (N_2431,In_238,In_1967);
and U2432 (N_2432,In_682,In_550);
nand U2433 (N_2433,In_1561,In_28);
nor U2434 (N_2434,In_1675,In_332);
nand U2435 (N_2435,In_895,In_1730);
and U2436 (N_2436,In_890,In_167);
nand U2437 (N_2437,In_1221,In_1035);
and U2438 (N_2438,In_1784,In_266);
xnor U2439 (N_2439,In_7,In_686);
nor U2440 (N_2440,In_1196,In_265);
nor U2441 (N_2441,In_1905,In_595);
and U2442 (N_2442,In_1217,In_611);
xor U2443 (N_2443,In_1278,In_1651);
xnor U2444 (N_2444,In_1897,In_677);
nand U2445 (N_2445,In_808,In_661);
or U2446 (N_2446,In_418,In_702);
or U2447 (N_2447,In_879,In_149);
nand U2448 (N_2448,In_1822,In_1995);
and U2449 (N_2449,In_795,In_1391);
and U2450 (N_2450,In_1648,In_1788);
nor U2451 (N_2451,In_1784,In_1227);
xor U2452 (N_2452,In_838,In_1496);
nor U2453 (N_2453,In_249,In_1932);
or U2454 (N_2454,In_1909,In_25);
xor U2455 (N_2455,In_364,In_329);
nand U2456 (N_2456,In_1987,In_1936);
and U2457 (N_2457,In_1001,In_1900);
xor U2458 (N_2458,In_1750,In_498);
nor U2459 (N_2459,In_630,In_386);
xnor U2460 (N_2460,In_1011,In_164);
or U2461 (N_2461,In_1000,In_366);
or U2462 (N_2462,In_946,In_617);
or U2463 (N_2463,In_1677,In_203);
and U2464 (N_2464,In_1044,In_272);
or U2465 (N_2465,In_1163,In_509);
nand U2466 (N_2466,In_992,In_611);
or U2467 (N_2467,In_1305,In_346);
nand U2468 (N_2468,In_1486,In_957);
nand U2469 (N_2469,In_257,In_1019);
xnor U2470 (N_2470,In_827,In_581);
or U2471 (N_2471,In_441,In_1835);
nand U2472 (N_2472,In_884,In_1982);
and U2473 (N_2473,In_1152,In_1533);
and U2474 (N_2474,In_559,In_995);
nor U2475 (N_2475,In_1081,In_1739);
or U2476 (N_2476,In_844,In_1625);
and U2477 (N_2477,In_241,In_37);
nand U2478 (N_2478,In_898,In_983);
and U2479 (N_2479,In_35,In_1335);
nand U2480 (N_2480,In_1694,In_1947);
xnor U2481 (N_2481,In_281,In_642);
nor U2482 (N_2482,In_579,In_888);
nand U2483 (N_2483,In_1418,In_408);
or U2484 (N_2484,In_1378,In_1090);
and U2485 (N_2485,In_36,In_933);
or U2486 (N_2486,In_245,In_336);
nor U2487 (N_2487,In_712,In_190);
or U2488 (N_2488,In_1218,In_1914);
and U2489 (N_2489,In_249,In_39);
and U2490 (N_2490,In_585,In_42);
or U2491 (N_2491,In_1460,In_1850);
xnor U2492 (N_2492,In_1467,In_895);
nand U2493 (N_2493,In_11,In_208);
xnor U2494 (N_2494,In_1622,In_1156);
and U2495 (N_2495,In_229,In_802);
nand U2496 (N_2496,In_343,In_1303);
or U2497 (N_2497,In_1798,In_1412);
or U2498 (N_2498,In_1380,In_484);
nor U2499 (N_2499,In_1441,In_1337);
nand U2500 (N_2500,In_854,In_1598);
or U2501 (N_2501,In_1057,In_799);
and U2502 (N_2502,In_1203,In_740);
or U2503 (N_2503,In_1934,In_1103);
or U2504 (N_2504,In_855,In_50);
and U2505 (N_2505,In_1017,In_1826);
and U2506 (N_2506,In_835,In_1775);
or U2507 (N_2507,In_1089,In_334);
nand U2508 (N_2508,In_989,In_1142);
or U2509 (N_2509,In_1304,In_1870);
or U2510 (N_2510,In_1966,In_438);
and U2511 (N_2511,In_1157,In_90);
and U2512 (N_2512,In_38,In_1967);
nand U2513 (N_2513,In_1997,In_1593);
or U2514 (N_2514,In_723,In_1733);
nand U2515 (N_2515,In_716,In_1050);
nand U2516 (N_2516,In_1625,In_971);
nor U2517 (N_2517,In_1666,In_1163);
nand U2518 (N_2518,In_1770,In_1056);
and U2519 (N_2519,In_1998,In_472);
nor U2520 (N_2520,In_93,In_998);
nand U2521 (N_2521,In_617,In_1219);
and U2522 (N_2522,In_588,In_1614);
nand U2523 (N_2523,In_219,In_1922);
or U2524 (N_2524,In_770,In_746);
and U2525 (N_2525,In_1753,In_1362);
nor U2526 (N_2526,In_998,In_1566);
or U2527 (N_2527,In_532,In_860);
and U2528 (N_2528,In_1619,In_378);
and U2529 (N_2529,In_856,In_1708);
nand U2530 (N_2530,In_260,In_1677);
xnor U2531 (N_2531,In_111,In_1225);
nand U2532 (N_2532,In_1915,In_1264);
or U2533 (N_2533,In_1649,In_1151);
or U2534 (N_2534,In_610,In_1341);
nand U2535 (N_2535,In_1279,In_669);
or U2536 (N_2536,In_877,In_1558);
or U2537 (N_2537,In_1232,In_1282);
nand U2538 (N_2538,In_1335,In_1209);
or U2539 (N_2539,In_868,In_1403);
nand U2540 (N_2540,In_1795,In_793);
nor U2541 (N_2541,In_1982,In_1654);
and U2542 (N_2542,In_1093,In_1361);
nor U2543 (N_2543,In_1516,In_353);
nand U2544 (N_2544,In_808,In_826);
or U2545 (N_2545,In_48,In_445);
or U2546 (N_2546,In_1681,In_1300);
nor U2547 (N_2547,In_128,In_342);
nor U2548 (N_2548,In_730,In_76);
and U2549 (N_2549,In_1568,In_1681);
nand U2550 (N_2550,In_1413,In_678);
nor U2551 (N_2551,In_1802,In_739);
or U2552 (N_2552,In_1897,In_1331);
xor U2553 (N_2553,In_942,In_902);
or U2554 (N_2554,In_641,In_55);
nor U2555 (N_2555,In_1693,In_1187);
or U2556 (N_2556,In_1613,In_380);
nor U2557 (N_2557,In_1343,In_22);
nor U2558 (N_2558,In_1156,In_614);
nand U2559 (N_2559,In_1209,In_1214);
xor U2560 (N_2560,In_1671,In_968);
nor U2561 (N_2561,In_832,In_1652);
and U2562 (N_2562,In_823,In_867);
or U2563 (N_2563,In_685,In_396);
nand U2564 (N_2564,In_208,In_1271);
or U2565 (N_2565,In_1828,In_1294);
nand U2566 (N_2566,In_499,In_415);
and U2567 (N_2567,In_78,In_223);
xor U2568 (N_2568,In_1545,In_1069);
nand U2569 (N_2569,In_1056,In_1009);
nor U2570 (N_2570,In_1337,In_215);
nor U2571 (N_2571,In_1586,In_628);
and U2572 (N_2572,In_580,In_1999);
and U2573 (N_2573,In_1576,In_1613);
or U2574 (N_2574,In_1297,In_1286);
nand U2575 (N_2575,In_1839,In_1319);
nor U2576 (N_2576,In_880,In_742);
or U2577 (N_2577,In_1779,In_134);
nand U2578 (N_2578,In_1024,In_1541);
nand U2579 (N_2579,In_1208,In_732);
and U2580 (N_2580,In_385,In_1333);
nand U2581 (N_2581,In_392,In_1691);
or U2582 (N_2582,In_1183,In_1540);
xnor U2583 (N_2583,In_1643,In_690);
nor U2584 (N_2584,In_1139,In_1276);
nor U2585 (N_2585,In_231,In_1958);
nor U2586 (N_2586,In_1350,In_979);
and U2587 (N_2587,In_142,In_1705);
xor U2588 (N_2588,In_1718,In_1474);
or U2589 (N_2589,In_1061,In_490);
nor U2590 (N_2590,In_366,In_685);
nand U2591 (N_2591,In_1932,In_1339);
or U2592 (N_2592,In_1379,In_205);
or U2593 (N_2593,In_1741,In_430);
nor U2594 (N_2594,In_1360,In_16);
nor U2595 (N_2595,In_1270,In_12);
nand U2596 (N_2596,In_566,In_1628);
nand U2597 (N_2597,In_1414,In_1867);
or U2598 (N_2598,In_115,In_216);
or U2599 (N_2599,In_1733,In_1333);
and U2600 (N_2600,In_1815,In_1964);
xor U2601 (N_2601,In_1352,In_376);
nand U2602 (N_2602,In_826,In_1154);
xor U2603 (N_2603,In_1953,In_436);
and U2604 (N_2604,In_1612,In_1552);
or U2605 (N_2605,In_291,In_724);
nor U2606 (N_2606,In_1212,In_607);
nor U2607 (N_2607,In_761,In_373);
nand U2608 (N_2608,In_152,In_754);
or U2609 (N_2609,In_1083,In_1092);
and U2610 (N_2610,In_512,In_705);
or U2611 (N_2611,In_569,In_1188);
and U2612 (N_2612,In_347,In_407);
and U2613 (N_2613,In_940,In_1981);
or U2614 (N_2614,In_943,In_699);
xnor U2615 (N_2615,In_441,In_587);
or U2616 (N_2616,In_1750,In_139);
or U2617 (N_2617,In_104,In_398);
and U2618 (N_2618,In_956,In_1652);
or U2619 (N_2619,In_978,In_1738);
xor U2620 (N_2620,In_657,In_1377);
or U2621 (N_2621,In_1570,In_342);
xnor U2622 (N_2622,In_1179,In_283);
and U2623 (N_2623,In_1125,In_1481);
nand U2624 (N_2624,In_394,In_745);
nand U2625 (N_2625,In_1379,In_1604);
and U2626 (N_2626,In_1411,In_1617);
nor U2627 (N_2627,In_1707,In_818);
nand U2628 (N_2628,In_1939,In_1187);
nand U2629 (N_2629,In_586,In_1223);
nor U2630 (N_2630,In_1793,In_1721);
or U2631 (N_2631,In_1076,In_1760);
nor U2632 (N_2632,In_402,In_923);
and U2633 (N_2633,In_392,In_655);
or U2634 (N_2634,In_1885,In_1066);
nor U2635 (N_2635,In_1572,In_1737);
or U2636 (N_2636,In_1373,In_1636);
and U2637 (N_2637,In_1348,In_883);
or U2638 (N_2638,In_1177,In_598);
or U2639 (N_2639,In_1463,In_1167);
nand U2640 (N_2640,In_125,In_384);
nor U2641 (N_2641,In_1783,In_1656);
nor U2642 (N_2642,In_445,In_1570);
nor U2643 (N_2643,In_335,In_1965);
nand U2644 (N_2644,In_800,In_1771);
nor U2645 (N_2645,In_1378,In_671);
nor U2646 (N_2646,In_1123,In_277);
and U2647 (N_2647,In_1160,In_212);
nand U2648 (N_2648,In_1510,In_1170);
and U2649 (N_2649,In_166,In_1903);
and U2650 (N_2650,In_314,In_735);
nor U2651 (N_2651,In_1440,In_67);
and U2652 (N_2652,In_1191,In_1477);
nand U2653 (N_2653,In_1191,In_1612);
xnor U2654 (N_2654,In_1674,In_267);
nor U2655 (N_2655,In_1876,In_301);
nor U2656 (N_2656,In_311,In_1847);
and U2657 (N_2657,In_1893,In_403);
xor U2658 (N_2658,In_775,In_1637);
and U2659 (N_2659,In_805,In_981);
xor U2660 (N_2660,In_993,In_481);
or U2661 (N_2661,In_1594,In_390);
xnor U2662 (N_2662,In_1115,In_87);
nand U2663 (N_2663,In_353,In_1807);
nand U2664 (N_2664,In_685,In_1240);
nor U2665 (N_2665,In_664,In_945);
nand U2666 (N_2666,In_166,In_1992);
nor U2667 (N_2667,In_560,In_955);
and U2668 (N_2668,In_1785,In_1896);
xor U2669 (N_2669,In_1127,In_1421);
nand U2670 (N_2670,In_1239,In_1413);
xor U2671 (N_2671,In_1161,In_1997);
or U2672 (N_2672,In_705,In_716);
or U2673 (N_2673,In_1274,In_1500);
or U2674 (N_2674,In_1584,In_1846);
nand U2675 (N_2675,In_905,In_1796);
and U2676 (N_2676,In_1103,In_296);
xnor U2677 (N_2677,In_110,In_416);
and U2678 (N_2678,In_533,In_178);
and U2679 (N_2679,In_1848,In_1187);
and U2680 (N_2680,In_1810,In_375);
or U2681 (N_2681,In_1614,In_992);
xor U2682 (N_2682,In_697,In_1698);
and U2683 (N_2683,In_848,In_1463);
nor U2684 (N_2684,In_1567,In_1865);
xnor U2685 (N_2685,In_1637,In_1007);
nand U2686 (N_2686,In_909,In_667);
nand U2687 (N_2687,In_1093,In_1863);
or U2688 (N_2688,In_851,In_1504);
nor U2689 (N_2689,In_329,In_1868);
or U2690 (N_2690,In_1504,In_274);
nand U2691 (N_2691,In_948,In_246);
nor U2692 (N_2692,In_1490,In_1906);
or U2693 (N_2693,In_1572,In_1041);
nand U2694 (N_2694,In_732,In_905);
nor U2695 (N_2695,In_1365,In_1054);
or U2696 (N_2696,In_777,In_1094);
nand U2697 (N_2697,In_1183,In_1276);
nand U2698 (N_2698,In_753,In_1783);
nor U2699 (N_2699,In_1361,In_1626);
xor U2700 (N_2700,In_890,In_376);
or U2701 (N_2701,In_1338,In_313);
xnor U2702 (N_2702,In_454,In_725);
or U2703 (N_2703,In_1033,In_21);
and U2704 (N_2704,In_635,In_245);
and U2705 (N_2705,In_165,In_1540);
or U2706 (N_2706,In_971,In_437);
and U2707 (N_2707,In_70,In_1738);
nor U2708 (N_2708,In_280,In_1415);
and U2709 (N_2709,In_30,In_598);
or U2710 (N_2710,In_618,In_1490);
nand U2711 (N_2711,In_1670,In_428);
nand U2712 (N_2712,In_1471,In_555);
or U2713 (N_2713,In_1892,In_331);
xnor U2714 (N_2714,In_1891,In_1928);
or U2715 (N_2715,In_1344,In_508);
xor U2716 (N_2716,In_413,In_133);
and U2717 (N_2717,In_203,In_1873);
nor U2718 (N_2718,In_1321,In_1738);
nand U2719 (N_2719,In_887,In_1782);
or U2720 (N_2720,In_213,In_1177);
nand U2721 (N_2721,In_510,In_1676);
nor U2722 (N_2722,In_825,In_212);
nand U2723 (N_2723,In_603,In_1997);
or U2724 (N_2724,In_1167,In_148);
or U2725 (N_2725,In_1816,In_751);
nand U2726 (N_2726,In_1202,In_949);
nand U2727 (N_2727,In_1905,In_396);
or U2728 (N_2728,In_858,In_1204);
and U2729 (N_2729,In_424,In_733);
or U2730 (N_2730,In_1381,In_12);
nand U2731 (N_2731,In_1454,In_1283);
xnor U2732 (N_2732,In_1734,In_99);
nor U2733 (N_2733,In_458,In_268);
nand U2734 (N_2734,In_1861,In_538);
nor U2735 (N_2735,In_1419,In_864);
xor U2736 (N_2736,In_280,In_1411);
nor U2737 (N_2737,In_568,In_1241);
xnor U2738 (N_2738,In_904,In_1549);
nand U2739 (N_2739,In_1823,In_294);
nor U2740 (N_2740,In_84,In_287);
nand U2741 (N_2741,In_1542,In_199);
nor U2742 (N_2742,In_660,In_1082);
nor U2743 (N_2743,In_860,In_1438);
nand U2744 (N_2744,In_244,In_1132);
or U2745 (N_2745,In_1323,In_1525);
nand U2746 (N_2746,In_1903,In_1725);
nor U2747 (N_2747,In_903,In_1569);
or U2748 (N_2748,In_1371,In_1863);
nand U2749 (N_2749,In_307,In_315);
nand U2750 (N_2750,In_201,In_1503);
or U2751 (N_2751,In_990,In_1021);
xor U2752 (N_2752,In_196,In_504);
nand U2753 (N_2753,In_422,In_1478);
or U2754 (N_2754,In_1021,In_1999);
nor U2755 (N_2755,In_516,In_608);
nand U2756 (N_2756,In_1169,In_63);
nor U2757 (N_2757,In_1248,In_1564);
and U2758 (N_2758,In_884,In_1238);
xnor U2759 (N_2759,In_178,In_1795);
or U2760 (N_2760,In_1688,In_1263);
nor U2761 (N_2761,In_1399,In_944);
and U2762 (N_2762,In_829,In_843);
nand U2763 (N_2763,In_754,In_1505);
nand U2764 (N_2764,In_1107,In_680);
and U2765 (N_2765,In_1537,In_1208);
and U2766 (N_2766,In_1954,In_1360);
and U2767 (N_2767,In_735,In_1806);
nand U2768 (N_2768,In_1526,In_1780);
and U2769 (N_2769,In_944,In_165);
and U2770 (N_2770,In_165,In_600);
xnor U2771 (N_2771,In_954,In_1865);
nor U2772 (N_2772,In_712,In_476);
nand U2773 (N_2773,In_109,In_1448);
xor U2774 (N_2774,In_1502,In_556);
or U2775 (N_2775,In_1006,In_326);
nor U2776 (N_2776,In_1663,In_1146);
nand U2777 (N_2777,In_1764,In_1603);
nand U2778 (N_2778,In_354,In_1270);
nand U2779 (N_2779,In_1985,In_1508);
and U2780 (N_2780,In_1822,In_403);
xor U2781 (N_2781,In_1715,In_1657);
and U2782 (N_2782,In_110,In_52);
nor U2783 (N_2783,In_1395,In_230);
nor U2784 (N_2784,In_800,In_1533);
or U2785 (N_2785,In_318,In_1779);
nand U2786 (N_2786,In_373,In_787);
nand U2787 (N_2787,In_1624,In_1875);
nor U2788 (N_2788,In_797,In_1315);
and U2789 (N_2789,In_202,In_885);
or U2790 (N_2790,In_455,In_959);
or U2791 (N_2791,In_1667,In_1444);
nand U2792 (N_2792,In_1488,In_698);
and U2793 (N_2793,In_855,In_1190);
or U2794 (N_2794,In_574,In_14);
nor U2795 (N_2795,In_1544,In_551);
nand U2796 (N_2796,In_984,In_550);
or U2797 (N_2797,In_1096,In_1004);
nor U2798 (N_2798,In_1394,In_1595);
nand U2799 (N_2799,In_1837,In_1890);
or U2800 (N_2800,In_1596,In_1410);
and U2801 (N_2801,In_834,In_1313);
nor U2802 (N_2802,In_92,In_605);
or U2803 (N_2803,In_1418,In_1361);
nand U2804 (N_2804,In_1579,In_1166);
nor U2805 (N_2805,In_1218,In_1342);
xor U2806 (N_2806,In_1846,In_1222);
nand U2807 (N_2807,In_1562,In_712);
and U2808 (N_2808,In_909,In_773);
and U2809 (N_2809,In_1615,In_1357);
and U2810 (N_2810,In_1136,In_1123);
nand U2811 (N_2811,In_1410,In_1666);
nor U2812 (N_2812,In_1281,In_390);
nor U2813 (N_2813,In_1600,In_262);
nor U2814 (N_2814,In_1411,In_94);
nor U2815 (N_2815,In_1937,In_201);
or U2816 (N_2816,In_1876,In_1644);
nor U2817 (N_2817,In_1426,In_336);
nand U2818 (N_2818,In_921,In_557);
or U2819 (N_2819,In_1997,In_1507);
and U2820 (N_2820,In_149,In_1870);
or U2821 (N_2821,In_1103,In_206);
or U2822 (N_2822,In_1954,In_366);
nor U2823 (N_2823,In_934,In_1251);
and U2824 (N_2824,In_528,In_811);
nand U2825 (N_2825,In_1078,In_244);
nand U2826 (N_2826,In_362,In_921);
xor U2827 (N_2827,In_331,In_515);
or U2828 (N_2828,In_811,In_1891);
and U2829 (N_2829,In_302,In_937);
or U2830 (N_2830,In_367,In_1873);
nand U2831 (N_2831,In_708,In_473);
nand U2832 (N_2832,In_111,In_1257);
or U2833 (N_2833,In_228,In_1490);
nand U2834 (N_2834,In_600,In_900);
xor U2835 (N_2835,In_454,In_75);
nand U2836 (N_2836,In_1284,In_1339);
and U2837 (N_2837,In_581,In_1383);
nor U2838 (N_2838,In_1260,In_1593);
and U2839 (N_2839,In_1117,In_659);
or U2840 (N_2840,In_1521,In_551);
or U2841 (N_2841,In_212,In_1890);
nand U2842 (N_2842,In_1457,In_123);
or U2843 (N_2843,In_161,In_1533);
nand U2844 (N_2844,In_1112,In_1938);
xor U2845 (N_2845,In_1833,In_1590);
nor U2846 (N_2846,In_1969,In_1321);
or U2847 (N_2847,In_1694,In_1397);
and U2848 (N_2848,In_1526,In_368);
or U2849 (N_2849,In_1970,In_865);
or U2850 (N_2850,In_1711,In_961);
nand U2851 (N_2851,In_1776,In_1767);
or U2852 (N_2852,In_333,In_370);
nor U2853 (N_2853,In_901,In_805);
nor U2854 (N_2854,In_1597,In_1669);
nor U2855 (N_2855,In_1744,In_1086);
nand U2856 (N_2856,In_107,In_621);
or U2857 (N_2857,In_265,In_896);
and U2858 (N_2858,In_243,In_371);
nor U2859 (N_2859,In_1861,In_1687);
nand U2860 (N_2860,In_1326,In_14);
xor U2861 (N_2861,In_1973,In_924);
or U2862 (N_2862,In_1032,In_1989);
nor U2863 (N_2863,In_299,In_556);
and U2864 (N_2864,In_1380,In_1515);
nand U2865 (N_2865,In_811,In_665);
or U2866 (N_2866,In_1240,In_1006);
or U2867 (N_2867,In_425,In_1485);
nor U2868 (N_2868,In_382,In_1329);
nor U2869 (N_2869,In_387,In_818);
nand U2870 (N_2870,In_1367,In_688);
and U2871 (N_2871,In_1482,In_1344);
nor U2872 (N_2872,In_1241,In_1385);
xnor U2873 (N_2873,In_1814,In_690);
xor U2874 (N_2874,In_704,In_1400);
nand U2875 (N_2875,In_1047,In_1346);
nand U2876 (N_2876,In_731,In_1345);
or U2877 (N_2877,In_1201,In_1998);
nor U2878 (N_2878,In_437,In_1200);
and U2879 (N_2879,In_381,In_112);
nor U2880 (N_2880,In_1838,In_136);
nand U2881 (N_2881,In_1802,In_491);
xnor U2882 (N_2882,In_1283,In_494);
nand U2883 (N_2883,In_553,In_249);
and U2884 (N_2884,In_100,In_1648);
or U2885 (N_2885,In_253,In_1807);
or U2886 (N_2886,In_1679,In_596);
nor U2887 (N_2887,In_1285,In_137);
or U2888 (N_2888,In_1661,In_1755);
or U2889 (N_2889,In_633,In_1786);
and U2890 (N_2890,In_1382,In_826);
nand U2891 (N_2891,In_572,In_591);
or U2892 (N_2892,In_246,In_1328);
and U2893 (N_2893,In_1329,In_1768);
and U2894 (N_2894,In_1232,In_382);
nor U2895 (N_2895,In_1334,In_169);
or U2896 (N_2896,In_1501,In_883);
nand U2897 (N_2897,In_334,In_94);
nor U2898 (N_2898,In_305,In_953);
nor U2899 (N_2899,In_446,In_381);
nand U2900 (N_2900,In_401,In_926);
or U2901 (N_2901,In_184,In_430);
or U2902 (N_2902,In_634,In_913);
xnor U2903 (N_2903,In_707,In_1939);
nand U2904 (N_2904,In_1131,In_1632);
and U2905 (N_2905,In_1427,In_811);
nor U2906 (N_2906,In_1368,In_240);
or U2907 (N_2907,In_681,In_1923);
or U2908 (N_2908,In_1414,In_524);
nand U2909 (N_2909,In_1715,In_598);
and U2910 (N_2910,In_598,In_751);
or U2911 (N_2911,In_793,In_1714);
and U2912 (N_2912,In_1481,In_1855);
and U2913 (N_2913,In_1415,In_1197);
nor U2914 (N_2914,In_1309,In_626);
or U2915 (N_2915,In_1259,In_1187);
and U2916 (N_2916,In_1968,In_1998);
nand U2917 (N_2917,In_1778,In_922);
nor U2918 (N_2918,In_439,In_535);
nand U2919 (N_2919,In_1200,In_187);
nand U2920 (N_2920,In_1563,In_828);
nand U2921 (N_2921,In_1011,In_1493);
xnor U2922 (N_2922,In_47,In_735);
xor U2923 (N_2923,In_609,In_1159);
xnor U2924 (N_2924,In_1336,In_395);
and U2925 (N_2925,In_1293,In_1130);
xor U2926 (N_2926,In_1035,In_1060);
and U2927 (N_2927,In_660,In_513);
nor U2928 (N_2928,In_53,In_104);
nand U2929 (N_2929,In_616,In_76);
nor U2930 (N_2930,In_397,In_1350);
or U2931 (N_2931,In_1221,In_1224);
xor U2932 (N_2932,In_1376,In_855);
or U2933 (N_2933,In_58,In_1581);
nand U2934 (N_2934,In_617,In_614);
nand U2935 (N_2935,In_1969,In_86);
nor U2936 (N_2936,In_1827,In_312);
nand U2937 (N_2937,In_25,In_254);
xor U2938 (N_2938,In_1491,In_993);
nand U2939 (N_2939,In_1816,In_661);
or U2940 (N_2940,In_234,In_555);
nor U2941 (N_2941,In_1499,In_847);
nor U2942 (N_2942,In_103,In_1594);
nor U2943 (N_2943,In_1167,In_1566);
or U2944 (N_2944,In_120,In_1702);
nand U2945 (N_2945,In_134,In_618);
xnor U2946 (N_2946,In_1615,In_213);
or U2947 (N_2947,In_257,In_1249);
nor U2948 (N_2948,In_1173,In_334);
nor U2949 (N_2949,In_609,In_1604);
nor U2950 (N_2950,In_1572,In_1863);
or U2951 (N_2951,In_599,In_405);
and U2952 (N_2952,In_973,In_355);
xnor U2953 (N_2953,In_1537,In_1222);
nand U2954 (N_2954,In_1238,In_1839);
and U2955 (N_2955,In_264,In_1384);
nand U2956 (N_2956,In_1728,In_1858);
nor U2957 (N_2957,In_321,In_1238);
xnor U2958 (N_2958,In_1685,In_997);
xor U2959 (N_2959,In_564,In_384);
nor U2960 (N_2960,In_280,In_907);
or U2961 (N_2961,In_1642,In_1212);
and U2962 (N_2962,In_1872,In_693);
nor U2963 (N_2963,In_936,In_1506);
nor U2964 (N_2964,In_221,In_874);
nand U2965 (N_2965,In_505,In_1740);
nor U2966 (N_2966,In_1044,In_1329);
and U2967 (N_2967,In_500,In_155);
and U2968 (N_2968,In_284,In_45);
and U2969 (N_2969,In_1446,In_856);
or U2970 (N_2970,In_1864,In_1168);
or U2971 (N_2971,In_131,In_218);
nor U2972 (N_2972,In_1619,In_432);
and U2973 (N_2973,In_106,In_942);
nor U2974 (N_2974,In_1747,In_1218);
nand U2975 (N_2975,In_1747,In_1801);
nand U2976 (N_2976,In_1387,In_764);
nand U2977 (N_2977,In_1970,In_698);
nand U2978 (N_2978,In_40,In_1454);
and U2979 (N_2979,In_1008,In_1540);
and U2980 (N_2980,In_15,In_339);
nand U2981 (N_2981,In_1892,In_1449);
and U2982 (N_2982,In_561,In_1807);
and U2983 (N_2983,In_616,In_1410);
and U2984 (N_2984,In_296,In_815);
and U2985 (N_2985,In_1411,In_233);
nor U2986 (N_2986,In_865,In_1670);
and U2987 (N_2987,In_1152,In_932);
or U2988 (N_2988,In_425,In_1543);
nor U2989 (N_2989,In_1407,In_689);
nor U2990 (N_2990,In_1879,In_1550);
nand U2991 (N_2991,In_1473,In_1976);
and U2992 (N_2992,In_1575,In_17);
nor U2993 (N_2993,In_1152,In_1807);
and U2994 (N_2994,In_1049,In_1067);
or U2995 (N_2995,In_1740,In_1463);
nand U2996 (N_2996,In_1571,In_394);
nor U2997 (N_2997,In_1509,In_714);
nand U2998 (N_2998,In_816,In_297);
or U2999 (N_2999,In_1290,In_541);
xor U3000 (N_3000,In_906,In_78);
nor U3001 (N_3001,In_974,In_41);
xnor U3002 (N_3002,In_712,In_1330);
or U3003 (N_3003,In_1905,In_1813);
nor U3004 (N_3004,In_1829,In_1650);
nor U3005 (N_3005,In_390,In_470);
nor U3006 (N_3006,In_1477,In_188);
and U3007 (N_3007,In_310,In_148);
and U3008 (N_3008,In_1017,In_1429);
or U3009 (N_3009,In_218,In_1058);
nor U3010 (N_3010,In_605,In_1642);
nand U3011 (N_3011,In_242,In_1981);
nor U3012 (N_3012,In_1481,In_198);
nand U3013 (N_3013,In_1587,In_1739);
nand U3014 (N_3014,In_1176,In_630);
nor U3015 (N_3015,In_999,In_1618);
and U3016 (N_3016,In_1929,In_1338);
and U3017 (N_3017,In_506,In_791);
and U3018 (N_3018,In_1024,In_646);
and U3019 (N_3019,In_135,In_1085);
xor U3020 (N_3020,In_1359,In_1397);
nand U3021 (N_3021,In_1488,In_1457);
xor U3022 (N_3022,In_550,In_137);
or U3023 (N_3023,In_1481,In_587);
nand U3024 (N_3024,In_1492,In_1059);
and U3025 (N_3025,In_1801,In_680);
nor U3026 (N_3026,In_1830,In_860);
nor U3027 (N_3027,In_824,In_815);
nand U3028 (N_3028,In_277,In_273);
xnor U3029 (N_3029,In_310,In_1394);
and U3030 (N_3030,In_1478,In_1136);
nor U3031 (N_3031,In_190,In_1436);
nand U3032 (N_3032,In_1358,In_731);
or U3033 (N_3033,In_1611,In_1088);
and U3034 (N_3034,In_1748,In_1782);
nand U3035 (N_3035,In_541,In_1210);
or U3036 (N_3036,In_1989,In_654);
and U3037 (N_3037,In_1364,In_797);
nor U3038 (N_3038,In_1433,In_1732);
or U3039 (N_3039,In_24,In_201);
nand U3040 (N_3040,In_1437,In_1826);
nand U3041 (N_3041,In_844,In_1097);
nand U3042 (N_3042,In_921,In_1454);
nand U3043 (N_3043,In_526,In_68);
nor U3044 (N_3044,In_1075,In_1997);
and U3045 (N_3045,In_1580,In_438);
or U3046 (N_3046,In_461,In_56);
and U3047 (N_3047,In_1157,In_446);
nor U3048 (N_3048,In_1443,In_1549);
nor U3049 (N_3049,In_928,In_583);
and U3050 (N_3050,In_1731,In_707);
and U3051 (N_3051,In_1718,In_733);
and U3052 (N_3052,In_1082,In_96);
nand U3053 (N_3053,In_296,In_1525);
xnor U3054 (N_3054,In_1390,In_908);
or U3055 (N_3055,In_229,In_897);
or U3056 (N_3056,In_462,In_29);
or U3057 (N_3057,In_522,In_1678);
and U3058 (N_3058,In_185,In_992);
xnor U3059 (N_3059,In_1436,In_1567);
and U3060 (N_3060,In_473,In_1968);
and U3061 (N_3061,In_1064,In_1950);
or U3062 (N_3062,In_125,In_997);
nand U3063 (N_3063,In_436,In_1255);
or U3064 (N_3064,In_1811,In_1169);
nand U3065 (N_3065,In_1087,In_241);
and U3066 (N_3066,In_1052,In_1888);
and U3067 (N_3067,In_1663,In_1319);
or U3068 (N_3068,In_382,In_1591);
and U3069 (N_3069,In_979,In_473);
and U3070 (N_3070,In_1207,In_1847);
nor U3071 (N_3071,In_175,In_912);
or U3072 (N_3072,In_1050,In_643);
nor U3073 (N_3073,In_1806,In_1744);
nor U3074 (N_3074,In_34,In_1596);
or U3075 (N_3075,In_1710,In_1673);
and U3076 (N_3076,In_476,In_1558);
nor U3077 (N_3077,In_1731,In_295);
nand U3078 (N_3078,In_372,In_568);
and U3079 (N_3079,In_278,In_1403);
nand U3080 (N_3080,In_1943,In_92);
or U3081 (N_3081,In_489,In_1089);
or U3082 (N_3082,In_960,In_724);
or U3083 (N_3083,In_60,In_1130);
and U3084 (N_3084,In_218,In_1274);
nor U3085 (N_3085,In_1330,In_1135);
or U3086 (N_3086,In_1481,In_1653);
nor U3087 (N_3087,In_1312,In_352);
nand U3088 (N_3088,In_1713,In_328);
or U3089 (N_3089,In_510,In_28);
and U3090 (N_3090,In_58,In_946);
or U3091 (N_3091,In_1538,In_872);
and U3092 (N_3092,In_396,In_484);
nand U3093 (N_3093,In_353,In_28);
nor U3094 (N_3094,In_1705,In_1703);
nor U3095 (N_3095,In_1059,In_441);
nor U3096 (N_3096,In_1226,In_1622);
nand U3097 (N_3097,In_1397,In_1210);
nor U3098 (N_3098,In_942,In_90);
or U3099 (N_3099,In_1604,In_711);
or U3100 (N_3100,In_526,In_821);
and U3101 (N_3101,In_1062,In_478);
nor U3102 (N_3102,In_1370,In_1421);
nand U3103 (N_3103,In_794,In_1438);
xor U3104 (N_3104,In_598,In_1843);
xnor U3105 (N_3105,In_228,In_100);
and U3106 (N_3106,In_1360,In_1514);
or U3107 (N_3107,In_117,In_548);
nor U3108 (N_3108,In_377,In_1573);
and U3109 (N_3109,In_1275,In_826);
or U3110 (N_3110,In_1552,In_47);
nand U3111 (N_3111,In_1928,In_790);
nand U3112 (N_3112,In_1763,In_1940);
and U3113 (N_3113,In_1852,In_275);
and U3114 (N_3114,In_987,In_85);
nor U3115 (N_3115,In_507,In_741);
or U3116 (N_3116,In_471,In_1410);
nand U3117 (N_3117,In_441,In_869);
nor U3118 (N_3118,In_1376,In_1899);
nor U3119 (N_3119,In_1909,In_1525);
nor U3120 (N_3120,In_393,In_131);
nor U3121 (N_3121,In_827,In_995);
or U3122 (N_3122,In_769,In_642);
xnor U3123 (N_3123,In_1899,In_667);
and U3124 (N_3124,In_1920,In_1182);
xnor U3125 (N_3125,In_1279,In_1362);
nor U3126 (N_3126,In_1642,In_672);
nand U3127 (N_3127,In_836,In_1547);
nand U3128 (N_3128,In_1128,In_823);
or U3129 (N_3129,In_705,In_768);
xnor U3130 (N_3130,In_733,In_241);
or U3131 (N_3131,In_1180,In_260);
nand U3132 (N_3132,In_1900,In_690);
nor U3133 (N_3133,In_1883,In_1125);
nor U3134 (N_3134,In_1546,In_990);
and U3135 (N_3135,In_1030,In_1044);
or U3136 (N_3136,In_1612,In_618);
or U3137 (N_3137,In_1149,In_1887);
nand U3138 (N_3138,In_1254,In_1649);
nor U3139 (N_3139,In_1427,In_1282);
or U3140 (N_3140,In_1932,In_1978);
nand U3141 (N_3141,In_454,In_1119);
nand U3142 (N_3142,In_384,In_1170);
xnor U3143 (N_3143,In_1050,In_324);
nor U3144 (N_3144,In_1718,In_356);
nand U3145 (N_3145,In_156,In_405);
nor U3146 (N_3146,In_901,In_269);
and U3147 (N_3147,In_1204,In_966);
and U3148 (N_3148,In_1532,In_1883);
and U3149 (N_3149,In_661,In_1066);
or U3150 (N_3150,In_232,In_1573);
nor U3151 (N_3151,In_303,In_1506);
nor U3152 (N_3152,In_17,In_1922);
or U3153 (N_3153,In_812,In_224);
nand U3154 (N_3154,In_43,In_601);
or U3155 (N_3155,In_1807,In_1606);
or U3156 (N_3156,In_815,In_267);
nand U3157 (N_3157,In_1096,In_1003);
nor U3158 (N_3158,In_811,In_868);
xor U3159 (N_3159,In_492,In_1725);
nand U3160 (N_3160,In_1743,In_1897);
nor U3161 (N_3161,In_1249,In_1015);
nand U3162 (N_3162,In_861,In_288);
or U3163 (N_3163,In_951,In_404);
or U3164 (N_3164,In_1701,In_753);
or U3165 (N_3165,In_1673,In_1877);
xnor U3166 (N_3166,In_92,In_931);
or U3167 (N_3167,In_252,In_1676);
and U3168 (N_3168,In_17,In_324);
nand U3169 (N_3169,In_373,In_1753);
nand U3170 (N_3170,In_1834,In_339);
or U3171 (N_3171,In_1888,In_1901);
nand U3172 (N_3172,In_607,In_219);
nand U3173 (N_3173,In_1498,In_993);
xnor U3174 (N_3174,In_469,In_1579);
nor U3175 (N_3175,In_1078,In_1711);
or U3176 (N_3176,In_392,In_681);
and U3177 (N_3177,In_412,In_1066);
nand U3178 (N_3178,In_1569,In_27);
and U3179 (N_3179,In_219,In_1978);
nand U3180 (N_3180,In_1979,In_1726);
nor U3181 (N_3181,In_1036,In_1463);
nor U3182 (N_3182,In_812,In_1773);
or U3183 (N_3183,In_1268,In_578);
nand U3184 (N_3184,In_1478,In_373);
and U3185 (N_3185,In_882,In_1618);
nand U3186 (N_3186,In_736,In_624);
nand U3187 (N_3187,In_1564,In_1907);
and U3188 (N_3188,In_1435,In_574);
nor U3189 (N_3189,In_452,In_98);
nand U3190 (N_3190,In_783,In_212);
nor U3191 (N_3191,In_1324,In_1621);
nor U3192 (N_3192,In_714,In_1739);
or U3193 (N_3193,In_493,In_1044);
nor U3194 (N_3194,In_1477,In_35);
nor U3195 (N_3195,In_1117,In_202);
and U3196 (N_3196,In_943,In_1352);
or U3197 (N_3197,In_962,In_1936);
and U3198 (N_3198,In_1687,In_457);
nand U3199 (N_3199,In_1939,In_1137);
nor U3200 (N_3200,In_99,In_805);
and U3201 (N_3201,In_730,In_48);
nand U3202 (N_3202,In_1301,In_670);
and U3203 (N_3203,In_1935,In_1190);
or U3204 (N_3204,In_161,In_167);
nor U3205 (N_3205,In_1891,In_1321);
xor U3206 (N_3206,In_1564,In_1578);
and U3207 (N_3207,In_1923,In_1547);
nor U3208 (N_3208,In_1865,In_1893);
nor U3209 (N_3209,In_405,In_411);
and U3210 (N_3210,In_194,In_1240);
and U3211 (N_3211,In_1084,In_1227);
xor U3212 (N_3212,In_138,In_606);
or U3213 (N_3213,In_333,In_1888);
xor U3214 (N_3214,In_613,In_1880);
nor U3215 (N_3215,In_1475,In_1455);
nor U3216 (N_3216,In_1914,In_1731);
xnor U3217 (N_3217,In_488,In_1023);
or U3218 (N_3218,In_992,In_45);
and U3219 (N_3219,In_1156,In_1719);
nand U3220 (N_3220,In_950,In_451);
nand U3221 (N_3221,In_347,In_594);
nand U3222 (N_3222,In_1216,In_1934);
nor U3223 (N_3223,In_379,In_526);
nand U3224 (N_3224,In_1812,In_1968);
nand U3225 (N_3225,In_1702,In_232);
or U3226 (N_3226,In_433,In_1210);
nor U3227 (N_3227,In_1354,In_1650);
xor U3228 (N_3228,In_200,In_1387);
nor U3229 (N_3229,In_446,In_1489);
and U3230 (N_3230,In_1334,In_1337);
and U3231 (N_3231,In_114,In_80);
and U3232 (N_3232,In_970,In_250);
nand U3233 (N_3233,In_598,In_179);
and U3234 (N_3234,In_655,In_1161);
nor U3235 (N_3235,In_1213,In_1613);
nor U3236 (N_3236,In_175,In_256);
nor U3237 (N_3237,In_519,In_131);
nand U3238 (N_3238,In_1696,In_1508);
and U3239 (N_3239,In_818,In_364);
or U3240 (N_3240,In_1335,In_514);
xnor U3241 (N_3241,In_1825,In_1083);
and U3242 (N_3242,In_1452,In_438);
or U3243 (N_3243,In_627,In_747);
nor U3244 (N_3244,In_830,In_323);
or U3245 (N_3245,In_932,In_1277);
or U3246 (N_3246,In_784,In_1396);
nor U3247 (N_3247,In_48,In_1971);
nor U3248 (N_3248,In_1868,In_1026);
xnor U3249 (N_3249,In_1924,In_1774);
nand U3250 (N_3250,In_1413,In_1490);
nor U3251 (N_3251,In_21,In_25);
and U3252 (N_3252,In_509,In_1551);
xnor U3253 (N_3253,In_118,In_305);
and U3254 (N_3254,In_781,In_46);
or U3255 (N_3255,In_1888,In_689);
and U3256 (N_3256,In_57,In_77);
nand U3257 (N_3257,In_1074,In_545);
nand U3258 (N_3258,In_1866,In_1852);
xnor U3259 (N_3259,In_719,In_699);
and U3260 (N_3260,In_669,In_634);
nor U3261 (N_3261,In_1896,In_1350);
and U3262 (N_3262,In_1191,In_1178);
or U3263 (N_3263,In_735,In_1495);
nand U3264 (N_3264,In_369,In_394);
or U3265 (N_3265,In_1271,In_37);
nand U3266 (N_3266,In_1969,In_1068);
and U3267 (N_3267,In_641,In_1457);
nor U3268 (N_3268,In_1607,In_1136);
and U3269 (N_3269,In_882,In_1576);
nand U3270 (N_3270,In_677,In_1819);
nor U3271 (N_3271,In_1472,In_173);
and U3272 (N_3272,In_300,In_317);
or U3273 (N_3273,In_1873,In_1746);
or U3274 (N_3274,In_1098,In_1725);
and U3275 (N_3275,In_1604,In_290);
or U3276 (N_3276,In_527,In_1900);
nand U3277 (N_3277,In_1837,In_1096);
nand U3278 (N_3278,In_1326,In_1180);
nand U3279 (N_3279,In_1623,In_314);
nor U3280 (N_3280,In_472,In_42);
or U3281 (N_3281,In_1169,In_819);
nand U3282 (N_3282,In_304,In_1223);
and U3283 (N_3283,In_1147,In_552);
or U3284 (N_3284,In_300,In_1002);
and U3285 (N_3285,In_1125,In_1732);
xor U3286 (N_3286,In_1091,In_789);
nand U3287 (N_3287,In_1834,In_1596);
nand U3288 (N_3288,In_1256,In_372);
or U3289 (N_3289,In_1619,In_780);
or U3290 (N_3290,In_511,In_1379);
and U3291 (N_3291,In_240,In_291);
or U3292 (N_3292,In_296,In_439);
nand U3293 (N_3293,In_434,In_760);
and U3294 (N_3294,In_680,In_359);
and U3295 (N_3295,In_566,In_1136);
xnor U3296 (N_3296,In_229,In_471);
xnor U3297 (N_3297,In_1609,In_1034);
and U3298 (N_3298,In_1173,In_1107);
nor U3299 (N_3299,In_1453,In_1788);
nand U3300 (N_3300,In_478,In_201);
nand U3301 (N_3301,In_602,In_1537);
and U3302 (N_3302,In_125,In_375);
and U3303 (N_3303,In_1375,In_778);
nor U3304 (N_3304,In_345,In_1156);
xnor U3305 (N_3305,In_1527,In_664);
or U3306 (N_3306,In_301,In_642);
nand U3307 (N_3307,In_404,In_1965);
or U3308 (N_3308,In_1232,In_928);
or U3309 (N_3309,In_1614,In_704);
nor U3310 (N_3310,In_339,In_1042);
or U3311 (N_3311,In_579,In_1855);
or U3312 (N_3312,In_1348,In_1392);
and U3313 (N_3313,In_1373,In_25);
or U3314 (N_3314,In_985,In_1355);
nand U3315 (N_3315,In_1724,In_1900);
or U3316 (N_3316,In_93,In_1700);
xnor U3317 (N_3317,In_656,In_846);
nand U3318 (N_3318,In_28,In_1893);
nand U3319 (N_3319,In_409,In_1444);
or U3320 (N_3320,In_1881,In_555);
and U3321 (N_3321,In_36,In_1624);
nor U3322 (N_3322,In_415,In_1298);
or U3323 (N_3323,In_728,In_820);
or U3324 (N_3324,In_161,In_1704);
and U3325 (N_3325,In_339,In_231);
nor U3326 (N_3326,In_1399,In_1010);
nand U3327 (N_3327,In_750,In_1587);
or U3328 (N_3328,In_1316,In_195);
nor U3329 (N_3329,In_1995,In_1839);
nor U3330 (N_3330,In_580,In_503);
nor U3331 (N_3331,In_800,In_1382);
nand U3332 (N_3332,In_1348,In_1065);
or U3333 (N_3333,In_974,In_922);
nand U3334 (N_3334,In_375,In_881);
nor U3335 (N_3335,In_368,In_830);
and U3336 (N_3336,In_1455,In_1072);
or U3337 (N_3337,In_1960,In_17);
or U3338 (N_3338,In_1637,In_497);
nand U3339 (N_3339,In_1338,In_970);
or U3340 (N_3340,In_245,In_812);
nand U3341 (N_3341,In_1792,In_200);
nand U3342 (N_3342,In_204,In_1073);
and U3343 (N_3343,In_766,In_1611);
nor U3344 (N_3344,In_438,In_1834);
nor U3345 (N_3345,In_1832,In_746);
or U3346 (N_3346,In_884,In_1116);
nand U3347 (N_3347,In_1674,In_627);
nand U3348 (N_3348,In_1239,In_185);
and U3349 (N_3349,In_612,In_307);
and U3350 (N_3350,In_176,In_1176);
nand U3351 (N_3351,In_1548,In_560);
nand U3352 (N_3352,In_994,In_1307);
xor U3353 (N_3353,In_1169,In_1741);
nor U3354 (N_3354,In_57,In_495);
and U3355 (N_3355,In_914,In_416);
nor U3356 (N_3356,In_157,In_607);
and U3357 (N_3357,In_470,In_774);
or U3358 (N_3358,In_1367,In_1960);
nor U3359 (N_3359,In_1691,In_1158);
or U3360 (N_3360,In_644,In_258);
and U3361 (N_3361,In_1549,In_1603);
nor U3362 (N_3362,In_1864,In_183);
or U3363 (N_3363,In_1879,In_1886);
xor U3364 (N_3364,In_513,In_1425);
or U3365 (N_3365,In_1932,In_1143);
and U3366 (N_3366,In_1221,In_1050);
and U3367 (N_3367,In_1166,In_1774);
or U3368 (N_3368,In_265,In_1603);
and U3369 (N_3369,In_719,In_1732);
or U3370 (N_3370,In_997,In_674);
and U3371 (N_3371,In_244,In_292);
and U3372 (N_3372,In_772,In_804);
xnor U3373 (N_3373,In_27,In_323);
and U3374 (N_3374,In_1487,In_1647);
or U3375 (N_3375,In_1737,In_5);
xnor U3376 (N_3376,In_1293,In_864);
and U3377 (N_3377,In_1883,In_1053);
nand U3378 (N_3378,In_746,In_1980);
or U3379 (N_3379,In_680,In_947);
or U3380 (N_3380,In_1900,In_1190);
or U3381 (N_3381,In_364,In_128);
xnor U3382 (N_3382,In_1488,In_1246);
or U3383 (N_3383,In_1643,In_791);
and U3384 (N_3384,In_789,In_164);
nand U3385 (N_3385,In_981,In_1195);
nand U3386 (N_3386,In_647,In_1610);
and U3387 (N_3387,In_4,In_1535);
or U3388 (N_3388,In_470,In_1371);
and U3389 (N_3389,In_1009,In_1586);
or U3390 (N_3390,In_739,In_993);
nand U3391 (N_3391,In_1525,In_1197);
or U3392 (N_3392,In_1467,In_1567);
nor U3393 (N_3393,In_1589,In_226);
xnor U3394 (N_3394,In_1410,In_583);
nand U3395 (N_3395,In_10,In_1345);
nor U3396 (N_3396,In_1631,In_122);
nor U3397 (N_3397,In_955,In_1572);
and U3398 (N_3398,In_1659,In_911);
or U3399 (N_3399,In_44,In_1935);
and U3400 (N_3400,In_1031,In_584);
nor U3401 (N_3401,In_249,In_1214);
or U3402 (N_3402,In_220,In_1161);
or U3403 (N_3403,In_1268,In_1846);
nand U3404 (N_3404,In_1332,In_1108);
xnor U3405 (N_3405,In_1118,In_503);
nor U3406 (N_3406,In_1923,In_55);
and U3407 (N_3407,In_1757,In_1468);
or U3408 (N_3408,In_345,In_1675);
or U3409 (N_3409,In_1574,In_1484);
or U3410 (N_3410,In_1732,In_966);
nor U3411 (N_3411,In_1789,In_69);
nand U3412 (N_3412,In_852,In_253);
and U3413 (N_3413,In_1857,In_1751);
and U3414 (N_3414,In_673,In_1941);
or U3415 (N_3415,In_1809,In_4);
nand U3416 (N_3416,In_611,In_1793);
or U3417 (N_3417,In_1920,In_1826);
and U3418 (N_3418,In_229,In_626);
nand U3419 (N_3419,In_560,In_934);
and U3420 (N_3420,In_249,In_355);
or U3421 (N_3421,In_562,In_1971);
nor U3422 (N_3422,In_820,In_872);
nand U3423 (N_3423,In_1301,In_157);
and U3424 (N_3424,In_724,In_987);
nand U3425 (N_3425,In_1779,In_1395);
nand U3426 (N_3426,In_871,In_1757);
nand U3427 (N_3427,In_1094,In_1747);
and U3428 (N_3428,In_1342,In_1322);
nor U3429 (N_3429,In_970,In_1380);
nor U3430 (N_3430,In_1557,In_1528);
nor U3431 (N_3431,In_1889,In_339);
nor U3432 (N_3432,In_91,In_1989);
nand U3433 (N_3433,In_433,In_355);
and U3434 (N_3434,In_205,In_497);
nor U3435 (N_3435,In_596,In_1798);
and U3436 (N_3436,In_487,In_327);
nand U3437 (N_3437,In_518,In_1243);
nand U3438 (N_3438,In_1478,In_1287);
nand U3439 (N_3439,In_730,In_640);
and U3440 (N_3440,In_1372,In_501);
nand U3441 (N_3441,In_1074,In_283);
and U3442 (N_3442,In_271,In_41);
nor U3443 (N_3443,In_1556,In_1593);
nand U3444 (N_3444,In_415,In_229);
and U3445 (N_3445,In_566,In_185);
nor U3446 (N_3446,In_544,In_1467);
or U3447 (N_3447,In_1102,In_1860);
xnor U3448 (N_3448,In_310,In_1920);
nor U3449 (N_3449,In_1747,In_1082);
xnor U3450 (N_3450,In_138,In_414);
or U3451 (N_3451,In_1840,In_827);
nor U3452 (N_3452,In_1413,In_1770);
nor U3453 (N_3453,In_209,In_1762);
nor U3454 (N_3454,In_1530,In_43);
or U3455 (N_3455,In_1501,In_230);
nand U3456 (N_3456,In_399,In_1697);
or U3457 (N_3457,In_778,In_937);
nor U3458 (N_3458,In_1545,In_631);
and U3459 (N_3459,In_1805,In_769);
xor U3460 (N_3460,In_1235,In_852);
nand U3461 (N_3461,In_1656,In_796);
and U3462 (N_3462,In_1624,In_666);
xnor U3463 (N_3463,In_1248,In_488);
and U3464 (N_3464,In_1532,In_1202);
and U3465 (N_3465,In_445,In_1808);
and U3466 (N_3466,In_622,In_756);
nor U3467 (N_3467,In_951,In_269);
nor U3468 (N_3468,In_729,In_362);
and U3469 (N_3469,In_402,In_1369);
nand U3470 (N_3470,In_1149,In_645);
nand U3471 (N_3471,In_1275,In_139);
nor U3472 (N_3472,In_1356,In_480);
or U3473 (N_3473,In_1919,In_395);
and U3474 (N_3474,In_1252,In_1214);
or U3475 (N_3475,In_374,In_1203);
xnor U3476 (N_3476,In_558,In_12);
nor U3477 (N_3477,In_1783,In_1911);
and U3478 (N_3478,In_1261,In_141);
and U3479 (N_3479,In_990,In_1728);
nor U3480 (N_3480,In_144,In_1901);
and U3481 (N_3481,In_1987,In_556);
nand U3482 (N_3482,In_1097,In_700);
xnor U3483 (N_3483,In_1145,In_1569);
nor U3484 (N_3484,In_1561,In_1805);
nand U3485 (N_3485,In_1442,In_180);
and U3486 (N_3486,In_256,In_1100);
or U3487 (N_3487,In_240,In_207);
or U3488 (N_3488,In_728,In_623);
nor U3489 (N_3489,In_193,In_484);
xor U3490 (N_3490,In_1180,In_981);
nand U3491 (N_3491,In_1391,In_299);
or U3492 (N_3492,In_408,In_1564);
and U3493 (N_3493,In_559,In_1176);
or U3494 (N_3494,In_898,In_436);
nand U3495 (N_3495,In_974,In_583);
nand U3496 (N_3496,In_1560,In_1284);
nand U3497 (N_3497,In_271,In_1338);
nand U3498 (N_3498,In_1080,In_1391);
or U3499 (N_3499,In_1009,In_1732);
or U3500 (N_3500,In_262,In_455);
or U3501 (N_3501,In_5,In_1828);
nand U3502 (N_3502,In_674,In_1856);
and U3503 (N_3503,In_525,In_439);
xnor U3504 (N_3504,In_1549,In_480);
nand U3505 (N_3505,In_143,In_727);
nand U3506 (N_3506,In_791,In_1837);
nand U3507 (N_3507,In_1459,In_1411);
or U3508 (N_3508,In_163,In_1931);
or U3509 (N_3509,In_1083,In_1899);
nand U3510 (N_3510,In_1758,In_1648);
nor U3511 (N_3511,In_1205,In_1098);
or U3512 (N_3512,In_497,In_1919);
or U3513 (N_3513,In_1759,In_1154);
nand U3514 (N_3514,In_1970,In_220);
nand U3515 (N_3515,In_86,In_1825);
or U3516 (N_3516,In_1762,In_390);
and U3517 (N_3517,In_1243,In_1691);
nand U3518 (N_3518,In_770,In_0);
nor U3519 (N_3519,In_1630,In_422);
xnor U3520 (N_3520,In_1576,In_917);
or U3521 (N_3521,In_565,In_51);
or U3522 (N_3522,In_214,In_98);
nand U3523 (N_3523,In_316,In_1838);
nand U3524 (N_3524,In_492,In_383);
or U3525 (N_3525,In_1234,In_1301);
nand U3526 (N_3526,In_447,In_1242);
and U3527 (N_3527,In_1248,In_1697);
or U3528 (N_3528,In_1408,In_91);
or U3529 (N_3529,In_1157,In_113);
nor U3530 (N_3530,In_1875,In_304);
nand U3531 (N_3531,In_605,In_1488);
nor U3532 (N_3532,In_1711,In_160);
nor U3533 (N_3533,In_877,In_1659);
and U3534 (N_3534,In_1261,In_829);
or U3535 (N_3535,In_569,In_906);
nor U3536 (N_3536,In_129,In_1381);
and U3537 (N_3537,In_527,In_551);
nor U3538 (N_3538,In_195,In_1661);
xor U3539 (N_3539,In_1030,In_915);
nand U3540 (N_3540,In_811,In_1806);
or U3541 (N_3541,In_189,In_1809);
and U3542 (N_3542,In_606,In_1397);
nor U3543 (N_3543,In_1897,In_482);
nand U3544 (N_3544,In_258,In_632);
nor U3545 (N_3545,In_1297,In_1756);
nor U3546 (N_3546,In_1506,In_783);
nor U3547 (N_3547,In_71,In_1135);
and U3548 (N_3548,In_1947,In_1640);
and U3549 (N_3549,In_82,In_1997);
and U3550 (N_3550,In_1620,In_894);
or U3551 (N_3551,In_246,In_1302);
nor U3552 (N_3552,In_1522,In_2);
nand U3553 (N_3553,In_1336,In_1829);
and U3554 (N_3554,In_892,In_1251);
xor U3555 (N_3555,In_1574,In_1673);
xor U3556 (N_3556,In_806,In_1376);
nor U3557 (N_3557,In_179,In_1265);
nor U3558 (N_3558,In_91,In_1480);
and U3559 (N_3559,In_662,In_365);
and U3560 (N_3560,In_685,In_277);
or U3561 (N_3561,In_1296,In_1011);
nor U3562 (N_3562,In_540,In_1501);
nor U3563 (N_3563,In_349,In_798);
or U3564 (N_3564,In_387,In_561);
nor U3565 (N_3565,In_1982,In_588);
nor U3566 (N_3566,In_1072,In_1232);
xnor U3567 (N_3567,In_886,In_149);
nor U3568 (N_3568,In_1439,In_9);
xor U3569 (N_3569,In_905,In_1738);
nand U3570 (N_3570,In_1582,In_500);
or U3571 (N_3571,In_801,In_1452);
xnor U3572 (N_3572,In_1123,In_810);
or U3573 (N_3573,In_1593,In_1235);
nand U3574 (N_3574,In_890,In_1618);
and U3575 (N_3575,In_67,In_1098);
nand U3576 (N_3576,In_1507,In_1965);
xnor U3577 (N_3577,In_63,In_941);
nand U3578 (N_3578,In_365,In_388);
nand U3579 (N_3579,In_1000,In_252);
and U3580 (N_3580,In_1714,In_470);
nand U3581 (N_3581,In_1353,In_1825);
and U3582 (N_3582,In_643,In_1869);
or U3583 (N_3583,In_864,In_1311);
nand U3584 (N_3584,In_68,In_1301);
or U3585 (N_3585,In_41,In_1324);
or U3586 (N_3586,In_993,In_1928);
and U3587 (N_3587,In_1599,In_1990);
and U3588 (N_3588,In_1043,In_170);
nor U3589 (N_3589,In_1217,In_1370);
or U3590 (N_3590,In_481,In_1314);
or U3591 (N_3591,In_1140,In_649);
and U3592 (N_3592,In_1377,In_679);
nor U3593 (N_3593,In_1184,In_828);
nor U3594 (N_3594,In_847,In_235);
nand U3595 (N_3595,In_219,In_66);
or U3596 (N_3596,In_1241,In_916);
xnor U3597 (N_3597,In_1496,In_1115);
nand U3598 (N_3598,In_391,In_988);
nand U3599 (N_3599,In_550,In_1300);
and U3600 (N_3600,In_1199,In_1367);
nand U3601 (N_3601,In_1664,In_1813);
or U3602 (N_3602,In_1574,In_1811);
or U3603 (N_3603,In_318,In_511);
nor U3604 (N_3604,In_698,In_1853);
and U3605 (N_3605,In_1442,In_1968);
xor U3606 (N_3606,In_539,In_165);
xor U3607 (N_3607,In_1286,In_434);
nor U3608 (N_3608,In_1058,In_796);
xnor U3609 (N_3609,In_768,In_1521);
and U3610 (N_3610,In_504,In_1155);
and U3611 (N_3611,In_159,In_1162);
nand U3612 (N_3612,In_1096,In_1112);
and U3613 (N_3613,In_889,In_290);
or U3614 (N_3614,In_422,In_403);
nand U3615 (N_3615,In_1624,In_1328);
nor U3616 (N_3616,In_196,In_621);
and U3617 (N_3617,In_1892,In_1174);
or U3618 (N_3618,In_1244,In_1233);
and U3619 (N_3619,In_408,In_1641);
and U3620 (N_3620,In_1148,In_320);
and U3621 (N_3621,In_1499,In_229);
nand U3622 (N_3622,In_197,In_516);
xnor U3623 (N_3623,In_1070,In_1981);
nor U3624 (N_3624,In_834,In_1272);
nand U3625 (N_3625,In_1922,In_1373);
nor U3626 (N_3626,In_276,In_1978);
nor U3627 (N_3627,In_1400,In_1615);
or U3628 (N_3628,In_995,In_903);
or U3629 (N_3629,In_1086,In_1628);
and U3630 (N_3630,In_503,In_1810);
nand U3631 (N_3631,In_1845,In_1662);
nor U3632 (N_3632,In_252,In_798);
nor U3633 (N_3633,In_984,In_1868);
xnor U3634 (N_3634,In_385,In_113);
or U3635 (N_3635,In_178,In_1912);
and U3636 (N_3636,In_1361,In_1362);
nor U3637 (N_3637,In_35,In_1391);
nand U3638 (N_3638,In_1098,In_174);
nand U3639 (N_3639,In_440,In_964);
and U3640 (N_3640,In_587,In_1256);
and U3641 (N_3641,In_1737,In_306);
xnor U3642 (N_3642,In_1750,In_837);
or U3643 (N_3643,In_424,In_1355);
nor U3644 (N_3644,In_5,In_1950);
and U3645 (N_3645,In_1477,In_1944);
nand U3646 (N_3646,In_477,In_1015);
nand U3647 (N_3647,In_1529,In_1893);
nor U3648 (N_3648,In_1102,In_198);
nor U3649 (N_3649,In_833,In_636);
or U3650 (N_3650,In_1448,In_877);
and U3651 (N_3651,In_758,In_677);
nand U3652 (N_3652,In_1399,In_1644);
nor U3653 (N_3653,In_1844,In_773);
nor U3654 (N_3654,In_207,In_252);
or U3655 (N_3655,In_1806,In_426);
and U3656 (N_3656,In_1334,In_1878);
nor U3657 (N_3657,In_1610,In_822);
nand U3658 (N_3658,In_371,In_1821);
nand U3659 (N_3659,In_647,In_859);
nor U3660 (N_3660,In_500,In_100);
and U3661 (N_3661,In_55,In_626);
nand U3662 (N_3662,In_920,In_1100);
or U3663 (N_3663,In_660,In_64);
xnor U3664 (N_3664,In_1905,In_1144);
or U3665 (N_3665,In_734,In_1767);
nand U3666 (N_3666,In_326,In_1724);
nor U3667 (N_3667,In_1054,In_1443);
nand U3668 (N_3668,In_720,In_604);
or U3669 (N_3669,In_344,In_632);
and U3670 (N_3670,In_451,In_1828);
nor U3671 (N_3671,In_559,In_226);
or U3672 (N_3672,In_579,In_1844);
nor U3673 (N_3673,In_1172,In_241);
or U3674 (N_3674,In_23,In_1714);
xnor U3675 (N_3675,In_1978,In_1944);
nor U3676 (N_3676,In_1214,In_1320);
nand U3677 (N_3677,In_261,In_1219);
and U3678 (N_3678,In_615,In_455);
nor U3679 (N_3679,In_1463,In_645);
and U3680 (N_3680,In_353,In_1521);
and U3681 (N_3681,In_548,In_1796);
and U3682 (N_3682,In_1798,In_1494);
nand U3683 (N_3683,In_1661,In_199);
or U3684 (N_3684,In_215,In_160);
nand U3685 (N_3685,In_1841,In_1174);
or U3686 (N_3686,In_1527,In_495);
nand U3687 (N_3687,In_1585,In_1774);
nand U3688 (N_3688,In_1944,In_806);
nor U3689 (N_3689,In_433,In_1362);
or U3690 (N_3690,In_145,In_1455);
or U3691 (N_3691,In_1337,In_1480);
nor U3692 (N_3692,In_1151,In_848);
nor U3693 (N_3693,In_1795,In_1140);
and U3694 (N_3694,In_1502,In_1453);
nand U3695 (N_3695,In_388,In_448);
and U3696 (N_3696,In_1317,In_998);
and U3697 (N_3697,In_1788,In_923);
and U3698 (N_3698,In_1624,In_1286);
and U3699 (N_3699,In_388,In_1687);
nand U3700 (N_3700,In_1998,In_1712);
and U3701 (N_3701,In_723,In_1915);
or U3702 (N_3702,In_484,In_892);
and U3703 (N_3703,In_1732,In_1752);
or U3704 (N_3704,In_1269,In_865);
nor U3705 (N_3705,In_1545,In_755);
or U3706 (N_3706,In_938,In_1120);
nor U3707 (N_3707,In_1466,In_1251);
xnor U3708 (N_3708,In_49,In_1052);
xor U3709 (N_3709,In_792,In_885);
nand U3710 (N_3710,In_342,In_600);
and U3711 (N_3711,In_1350,In_1407);
nor U3712 (N_3712,In_667,In_411);
xor U3713 (N_3713,In_976,In_1060);
or U3714 (N_3714,In_1121,In_1779);
xor U3715 (N_3715,In_980,In_974);
nor U3716 (N_3716,In_1846,In_1358);
nor U3717 (N_3717,In_1753,In_1161);
or U3718 (N_3718,In_208,In_1078);
xor U3719 (N_3719,In_331,In_986);
nand U3720 (N_3720,In_1100,In_1935);
nor U3721 (N_3721,In_238,In_1584);
or U3722 (N_3722,In_1946,In_1100);
xor U3723 (N_3723,In_375,In_1636);
nand U3724 (N_3724,In_1785,In_39);
or U3725 (N_3725,In_1219,In_380);
nand U3726 (N_3726,In_465,In_1086);
nand U3727 (N_3727,In_406,In_346);
or U3728 (N_3728,In_966,In_489);
or U3729 (N_3729,In_1825,In_376);
or U3730 (N_3730,In_593,In_599);
or U3731 (N_3731,In_1955,In_715);
and U3732 (N_3732,In_654,In_1635);
nor U3733 (N_3733,In_1871,In_588);
and U3734 (N_3734,In_181,In_1254);
nand U3735 (N_3735,In_1382,In_1815);
and U3736 (N_3736,In_154,In_1956);
xor U3737 (N_3737,In_1566,In_1869);
or U3738 (N_3738,In_1796,In_215);
nand U3739 (N_3739,In_201,In_84);
xnor U3740 (N_3740,In_1787,In_712);
and U3741 (N_3741,In_1616,In_1459);
nor U3742 (N_3742,In_191,In_632);
nand U3743 (N_3743,In_1535,In_1478);
and U3744 (N_3744,In_617,In_1448);
xnor U3745 (N_3745,In_796,In_874);
nand U3746 (N_3746,In_299,In_491);
and U3747 (N_3747,In_582,In_656);
nor U3748 (N_3748,In_621,In_1629);
or U3749 (N_3749,In_787,In_1908);
xor U3750 (N_3750,In_1094,In_288);
and U3751 (N_3751,In_1766,In_978);
or U3752 (N_3752,In_83,In_561);
nand U3753 (N_3753,In_801,In_1883);
and U3754 (N_3754,In_709,In_416);
and U3755 (N_3755,In_1506,In_1153);
xor U3756 (N_3756,In_740,In_427);
or U3757 (N_3757,In_1097,In_1516);
nand U3758 (N_3758,In_398,In_223);
and U3759 (N_3759,In_259,In_1856);
and U3760 (N_3760,In_1788,In_1071);
or U3761 (N_3761,In_1555,In_674);
xnor U3762 (N_3762,In_621,In_387);
nand U3763 (N_3763,In_1439,In_1585);
or U3764 (N_3764,In_733,In_1586);
nor U3765 (N_3765,In_501,In_1719);
and U3766 (N_3766,In_510,In_562);
nand U3767 (N_3767,In_1944,In_621);
or U3768 (N_3768,In_1969,In_757);
nand U3769 (N_3769,In_103,In_1522);
and U3770 (N_3770,In_1663,In_290);
nor U3771 (N_3771,In_1787,In_261);
nand U3772 (N_3772,In_1890,In_1545);
nor U3773 (N_3773,In_936,In_722);
nand U3774 (N_3774,In_763,In_1274);
nand U3775 (N_3775,In_923,In_1171);
nor U3776 (N_3776,In_1983,In_406);
or U3777 (N_3777,In_789,In_641);
or U3778 (N_3778,In_632,In_1929);
nor U3779 (N_3779,In_567,In_1338);
nand U3780 (N_3780,In_312,In_97);
nor U3781 (N_3781,In_1280,In_1320);
nand U3782 (N_3782,In_356,In_165);
nor U3783 (N_3783,In_1859,In_1766);
and U3784 (N_3784,In_1169,In_1145);
nor U3785 (N_3785,In_1499,In_710);
nand U3786 (N_3786,In_874,In_713);
or U3787 (N_3787,In_990,In_14);
xnor U3788 (N_3788,In_1116,In_1534);
and U3789 (N_3789,In_274,In_154);
and U3790 (N_3790,In_679,In_934);
nand U3791 (N_3791,In_862,In_265);
nor U3792 (N_3792,In_476,In_189);
and U3793 (N_3793,In_1347,In_1465);
or U3794 (N_3794,In_969,In_1664);
nand U3795 (N_3795,In_1029,In_937);
or U3796 (N_3796,In_1864,In_1469);
nand U3797 (N_3797,In_989,In_391);
or U3798 (N_3798,In_922,In_634);
nor U3799 (N_3799,In_1449,In_1438);
nand U3800 (N_3800,In_644,In_1284);
nor U3801 (N_3801,In_943,In_948);
or U3802 (N_3802,In_1785,In_634);
or U3803 (N_3803,In_138,In_726);
nor U3804 (N_3804,In_260,In_1965);
nand U3805 (N_3805,In_1635,In_1993);
and U3806 (N_3806,In_635,In_43);
xnor U3807 (N_3807,In_1241,In_1195);
nor U3808 (N_3808,In_4,In_538);
nor U3809 (N_3809,In_988,In_932);
nand U3810 (N_3810,In_153,In_1412);
or U3811 (N_3811,In_812,In_1918);
or U3812 (N_3812,In_1344,In_1448);
or U3813 (N_3813,In_531,In_244);
and U3814 (N_3814,In_1780,In_635);
nor U3815 (N_3815,In_118,In_1660);
and U3816 (N_3816,In_994,In_728);
and U3817 (N_3817,In_764,In_713);
or U3818 (N_3818,In_1740,In_984);
xor U3819 (N_3819,In_1008,In_1430);
and U3820 (N_3820,In_783,In_449);
or U3821 (N_3821,In_1817,In_189);
and U3822 (N_3822,In_1417,In_1080);
and U3823 (N_3823,In_1833,In_1846);
nand U3824 (N_3824,In_321,In_1601);
or U3825 (N_3825,In_1728,In_1757);
nand U3826 (N_3826,In_590,In_856);
nand U3827 (N_3827,In_829,In_1006);
and U3828 (N_3828,In_1963,In_505);
nor U3829 (N_3829,In_1636,In_53);
or U3830 (N_3830,In_818,In_1167);
and U3831 (N_3831,In_1010,In_40);
nand U3832 (N_3832,In_514,In_1660);
nand U3833 (N_3833,In_1653,In_95);
and U3834 (N_3834,In_187,In_1762);
or U3835 (N_3835,In_365,In_42);
or U3836 (N_3836,In_123,In_417);
nor U3837 (N_3837,In_1879,In_1687);
nor U3838 (N_3838,In_598,In_645);
nand U3839 (N_3839,In_1286,In_989);
or U3840 (N_3840,In_327,In_765);
nor U3841 (N_3841,In_646,In_546);
and U3842 (N_3842,In_1608,In_159);
and U3843 (N_3843,In_1941,In_613);
nand U3844 (N_3844,In_434,In_1916);
xnor U3845 (N_3845,In_746,In_315);
nand U3846 (N_3846,In_519,In_1967);
nor U3847 (N_3847,In_919,In_707);
nor U3848 (N_3848,In_439,In_124);
nand U3849 (N_3849,In_864,In_1636);
xnor U3850 (N_3850,In_1111,In_93);
or U3851 (N_3851,In_307,In_1608);
nand U3852 (N_3852,In_917,In_1428);
or U3853 (N_3853,In_1254,In_162);
nand U3854 (N_3854,In_883,In_765);
xnor U3855 (N_3855,In_959,In_1240);
or U3856 (N_3856,In_109,In_768);
nor U3857 (N_3857,In_1056,In_1943);
xnor U3858 (N_3858,In_1594,In_448);
xnor U3859 (N_3859,In_785,In_1543);
or U3860 (N_3860,In_1782,In_434);
nor U3861 (N_3861,In_1651,In_1491);
and U3862 (N_3862,In_758,In_1056);
nand U3863 (N_3863,In_1735,In_1424);
and U3864 (N_3864,In_187,In_1774);
nand U3865 (N_3865,In_731,In_1306);
nor U3866 (N_3866,In_308,In_460);
and U3867 (N_3867,In_507,In_1455);
nor U3868 (N_3868,In_337,In_620);
nand U3869 (N_3869,In_1360,In_1656);
or U3870 (N_3870,In_87,In_374);
or U3871 (N_3871,In_1115,In_1425);
or U3872 (N_3872,In_260,In_466);
or U3873 (N_3873,In_471,In_1946);
nand U3874 (N_3874,In_1519,In_999);
nor U3875 (N_3875,In_1590,In_1697);
nor U3876 (N_3876,In_78,In_1206);
nand U3877 (N_3877,In_729,In_1104);
nand U3878 (N_3878,In_1968,In_1753);
nor U3879 (N_3879,In_95,In_765);
nand U3880 (N_3880,In_1112,In_716);
nand U3881 (N_3881,In_167,In_537);
or U3882 (N_3882,In_1411,In_461);
xnor U3883 (N_3883,In_1510,In_1406);
nor U3884 (N_3884,In_979,In_1573);
and U3885 (N_3885,In_842,In_37);
nor U3886 (N_3886,In_898,In_538);
nor U3887 (N_3887,In_241,In_1340);
nand U3888 (N_3888,In_1592,In_1637);
nor U3889 (N_3889,In_461,In_216);
nand U3890 (N_3890,In_1740,In_822);
and U3891 (N_3891,In_56,In_581);
nor U3892 (N_3892,In_1291,In_150);
or U3893 (N_3893,In_1263,In_1061);
or U3894 (N_3894,In_1638,In_21);
or U3895 (N_3895,In_172,In_896);
and U3896 (N_3896,In_401,In_1041);
nand U3897 (N_3897,In_1050,In_1420);
nand U3898 (N_3898,In_99,In_1460);
nor U3899 (N_3899,In_635,In_800);
nor U3900 (N_3900,In_1039,In_426);
nor U3901 (N_3901,In_944,In_799);
and U3902 (N_3902,In_1392,In_1561);
nor U3903 (N_3903,In_200,In_395);
or U3904 (N_3904,In_1174,In_624);
and U3905 (N_3905,In_1707,In_591);
or U3906 (N_3906,In_487,In_1547);
nand U3907 (N_3907,In_1632,In_1081);
and U3908 (N_3908,In_352,In_636);
nand U3909 (N_3909,In_785,In_1318);
nor U3910 (N_3910,In_101,In_894);
or U3911 (N_3911,In_41,In_669);
xor U3912 (N_3912,In_1299,In_1053);
xnor U3913 (N_3913,In_700,In_502);
nor U3914 (N_3914,In_1055,In_82);
xor U3915 (N_3915,In_695,In_1399);
and U3916 (N_3916,In_1834,In_539);
or U3917 (N_3917,In_1541,In_421);
nor U3918 (N_3918,In_128,In_346);
or U3919 (N_3919,In_142,In_596);
and U3920 (N_3920,In_1302,In_669);
nand U3921 (N_3921,In_1647,In_1408);
and U3922 (N_3922,In_427,In_688);
or U3923 (N_3923,In_399,In_1298);
or U3924 (N_3924,In_185,In_803);
nand U3925 (N_3925,In_1087,In_989);
or U3926 (N_3926,In_1770,In_321);
and U3927 (N_3927,In_643,In_1514);
and U3928 (N_3928,In_768,In_1273);
or U3929 (N_3929,In_1934,In_1713);
nor U3930 (N_3930,In_1902,In_1969);
nor U3931 (N_3931,In_1796,In_1637);
nand U3932 (N_3932,In_1420,In_944);
or U3933 (N_3933,In_1469,In_1274);
and U3934 (N_3934,In_1307,In_244);
and U3935 (N_3935,In_1017,In_1384);
nand U3936 (N_3936,In_1921,In_68);
or U3937 (N_3937,In_1673,In_1291);
xor U3938 (N_3938,In_648,In_110);
or U3939 (N_3939,In_1302,In_1138);
or U3940 (N_3940,In_1269,In_34);
nand U3941 (N_3941,In_445,In_264);
and U3942 (N_3942,In_604,In_976);
nand U3943 (N_3943,In_343,In_36);
nor U3944 (N_3944,In_173,In_634);
or U3945 (N_3945,In_102,In_1072);
or U3946 (N_3946,In_1259,In_1069);
nor U3947 (N_3947,In_422,In_964);
nand U3948 (N_3948,In_831,In_1682);
nor U3949 (N_3949,In_1033,In_1221);
nand U3950 (N_3950,In_759,In_1134);
and U3951 (N_3951,In_1617,In_1727);
nor U3952 (N_3952,In_146,In_72);
nand U3953 (N_3953,In_561,In_1833);
xor U3954 (N_3954,In_1823,In_985);
or U3955 (N_3955,In_1287,In_1309);
and U3956 (N_3956,In_1244,In_1062);
xnor U3957 (N_3957,In_910,In_277);
or U3958 (N_3958,In_453,In_663);
and U3959 (N_3959,In_985,In_667);
and U3960 (N_3960,In_1429,In_328);
and U3961 (N_3961,In_172,In_491);
and U3962 (N_3962,In_1662,In_580);
nor U3963 (N_3963,In_52,In_80);
nor U3964 (N_3964,In_309,In_630);
xor U3965 (N_3965,In_627,In_821);
or U3966 (N_3966,In_789,In_751);
nand U3967 (N_3967,In_1590,In_1181);
and U3968 (N_3968,In_1315,In_61);
and U3969 (N_3969,In_540,In_1077);
or U3970 (N_3970,In_272,In_1920);
nor U3971 (N_3971,In_1859,In_1120);
nor U3972 (N_3972,In_208,In_581);
or U3973 (N_3973,In_925,In_1121);
and U3974 (N_3974,In_598,In_1164);
xor U3975 (N_3975,In_581,In_1530);
nor U3976 (N_3976,In_535,In_1464);
nand U3977 (N_3977,In_1399,In_1880);
nor U3978 (N_3978,In_970,In_1187);
nand U3979 (N_3979,In_253,In_1621);
nand U3980 (N_3980,In_522,In_555);
nor U3981 (N_3981,In_1530,In_1495);
and U3982 (N_3982,In_1521,In_447);
nand U3983 (N_3983,In_1462,In_342);
and U3984 (N_3984,In_546,In_1387);
nand U3985 (N_3985,In_1464,In_1056);
and U3986 (N_3986,In_1605,In_908);
or U3987 (N_3987,In_1337,In_17);
nand U3988 (N_3988,In_1129,In_615);
and U3989 (N_3989,In_563,In_1211);
nor U3990 (N_3990,In_102,In_760);
and U3991 (N_3991,In_1813,In_269);
nand U3992 (N_3992,In_1289,In_158);
nor U3993 (N_3993,In_1474,In_1886);
or U3994 (N_3994,In_56,In_1719);
nand U3995 (N_3995,In_1811,In_1718);
nor U3996 (N_3996,In_1054,In_1039);
nand U3997 (N_3997,In_1904,In_1496);
nor U3998 (N_3998,In_265,In_1982);
nand U3999 (N_3999,In_987,In_840);
nand U4000 (N_4000,N_3849,N_3621);
or U4001 (N_4001,N_1678,N_1742);
nor U4002 (N_4002,N_3764,N_3600);
nand U4003 (N_4003,N_316,N_3826);
nand U4004 (N_4004,N_1839,N_3444);
xnor U4005 (N_4005,N_122,N_2847);
and U4006 (N_4006,N_1295,N_739);
nor U4007 (N_4007,N_1621,N_3098);
nor U4008 (N_4008,N_1233,N_250);
and U4009 (N_4009,N_3582,N_2247);
or U4010 (N_4010,N_2448,N_3180);
and U4011 (N_4011,N_2100,N_931);
or U4012 (N_4012,N_1904,N_2580);
and U4013 (N_4013,N_873,N_804);
xnor U4014 (N_4014,N_3193,N_1712);
nor U4015 (N_4015,N_3378,N_2432);
nor U4016 (N_4016,N_3191,N_726);
or U4017 (N_4017,N_447,N_2749);
and U4018 (N_4018,N_415,N_1326);
nand U4019 (N_4019,N_1642,N_3711);
and U4020 (N_4020,N_3596,N_3768);
nand U4021 (N_4021,N_2829,N_2615);
nand U4022 (N_4022,N_233,N_3588);
and U4023 (N_4023,N_3623,N_685);
nor U4024 (N_4024,N_745,N_1408);
nand U4025 (N_4025,N_575,N_3151);
nand U4026 (N_4026,N_1555,N_2519);
xnor U4027 (N_4027,N_290,N_917);
and U4028 (N_4028,N_2628,N_3552);
nor U4029 (N_4029,N_3274,N_2154);
nand U4030 (N_4030,N_2608,N_178);
and U4031 (N_4031,N_2697,N_2449);
and U4032 (N_4032,N_2709,N_3377);
or U4033 (N_4033,N_1434,N_1545);
nor U4034 (N_4034,N_1231,N_1360);
or U4035 (N_4035,N_2277,N_835);
or U4036 (N_4036,N_3092,N_274);
xor U4037 (N_4037,N_2031,N_3078);
nor U4038 (N_4038,N_2024,N_1673);
nor U4039 (N_4039,N_2422,N_1818);
or U4040 (N_4040,N_1021,N_1467);
and U4041 (N_4041,N_3341,N_433);
and U4042 (N_4042,N_3519,N_1169);
xnor U4043 (N_4043,N_2579,N_3490);
nor U4044 (N_4044,N_3023,N_3941);
and U4045 (N_4045,N_949,N_487);
nor U4046 (N_4046,N_3505,N_819);
or U4047 (N_4047,N_1575,N_136);
or U4048 (N_4048,N_3494,N_1289);
or U4049 (N_4049,N_3999,N_1596);
nand U4050 (N_4050,N_573,N_3113);
nor U4051 (N_4051,N_544,N_183);
nor U4052 (N_4052,N_2332,N_1628);
xor U4053 (N_4053,N_1574,N_891);
nor U4054 (N_4054,N_2503,N_2101);
nand U4055 (N_4055,N_1014,N_77);
nor U4056 (N_4056,N_3889,N_3610);
and U4057 (N_4057,N_2178,N_3190);
and U4058 (N_4058,N_3453,N_904);
xor U4059 (N_4059,N_3607,N_1722);
nor U4060 (N_4060,N_1861,N_2092);
or U4061 (N_4061,N_3026,N_2284);
xnor U4062 (N_4062,N_128,N_2870);
and U4063 (N_4063,N_650,N_3844);
nand U4064 (N_4064,N_1209,N_2496);
or U4065 (N_4065,N_1862,N_3467);
or U4066 (N_4066,N_1812,N_2581);
or U4067 (N_4067,N_1849,N_3192);
or U4068 (N_4068,N_3967,N_1114);
and U4069 (N_4069,N_3995,N_2116);
and U4070 (N_4070,N_1824,N_3181);
nor U4071 (N_4071,N_2714,N_2254);
xor U4072 (N_4072,N_1670,N_1653);
and U4073 (N_4073,N_2766,N_3627);
nor U4074 (N_4074,N_1842,N_2688);
nor U4075 (N_4075,N_3514,N_3038);
xor U4076 (N_4076,N_74,N_2785);
xnor U4077 (N_4077,N_3950,N_2699);
or U4078 (N_4078,N_571,N_3501);
nor U4079 (N_4079,N_1676,N_2691);
and U4080 (N_4080,N_764,N_3470);
nor U4081 (N_4081,N_2602,N_2864);
nor U4082 (N_4082,N_1539,N_354);
nand U4083 (N_4083,N_1112,N_1896);
and U4084 (N_4084,N_1763,N_2658);
or U4085 (N_4085,N_2755,N_847);
xor U4086 (N_4086,N_3899,N_2427);
xnor U4087 (N_4087,N_1113,N_1310);
nor U4088 (N_4088,N_2337,N_349);
or U4089 (N_4089,N_2372,N_645);
nand U4090 (N_4090,N_1221,N_1605);
or U4091 (N_4091,N_2931,N_768);
nand U4092 (N_4092,N_2086,N_1106);
nor U4093 (N_4093,N_563,N_2975);
nor U4094 (N_4094,N_3635,N_2486);
xnor U4095 (N_4095,N_3604,N_699);
nand U4096 (N_4096,N_1695,N_386);
or U4097 (N_4097,N_2308,N_2052);
nor U4098 (N_4098,N_476,N_1174);
nand U4099 (N_4099,N_2523,N_3441);
and U4100 (N_4100,N_1424,N_159);
nor U4101 (N_4101,N_698,N_2919);
nand U4102 (N_4102,N_149,N_3808);
nor U4103 (N_4103,N_1941,N_3553);
or U4104 (N_4104,N_3175,N_515);
nand U4105 (N_4105,N_630,N_1521);
or U4106 (N_4106,N_1238,N_3935);
nand U4107 (N_4107,N_121,N_1751);
nand U4108 (N_4108,N_384,N_3442);
nor U4109 (N_4109,N_1547,N_1980);
nor U4110 (N_4110,N_1368,N_1131);
and U4111 (N_4111,N_2767,N_559);
nand U4112 (N_4112,N_695,N_3060);
xor U4113 (N_4113,N_3801,N_2787);
nand U4114 (N_4114,N_1503,N_2941);
nor U4115 (N_4115,N_1156,N_3154);
nand U4116 (N_4116,N_3919,N_662);
nand U4117 (N_4117,N_1070,N_1506);
and U4118 (N_4118,N_1510,N_2543);
nor U4119 (N_4119,N_1256,N_1648);
nor U4120 (N_4120,N_3250,N_2992);
or U4121 (N_4121,N_2409,N_3882);
nand U4122 (N_4122,N_689,N_3533);
nor U4123 (N_4123,N_2853,N_1500);
or U4124 (N_4124,N_2062,N_402);
or U4125 (N_4125,N_3946,N_2330);
or U4126 (N_4126,N_2637,N_3408);
and U4127 (N_4127,N_3286,N_356);
and U4128 (N_4128,N_1723,N_3759);
nor U4129 (N_4129,N_3160,N_3485);
and U4130 (N_4130,N_2612,N_2158);
and U4131 (N_4131,N_692,N_694);
nand U4132 (N_4132,N_2609,N_378);
nor U4133 (N_4133,N_2266,N_269);
nand U4134 (N_4134,N_738,N_3318);
or U4135 (N_4135,N_852,N_1755);
or U4136 (N_4136,N_185,N_3856);
xnor U4137 (N_4137,N_2732,N_1453);
xor U4138 (N_4138,N_3474,N_814);
or U4139 (N_4139,N_2573,N_2544);
nor U4140 (N_4140,N_3987,N_581);
nor U4141 (N_4141,N_2892,N_1475);
or U4142 (N_4142,N_3997,N_3932);
nor U4143 (N_4143,N_1840,N_1227);
nor U4144 (N_4144,N_382,N_2899);
or U4145 (N_4145,N_1171,N_3232);
nand U4146 (N_4146,N_3165,N_3710);
nand U4147 (N_4147,N_3345,N_1418);
nor U4148 (N_4148,N_421,N_3930);
nand U4149 (N_4149,N_1721,N_3030);
and U4150 (N_4150,N_3806,N_3022);
xor U4151 (N_4151,N_2272,N_3745);
nor U4152 (N_4152,N_305,N_1054);
or U4153 (N_4153,N_1945,N_2420);
or U4154 (N_4154,N_989,N_2090);
nand U4155 (N_4155,N_1313,N_3169);
nor U4156 (N_4156,N_3230,N_230);
nand U4157 (N_4157,N_3668,N_2061);
nor U4158 (N_4158,N_1271,N_211);
nand U4159 (N_4159,N_2351,N_1650);
nor U4160 (N_4160,N_1457,N_913);
nand U4161 (N_4161,N_686,N_1656);
xnor U4162 (N_4162,N_282,N_2171);
nor U4163 (N_4163,N_350,N_625);
and U4164 (N_4164,N_3460,N_2526);
nor U4165 (N_4165,N_3829,N_3951);
xnor U4166 (N_4166,N_1397,N_3456);
and U4167 (N_4167,N_2151,N_900);
and U4168 (N_4168,N_984,N_1699);
nor U4169 (N_4169,N_1957,N_1924);
and U4170 (N_4170,N_2226,N_756);
or U4171 (N_4171,N_3753,N_2190);
or U4172 (N_4172,N_787,N_3497);
xor U4173 (N_4173,N_3721,N_1761);
nor U4174 (N_4174,N_1459,N_1556);
and U4175 (N_4175,N_2321,N_3222);
and U4176 (N_4176,N_1180,N_1191);
or U4177 (N_4177,N_2704,N_1549);
or U4178 (N_4178,N_2618,N_2730);
or U4179 (N_4179,N_147,N_1659);
and U4180 (N_4180,N_219,N_3001);
xor U4181 (N_4181,N_890,N_658);
or U4182 (N_4182,N_3472,N_3793);
nor U4183 (N_4183,N_295,N_2912);
nand U4184 (N_4184,N_3320,N_3924);
and U4185 (N_4185,N_1009,N_2459);
xnor U4186 (N_4186,N_3097,N_718);
xnor U4187 (N_4187,N_3064,N_657);
nand U4188 (N_4188,N_868,N_2323);
xnor U4189 (N_4189,N_864,N_1585);
and U4190 (N_4190,N_3564,N_2072);
or U4191 (N_4191,N_1303,N_1955);
or U4192 (N_4192,N_376,N_3658);
nand U4193 (N_4193,N_1882,N_1765);
and U4194 (N_4194,N_3788,N_3067);
or U4195 (N_4195,N_1305,N_2130);
or U4196 (N_4196,N_951,N_2725);
nor U4197 (N_4197,N_1858,N_2595);
nor U4198 (N_4198,N_73,N_3928);
and U4199 (N_4199,N_895,N_3700);
and U4200 (N_4200,N_1463,N_3381);
and U4201 (N_4201,N_1655,N_1287);
nand U4202 (N_4202,N_458,N_1683);
nand U4203 (N_4203,N_823,N_2124);
nand U4204 (N_4204,N_1377,N_1876);
nand U4205 (N_4205,N_3331,N_1996);
and U4206 (N_4206,N_3295,N_1728);
or U4207 (N_4207,N_3210,N_1880);
and U4208 (N_4208,N_4,N_2669);
nand U4209 (N_4209,N_3150,N_3188);
nor U4210 (N_4210,N_3428,N_2363);
or U4211 (N_4211,N_102,N_80);
nor U4212 (N_4212,N_906,N_3651);
nand U4213 (N_4213,N_65,N_970);
nand U4214 (N_4214,N_1123,N_398);
nor U4215 (N_4215,N_908,N_2307);
nand U4216 (N_4216,N_1454,N_1879);
or U4217 (N_4217,N_5,N_2832);
nand U4218 (N_4218,N_2001,N_1580);
and U4219 (N_4219,N_2378,N_505);
xnor U4220 (N_4220,N_2642,N_3732);
or U4221 (N_4221,N_2937,N_2487);
nor U4222 (N_4222,N_1081,N_27);
or U4223 (N_4223,N_2902,N_1373);
nand U4224 (N_4224,N_2067,N_2930);
nand U4225 (N_4225,N_3090,N_38);
nand U4226 (N_4226,N_1601,N_1778);
and U4227 (N_4227,N_3525,N_3775);
or U4228 (N_4228,N_1914,N_2655);
xnor U4229 (N_4229,N_1176,N_1530);
or U4230 (N_4230,N_3041,N_60);
nor U4231 (N_4231,N_1793,N_1959);
and U4232 (N_4232,N_574,N_772);
nor U4233 (N_4233,N_1967,N_2071);
or U4234 (N_4234,N_1348,N_3632);
nand U4235 (N_4235,N_3595,N_1988);
nand U4236 (N_4236,N_3702,N_140);
nand U4237 (N_4237,N_1323,N_2451);
or U4238 (N_4238,N_2694,N_1590);
and U4239 (N_4239,N_1175,N_1711);
and U4240 (N_4240,N_3128,N_2080);
or U4241 (N_4241,N_262,N_1860);
or U4242 (N_4242,N_2860,N_1265);
and U4243 (N_4243,N_3224,N_3937);
nor U4244 (N_4244,N_547,N_198);
nor U4245 (N_4245,N_1104,N_380);
nor U4246 (N_4246,N_3529,N_2053);
and U4247 (N_4247,N_2365,N_508);
nor U4248 (N_4248,N_2150,N_1432);
nor U4249 (N_4249,N_3068,N_2993);
or U4250 (N_4250,N_3599,N_855);
nor U4251 (N_4251,N_3332,N_3736);
or U4252 (N_4252,N_1207,N_2155);
nor U4253 (N_4253,N_3061,N_1269);
nand U4254 (N_4254,N_3449,N_3750);
nor U4255 (N_4255,N_1963,N_2495);
and U4256 (N_4256,N_2267,N_2157);
nand U4257 (N_4257,N_953,N_1756);
nand U4258 (N_4258,N_3316,N_3409);
or U4259 (N_4259,N_1272,N_176);
and U4260 (N_4260,N_3045,N_1312);
nor U4261 (N_4261,N_3847,N_760);
nand U4262 (N_4262,N_2692,N_2461);
or U4263 (N_4263,N_1263,N_462);
or U4264 (N_4264,N_3290,N_3130);
nor U4265 (N_4265,N_2835,N_1629);
nand U4266 (N_4266,N_606,N_1046);
and U4267 (N_4267,N_3258,N_3585);
or U4268 (N_4268,N_860,N_1056);
nor U4269 (N_4269,N_1552,N_213);
nor U4270 (N_4270,N_2933,N_2903);
nand U4271 (N_4271,N_319,N_3382);
nor U4272 (N_4272,N_3254,N_100);
and U4273 (N_4273,N_2474,N_1713);
nand U4274 (N_4274,N_2536,N_2672);
xor U4275 (N_4275,N_2118,N_1570);
nand U4276 (N_4276,N_138,N_1551);
nand U4277 (N_4277,N_2586,N_2837);
or U4278 (N_4278,N_1359,N_330);
nand U4279 (N_4279,N_3571,N_1385);
and U4280 (N_4280,N_287,N_598);
or U4281 (N_4281,N_2574,N_2589);
nand U4282 (N_4282,N_388,N_961);
or U4283 (N_4283,N_3065,N_733);
nand U4284 (N_4284,N_3147,N_1871);
or U4285 (N_4285,N_767,N_2188);
nor U4286 (N_4286,N_212,N_569);
or U4287 (N_4287,N_2865,N_786);
nand U4288 (N_4288,N_2007,N_3731);
nand U4289 (N_4289,N_968,N_2850);
nand U4290 (N_4290,N_3390,N_96);
and U4291 (N_4291,N_1498,N_3686);
nor U4292 (N_4292,N_2388,N_2973);
and U4293 (N_4293,N_460,N_3953);
and U4294 (N_4294,N_1685,N_1883);
xnor U4295 (N_4295,N_2738,N_2506);
and U4296 (N_4296,N_1679,N_1304);
and U4297 (N_4297,N_3330,N_3207);
or U4298 (N_4298,N_493,N_729);
xnor U4299 (N_4299,N_1491,N_706);
nor U4300 (N_4300,N_1384,N_1768);
nor U4301 (N_4301,N_3241,N_182);
or U4302 (N_4302,N_1400,N_646);
and U4303 (N_4303,N_2208,N_1476);
and U4304 (N_4304,N_221,N_2197);
nor U4305 (N_4305,N_2491,N_1565);
nor U4306 (N_4306,N_1328,N_2048);
or U4307 (N_4307,N_2398,N_2789);
nand U4308 (N_4308,N_3412,N_580);
nand U4309 (N_4309,N_558,N_3215);
or U4310 (N_4310,N_1414,N_1594);
and U4311 (N_4311,N_3372,N_144);
nand U4312 (N_4312,N_3563,N_3637);
nand U4313 (N_4313,N_2074,N_1609);
and U4314 (N_4314,N_43,N_2839);
nor U4315 (N_4315,N_1477,N_3407);
nand U4316 (N_4316,N_51,N_3597);
and U4317 (N_4317,N_3179,N_2056);
xnor U4318 (N_4318,N_666,N_62);
nor U4319 (N_4319,N_3539,N_162);
nand U4320 (N_4320,N_1935,N_1012);
nor U4321 (N_4321,N_3725,N_2161);
nand U4322 (N_4322,N_3542,N_2356);
nor U4323 (N_4323,N_3112,N_1341);
xor U4324 (N_4324,N_3285,N_3433);
or U4325 (N_4325,N_1439,N_548);
and U4326 (N_4326,N_3839,N_85);
and U4327 (N_4327,N_347,N_550);
xor U4328 (N_4328,N_2162,N_2112);
nor U4329 (N_4329,N_56,N_2379);
and U4330 (N_4330,N_2967,N_3548);
and U4331 (N_4331,N_3703,N_2035);
nand U4332 (N_4332,N_1952,N_3189);
nand U4333 (N_4333,N_1610,N_986);
nand U4334 (N_4334,N_597,N_877);
nand U4335 (N_4335,N_3202,N_297);
xor U4336 (N_4336,N_927,N_1878);
xnor U4337 (N_4337,N_466,N_2);
xnor U4338 (N_4338,N_2868,N_3777);
or U4339 (N_4339,N_791,N_461);
nand U4340 (N_4340,N_1750,N_2107);
nand U4341 (N_4341,N_977,N_419);
and U4342 (N_4342,N_214,N_2088);
xor U4343 (N_4343,N_3103,N_1342);
or U4344 (N_4344,N_3360,N_712);
and U4345 (N_4345,N_94,N_2006);
or U4346 (N_4346,N_2055,N_36);
or U4347 (N_4347,N_2346,N_2959);
nor U4348 (N_4348,N_2610,N_3493);
nor U4349 (N_4349,N_1471,N_800);
nor U4350 (N_4350,N_3834,N_2596);
xnor U4351 (N_4351,N_2751,N_3706);
and U4352 (N_4352,N_3153,N_2783);
nand U4353 (N_4353,N_759,N_435);
or U4354 (N_4354,N_134,N_1835);
nand U4355 (N_4355,N_952,N_152);
and U4356 (N_4356,N_1979,N_1415);
and U4357 (N_4357,N_3495,N_474);
and U4358 (N_4358,N_3852,N_1644);
and U4359 (N_4359,N_3864,N_2265);
nand U4360 (N_4360,N_101,N_3247);
nand U4361 (N_4361,N_3991,N_1646);
nand U4362 (N_4362,N_2668,N_263);
and U4363 (N_4363,N_1888,N_2301);
nor U4364 (N_4364,N_987,N_602);
xnor U4365 (N_4365,N_2408,N_2675);
nor U4366 (N_4366,N_1474,N_627);
or U4367 (N_4367,N_1607,N_3507);
nor U4368 (N_4368,N_2381,N_3530);
nor U4369 (N_4369,N_922,N_3681);
and U4370 (N_4370,N_3968,N_2022);
xor U4371 (N_4371,N_1270,N_1354);
nor U4372 (N_4372,N_372,N_1257);
and U4373 (N_4373,N_2530,N_3133);
nor U4374 (N_4374,N_3439,N_232);
nor U4375 (N_4375,N_616,N_640);
nand U4376 (N_4376,N_3079,N_1406);
nor U4377 (N_4377,N_2854,N_2948);
nor U4378 (N_4378,N_3905,N_2624);
and U4379 (N_4379,N_1785,N_1950);
and U4380 (N_4380,N_286,N_2759);
or U4381 (N_4381,N_3149,N_1402);
nand U4382 (N_4382,N_1108,N_1752);
or U4383 (N_4383,N_2040,N_3323);
or U4384 (N_4384,N_3954,N_849);
and U4385 (N_4385,N_42,N_2559);
or U4386 (N_4386,N_3975,N_1897);
nor U4387 (N_4387,N_715,N_3716);
nand U4388 (N_4388,N_3343,N_2261);
nor U4389 (N_4389,N_271,N_3237);
nand U4390 (N_4390,N_582,N_3796);
xor U4391 (N_4391,N_1355,N_614);
nand U4392 (N_4392,N_3959,N_3741);
nor U4393 (N_4393,N_945,N_1564);
or U4394 (N_4394,N_1863,N_1480);
nand U4395 (N_4395,N_1753,N_2594);
nor U4396 (N_4396,N_167,N_1844);
and U4397 (N_4397,N_3367,N_1515);
nor U4398 (N_4398,N_1573,N_2889);
or U4399 (N_4399,N_2840,N_1090);
nand U4400 (N_4400,N_3347,N_1969);
or U4401 (N_4401,N_1118,N_2677);
nand U4402 (N_4402,N_3508,N_2493);
nand U4403 (N_4403,N_307,N_1314);
and U4404 (N_4404,N_1731,N_1968);
or U4405 (N_4405,N_2507,N_399);
or U4406 (N_4406,N_2798,N_1909);
nor U4407 (N_4407,N_3717,N_1604);
nor U4408 (N_4408,N_3021,N_3811);
and U4409 (N_4409,N_663,N_3368);
nand U4410 (N_4410,N_2654,N_1072);
or U4411 (N_4411,N_3294,N_3476);
nand U4412 (N_4412,N_2890,N_1518);
nor U4413 (N_4413,N_1630,N_2721);
and U4414 (N_4414,N_1005,N_636);
and U4415 (N_4415,N_2623,N_3837);
or U4416 (N_4416,N_1083,N_2129);
nor U4417 (N_4417,N_3559,N_2932);
or U4418 (N_4418,N_3846,N_1177);
nor U4419 (N_4419,N_1769,N_95);
nor U4420 (N_4420,N_453,N_1382);
or U4421 (N_4421,N_2095,N_2211);
xnor U4422 (N_4422,N_2399,N_2204);
or U4423 (N_4423,N_1661,N_408);
and U4424 (N_4424,N_2653,N_3733);
nor U4425 (N_4425,N_2236,N_2760);
and U4426 (N_4426,N_3088,N_2371);
and U4427 (N_4427,N_41,N_2384);
nand U4428 (N_4428,N_1597,N_3399);
nand U4429 (N_4429,N_3277,N_2029);
or U4430 (N_4430,N_2974,N_2517);
nand U4431 (N_4431,N_1001,N_3615);
or U4432 (N_4432,N_2075,N_1220);
xnor U4433 (N_4433,N_68,N_3860);
and U4434 (N_4434,N_3255,N_3252);
nor U4435 (N_4435,N_1433,N_397);
nand U4436 (N_4436,N_1210,N_2357);
xnor U4437 (N_4437,N_3281,N_482);
and U4438 (N_4438,N_2680,N_3520);
nor U4439 (N_4439,N_3724,N_1300);
nand U4440 (N_4440,N_2415,N_3326);
nor U4441 (N_4441,N_137,N_1986);
and U4442 (N_4442,N_3364,N_3475);
or U4443 (N_4443,N_1803,N_1984);
nor U4444 (N_4444,N_2401,N_3223);
and U4445 (N_4445,N_1120,N_2845);
and U4446 (N_4446,N_3009,N_2455);
nor U4447 (N_4447,N_3404,N_3532);
xnor U4448 (N_4448,N_2111,N_404);
or U4449 (N_4449,N_2166,N_3857);
nor U4450 (N_4450,N_55,N_3929);
nand U4451 (N_4451,N_1478,N_2622);
nand U4452 (N_4452,N_15,N_696);
and U4453 (N_4453,N_2028,N_2470);
nor U4454 (N_4454,N_1692,N_2548);
nand U4455 (N_4455,N_2737,N_3251);
or U4456 (N_4456,N_2400,N_1484);
nand U4457 (N_4457,N_2103,N_941);
nand U4458 (N_4458,N_3394,N_2911);
xnor U4459 (N_4459,N_291,N_2057);
or U4460 (N_4460,N_2032,N_3303);
or U4461 (N_4461,N_1291,N_939);
nand U4462 (N_4462,N_876,N_1838);
nand U4463 (N_4463,N_2172,N_2505);
nor U4464 (N_4464,N_3746,N_265);
nand U4465 (N_4465,N_3036,N_3772);
nor U4466 (N_4466,N_533,N_3707);
xor U4467 (N_4467,N_352,N_465);
nand U4468 (N_4468,N_1528,N_3871);
xor U4469 (N_4469,N_2206,N_912);
and U4470 (N_4470,N_2434,N_2393);
or U4471 (N_4471,N_3964,N_3638);
nand U4472 (N_4472,N_850,N_387);
nor U4473 (N_4473,N_84,N_1325);
xor U4474 (N_4474,N_687,N_2259);
nand U4475 (N_4475,N_1625,N_3749);
nor U4476 (N_4476,N_2687,N_190);
or U4477 (N_4477,N_2070,N_2089);
nand U4478 (N_4478,N_2910,N_3757);
or U4479 (N_4479,N_3402,N_2186);
or U4480 (N_4480,N_2336,N_1111);
and U4481 (N_4481,N_3781,N_1790);
nor U4482 (N_4482,N_1143,N_536);
and U4483 (N_4483,N_3389,N_862);
or U4484 (N_4484,N_126,N_1153);
or U4485 (N_4485,N_1561,N_2765);
nor U4486 (N_4486,N_1004,N_2898);
and U4487 (N_4487,N_1544,N_1493);
nand U4488 (N_4488,N_3897,N_3071);
nor U4489 (N_4489,N_817,N_2620);
nor U4490 (N_4490,N_3767,N_1214);
nand U4491 (N_4491,N_1026,N_1837);
nor U4492 (N_4492,N_346,N_3297);
xor U4493 (N_4493,N_2113,N_2681);
nand U4494 (N_4494,N_86,N_2812);
and U4495 (N_4495,N_1563,N_337);
and U4496 (N_4496,N_206,N_1852);
nor U4497 (N_4497,N_708,N_518);
and U4498 (N_4498,N_1389,N_2913);
xnor U4499 (N_4499,N_3662,N_751);
or U4500 (N_4500,N_3170,N_2010);
or U4501 (N_4501,N_2221,N_3410);
and U4502 (N_4502,N_2156,N_918);
nand U4503 (N_4503,N_1076,N_3673);
nor U4504 (N_4504,N_2786,N_2958);
and U4505 (N_4505,N_464,N_401);
or U4506 (N_4506,N_1351,N_1928);
or U4507 (N_4507,N_2141,N_1627);
nor U4508 (N_4508,N_811,N_498);
xnor U4509 (N_4509,N_1981,N_2466);
xor U4510 (N_4510,N_3157,N_866);
and U4511 (N_4511,N_3084,N_669);
and U4512 (N_4512,N_2736,N_3916);
nor U4513 (N_4513,N_1181,N_3225);
and U4514 (N_4514,N_3312,N_264);
nand U4515 (N_4515,N_719,N_3728);
nand U4516 (N_4516,N_2676,N_267);
nor U4517 (N_4517,N_3123,N_1229);
and U4518 (N_4518,N_3862,N_1002);
nand U4519 (N_4519,N_3371,N_2708);
or U4520 (N_4520,N_1178,N_829);
or U4521 (N_4521,N_2000,N_1828);
and U4522 (N_4522,N_1006,N_1944);
xnor U4523 (N_4523,N_3661,N_1912);
or U4524 (N_4524,N_2756,N_1050);
xor U4525 (N_4525,N_1730,N_3957);
nor U4526 (N_4526,N_413,N_3445);
nor U4527 (N_4527,N_3840,N_3634);
nor U4528 (N_4528,N_1501,N_3690);
xor U4529 (N_4529,N_2533,N_393);
nor U4530 (N_4530,N_1363,N_3926);
or U4531 (N_4531,N_3538,N_1042);
nor U4532 (N_4532,N_3522,N_3070);
and U4533 (N_4533,N_1365,N_1386);
nor U4534 (N_4534,N_3664,N_1172);
nor U4535 (N_4535,N_1932,N_3118);
and U4536 (N_4536,N_2138,N_972);
nand U4537 (N_4537,N_2489,N_3116);
nand U4538 (N_4538,N_2406,N_2324);
and U4539 (N_4539,N_2570,N_2830);
nand U4540 (N_4540,N_342,N_2471);
nand U4541 (N_4541,N_2046,N_1358);
or U4542 (N_4542,N_37,N_1437);
nand U4543 (N_4543,N_592,N_1456);
xor U4544 (N_4544,N_2479,N_1183);
or U4545 (N_4545,N_180,N_1110);
nor U4546 (N_4546,N_2939,N_1319);
xnor U4547 (N_4547,N_2790,N_2051);
nand U4548 (N_4548,N_1636,N_2182);
nor U4549 (N_4549,N_1069,N_1145);
nor U4550 (N_4550,N_2818,N_762);
nor U4551 (N_4551,N_2639,N_2285);
or U4552 (N_4552,N_810,N_2354);
nand U4553 (N_4553,N_3671,N_1133);
and U4554 (N_4554,N_2861,N_1576);
xnor U4555 (N_4555,N_2179,N_1921);
nor U4556 (N_4556,N_1,N_3498);
nor U4557 (N_4557,N_2524,N_3835);
nand U4558 (N_4558,N_3059,N_2304);
xor U4559 (N_4559,N_1960,N_2355);
nand U4560 (N_4560,N_3208,N_1985);
nor U4561 (N_4561,N_993,N_3523);
xor U4562 (N_4562,N_2633,N_3903);
and U4563 (N_4563,N_3629,N_418);
and U4564 (N_4564,N_2177,N_3426);
and U4565 (N_4565,N_234,N_3033);
nand U4566 (N_4566,N_2528,N_1211);
nor U4567 (N_4567,N_3244,N_3162);
or U4568 (N_4568,N_1983,N_578);
nor U4569 (N_4569,N_1275,N_2331);
nor U4570 (N_4570,N_2248,N_2445);
or U4571 (N_4571,N_519,N_3385);
nand U4572 (N_4572,N_3008,N_2532);
and U4573 (N_4573,N_1065,N_1649);
or U4574 (N_4574,N_3755,N_3122);
nand U4575 (N_4575,N_2404,N_490);
or U4576 (N_4576,N_2258,N_361);
nand U4577 (N_4577,N_3898,N_2271);
or U4578 (N_4578,N_710,N_1419);
xnor U4579 (N_4579,N_2978,N_887);
nor U4580 (N_4580,N_967,N_727);
nand U4581 (N_4581,N_1698,N_2325);
nand U4582 (N_4582,N_2412,N_2475);
xnor U4583 (N_4583,N_1834,N_1872);
or U4584 (N_4584,N_1485,N_3212);
and U4585 (N_4585,N_3655,N_488);
xor U4586 (N_4586,N_2878,N_3362);
nand U4587 (N_4587,N_78,N_164);
nor U4588 (N_4588,N_1993,N_3578);
and U4589 (N_4589,N_2081,N_1949);
nand U4590 (N_4590,N_3365,N_1103);
nand U4591 (N_4591,N_2689,N_1075);
nor U4592 (N_4592,N_2037,N_459);
nor U4593 (N_4593,N_1489,N_2643);
nor U4594 (N_4594,N_3486,N_2134);
and U4595 (N_4595,N_3400,N_2953);
or U4596 (N_4596,N_2279,N_1311);
nor U4597 (N_4597,N_2299,N_843);
nor U4598 (N_4598,N_3752,N_2096);
nor U4599 (N_4599,N_2215,N_1147);
nor U4600 (N_4600,N_1322,N_133);
and U4601 (N_4601,N_2945,N_528);
nor U4602 (N_4602,N_3984,N_306);
and U4603 (N_4603,N_2841,N_3780);
and U4604 (N_4604,N_1331,N_426);
or U4605 (N_4605,N_3841,N_2472);
nand U4606 (N_4606,N_1900,N_132);
nor U4607 (N_4607,N_1965,N_3884);
nor U4608 (N_4608,N_1308,N_966);
or U4609 (N_4609,N_2435,N_2314);
and U4610 (N_4610,N_3354,N_2552);
nand U4611 (N_4611,N_3473,N_2908);
nand U4612 (N_4612,N_3691,N_1749);
xor U4613 (N_4613,N_2352,N_2465);
nand U4614 (N_4614,N_3901,N_1243);
or U4615 (N_4615,N_617,N_1893);
and U4616 (N_4616,N_2490,N_2255);
or U4617 (N_4617,N_881,N_424);
xor U4618 (N_4618,N_534,N_1531);
or U4619 (N_4619,N_3173,N_3159);
nand U4620 (N_4620,N_1068,N_1885);
and U4621 (N_4621,N_795,N_400);
or U4622 (N_4622,N_261,N_3863);
nand U4623 (N_4623,N_2605,N_2696);
nand U4624 (N_4624,N_1247,N_3013);
or U4625 (N_4625,N_2720,N_2954);
and U4626 (N_4626,N_572,N_3649);
xor U4627 (N_4627,N_1372,N_18);
and U4628 (N_4628,N_3537,N_2327);
or U4629 (N_4629,N_46,N_2641);
nand U4630 (N_4630,N_2666,N_2453);
nand U4631 (N_4631,N_1208,N_2722);
and U4632 (N_4632,N_1892,N_929);
xnor U4633 (N_4633,N_3962,N_2023);
xnor U4634 (N_4634,N_1235,N_2430);
nand U4635 (N_4635,N_1708,N_1813);
nor U4636 (N_4636,N_684,N_2360);
xnor U4637 (N_4637,N_594,N_3972);
or U4638 (N_4638,N_3447,N_300);
and U4639 (N_4639,N_3797,N_2083);
nand U4640 (N_4640,N_313,N_1737);
nor U4641 (N_4641,N_470,N_1619);
or U4642 (N_4642,N_1017,N_257);
or U4643 (N_4643,N_3545,N_2143);
nor U4644 (N_4644,N_69,N_3653);
nor U4645 (N_4645,N_1159,N_2851);
or U4646 (N_4646,N_2823,N_3146);
or U4647 (N_4647,N_2233,N_2678);
nor U4648 (N_4648,N_3506,N_2525);
or U4649 (N_4649,N_1745,N_3694);
xnor U4650 (N_4650,N_809,N_1279);
xor U4651 (N_4651,N_1022,N_3744);
nor U4652 (N_4652,N_445,N_3327);
and U4653 (N_4653,N_1706,N_886);
nor U4654 (N_4654,N_2064,N_516);
xor U4655 (N_4655,N_3823,N_2659);
nor U4656 (N_4656,N_296,N_1333);
xnor U4657 (N_4657,N_1534,N_1977);
nor U4658 (N_4658,N_2894,N_2502);
nand U4659 (N_4659,N_2690,N_1197);
and U4660 (N_4660,N_2587,N_438);
and U4661 (N_4661,N_693,N_2813);
nor U4662 (N_4662,N_3735,N_325);
nand U4663 (N_4663,N_2246,N_2729);
nor U4664 (N_4664,N_2433,N_3174);
nor U4665 (N_4665,N_590,N_982);
or U4666 (N_4666,N_1013,N_1219);
and U4667 (N_4667,N_2557,N_957);
and U4668 (N_4668,N_872,N_2091);
nor U4669 (N_4669,N_3053,N_1595);
nor U4670 (N_4670,N_1201,N_1859);
or U4671 (N_4671,N_1000,N_2588);
nand U4672 (N_4672,N_660,N_3342);
nor U4673 (N_4673,N_511,N_284);
nor U4674 (N_4674,N_345,N_507);
nor U4675 (N_4675,N_1066,N_362);
and U4676 (N_4676,N_103,N_3677);
nor U4677 (N_4677,N_2647,N_485);
or U4678 (N_4678,N_2125,N_1425);
nand U4679 (N_4679,N_1908,N_1317);
nor U4680 (N_4680,N_3479,N_2460);
xnor U4681 (N_4681,N_57,N_1875);
nand U4682 (N_4682,N_3308,N_3865);
xnor U4683 (N_4683,N_1660,N_2583);
or U4684 (N_4684,N_3106,N_2292);
or U4685 (N_4685,N_2598,N_1007);
nor U4686 (N_4686,N_856,N_3043);
nor U4687 (N_4687,N_166,N_1867);
or U4688 (N_4688,N_3892,N_1634);
nor U4689 (N_4689,N_1438,N_659);
nand U4690 (N_4690,N_3813,N_2987);
nor U4691 (N_4691,N_2322,N_3550);
nand U4692 (N_4692,N_3727,N_2087);
nor U4693 (N_4693,N_3226,N_3612);
nand U4694 (N_4694,N_1086,N_2446);
nor U4695 (N_4695,N_1023,N_1041);
nor U4696 (N_4696,N_1185,N_1865);
nand U4697 (N_4697,N_3040,N_1796);
nand U4698 (N_4698,N_1626,N_3292);
nand U4699 (N_4699,N_3874,N_1262);
nand U4700 (N_4700,N_31,N_3374);
nand U4701 (N_4701,N_2066,N_2005);
nor U4702 (N_4702,N_608,N_3214);
nor U4703 (N_4703,N_1251,N_506);
or U4704 (N_4704,N_1390,N_964);
nor U4705 (N_4705,N_794,N_618);
nor U4706 (N_4706,N_3129,N_2891);
nand U4707 (N_4707,N_3016,N_2537);
or U4708 (N_4708,N_3760,N_2673);
or U4709 (N_4709,N_2859,N_564);
nor U4710 (N_4710,N_3379,N_2777);
nand U4711 (N_4711,N_937,N_2976);
or U4712 (N_4712,N_1301,N_3574);
nand U4713 (N_4713,N_392,N_1799);
nor U4714 (N_4714,N_428,N_1910);
and U4715 (N_4715,N_3618,N_728);
xor U4716 (N_4716,N_2972,N_285);
and U4717 (N_4717,N_2428,N_775);
nand U4718 (N_4718,N_750,N_315);
xnor U4719 (N_4719,N_732,N_1117);
and U4720 (N_4720,N_3152,N_1807);
xnor U4721 (N_4721,N_1637,N_109);
and U4722 (N_4722,N_2863,N_3457);
or U4723 (N_4723,N_11,N_3751);
xnor U4724 (N_4724,N_331,N_1781);
nor U4725 (N_4725,N_1975,N_3556);
nor U4726 (N_4726,N_607,N_3560);
and U4727 (N_4727,N_1230,N_3256);
nand U4728 (N_4728,N_683,N_2752);
or U4729 (N_4729,N_2217,N_1309);
nand U4730 (N_4730,N_1948,N_629);
and U4731 (N_4731,N_1620,N_2980);
or U4732 (N_4732,N_1296,N_3011);
nand U4733 (N_4733,N_341,N_1931);
and U4734 (N_4734,N_1062,N_2425);
and U4735 (N_4735,N_671,N_915);
or U4736 (N_4736,N_538,N_123);
and U4737 (N_4737,N_1073,N_1492);
nor U4738 (N_4738,N_79,N_3054);
nor U4739 (N_4739,N_2969,N_3454);
nor U4740 (N_4740,N_3114,N_2026);
nor U4741 (N_4741,N_3046,N_114);
and U4742 (N_4742,N_3576,N_3435);
or U4743 (N_4743,N_2716,N_3566);
or U4744 (N_4744,N_2734,N_248);
and U4745 (N_4745,N_1973,N_371);
nand U4746 (N_4746,N_3998,N_1195);
xnor U4747 (N_4747,N_1030,N_3602);
nand U4748 (N_4748,N_985,N_2163);
and U4749 (N_4749,N_2383,N_2743);
nand U4750 (N_4750,N_3881,N_1499);
xor U4751 (N_4751,N_1376,N_1946);
xnor U4752 (N_4752,N_637,N_1058);
and U4753 (N_4753,N_2334,N_2450);
or U4754 (N_4754,N_2367,N_3895);
nand U4755 (N_4755,N_3095,N_2771);
nor U4756 (N_4756,N_2160,N_3282);
nor U4757 (N_4757,N_3168,N_3311);
xnor U4758 (N_4758,N_81,N_869);
nand U4759 (N_4759,N_2176,N_3783);
and U4760 (N_4760,N_90,N_3267);
and U4761 (N_4761,N_1297,N_2345);
xnor U4762 (N_4762,N_2719,N_1821);
nor U4763 (N_4763,N_3771,N_724);
nor U4764 (N_4764,N_2468,N_143);
xor U4765 (N_4765,N_1869,N_3791);
and U4766 (N_4766,N_3171,N_3657);
nand U4767 (N_4767,N_2657,N_2076);
and U4768 (N_4768,N_3131,N_2842);
nand U4769 (N_4769,N_3055,N_427);
and U4770 (N_4770,N_2041,N_2108);
nor U4771 (N_4771,N_3696,N_999);
nor U4772 (N_4772,N_3541,N_2058);
and U4773 (N_4773,N_3358,N_1222);
and U4774 (N_4774,N_1452,N_1087);
and U4775 (N_4775,N_2607,N_761);
xor U4776 (N_4776,N_3712,N_2362);
nand U4777 (N_4777,N_3462,N_1587);
xnor U4778 (N_4778,N_641,N_3931);
nand U4779 (N_4779,N_3086,N_1024);
and U4780 (N_4780,N_2644,N_593);
nand U4781 (N_4781,N_1766,N_1031);
nor U4782 (N_4782,N_1523,N_981);
nor U4783 (N_4783,N_2656,N_2413);
or U4784 (N_4784,N_108,N_2223);
nand U4785 (N_4785,N_2872,N_789);
nor U4786 (N_4786,N_3348,N_481);
or U4787 (N_4787,N_209,N_328);
nor U4788 (N_4788,N_623,N_779);
nand U4789 (N_4789,N_3516,N_1738);
xnor U4790 (N_4790,N_1990,N_1690);
nor U4791 (N_4791,N_3099,N_1427);
or U4792 (N_4792,N_771,N_568);
or U4793 (N_4793,N_806,N_2682);
and U4794 (N_4794,N_1374,N_1667);
nor U4795 (N_4795,N_2370,N_831);
and U4796 (N_4796,N_1252,N_2185);
or U4797 (N_4797,N_2833,N_2152);
or U4798 (N_4798,N_542,N_54);
and U4799 (N_4799,N_3184,N_2547);
and U4800 (N_4800,N_3265,N_1947);
nor U4801 (N_4801,N_3234,N_2175);
nand U4802 (N_4802,N_959,N_268);
nand U4803 (N_4803,N_3069,N_1163);
nor U4804 (N_4804,N_3395,N_612);
nand U4805 (N_4805,N_2286,N_2565);
nand U4806 (N_4806,N_91,N_2923);
and U4807 (N_4807,N_839,N_844);
nor U4808 (N_4808,N_3384,N_2280);
or U4809 (N_4809,N_537,N_1194);
nand U4810 (N_4810,N_2698,N_3977);
and U4811 (N_4811,N_1733,N_1098);
and U4812 (N_4812,N_2935,N_1582);
and U4813 (N_4813,N_3272,N_587);
nand U4814 (N_4814,N_2106,N_910);
nand U4815 (N_4815,N_222,N_1744);
nor U4816 (N_4816,N_1703,N_1138);
nand U4817 (N_4817,N_2136,N_410);
or U4818 (N_4818,N_3111,N_3934);
nand U4819 (N_4819,N_1819,N_3726);
or U4820 (N_4820,N_2996,N_1907);
and U4821 (N_4821,N_239,N_1734);
or U4822 (N_4822,N_3422,N_1435);
or U4823 (N_4823,N_2174,N_3438);
or U4824 (N_4824,N_2648,N_3587);
or U4825 (N_4825,N_33,N_1617);
or U4826 (N_4826,N_2849,N_545);
nor U4827 (N_4827,N_717,N_3182);
nand U4828 (N_4828,N_577,N_3073);
or U4829 (N_4829,N_1808,N_1061);
nor U4830 (N_4830,N_442,N_2794);
xnor U4831 (N_4831,N_543,N_2410);
nor U4832 (N_4832,N_2047,N_2376);
and U4833 (N_4833,N_1583,N_1224);
nor U4834 (N_4834,N_279,N_3275);
nor U4835 (N_4835,N_1152,N_2982);
nor U4836 (N_4836,N_1727,N_1726);
nor U4837 (N_4837,N_3645,N_236);
nand U4838 (N_4838,N_2600,N_1027);
nand U4839 (N_4839,N_2795,N_2928);
nand U4840 (N_4840,N_443,N_3993);
xor U4841 (N_4841,N_412,N_2281);
or U4842 (N_4842,N_591,N_298);
or U4843 (N_4843,N_865,N_2739);
nand U4844 (N_4844,N_1868,N_2002);
nand U4845 (N_4845,N_441,N_3963);
nor U4846 (N_4846,N_1399,N_3510);
xor U4847 (N_4847,N_2073,N_432);
nor U4848 (N_4848,N_2929,N_3943);
or U4849 (N_4849,N_329,N_2801);
and U4850 (N_4850,N_975,N_3546);
nand U4851 (N_4851,N_340,N_299);
nand U4852 (N_4852,N_1088,N_3827);
and U4853 (N_4853,N_737,N_118);
nand U4854 (N_4854,N_3980,N_1417);
and U4855 (N_4855,N_29,N_1671);
nor U4856 (N_4856,N_797,N_2219);
and U4857 (N_4857,N_1278,N_2661);
or U4858 (N_4858,N_1125,N_1450);
or U4859 (N_4859,N_2452,N_92);
and U4860 (N_4860,N_1718,N_2784);
nor U4861 (N_4861,N_2043,N_3039);
and U4862 (N_4862,N_2855,N_2550);
nand U4863 (N_4863,N_2431,N_3280);
xnor U4864 (N_4864,N_1529,N_1124);
and U4865 (N_4865,N_2917,N_3656);
and U4866 (N_4866,N_3489,N_1466);
or U4867 (N_4867,N_3792,N_3723);
and U4868 (N_4868,N_2164,N_2800);
nor U4869 (N_4869,N_3437,N_370);
nor U4870 (N_4870,N_168,N_3213);
or U4871 (N_4871,N_824,N_1011);
and U4872 (N_4872,N_3145,N_2213);
or U4873 (N_4873,N_336,N_3393);
nor U4874 (N_4874,N_3136,N_2313);
or U4875 (N_4875,N_3594,N_714);
xor U4876 (N_4876,N_1212,N_2497);
nor U4877 (N_4877,N_1512,N_3584);
xnor U4878 (N_4878,N_1797,N_1407);
nand U4879 (N_4879,N_1956,N_3351);
xor U4880 (N_4880,N_2616,N_150);
xor U4881 (N_4881,N_3034,N_2282);
and U4882 (N_4882,N_2621,N_1504);
or U4883 (N_4883,N_294,N_3648);
or U4884 (N_4884,N_1364,N_497);
and U4885 (N_4885,N_3877,N_2906);
xor U4886 (N_4886,N_570,N_1294);
xnor U4887 (N_4887,N_2509,N_3499);
nand U4888 (N_4888,N_2456,N_2287);
nand U4889 (N_4889,N_3858,N_1550);
and U4890 (N_4890,N_556,N_502);
nand U4891 (N_4891,N_3236,N_3699);
or U4892 (N_4892,N_2572,N_48);
nor U4893 (N_4893,N_3812,N_2283);
and U4894 (N_4894,N_255,N_670);
and U4895 (N_4895,N_755,N_2914);
nand U4896 (N_4896,N_2335,N_1481);
xnor U4897 (N_4897,N_3540,N_1877);
and U4898 (N_4898,N_3737,N_3855);
and U4899 (N_4899,N_2209,N_583);
and U4900 (N_4900,N_3357,N_2191);
nor U4901 (N_4901,N_504,N_3614);
nand U4902 (N_4902,N_1611,N_1999);
nand U4903 (N_4903,N_3670,N_1829);
xnor U4904 (N_4904,N_2234,N_3203);
nor U4905 (N_4905,N_437,N_478);
or U4906 (N_4906,N_2741,N_1546);
nor U4907 (N_4907,N_2625,N_2726);
and U4908 (N_4908,N_3766,N_1811);
or U4909 (N_4909,N_2303,N_697);
and U4910 (N_4910,N_3795,N_766);
or U4911 (N_4911,N_1663,N_976);
nor U4912 (N_4912,N_1395,N_2754);
and U4913 (N_4913,N_812,N_3229);
nand U4914 (N_4914,N_3020,N_3944);
and U4915 (N_4915,N_2989,N_2059);
or U4916 (N_4916,N_3010,N_3076);
or U4917 (N_4917,N_3814,N_3816);
or U4918 (N_4918,N_3488,N_1855);
nand U4919 (N_4919,N_595,N_2897);
xor U4920 (N_4920,N_3970,N_2180);
nand U4921 (N_4921,N_628,N_1714);
or U4922 (N_4922,N_2807,N_3952);
or U4923 (N_4923,N_3748,N_3682);
xor U4924 (N_4924,N_711,N_3734);
or U4925 (N_4925,N_429,N_557);
or U4926 (N_4926,N_1109,N_1396);
and U4927 (N_4927,N_2419,N_672);
nor U4928 (N_4928,N_871,N_32);
and U4929 (N_4929,N_449,N_2770);
and U4930 (N_4930,N_1930,N_1206);
nand U4931 (N_4931,N_3922,N_1495);
or U4932 (N_4932,N_757,N_2054);
nand U4933 (N_4933,N_2991,N_1121);
nand U4934 (N_4934,N_172,N_3328);
or U4935 (N_4935,N_1010,N_2121);
nor U4936 (N_4936,N_613,N_2946);
nand U4937 (N_4937,N_777,N_3329);
or U4938 (N_4938,N_2924,N_2225);
nor U4939 (N_4939,N_3205,N_266);
or U4940 (N_4940,N_1635,N_2955);
nand U4941 (N_4941,N_3921,N_1792);
nor U4942 (N_4942,N_3459,N_204);
and U4943 (N_4943,N_355,N_2205);
xnor U4944 (N_4944,N_1055,N_3617);
nor U4945 (N_4945,N_2252,N_584);
xor U4946 (N_4946,N_2196,N_1236);
or U4947 (N_4947,N_1918,N_3701);
and U4948 (N_4948,N_2260,N_416);
nor U4949 (N_4949,N_3465,N_3983);
nor U4950 (N_4950,N_3333,N_705);
and U4951 (N_4951,N_1199,N_3570);
nor U4952 (N_4952,N_631,N_1830);
nand U4953 (N_4953,N_3427,N_1505);
or U4954 (N_4954,N_652,N_3227);
nor U4955 (N_4955,N_1687,N_971);
nand U4956 (N_4956,N_2013,N_289);
xor U4957 (N_4957,N_924,N_3413);
and U4958 (N_4958,N_3973,N_2386);
or U4959 (N_4959,N_333,N_3579);
nand U4960 (N_4960,N_326,N_1884);
or U4961 (N_4961,N_1729,N_1758);
nor U4962 (N_4962,N_2501,N_1923);
and U4963 (N_4963,N_2888,N_632);
and U4964 (N_4964,N_3144,N_3960);
nor U4965 (N_4965,N_690,N_3549);
and U4966 (N_4966,N_3451,N_3586);
xnor U4967 (N_4967,N_1569,N_2097);
xor U4968 (N_4968,N_2044,N_1915);
nor U4969 (N_4969,N_834,N_979);
and U4970 (N_4970,N_2119,N_2302);
nand U4971 (N_4971,N_780,N_139);
xor U4972 (N_4972,N_231,N_1160);
or U4973 (N_4973,N_2218,N_2133);
or U4974 (N_4974,N_173,N_3167);
or U4975 (N_4975,N_191,N_1401);
nor U4976 (N_4976,N_532,N_153);
nor U4977 (N_4977,N_3177,N_2222);
nor U4978 (N_4978,N_2347,N_503);
or U4979 (N_4979,N_1460,N_2569);
nor U4980 (N_4980,N_2288,N_3971);
xor U4981 (N_4981,N_1059,N_3143);
nor U4982 (N_4982,N_64,N_2920);
nor U4983 (N_4983,N_2883,N_2988);
or U4984 (N_4984,N_2896,N_3769);
xor U4985 (N_4985,N_3014,N_1809);
or U4986 (N_4986,N_3714,N_2375);
or U4987 (N_4987,N_2630,N_1553);
and U4988 (N_4988,N_3121,N_1388);
or U4989 (N_4989,N_514,N_2159);
or U4990 (N_4990,N_892,N_375);
xor U4991 (N_4991,N_3740,N_2561);
or U4992 (N_4992,N_1370,N_3822);
or U4993 (N_4993,N_3630,N_1978);
nand U4994 (N_4994,N_3049,N_3417);
or U4995 (N_4995,N_549,N_1043);
and U4996 (N_4996,N_1254,N_141);
and U4997 (N_4997,N_1557,N_1874);
or U4998 (N_4998,N_195,N_1464);
and U4999 (N_4999,N_2857,N_3388);
and U5000 (N_5000,N_3194,N_1638);
nand U5001 (N_5001,N_2416,N_477);
and U5002 (N_5002,N_1451,N_2599);
xnor U5003 (N_5003,N_2592,N_3117);
nor U5004 (N_5004,N_1705,N_725);
nand U5005 (N_5005,N_673,N_310);
nand U5006 (N_5006,N_3336,N_2369);
nand U5007 (N_5007,N_916,N_357);
and U5008 (N_5008,N_66,N_3718);
nor U5009 (N_5009,N_2132,N_815);
nand U5010 (N_5010,N_2646,N_3641);
nand U5011 (N_5011,N_1375,N_773);
or U5012 (N_5012,N_1280,N_3674);
nor U5013 (N_5013,N_920,N_2230);
or U5014 (N_5014,N_3562,N_1033);
and U5015 (N_5015,N_3109,N_1937);
or U5016 (N_5016,N_500,N_174);
nand U5017 (N_5017,N_2480,N_713);
or U5018 (N_5018,N_1095,N_1164);
nand U5019 (N_5019,N_2814,N_3986);
nand U5020 (N_5020,N_3271,N_599);
and U5021 (N_5021,N_2458,N_2578);
or U5022 (N_5022,N_807,N_1559);
or U5023 (N_5023,N_3705,N_3961);
nor U5024 (N_5024,N_882,N_3536);
nand U5025 (N_5025,N_1091,N_2884);
xnor U5026 (N_5026,N_770,N_596);
or U5027 (N_5027,N_3019,N_3869);
and U5028 (N_5028,N_3082,N_2391);
nand U5029 (N_5029,N_2753,N_3340);
xor U5030 (N_5030,N_6,N_781);
nand U5031 (N_5031,N_1548,N_14);
and U5032 (N_5032,N_1409,N_1640);
nand U5033 (N_5033,N_2649,N_647);
or U5034 (N_5034,N_3820,N_3127);
or U5035 (N_5035,N_2008,N_469);
and U5036 (N_5036,N_3660,N_2239);
or U5037 (N_5037,N_1468,N_3471);
and U5038 (N_5038,N_2315,N_2723);
nor U5039 (N_5039,N_3936,N_1443);
nand U5040 (N_5040,N_3958,N_2895);
nor U5041 (N_5041,N_3463,N_2068);
nand U5042 (N_5042,N_3186,N_3504);
or U5043 (N_5043,N_603,N_1440);
nand U5044 (N_5044,N_281,N_3800);
nand U5045 (N_5045,N_1379,N_324);
xor U5046 (N_5046,N_23,N_748);
nor U5047 (N_5047,N_2909,N_2705);
and U5048 (N_5048,N_3148,N_1391);
nand U5049 (N_5049,N_3273,N_3139);
or U5050 (N_5050,N_517,N_468);
or U5051 (N_5051,N_1789,N_3643);
or U5052 (N_5052,N_2998,N_3909);
or U5053 (N_5053,N_2250,N_472);
nand U5054 (N_5054,N_702,N_1657);
or U5055 (N_5055,N_826,N_799);
nor U5056 (N_5056,N_2685,N_2604);
or U5057 (N_5057,N_531,N_3455);
or U5058 (N_5058,N_846,N_1538);
xor U5059 (N_5059,N_2195,N_3132);
xnor U5060 (N_5060,N_1264,N_2511);
nand U5061 (N_5061,N_958,N_2856);
xnor U5062 (N_5062,N_3228,N_744);
xnor U5063 (N_5063,N_3324,N_3380);
or U5064 (N_5064,N_2341,N_1292);
nor U5065 (N_5065,N_2663,N_2273);
and U5066 (N_5066,N_3429,N_1253);
nand U5067 (N_5067,N_734,N_854);
or U5068 (N_5068,N_3678,N_2724);
nor U5069 (N_5069,N_423,N_2144);
and U5070 (N_5070,N_1350,N_2464);
or U5071 (N_5071,N_973,N_2019);
or U5072 (N_5072,N_753,N_275);
and U5073 (N_5073,N_303,N_1586);
nor U5074 (N_5074,N_2793,N_3575);
and U5075 (N_5075,N_2862,N_3334);
nor U5076 (N_5076,N_3900,N_980);
or U5077 (N_5077,N_909,N_1213);
nor U5078 (N_5078,N_440,N_2018);
nand U5079 (N_5079,N_679,N_653);
nand U5080 (N_5080,N_479,N_2319);
and U5081 (N_5081,N_3135,N_3338);
nand U5082 (N_5082,N_1198,N_1927);
or U5083 (N_5083,N_3196,N_2821);
nand U5084 (N_5084,N_1593,N_1154);
nand U5085 (N_5085,N_3754,N_1940);
nand U5086 (N_5086,N_1337,N_2918);
and U5087 (N_5087,N_731,N_1165);
nor U5088 (N_5088,N_3278,N_3815);
or U5089 (N_5089,N_828,N_1903);
xor U5090 (N_5090,N_3344,N_3573);
or U5091 (N_5091,N_2652,N_244);
and U5092 (N_5092,N_3885,N_3784);
nor U5093 (N_5093,N_1603,N_3058);
or U5094 (N_5094,N_2102,N_3913);
xnor U5095 (N_5095,N_1815,N_1018);
and U5096 (N_5096,N_202,N_3555);
xnor U5097 (N_5097,N_1412,N_2877);
nand U5098 (N_5098,N_220,N_3628);
or U5099 (N_5099,N_3313,N_3589);
and U5100 (N_5100,N_2826,N_1786);
nand U5101 (N_5101,N_2473,N_2344);
nor U5102 (N_5102,N_446,N_1772);
nand U5103 (N_5103,N_509,N_2454);
or U5104 (N_5104,N_3956,N_3654);
nor U5105 (N_5105,N_2999,N_3698);
and U5106 (N_5106,N_664,N_3051);
xnor U5107 (N_5107,N_2516,N_3141);
and U5108 (N_5108,N_1740,N_1273);
nor U5109 (N_5109,N_3832,N_2828);
nor U5110 (N_5110,N_3683,N_146);
or U5111 (N_5111,N_1994,N_3004);
nor U5112 (N_5112,N_2417,N_1122);
or U5113 (N_5113,N_898,N_2665);
or U5114 (N_5114,N_2773,N_3531);
nor U5115 (N_5115,N_1431,N_1387);
nand U5116 (N_5116,N_425,N_2542);
or U5117 (N_5117,N_3468,N_674);
and U5118 (N_5118,N_3406,N_991);
nand U5119 (N_5119,N_3619,N_2563);
or U5120 (N_5120,N_611,N_2713);
and U5121 (N_5121,N_58,N_1428);
xor U5122 (N_5122,N_3535,N_1393);
nand U5123 (N_5123,N_3756,N_3613);
and U5124 (N_5124,N_451,N_3201);
or U5125 (N_5125,N_2634,N_2291);
or U5126 (N_5126,N_3134,N_2228);
or U5127 (N_5127,N_3616,N_1085);
nand U5128 (N_5128,N_700,N_1672);
nand U5129 (N_5129,N_369,N_2207);
and U5130 (N_5130,N_1866,N_3);
nor U5131 (N_5131,N_3421,N_1245);
nand U5132 (N_5132,N_1911,N_2733);
xnor U5133 (N_5133,N_89,N_1632);
nand U5134 (N_5134,N_3074,N_1411);
or U5135 (N_5135,N_1654,N_1047);
nor U5136 (N_5136,N_3301,N_1936);
or U5137 (N_5137,N_3142,N_1773);
or U5138 (N_5138,N_348,N_1886);
and U5139 (N_5139,N_161,N_1232);
nand U5140 (N_5140,N_3513,N_3590);
nand U5141 (N_5141,N_3325,N_1933);
or U5142 (N_5142,N_3235,N_1064);
nor U5143 (N_5143,N_2808,N_654);
or U5144 (N_5144,N_2822,N_1421);
nand U5145 (N_5145,N_2632,N_1413);
nor U5146 (N_5146,N_381,N_2342);
and U5147 (N_5147,N_1913,N_1242);
xnor U5148 (N_5148,N_1101,N_3593);
nand U5149 (N_5149,N_407,N_1567);
nand U5150 (N_5150,N_1276,N_3810);
nor U5151 (N_5151,N_2782,N_3204);
nor U5152 (N_5152,N_98,N_1416);
xor U5153 (N_5153,N_527,N_3873);
and U5154 (N_5154,N_1003,N_2099);
xor U5155 (N_5155,N_763,N_1334);
or U5156 (N_5156,N_2294,N_1942);
or U5157 (N_5157,N_3350,N_902);
nand U5158 (N_5158,N_3478,N_389);
and U5159 (N_5159,N_1132,N_2747);
or U5160 (N_5160,N_1290,N_323);
xnor U5161 (N_5161,N_3715,N_897);
nand U5162 (N_5162,N_3322,N_3558);
or U5163 (N_5163,N_480,N_1526);
xor U5164 (N_5164,N_2009,N_1345);
nor U5165 (N_5165,N_1823,N_940);
xnor U5166 (N_5166,N_245,N_327);
and U5167 (N_5167,N_3432,N_1589);
and U5168 (N_5168,N_2571,N_3790);
or U5169 (N_5169,N_3875,N_3838);
or U5170 (N_5170,N_171,N_3945);
xnor U5171 (N_5171,N_3761,N_2411);
and U5172 (N_5172,N_1759,N_19);
nor U5173 (N_5173,N_889,N_2585);
nand U5174 (N_5174,N_2358,N_680);
xnor U5175 (N_5175,N_3339,N_1951);
nand U5176 (N_5176,N_1092,N_793);
nand U5177 (N_5177,N_2820,N_2774);
and U5178 (N_5178,N_194,N_3830);
xnor U5179 (N_5179,N_431,N_344);
nor U5180 (N_5180,N_2703,N_1507);
nor U5181 (N_5181,N_1715,N_13);
or U5182 (N_5182,N_2389,N_2584);
nand U5183 (N_5183,N_160,N_784);
or U5184 (N_5184,N_896,N_3509);
or U5185 (N_5185,N_1917,N_1161);
nand U5186 (N_5186,N_2776,N_186);
nand U5187 (N_5187,N_129,N_3543);
nor U5188 (N_5188,N_1259,N_3209);
or U5189 (N_5189,N_853,N_1599);
nor U5190 (N_5190,N_2114,N_196);
nand U5191 (N_5191,N_749,N_649);
or U5192 (N_5192,N_2508,N_928);
and U5193 (N_5193,N_2990,N_2038);
nand U5194 (N_5194,N_181,N_1929);
or U5195 (N_5195,N_2210,N_3675);
and U5196 (N_5196,N_3138,N_373);
nor U5197 (N_5197,N_3974,N_2568);
or U5198 (N_5198,N_2310,N_1028);
or U5199 (N_5199,N_1919,N_2149);
nand U5200 (N_5200,N_2390,N_2120);
xor U5201 (N_5201,N_551,N_651);
and U5202 (N_5202,N_3464,N_2123);
nor U5203 (N_5203,N_3665,N_499);
nand U5204 (N_5204,N_2512,N_2153);
or U5205 (N_5205,N_318,N_1025);
nor U5206 (N_5206,N_3291,N_70);
xnor U5207 (N_5207,N_125,N_948);
or U5208 (N_5208,N_944,N_1681);
xnor U5209 (N_5209,N_3557,N_701);
and U5210 (N_5210,N_1664,N_2901);
nand U5211 (N_5211,N_201,N_851);
or U5212 (N_5212,N_3779,N_2039);
nor U5213 (N_5213,N_541,N_2712);
nand U5214 (N_5214,N_703,N_277);
or U5215 (N_5215,N_2276,N_179);
and U5216 (N_5216,N_2638,N_2626);
nor U5217 (N_5217,N_1020,N_359);
or U5218 (N_5218,N_3988,N_3155);
nor U5219 (N_5219,N_3719,N_170);
or U5220 (N_5220,N_2949,N_1045);
nor U5221 (N_5221,N_1541,N_888);
nor U5222 (N_5222,N_3452,N_308);
or U5223 (N_5223,N_1140,N_1016);
nand U5224 (N_5224,N_3346,N_2873);
nor U5225 (N_5225,N_2943,N_2249);
and U5226 (N_5226,N_3018,N_682);
or U5227 (N_5227,N_3636,N_131);
or U5228 (N_5228,N_586,N_601);
nand U5229 (N_5229,N_2243,N_3500);
or U5230 (N_5230,N_1306,N_1788);
and U5231 (N_5231,N_2700,N_3240);
and U5232 (N_5232,N_3985,N_1847);
or U5233 (N_5233,N_2963,N_2535);
nand U5234 (N_5234,N_3554,N_2824);
xnor U5235 (N_5235,N_3515,N_3029);
nand U5236 (N_5236,N_1666,N_335);
or U5237 (N_5237,N_3335,N_2127);
nor U5238 (N_5238,N_1187,N_317);
xor U5239 (N_5239,N_3782,N_1810);
and U5240 (N_5240,N_1082,N_874);
or U5241 (N_5241,N_2045,N_769);
or U5242 (N_5242,N_691,N_2791);
nand U5243 (N_5243,N_3802,N_3469);
nor U5244 (N_5244,N_1283,N_3183);
nor U5245 (N_5245,N_704,N_1517);
nand U5246 (N_5246,N_524,N_2555);
nor U5247 (N_5247,N_3310,N_3906);
or U5248 (N_5248,N_1261,N_934);
nand U5249 (N_5249,N_243,N_3893);
or U5250 (N_5250,N_3246,N_3583);
nand U5251 (N_5251,N_2701,N_923);
nor U5252 (N_5252,N_3300,N_2879);
nor U5253 (N_5253,N_2395,N_848);
or U5254 (N_5254,N_207,N_1329);
and U5255 (N_5255,N_1645,N_1067);
nand U5256 (N_5256,N_2981,N_3431);
nor U5257 (N_5257,N_878,N_1078);
nand U5258 (N_5258,N_1250,N_110);
and U5259 (N_5259,N_1748,N_3007);
and U5260 (N_5260,N_983,N_1697);
nor U5261 (N_5261,N_1513,N_2025);
nor U5262 (N_5262,N_1696,N_520);
nor U5263 (N_5263,N_740,N_723);
nor U5264 (N_5264,N_1787,N_2942);
and U5265 (N_5265,N_2926,N_2326);
xor U5266 (N_5266,N_2309,N_366);
or U5267 (N_5267,N_661,N_2764);
xor U5268 (N_5268,N_3178,N_1040);
nor U5269 (N_5269,N_1764,N_2423);
or U5270 (N_5270,N_3105,N_678);
nand U5271 (N_5271,N_3481,N_2394);
nor U5272 (N_5272,N_1204,N_2194);
nand U5273 (N_5273,N_3709,N_859);
nand U5274 (N_5274,N_2264,N_2135);
or U5275 (N_5275,N_260,N_99);
nor U5276 (N_5276,N_3239,N_840);
and U5277 (N_5277,N_1962,N_1606);
or U5278 (N_5278,N_339,N_1470);
xor U5279 (N_5279,N_3187,N_1554);
and U5280 (N_5280,N_1260,N_2718);
xor U5281 (N_5281,N_1675,N_1179);
and U5282 (N_5282,N_2804,N_1724);
nor U5283 (N_5283,N_540,N_1188);
nor U5284 (N_5284,N_396,N_53);
and U5285 (N_5285,N_3081,N_3063);
nor U5286 (N_5286,N_3458,N_1107);
nand U5287 (N_5287,N_2916,N_2289);
and U5288 (N_5288,N_1669,N_30);
or U5289 (N_5289,N_808,N_1479);
or U5290 (N_5290,N_2606,N_1833);
nor U5291 (N_5291,N_1226,N_2645);
and U5292 (N_5292,N_1870,N_1746);
nand U5293 (N_5293,N_2858,N_2082);
and U5294 (N_5294,N_838,N_620);
nand U5295 (N_5295,N_1248,N_818);
or U5296 (N_5296,N_1825,N_576);
or U5297 (N_5297,N_135,N_1115);
nor U5298 (N_5298,N_589,N_513);
or U5299 (N_5299,N_2482,N_1560);
nor U5300 (N_5300,N_1966,N_1688);
nand U5301 (N_5301,N_3137,N_3799);
or U5302 (N_5302,N_2229,N_3298);
nand U5303 (N_5303,N_1158,N_3261);
or U5304 (N_5304,N_2964,N_774);
or U5305 (N_5305,N_1249,N_2887);
nor U5306 (N_5306,N_1592,N_3056);
nor U5307 (N_5307,N_1338,N_1284);
nand U5308 (N_5308,N_430,N_3172);
nand U5309 (N_5309,N_3195,N_3466);
or U5310 (N_5310,N_83,N_2539);
nand U5311 (N_5311,N_2003,N_1340);
and U5312 (N_5312,N_845,N_3669);
and U5313 (N_5313,N_50,N_1128);
nand U5314 (N_5314,N_562,N_3679);
nand U5315 (N_5315,N_3561,N_276);
and U5316 (N_5316,N_1446,N_2966);
nand U5317 (N_5317,N_522,N_3483);
nor U5318 (N_5318,N_1381,N_2269);
or U5319 (N_5319,N_3518,N_1403);
or U5320 (N_5320,N_1394,N_2012);
nor U5321 (N_5321,N_309,N_71);
nand U5322 (N_5322,N_3625,N_2244);
or U5323 (N_5323,N_2836,N_3126);
nor U5324 (N_5324,N_3249,N_1134);
nor U5325 (N_5325,N_765,N_1845);
nor U5326 (N_5326,N_3917,N_2631);
nand U5327 (N_5327,N_374,N_2436);
nand U5328 (N_5328,N_288,N_3383);
nor U5329 (N_5329,N_2750,N_3305);
nand U5330 (N_5330,N_496,N_1578);
or U5331 (N_5331,N_390,N_1832);
nand U5332 (N_5332,N_3415,N_2597);
nor U5333 (N_5333,N_1136,N_884);
nor U5334 (N_5334,N_3100,N_857);
nor U5335 (N_5335,N_3646,N_2674);
xnor U5336 (N_5336,N_302,N_2838);
xnor U5337 (N_5337,N_1616,N_2640);
nor U5338 (N_5338,N_116,N_2426);
nor U5339 (N_5339,N_107,N_1094);
or U5340 (N_5340,N_2591,N_20);
xnor U5341 (N_5341,N_2488,N_199);
and U5342 (N_5342,N_1806,N_253);
and U5343 (N_5343,N_3902,N_2349);
and U5344 (N_5344,N_3845,N_688);
nand U5345 (N_5345,N_2184,N_1954);
and U5346 (N_5346,N_1410,N_1643);
nor U5347 (N_5347,N_1015,N_526);
and U5348 (N_5348,N_2702,N_656);
nor U5349 (N_5349,N_2500,N_1762);
nor U5350 (N_5350,N_1483,N_364);
xor U5351 (N_5351,N_741,N_320);
nor U5352 (N_5352,N_1079,N_1794);
xor U5353 (N_5353,N_2220,N_2231);
or U5354 (N_5354,N_3569,N_805);
or U5355 (N_5355,N_1330,N_3104);
and U5356 (N_5356,N_1099,N_105);
and U5357 (N_5357,N_3568,N_3888);
nand U5358 (N_5358,N_3738,N_1237);
and U5359 (N_5359,N_3776,N_885);
or U5360 (N_5360,N_1943,N_217);
nand U5361 (N_5361,N_2104,N_867);
nand U5362 (N_5362,N_2940,N_1674);
nor U5363 (N_5363,N_2806,N_2944);
or U5364 (N_5364,N_208,N_2601);
nand U5365 (N_5365,N_1039,N_1105);
nor U5366 (N_5366,N_2348,N_3396);
nand U5367 (N_5367,N_3140,N_3870);
and U5368 (N_5368,N_270,N_2444);
nor U5369 (N_5369,N_1864,N_3221);
nand U5370 (N_5370,N_721,N_2397);
or U5371 (N_5371,N_1916,N_3199);
and U5372 (N_5372,N_3089,N_450);
and U5373 (N_5373,N_1743,N_1608);
nor U5374 (N_5374,N_2852,N_1906);
or U5375 (N_5375,N_2549,N_1719);
or U5376 (N_5376,N_3434,N_3198);
xor U5377 (N_5377,N_655,N_1441);
and U5378 (N_5378,N_2169,N_955);
nor U5379 (N_5379,N_2846,N_3262);
or U5380 (N_5380,N_22,N_3353);
xor U5381 (N_5381,N_439,N_3697);
nor U5382 (N_5382,N_1129,N_1282);
and U5383 (N_5383,N_1266,N_2262);
and U5384 (N_5384,N_343,N_1964);
xnor U5385 (N_5385,N_237,N_825);
xor U5386 (N_5386,N_3031,N_3403);
and U5387 (N_5387,N_2556,N_1429);
or U5388 (N_5388,N_59,N_1725);
or U5389 (N_5389,N_956,N_926);
nand U5390 (N_5390,N_2316,N_2485);
or U5391 (N_5391,N_3626,N_919);
nand U5392 (N_5392,N_3890,N_2110);
nand U5393 (N_5393,N_3831,N_3887);
and U5394 (N_5394,N_1490,N_1520);
nor U5395 (N_5395,N_735,N_1298);
nor U5396 (N_5396,N_2534,N_3200);
nand U5397 (N_5397,N_3938,N_1436);
nor U5398 (N_5398,N_2907,N_978);
or U5399 (N_5399,N_2224,N_3425);
or U5400 (N_5400,N_215,N_2551);
or U5401 (N_5401,N_3904,N_1063);
or U5402 (N_5402,N_16,N_947);
nor U5403 (N_5403,N_251,N_1246);
nor U5404 (N_5404,N_1511,N_120);
or U5405 (N_5405,N_1034,N_1029);
or U5406 (N_5406,N_554,N_1469);
xnor U5407 (N_5407,N_914,N_3692);
and U5408 (N_5408,N_2560,N_63);
xnor U5409 (N_5409,N_1142,N_1618);
nand U5410 (N_5410,N_604,N_3896);
nor U5411 (N_5411,N_3526,N_1776);
or U5412 (N_5412,N_3355,N_716);
nand U5413 (N_5413,N_1717,N_3387);
and U5414 (N_5414,N_1234,N_3680);
nor U5415 (N_5415,N_1856,N_1482);
and U5416 (N_5416,N_1218,N_3503);
or U5417 (N_5417,N_1600,N_1716);
nand U5418 (N_5418,N_1579,N_2757);
and U5419 (N_5419,N_2965,N_301);
nor U5420 (N_5420,N_252,N_1286);
or U5421 (N_5421,N_1277,N_2529);
nand U5422 (N_5422,N_2775,N_368);
nand U5423 (N_5423,N_1961,N_2438);
or U5424 (N_5424,N_104,N_816);
and U5425 (N_5425,N_2311,N_2439);
xnor U5426 (N_5426,N_2306,N_1502);
nor U5427 (N_5427,N_2168,N_3608);
or U5428 (N_5428,N_3891,N_2245);
nand U5429 (N_5429,N_3416,N_3824);
nor U5430 (N_5430,N_471,N_3317);
nor U5431 (N_5431,N_1805,N_1349);
and U5432 (N_5432,N_1691,N_782);
xnor U5433 (N_5433,N_798,N_242);
or U5434 (N_5434,N_1639,N_2329);
nand U5435 (N_5435,N_2181,N_2876);
xnor U5436 (N_5436,N_2746,N_1827);
nor U5437 (N_5437,N_1093,N_3337);
or U5438 (N_5438,N_707,N_1598);
nand U5439 (N_5439,N_1767,N_962);
xor U5440 (N_5440,N_1077,N_12);
xor U5441 (N_5441,N_3370,N_565);
or U5442 (N_5442,N_2139,N_2827);
or U5443 (N_5443,N_995,N_2084);
or U5444 (N_5444,N_610,N_3176);
nand U5445 (N_5445,N_483,N_722);
and U5446 (N_5446,N_240,N_2015);
nand U5447 (N_5447,N_273,N_820);
or U5448 (N_5448,N_2004,N_2034);
nor U5449 (N_5449,N_2968,N_3966);
and U5450 (N_5450,N_1841,N_93);
nand U5451 (N_5451,N_3611,N_2328);
nand U5452 (N_5452,N_1920,N_2385);
or U5453 (N_5453,N_2629,N_1694);
or U5454 (N_5454,N_3720,N_3933);
and U5455 (N_5455,N_3096,N_3461);
nor U5456 (N_5456,N_911,N_1581);
xnor U5457 (N_5457,N_1422,N_1102);
nand U5458 (N_5458,N_3279,N_2670);
or U5459 (N_5459,N_2983,N_2815);
or U5460 (N_5460,N_2492,N_2520);
or U5461 (N_5461,N_2769,N_3851);
xnor U5462 (N_5462,N_2407,N_2962);
and U5463 (N_5463,N_2060,N_842);
nand U5464 (N_5464,N_2418,N_3443);
nor U5465 (N_5465,N_1798,N_2513);
and U5466 (N_5466,N_2627,N_2192);
nand U5467 (N_5467,N_792,N_1516);
nor U5468 (N_5468,N_3803,N_1817);
nor U5469 (N_5469,N_3747,N_2145);
and U5470 (N_5470,N_254,N_681);
nand U5471 (N_5471,N_2020,N_2843);
nor U5472 (N_5472,N_3676,N_2684);
xnor U5473 (N_5473,N_3598,N_3807);
nor U5474 (N_5474,N_2317,N_2772);
or U5475 (N_5475,N_2504,N_417);
nand U5476 (N_5476,N_1992,N_3770);
or U5477 (N_5477,N_1157,N_2951);
nand U5478 (N_5478,N_3072,N_2203);
nand U5479 (N_5479,N_863,N_2098);
and U5480 (N_5480,N_1571,N_1816);
nor U5481 (N_5481,N_841,N_1203);
nand U5482 (N_5482,N_1848,N_363);
or U5483 (N_5483,N_1971,N_1274);
nand U5484 (N_5484,N_3818,N_2900);
and U5485 (N_5485,N_1258,N_1426);
nor U5486 (N_5486,N_2305,N_3405);
or U5487 (N_5487,N_2803,N_1820);
nor U5488 (N_5488,N_2762,N_3672);
and U5489 (N_5489,N_3577,N_2603);
nor U5490 (N_5490,N_1677,N_1019);
or U5491 (N_5491,N_2011,N_936);
xor U5492 (N_5492,N_3923,N_788);
nor U5493 (N_5493,N_1514,N_3066);
nand U5494 (N_5494,N_3245,N_801);
nand U5495 (N_5495,N_44,N_2619);
and U5496 (N_5496,N_2373,N_1925);
or U5497 (N_5497,N_3601,N_456);
nor U5498 (N_5498,N_2498,N_1647);
or U5499 (N_5499,N_1591,N_3448);
nor U5500 (N_5500,N_2936,N_241);
nand U5501 (N_5501,N_879,N_3238);
nand U5502 (N_5502,N_272,N_3765);
nand U5503 (N_5503,N_457,N_2521);
nand U5504 (N_5504,N_1462,N_2904);
or U5505 (N_5505,N_1193,N_1449);
and U5506 (N_5506,N_3687,N_883);
nand U5507 (N_5507,N_943,N_1891);
nand U5508 (N_5508,N_561,N_224);
or U5509 (N_5509,N_2202,N_1775);
and U5510 (N_5510,N_1800,N_709);
and U5511 (N_5511,N_894,N_2297);
nand U5512 (N_5512,N_1455,N_2662);
nand U5513 (N_5513,N_2763,N_1826);
nor U5514 (N_5514,N_2128,N_2033);
nor U5515 (N_5515,N_1215,N_1651);
and U5516 (N_5516,N_3309,N_2740);
or U5517 (N_5517,N_2173,N_969);
or U5518 (N_5518,N_3419,N_3484);
or U5519 (N_5519,N_2995,N_1568);
and U5520 (N_5520,N_1281,N_28);
nor U5521 (N_5521,N_1873,N_1038);
and U5522 (N_5522,N_2421,N_3786);
and U5523 (N_5523,N_3609,N_3037);
nand U5524 (N_5524,N_1267,N_2017);
nand U5525 (N_5525,N_2527,N_2268);
nand U5526 (N_5526,N_3729,N_40);
nor U5527 (N_5527,N_2238,N_2875);
nor U5528 (N_5528,N_2831,N_223);
or U5529 (N_5529,N_2270,N_3742);
and U5530 (N_5530,N_1137,N_246);
nor U5531 (N_5531,N_1383,N_1602);
nand U5532 (N_5532,N_903,N_2476);
nand U5533 (N_5533,N_3939,N_3940);
nand U5534 (N_5534,N_1146,N_1701);
nand U5535 (N_5535,N_2442,N_830);
xor U5536 (N_5536,N_406,N_1631);
nor U5537 (N_5537,N_2515,N_539);
nand U5538 (N_5538,N_3161,N_3006);
or U5539 (N_5539,N_117,N_1804);
and U5540 (N_5540,N_3622,N_2478);
and U5541 (N_5541,N_1542,N_752);
or U5542 (N_5542,N_165,N_2200);
or U5543 (N_5543,N_3947,N_334);
nor U5544 (N_5544,N_3773,N_1241);
and U5545 (N_5545,N_111,N_210);
and U5546 (N_5546,N_3077,N_130);
xnor U5547 (N_5547,N_256,N_1540);
nor U5548 (N_5548,N_2392,N_3216);
nor U5549 (N_5549,N_3642,N_2115);
or U5550 (N_5550,N_188,N_235);
nand U5551 (N_5551,N_2183,N_1613);
nand U5552 (N_5552,N_1356,N_942);
nor U5553 (N_5553,N_1895,N_156);
or U5554 (N_5554,N_2242,N_3233);
and U5555 (N_5555,N_3048,N_2036);
nor U5556 (N_5556,N_3052,N_2816);
or U5557 (N_5557,N_2614,N_529);
xnor U5558 (N_5558,N_1299,N_1791);
or U5559 (N_5559,N_2577,N_3965);
nor U5560 (N_5560,N_2809,N_736);
nor U5561 (N_5561,N_26,N_2817);
nor U5562 (N_5562,N_2886,N_2667);
nand U5563 (N_5563,N_2882,N_609);
or U5564 (N_5564,N_142,N_2147);
and U5565 (N_5565,N_3299,N_1508);
and U5566 (N_5566,N_454,N_938);
or U5567 (N_5567,N_1995,N_127);
nor U5568 (N_5568,N_2069,N_1802);
or U5569 (N_5569,N_2952,N_2927);
and U5570 (N_5570,N_3592,N_3911);
xor U5571 (N_5571,N_1795,N_1049);
or U5572 (N_5572,N_2576,N_2078);
and U5573 (N_5573,N_2441,N_720);
nor U5574 (N_5574,N_1997,N_2256);
or U5575 (N_5575,N_3032,N_1405);
nand U5576 (N_5576,N_3927,N_2199);
or U5577 (N_5577,N_1228,N_3825);
and U5578 (N_5578,N_395,N_2590);
nor U5579 (N_5579,N_2137,N_639);
xor U5580 (N_5580,N_3912,N_124);
nand U5581 (N_5581,N_158,N_3572);
nand U5582 (N_5582,N_473,N_1318);
or U5583 (N_5583,N_45,N_216);
xor U5584 (N_5584,N_3110,N_3220);
and U5585 (N_5585,N_2105,N_988);
and U5586 (N_5586,N_175,N_1982);
or U5587 (N_5587,N_1710,N_332);
and U5588 (N_5588,N_2728,N_813);
or U5589 (N_5589,N_965,N_3319);
xnor U5590 (N_5590,N_1488,N_3603);
or U5591 (N_5591,N_3996,N_1881);
nand U5592 (N_5592,N_1771,N_3124);
nor U5593 (N_5593,N_585,N_1051);
nand U5594 (N_5594,N_992,N_311);
or U5595 (N_5595,N_1934,N_1926);
and U5596 (N_5596,N_2353,N_2660);
nor U5597 (N_5597,N_1162,N_1445);
nor U5598 (N_5598,N_1533,N_1588);
nor U5599 (N_5599,N_1739,N_2193);
nor U5600 (N_5600,N_3695,N_2312);
and U5601 (N_5601,N_3685,N_1202);
xnor U5602 (N_5602,N_998,N_1509);
and U5603 (N_5603,N_3361,N_954);
nor U5604 (N_5604,N_1053,N_1851);
nor U5605 (N_5605,N_1458,N_3955);
nor U5606 (N_5606,N_1537,N_2971);
nor U5607 (N_5607,N_3101,N_495);
or U5608 (N_5608,N_1044,N_82);
or U5609 (N_5609,N_436,N_3050);
nand U5610 (N_5610,N_3978,N_1473);
or U5611 (N_5611,N_1268,N_2340);
nand U5612 (N_5612,N_1339,N_2463);
or U5613 (N_5613,N_1889,N_1398);
or U5614 (N_5614,N_184,N_1822);
and U5615 (N_5615,N_3307,N_3708);
or U5616 (N_5616,N_2065,N_2403);
and U5617 (N_5617,N_475,N_1735);
or U5618 (N_5618,N_3083,N_2457);
nor U5619 (N_5619,N_3867,N_822);
or U5620 (N_5620,N_2050,N_1186);
or U5621 (N_5621,N_434,N_25);
and U5622 (N_5622,N_193,N_2142);
nor U5623 (N_5623,N_3534,N_3861);
nor U5624 (N_5624,N_1135,N_2251);
or U5625 (N_5625,N_1732,N_1854);
or U5626 (N_5626,N_3259,N_1774);
nor U5627 (N_5627,N_1336,N_2201);
and U5628 (N_5628,N_155,N_3257);
xor U5629 (N_5629,N_2424,N_933);
nand U5630 (N_5630,N_3633,N_2825);
nand U5631 (N_5631,N_2483,N_3713);
and U5632 (N_5632,N_3693,N_1853);
or U5633 (N_5633,N_3085,N_1052);
or U5634 (N_5634,N_3411,N_832);
and U5635 (N_5635,N_3942,N_2977);
xnor U5636 (N_5636,N_837,N_3994);
nor U5637 (N_5637,N_3631,N_2531);
nand U5638 (N_5638,N_588,N_668);
nand U5639 (N_5639,N_2109,N_106);
and U5640 (N_5640,N_1200,N_2707);
or U5641 (N_5641,N_605,N_2447);
nand U5642 (N_5642,N_3482,N_3524);
or U5643 (N_5643,N_39,N_2617);
nand U5644 (N_5644,N_1519,N_3283);
or U5645 (N_5645,N_1343,N_1244);
nand U5646 (N_5646,N_3990,N_747);
nand U5647 (N_5647,N_2240,N_3028);
nor U5648 (N_5648,N_555,N_3949);
or U5649 (N_5649,N_2085,N_1423);
nor U5650 (N_5650,N_1089,N_3730);
and U5651 (N_5651,N_2518,N_776);
nor U5652 (N_5652,N_2947,N_2593);
and U5653 (N_5653,N_621,N_3446);
and U5654 (N_5654,N_1857,N_1119);
and U5655 (N_5655,N_3401,N_2994);
nand U5656 (N_5656,N_3979,N_2227);
and U5657 (N_5657,N_409,N_803);
and U5658 (N_5658,N_3242,N_3217);
or U5659 (N_5659,N_1127,N_1057);
nor U5660 (N_5660,N_644,N_3035);
or U5661 (N_5661,N_2263,N_3848);
or U5662 (N_5662,N_2921,N_3684);
xnor U5663 (N_5663,N_3809,N_3910);
and U5664 (N_5664,N_157,N_3704);
and U5665 (N_5665,N_3981,N_3591);
or U5666 (N_5666,N_2117,N_3440);
or U5667 (N_5667,N_3206,N_2290);
or U5668 (N_5668,N_2437,N_2671);
and U5669 (N_5669,N_467,N_148);
nor U5670 (N_5670,N_1332,N_930);
nand U5671 (N_5671,N_9,N_1641);
and U5672 (N_5672,N_1196,N_1320);
nand U5673 (N_5673,N_3120,N_2984);
xnor U5674 (N_5674,N_2717,N_3306);
nand U5675 (N_5675,N_2848,N_3398);
and U5676 (N_5676,N_1225,N_3218);
nand U5677 (N_5677,N_3652,N_2961);
nor U5678 (N_5678,N_3107,N_1465);
nand U5679 (N_5679,N_3366,N_49);
nor U5680 (N_5680,N_827,N_1682);
or U5681 (N_5681,N_1958,N_3119);
nand U5682 (N_5682,N_1380,N_2950);
nand U5683 (N_5683,N_314,N_2997);
or U5684 (N_5684,N_2368,N_293);
and U5685 (N_5685,N_3739,N_921);
or U5686 (N_5686,N_3620,N_523);
or U5687 (N_5687,N_2214,N_385);
nand U5688 (N_5688,N_3044,N_3197);
and U5689 (N_5689,N_3094,N_2695);
nand U5690 (N_5690,N_1316,N_2683);
or U5691 (N_5691,N_3042,N_2715);
xor U5692 (N_5692,N_1369,N_1141);
nand U5693 (N_5693,N_2093,N_1939);
nand U5694 (N_5694,N_525,N_870);
nand U5695 (N_5695,N_379,N_3352);
nor U5696 (N_5696,N_192,N_3663);
nand U5697 (N_5697,N_3268,N_2546);
or U5698 (N_5698,N_2553,N_3260);
or U5699 (N_5699,N_3565,N_2364);
nand U5700 (N_5700,N_3002,N_2467);
or U5701 (N_5701,N_238,N_2582);
nor U5702 (N_5702,N_228,N_3296);
nor U5703 (N_5703,N_3231,N_1707);
nand U5704 (N_5704,N_643,N_899);
nand U5705 (N_5705,N_1686,N_3878);
nor U5706 (N_5706,N_1173,N_2462);
nor U5707 (N_5707,N_2575,N_2735);
xor U5708 (N_5708,N_1989,N_1496);
or U5709 (N_5709,N_3276,N_858);
nor U5710 (N_5710,N_996,N_2350);
nand U5711 (N_5711,N_1150,N_3859);
xnor U5712 (N_5712,N_3787,N_2819);
nor U5713 (N_5713,N_87,N_1747);
nor U5714 (N_5714,N_1315,N_1240);
nor U5715 (N_5715,N_2296,N_907);
nor U5716 (N_5716,N_1991,N_2885);
or U5717 (N_5717,N_730,N_1836);
nor U5718 (N_5718,N_626,N_1216);
nand U5719 (N_5719,N_1702,N_3288);
and U5720 (N_5720,N_3491,N_1902);
or U5721 (N_5721,N_2396,N_619);
nor U5722 (N_5722,N_946,N_2126);
and U5723 (N_5723,N_3080,N_2298);
xnor U5724 (N_5724,N_2778,N_35);
and U5725 (N_5725,N_491,N_3805);
or U5726 (N_5726,N_1148,N_1060);
and U5727 (N_5727,N_3315,N_145);
xnor U5728 (N_5728,N_821,N_2094);
nand U5729 (N_5729,N_1566,N_2788);
and U5730 (N_5730,N_3688,N_1361);
or U5731 (N_5731,N_1976,N_3102);
nor U5732 (N_5732,N_405,N_3477);
xnor U5733 (N_5733,N_875,N_1321);
or U5734 (N_5734,N_2731,N_2253);
or U5735 (N_5735,N_1704,N_2361);
nor U5736 (N_5736,N_2377,N_163);
or U5737 (N_5737,N_2985,N_3436);
nand U5738 (N_5738,N_783,N_3219);
or U5739 (N_5739,N_3289,N_1680);
or U5740 (N_5740,N_3164,N_486);
and U5741 (N_5741,N_119,N_1899);
and U5742 (N_5742,N_321,N_1497);
nand U5743 (N_5743,N_1532,N_2237);
nand U5744 (N_5744,N_1205,N_3075);
or U5745 (N_5745,N_2562,N_2165);
nand U5746 (N_5746,N_1116,N_3156);
and U5747 (N_5747,N_1524,N_2957);
nand U5748 (N_5748,N_2469,N_3722);
or U5749 (N_5749,N_1898,N_501);
nand U5750 (N_5750,N_3057,N_2925);
or U5751 (N_5751,N_2278,N_3817);
or U5752 (N_5752,N_3914,N_1307);
xor U5753 (N_5753,N_1543,N_1037);
and U5754 (N_5754,N_3907,N_3015);
nor U5755 (N_5755,N_1032,N_3512);
or U5756 (N_5756,N_3450,N_3689);
and U5757 (N_5757,N_2122,N_112);
xnor U5758 (N_5758,N_3321,N_600);
and U5759 (N_5759,N_3763,N_2554);
nor U5760 (N_5760,N_7,N_2257);
and U5761 (N_5761,N_2318,N_67);
and U5762 (N_5762,N_2844,N_994);
nor U5763 (N_5763,N_1217,N_2781);
xor U5764 (N_5764,N_1535,N_1622);
nand U5765 (N_5765,N_3005,N_2216);
nand U5766 (N_5766,N_3639,N_76);
nor U5767 (N_5767,N_1182,N_3185);
nor U5768 (N_5768,N_3908,N_1887);
or U5769 (N_5769,N_2871,N_1922);
nor U5770 (N_5770,N_1623,N_2679);
or U5771 (N_5771,N_3373,N_677);
or U5772 (N_5772,N_2063,N_2380);
or U5773 (N_5773,N_1189,N_3414);
xnor U5774 (N_5774,N_3369,N_151);
nor U5775 (N_5775,N_1293,N_3789);
or U5776 (N_5776,N_3391,N_2805);
or U5777 (N_5777,N_2293,N_3879);
nand U5778 (N_5778,N_3211,N_3918);
xor U5779 (N_5779,N_1777,N_3989);
or U5780 (N_5780,N_1709,N_2867);
xor U5781 (N_5781,N_1461,N_2834);
nor U5782 (N_5782,N_3774,N_444);
nand U5783 (N_5783,N_1572,N_3517);
and U5784 (N_5784,N_901,N_3376);
and U5785 (N_5785,N_2635,N_635);
and U5786 (N_5786,N_1536,N_452);
xnor U5787 (N_5787,N_403,N_52);
and U5788 (N_5788,N_2198,N_1850);
nor U5789 (N_5789,N_3115,N_2758);
nor U5790 (N_5790,N_3243,N_2744);
nand U5791 (N_5791,N_1404,N_1420);
or U5792 (N_5792,N_2796,N_3833);
nand U5793 (N_5793,N_2167,N_1736);
or U5794 (N_5794,N_2664,N_642);
or U5795 (N_5795,N_72,N_2232);
nand U5796 (N_5796,N_2187,N_411);
nor U5797 (N_5797,N_546,N_665);
and U5798 (N_5798,N_2748,N_365);
xnor U5799 (N_5799,N_3778,N_1151);
nand U5800 (N_5800,N_169,N_3850);
nor U5801 (N_5801,N_2235,N_3253);
and U5802 (N_5802,N_1144,N_367);
and U5803 (N_5803,N_1624,N_1693);
and U5804 (N_5804,N_3528,N_3418);
nand U5805 (N_5805,N_1700,N_1362);
and U5806 (N_5806,N_2727,N_2650);
and U5807 (N_5807,N_3580,N_2170);
or U5808 (N_5808,N_1371,N_218);
xnor U5809 (N_5809,N_2443,N_1255);
and U5810 (N_5810,N_3270,N_1890);
xor U5811 (N_5811,N_2566,N_667);
or U5812 (N_5812,N_3948,N_492);
and U5813 (N_5813,N_2320,N_1905);
or U5814 (N_5814,N_203,N_3547);
or U5815 (N_5815,N_1353,N_1831);
nand U5816 (N_5816,N_2140,N_197);
or U5817 (N_5817,N_1288,N_1527);
nor U5818 (N_5818,N_351,N_3843);
or U5819 (N_5819,N_3108,N_2611);
or U5820 (N_5820,N_1783,N_3047);
nor U5821 (N_5821,N_3880,N_3976);
xor U5822 (N_5822,N_2934,N_2799);
nand U5823 (N_5823,N_1324,N_1036);
nand U5824 (N_5824,N_2567,N_2558);
nand U5825 (N_5825,N_3883,N_2693);
nand U5826 (N_5826,N_3798,N_3397);
xor U5827 (N_5827,N_3762,N_2960);
and U5828 (N_5828,N_2742,N_833);
and U5829 (N_5829,N_1048,N_47);
nand U5830 (N_5830,N_2295,N_2148);
or U5831 (N_5831,N_1577,N_3087);
nand U5832 (N_5832,N_1167,N_1754);
and U5833 (N_5833,N_3502,N_1814);
xnor U5834 (N_5834,N_510,N_2030);
and U5835 (N_5835,N_560,N_3024);
and U5836 (N_5836,N_377,N_1668);
nor U5837 (N_5837,N_3359,N_1846);
nand U5838 (N_5838,N_3430,N_2710);
or U5839 (N_5839,N_1184,N_75);
nor U5840 (N_5840,N_3758,N_553);
nor U5841 (N_5841,N_3567,N_2077);
and U5842 (N_5842,N_227,N_3480);
nor U5843 (N_5843,N_3982,N_1100);
nand U5844 (N_5844,N_113,N_622);
nor U5845 (N_5845,N_247,N_785);
and U5846 (N_5846,N_2484,N_3544);
or U5847 (N_5847,N_3163,N_2146);
nand U5848 (N_5848,N_205,N_154);
nand U5849 (N_5849,N_2300,N_2564);
and U5850 (N_5850,N_2651,N_790);
nand U5851 (N_5851,N_200,N_489);
nand U5852 (N_5852,N_1378,N_3647);
nor U5853 (N_5853,N_455,N_3423);
nand U5854 (N_5854,N_3992,N_1472);
and U5855 (N_5855,N_1894,N_676);
nor U5856 (N_5856,N_2189,N_3666);
nor U5857 (N_5857,N_3487,N_1442);
nor U5858 (N_5858,N_1525,N_3158);
nand U5859 (N_5859,N_3854,N_1558);
nand U5860 (N_5860,N_935,N_2970);
or U5861 (N_5861,N_1285,N_950);
nor U5862 (N_5862,N_2792,N_1071);
nand U5863 (N_5863,N_1782,N_1652);
or U5864 (N_5864,N_414,N_3920);
nor U5865 (N_5865,N_2402,N_1741);
xor U5866 (N_5866,N_1757,N_3551);
and U5867 (N_5867,N_2938,N_278);
or U5868 (N_5868,N_3804,N_2797);
nand U5869 (N_5869,N_2414,N_187);
or U5870 (N_5870,N_3821,N_2499);
nand U5871 (N_5871,N_3091,N_1080);
and U5872 (N_5872,N_754,N_3093);
and U5873 (N_5873,N_2477,N_3606);
nand U5874 (N_5874,N_3266,N_3062);
and U5875 (N_5875,N_226,N_1720);
xor U5876 (N_5876,N_521,N_2514);
or U5877 (N_5877,N_292,N_530);
nor U5878 (N_5878,N_2979,N_1612);
or U5879 (N_5879,N_1239,N_2874);
nand U5880 (N_5880,N_2014,N_2880);
nor U5881 (N_5881,N_1302,N_2374);
or U5882 (N_5882,N_2212,N_391);
or U5883 (N_5883,N_2405,N_742);
nand U5884 (N_5884,N_1938,N_1008);
nor U5885 (N_5885,N_3125,N_990);
and U5886 (N_5886,N_1972,N_3349);
nand U5887 (N_5887,N_2922,N_1346);
nor U5888 (N_5888,N_229,N_648);
nand U5889 (N_5889,N_2780,N_1448);
xor U5890 (N_5890,N_2541,N_17);
and U5891 (N_5891,N_3496,N_3000);
nor U5892 (N_5892,N_2343,N_1684);
and U5893 (N_5893,N_535,N_3872);
and U5894 (N_5894,N_2049,N_304);
nand U5895 (N_5895,N_10,N_2494);
nand U5896 (N_5896,N_1970,N_2339);
and U5897 (N_5897,N_3605,N_1615);
or U5898 (N_5898,N_880,N_3819);
xnor U5899 (N_5899,N_2359,N_2811);
or U5900 (N_5900,N_2079,N_2956);
xor U5901 (N_5901,N_566,N_3785);
nand U5902 (N_5902,N_3027,N_1170);
nor U5903 (N_5903,N_3876,N_675);
nand U5904 (N_5904,N_1166,N_383);
and U5905 (N_5905,N_1126,N_394);
and U5906 (N_5906,N_3420,N_552);
and U5907 (N_5907,N_283,N_24);
and U5908 (N_5908,N_2241,N_1130);
nand U5909 (N_5909,N_567,N_1392);
xor U5910 (N_5910,N_312,N_3363);
and U5911 (N_5911,N_3624,N_3743);
nor U5912 (N_5912,N_1035,N_2440);
or U5913 (N_5913,N_802,N_3521);
or U5914 (N_5914,N_3836,N_1784);
nor U5915 (N_5915,N_743,N_280);
or U5916 (N_5916,N_1192,N_3969);
or U5917 (N_5917,N_905,N_2866);
nor U5918 (N_5918,N_1168,N_836);
nor U5919 (N_5919,N_1584,N_1074);
nor U5920 (N_5920,N_1149,N_893);
nand U5921 (N_5921,N_422,N_2686);
nor U5922 (N_5922,N_1335,N_758);
and U5923 (N_5923,N_1843,N_2016);
and U5924 (N_5924,N_2905,N_3925);
xor U5925 (N_5925,N_1139,N_1352);
nand U5926 (N_5926,N_2881,N_21);
or U5927 (N_5927,N_963,N_3581);
nor U5928 (N_5928,N_1096,N_633);
nand U5929 (N_5929,N_2338,N_1633);
xnor U5930 (N_5930,N_615,N_1614);
xnor U5931 (N_5931,N_1689,N_2745);
nand U5932 (N_5932,N_3392,N_925);
or U5933 (N_5933,N_61,N_3314);
nor U5934 (N_5934,N_624,N_2021);
xor U5935 (N_5935,N_1487,N_3866);
nor U5936 (N_5936,N_3894,N_579);
and U5937 (N_5937,N_960,N_258);
or U5938 (N_5938,N_1953,N_2711);
or U5939 (N_5939,N_1779,N_1444);
nand U5940 (N_5940,N_2027,N_2366);
nand U5941 (N_5941,N_1327,N_2768);
nand U5942 (N_5942,N_259,N_2545);
and U5943 (N_5943,N_3025,N_2636);
nor U5944 (N_5944,N_1190,N_1522);
or U5945 (N_5945,N_3166,N_484);
or U5946 (N_5946,N_3302,N_420);
nor U5947 (N_5947,N_3248,N_1447);
xor U5948 (N_5948,N_97,N_249);
xnor U5949 (N_5949,N_778,N_3269);
or U5950 (N_5950,N_1974,N_2986);
and U5951 (N_5951,N_997,N_494);
nand U5952 (N_5952,N_1987,N_512);
nor U5953 (N_5953,N_1430,N_3003);
or U5954 (N_5954,N_2429,N_1760);
nor U5955 (N_5955,N_3853,N_3527);
xnor U5956 (N_5956,N_1155,N_1562);
and U5957 (N_5957,N_177,N_2613);
nor U5958 (N_5958,N_2510,N_1662);
nor U5959 (N_5959,N_8,N_34);
nand U5960 (N_5960,N_1366,N_746);
or U5961 (N_5961,N_796,N_1084);
xor U5962 (N_5962,N_932,N_3287);
nand U5963 (N_5963,N_1801,N_1486);
nor U5964 (N_5964,N_3017,N_3659);
or U5965 (N_5965,N_1665,N_2893);
and U5966 (N_5966,N_2761,N_1347);
nand U5967 (N_5967,N_2706,N_634);
nand U5968 (N_5968,N_353,N_1998);
xnor U5969 (N_5969,N_463,N_861);
nand U5970 (N_5970,N_115,N_3263);
and U5971 (N_5971,N_3293,N_1770);
nand U5972 (N_5972,N_2522,N_3012);
and U5973 (N_5973,N_3667,N_3284);
and U5974 (N_5974,N_1357,N_2540);
xnor U5975 (N_5975,N_3828,N_2042);
nor U5976 (N_5976,N_3356,N_1367);
and U5977 (N_5977,N_2131,N_3842);
or U5978 (N_5978,N_88,N_2538);
or U5979 (N_5979,N_2869,N_1344);
nor U5980 (N_5980,N_0,N_2915);
or U5981 (N_5981,N_3915,N_2382);
and U5982 (N_5982,N_3386,N_1780);
nand U5983 (N_5983,N_322,N_3264);
xnor U5984 (N_5984,N_3886,N_974);
and U5985 (N_5985,N_3304,N_1223);
and U5986 (N_5986,N_358,N_3492);
and U5987 (N_5987,N_2387,N_338);
or U5988 (N_5988,N_2810,N_1658);
nand U5989 (N_5989,N_2802,N_3644);
nand U5990 (N_5990,N_1494,N_189);
and U5991 (N_5991,N_2275,N_3650);
and U5992 (N_5992,N_2274,N_1097);
and U5993 (N_5993,N_3794,N_225);
xnor U5994 (N_5994,N_448,N_2481);
nand U5995 (N_5995,N_638,N_2333);
and U5996 (N_5996,N_1901,N_2779);
or U5997 (N_5997,N_3868,N_3511);
and U5998 (N_5998,N_3640,N_360);
or U5999 (N_5999,N_3375,N_3424);
nand U6000 (N_6000,N_2345,N_84);
nand U6001 (N_6001,N_309,N_2378);
or U6002 (N_6002,N_802,N_1750);
and U6003 (N_6003,N_407,N_2506);
nand U6004 (N_6004,N_2533,N_3494);
or U6005 (N_6005,N_634,N_3184);
or U6006 (N_6006,N_2211,N_1098);
or U6007 (N_6007,N_1155,N_1448);
nand U6008 (N_6008,N_252,N_736);
or U6009 (N_6009,N_2481,N_2905);
or U6010 (N_6010,N_3439,N_2771);
or U6011 (N_6011,N_2224,N_2400);
and U6012 (N_6012,N_2150,N_1531);
and U6013 (N_6013,N_761,N_1006);
or U6014 (N_6014,N_2382,N_29);
nand U6015 (N_6015,N_1464,N_905);
nand U6016 (N_6016,N_3899,N_2789);
or U6017 (N_6017,N_3890,N_2234);
and U6018 (N_6018,N_174,N_2463);
nand U6019 (N_6019,N_1922,N_3349);
and U6020 (N_6020,N_2935,N_1070);
nand U6021 (N_6021,N_2391,N_120);
nor U6022 (N_6022,N_215,N_2197);
or U6023 (N_6023,N_1857,N_1893);
or U6024 (N_6024,N_1268,N_3858);
and U6025 (N_6025,N_2101,N_2738);
and U6026 (N_6026,N_180,N_2169);
and U6027 (N_6027,N_2499,N_702);
nor U6028 (N_6028,N_3539,N_800);
and U6029 (N_6029,N_3499,N_344);
nand U6030 (N_6030,N_3046,N_304);
and U6031 (N_6031,N_2010,N_1359);
nand U6032 (N_6032,N_2024,N_2795);
or U6033 (N_6033,N_325,N_2387);
and U6034 (N_6034,N_1572,N_2986);
or U6035 (N_6035,N_1142,N_3110);
or U6036 (N_6036,N_1144,N_2206);
or U6037 (N_6037,N_2034,N_1286);
nand U6038 (N_6038,N_3935,N_912);
xnor U6039 (N_6039,N_629,N_2720);
or U6040 (N_6040,N_1,N_1388);
or U6041 (N_6041,N_1986,N_488);
nor U6042 (N_6042,N_3032,N_3620);
nand U6043 (N_6043,N_3607,N_721);
or U6044 (N_6044,N_1580,N_390);
nand U6045 (N_6045,N_2915,N_3834);
nand U6046 (N_6046,N_1625,N_3231);
xor U6047 (N_6047,N_1936,N_301);
and U6048 (N_6048,N_1611,N_3913);
nand U6049 (N_6049,N_3899,N_2904);
nand U6050 (N_6050,N_1228,N_2728);
or U6051 (N_6051,N_3562,N_2149);
nor U6052 (N_6052,N_3408,N_641);
and U6053 (N_6053,N_3061,N_3960);
or U6054 (N_6054,N_904,N_2177);
nand U6055 (N_6055,N_3328,N_3378);
or U6056 (N_6056,N_2797,N_2);
xnor U6057 (N_6057,N_2781,N_425);
nand U6058 (N_6058,N_369,N_815);
nor U6059 (N_6059,N_3509,N_2733);
and U6060 (N_6060,N_648,N_3773);
nand U6061 (N_6061,N_469,N_1055);
or U6062 (N_6062,N_1895,N_3901);
and U6063 (N_6063,N_3200,N_2555);
and U6064 (N_6064,N_2039,N_1257);
or U6065 (N_6065,N_3234,N_1194);
or U6066 (N_6066,N_2705,N_2917);
nand U6067 (N_6067,N_686,N_2857);
nand U6068 (N_6068,N_3489,N_500);
and U6069 (N_6069,N_3720,N_600);
and U6070 (N_6070,N_3522,N_1129);
and U6071 (N_6071,N_279,N_3605);
and U6072 (N_6072,N_3699,N_997);
or U6073 (N_6073,N_1200,N_2209);
nand U6074 (N_6074,N_2835,N_3893);
nand U6075 (N_6075,N_2593,N_1578);
nor U6076 (N_6076,N_3998,N_3296);
nand U6077 (N_6077,N_3686,N_1500);
nand U6078 (N_6078,N_2396,N_3400);
xnor U6079 (N_6079,N_2520,N_693);
or U6080 (N_6080,N_108,N_2428);
nor U6081 (N_6081,N_3791,N_306);
xor U6082 (N_6082,N_2319,N_2023);
xor U6083 (N_6083,N_654,N_1239);
and U6084 (N_6084,N_2157,N_689);
or U6085 (N_6085,N_345,N_2532);
and U6086 (N_6086,N_2785,N_1563);
and U6087 (N_6087,N_2701,N_3862);
or U6088 (N_6088,N_3769,N_3739);
nor U6089 (N_6089,N_2614,N_584);
xnor U6090 (N_6090,N_2523,N_1210);
or U6091 (N_6091,N_3518,N_1780);
nand U6092 (N_6092,N_201,N_2968);
nand U6093 (N_6093,N_722,N_2340);
nor U6094 (N_6094,N_150,N_3578);
nand U6095 (N_6095,N_2035,N_1415);
nor U6096 (N_6096,N_2433,N_1224);
and U6097 (N_6097,N_2096,N_2915);
nand U6098 (N_6098,N_774,N_979);
or U6099 (N_6099,N_3227,N_140);
nor U6100 (N_6100,N_467,N_3867);
or U6101 (N_6101,N_2036,N_1606);
nand U6102 (N_6102,N_1264,N_2850);
or U6103 (N_6103,N_3768,N_749);
nand U6104 (N_6104,N_1111,N_924);
nor U6105 (N_6105,N_1468,N_3574);
and U6106 (N_6106,N_3357,N_3150);
nand U6107 (N_6107,N_2524,N_2885);
nand U6108 (N_6108,N_2433,N_2513);
and U6109 (N_6109,N_3386,N_743);
nand U6110 (N_6110,N_2224,N_3545);
nand U6111 (N_6111,N_1647,N_1687);
xnor U6112 (N_6112,N_3178,N_2064);
nand U6113 (N_6113,N_3473,N_2565);
nor U6114 (N_6114,N_1839,N_2666);
nand U6115 (N_6115,N_2423,N_2097);
nor U6116 (N_6116,N_2203,N_906);
nor U6117 (N_6117,N_3443,N_2731);
and U6118 (N_6118,N_210,N_1723);
and U6119 (N_6119,N_672,N_2591);
nor U6120 (N_6120,N_573,N_2037);
nor U6121 (N_6121,N_3847,N_550);
and U6122 (N_6122,N_1725,N_1086);
nand U6123 (N_6123,N_2226,N_2373);
nor U6124 (N_6124,N_270,N_64);
nor U6125 (N_6125,N_67,N_2640);
nor U6126 (N_6126,N_707,N_134);
or U6127 (N_6127,N_527,N_136);
nor U6128 (N_6128,N_750,N_529);
nand U6129 (N_6129,N_2222,N_2895);
nand U6130 (N_6130,N_1742,N_3785);
and U6131 (N_6131,N_1610,N_973);
xor U6132 (N_6132,N_623,N_1702);
nand U6133 (N_6133,N_2510,N_2440);
xor U6134 (N_6134,N_3350,N_3425);
nand U6135 (N_6135,N_1764,N_1991);
nor U6136 (N_6136,N_753,N_1562);
nor U6137 (N_6137,N_3660,N_992);
and U6138 (N_6138,N_1613,N_96);
nor U6139 (N_6139,N_3243,N_3458);
nor U6140 (N_6140,N_1364,N_3555);
nand U6141 (N_6141,N_1530,N_779);
or U6142 (N_6142,N_1305,N_3034);
and U6143 (N_6143,N_892,N_594);
and U6144 (N_6144,N_3477,N_1546);
xor U6145 (N_6145,N_542,N_449);
and U6146 (N_6146,N_3411,N_1087);
nor U6147 (N_6147,N_2730,N_182);
nor U6148 (N_6148,N_1963,N_1508);
and U6149 (N_6149,N_3262,N_3578);
or U6150 (N_6150,N_3986,N_935);
nor U6151 (N_6151,N_1856,N_433);
or U6152 (N_6152,N_2974,N_1212);
nor U6153 (N_6153,N_2703,N_2426);
xnor U6154 (N_6154,N_1741,N_3182);
xor U6155 (N_6155,N_531,N_1748);
and U6156 (N_6156,N_2333,N_537);
xnor U6157 (N_6157,N_1899,N_24);
or U6158 (N_6158,N_3742,N_1137);
and U6159 (N_6159,N_2162,N_95);
and U6160 (N_6160,N_3347,N_3584);
nor U6161 (N_6161,N_785,N_1959);
nor U6162 (N_6162,N_2447,N_2509);
or U6163 (N_6163,N_2242,N_1527);
nor U6164 (N_6164,N_727,N_1356);
nor U6165 (N_6165,N_719,N_1890);
and U6166 (N_6166,N_3125,N_3986);
and U6167 (N_6167,N_2847,N_2989);
and U6168 (N_6168,N_2176,N_3501);
nand U6169 (N_6169,N_1756,N_2586);
nand U6170 (N_6170,N_225,N_531);
xnor U6171 (N_6171,N_2929,N_150);
nor U6172 (N_6172,N_33,N_3272);
and U6173 (N_6173,N_2424,N_1937);
nand U6174 (N_6174,N_1089,N_3676);
or U6175 (N_6175,N_793,N_487);
xor U6176 (N_6176,N_1845,N_3352);
xor U6177 (N_6177,N_493,N_2799);
nor U6178 (N_6178,N_344,N_1493);
nand U6179 (N_6179,N_138,N_3189);
nand U6180 (N_6180,N_3636,N_183);
xnor U6181 (N_6181,N_2157,N_526);
xnor U6182 (N_6182,N_1860,N_3537);
and U6183 (N_6183,N_2630,N_3391);
nand U6184 (N_6184,N_206,N_156);
nor U6185 (N_6185,N_447,N_3369);
and U6186 (N_6186,N_2852,N_3156);
or U6187 (N_6187,N_73,N_2659);
xnor U6188 (N_6188,N_2469,N_3820);
nor U6189 (N_6189,N_3792,N_1027);
nand U6190 (N_6190,N_483,N_1252);
nand U6191 (N_6191,N_3227,N_2230);
or U6192 (N_6192,N_1580,N_2737);
and U6193 (N_6193,N_3963,N_1428);
or U6194 (N_6194,N_3133,N_198);
xnor U6195 (N_6195,N_2718,N_1982);
nor U6196 (N_6196,N_946,N_254);
nand U6197 (N_6197,N_3666,N_1198);
nor U6198 (N_6198,N_3192,N_2289);
nand U6199 (N_6199,N_3955,N_1994);
xnor U6200 (N_6200,N_1851,N_1955);
nor U6201 (N_6201,N_3373,N_2388);
nand U6202 (N_6202,N_2088,N_575);
and U6203 (N_6203,N_2682,N_311);
nand U6204 (N_6204,N_1920,N_1214);
nand U6205 (N_6205,N_695,N_1743);
nor U6206 (N_6206,N_824,N_3710);
or U6207 (N_6207,N_12,N_1590);
nor U6208 (N_6208,N_2359,N_425);
nand U6209 (N_6209,N_2147,N_1909);
nor U6210 (N_6210,N_3823,N_2749);
nor U6211 (N_6211,N_3395,N_1583);
and U6212 (N_6212,N_2938,N_2893);
nor U6213 (N_6213,N_2535,N_227);
nor U6214 (N_6214,N_3442,N_3600);
or U6215 (N_6215,N_3819,N_286);
or U6216 (N_6216,N_804,N_3231);
nand U6217 (N_6217,N_1907,N_3623);
or U6218 (N_6218,N_3148,N_395);
nor U6219 (N_6219,N_3094,N_3140);
nand U6220 (N_6220,N_3235,N_2561);
nand U6221 (N_6221,N_1392,N_3845);
or U6222 (N_6222,N_1441,N_191);
xor U6223 (N_6223,N_3202,N_3059);
or U6224 (N_6224,N_2526,N_1529);
and U6225 (N_6225,N_3430,N_1872);
xnor U6226 (N_6226,N_2558,N_1836);
and U6227 (N_6227,N_1967,N_119);
and U6228 (N_6228,N_837,N_707);
or U6229 (N_6229,N_32,N_1299);
and U6230 (N_6230,N_733,N_3732);
and U6231 (N_6231,N_530,N_674);
or U6232 (N_6232,N_3748,N_3649);
nor U6233 (N_6233,N_3186,N_2324);
nand U6234 (N_6234,N_3494,N_1738);
xnor U6235 (N_6235,N_2780,N_2686);
or U6236 (N_6236,N_3343,N_966);
or U6237 (N_6237,N_3214,N_2882);
nor U6238 (N_6238,N_997,N_2225);
nor U6239 (N_6239,N_2323,N_486);
and U6240 (N_6240,N_2562,N_1453);
nor U6241 (N_6241,N_291,N_2832);
xor U6242 (N_6242,N_3265,N_2944);
or U6243 (N_6243,N_3661,N_2894);
and U6244 (N_6244,N_569,N_3361);
xnor U6245 (N_6245,N_1007,N_3579);
nor U6246 (N_6246,N_1203,N_38);
or U6247 (N_6247,N_3575,N_2341);
nand U6248 (N_6248,N_3855,N_2872);
nor U6249 (N_6249,N_3326,N_3798);
xor U6250 (N_6250,N_1836,N_16);
xor U6251 (N_6251,N_851,N_335);
or U6252 (N_6252,N_2525,N_3553);
nor U6253 (N_6253,N_3737,N_2684);
and U6254 (N_6254,N_616,N_3254);
nor U6255 (N_6255,N_3684,N_3493);
nand U6256 (N_6256,N_1868,N_1245);
nor U6257 (N_6257,N_3233,N_1362);
nor U6258 (N_6258,N_3319,N_618);
xor U6259 (N_6259,N_1578,N_3385);
nor U6260 (N_6260,N_3721,N_2845);
or U6261 (N_6261,N_1952,N_1918);
nor U6262 (N_6262,N_3415,N_1103);
and U6263 (N_6263,N_368,N_1062);
and U6264 (N_6264,N_2805,N_1821);
or U6265 (N_6265,N_97,N_3685);
nand U6266 (N_6266,N_1285,N_289);
xor U6267 (N_6267,N_473,N_2991);
or U6268 (N_6268,N_2770,N_1533);
nand U6269 (N_6269,N_2968,N_3943);
nor U6270 (N_6270,N_1871,N_3713);
and U6271 (N_6271,N_1738,N_3061);
nor U6272 (N_6272,N_498,N_1526);
nand U6273 (N_6273,N_1918,N_559);
and U6274 (N_6274,N_1160,N_730);
nor U6275 (N_6275,N_847,N_835);
nand U6276 (N_6276,N_2157,N_2390);
or U6277 (N_6277,N_1451,N_3621);
xnor U6278 (N_6278,N_1665,N_228);
or U6279 (N_6279,N_3310,N_1354);
or U6280 (N_6280,N_2722,N_715);
and U6281 (N_6281,N_1916,N_1766);
nand U6282 (N_6282,N_2975,N_2276);
or U6283 (N_6283,N_846,N_2260);
or U6284 (N_6284,N_39,N_389);
and U6285 (N_6285,N_737,N_1547);
and U6286 (N_6286,N_3460,N_2525);
xor U6287 (N_6287,N_41,N_1343);
or U6288 (N_6288,N_3104,N_1437);
xor U6289 (N_6289,N_1950,N_142);
and U6290 (N_6290,N_2704,N_2583);
xnor U6291 (N_6291,N_3318,N_1477);
nand U6292 (N_6292,N_740,N_422);
nand U6293 (N_6293,N_1900,N_1001);
nand U6294 (N_6294,N_1384,N_3657);
nor U6295 (N_6295,N_2982,N_69);
nand U6296 (N_6296,N_1808,N_2860);
or U6297 (N_6297,N_3290,N_2653);
nand U6298 (N_6298,N_2943,N_3221);
nor U6299 (N_6299,N_379,N_589);
or U6300 (N_6300,N_3336,N_2837);
nand U6301 (N_6301,N_1504,N_644);
and U6302 (N_6302,N_1273,N_1458);
and U6303 (N_6303,N_3568,N_2623);
nor U6304 (N_6304,N_2598,N_3629);
or U6305 (N_6305,N_877,N_2315);
nand U6306 (N_6306,N_2212,N_3732);
nor U6307 (N_6307,N_3149,N_2925);
xor U6308 (N_6308,N_1675,N_2731);
or U6309 (N_6309,N_2209,N_29);
nor U6310 (N_6310,N_2773,N_678);
xor U6311 (N_6311,N_3054,N_3996);
nand U6312 (N_6312,N_2778,N_3293);
nand U6313 (N_6313,N_2306,N_781);
or U6314 (N_6314,N_2126,N_2366);
nor U6315 (N_6315,N_3076,N_822);
nor U6316 (N_6316,N_1283,N_82);
or U6317 (N_6317,N_3482,N_2658);
and U6318 (N_6318,N_3645,N_3740);
and U6319 (N_6319,N_139,N_1191);
and U6320 (N_6320,N_3890,N_716);
nand U6321 (N_6321,N_2641,N_467);
or U6322 (N_6322,N_910,N_2046);
or U6323 (N_6323,N_1158,N_2443);
and U6324 (N_6324,N_2791,N_1740);
and U6325 (N_6325,N_3223,N_2223);
nor U6326 (N_6326,N_431,N_1379);
and U6327 (N_6327,N_1182,N_1858);
and U6328 (N_6328,N_2175,N_2225);
xor U6329 (N_6329,N_1529,N_2681);
and U6330 (N_6330,N_2896,N_2353);
nor U6331 (N_6331,N_3799,N_1470);
nand U6332 (N_6332,N_1217,N_2409);
or U6333 (N_6333,N_337,N_1100);
or U6334 (N_6334,N_2354,N_455);
nand U6335 (N_6335,N_886,N_1639);
nor U6336 (N_6336,N_2270,N_988);
or U6337 (N_6337,N_1843,N_976);
and U6338 (N_6338,N_1345,N_1571);
nand U6339 (N_6339,N_954,N_977);
or U6340 (N_6340,N_2586,N_2744);
nor U6341 (N_6341,N_986,N_3887);
or U6342 (N_6342,N_1179,N_2996);
nor U6343 (N_6343,N_3298,N_481);
xnor U6344 (N_6344,N_2085,N_2603);
xnor U6345 (N_6345,N_92,N_1122);
or U6346 (N_6346,N_2806,N_1594);
xor U6347 (N_6347,N_1932,N_3148);
nand U6348 (N_6348,N_2719,N_812);
nor U6349 (N_6349,N_3088,N_1288);
or U6350 (N_6350,N_3369,N_3551);
or U6351 (N_6351,N_3054,N_1998);
nor U6352 (N_6352,N_1889,N_485);
nand U6353 (N_6353,N_3667,N_3871);
or U6354 (N_6354,N_2995,N_168);
xor U6355 (N_6355,N_3737,N_1717);
or U6356 (N_6356,N_2127,N_402);
nand U6357 (N_6357,N_1594,N_2656);
and U6358 (N_6358,N_119,N_1803);
nand U6359 (N_6359,N_2417,N_1236);
nor U6360 (N_6360,N_2324,N_237);
or U6361 (N_6361,N_132,N_3205);
nand U6362 (N_6362,N_435,N_3241);
and U6363 (N_6363,N_306,N_3329);
nor U6364 (N_6364,N_99,N_1413);
nor U6365 (N_6365,N_2271,N_1171);
and U6366 (N_6366,N_2195,N_1507);
nor U6367 (N_6367,N_2668,N_460);
or U6368 (N_6368,N_623,N_2435);
nor U6369 (N_6369,N_1415,N_1871);
or U6370 (N_6370,N_1851,N_597);
nor U6371 (N_6371,N_2169,N_1936);
or U6372 (N_6372,N_2,N_3532);
nand U6373 (N_6373,N_3950,N_3458);
and U6374 (N_6374,N_564,N_2549);
and U6375 (N_6375,N_1961,N_1450);
nor U6376 (N_6376,N_2465,N_764);
or U6377 (N_6377,N_3852,N_958);
and U6378 (N_6378,N_2712,N_3370);
and U6379 (N_6379,N_1634,N_1093);
nand U6380 (N_6380,N_784,N_326);
or U6381 (N_6381,N_1576,N_249);
and U6382 (N_6382,N_507,N_2639);
nor U6383 (N_6383,N_2812,N_2876);
xnor U6384 (N_6384,N_1536,N_653);
nor U6385 (N_6385,N_2082,N_2730);
xnor U6386 (N_6386,N_2535,N_956);
xnor U6387 (N_6387,N_1784,N_2084);
or U6388 (N_6388,N_2683,N_3081);
xnor U6389 (N_6389,N_2308,N_2359);
or U6390 (N_6390,N_198,N_2234);
nand U6391 (N_6391,N_16,N_1734);
nand U6392 (N_6392,N_1383,N_2131);
nand U6393 (N_6393,N_2081,N_2387);
and U6394 (N_6394,N_3148,N_3839);
and U6395 (N_6395,N_486,N_2392);
or U6396 (N_6396,N_3420,N_1302);
and U6397 (N_6397,N_466,N_2402);
and U6398 (N_6398,N_1875,N_2762);
xor U6399 (N_6399,N_65,N_3928);
or U6400 (N_6400,N_3211,N_2869);
nor U6401 (N_6401,N_1830,N_782);
nand U6402 (N_6402,N_2664,N_3521);
nand U6403 (N_6403,N_865,N_1680);
nor U6404 (N_6404,N_496,N_893);
nor U6405 (N_6405,N_915,N_2662);
nand U6406 (N_6406,N_143,N_1837);
xnor U6407 (N_6407,N_158,N_2114);
and U6408 (N_6408,N_3969,N_3583);
or U6409 (N_6409,N_2246,N_3724);
nor U6410 (N_6410,N_365,N_3908);
nor U6411 (N_6411,N_1822,N_1297);
or U6412 (N_6412,N_3387,N_1856);
and U6413 (N_6413,N_2614,N_3337);
and U6414 (N_6414,N_1302,N_593);
xor U6415 (N_6415,N_2748,N_3499);
and U6416 (N_6416,N_1280,N_3773);
nor U6417 (N_6417,N_3491,N_2300);
and U6418 (N_6418,N_1371,N_2288);
nand U6419 (N_6419,N_3094,N_260);
nand U6420 (N_6420,N_3338,N_601);
nor U6421 (N_6421,N_2298,N_2414);
and U6422 (N_6422,N_2908,N_3552);
nor U6423 (N_6423,N_3339,N_1707);
or U6424 (N_6424,N_2500,N_3212);
nand U6425 (N_6425,N_147,N_1752);
nand U6426 (N_6426,N_54,N_2583);
nor U6427 (N_6427,N_1571,N_1982);
or U6428 (N_6428,N_419,N_504);
nand U6429 (N_6429,N_1217,N_2317);
nand U6430 (N_6430,N_1397,N_397);
nor U6431 (N_6431,N_3203,N_1195);
nor U6432 (N_6432,N_807,N_202);
and U6433 (N_6433,N_2824,N_529);
or U6434 (N_6434,N_1347,N_1432);
and U6435 (N_6435,N_759,N_1795);
nor U6436 (N_6436,N_2427,N_3462);
nor U6437 (N_6437,N_1794,N_3112);
nand U6438 (N_6438,N_42,N_925);
nand U6439 (N_6439,N_2266,N_815);
nor U6440 (N_6440,N_3705,N_1557);
nand U6441 (N_6441,N_480,N_406);
and U6442 (N_6442,N_2415,N_3780);
nor U6443 (N_6443,N_3750,N_1370);
nand U6444 (N_6444,N_3465,N_3770);
or U6445 (N_6445,N_1060,N_2621);
or U6446 (N_6446,N_2808,N_256);
nand U6447 (N_6447,N_3605,N_906);
xor U6448 (N_6448,N_2256,N_386);
xor U6449 (N_6449,N_2426,N_2891);
or U6450 (N_6450,N_3922,N_105);
nor U6451 (N_6451,N_3575,N_1252);
or U6452 (N_6452,N_1637,N_2516);
and U6453 (N_6453,N_2278,N_1837);
or U6454 (N_6454,N_1744,N_2723);
nor U6455 (N_6455,N_3256,N_2458);
nand U6456 (N_6456,N_930,N_2979);
nand U6457 (N_6457,N_2048,N_3816);
xor U6458 (N_6458,N_117,N_2936);
and U6459 (N_6459,N_3038,N_1368);
nand U6460 (N_6460,N_3249,N_703);
or U6461 (N_6461,N_1582,N_3826);
nor U6462 (N_6462,N_1558,N_653);
or U6463 (N_6463,N_2957,N_3622);
nor U6464 (N_6464,N_2795,N_2437);
nor U6465 (N_6465,N_701,N_922);
nand U6466 (N_6466,N_2591,N_1534);
nand U6467 (N_6467,N_2877,N_57);
or U6468 (N_6468,N_1400,N_3648);
nor U6469 (N_6469,N_2862,N_526);
or U6470 (N_6470,N_1106,N_2556);
and U6471 (N_6471,N_3244,N_2952);
and U6472 (N_6472,N_2913,N_3356);
xor U6473 (N_6473,N_1040,N_3702);
xnor U6474 (N_6474,N_288,N_2615);
and U6475 (N_6475,N_3533,N_3853);
nor U6476 (N_6476,N_1318,N_1109);
xor U6477 (N_6477,N_186,N_1366);
xnor U6478 (N_6478,N_684,N_2876);
nor U6479 (N_6479,N_924,N_1275);
nand U6480 (N_6480,N_3511,N_1203);
or U6481 (N_6481,N_2244,N_347);
or U6482 (N_6482,N_2452,N_1535);
and U6483 (N_6483,N_3749,N_2011);
nor U6484 (N_6484,N_3418,N_789);
or U6485 (N_6485,N_1137,N_1447);
nand U6486 (N_6486,N_1850,N_515);
nand U6487 (N_6487,N_760,N_909);
nand U6488 (N_6488,N_1398,N_2861);
and U6489 (N_6489,N_1641,N_394);
or U6490 (N_6490,N_2342,N_1295);
nand U6491 (N_6491,N_2630,N_124);
nor U6492 (N_6492,N_3780,N_2286);
or U6493 (N_6493,N_185,N_177);
xor U6494 (N_6494,N_382,N_28);
nor U6495 (N_6495,N_1493,N_1560);
nand U6496 (N_6496,N_2996,N_2382);
nor U6497 (N_6497,N_2338,N_3476);
and U6498 (N_6498,N_2990,N_69);
nor U6499 (N_6499,N_3496,N_2523);
nor U6500 (N_6500,N_1825,N_2985);
nor U6501 (N_6501,N_1913,N_3787);
nand U6502 (N_6502,N_3681,N_2682);
or U6503 (N_6503,N_1540,N_1715);
or U6504 (N_6504,N_1512,N_2614);
and U6505 (N_6505,N_2595,N_2587);
and U6506 (N_6506,N_3231,N_3463);
xnor U6507 (N_6507,N_3743,N_2978);
and U6508 (N_6508,N_2026,N_2177);
nor U6509 (N_6509,N_3857,N_3776);
nor U6510 (N_6510,N_518,N_2765);
or U6511 (N_6511,N_602,N_495);
nor U6512 (N_6512,N_3141,N_1656);
nand U6513 (N_6513,N_890,N_1461);
nand U6514 (N_6514,N_2663,N_2054);
or U6515 (N_6515,N_1742,N_3628);
nand U6516 (N_6516,N_2360,N_3076);
nor U6517 (N_6517,N_1995,N_935);
nor U6518 (N_6518,N_3055,N_373);
or U6519 (N_6519,N_3046,N_583);
or U6520 (N_6520,N_2211,N_498);
nor U6521 (N_6521,N_606,N_2927);
nor U6522 (N_6522,N_2799,N_481);
nor U6523 (N_6523,N_2290,N_13);
nor U6524 (N_6524,N_1746,N_2302);
nor U6525 (N_6525,N_2930,N_3928);
nand U6526 (N_6526,N_640,N_1465);
or U6527 (N_6527,N_3366,N_1821);
nor U6528 (N_6528,N_1213,N_2148);
and U6529 (N_6529,N_2769,N_2931);
nor U6530 (N_6530,N_2113,N_1634);
nand U6531 (N_6531,N_3015,N_598);
nand U6532 (N_6532,N_3504,N_2822);
nor U6533 (N_6533,N_933,N_1938);
nand U6534 (N_6534,N_1009,N_3640);
xor U6535 (N_6535,N_2674,N_117);
and U6536 (N_6536,N_2791,N_3673);
nand U6537 (N_6537,N_3956,N_1637);
and U6538 (N_6538,N_2461,N_1013);
nor U6539 (N_6539,N_1807,N_656);
or U6540 (N_6540,N_1342,N_2061);
nand U6541 (N_6541,N_1549,N_1402);
or U6542 (N_6542,N_2629,N_3735);
or U6543 (N_6543,N_1448,N_885);
nor U6544 (N_6544,N_554,N_266);
or U6545 (N_6545,N_1001,N_795);
nand U6546 (N_6546,N_1785,N_3162);
nor U6547 (N_6547,N_910,N_1182);
nand U6548 (N_6548,N_775,N_647);
nor U6549 (N_6549,N_1561,N_2075);
nand U6550 (N_6550,N_1820,N_538);
xnor U6551 (N_6551,N_894,N_3003);
or U6552 (N_6552,N_3937,N_3809);
and U6553 (N_6553,N_575,N_3602);
or U6554 (N_6554,N_1014,N_2603);
and U6555 (N_6555,N_3777,N_1381);
nand U6556 (N_6556,N_1525,N_394);
nand U6557 (N_6557,N_3008,N_1803);
and U6558 (N_6558,N_3146,N_2616);
nand U6559 (N_6559,N_2988,N_3897);
or U6560 (N_6560,N_2800,N_3676);
nor U6561 (N_6561,N_1725,N_3398);
or U6562 (N_6562,N_915,N_3396);
and U6563 (N_6563,N_605,N_3704);
nor U6564 (N_6564,N_3429,N_332);
and U6565 (N_6565,N_3603,N_3515);
nor U6566 (N_6566,N_2109,N_2216);
nand U6567 (N_6567,N_1978,N_4);
or U6568 (N_6568,N_3697,N_3419);
xor U6569 (N_6569,N_848,N_512);
and U6570 (N_6570,N_1550,N_1954);
nand U6571 (N_6571,N_3481,N_53);
and U6572 (N_6572,N_2004,N_1518);
and U6573 (N_6573,N_3455,N_1197);
and U6574 (N_6574,N_1061,N_2592);
nand U6575 (N_6575,N_282,N_1725);
and U6576 (N_6576,N_2412,N_2827);
and U6577 (N_6577,N_2782,N_1673);
or U6578 (N_6578,N_3788,N_3292);
nand U6579 (N_6579,N_673,N_2405);
or U6580 (N_6580,N_616,N_2431);
nand U6581 (N_6581,N_2178,N_3150);
and U6582 (N_6582,N_741,N_3907);
nand U6583 (N_6583,N_1541,N_2033);
nor U6584 (N_6584,N_2939,N_3667);
or U6585 (N_6585,N_1251,N_3860);
nand U6586 (N_6586,N_1482,N_549);
and U6587 (N_6587,N_573,N_3742);
or U6588 (N_6588,N_1288,N_2305);
nand U6589 (N_6589,N_2106,N_3046);
xnor U6590 (N_6590,N_1036,N_2713);
nor U6591 (N_6591,N_1013,N_2293);
or U6592 (N_6592,N_1422,N_2392);
nor U6593 (N_6593,N_854,N_2908);
or U6594 (N_6594,N_2258,N_1016);
nand U6595 (N_6595,N_2510,N_2736);
nor U6596 (N_6596,N_1582,N_581);
nor U6597 (N_6597,N_2090,N_3445);
and U6598 (N_6598,N_1548,N_3341);
nand U6599 (N_6599,N_178,N_2626);
nor U6600 (N_6600,N_3688,N_881);
and U6601 (N_6601,N_636,N_3968);
and U6602 (N_6602,N_3113,N_3292);
nor U6603 (N_6603,N_925,N_509);
and U6604 (N_6604,N_3259,N_1083);
or U6605 (N_6605,N_2835,N_2660);
or U6606 (N_6606,N_1482,N_3996);
xor U6607 (N_6607,N_973,N_2989);
nand U6608 (N_6608,N_139,N_2773);
nor U6609 (N_6609,N_3545,N_677);
nand U6610 (N_6610,N_3330,N_1395);
and U6611 (N_6611,N_2726,N_1561);
or U6612 (N_6612,N_2967,N_1180);
and U6613 (N_6613,N_2441,N_267);
or U6614 (N_6614,N_3708,N_3503);
or U6615 (N_6615,N_3211,N_2472);
or U6616 (N_6616,N_3371,N_3702);
or U6617 (N_6617,N_930,N_3878);
nor U6618 (N_6618,N_2373,N_1329);
and U6619 (N_6619,N_2769,N_2138);
or U6620 (N_6620,N_2540,N_8);
and U6621 (N_6621,N_3999,N_1167);
or U6622 (N_6622,N_2444,N_363);
or U6623 (N_6623,N_2718,N_2389);
nand U6624 (N_6624,N_1377,N_667);
and U6625 (N_6625,N_668,N_3959);
nand U6626 (N_6626,N_1538,N_2633);
nand U6627 (N_6627,N_279,N_1954);
nand U6628 (N_6628,N_2316,N_60);
nor U6629 (N_6629,N_3854,N_2074);
nand U6630 (N_6630,N_3506,N_460);
or U6631 (N_6631,N_2758,N_1935);
xor U6632 (N_6632,N_1845,N_3369);
nand U6633 (N_6633,N_1488,N_1316);
and U6634 (N_6634,N_2441,N_509);
or U6635 (N_6635,N_2045,N_135);
and U6636 (N_6636,N_3553,N_1904);
nand U6637 (N_6637,N_3169,N_386);
and U6638 (N_6638,N_1085,N_607);
nor U6639 (N_6639,N_3621,N_1529);
nor U6640 (N_6640,N_1182,N_2582);
or U6641 (N_6641,N_2165,N_365);
nand U6642 (N_6642,N_634,N_969);
and U6643 (N_6643,N_3308,N_1117);
and U6644 (N_6644,N_2013,N_2079);
nor U6645 (N_6645,N_486,N_3964);
nor U6646 (N_6646,N_3249,N_1299);
nor U6647 (N_6647,N_129,N_527);
nand U6648 (N_6648,N_174,N_171);
nand U6649 (N_6649,N_3860,N_2271);
nor U6650 (N_6650,N_81,N_2422);
nor U6651 (N_6651,N_2830,N_2623);
nor U6652 (N_6652,N_285,N_1020);
and U6653 (N_6653,N_2931,N_424);
or U6654 (N_6654,N_854,N_2896);
nand U6655 (N_6655,N_1305,N_1092);
nor U6656 (N_6656,N_3964,N_932);
xnor U6657 (N_6657,N_1405,N_2397);
or U6658 (N_6658,N_592,N_437);
xor U6659 (N_6659,N_3264,N_3915);
nand U6660 (N_6660,N_863,N_3544);
and U6661 (N_6661,N_3631,N_1946);
or U6662 (N_6662,N_658,N_70);
nand U6663 (N_6663,N_3913,N_3731);
and U6664 (N_6664,N_685,N_1960);
nand U6665 (N_6665,N_844,N_1961);
nand U6666 (N_6666,N_1399,N_1073);
nand U6667 (N_6667,N_2575,N_3489);
nor U6668 (N_6668,N_1495,N_1501);
nand U6669 (N_6669,N_1293,N_3787);
nor U6670 (N_6670,N_2366,N_3948);
nor U6671 (N_6671,N_2845,N_3069);
xnor U6672 (N_6672,N_1868,N_803);
xor U6673 (N_6673,N_1185,N_1412);
and U6674 (N_6674,N_368,N_290);
nor U6675 (N_6675,N_375,N_635);
nand U6676 (N_6676,N_3871,N_3686);
nand U6677 (N_6677,N_231,N_3558);
nor U6678 (N_6678,N_1389,N_3194);
or U6679 (N_6679,N_3598,N_2777);
xnor U6680 (N_6680,N_1630,N_1850);
nand U6681 (N_6681,N_2688,N_3869);
nor U6682 (N_6682,N_107,N_3027);
and U6683 (N_6683,N_1062,N_2426);
nand U6684 (N_6684,N_36,N_1559);
or U6685 (N_6685,N_1131,N_740);
nand U6686 (N_6686,N_482,N_1381);
nand U6687 (N_6687,N_2690,N_2200);
nand U6688 (N_6688,N_507,N_634);
nand U6689 (N_6689,N_3052,N_2118);
and U6690 (N_6690,N_2296,N_3552);
xor U6691 (N_6691,N_3608,N_384);
and U6692 (N_6692,N_30,N_3009);
or U6693 (N_6693,N_1399,N_558);
nor U6694 (N_6694,N_2013,N_23);
nand U6695 (N_6695,N_1756,N_1578);
nand U6696 (N_6696,N_603,N_942);
nand U6697 (N_6697,N_2321,N_2799);
nor U6698 (N_6698,N_3738,N_669);
nand U6699 (N_6699,N_338,N_1478);
and U6700 (N_6700,N_1483,N_711);
or U6701 (N_6701,N_3391,N_1623);
and U6702 (N_6702,N_2738,N_3172);
or U6703 (N_6703,N_623,N_852);
nor U6704 (N_6704,N_3391,N_2722);
nand U6705 (N_6705,N_2321,N_2298);
nand U6706 (N_6706,N_3073,N_3804);
xor U6707 (N_6707,N_1385,N_846);
nor U6708 (N_6708,N_3956,N_179);
nand U6709 (N_6709,N_3019,N_2071);
nand U6710 (N_6710,N_3411,N_188);
nand U6711 (N_6711,N_2277,N_3951);
and U6712 (N_6712,N_2529,N_3684);
nand U6713 (N_6713,N_1796,N_3552);
or U6714 (N_6714,N_3812,N_2452);
nand U6715 (N_6715,N_1549,N_1035);
nand U6716 (N_6716,N_268,N_1786);
nor U6717 (N_6717,N_1464,N_2626);
and U6718 (N_6718,N_855,N_763);
nand U6719 (N_6719,N_1155,N_1252);
and U6720 (N_6720,N_2411,N_3561);
or U6721 (N_6721,N_1955,N_1045);
or U6722 (N_6722,N_1746,N_2711);
or U6723 (N_6723,N_1114,N_2525);
or U6724 (N_6724,N_739,N_3714);
nand U6725 (N_6725,N_487,N_3331);
xor U6726 (N_6726,N_220,N_1314);
nor U6727 (N_6727,N_767,N_1111);
nor U6728 (N_6728,N_578,N_2652);
and U6729 (N_6729,N_3586,N_791);
xnor U6730 (N_6730,N_3287,N_3532);
or U6731 (N_6731,N_1109,N_1661);
nand U6732 (N_6732,N_552,N_1807);
nand U6733 (N_6733,N_1852,N_3880);
xnor U6734 (N_6734,N_1716,N_3008);
and U6735 (N_6735,N_3279,N_3332);
and U6736 (N_6736,N_3704,N_153);
nor U6737 (N_6737,N_1751,N_1236);
or U6738 (N_6738,N_3620,N_941);
nand U6739 (N_6739,N_3407,N_2300);
nor U6740 (N_6740,N_983,N_702);
and U6741 (N_6741,N_1826,N_2925);
xnor U6742 (N_6742,N_1008,N_3314);
and U6743 (N_6743,N_3246,N_1005);
nand U6744 (N_6744,N_3907,N_329);
nand U6745 (N_6745,N_2457,N_558);
xor U6746 (N_6746,N_1850,N_3092);
and U6747 (N_6747,N_3054,N_864);
and U6748 (N_6748,N_3005,N_3284);
and U6749 (N_6749,N_3095,N_1348);
nor U6750 (N_6750,N_2187,N_1052);
nand U6751 (N_6751,N_817,N_274);
nand U6752 (N_6752,N_2954,N_3724);
or U6753 (N_6753,N_1481,N_1721);
nor U6754 (N_6754,N_2083,N_592);
nor U6755 (N_6755,N_3783,N_41);
xor U6756 (N_6756,N_1488,N_1052);
xor U6757 (N_6757,N_2505,N_2018);
and U6758 (N_6758,N_573,N_950);
or U6759 (N_6759,N_3060,N_183);
and U6760 (N_6760,N_3403,N_1943);
nor U6761 (N_6761,N_1154,N_908);
and U6762 (N_6762,N_987,N_2634);
nor U6763 (N_6763,N_2167,N_1685);
or U6764 (N_6764,N_1525,N_2064);
or U6765 (N_6765,N_3838,N_1724);
nand U6766 (N_6766,N_210,N_644);
nand U6767 (N_6767,N_2686,N_135);
xnor U6768 (N_6768,N_1496,N_629);
nand U6769 (N_6769,N_1595,N_1378);
nor U6770 (N_6770,N_418,N_3157);
nor U6771 (N_6771,N_3432,N_2338);
nand U6772 (N_6772,N_1372,N_3731);
or U6773 (N_6773,N_1637,N_3213);
or U6774 (N_6774,N_2077,N_1504);
and U6775 (N_6775,N_139,N_537);
and U6776 (N_6776,N_842,N_3241);
nand U6777 (N_6777,N_1108,N_3574);
nor U6778 (N_6778,N_2480,N_3696);
or U6779 (N_6779,N_3624,N_2914);
and U6780 (N_6780,N_853,N_413);
xnor U6781 (N_6781,N_50,N_106);
nor U6782 (N_6782,N_871,N_2220);
nand U6783 (N_6783,N_2229,N_1887);
xnor U6784 (N_6784,N_3508,N_453);
nand U6785 (N_6785,N_2009,N_249);
xor U6786 (N_6786,N_32,N_1763);
or U6787 (N_6787,N_116,N_1827);
and U6788 (N_6788,N_2131,N_1160);
and U6789 (N_6789,N_1572,N_1015);
nand U6790 (N_6790,N_1024,N_3437);
nor U6791 (N_6791,N_2807,N_2659);
nand U6792 (N_6792,N_3886,N_1782);
xnor U6793 (N_6793,N_2456,N_212);
nand U6794 (N_6794,N_3642,N_1562);
or U6795 (N_6795,N_1615,N_1304);
nand U6796 (N_6796,N_1545,N_1589);
xnor U6797 (N_6797,N_1709,N_3743);
nand U6798 (N_6798,N_1463,N_3095);
and U6799 (N_6799,N_2811,N_276);
and U6800 (N_6800,N_3744,N_3961);
and U6801 (N_6801,N_3807,N_746);
nand U6802 (N_6802,N_1490,N_1950);
nand U6803 (N_6803,N_1114,N_1662);
xor U6804 (N_6804,N_3963,N_923);
nor U6805 (N_6805,N_247,N_1957);
and U6806 (N_6806,N_1127,N_3834);
xor U6807 (N_6807,N_1728,N_2425);
nand U6808 (N_6808,N_1834,N_3000);
and U6809 (N_6809,N_3333,N_1628);
or U6810 (N_6810,N_3982,N_1383);
and U6811 (N_6811,N_842,N_3247);
or U6812 (N_6812,N_677,N_568);
or U6813 (N_6813,N_3913,N_1191);
and U6814 (N_6814,N_3941,N_1899);
nor U6815 (N_6815,N_943,N_1118);
nand U6816 (N_6816,N_262,N_3660);
nand U6817 (N_6817,N_3289,N_477);
or U6818 (N_6818,N_2325,N_3951);
or U6819 (N_6819,N_2067,N_3284);
or U6820 (N_6820,N_572,N_2033);
or U6821 (N_6821,N_3923,N_3467);
and U6822 (N_6822,N_599,N_1904);
or U6823 (N_6823,N_3585,N_2950);
nor U6824 (N_6824,N_3788,N_2465);
or U6825 (N_6825,N_3595,N_1331);
or U6826 (N_6826,N_2802,N_2931);
nor U6827 (N_6827,N_3179,N_3117);
nor U6828 (N_6828,N_1504,N_2763);
nor U6829 (N_6829,N_3031,N_1176);
or U6830 (N_6830,N_856,N_1082);
and U6831 (N_6831,N_1880,N_2656);
nand U6832 (N_6832,N_2300,N_3985);
or U6833 (N_6833,N_133,N_2396);
nand U6834 (N_6834,N_793,N_540);
nor U6835 (N_6835,N_3478,N_890);
nand U6836 (N_6836,N_2349,N_1247);
nand U6837 (N_6837,N_1480,N_3894);
nand U6838 (N_6838,N_3367,N_2735);
and U6839 (N_6839,N_1743,N_2300);
and U6840 (N_6840,N_2103,N_3454);
or U6841 (N_6841,N_3280,N_1785);
and U6842 (N_6842,N_521,N_1265);
nand U6843 (N_6843,N_561,N_3693);
nor U6844 (N_6844,N_2813,N_1446);
and U6845 (N_6845,N_773,N_700);
and U6846 (N_6846,N_696,N_885);
and U6847 (N_6847,N_2564,N_771);
and U6848 (N_6848,N_2300,N_43);
nor U6849 (N_6849,N_1168,N_521);
or U6850 (N_6850,N_1332,N_1313);
nor U6851 (N_6851,N_2954,N_1009);
or U6852 (N_6852,N_574,N_3171);
or U6853 (N_6853,N_2199,N_2044);
nor U6854 (N_6854,N_1417,N_942);
or U6855 (N_6855,N_1646,N_3505);
nand U6856 (N_6856,N_2738,N_2438);
or U6857 (N_6857,N_867,N_2662);
or U6858 (N_6858,N_139,N_584);
or U6859 (N_6859,N_414,N_352);
or U6860 (N_6860,N_1085,N_1357);
xor U6861 (N_6861,N_2504,N_3466);
nor U6862 (N_6862,N_281,N_1181);
xnor U6863 (N_6863,N_3735,N_1058);
nor U6864 (N_6864,N_3172,N_478);
and U6865 (N_6865,N_3648,N_3456);
and U6866 (N_6866,N_2337,N_3133);
xor U6867 (N_6867,N_1015,N_471);
nor U6868 (N_6868,N_476,N_1526);
and U6869 (N_6869,N_1573,N_404);
nand U6870 (N_6870,N_660,N_3723);
nand U6871 (N_6871,N_3724,N_500);
nor U6872 (N_6872,N_1315,N_3733);
nor U6873 (N_6873,N_2873,N_2374);
nor U6874 (N_6874,N_276,N_1546);
and U6875 (N_6875,N_3394,N_349);
or U6876 (N_6876,N_1747,N_3480);
nand U6877 (N_6877,N_674,N_3861);
and U6878 (N_6878,N_630,N_1399);
nor U6879 (N_6879,N_3558,N_1430);
xnor U6880 (N_6880,N_2527,N_1634);
and U6881 (N_6881,N_2529,N_488);
and U6882 (N_6882,N_3896,N_3222);
and U6883 (N_6883,N_2934,N_1440);
and U6884 (N_6884,N_3922,N_3578);
nand U6885 (N_6885,N_1107,N_2877);
nand U6886 (N_6886,N_2532,N_1120);
and U6887 (N_6887,N_1214,N_1923);
nand U6888 (N_6888,N_46,N_3432);
and U6889 (N_6889,N_2810,N_387);
nor U6890 (N_6890,N_3833,N_3306);
xnor U6891 (N_6891,N_1397,N_830);
and U6892 (N_6892,N_3403,N_650);
nor U6893 (N_6893,N_3557,N_86);
nor U6894 (N_6894,N_2296,N_2538);
or U6895 (N_6895,N_3165,N_1101);
nand U6896 (N_6896,N_262,N_2092);
or U6897 (N_6897,N_1323,N_1745);
and U6898 (N_6898,N_1710,N_1384);
xnor U6899 (N_6899,N_1293,N_3205);
or U6900 (N_6900,N_2056,N_241);
xnor U6901 (N_6901,N_918,N_654);
nand U6902 (N_6902,N_2130,N_1482);
and U6903 (N_6903,N_1288,N_667);
and U6904 (N_6904,N_2105,N_1344);
nand U6905 (N_6905,N_1856,N_3180);
nand U6906 (N_6906,N_2475,N_3787);
nor U6907 (N_6907,N_1501,N_1316);
xor U6908 (N_6908,N_244,N_3777);
xor U6909 (N_6909,N_3877,N_854);
nor U6910 (N_6910,N_1182,N_3633);
or U6911 (N_6911,N_3577,N_126);
or U6912 (N_6912,N_3900,N_2482);
nand U6913 (N_6913,N_737,N_2108);
nor U6914 (N_6914,N_1542,N_2938);
or U6915 (N_6915,N_153,N_498);
nor U6916 (N_6916,N_256,N_3675);
nor U6917 (N_6917,N_137,N_3168);
and U6918 (N_6918,N_3678,N_1737);
or U6919 (N_6919,N_571,N_124);
xnor U6920 (N_6920,N_1089,N_1319);
nand U6921 (N_6921,N_538,N_1320);
or U6922 (N_6922,N_281,N_968);
and U6923 (N_6923,N_244,N_2368);
nand U6924 (N_6924,N_3050,N_2665);
nand U6925 (N_6925,N_2926,N_2871);
or U6926 (N_6926,N_2676,N_2909);
nand U6927 (N_6927,N_2066,N_3140);
or U6928 (N_6928,N_1864,N_3810);
or U6929 (N_6929,N_1491,N_1742);
nand U6930 (N_6930,N_2643,N_753);
xor U6931 (N_6931,N_2435,N_3308);
or U6932 (N_6932,N_2742,N_3356);
nor U6933 (N_6933,N_1069,N_2569);
or U6934 (N_6934,N_3388,N_2943);
and U6935 (N_6935,N_2280,N_193);
nor U6936 (N_6936,N_3305,N_1911);
or U6937 (N_6937,N_2942,N_389);
nand U6938 (N_6938,N_690,N_1253);
xnor U6939 (N_6939,N_1637,N_1083);
nand U6940 (N_6940,N_3566,N_2324);
nand U6941 (N_6941,N_907,N_1193);
nor U6942 (N_6942,N_1143,N_565);
nor U6943 (N_6943,N_1492,N_3181);
nand U6944 (N_6944,N_113,N_3160);
nor U6945 (N_6945,N_2676,N_862);
xnor U6946 (N_6946,N_575,N_2077);
or U6947 (N_6947,N_438,N_1079);
or U6948 (N_6948,N_3880,N_1196);
or U6949 (N_6949,N_995,N_3391);
and U6950 (N_6950,N_3386,N_1070);
or U6951 (N_6951,N_1728,N_3303);
or U6952 (N_6952,N_2730,N_1860);
nand U6953 (N_6953,N_3151,N_2981);
xor U6954 (N_6954,N_1102,N_3761);
and U6955 (N_6955,N_2919,N_1511);
nor U6956 (N_6956,N_276,N_823);
nand U6957 (N_6957,N_118,N_2469);
nand U6958 (N_6958,N_864,N_1240);
nand U6959 (N_6959,N_2306,N_2625);
nor U6960 (N_6960,N_2579,N_403);
and U6961 (N_6961,N_1960,N_3935);
nand U6962 (N_6962,N_3791,N_915);
or U6963 (N_6963,N_1356,N_1726);
or U6964 (N_6964,N_391,N_2209);
and U6965 (N_6965,N_2507,N_1743);
nor U6966 (N_6966,N_3382,N_3384);
and U6967 (N_6967,N_3691,N_1713);
nor U6968 (N_6968,N_3957,N_2256);
nor U6969 (N_6969,N_436,N_2262);
xnor U6970 (N_6970,N_2625,N_348);
or U6971 (N_6971,N_948,N_3297);
nor U6972 (N_6972,N_3507,N_1328);
and U6973 (N_6973,N_3105,N_1433);
or U6974 (N_6974,N_3252,N_2165);
nand U6975 (N_6975,N_2790,N_1018);
nand U6976 (N_6976,N_2141,N_3561);
nand U6977 (N_6977,N_3837,N_436);
and U6978 (N_6978,N_1102,N_849);
nor U6979 (N_6979,N_1684,N_3640);
and U6980 (N_6980,N_2674,N_420);
xnor U6981 (N_6981,N_3416,N_3286);
nor U6982 (N_6982,N_983,N_1078);
nor U6983 (N_6983,N_1124,N_2961);
nand U6984 (N_6984,N_1727,N_2677);
xor U6985 (N_6985,N_1415,N_2348);
nor U6986 (N_6986,N_96,N_2745);
nand U6987 (N_6987,N_1123,N_2235);
or U6988 (N_6988,N_399,N_3809);
nand U6989 (N_6989,N_2054,N_3232);
or U6990 (N_6990,N_2935,N_422);
nor U6991 (N_6991,N_141,N_3823);
nand U6992 (N_6992,N_2854,N_1584);
nand U6993 (N_6993,N_2212,N_12);
nor U6994 (N_6994,N_32,N_9);
nor U6995 (N_6995,N_2500,N_2067);
nor U6996 (N_6996,N_3585,N_3521);
nand U6997 (N_6997,N_1270,N_1867);
nor U6998 (N_6998,N_3269,N_1333);
xor U6999 (N_6999,N_1300,N_2817);
and U7000 (N_7000,N_3460,N_2130);
xor U7001 (N_7001,N_3712,N_3071);
nand U7002 (N_7002,N_3868,N_1268);
and U7003 (N_7003,N_2507,N_3335);
nor U7004 (N_7004,N_3716,N_1312);
nor U7005 (N_7005,N_3182,N_3392);
nor U7006 (N_7006,N_2694,N_2279);
nor U7007 (N_7007,N_1964,N_2720);
or U7008 (N_7008,N_2269,N_1460);
nor U7009 (N_7009,N_2498,N_1940);
nor U7010 (N_7010,N_848,N_14);
nor U7011 (N_7011,N_2989,N_305);
xor U7012 (N_7012,N_1751,N_2441);
nand U7013 (N_7013,N_270,N_3561);
nor U7014 (N_7014,N_2567,N_1233);
or U7015 (N_7015,N_3887,N_1415);
and U7016 (N_7016,N_1776,N_3412);
or U7017 (N_7017,N_167,N_164);
nor U7018 (N_7018,N_2286,N_1016);
nand U7019 (N_7019,N_1875,N_2343);
xnor U7020 (N_7020,N_1999,N_2620);
and U7021 (N_7021,N_2470,N_2727);
nand U7022 (N_7022,N_648,N_3032);
and U7023 (N_7023,N_2396,N_2859);
nand U7024 (N_7024,N_1826,N_3778);
and U7025 (N_7025,N_3524,N_3303);
or U7026 (N_7026,N_3979,N_1939);
xor U7027 (N_7027,N_963,N_664);
or U7028 (N_7028,N_1771,N_39);
nand U7029 (N_7029,N_300,N_1101);
nand U7030 (N_7030,N_3905,N_2729);
nor U7031 (N_7031,N_2024,N_3995);
and U7032 (N_7032,N_1195,N_129);
or U7033 (N_7033,N_2997,N_1483);
nand U7034 (N_7034,N_2752,N_2849);
xor U7035 (N_7035,N_181,N_2523);
and U7036 (N_7036,N_567,N_125);
and U7037 (N_7037,N_1011,N_1841);
nand U7038 (N_7038,N_1129,N_2821);
or U7039 (N_7039,N_1257,N_1768);
nor U7040 (N_7040,N_3001,N_3859);
nor U7041 (N_7041,N_613,N_2028);
and U7042 (N_7042,N_2666,N_3018);
or U7043 (N_7043,N_1767,N_3596);
nor U7044 (N_7044,N_2349,N_1103);
nor U7045 (N_7045,N_1908,N_1649);
nand U7046 (N_7046,N_2073,N_2100);
or U7047 (N_7047,N_1679,N_2688);
nor U7048 (N_7048,N_3576,N_121);
nand U7049 (N_7049,N_655,N_3272);
nand U7050 (N_7050,N_3640,N_709);
nand U7051 (N_7051,N_3472,N_2860);
or U7052 (N_7052,N_3985,N_3905);
nand U7053 (N_7053,N_1773,N_1463);
xnor U7054 (N_7054,N_3317,N_2245);
and U7055 (N_7055,N_1234,N_2247);
nand U7056 (N_7056,N_1497,N_1475);
and U7057 (N_7057,N_495,N_3430);
nor U7058 (N_7058,N_1069,N_358);
or U7059 (N_7059,N_2621,N_2095);
nor U7060 (N_7060,N_1540,N_774);
xnor U7061 (N_7061,N_1030,N_53);
nand U7062 (N_7062,N_3745,N_1764);
nand U7063 (N_7063,N_2988,N_889);
nor U7064 (N_7064,N_2863,N_3688);
or U7065 (N_7065,N_538,N_1478);
nand U7066 (N_7066,N_1422,N_745);
xor U7067 (N_7067,N_933,N_3812);
nand U7068 (N_7068,N_3354,N_923);
and U7069 (N_7069,N_3828,N_3579);
nor U7070 (N_7070,N_1869,N_2047);
nor U7071 (N_7071,N_1128,N_3554);
and U7072 (N_7072,N_1468,N_1048);
or U7073 (N_7073,N_2608,N_3636);
nor U7074 (N_7074,N_557,N_3232);
or U7075 (N_7075,N_2094,N_1712);
or U7076 (N_7076,N_2750,N_3045);
nor U7077 (N_7077,N_54,N_1384);
or U7078 (N_7078,N_3588,N_1029);
nand U7079 (N_7079,N_2759,N_3472);
xor U7080 (N_7080,N_3150,N_1413);
or U7081 (N_7081,N_3691,N_1197);
nand U7082 (N_7082,N_811,N_1992);
or U7083 (N_7083,N_2225,N_2081);
nor U7084 (N_7084,N_1081,N_3589);
nor U7085 (N_7085,N_452,N_1107);
and U7086 (N_7086,N_221,N_3183);
nor U7087 (N_7087,N_479,N_85);
or U7088 (N_7088,N_171,N_3980);
or U7089 (N_7089,N_487,N_2282);
nand U7090 (N_7090,N_3025,N_3725);
and U7091 (N_7091,N_559,N_1720);
nand U7092 (N_7092,N_2068,N_1063);
xnor U7093 (N_7093,N_93,N_905);
xnor U7094 (N_7094,N_3589,N_3610);
or U7095 (N_7095,N_198,N_3425);
and U7096 (N_7096,N_2056,N_3350);
nand U7097 (N_7097,N_3650,N_1874);
nand U7098 (N_7098,N_306,N_3602);
and U7099 (N_7099,N_2713,N_3769);
nand U7100 (N_7100,N_1033,N_1377);
or U7101 (N_7101,N_3327,N_289);
xnor U7102 (N_7102,N_364,N_3364);
and U7103 (N_7103,N_1798,N_3436);
and U7104 (N_7104,N_1978,N_825);
nor U7105 (N_7105,N_544,N_1179);
or U7106 (N_7106,N_103,N_85);
nand U7107 (N_7107,N_1037,N_729);
or U7108 (N_7108,N_3697,N_959);
xnor U7109 (N_7109,N_3159,N_1776);
nor U7110 (N_7110,N_169,N_2504);
and U7111 (N_7111,N_1707,N_3821);
nor U7112 (N_7112,N_64,N_1787);
xnor U7113 (N_7113,N_818,N_906);
and U7114 (N_7114,N_1711,N_1958);
or U7115 (N_7115,N_3270,N_243);
nand U7116 (N_7116,N_2164,N_1093);
xor U7117 (N_7117,N_3693,N_3881);
nor U7118 (N_7118,N_1140,N_828);
or U7119 (N_7119,N_2571,N_547);
nor U7120 (N_7120,N_2400,N_2829);
and U7121 (N_7121,N_2774,N_2233);
or U7122 (N_7122,N_2466,N_2566);
nor U7123 (N_7123,N_336,N_2575);
and U7124 (N_7124,N_2319,N_914);
xnor U7125 (N_7125,N_1006,N_2469);
nand U7126 (N_7126,N_1085,N_1333);
or U7127 (N_7127,N_638,N_654);
or U7128 (N_7128,N_2236,N_1909);
and U7129 (N_7129,N_1710,N_643);
nand U7130 (N_7130,N_1066,N_3095);
nor U7131 (N_7131,N_526,N_373);
nand U7132 (N_7132,N_3218,N_3121);
xor U7133 (N_7133,N_1376,N_75);
nand U7134 (N_7134,N_612,N_1923);
and U7135 (N_7135,N_2413,N_1461);
and U7136 (N_7136,N_1290,N_1494);
nand U7137 (N_7137,N_1702,N_3393);
nand U7138 (N_7138,N_3377,N_3786);
nand U7139 (N_7139,N_378,N_921);
nor U7140 (N_7140,N_458,N_889);
or U7141 (N_7141,N_616,N_2440);
nor U7142 (N_7142,N_361,N_3236);
nor U7143 (N_7143,N_362,N_3709);
nor U7144 (N_7144,N_2626,N_292);
xnor U7145 (N_7145,N_175,N_3409);
nor U7146 (N_7146,N_2092,N_1350);
or U7147 (N_7147,N_3717,N_2260);
and U7148 (N_7148,N_2604,N_3280);
nor U7149 (N_7149,N_2846,N_2737);
nor U7150 (N_7150,N_3216,N_2212);
nor U7151 (N_7151,N_2189,N_1736);
nor U7152 (N_7152,N_1245,N_1764);
and U7153 (N_7153,N_655,N_1423);
nand U7154 (N_7154,N_3933,N_3640);
or U7155 (N_7155,N_1855,N_1457);
nand U7156 (N_7156,N_1520,N_3051);
and U7157 (N_7157,N_2055,N_1740);
nand U7158 (N_7158,N_627,N_1785);
or U7159 (N_7159,N_552,N_3341);
and U7160 (N_7160,N_463,N_622);
xnor U7161 (N_7161,N_1399,N_161);
nor U7162 (N_7162,N_450,N_1243);
nand U7163 (N_7163,N_1306,N_153);
or U7164 (N_7164,N_801,N_2795);
nand U7165 (N_7165,N_2229,N_2834);
nand U7166 (N_7166,N_363,N_1676);
xnor U7167 (N_7167,N_962,N_3579);
nor U7168 (N_7168,N_36,N_1426);
nand U7169 (N_7169,N_3522,N_3104);
and U7170 (N_7170,N_706,N_2251);
nand U7171 (N_7171,N_1370,N_1979);
xor U7172 (N_7172,N_2607,N_664);
or U7173 (N_7173,N_3914,N_2963);
nand U7174 (N_7174,N_2552,N_2096);
and U7175 (N_7175,N_2690,N_2043);
or U7176 (N_7176,N_2558,N_1999);
and U7177 (N_7177,N_1383,N_36);
nor U7178 (N_7178,N_2261,N_3244);
or U7179 (N_7179,N_1349,N_1266);
nand U7180 (N_7180,N_2951,N_987);
and U7181 (N_7181,N_1610,N_361);
or U7182 (N_7182,N_1832,N_176);
and U7183 (N_7183,N_1388,N_3890);
or U7184 (N_7184,N_2976,N_240);
and U7185 (N_7185,N_2748,N_3425);
nand U7186 (N_7186,N_3092,N_1604);
nor U7187 (N_7187,N_78,N_122);
nand U7188 (N_7188,N_421,N_804);
and U7189 (N_7189,N_3725,N_578);
or U7190 (N_7190,N_1693,N_637);
nor U7191 (N_7191,N_3016,N_986);
nand U7192 (N_7192,N_1292,N_1337);
xor U7193 (N_7193,N_3146,N_2627);
and U7194 (N_7194,N_476,N_1748);
or U7195 (N_7195,N_328,N_3794);
and U7196 (N_7196,N_22,N_3132);
xnor U7197 (N_7197,N_669,N_3535);
or U7198 (N_7198,N_2643,N_960);
nand U7199 (N_7199,N_2513,N_3955);
nor U7200 (N_7200,N_1033,N_2423);
nand U7201 (N_7201,N_2937,N_25);
nand U7202 (N_7202,N_2257,N_136);
and U7203 (N_7203,N_2299,N_3021);
nand U7204 (N_7204,N_2677,N_1040);
nand U7205 (N_7205,N_1705,N_3808);
nand U7206 (N_7206,N_2670,N_3108);
nor U7207 (N_7207,N_2573,N_3612);
and U7208 (N_7208,N_1841,N_456);
and U7209 (N_7209,N_3308,N_1048);
nand U7210 (N_7210,N_3606,N_2740);
nor U7211 (N_7211,N_1866,N_1725);
and U7212 (N_7212,N_3659,N_2243);
and U7213 (N_7213,N_188,N_1324);
and U7214 (N_7214,N_1032,N_1325);
and U7215 (N_7215,N_2400,N_704);
or U7216 (N_7216,N_3603,N_86);
or U7217 (N_7217,N_3549,N_965);
nor U7218 (N_7218,N_56,N_108);
nor U7219 (N_7219,N_2300,N_2885);
xnor U7220 (N_7220,N_3204,N_3711);
or U7221 (N_7221,N_3327,N_595);
nor U7222 (N_7222,N_2488,N_3827);
or U7223 (N_7223,N_637,N_573);
or U7224 (N_7224,N_2886,N_3062);
xor U7225 (N_7225,N_3589,N_3639);
or U7226 (N_7226,N_33,N_109);
nand U7227 (N_7227,N_3512,N_3253);
and U7228 (N_7228,N_2125,N_1128);
nand U7229 (N_7229,N_2688,N_2118);
or U7230 (N_7230,N_360,N_3608);
or U7231 (N_7231,N_2587,N_2253);
nor U7232 (N_7232,N_359,N_2198);
or U7233 (N_7233,N_1900,N_33);
nor U7234 (N_7234,N_613,N_3786);
nor U7235 (N_7235,N_413,N_1921);
or U7236 (N_7236,N_1130,N_2129);
or U7237 (N_7237,N_2147,N_1728);
or U7238 (N_7238,N_714,N_628);
nand U7239 (N_7239,N_1303,N_3665);
and U7240 (N_7240,N_1006,N_1338);
nor U7241 (N_7241,N_3544,N_430);
nor U7242 (N_7242,N_1668,N_1105);
or U7243 (N_7243,N_3077,N_606);
nor U7244 (N_7244,N_3649,N_298);
nor U7245 (N_7245,N_85,N_2980);
or U7246 (N_7246,N_2851,N_3690);
nor U7247 (N_7247,N_3833,N_372);
and U7248 (N_7248,N_3370,N_391);
nand U7249 (N_7249,N_815,N_1324);
nand U7250 (N_7250,N_424,N_260);
or U7251 (N_7251,N_1405,N_898);
nand U7252 (N_7252,N_396,N_2022);
nand U7253 (N_7253,N_3463,N_2055);
nor U7254 (N_7254,N_3454,N_1425);
or U7255 (N_7255,N_1158,N_3495);
or U7256 (N_7256,N_1532,N_2418);
nor U7257 (N_7257,N_3143,N_3660);
or U7258 (N_7258,N_2738,N_3963);
or U7259 (N_7259,N_609,N_1045);
nand U7260 (N_7260,N_3917,N_3066);
or U7261 (N_7261,N_508,N_2605);
or U7262 (N_7262,N_1391,N_3644);
and U7263 (N_7263,N_2629,N_3358);
nor U7264 (N_7264,N_1839,N_1298);
nand U7265 (N_7265,N_1154,N_709);
nor U7266 (N_7266,N_3761,N_2615);
xnor U7267 (N_7267,N_2931,N_1940);
nand U7268 (N_7268,N_2151,N_2934);
or U7269 (N_7269,N_404,N_2629);
nand U7270 (N_7270,N_3606,N_2994);
xor U7271 (N_7271,N_3479,N_2958);
nor U7272 (N_7272,N_2195,N_119);
and U7273 (N_7273,N_1518,N_743);
and U7274 (N_7274,N_2614,N_3025);
nor U7275 (N_7275,N_3065,N_3452);
and U7276 (N_7276,N_1119,N_3350);
nor U7277 (N_7277,N_3767,N_718);
and U7278 (N_7278,N_1411,N_430);
or U7279 (N_7279,N_2236,N_3457);
xnor U7280 (N_7280,N_3079,N_3057);
nand U7281 (N_7281,N_3274,N_719);
nor U7282 (N_7282,N_227,N_1028);
nand U7283 (N_7283,N_1130,N_2395);
nor U7284 (N_7284,N_3670,N_2418);
nand U7285 (N_7285,N_2554,N_3921);
xnor U7286 (N_7286,N_93,N_3871);
nor U7287 (N_7287,N_191,N_278);
nand U7288 (N_7288,N_2253,N_3628);
nand U7289 (N_7289,N_1582,N_2106);
nand U7290 (N_7290,N_2185,N_3022);
and U7291 (N_7291,N_3440,N_2023);
nor U7292 (N_7292,N_1331,N_1370);
or U7293 (N_7293,N_1874,N_932);
nand U7294 (N_7294,N_2679,N_51);
or U7295 (N_7295,N_2894,N_303);
and U7296 (N_7296,N_1655,N_3828);
xor U7297 (N_7297,N_2119,N_969);
nand U7298 (N_7298,N_1250,N_2815);
nor U7299 (N_7299,N_2965,N_1859);
nor U7300 (N_7300,N_1877,N_3053);
nor U7301 (N_7301,N_3744,N_1244);
xor U7302 (N_7302,N_1459,N_1794);
or U7303 (N_7303,N_1776,N_205);
nor U7304 (N_7304,N_2691,N_2584);
xor U7305 (N_7305,N_2073,N_1864);
and U7306 (N_7306,N_1653,N_936);
and U7307 (N_7307,N_418,N_1236);
nand U7308 (N_7308,N_1863,N_3752);
nor U7309 (N_7309,N_102,N_3096);
nand U7310 (N_7310,N_2411,N_2974);
nand U7311 (N_7311,N_920,N_1513);
or U7312 (N_7312,N_1225,N_381);
or U7313 (N_7313,N_1736,N_751);
xnor U7314 (N_7314,N_236,N_3710);
or U7315 (N_7315,N_1945,N_665);
nand U7316 (N_7316,N_3409,N_1404);
and U7317 (N_7317,N_1970,N_3548);
nand U7318 (N_7318,N_3767,N_1023);
and U7319 (N_7319,N_1772,N_3598);
and U7320 (N_7320,N_3753,N_2860);
nand U7321 (N_7321,N_1530,N_2500);
and U7322 (N_7322,N_1884,N_307);
or U7323 (N_7323,N_3455,N_113);
xor U7324 (N_7324,N_1910,N_3734);
or U7325 (N_7325,N_1469,N_2554);
nand U7326 (N_7326,N_1900,N_3945);
xor U7327 (N_7327,N_512,N_700);
nand U7328 (N_7328,N_737,N_2270);
and U7329 (N_7329,N_1506,N_2652);
nor U7330 (N_7330,N_1821,N_2091);
xor U7331 (N_7331,N_1428,N_3606);
or U7332 (N_7332,N_2743,N_2097);
and U7333 (N_7333,N_1529,N_197);
nand U7334 (N_7334,N_150,N_377);
or U7335 (N_7335,N_3640,N_1683);
nand U7336 (N_7336,N_1324,N_603);
nor U7337 (N_7337,N_2274,N_2628);
or U7338 (N_7338,N_3091,N_2545);
or U7339 (N_7339,N_2613,N_2799);
and U7340 (N_7340,N_2378,N_2933);
nor U7341 (N_7341,N_1515,N_3084);
and U7342 (N_7342,N_1083,N_2871);
and U7343 (N_7343,N_593,N_3390);
xnor U7344 (N_7344,N_304,N_1915);
nand U7345 (N_7345,N_563,N_2965);
nor U7346 (N_7346,N_2569,N_2171);
nand U7347 (N_7347,N_578,N_2225);
or U7348 (N_7348,N_2307,N_3782);
nor U7349 (N_7349,N_959,N_8);
nand U7350 (N_7350,N_3350,N_437);
and U7351 (N_7351,N_2983,N_1359);
nand U7352 (N_7352,N_1641,N_2151);
nor U7353 (N_7353,N_305,N_2933);
and U7354 (N_7354,N_975,N_2551);
and U7355 (N_7355,N_1601,N_3944);
nand U7356 (N_7356,N_1327,N_1378);
nor U7357 (N_7357,N_3551,N_832);
nor U7358 (N_7358,N_1343,N_3514);
nand U7359 (N_7359,N_3720,N_2823);
or U7360 (N_7360,N_605,N_2528);
xnor U7361 (N_7361,N_2574,N_396);
xor U7362 (N_7362,N_2943,N_3666);
or U7363 (N_7363,N_1150,N_590);
nor U7364 (N_7364,N_1954,N_1361);
and U7365 (N_7365,N_2828,N_2278);
nor U7366 (N_7366,N_3052,N_1084);
and U7367 (N_7367,N_1139,N_2720);
nor U7368 (N_7368,N_1912,N_1359);
nand U7369 (N_7369,N_2714,N_1302);
and U7370 (N_7370,N_910,N_1782);
and U7371 (N_7371,N_304,N_2932);
or U7372 (N_7372,N_1243,N_2061);
xor U7373 (N_7373,N_1097,N_2329);
or U7374 (N_7374,N_300,N_3424);
nand U7375 (N_7375,N_20,N_2191);
and U7376 (N_7376,N_2031,N_3859);
and U7377 (N_7377,N_831,N_1916);
nor U7378 (N_7378,N_1223,N_611);
and U7379 (N_7379,N_3431,N_3635);
and U7380 (N_7380,N_3494,N_128);
and U7381 (N_7381,N_3573,N_3840);
or U7382 (N_7382,N_3615,N_2793);
or U7383 (N_7383,N_3829,N_3581);
and U7384 (N_7384,N_89,N_2879);
nand U7385 (N_7385,N_2093,N_1278);
nand U7386 (N_7386,N_88,N_2676);
xor U7387 (N_7387,N_1761,N_1097);
or U7388 (N_7388,N_3222,N_3343);
xor U7389 (N_7389,N_2143,N_3040);
and U7390 (N_7390,N_2002,N_1367);
or U7391 (N_7391,N_3333,N_1553);
and U7392 (N_7392,N_1254,N_2270);
nand U7393 (N_7393,N_1125,N_2197);
xor U7394 (N_7394,N_648,N_3609);
nand U7395 (N_7395,N_1501,N_1469);
and U7396 (N_7396,N_353,N_886);
nor U7397 (N_7397,N_3508,N_2442);
and U7398 (N_7398,N_2839,N_1627);
or U7399 (N_7399,N_3197,N_3141);
and U7400 (N_7400,N_3945,N_3629);
nand U7401 (N_7401,N_1546,N_2344);
or U7402 (N_7402,N_3719,N_1211);
or U7403 (N_7403,N_267,N_473);
and U7404 (N_7404,N_2639,N_1588);
or U7405 (N_7405,N_2700,N_3526);
nor U7406 (N_7406,N_2799,N_3154);
and U7407 (N_7407,N_439,N_2842);
or U7408 (N_7408,N_1416,N_954);
nor U7409 (N_7409,N_1119,N_1821);
nand U7410 (N_7410,N_2457,N_3009);
and U7411 (N_7411,N_691,N_2281);
nand U7412 (N_7412,N_2398,N_2651);
nand U7413 (N_7413,N_3240,N_1944);
or U7414 (N_7414,N_1103,N_1431);
nand U7415 (N_7415,N_3756,N_3462);
or U7416 (N_7416,N_2306,N_125);
nor U7417 (N_7417,N_1890,N_1928);
or U7418 (N_7418,N_2698,N_2067);
nor U7419 (N_7419,N_451,N_1513);
and U7420 (N_7420,N_2789,N_3723);
and U7421 (N_7421,N_2580,N_2024);
and U7422 (N_7422,N_237,N_2540);
nor U7423 (N_7423,N_3698,N_3915);
or U7424 (N_7424,N_1892,N_652);
and U7425 (N_7425,N_2487,N_931);
or U7426 (N_7426,N_3808,N_2052);
or U7427 (N_7427,N_3908,N_3588);
nor U7428 (N_7428,N_971,N_567);
or U7429 (N_7429,N_2187,N_3165);
or U7430 (N_7430,N_3536,N_3885);
and U7431 (N_7431,N_1487,N_3936);
nand U7432 (N_7432,N_3670,N_1039);
nand U7433 (N_7433,N_160,N_907);
or U7434 (N_7434,N_3320,N_2443);
and U7435 (N_7435,N_3532,N_1596);
or U7436 (N_7436,N_2902,N_2278);
nand U7437 (N_7437,N_3551,N_2305);
or U7438 (N_7438,N_2424,N_3786);
or U7439 (N_7439,N_1487,N_3146);
nor U7440 (N_7440,N_3387,N_3213);
nor U7441 (N_7441,N_1788,N_182);
or U7442 (N_7442,N_1739,N_2296);
xor U7443 (N_7443,N_1643,N_1836);
or U7444 (N_7444,N_2687,N_1857);
nor U7445 (N_7445,N_95,N_2762);
nor U7446 (N_7446,N_3839,N_3245);
and U7447 (N_7447,N_3688,N_3227);
or U7448 (N_7448,N_1240,N_2618);
nor U7449 (N_7449,N_3921,N_1713);
or U7450 (N_7450,N_213,N_3542);
and U7451 (N_7451,N_887,N_1256);
nor U7452 (N_7452,N_3940,N_600);
xor U7453 (N_7453,N_3767,N_525);
nor U7454 (N_7454,N_3950,N_1707);
or U7455 (N_7455,N_1073,N_2846);
nor U7456 (N_7456,N_3537,N_2288);
and U7457 (N_7457,N_3651,N_3610);
and U7458 (N_7458,N_3708,N_2393);
nor U7459 (N_7459,N_333,N_3887);
nor U7460 (N_7460,N_3974,N_2500);
or U7461 (N_7461,N_2684,N_3839);
nor U7462 (N_7462,N_3148,N_22);
nor U7463 (N_7463,N_1028,N_76);
or U7464 (N_7464,N_2925,N_3622);
nand U7465 (N_7465,N_590,N_3119);
nand U7466 (N_7466,N_931,N_2900);
nor U7467 (N_7467,N_2837,N_2940);
nand U7468 (N_7468,N_2570,N_2752);
nand U7469 (N_7469,N_2130,N_2459);
nor U7470 (N_7470,N_2438,N_2468);
nand U7471 (N_7471,N_1512,N_494);
nor U7472 (N_7472,N_1224,N_3689);
nor U7473 (N_7473,N_1078,N_2795);
or U7474 (N_7474,N_2078,N_1839);
nand U7475 (N_7475,N_3840,N_1135);
nand U7476 (N_7476,N_3846,N_1229);
nand U7477 (N_7477,N_1918,N_2462);
nor U7478 (N_7478,N_3661,N_3695);
nor U7479 (N_7479,N_1684,N_2844);
nand U7480 (N_7480,N_2098,N_2872);
nand U7481 (N_7481,N_2476,N_2182);
nand U7482 (N_7482,N_3155,N_1621);
and U7483 (N_7483,N_1399,N_1832);
or U7484 (N_7484,N_3783,N_3663);
and U7485 (N_7485,N_2933,N_690);
nor U7486 (N_7486,N_3695,N_777);
and U7487 (N_7487,N_655,N_950);
nor U7488 (N_7488,N_779,N_3670);
nor U7489 (N_7489,N_1861,N_12);
nand U7490 (N_7490,N_24,N_3891);
and U7491 (N_7491,N_637,N_246);
or U7492 (N_7492,N_1135,N_2451);
nand U7493 (N_7493,N_2172,N_239);
and U7494 (N_7494,N_812,N_125);
or U7495 (N_7495,N_3428,N_3079);
and U7496 (N_7496,N_836,N_1001);
xnor U7497 (N_7497,N_1279,N_2879);
nor U7498 (N_7498,N_1895,N_653);
and U7499 (N_7499,N_3478,N_376);
or U7500 (N_7500,N_1872,N_1190);
nand U7501 (N_7501,N_3415,N_1910);
xnor U7502 (N_7502,N_698,N_3041);
nand U7503 (N_7503,N_1584,N_2348);
and U7504 (N_7504,N_3301,N_1897);
nor U7505 (N_7505,N_1172,N_3567);
nand U7506 (N_7506,N_3445,N_2984);
nand U7507 (N_7507,N_3928,N_437);
nand U7508 (N_7508,N_3432,N_130);
and U7509 (N_7509,N_3038,N_1481);
xnor U7510 (N_7510,N_3321,N_2062);
and U7511 (N_7511,N_2667,N_1979);
or U7512 (N_7512,N_3441,N_2331);
and U7513 (N_7513,N_3870,N_3);
xnor U7514 (N_7514,N_3124,N_459);
and U7515 (N_7515,N_1742,N_1889);
or U7516 (N_7516,N_792,N_1511);
nand U7517 (N_7517,N_3651,N_1633);
or U7518 (N_7518,N_3873,N_1194);
or U7519 (N_7519,N_2254,N_2660);
nand U7520 (N_7520,N_2034,N_2280);
nand U7521 (N_7521,N_1486,N_2031);
nor U7522 (N_7522,N_3205,N_235);
nor U7523 (N_7523,N_2689,N_1828);
and U7524 (N_7524,N_2575,N_3511);
xor U7525 (N_7525,N_2371,N_515);
or U7526 (N_7526,N_1586,N_1673);
nor U7527 (N_7527,N_1442,N_178);
and U7528 (N_7528,N_3413,N_2854);
and U7529 (N_7529,N_740,N_2895);
and U7530 (N_7530,N_2435,N_515);
xor U7531 (N_7531,N_233,N_1369);
nor U7532 (N_7532,N_1228,N_733);
nand U7533 (N_7533,N_737,N_3306);
xnor U7534 (N_7534,N_346,N_2395);
and U7535 (N_7535,N_244,N_2122);
nand U7536 (N_7536,N_112,N_856);
nor U7537 (N_7537,N_1629,N_1636);
nand U7538 (N_7538,N_706,N_969);
or U7539 (N_7539,N_3871,N_3053);
nand U7540 (N_7540,N_1673,N_2619);
and U7541 (N_7541,N_2398,N_425);
or U7542 (N_7542,N_1668,N_3070);
and U7543 (N_7543,N_3560,N_2755);
or U7544 (N_7544,N_936,N_1781);
nor U7545 (N_7545,N_1912,N_2117);
or U7546 (N_7546,N_2350,N_1442);
or U7547 (N_7547,N_219,N_3824);
and U7548 (N_7548,N_419,N_2203);
nand U7549 (N_7549,N_3831,N_2432);
nand U7550 (N_7550,N_1950,N_3191);
nand U7551 (N_7551,N_367,N_1987);
nor U7552 (N_7552,N_670,N_3227);
nor U7553 (N_7553,N_3255,N_1541);
nor U7554 (N_7554,N_2377,N_2610);
nand U7555 (N_7555,N_1733,N_1167);
nand U7556 (N_7556,N_1903,N_3749);
nor U7557 (N_7557,N_1703,N_2801);
and U7558 (N_7558,N_3335,N_1903);
nand U7559 (N_7559,N_19,N_1037);
xor U7560 (N_7560,N_423,N_756);
or U7561 (N_7561,N_2288,N_3703);
nor U7562 (N_7562,N_2461,N_3200);
and U7563 (N_7563,N_2110,N_1550);
and U7564 (N_7564,N_424,N_3988);
and U7565 (N_7565,N_3377,N_1773);
nand U7566 (N_7566,N_3494,N_101);
or U7567 (N_7567,N_2880,N_516);
or U7568 (N_7568,N_2982,N_3488);
and U7569 (N_7569,N_2174,N_1394);
xor U7570 (N_7570,N_2192,N_3048);
nand U7571 (N_7571,N_319,N_2597);
xnor U7572 (N_7572,N_3187,N_2915);
nand U7573 (N_7573,N_1615,N_1944);
nor U7574 (N_7574,N_3521,N_11);
or U7575 (N_7575,N_1199,N_2513);
or U7576 (N_7576,N_1166,N_3061);
xor U7577 (N_7577,N_105,N_1214);
nor U7578 (N_7578,N_2235,N_652);
and U7579 (N_7579,N_2383,N_1305);
and U7580 (N_7580,N_1643,N_3331);
and U7581 (N_7581,N_2822,N_975);
or U7582 (N_7582,N_177,N_3009);
or U7583 (N_7583,N_1397,N_1825);
nor U7584 (N_7584,N_2481,N_3674);
or U7585 (N_7585,N_3129,N_2243);
nor U7586 (N_7586,N_1324,N_3256);
or U7587 (N_7587,N_2647,N_993);
nor U7588 (N_7588,N_1838,N_3942);
nor U7589 (N_7589,N_462,N_529);
nor U7590 (N_7590,N_1865,N_2267);
or U7591 (N_7591,N_3559,N_2375);
nor U7592 (N_7592,N_1383,N_3584);
nand U7593 (N_7593,N_491,N_1623);
nand U7594 (N_7594,N_975,N_1535);
nand U7595 (N_7595,N_258,N_2788);
and U7596 (N_7596,N_1362,N_2116);
nor U7597 (N_7597,N_3284,N_448);
nand U7598 (N_7598,N_3221,N_2988);
or U7599 (N_7599,N_1980,N_1207);
or U7600 (N_7600,N_226,N_1325);
nand U7601 (N_7601,N_105,N_1447);
and U7602 (N_7602,N_1184,N_909);
nor U7603 (N_7603,N_210,N_951);
or U7604 (N_7604,N_2156,N_2956);
xnor U7605 (N_7605,N_2429,N_3964);
nand U7606 (N_7606,N_2168,N_3617);
nand U7607 (N_7607,N_3787,N_1901);
and U7608 (N_7608,N_434,N_1066);
nor U7609 (N_7609,N_150,N_1595);
or U7610 (N_7610,N_3980,N_3792);
or U7611 (N_7611,N_3315,N_116);
and U7612 (N_7612,N_133,N_3605);
and U7613 (N_7613,N_685,N_2443);
and U7614 (N_7614,N_2469,N_1240);
or U7615 (N_7615,N_2759,N_3329);
nand U7616 (N_7616,N_2996,N_2250);
xor U7617 (N_7617,N_447,N_526);
nor U7618 (N_7618,N_49,N_3097);
nand U7619 (N_7619,N_1190,N_782);
nand U7620 (N_7620,N_3694,N_1191);
or U7621 (N_7621,N_1963,N_2668);
nor U7622 (N_7622,N_2802,N_660);
nor U7623 (N_7623,N_1219,N_42);
nor U7624 (N_7624,N_2111,N_1379);
and U7625 (N_7625,N_1301,N_3908);
nor U7626 (N_7626,N_3371,N_3756);
nand U7627 (N_7627,N_1049,N_1861);
nor U7628 (N_7628,N_461,N_2897);
nor U7629 (N_7629,N_2578,N_3254);
nor U7630 (N_7630,N_3062,N_1815);
nand U7631 (N_7631,N_1452,N_241);
xnor U7632 (N_7632,N_1481,N_1665);
and U7633 (N_7633,N_1347,N_109);
xnor U7634 (N_7634,N_758,N_634);
nor U7635 (N_7635,N_3269,N_3073);
nand U7636 (N_7636,N_545,N_1528);
and U7637 (N_7637,N_2819,N_523);
and U7638 (N_7638,N_91,N_1391);
nand U7639 (N_7639,N_531,N_3030);
or U7640 (N_7640,N_3523,N_1387);
nand U7641 (N_7641,N_454,N_1769);
nor U7642 (N_7642,N_3497,N_1363);
xor U7643 (N_7643,N_1915,N_3068);
nor U7644 (N_7644,N_2884,N_1172);
or U7645 (N_7645,N_1293,N_2443);
and U7646 (N_7646,N_1114,N_3152);
and U7647 (N_7647,N_1822,N_1574);
xor U7648 (N_7648,N_3491,N_1229);
and U7649 (N_7649,N_1774,N_2407);
and U7650 (N_7650,N_2929,N_747);
and U7651 (N_7651,N_2468,N_712);
nor U7652 (N_7652,N_3956,N_3458);
nor U7653 (N_7653,N_346,N_3835);
and U7654 (N_7654,N_3858,N_916);
xnor U7655 (N_7655,N_1193,N_1509);
or U7656 (N_7656,N_1032,N_794);
or U7657 (N_7657,N_1638,N_2354);
nor U7658 (N_7658,N_1089,N_1165);
and U7659 (N_7659,N_934,N_1534);
or U7660 (N_7660,N_506,N_2203);
or U7661 (N_7661,N_1053,N_1061);
or U7662 (N_7662,N_463,N_39);
or U7663 (N_7663,N_1791,N_845);
or U7664 (N_7664,N_3256,N_1758);
or U7665 (N_7665,N_3854,N_3099);
xnor U7666 (N_7666,N_3159,N_3436);
or U7667 (N_7667,N_744,N_3244);
nor U7668 (N_7668,N_825,N_3169);
xor U7669 (N_7669,N_2203,N_479);
and U7670 (N_7670,N_1980,N_3563);
or U7671 (N_7671,N_2244,N_3879);
and U7672 (N_7672,N_1548,N_1620);
or U7673 (N_7673,N_2674,N_3313);
and U7674 (N_7674,N_1264,N_1022);
or U7675 (N_7675,N_1931,N_2090);
and U7676 (N_7676,N_1215,N_3455);
nand U7677 (N_7677,N_3606,N_2815);
or U7678 (N_7678,N_801,N_1636);
or U7679 (N_7679,N_1154,N_3626);
and U7680 (N_7680,N_1747,N_2436);
nand U7681 (N_7681,N_3110,N_1117);
or U7682 (N_7682,N_2080,N_1325);
and U7683 (N_7683,N_1669,N_1454);
or U7684 (N_7684,N_447,N_442);
xnor U7685 (N_7685,N_2748,N_3349);
and U7686 (N_7686,N_2319,N_3946);
nand U7687 (N_7687,N_775,N_3845);
nand U7688 (N_7688,N_504,N_2191);
nor U7689 (N_7689,N_896,N_945);
or U7690 (N_7690,N_857,N_1554);
nand U7691 (N_7691,N_3144,N_190);
nor U7692 (N_7692,N_465,N_3338);
nand U7693 (N_7693,N_868,N_505);
and U7694 (N_7694,N_3097,N_1219);
nor U7695 (N_7695,N_2242,N_3458);
nor U7696 (N_7696,N_2872,N_859);
or U7697 (N_7697,N_2457,N_2635);
or U7698 (N_7698,N_1405,N_2912);
and U7699 (N_7699,N_99,N_2679);
nor U7700 (N_7700,N_3389,N_2153);
and U7701 (N_7701,N_1161,N_2250);
nand U7702 (N_7702,N_3770,N_2000);
nor U7703 (N_7703,N_2060,N_648);
or U7704 (N_7704,N_3448,N_3057);
nor U7705 (N_7705,N_2383,N_2392);
nor U7706 (N_7706,N_3398,N_1943);
and U7707 (N_7707,N_1014,N_646);
nor U7708 (N_7708,N_657,N_980);
nor U7709 (N_7709,N_761,N_83);
and U7710 (N_7710,N_399,N_1921);
nand U7711 (N_7711,N_690,N_857);
nand U7712 (N_7712,N_1197,N_3626);
xnor U7713 (N_7713,N_1680,N_2634);
nand U7714 (N_7714,N_1761,N_2915);
nand U7715 (N_7715,N_2616,N_1308);
xnor U7716 (N_7716,N_1276,N_2234);
or U7717 (N_7717,N_457,N_3328);
and U7718 (N_7718,N_773,N_2882);
or U7719 (N_7719,N_3835,N_1833);
and U7720 (N_7720,N_2211,N_1649);
and U7721 (N_7721,N_1027,N_480);
and U7722 (N_7722,N_728,N_1775);
nor U7723 (N_7723,N_1871,N_2982);
or U7724 (N_7724,N_1871,N_1764);
nor U7725 (N_7725,N_1425,N_481);
xnor U7726 (N_7726,N_3122,N_3419);
nor U7727 (N_7727,N_2953,N_2697);
or U7728 (N_7728,N_3393,N_2077);
or U7729 (N_7729,N_3935,N_2258);
nor U7730 (N_7730,N_2421,N_428);
and U7731 (N_7731,N_1381,N_2414);
nand U7732 (N_7732,N_3059,N_3879);
nand U7733 (N_7733,N_1346,N_2417);
or U7734 (N_7734,N_1730,N_2077);
and U7735 (N_7735,N_2073,N_760);
and U7736 (N_7736,N_744,N_1238);
nand U7737 (N_7737,N_763,N_3955);
and U7738 (N_7738,N_2709,N_2568);
and U7739 (N_7739,N_3059,N_219);
and U7740 (N_7740,N_3097,N_2778);
or U7741 (N_7741,N_2681,N_1815);
nand U7742 (N_7742,N_1318,N_2227);
nand U7743 (N_7743,N_221,N_104);
and U7744 (N_7744,N_1559,N_2378);
nor U7745 (N_7745,N_770,N_3815);
xnor U7746 (N_7746,N_2960,N_862);
or U7747 (N_7747,N_2279,N_295);
nand U7748 (N_7748,N_1921,N_1260);
and U7749 (N_7749,N_2082,N_3433);
and U7750 (N_7750,N_1231,N_2532);
or U7751 (N_7751,N_3607,N_568);
and U7752 (N_7752,N_2377,N_2014);
xnor U7753 (N_7753,N_372,N_1152);
nor U7754 (N_7754,N_3412,N_1645);
and U7755 (N_7755,N_2409,N_1251);
xor U7756 (N_7756,N_2945,N_53);
nand U7757 (N_7757,N_339,N_1314);
xnor U7758 (N_7758,N_1560,N_3602);
or U7759 (N_7759,N_3451,N_3801);
nand U7760 (N_7760,N_1321,N_607);
xnor U7761 (N_7761,N_2778,N_1395);
or U7762 (N_7762,N_700,N_2595);
or U7763 (N_7763,N_818,N_3918);
or U7764 (N_7764,N_1783,N_3133);
or U7765 (N_7765,N_1099,N_87);
and U7766 (N_7766,N_2726,N_3258);
or U7767 (N_7767,N_3698,N_2436);
nand U7768 (N_7768,N_1487,N_94);
and U7769 (N_7769,N_3731,N_3820);
or U7770 (N_7770,N_3976,N_1712);
and U7771 (N_7771,N_654,N_2007);
xor U7772 (N_7772,N_3257,N_506);
xnor U7773 (N_7773,N_820,N_731);
and U7774 (N_7774,N_654,N_3285);
and U7775 (N_7775,N_1667,N_2211);
and U7776 (N_7776,N_674,N_3618);
and U7777 (N_7777,N_355,N_1370);
nor U7778 (N_7778,N_2424,N_3648);
nand U7779 (N_7779,N_2631,N_295);
or U7780 (N_7780,N_1082,N_2520);
or U7781 (N_7781,N_251,N_3416);
and U7782 (N_7782,N_262,N_2486);
and U7783 (N_7783,N_327,N_2777);
nor U7784 (N_7784,N_2550,N_1577);
or U7785 (N_7785,N_1917,N_3886);
or U7786 (N_7786,N_3758,N_2940);
nand U7787 (N_7787,N_2219,N_3491);
nor U7788 (N_7788,N_3914,N_2032);
nor U7789 (N_7789,N_281,N_1935);
nand U7790 (N_7790,N_1644,N_854);
or U7791 (N_7791,N_2289,N_3374);
nor U7792 (N_7792,N_3145,N_3107);
nand U7793 (N_7793,N_2270,N_2500);
nand U7794 (N_7794,N_347,N_670);
nand U7795 (N_7795,N_2568,N_1696);
and U7796 (N_7796,N_130,N_1312);
nand U7797 (N_7797,N_408,N_876);
or U7798 (N_7798,N_3537,N_1275);
and U7799 (N_7799,N_1647,N_3646);
nor U7800 (N_7800,N_1107,N_3366);
nor U7801 (N_7801,N_3183,N_454);
nor U7802 (N_7802,N_2943,N_2978);
or U7803 (N_7803,N_486,N_1725);
and U7804 (N_7804,N_1271,N_3025);
nor U7805 (N_7805,N_563,N_2568);
and U7806 (N_7806,N_660,N_3967);
and U7807 (N_7807,N_2257,N_71);
nand U7808 (N_7808,N_1244,N_1907);
nor U7809 (N_7809,N_3395,N_2261);
or U7810 (N_7810,N_223,N_2804);
or U7811 (N_7811,N_3544,N_3792);
nor U7812 (N_7812,N_231,N_1318);
nand U7813 (N_7813,N_230,N_296);
and U7814 (N_7814,N_1303,N_3645);
nand U7815 (N_7815,N_3779,N_2514);
nand U7816 (N_7816,N_3282,N_970);
and U7817 (N_7817,N_2486,N_3350);
nor U7818 (N_7818,N_817,N_2594);
and U7819 (N_7819,N_2136,N_2235);
and U7820 (N_7820,N_2005,N_3121);
and U7821 (N_7821,N_38,N_2269);
and U7822 (N_7822,N_524,N_205);
nor U7823 (N_7823,N_1061,N_1555);
nor U7824 (N_7824,N_1528,N_3869);
and U7825 (N_7825,N_1960,N_1712);
or U7826 (N_7826,N_2068,N_3859);
or U7827 (N_7827,N_2823,N_2752);
or U7828 (N_7828,N_3573,N_1908);
or U7829 (N_7829,N_1249,N_2586);
or U7830 (N_7830,N_1300,N_3098);
nor U7831 (N_7831,N_961,N_3376);
or U7832 (N_7832,N_2771,N_867);
or U7833 (N_7833,N_2734,N_3176);
nor U7834 (N_7834,N_41,N_9);
nor U7835 (N_7835,N_1532,N_3580);
or U7836 (N_7836,N_3074,N_2913);
or U7837 (N_7837,N_74,N_467);
and U7838 (N_7838,N_1635,N_3905);
and U7839 (N_7839,N_2694,N_3314);
and U7840 (N_7840,N_528,N_1619);
nor U7841 (N_7841,N_2478,N_3296);
and U7842 (N_7842,N_1788,N_2249);
xnor U7843 (N_7843,N_3269,N_1692);
and U7844 (N_7844,N_2421,N_2235);
or U7845 (N_7845,N_734,N_3058);
or U7846 (N_7846,N_1550,N_301);
or U7847 (N_7847,N_1960,N_1411);
nand U7848 (N_7848,N_1195,N_1064);
xor U7849 (N_7849,N_2575,N_3504);
nor U7850 (N_7850,N_897,N_1335);
nand U7851 (N_7851,N_1995,N_3184);
nand U7852 (N_7852,N_2128,N_2487);
and U7853 (N_7853,N_1110,N_2842);
nand U7854 (N_7854,N_1376,N_2153);
or U7855 (N_7855,N_2067,N_708);
nand U7856 (N_7856,N_2701,N_20);
and U7857 (N_7857,N_2647,N_2991);
or U7858 (N_7858,N_828,N_55);
nor U7859 (N_7859,N_3859,N_2350);
xnor U7860 (N_7860,N_847,N_1151);
and U7861 (N_7861,N_3358,N_1101);
and U7862 (N_7862,N_3693,N_3807);
and U7863 (N_7863,N_3317,N_3951);
or U7864 (N_7864,N_2926,N_1551);
or U7865 (N_7865,N_2487,N_2963);
or U7866 (N_7866,N_3531,N_2789);
or U7867 (N_7867,N_2982,N_2845);
or U7868 (N_7868,N_234,N_3339);
xor U7869 (N_7869,N_807,N_2159);
xnor U7870 (N_7870,N_2297,N_3274);
nor U7871 (N_7871,N_2704,N_963);
nor U7872 (N_7872,N_397,N_828);
nand U7873 (N_7873,N_3477,N_391);
nor U7874 (N_7874,N_3749,N_372);
nand U7875 (N_7875,N_3955,N_3437);
nor U7876 (N_7876,N_1143,N_1585);
nand U7877 (N_7877,N_2489,N_2143);
nand U7878 (N_7878,N_3150,N_2348);
nor U7879 (N_7879,N_2306,N_2177);
nand U7880 (N_7880,N_3485,N_368);
and U7881 (N_7881,N_678,N_1648);
xnor U7882 (N_7882,N_3024,N_1928);
nand U7883 (N_7883,N_1229,N_2484);
or U7884 (N_7884,N_2055,N_24);
and U7885 (N_7885,N_1815,N_1549);
nand U7886 (N_7886,N_2292,N_2157);
nand U7887 (N_7887,N_680,N_591);
nand U7888 (N_7888,N_1076,N_2982);
or U7889 (N_7889,N_1029,N_3835);
and U7890 (N_7890,N_3264,N_3556);
and U7891 (N_7891,N_2506,N_2400);
nor U7892 (N_7892,N_3288,N_1748);
nor U7893 (N_7893,N_297,N_3794);
nand U7894 (N_7894,N_2191,N_2348);
and U7895 (N_7895,N_578,N_2848);
and U7896 (N_7896,N_3650,N_699);
xor U7897 (N_7897,N_2605,N_2232);
nor U7898 (N_7898,N_3827,N_2786);
or U7899 (N_7899,N_623,N_1726);
or U7900 (N_7900,N_894,N_928);
nor U7901 (N_7901,N_2775,N_2431);
nand U7902 (N_7902,N_897,N_3194);
nor U7903 (N_7903,N_1974,N_2061);
xor U7904 (N_7904,N_2266,N_2208);
or U7905 (N_7905,N_643,N_3087);
nor U7906 (N_7906,N_3323,N_507);
and U7907 (N_7907,N_2480,N_218);
or U7908 (N_7908,N_3862,N_624);
or U7909 (N_7909,N_3155,N_3779);
nor U7910 (N_7910,N_1557,N_596);
nand U7911 (N_7911,N_948,N_2933);
nor U7912 (N_7912,N_2607,N_1118);
nor U7913 (N_7913,N_1973,N_2133);
nor U7914 (N_7914,N_529,N_3471);
and U7915 (N_7915,N_3715,N_392);
nor U7916 (N_7916,N_3269,N_3079);
and U7917 (N_7917,N_2731,N_498);
nand U7918 (N_7918,N_3086,N_1823);
nand U7919 (N_7919,N_389,N_80);
nor U7920 (N_7920,N_2804,N_3199);
or U7921 (N_7921,N_2442,N_3194);
and U7922 (N_7922,N_875,N_1483);
nor U7923 (N_7923,N_2017,N_2930);
nand U7924 (N_7924,N_1356,N_1316);
and U7925 (N_7925,N_283,N_3716);
nor U7926 (N_7926,N_3923,N_235);
nand U7927 (N_7927,N_641,N_445);
nand U7928 (N_7928,N_3849,N_2052);
nor U7929 (N_7929,N_2307,N_1698);
nor U7930 (N_7930,N_3855,N_717);
nand U7931 (N_7931,N_1075,N_3547);
nand U7932 (N_7932,N_3131,N_1709);
nand U7933 (N_7933,N_806,N_3852);
or U7934 (N_7934,N_1719,N_235);
nand U7935 (N_7935,N_1971,N_3038);
and U7936 (N_7936,N_2700,N_3319);
nand U7937 (N_7937,N_2242,N_3554);
xor U7938 (N_7938,N_2284,N_1248);
and U7939 (N_7939,N_2204,N_2173);
nand U7940 (N_7940,N_2982,N_2596);
and U7941 (N_7941,N_615,N_2221);
nor U7942 (N_7942,N_2100,N_1487);
or U7943 (N_7943,N_186,N_1009);
and U7944 (N_7944,N_1413,N_963);
or U7945 (N_7945,N_321,N_633);
nand U7946 (N_7946,N_1960,N_2368);
nand U7947 (N_7947,N_3900,N_414);
xnor U7948 (N_7948,N_3217,N_1531);
nand U7949 (N_7949,N_879,N_3629);
or U7950 (N_7950,N_1443,N_413);
or U7951 (N_7951,N_3806,N_39);
nand U7952 (N_7952,N_3284,N_3571);
nand U7953 (N_7953,N_1130,N_1131);
nor U7954 (N_7954,N_2363,N_3563);
nand U7955 (N_7955,N_3710,N_1937);
or U7956 (N_7956,N_975,N_801);
nand U7957 (N_7957,N_420,N_2);
nor U7958 (N_7958,N_872,N_451);
or U7959 (N_7959,N_3709,N_1290);
nor U7960 (N_7960,N_1117,N_381);
and U7961 (N_7961,N_3440,N_1467);
and U7962 (N_7962,N_305,N_3866);
nand U7963 (N_7963,N_3719,N_428);
and U7964 (N_7964,N_1307,N_2124);
nor U7965 (N_7965,N_3936,N_1983);
nor U7966 (N_7966,N_2436,N_2002);
and U7967 (N_7967,N_2819,N_1826);
xor U7968 (N_7968,N_340,N_860);
nor U7969 (N_7969,N_759,N_683);
nand U7970 (N_7970,N_2525,N_3288);
or U7971 (N_7971,N_739,N_2417);
nor U7972 (N_7972,N_2677,N_699);
nor U7973 (N_7973,N_1960,N_2677);
xor U7974 (N_7974,N_2323,N_3637);
xnor U7975 (N_7975,N_1536,N_576);
nand U7976 (N_7976,N_3638,N_3266);
nor U7977 (N_7977,N_1567,N_2843);
nand U7978 (N_7978,N_1451,N_1637);
nor U7979 (N_7979,N_2974,N_1077);
or U7980 (N_7980,N_1638,N_3231);
nor U7981 (N_7981,N_697,N_1460);
and U7982 (N_7982,N_926,N_3443);
and U7983 (N_7983,N_2023,N_1273);
or U7984 (N_7984,N_1707,N_3105);
nand U7985 (N_7985,N_3987,N_787);
or U7986 (N_7986,N_806,N_3509);
nor U7987 (N_7987,N_79,N_2041);
xnor U7988 (N_7988,N_395,N_20);
or U7989 (N_7989,N_3576,N_3281);
or U7990 (N_7990,N_1527,N_1649);
nand U7991 (N_7991,N_1019,N_1305);
nor U7992 (N_7992,N_2148,N_1458);
nand U7993 (N_7993,N_995,N_743);
and U7994 (N_7994,N_2655,N_1424);
nor U7995 (N_7995,N_3887,N_1815);
xor U7996 (N_7996,N_366,N_1507);
nand U7997 (N_7997,N_2602,N_3350);
nor U7998 (N_7998,N_1646,N_357);
nand U7999 (N_7999,N_2130,N_896);
xor U8000 (N_8000,N_4727,N_5332);
nand U8001 (N_8001,N_4259,N_5572);
nand U8002 (N_8002,N_7708,N_7140);
nand U8003 (N_8003,N_5219,N_7567);
and U8004 (N_8004,N_6359,N_7644);
xnor U8005 (N_8005,N_5882,N_6943);
nand U8006 (N_8006,N_6516,N_5656);
nand U8007 (N_8007,N_5611,N_4758);
xor U8008 (N_8008,N_4933,N_5166);
or U8009 (N_8009,N_4627,N_6745);
xnor U8010 (N_8010,N_6729,N_4281);
and U8011 (N_8011,N_6555,N_6707);
nor U8012 (N_8012,N_7966,N_4846);
and U8013 (N_8013,N_4269,N_7339);
or U8014 (N_8014,N_4570,N_4887);
and U8015 (N_8015,N_7700,N_4548);
nand U8016 (N_8016,N_6142,N_6891);
or U8017 (N_8017,N_7715,N_5457);
or U8018 (N_8018,N_4728,N_6438);
or U8019 (N_8019,N_5187,N_5379);
and U8020 (N_8020,N_5072,N_6921);
or U8021 (N_8021,N_5136,N_5463);
nor U8022 (N_8022,N_4677,N_6515);
and U8023 (N_8023,N_4113,N_5751);
nor U8024 (N_8024,N_7607,N_7139);
nor U8025 (N_8025,N_6217,N_4990);
or U8026 (N_8026,N_5058,N_7892);
nand U8027 (N_8027,N_7366,N_6846);
or U8028 (N_8028,N_4640,N_4424);
and U8029 (N_8029,N_6650,N_4367);
nand U8030 (N_8030,N_7394,N_7243);
nor U8031 (N_8031,N_6063,N_5631);
nand U8032 (N_8032,N_5423,N_6081);
or U8033 (N_8033,N_7372,N_7904);
and U8034 (N_8034,N_5771,N_7401);
nor U8035 (N_8035,N_5552,N_6839);
or U8036 (N_8036,N_6412,N_7743);
nand U8037 (N_8037,N_6638,N_4089);
xor U8038 (N_8038,N_7436,N_6875);
and U8039 (N_8039,N_6518,N_4106);
and U8040 (N_8040,N_4969,N_7894);
or U8041 (N_8041,N_5180,N_4672);
nor U8042 (N_8042,N_6051,N_4467);
or U8043 (N_8043,N_6461,N_4476);
nand U8044 (N_8044,N_7909,N_5218);
xor U8045 (N_8045,N_6117,N_6273);
or U8046 (N_8046,N_7256,N_6576);
nor U8047 (N_8047,N_4870,N_7374);
nor U8048 (N_8048,N_7963,N_6727);
and U8049 (N_8049,N_5562,N_4218);
and U8050 (N_8050,N_5617,N_4085);
xor U8051 (N_8051,N_5803,N_6353);
nand U8052 (N_8052,N_5723,N_4927);
nor U8053 (N_8053,N_6733,N_7893);
nor U8054 (N_8054,N_6648,N_6199);
and U8055 (N_8055,N_6041,N_7876);
or U8056 (N_8056,N_6102,N_6811);
xnor U8057 (N_8057,N_4357,N_4837);
nand U8058 (N_8058,N_5564,N_5862);
and U8059 (N_8059,N_7674,N_7886);
and U8060 (N_8060,N_6929,N_7479);
and U8061 (N_8061,N_4282,N_5889);
and U8062 (N_8062,N_6378,N_6455);
nor U8063 (N_8063,N_5306,N_6528);
nand U8064 (N_8064,N_4148,N_4434);
nor U8065 (N_8065,N_4585,N_4234);
or U8066 (N_8066,N_6284,N_6252);
nor U8067 (N_8067,N_5814,N_7947);
and U8068 (N_8068,N_6620,N_4690);
nand U8069 (N_8069,N_5436,N_4231);
or U8070 (N_8070,N_6456,N_6385);
or U8071 (N_8071,N_4545,N_7885);
xor U8072 (N_8072,N_6523,N_4670);
nor U8073 (N_8073,N_4723,N_4461);
and U8074 (N_8074,N_6519,N_4201);
nand U8075 (N_8075,N_6077,N_4731);
nor U8076 (N_8076,N_5581,N_4756);
nand U8077 (N_8077,N_6613,N_5311);
nor U8078 (N_8078,N_6094,N_7248);
and U8079 (N_8079,N_4492,N_5856);
nor U8080 (N_8080,N_6469,N_5654);
nand U8081 (N_8081,N_7847,N_7046);
or U8082 (N_8082,N_7203,N_4563);
nand U8083 (N_8083,N_6833,N_6335);
nand U8084 (N_8084,N_6610,N_6828);
or U8085 (N_8085,N_7848,N_4253);
nor U8086 (N_8086,N_7121,N_5874);
and U8087 (N_8087,N_7252,N_7581);
and U8088 (N_8088,N_7433,N_5975);
nor U8089 (N_8089,N_6158,N_5308);
nand U8090 (N_8090,N_7821,N_6192);
or U8091 (N_8091,N_4543,N_7703);
nand U8092 (N_8092,N_7096,N_4918);
or U8093 (N_8093,N_7419,N_7962);
nor U8094 (N_8094,N_5104,N_5259);
nor U8095 (N_8095,N_5150,N_7397);
nor U8096 (N_8096,N_5431,N_7317);
nand U8097 (N_8097,N_4027,N_7450);
or U8098 (N_8098,N_6622,N_4591);
or U8099 (N_8099,N_4811,N_6468);
and U8100 (N_8100,N_5993,N_6511);
nor U8101 (N_8101,N_5710,N_6730);
or U8102 (N_8102,N_7167,N_4354);
nor U8103 (N_8103,N_6577,N_4043);
nor U8104 (N_8104,N_4505,N_5555);
and U8105 (N_8105,N_7437,N_5348);
nor U8106 (N_8106,N_4227,N_4749);
or U8107 (N_8107,N_6358,N_7090);
nor U8108 (N_8108,N_6147,N_5858);
and U8109 (N_8109,N_5094,N_5542);
or U8110 (N_8110,N_4488,N_7679);
or U8111 (N_8111,N_4834,N_6920);
nand U8112 (N_8112,N_6799,N_7763);
and U8113 (N_8113,N_7126,N_7988);
nor U8114 (N_8114,N_7742,N_6782);
nand U8115 (N_8115,N_7497,N_6123);
nand U8116 (N_8116,N_5155,N_5647);
nor U8117 (N_8117,N_7625,N_5984);
xnor U8118 (N_8118,N_4560,N_5076);
or U8119 (N_8119,N_5322,N_7074);
and U8120 (N_8120,N_5604,N_7737);
or U8121 (N_8121,N_6957,N_5794);
nand U8122 (N_8122,N_5454,N_5154);
nor U8123 (N_8123,N_6323,N_6746);
xnor U8124 (N_8124,N_5836,N_5488);
nor U8125 (N_8125,N_4872,N_4735);
nand U8126 (N_8126,N_6661,N_6665);
nor U8127 (N_8127,N_6960,N_5990);
or U8128 (N_8128,N_6763,N_6114);
nor U8129 (N_8129,N_6810,N_5110);
xnor U8130 (N_8130,N_6011,N_7113);
nor U8131 (N_8131,N_6592,N_7949);
nand U8132 (N_8132,N_6067,N_7422);
nand U8133 (N_8133,N_7910,N_4320);
nand U8134 (N_8134,N_5062,N_4150);
and U8135 (N_8135,N_6475,N_5184);
or U8136 (N_8136,N_6531,N_6925);
or U8137 (N_8137,N_6294,N_4378);
nor U8138 (N_8138,N_7758,N_4428);
nor U8139 (N_8139,N_5997,N_5788);
and U8140 (N_8140,N_6495,N_6279);
nor U8141 (N_8141,N_7764,N_5842);
or U8142 (N_8142,N_4348,N_4950);
xor U8143 (N_8143,N_5810,N_6521);
and U8144 (N_8144,N_7722,N_6172);
xor U8145 (N_8145,N_4484,N_7650);
xor U8146 (N_8146,N_6202,N_6107);
and U8147 (N_8147,N_4986,N_4494);
or U8148 (N_8148,N_4205,N_6179);
or U8149 (N_8149,N_7075,N_7373);
xnor U8150 (N_8150,N_7595,N_6243);
nor U8151 (N_8151,N_7311,N_6564);
and U8152 (N_8152,N_5780,N_5355);
or U8153 (N_8153,N_7026,N_6964);
and U8154 (N_8154,N_6429,N_5782);
nor U8155 (N_8155,N_7820,N_5493);
xnor U8156 (N_8156,N_4318,N_7721);
nand U8157 (N_8157,N_4370,N_6291);
nor U8158 (N_8158,N_4911,N_6914);
or U8159 (N_8159,N_7235,N_6220);
xnor U8160 (N_8160,N_5199,N_4557);
and U8161 (N_8161,N_7440,N_5361);
or U8162 (N_8162,N_5805,N_6772);
and U8163 (N_8163,N_6274,N_7453);
or U8164 (N_8164,N_7955,N_6075);
nand U8165 (N_8165,N_4626,N_5663);
and U8166 (N_8166,N_7297,N_7180);
and U8167 (N_8167,N_6022,N_4663);
nand U8168 (N_8168,N_7196,N_5607);
nand U8169 (N_8169,N_6987,N_5586);
nor U8170 (N_8170,N_6227,N_5280);
nor U8171 (N_8171,N_4805,N_4339);
or U8172 (N_8172,N_4708,N_5535);
or U8173 (N_8173,N_5574,N_4779);
nand U8174 (N_8174,N_4130,N_6779);
nor U8175 (N_8175,N_4571,N_6320);
xnor U8176 (N_8176,N_5134,N_4725);
or U8177 (N_8177,N_5050,N_4953);
or U8178 (N_8178,N_7411,N_7699);
or U8179 (N_8179,N_6787,N_4820);
nand U8180 (N_8180,N_5066,N_7669);
or U8181 (N_8181,N_5353,N_5670);
nand U8182 (N_8182,N_7386,N_4510);
xnor U8183 (N_8183,N_5045,N_5823);
xnor U8184 (N_8184,N_5692,N_7534);
or U8185 (N_8185,N_6362,N_7124);
or U8186 (N_8186,N_5445,N_4018);
nand U8187 (N_8187,N_7940,N_7593);
or U8188 (N_8188,N_7670,N_5272);
or U8189 (N_8189,N_4595,N_4399);
and U8190 (N_8190,N_4896,N_5824);
or U8191 (N_8191,N_6853,N_5225);
and U8192 (N_8192,N_4624,N_4272);
nand U8193 (N_8193,N_4458,N_7579);
nor U8194 (N_8194,N_7580,N_6175);
nand U8195 (N_8195,N_6512,N_4246);
and U8196 (N_8196,N_4900,N_4256);
nand U8197 (N_8197,N_6904,N_7059);
nand U8198 (N_8198,N_7620,N_4160);
nor U8199 (N_8199,N_5000,N_6056);
or U8200 (N_8200,N_4120,N_6367);
nor U8201 (N_8201,N_5389,N_4631);
and U8202 (N_8202,N_7563,N_6292);
and U8203 (N_8203,N_5674,N_4766);
nand U8204 (N_8204,N_5662,N_6931);
or U8205 (N_8205,N_7470,N_4744);
nand U8206 (N_8206,N_5783,N_4333);
nor U8207 (N_8207,N_5174,N_6397);
and U8208 (N_8208,N_6024,N_4082);
nor U8209 (N_8209,N_6913,N_5914);
nor U8210 (N_8210,N_4792,N_4610);
nand U8211 (N_8211,N_4014,N_6149);
or U8212 (N_8212,N_5629,N_7467);
and U8213 (N_8213,N_5727,N_6000);
or U8214 (N_8214,N_4981,N_6723);
xor U8215 (N_8215,N_5750,N_6888);
nor U8216 (N_8216,N_7618,N_6491);
xor U8217 (N_8217,N_5244,N_5478);
and U8218 (N_8218,N_7251,N_5636);
and U8219 (N_8219,N_7306,N_4460);
or U8220 (N_8220,N_5729,N_5017);
xnor U8221 (N_8221,N_5525,N_7941);
nand U8222 (N_8222,N_5011,N_4429);
or U8223 (N_8223,N_4643,N_4974);
and U8224 (N_8224,N_6470,N_6735);
nand U8225 (N_8225,N_4678,N_7844);
nand U8226 (N_8226,N_5521,N_4935);
nor U8227 (N_8227,N_4877,N_7056);
and U8228 (N_8228,N_5934,N_5015);
nand U8229 (N_8229,N_6579,N_7521);
and U8230 (N_8230,N_4155,N_7286);
or U8231 (N_8231,N_6448,N_7207);
nand U8232 (N_8232,N_7877,N_7443);
or U8233 (N_8233,N_7514,N_4387);
nor U8234 (N_8234,N_6152,N_4906);
xnor U8235 (N_8235,N_6109,N_6878);
and U8236 (N_8236,N_4891,N_6605);
nor U8237 (N_8237,N_6507,N_4016);
nor U8238 (N_8238,N_4304,N_7690);
or U8239 (N_8239,N_7740,N_6593);
and U8240 (N_8240,N_4258,N_6380);
xor U8241 (N_8241,N_4843,N_4867);
and U8242 (N_8242,N_5440,N_4045);
or U8243 (N_8243,N_7486,N_4451);
xor U8244 (N_8244,N_4369,N_7431);
nand U8245 (N_8245,N_5433,N_5653);
or U8246 (N_8246,N_6601,N_7783);
and U8247 (N_8247,N_6183,N_5452);
nand U8248 (N_8248,N_5693,N_5769);
nand U8249 (N_8249,N_4329,N_7772);
xor U8250 (N_8250,N_7672,N_7184);
nor U8251 (N_8251,N_6406,N_7613);
xnor U8252 (N_8252,N_4868,N_7070);
nor U8253 (N_8253,N_6414,N_5953);
and U8254 (N_8254,N_5917,N_4252);
or U8255 (N_8255,N_7500,N_5964);
nor U8256 (N_8256,N_4902,N_7540);
nor U8257 (N_8257,N_7435,N_7427);
and U8258 (N_8258,N_5981,N_4948);
and U8259 (N_8259,N_7232,N_5561);
or U8260 (N_8260,N_7066,N_6681);
or U8261 (N_8261,N_4733,N_7723);
xor U8262 (N_8262,N_7092,N_5989);
nand U8263 (N_8263,N_4794,N_6127);
nand U8264 (N_8264,N_5969,N_5303);
nand U8265 (N_8265,N_6611,N_7601);
nand U8266 (N_8266,N_7757,N_4815);
and U8267 (N_8267,N_7079,N_5732);
nor U8268 (N_8268,N_4709,N_5132);
nor U8269 (N_8269,N_5667,N_4288);
nor U8270 (N_8270,N_4411,N_4167);
nor U8271 (N_8271,N_6316,N_7418);
or U8272 (N_8272,N_7901,N_4674);
and U8273 (N_8273,N_6234,N_5986);
xor U8274 (N_8274,N_4292,N_4904);
nand U8275 (N_8275,N_5724,N_4736);
nor U8276 (N_8276,N_7466,N_7045);
and U8277 (N_8277,N_6285,N_7314);
and U8278 (N_8278,N_7905,N_5567);
and U8279 (N_8279,N_7028,N_5203);
nand U8280 (N_8280,N_5372,N_7344);
and U8281 (N_8281,N_7770,N_6971);
xnor U8282 (N_8282,N_7602,N_7920);
and U8283 (N_8283,N_4023,N_7388);
nand U8284 (N_8284,N_6485,N_6652);
and U8285 (N_8285,N_7998,N_7819);
nand U8286 (N_8286,N_5888,N_4019);
and U8287 (N_8287,N_5784,N_4004);
nor U8288 (N_8288,N_5241,N_7355);
and U8289 (N_8289,N_4149,N_5140);
and U8290 (N_8290,N_4195,N_6460);
or U8291 (N_8291,N_5164,N_4208);
nor U8292 (N_8292,N_6071,N_5714);
nor U8293 (N_8293,N_4241,N_5296);
nand U8294 (N_8294,N_6629,N_4402);
and U8295 (N_8295,N_7342,N_4053);
or U8296 (N_8296,N_6053,N_5226);
or U8297 (N_8297,N_6118,N_7762);
xor U8298 (N_8298,N_6260,N_4214);
or U8299 (N_8299,N_6831,N_5412);
nor U8300 (N_8300,N_6578,N_5312);
and U8301 (N_8301,N_5143,N_4250);
nand U8302 (N_8302,N_7282,N_5720);
nor U8303 (N_8303,N_6883,N_5301);
and U8304 (N_8304,N_5234,N_5566);
or U8305 (N_8305,N_7425,N_7035);
or U8306 (N_8306,N_6884,N_6843);
nor U8307 (N_8307,N_5991,N_5494);
or U8308 (N_8308,N_6842,N_7768);
nor U8309 (N_8309,N_6841,N_5165);
xnor U8310 (N_8310,N_4912,N_5047);
and U8311 (N_8311,N_7632,N_7993);
or U8312 (N_8312,N_5201,N_7930);
or U8313 (N_8313,N_4928,N_6504);
xor U8314 (N_8314,N_5735,N_4553);
xor U8315 (N_8315,N_4238,N_7089);
or U8316 (N_8316,N_6893,N_4230);
nor U8317 (N_8317,N_7034,N_5923);
or U8318 (N_8318,N_5640,N_4337);
nand U8319 (N_8319,N_4752,N_6349);
or U8320 (N_8320,N_6719,N_5401);
or U8321 (N_8321,N_5338,N_6876);
nand U8322 (N_8322,N_7839,N_6407);
nor U8323 (N_8323,N_7274,N_6825);
or U8324 (N_8324,N_5922,N_5779);
or U8325 (N_8325,N_4580,N_7171);
and U8326 (N_8326,N_6138,N_4831);
and U8327 (N_8327,N_6129,N_5407);
and U8328 (N_8328,N_6662,N_5026);
and U8329 (N_8329,N_5031,N_4539);
nor U8330 (N_8330,N_7211,N_7986);
and U8331 (N_8331,N_7850,N_7189);
or U8332 (N_8332,N_4721,N_4828);
nand U8333 (N_8333,N_6814,N_5868);
nand U8334 (N_8334,N_6027,N_4699);
or U8335 (N_8335,N_4651,N_7493);
or U8336 (N_8336,N_5235,N_4717);
nor U8337 (N_8337,N_5756,N_7649);
or U8338 (N_8338,N_4030,N_5666);
nand U8339 (N_8339,N_6736,N_4943);
and U8340 (N_8340,N_6439,N_7532);
and U8341 (N_8341,N_5686,N_5243);
nor U8342 (N_8342,N_7190,N_4224);
xnor U8343 (N_8343,N_4042,N_6422);
xnor U8344 (N_8344,N_4655,N_4937);
nand U8345 (N_8345,N_5851,N_6326);
nand U8346 (N_8346,N_7350,N_4186);
and U8347 (N_8347,N_4547,N_6386);
nor U8348 (N_8348,N_6757,N_7570);
nand U8349 (N_8349,N_5977,N_4200);
nor U8350 (N_8350,N_7677,N_5876);
or U8351 (N_8351,N_7914,N_4842);
or U8352 (N_8352,N_4894,N_6901);
or U8353 (N_8353,N_6890,N_5119);
nor U8354 (N_8354,N_6715,N_7799);
or U8355 (N_8355,N_6264,N_6098);
and U8356 (N_8356,N_5305,N_4170);
or U8357 (N_8357,N_7400,N_6038);
xor U8358 (N_8358,N_6848,N_4142);
or U8359 (N_8359,N_6144,N_7230);
nand U8360 (N_8360,N_7424,N_6540);
or U8361 (N_8361,N_5787,N_5341);
nor U8362 (N_8362,N_4009,N_4518);
nor U8363 (N_8363,N_6623,N_7329);
nor U8364 (N_8364,N_4884,N_4345);
nand U8365 (N_8365,N_5281,N_7814);
and U8366 (N_8366,N_6031,N_6801);
or U8367 (N_8367,N_5696,N_4261);
and U8368 (N_8368,N_7489,N_4818);
nor U8369 (N_8369,N_5250,N_4131);
nor U8370 (N_8370,N_5786,N_4420);
nand U8371 (N_8371,N_4742,N_7365);
and U8372 (N_8372,N_4930,N_6936);
nor U8373 (N_8373,N_7911,N_6140);
nor U8374 (N_8374,N_6263,N_4295);
or U8375 (N_8375,N_7574,N_4645);
and U8376 (N_8376,N_5485,N_6125);
nor U8377 (N_8377,N_4423,N_6716);
nor U8378 (N_8378,N_4021,N_7392);
or U8379 (N_8379,N_6724,N_4916);
nor U8380 (N_8380,N_5210,N_7343);
or U8381 (N_8381,N_5375,N_6298);
nand U8382 (N_8382,N_7137,N_7865);
nor U8383 (N_8383,N_4477,N_6807);
or U8384 (N_8384,N_4235,N_7875);
and U8385 (N_8385,N_5123,N_4134);
or U8386 (N_8386,N_5253,N_7651);
or U8387 (N_8387,N_4983,N_4632);
nand U8388 (N_8388,N_4101,N_4342);
xnor U8389 (N_8389,N_7064,N_4144);
nor U8390 (N_8390,N_6043,N_4889);
or U8391 (N_8391,N_5288,N_6850);
or U8392 (N_8392,N_7899,N_6411);
nor U8393 (N_8393,N_7362,N_6795);
and U8394 (N_8394,N_7163,N_4715);
xor U8395 (N_8395,N_4438,N_7221);
xnor U8396 (N_8396,N_5852,N_4412);
nor U8397 (N_8397,N_5916,N_4588);
and U8398 (N_8398,N_7114,N_7360);
nor U8399 (N_8399,N_7788,N_5643);
nor U8400 (N_8400,N_4020,N_5726);
nor U8401 (N_8401,N_6995,N_5548);
xnor U8402 (N_8402,N_4642,N_4978);
xor U8403 (N_8403,N_4897,N_6044);
nand U8404 (N_8404,N_5595,N_7145);
or U8405 (N_8405,N_6151,N_7451);
or U8406 (N_8406,N_6200,N_5350);
nor U8407 (N_8407,N_4864,N_6992);
nand U8408 (N_8408,N_5684,N_7827);
nand U8409 (N_8409,N_4844,N_7543);
nand U8410 (N_8410,N_5351,N_5963);
nor U8411 (N_8411,N_7793,N_5825);
and U8412 (N_8412,N_4661,N_5509);
nor U8413 (N_8413,N_7507,N_5685);
nor U8414 (N_8414,N_6539,N_6166);
nand U8415 (N_8415,N_7148,N_5349);
nor U8416 (N_8416,N_5680,N_7193);
and U8417 (N_8417,N_4379,N_4078);
or U8418 (N_8418,N_5483,N_7561);
nor U8419 (N_8419,N_5317,N_4757);
xor U8420 (N_8420,N_4096,N_6953);
or U8421 (N_8421,N_6944,N_5264);
and U8422 (N_8422,N_7741,N_6206);
nor U8423 (N_8423,N_6877,N_7661);
nor U8424 (N_8424,N_6262,N_4255);
nand U8425 (N_8425,N_7659,N_7160);
nand U8426 (N_8426,N_5523,N_4297);
nor U8427 (N_8427,N_4682,N_5419);
and U8428 (N_8428,N_4450,N_5920);
nand U8429 (N_8429,N_4526,N_5554);
xnor U8430 (N_8430,N_5153,N_4776);
nor U8431 (N_8431,N_4762,N_7261);
or U8432 (N_8432,N_4540,N_6281);
or U8433 (N_8433,N_7556,N_5614);
or U8434 (N_8434,N_7597,N_7027);
nor U8435 (N_8435,N_7442,N_4123);
xnor U8436 (N_8436,N_7179,N_7224);
and U8437 (N_8437,N_7849,N_4349);
nand U8438 (N_8438,N_7951,N_4181);
or U8439 (N_8439,N_6947,N_4737);
and U8440 (N_8440,N_5334,N_4895);
nand U8441 (N_8441,N_5775,N_6722);
nor U8442 (N_8442,N_7001,N_5945);
nand U8443 (N_8443,N_5837,N_4503);
nand U8444 (N_8444,N_7313,N_4809);
nor U8445 (N_8445,N_7895,N_4444);
nor U8446 (N_8446,N_5893,N_5829);
or U8447 (N_8447,N_7276,N_6054);
nor U8448 (N_8448,N_6072,N_7859);
and U8449 (N_8449,N_4433,N_5745);
and U8450 (N_8450,N_4069,N_7606);
nor U8451 (N_8451,N_7277,N_4471);
and U8452 (N_8452,N_5755,N_4628);
and U8453 (N_8453,N_7695,N_4139);
nor U8454 (N_8454,N_7665,N_7776);
nand U8455 (N_8455,N_5426,N_7604);
and U8456 (N_8456,N_5757,N_4922);
or U8457 (N_8457,N_4210,N_6889);
xnor U8458 (N_8458,N_4949,N_4194);
nor U8459 (N_8459,N_6136,N_4482);
nor U8460 (N_8460,N_7057,N_6749);
or U8461 (N_8461,N_5507,N_7958);
nand U8462 (N_8462,N_7100,N_4365);
xor U8463 (N_8463,N_6786,N_5499);
nor U8464 (N_8464,N_5875,N_7809);
and U8465 (N_8465,N_6447,N_4513);
or U8466 (N_8466,N_4136,N_6421);
xor U8467 (N_8467,N_4786,N_4747);
nor U8468 (N_8468,N_5282,N_5085);
or U8469 (N_8469,N_7870,N_4984);
nand U8470 (N_8470,N_4913,N_6671);
nor U8471 (N_8471,N_5221,N_4037);
and U8472 (N_8472,N_4070,N_7692);
and U8473 (N_8473,N_6597,N_5496);
nand U8474 (N_8474,N_7278,N_7976);
xnor U8475 (N_8475,N_7959,N_7072);
or U8476 (N_8476,N_5839,N_7291);
nor U8477 (N_8477,N_4855,N_5034);
nor U8478 (N_8478,N_5879,N_6618);
and U8479 (N_8479,N_7950,N_4671);
nor U8480 (N_8480,N_6310,N_6935);
and U8481 (N_8481,N_4940,N_6478);
and U8482 (N_8482,N_5293,N_4022);
and U8483 (N_8483,N_4988,N_4326);
nor U8484 (N_8484,N_7663,N_6951);
and U8485 (N_8485,N_6493,N_4359);
nand U8486 (N_8486,N_5248,N_7073);
nand U8487 (N_8487,N_7609,N_6211);
nor U8488 (N_8488,N_6388,N_5059);
or U8489 (N_8489,N_4172,N_4804);
or U8490 (N_8490,N_7681,N_5952);
or U8491 (N_8491,N_7099,N_5637);
and U8492 (N_8492,N_6402,N_6743);
and U8493 (N_8493,N_4689,N_4088);
or U8494 (N_8494,N_4276,N_5767);
and U8495 (N_8495,N_5596,N_7492);
and U8496 (N_8496,N_7351,N_4781);
nand U8497 (N_8497,N_7880,N_5146);
xor U8498 (N_8498,N_4646,N_7972);
or U8499 (N_8499,N_4457,N_7444);
or U8500 (N_8500,N_4952,N_6905);
nor U8501 (N_8501,N_4473,N_6235);
and U8502 (N_8502,N_7022,N_4388);
and U8503 (N_8503,N_7919,N_5115);
and U8504 (N_8504,N_5133,N_5498);
or U8505 (N_8505,N_6346,N_4609);
or U8506 (N_8506,N_7013,N_5196);
and U8507 (N_8507,N_5690,N_6222);
or U8508 (N_8508,N_5135,N_7214);
nor U8509 (N_8509,N_4803,N_7116);
and U8510 (N_8510,N_5532,N_5247);
or U8511 (N_8511,N_5815,N_7068);
and U8512 (N_8512,N_4569,N_4861);
and U8513 (N_8513,N_5042,N_4619);
nand U8514 (N_8514,N_7104,N_7406);
nor U8515 (N_8515,N_6297,N_4669);
nand U8516 (N_8516,N_5130,N_5772);
and U8517 (N_8517,N_6128,N_5477);
nor U8518 (N_8518,N_6375,N_7780);
nor U8519 (N_8519,N_5216,N_5382);
nand U8520 (N_8520,N_6196,N_5137);
nand U8521 (N_8521,N_6980,N_5954);
or U8522 (N_8522,N_7155,N_7417);
xnor U8523 (N_8523,N_4903,N_7322);
nor U8524 (N_8524,N_5960,N_6695);
xnor U8525 (N_8525,N_7873,N_4615);
nor U8526 (N_8526,N_5678,N_6910);
nor U8527 (N_8527,N_5763,N_6649);
nor U8528 (N_8528,N_6171,N_7295);
nor U8529 (N_8529,N_5028,N_5206);
or U8530 (N_8530,N_5753,N_6974);
nand U8531 (N_8531,N_7903,N_6497);
and U8532 (N_8532,N_6858,N_4611);
nand U8533 (N_8533,N_4858,N_7263);
or U8534 (N_8534,N_6823,N_6173);
or U8535 (N_8535,N_4649,N_7200);
and U8536 (N_8536,N_7071,N_6499);
nor U8537 (N_8537,N_4071,N_7367);
or U8538 (N_8538,N_4386,N_6911);
or U8539 (N_8539,N_6549,N_5005);
nand U8540 (N_8540,N_7594,N_5832);
or U8541 (N_8541,N_6400,N_6619);
and U8542 (N_8542,N_6064,N_7302);
nor U8543 (N_8543,N_4141,N_7348);
xor U8544 (N_8544,N_5327,N_5808);
and U8545 (N_8545,N_7913,N_6633);
nor U8546 (N_8546,N_6721,N_4561);
nor U8547 (N_8547,N_5231,N_7979);
xor U8548 (N_8548,N_5676,N_5309);
nand U8549 (N_8549,N_6948,N_5929);
and U8550 (N_8550,N_5970,N_4520);
and U8551 (N_8551,N_4244,N_6481);
nand U8552 (N_8552,N_6069,N_5537);
nor U8553 (N_8553,N_6741,N_5887);
and U8554 (N_8554,N_7040,N_6463);
nand U8555 (N_8555,N_4327,N_5967);
nand U8556 (N_8556,N_5071,N_6760);
xnor U8557 (N_8557,N_5510,N_7520);
and U8558 (N_8558,N_5682,N_6899);
and U8559 (N_8559,N_6080,N_6443);
nor U8560 (N_8560,N_4633,N_5501);
or U8561 (N_8561,N_7219,N_6258);
or U8562 (N_8562,N_4614,N_7846);
or U8563 (N_8563,N_5869,N_6813);
or U8564 (N_8564,N_5819,N_5845);
or U8565 (N_8565,N_4302,N_5634);
xnor U8566 (N_8566,N_4344,N_6387);
and U8567 (N_8567,N_4777,N_6898);
nand U8568 (N_8568,N_4807,N_5087);
or U8569 (N_8569,N_6986,N_5655);
xnor U8570 (N_8570,N_6712,N_6394);
nor U8571 (N_8571,N_4687,N_7710);
nand U8572 (N_8572,N_7822,N_6486);
nor U8573 (N_8573,N_7050,N_5563);
and U8574 (N_8574,N_4338,N_5343);
xnor U8575 (N_8575,N_4159,N_5592);
nand U8576 (N_8576,N_4446,N_5475);
nand U8577 (N_8577,N_4140,N_6510);
nor U8578 (N_8578,N_7005,N_6886);
or U8579 (N_8579,N_6675,N_5754);
nand U8580 (N_8580,N_6720,N_6557);
and U8581 (N_8581,N_6547,N_5597);
nor U8582 (N_8582,N_5195,N_6120);
nand U8583 (N_8583,N_4350,N_4343);
nand U8584 (N_8584,N_5939,N_5222);
and U8585 (N_8585,N_6690,N_4228);
xor U8586 (N_8586,N_6973,N_7924);
or U8587 (N_8587,N_7455,N_5821);
nor U8588 (N_8588,N_7447,N_6517);
nor U8589 (N_8589,N_6635,N_4376);
nand U8590 (N_8590,N_5816,N_6879);
or U8591 (N_8591,N_5314,N_7791);
or U8592 (N_8592,N_4495,N_5441);
nand U8593 (N_8593,N_7812,N_4966);
xor U8594 (N_8594,N_4886,N_6774);
or U8595 (N_8595,N_7738,N_5202);
nand U8596 (N_8596,N_5764,N_7363);
or U8597 (N_8597,N_4010,N_6410);
xnor U8598 (N_8598,N_4963,N_7458);
or U8599 (N_8599,N_4597,N_7803);
nor U8600 (N_8600,N_7541,N_6972);
xnor U8601 (N_8601,N_7879,N_7942);
nor U8602 (N_8602,N_7310,N_7448);
and U8603 (N_8603,N_5704,N_7107);
nor U8604 (N_8604,N_4145,N_5618);
nor U8605 (N_8605,N_5186,N_7638);
or U8606 (N_8606,N_6568,N_6032);
xnor U8607 (N_8607,N_7257,N_7832);
or U8608 (N_8608,N_5612,N_6266);
and U8609 (N_8609,N_6554,N_5513);
or U8610 (N_8610,N_5943,N_4264);
nor U8611 (N_8611,N_4418,N_7012);
and U8612 (N_8612,N_5051,N_7004);
nand U8613 (N_8613,N_7141,N_5818);
nand U8614 (N_8614,N_4385,N_4915);
or U8615 (N_8615,N_6533,N_6023);
or U8616 (N_8616,N_7616,N_5270);
nor U8617 (N_8617,N_5079,N_5193);
or U8618 (N_8618,N_5739,N_7502);
nor U8619 (N_8619,N_7836,N_6057);
nor U8620 (N_8620,N_4055,N_4286);
nor U8621 (N_8621,N_7020,N_6083);
and U8622 (N_8622,N_6574,N_7385);
xnor U8623 (N_8623,N_7615,N_5886);
and U8624 (N_8624,N_7851,N_4572);
and U8625 (N_8625,N_7575,N_4519);
nor U8626 (N_8626,N_5242,N_5386);
and U8627 (N_8627,N_4033,N_4760);
xnor U8628 (N_8628,N_7739,N_4392);
xor U8629 (N_8629,N_7359,N_4242);
and U8630 (N_8630,N_5149,N_7229);
or U8631 (N_8631,N_5122,N_6740);
nand U8632 (N_8632,N_7003,N_7852);
nor U8633 (N_8633,N_4005,N_6657);
and U8634 (N_8634,N_7749,N_6734);
xor U8635 (N_8635,N_7051,N_5905);
nand U8636 (N_8636,N_7952,N_5330);
or U8637 (N_8637,N_4497,N_7671);
nor U8638 (N_8638,N_7228,N_5204);
or U8639 (N_8639,N_7529,N_6132);
or U8640 (N_8640,N_6867,N_4688);
or U8641 (N_8641,N_5743,N_6857);
and U8642 (N_8642,N_5194,N_5961);
nand U8643 (N_8643,N_5996,N_5070);
nand U8644 (N_8644,N_7460,N_5919);
and U8645 (N_8645,N_4188,N_5473);
nand U8646 (N_8646,N_6203,N_7874);
nor U8647 (N_8647,N_4700,N_6990);
or U8648 (N_8648,N_4448,N_7173);
nor U8649 (N_8649,N_4417,N_4961);
nor U8650 (N_8650,N_4801,N_4932);
nand U8651 (N_8651,N_6546,N_6318);
nor U8652 (N_8652,N_4654,N_7591);
nor U8653 (N_8653,N_4701,N_4233);
nand U8654 (N_8654,N_6017,N_6477);
and U8655 (N_8655,N_5459,N_7463);
xor U8656 (N_8656,N_5752,N_5316);
or U8657 (N_8657,N_5486,N_7519);
or U8658 (N_8658,N_7415,N_5041);
nand U8659 (N_8659,N_6949,N_7735);
nor U8660 (N_8660,N_6494,N_4813);
xor U8661 (N_8661,N_5848,N_7662);
and U8662 (N_8662,N_6703,N_5591);
or U8663 (N_8663,N_6565,N_5329);
nor U8664 (N_8664,N_7202,N_5950);
xor U8665 (N_8665,N_6401,N_7161);
xnor U8666 (N_8666,N_5526,N_5539);
or U8667 (N_8667,N_7571,N_6325);
and U8668 (N_8668,N_4923,N_6253);
or U8669 (N_8669,N_4355,N_7087);
or U8670 (N_8670,N_5575,N_4726);
nand U8671 (N_8671,N_5665,N_5826);
and U8672 (N_8672,N_5176,N_6501);
nor U8673 (N_8673,N_4462,N_5465);
xor U8674 (N_8674,N_7584,N_6324);
and U8675 (N_8675,N_4374,N_4964);
nor U8676 (N_8676,N_4823,N_5476);
nand U8677 (N_8677,N_4664,N_5602);
and U8678 (N_8678,N_7380,N_5101);
nor U8679 (N_8679,N_7935,N_7399);
or U8680 (N_8680,N_4882,N_5116);
nor U8681 (N_8681,N_4135,N_5691);
nand U8682 (N_8682,N_5345,N_5471);
nor U8683 (N_8683,N_5455,N_5453);
nand U8684 (N_8684,N_5318,N_5258);
nand U8685 (N_8685,N_4622,N_5702);
and U8686 (N_8686,N_5627,N_5812);
nor U8687 (N_8687,N_4841,N_7653);
nand U8688 (N_8688,N_6945,N_5622);
xnor U8689 (N_8689,N_6241,N_5291);
nand U8690 (N_8690,N_7340,N_7049);
nor U8691 (N_8691,N_6392,N_6829);
and U8692 (N_8692,N_7298,N_6453);
nand U8693 (N_8693,N_5249,N_7927);
xnor U8694 (N_8694,N_4946,N_5434);
or U8695 (N_8695,N_4934,N_7726);
nor U8696 (N_8696,N_6134,N_7610);
xor U8697 (N_8697,N_7805,N_7376);
nor U8698 (N_8698,N_4171,N_5860);
nand U8699 (N_8699,N_4929,N_5728);
or U8700 (N_8700,N_4732,N_7637);
or U8701 (N_8701,N_4730,N_5551);
nor U8702 (N_8702,N_6299,N_6988);
nand U8703 (N_8703,N_5610,N_5623);
nand U8704 (N_8704,N_5624,N_4408);
xnor U8705 (N_8705,N_7098,N_6639);
or U8706 (N_8706,N_6238,N_4128);
nor U8707 (N_8707,N_6785,N_5001);
nand U8708 (N_8708,N_7775,N_5511);
xnor U8709 (N_8709,N_4791,N_7504);
or U8710 (N_8710,N_7402,N_7513);
nor U8711 (N_8711,N_4802,N_4798);
nand U8712 (N_8712,N_5672,N_7693);
xnor U8713 (N_8713,N_4871,N_7777);
xor U8714 (N_8714,N_5900,N_6216);
nand U8715 (N_8715,N_5012,N_7330);
and U8716 (N_8716,N_7398,N_6465);
or U8717 (N_8717,N_5376,N_7323);
nand U8718 (N_8718,N_5599,N_4278);
nor U8719 (N_8719,N_5645,N_4064);
xnor U8720 (N_8720,N_5360,N_4531);
or U8721 (N_8721,N_7864,N_7128);
or U8722 (N_8722,N_6737,N_7010);
nand U8723 (N_8723,N_4740,N_4093);
and U8724 (N_8724,N_7792,N_4154);
nand U8725 (N_8725,N_4303,N_4782);
and U8726 (N_8726,N_4262,N_5987);
nand U8727 (N_8727,N_4722,N_4602);
nor U8728 (N_8728,N_7206,N_4452);
nor U8729 (N_8729,N_5785,N_4652);
or U8730 (N_8730,N_4771,N_6940);
nand U8731 (N_8731,N_7553,N_5982);
or U8732 (N_8732,N_7969,N_4296);
and U8733 (N_8733,N_4556,N_5082);
and U8734 (N_8734,N_7990,N_7044);
and U8735 (N_8735,N_5962,N_6765);
nor U8736 (N_8736,N_4854,N_5576);
xor U8737 (N_8737,N_7983,N_6288);
or U8738 (N_8738,N_6368,N_5181);
nor U8739 (N_8739,N_4550,N_6003);
and U8740 (N_8740,N_5044,N_5582);
nand U8741 (N_8741,N_4158,N_4552);
or U8742 (N_8742,N_6246,N_5046);
nor U8743 (N_8743,N_5021,N_5108);
and U8744 (N_8744,N_6869,N_7730);
nor U8745 (N_8745,N_4724,N_7352);
nor U8746 (N_8746,N_5942,N_6100);
xnor U8747 (N_8747,N_6305,N_4098);
and U8748 (N_8748,N_4361,N_5883);
nand U8749 (N_8749,N_5438,N_4653);
nand U8750 (N_8750,N_4592,N_7997);
nand U8751 (N_8751,N_6006,N_4100);
nor U8752 (N_8752,N_6520,N_6699);
and U8753 (N_8753,N_6420,N_5141);
nand U8754 (N_8754,N_5859,N_4507);
or U8755 (N_8755,N_7264,N_7621);
and U8756 (N_8756,N_5765,N_6308);
nor U8757 (N_8757,N_6847,N_6781);
and U8758 (N_8758,N_4695,N_4493);
or U8759 (N_8759,N_7569,N_4827);
xnor U8760 (N_8760,N_4586,N_4416);
nand U8761 (N_8761,N_7213,N_7142);
and U8762 (N_8762,N_4351,N_4741);
nand U8763 (N_8763,N_5245,N_5430);
nor U8764 (N_8764,N_4092,N_4251);
nand U8765 (N_8765,N_4185,N_5545);
or U8766 (N_8766,N_7408,N_4504);
nand U8767 (N_8767,N_6626,N_6892);
nand U8768 (N_8768,N_4271,N_7191);
or U8769 (N_8769,N_5553,N_7198);
or U8770 (N_8770,N_5872,N_4017);
nor U8771 (N_8771,N_7186,N_5084);
and U8772 (N_8772,N_7530,N_6933);
nand U8773 (N_8773,N_6537,N_6530);
nor U8774 (N_8774,N_6372,N_4814);
and U8775 (N_8775,N_4713,N_4217);
nor U8776 (N_8776,N_5841,N_7432);
and U8777 (N_8777,N_7957,N_7019);
or U8778 (N_8778,N_7147,N_7943);
and U8779 (N_8779,N_7195,N_4368);
nor U8780 (N_8780,N_7308,N_7041);
nor U8781 (N_8781,N_6427,N_6808);
or U8782 (N_8782,N_7779,N_6121);
xor U8783 (N_8783,N_4353,N_5023);
nor U8784 (N_8784,N_7434,N_6607);
xnor U8785 (N_8785,N_4475,N_7105);
or U8786 (N_8786,N_7108,N_4090);
and U8787 (N_8787,N_6500,N_5271);
or U8788 (N_8788,N_7866,N_5069);
nor U8789 (N_8789,N_7857,N_6340);
nor U8790 (N_8790,N_7552,N_7588);
or U8791 (N_8791,N_6487,N_7817);
xor U8792 (N_8792,N_7731,N_5980);
or U8793 (N_8793,N_7081,N_7259);
nand U8794 (N_8794,N_4879,N_6314);
and U8795 (N_8795,N_5870,N_6268);
nand U8796 (N_8796,N_5362,N_5834);
nand U8797 (N_8797,N_6525,N_7129);
and U8798 (N_8798,N_7109,N_7713);
and U8799 (N_8799,N_4517,N_5238);
nand U8800 (N_8800,N_7215,N_4559);
nand U8801 (N_8801,N_6490,N_5688);
and U8802 (N_8802,N_4321,N_6780);
xnor U8803 (N_8803,N_5408,N_6604);
and U8804 (N_8804,N_4873,N_5804);
nand U8805 (N_8805,N_4048,N_6894);
or U8806 (N_8806,N_7985,N_7590);
xnor U8807 (N_8807,N_5255,N_7389);
nand U8808 (N_8808,N_5651,N_6404);
nor U8809 (N_8809,N_5978,N_5061);
xnor U8810 (N_8810,N_7682,N_5514);
nor U8811 (N_8811,N_4824,N_7527);
nand U8812 (N_8812,N_7292,N_5946);
or U8813 (N_8813,N_4322,N_4826);
nor U8814 (N_8814,N_6015,N_7430);
and U8815 (N_8815,N_4083,N_7897);
nand U8816 (N_8816,N_6742,N_4435);
or U8817 (N_8817,N_6312,N_6963);
nor U8818 (N_8818,N_6625,N_5057);
nor U8819 (N_8819,N_7391,N_7510);
or U8820 (N_8820,N_4529,N_5937);
or U8821 (N_8821,N_7241,N_4711);
or U8822 (N_8822,N_4441,N_5100);
nand U8823 (N_8823,N_5370,N_6676);
nand U8824 (N_8824,N_7216,N_4850);
and U8825 (N_8825,N_6838,N_6508);
nand U8826 (N_8826,N_4996,N_5236);
nand U8827 (N_8827,N_5838,N_7112);
and U8828 (N_8828,N_5971,N_7576);
nor U8829 (N_8829,N_6701,N_7000);
nand U8830 (N_8830,N_4523,N_5416);
nand U8831 (N_8831,N_5106,N_4676);
xor U8832 (N_8832,N_6560,N_5846);
nand U8833 (N_8833,N_7868,N_4917);
nor U8834 (N_8834,N_7729,N_5994);
nor U8835 (N_8835,N_5632,N_6514);
nand U8836 (N_8836,N_6033,N_6163);
nor U8837 (N_8837,N_6384,N_7438);
nor U8838 (N_8838,N_4767,N_4635);
or U8839 (N_8839,N_7890,N_7452);
nor U8840 (N_8840,N_7781,N_7414);
and U8841 (N_8841,N_5027,N_5768);
or U8842 (N_8842,N_5625,N_6393);
and U8843 (N_8843,N_4206,N_6924);
nor U8844 (N_8844,N_6818,N_4275);
or U8845 (N_8845,N_6820,N_5266);
and U8846 (N_8846,N_7908,N_4143);
xor U8847 (N_8847,N_4146,N_6840);
or U8848 (N_8848,N_6021,N_4590);
xor U8849 (N_8849,N_6775,N_5262);
and U8850 (N_8850,N_7021,N_4657);
or U8851 (N_8851,N_4449,N_7039);
and U8852 (N_8852,N_6939,N_5944);
or U8853 (N_8853,N_5009,N_7325);
and U8854 (N_8854,N_4166,N_7756);
nand U8855 (N_8855,N_7766,N_6750);
and U8856 (N_8856,N_5903,N_5791);
or U8857 (N_8857,N_7454,N_4265);
xor U8858 (N_8858,N_7247,N_5256);
xnor U8859 (N_8859,N_4328,N_5613);
xnor U8860 (N_8860,N_6020,N_6553);
or U8861 (N_8861,N_6177,N_6900);
nand U8862 (N_8862,N_6309,N_5725);
nand U8863 (N_8863,N_7837,N_6962);
xnor U8864 (N_8864,N_4783,N_4573);
xnor U8865 (N_8865,N_4491,N_5940);
nor U8866 (N_8866,N_7279,N_6922);
nor U8867 (N_8867,N_4400,N_5850);
nor U8868 (N_8868,N_4898,N_6643);
nand U8869 (N_8869,N_4958,N_7077);
nand U8870 (N_8870,N_4976,N_5687);
nor U8871 (N_8871,N_4191,N_4956);
nand U8872 (N_8872,N_4204,N_5347);
nand U8873 (N_8873,N_6770,N_5365);
or U8874 (N_8874,N_6218,N_5557);
nor U8875 (N_8875,N_4533,N_7572);
xor U8876 (N_8876,N_4052,N_6342);
nand U8877 (N_8877,N_5078,N_4739);
or U8878 (N_8878,N_4860,N_5603);
xnor U8879 (N_8879,N_4836,N_6327);
xnor U8880 (N_8880,N_7354,N_4164);
nand U8881 (N_8881,N_7673,N_4193);
nand U8882 (N_8882,N_7086,N_4347);
nand U8883 (N_8883,N_5861,N_7683);
nand U8884 (N_8884,N_4565,N_6702);
or U8885 (N_8885,N_6860,N_4175);
or U8886 (N_8886,N_6269,N_4888);
nand U8887 (N_8887,N_6205,N_6959);
nand U8888 (N_8888,N_4521,N_6502);
and U8889 (N_8889,N_4769,N_7205);
or U8890 (N_8890,N_6329,N_6265);
nor U8891 (N_8891,N_7646,N_6656);
nand U8892 (N_8892,N_4094,N_6307);
nand U8893 (N_8893,N_6339,N_7746);
nor U8894 (N_8894,N_6197,N_7024);
nand U8895 (N_8895,N_5460,N_6627);
and U8896 (N_8896,N_6513,N_6536);
and U8897 (N_8897,N_4443,N_6827);
nor U8898 (N_8898,N_4907,N_5230);
or U8899 (N_8899,N_7426,N_7387);
nand U8900 (N_8900,N_5336,N_6289);
or U8901 (N_8901,N_6207,N_6219);
nor U8902 (N_8902,N_6642,N_7640);
nor U8903 (N_8903,N_5749,N_7158);
and U8904 (N_8904,N_6573,N_7018);
xor U8905 (N_8905,N_5911,N_6682);
or U8906 (N_8906,N_7138,N_5520);
and U8907 (N_8907,N_6766,N_7307);
or U8908 (N_8908,N_6696,N_6768);
or U8909 (N_8909,N_5733,N_4003);
xnor U8910 (N_8910,N_7926,N_5706);
nand U8911 (N_8911,N_4413,N_4509);
xor U8912 (N_8912,N_4839,N_4317);
nor U8913 (N_8913,N_5326,N_6615);
xnor U8914 (N_8914,N_5801,N_7242);
or U8915 (N_8915,N_7119,N_7944);
or U8916 (N_8916,N_6062,N_5973);
nand U8917 (N_8917,N_7305,N_5462);
xnor U8918 (N_8918,N_7094,N_5506);
and U8919 (N_8919,N_6835,N_5289);
and U8920 (N_8920,N_4397,N_6667);
or U8921 (N_8921,N_6941,N_7091);
nand U8922 (N_8922,N_6492,N_5972);
and U8923 (N_8923,N_5215,N_5500);
nand U8924 (N_8924,N_5921,N_4124);
xor U8925 (N_8925,N_7197,N_4222);
or U8926 (N_8926,N_5867,N_6778);
or U8927 (N_8927,N_7718,N_6287);
nor U8928 (N_8928,N_6655,N_5277);
nor U8929 (N_8929,N_6169,N_4613);
and U8930 (N_8930,N_7111,N_6793);
and U8931 (N_8931,N_7538,N_6503);
or U8932 (N_8932,N_5820,N_5073);
nor U8933 (N_8933,N_4658,N_7813);
nor U8934 (N_8934,N_7697,N_5731);
nor U8935 (N_8935,N_4325,N_7503);
or U8936 (N_8936,N_5188,N_7037);
or U8937 (N_8937,N_4859,N_6159);
or U8938 (N_8938,N_4132,N_5738);
xnor U8939 (N_8939,N_4056,N_7281);
and U8940 (N_8940,N_7181,N_5795);
nor U8941 (N_8941,N_6150,N_4274);
nand U8942 (N_8942,N_6868,N_6673);
or U8943 (N_8943,N_7754,N_7101);
or U8944 (N_8944,N_4656,N_6364);
and U8945 (N_8945,N_7006,N_4395);
and U8946 (N_8946,N_5354,N_7714);
nor U8947 (N_8947,N_5447,N_4581);
or U8948 (N_8948,N_4249,N_5109);
nor U8949 (N_8949,N_7125,N_4031);
and U8950 (N_8950,N_7143,N_7915);
nor U8951 (N_8951,N_4665,N_4968);
and U8952 (N_8952,N_5105,N_6088);
nand U8953 (N_8953,N_5709,N_7378);
and U8954 (N_8954,N_7464,N_4464);
nand U8955 (N_8955,N_5356,N_4971);
nor U8956 (N_8956,N_4987,N_4598);
nand U8957 (N_8957,N_5118,N_7381);
nor U8958 (N_8958,N_4196,N_6694);
or U8959 (N_8959,N_5340,N_5827);
nand U8960 (N_8960,N_5337,N_5559);
nor U8961 (N_8961,N_4780,N_5482);
nor U8962 (N_8962,N_7861,N_7932);
or U8963 (N_8963,N_7301,N_4909);
nand U8964 (N_8964,N_4119,N_4215);
nand U8965 (N_8965,N_5152,N_5588);
and U8966 (N_8966,N_6112,N_7496);
and U8967 (N_8967,N_4202,N_5285);
xor U8968 (N_8968,N_5577,N_4277);
nor U8969 (N_8969,N_6473,N_5522);
xor U8970 (N_8970,N_4755,N_5006);
nor U8971 (N_8971,N_4300,N_5849);
nand U8972 (N_8972,N_4168,N_5126);
and U8973 (N_8973,N_4436,N_6753);
nand U8974 (N_8974,N_7536,N_5037);
or U8975 (N_8975,N_7863,N_4373);
nor U8976 (N_8976,N_6366,N_7872);
and U8977 (N_8977,N_6725,N_6039);
nand U8978 (N_8978,N_6198,N_7154);
and U8979 (N_8979,N_5956,N_5467);
nand U8980 (N_8980,N_5450,N_6283);
nor U8981 (N_8981,N_7537,N_6830);
xnor U8982 (N_8982,N_5516,N_4192);
and U8983 (N_8983,N_7118,N_5405);
nand U8984 (N_8984,N_5448,N_6275);
nor U8985 (N_8985,N_7968,N_6824);
nand U8986 (N_8986,N_5213,N_4383);
nand U8987 (N_8987,N_5609,N_4704);
and U8988 (N_8988,N_7361,N_7883);
xnor U8989 (N_8989,N_7368,N_5144);
nor U8990 (N_8990,N_4502,N_5585);
nand U8991 (N_8991,N_4576,N_4522);
xnor U8992 (N_8992,N_5528,N_5833);
or U8993 (N_8993,N_4138,N_5310);
and U8994 (N_8994,N_7290,N_4593);
or U8995 (N_8995,N_4223,N_6912);
nand U8996 (N_8996,N_5054,N_5112);
or U8997 (N_8997,N_5413,N_7828);
xnor U8998 (N_8998,N_4532,N_7589);
or U8999 (N_8999,N_6663,N_4479);
nand U9000 (N_9000,N_4240,N_6111);
and U9001 (N_9001,N_7995,N_7225);
nand U9002 (N_9002,N_6621,N_7482);
and U9003 (N_9003,N_4079,N_7900);
nand U9004 (N_9004,N_6113,N_5456);
nor U9005 (N_9005,N_4310,N_4880);
and U9006 (N_9006,N_5458,N_6369);
and U9007 (N_9007,N_5935,N_4456);
nor U9008 (N_9008,N_6602,N_5683);
nor U9009 (N_9009,N_6738,N_4439);
nor U9010 (N_9010,N_7316,N_7175);
or U9011 (N_9011,N_7664,N_5828);
or U9012 (N_9012,N_4866,N_7634);
xnor U9013 (N_9013,N_7315,N_5292);
and U9014 (N_9014,N_7159,N_4920);
and U9015 (N_9015,N_4599,N_7146);
nor U9016 (N_9016,N_5113,N_4219);
nor U9017 (N_9017,N_7964,N_6374);
nand U9018 (N_9018,N_6045,N_4180);
and U9019 (N_9019,N_7371,N_7999);
and U9020 (N_9020,N_6398,N_4942);
and U9021 (N_9021,N_6373,N_4483);
or U9022 (N_9022,N_6242,N_7403);
or U9023 (N_9023,N_5161,N_6457);
nand U9024 (N_9024,N_7921,N_5713);
nand U9025 (N_9025,N_4562,N_4486);
nor U9026 (N_9026,N_7918,N_5363);
nor U9027 (N_9027,N_6315,N_7347);
or U9028 (N_9028,N_7312,N_4589);
nand U9029 (N_9029,N_5891,N_6764);
and U9030 (N_9030,N_6548,N_5422);
and U9031 (N_9031,N_7675,N_7237);
nand U9032 (N_9032,N_4032,N_7810);
nor U9033 (N_9033,N_4283,N_5480);
or U9034 (N_9034,N_6377,N_5715);
or U9035 (N_9035,N_6970,N_5573);
and U9036 (N_9036,N_6188,N_6614);
nand U9037 (N_9037,N_6130,N_4468);
nand U9038 (N_9038,N_6035,N_4453);
and U9039 (N_9039,N_5313,N_5484);
xnor U9040 (N_9040,N_7007,N_5364);
nand U9041 (N_9041,N_6066,N_7666);
or U9042 (N_9042,N_6413,N_4177);
xor U9043 (N_9043,N_7287,N_4319);
nor U9044 (N_9044,N_5781,N_4480);
or U9045 (N_9045,N_7807,N_7254);
and U9046 (N_9046,N_5844,N_7840);
or U9047 (N_9047,N_7929,N_7468);
and U9048 (N_9048,N_4830,N_4115);
and U9049 (N_9049,N_5705,N_6226);
or U9050 (N_9050,N_6984,N_5391);
or U9051 (N_9051,N_5089,N_6096);
xor U9052 (N_9052,N_5128,N_5877);
and U9053 (N_9053,N_5616,N_6276);
nand U9054 (N_9054,N_7518,N_7250);
or U9055 (N_9055,N_6459,N_6271);
or U9056 (N_9056,N_4406,N_4285);
and U9057 (N_9057,N_6934,N_7199);
nand U9058 (N_9058,N_5527,N_5855);
or U9059 (N_9059,N_6863,N_5697);
nor U9060 (N_9060,N_7309,N_5556);
nand U9061 (N_9061,N_7227,N_7349);
nor U9062 (N_9062,N_4784,N_4151);
nand U9063 (N_9063,N_7471,N_4381);
nand U9064 (N_9064,N_5162,N_4270);
nor U9065 (N_9065,N_6773,N_4746);
and U9066 (N_9066,N_7273,N_6583);
and U9067 (N_9067,N_7055,N_6257);
xnor U9068 (N_9068,N_6969,N_6849);
nand U9069 (N_9069,N_6110,N_6550);
xnor U9070 (N_9070,N_5179,N_4962);
or U9071 (N_9071,N_6566,N_6822);
nor U9072 (N_9072,N_4869,N_4263);
nand U9073 (N_9073,N_6754,N_6018);
and U9074 (N_9074,N_7333,N_5142);
nand U9075 (N_9075,N_5884,N_7194);
xor U9076 (N_9076,N_6861,N_7624);
xor U9077 (N_9077,N_5958,N_6417);
nand U9078 (N_9078,N_5008,N_4232);
and U9079 (N_9079,N_5621,N_6103);
nor U9080 (N_9080,N_6419,N_4993);
and U9081 (N_9081,N_7320,N_6660);
and U9082 (N_9082,N_6319,N_7887);
and U9083 (N_9083,N_4554,N_5013);
and U9084 (N_9084,N_5223,N_4840);
or U9085 (N_9085,N_7733,N_6007);
nor U9086 (N_9086,N_7201,N_7984);
and U9087 (N_9087,N_4068,N_4706);
nand U9088 (N_9088,N_5495,N_5966);
nand U9089 (N_9089,N_6591,N_6232);
and U9090 (N_9090,N_6333,N_5232);
nor U9091 (N_9091,N_7011,N_4936);
nand U9092 (N_9092,N_4157,N_6155);
and U9093 (N_9093,N_7524,N_5531);
nand U9094 (N_9094,N_5583,N_6382);
nand U9095 (N_9095,N_4380,N_7284);
and U9096 (N_9096,N_4216,N_7896);
and U9097 (N_9097,N_4454,N_6641);
or U9098 (N_9098,N_6646,N_7014);
nor U9099 (N_9099,N_5380,N_6249);
and U9100 (N_9100,N_6798,N_5974);
and U9101 (N_9101,N_6979,N_7752);
nor U9102 (N_9102,N_6376,N_6965);
or U9103 (N_9103,N_6976,N_7226);
nand U9104 (N_9104,N_5504,N_5949);
and U9105 (N_9105,N_7994,N_4705);
or U9106 (N_9106,N_6157,N_4582);
or U9107 (N_9107,N_5695,N_6162);
and U9108 (N_9108,N_6596,N_6852);
nand U9109 (N_9109,N_4273,N_6654);
nand U9110 (N_9110,N_5267,N_7506);
or U9111 (N_9111,N_5742,N_4848);
nor U9112 (N_9112,N_5908,N_5789);
and U9113 (N_9113,N_7745,N_5278);
or U9114 (N_9114,N_4290,N_5056);
or U9115 (N_9115,N_6480,N_4825);
nor U9116 (N_9116,N_4314,N_4555);
nor U9117 (N_9117,N_7614,N_6836);
and U9118 (N_9118,N_4212,N_5979);
nand U9119 (N_9119,N_7928,N_6282);
nor U9120 (N_9120,N_5881,N_7293);
or U9121 (N_9121,N_5524,N_4087);
nor U9122 (N_9122,N_6355,N_4992);
or U9123 (N_9123,N_4761,N_7244);
nand U9124 (N_9124,N_4883,N_4558);
nand U9125 (N_9125,N_4965,N_7578);
nand U9126 (N_9126,N_7728,N_4012);
xnor U9127 (N_9127,N_7657,N_7054);
and U9128 (N_9128,N_6084,N_5721);
or U9129 (N_9129,N_4459,N_7560);
xor U9130 (N_9130,N_6685,N_7168);
or U9131 (N_9131,N_6304,N_7619);
and U9132 (N_9132,N_4335,N_7223);
xnor U9133 (N_9133,N_7508,N_4372);
nand U9134 (N_9134,N_7946,N_7583);
or U9135 (N_9135,N_5065,N_5442);
and U9136 (N_9136,N_5570,N_4364);
nand U9137 (N_9137,N_4315,N_6999);
nor U9138 (N_9138,N_6185,N_5002);
nor U9139 (N_9139,N_7465,N_4046);
nand U9140 (N_9140,N_6688,N_4084);
and U9141 (N_9141,N_6535,N_4189);
and U9142 (N_9142,N_4544,N_4332);
or U9143 (N_9143,N_4394,N_4881);
nor U9144 (N_9144,N_7691,N_4178);
nand U9145 (N_9145,N_5747,N_7906);
and U9146 (N_9146,N_4541,N_5208);
or U9147 (N_9147,N_6871,N_4680);
nand U9148 (N_9148,N_5549,N_6225);
and U9149 (N_9149,N_7639,N_6726);
nor U9150 (N_9150,N_6761,N_7794);
and U9151 (N_9151,N_7156,N_7795);
and U9152 (N_9152,N_7067,N_6896);
or U9153 (N_9153,N_6148,N_7727);
and U9154 (N_9154,N_7299,N_6446);
nand U9155 (N_9155,N_7331,N_7088);
or U9156 (N_9156,N_6371,N_6005);
and U9157 (N_9157,N_6278,N_5220);
nand U9158 (N_9158,N_4515,N_5840);
nor U9159 (N_9159,N_5025,N_6049);
and U9160 (N_9160,N_5315,N_7480);
and U9161 (N_9161,N_7599,N_4899);
and U9162 (N_9162,N_5543,N_4163);
or U9163 (N_9163,N_5766,N_6628);
nor U9164 (N_9164,N_6409,N_6001);
xor U9165 (N_9165,N_4247,N_5157);
or U9166 (N_9166,N_4061,N_7992);
and U9167 (N_9167,N_5871,N_6239);
or U9168 (N_9168,N_6630,N_7680);
nand U9169 (N_9169,N_4197,N_6937);
or U9170 (N_9170,N_5807,N_6013);
and U9171 (N_9171,N_7771,N_6010);
xor U9172 (N_9172,N_6290,N_4977);
nand U9173 (N_9173,N_6058,N_4183);
and U9174 (N_9174,N_5287,N_6416);
nor U9175 (N_9175,N_6082,N_7262);
nor U9176 (N_9176,N_6631,N_4600);
and U9177 (N_9177,N_4773,N_5403);
and U9178 (N_9178,N_6357,N_5205);
nor U9179 (N_9179,N_7782,N_6684);
or U9180 (N_9180,N_7798,N_5040);
or U9181 (N_9181,N_6060,N_5394);
or U9182 (N_9182,N_5778,N_4578);
xor U9183 (N_9183,N_7258,N_6441);
nand U9184 (N_9184,N_5959,N_6866);
or U9185 (N_9185,N_5560,N_6710);
nand U9186 (N_9186,N_7353,N_4182);
nor U9187 (N_9187,N_4024,N_5470);
xnor U9188 (N_9188,N_7925,N_7592);
xor U9189 (N_9189,N_7218,N_7642);
nand U9190 (N_9190,N_7856,N_5254);
nor U9191 (N_9191,N_6612,N_6352);
and U9192 (N_9192,N_4324,N_5601);
nand U9193 (N_9193,N_7755,N_7265);
and U9194 (N_9194,N_6311,N_5381);
and U9195 (N_9195,N_6137,N_5269);
and U9196 (N_9196,N_6581,N_4073);
nor U9197 (N_9197,N_4220,N_6791);
and U9198 (N_9198,N_4745,N_6215);
or U9199 (N_9199,N_5092,N_6488);
and U9200 (N_9200,N_7853,N_5661);
nor U9201 (N_9201,N_5429,N_7939);
nand U9202 (N_9202,N_7975,N_6028);
and U9203 (N_9203,N_6777,N_4336);
nor U9204 (N_9204,N_4694,N_6433);
or U9205 (N_9205,N_4810,N_5831);
nor U9206 (N_9206,N_7475,N_5968);
nand U9207 (N_9207,N_7267,N_6361);
nand U9208 (N_9208,N_4051,N_5103);
and U9209 (N_9209,N_4209,N_5547);
nor U9210 (N_9210,N_6603,N_4041);
or U9211 (N_9211,N_4793,N_4306);
and U9212 (N_9212,N_5594,N_4954);
nor U9213 (N_9213,N_4371,N_5897);
or U9214 (N_9214,N_4577,N_7499);
nand U9215 (N_9215,N_7725,N_7058);
or U9216 (N_9216,N_6440,N_7157);
nand U9217 (N_9217,N_6034,N_4077);
nand U9218 (N_9218,N_6758,N_7334);
or U9219 (N_9219,N_7808,N_4490);
xnor U9220 (N_9220,N_5049,N_5064);
or U9221 (N_9221,N_6804,N_4179);
and U9222 (N_9222,N_7236,N_4284);
nor U9223 (N_9223,N_4914,N_6788);
and U9224 (N_9224,N_6958,N_6016);
xor U9225 (N_9225,N_7834,N_7517);
and U9226 (N_9226,N_7421,N_4567);
nand U9227 (N_9227,N_6594,N_6370);
and U9228 (N_9228,N_7405,N_4617);
nor U9229 (N_9229,N_6087,N_5402);
or U9230 (N_9230,N_5265,N_6167);
nor U9231 (N_9231,N_7174,N_7523);
nand U9232 (N_9232,N_7582,N_4111);
nand U9233 (N_9233,N_5497,N_6551);
or U9234 (N_9234,N_6932,N_5320);
nand U9235 (N_9235,N_4865,N_5156);
or U9236 (N_9236,N_7182,N_6143);
nand U9237 (N_9237,N_7177,N_6844);
nand U9238 (N_9238,N_4396,N_5016);
nor U9239 (N_9239,N_5650,N_4445);
or U9240 (N_9240,N_6408,N_4684);
or U9241 (N_9241,N_4161,N_5529);
nand U9242 (N_9242,N_5229,N_7608);
or U9243 (N_9243,N_6918,N_5373);
or U9244 (N_9244,N_5505,N_4957);
or U9245 (N_9245,N_4301,N_6930);
xor U9246 (N_9246,N_6651,N_5928);
or U9247 (N_9247,N_4579,N_4584);
nor U9248 (N_9248,N_7240,N_5608);
or U9249 (N_9249,N_5406,N_5098);
or U9250 (N_9250,N_7130,N_4207);
nor U9251 (N_9251,N_6099,N_5159);
nor U9252 (N_9252,N_6569,N_4662);
or U9253 (N_9253,N_6012,N_6796);
or U9254 (N_9254,N_5035,N_6391);
nor U9255 (N_9255,N_4778,N_7558);
and U9256 (N_9256,N_4691,N_4346);
or U9257 (N_9257,N_7512,N_5748);
nand U9258 (N_9258,N_4989,N_4312);
and U9259 (N_9259,N_4426,N_7790);
or U9260 (N_9260,N_5633,N_5446);
or U9261 (N_9261,N_5227,N_4062);
nand U9262 (N_9262,N_5734,N_7888);
or U9263 (N_9263,N_7631,N_7170);
nor U9264 (N_9264,N_6418,N_5830);
or U9265 (N_9265,N_6975,N_7210);
nor U9266 (N_9266,N_6670,N_7289);
nand U9267 (N_9267,N_4710,N_4876);
and U9268 (N_9268,N_7255,N_4422);
and U9269 (N_9269,N_6078,N_7357);
and U9270 (N_9270,N_4137,N_6789);
nand U9271 (N_9271,N_4718,N_4401);
xor U9272 (N_9272,N_4266,N_5224);
nand U9273 (N_9273,N_7636,N_4905);
and U9274 (N_9274,N_7551,N_5642);
and U9275 (N_9275,N_5411,N_5290);
or U9276 (N_9276,N_7327,N_6991);
nor U9277 (N_9277,N_6434,N_6728);
xnor U9278 (N_9278,N_5550,N_5163);
nor U9279 (N_9279,N_5813,N_6698);
or U9280 (N_9280,N_7383,N_6425);
nand U9281 (N_9281,N_5138,N_7498);
xnor U9282 (N_9282,N_6541,N_6002);
nor U9283 (N_9283,N_5410,N_4243);
or U9284 (N_9284,N_4432,N_7938);
or U9285 (N_9285,N_4384,N_5864);
nor U9286 (N_9286,N_4118,N_7036);
and U9287 (N_9287,N_5806,N_5125);
xor U9288 (N_9288,N_4542,N_7823);
and U9289 (N_9289,N_7596,N_7153);
or U9290 (N_9290,N_4692,N_4129);
nand U9291 (N_9291,N_5770,N_5936);
nor U9292 (N_9292,N_7319,N_7420);
nor U9293 (N_9293,N_6767,N_5626);
nor U9294 (N_9294,N_7526,N_4608);
nor U9295 (N_9295,N_7009,N_7283);
or U9296 (N_9296,N_4686,N_4673);
nand U9297 (N_9297,N_5298,N_6803);
and U9298 (N_9298,N_4036,N_5580);
nor U9299 (N_9299,N_7786,N_5240);
xnor U9300 (N_9300,N_5907,N_4110);
and U9301 (N_9301,N_4546,N_7577);
or U9302 (N_9302,N_5530,N_5668);
and U9303 (N_9303,N_4551,N_4994);
or U9304 (N_9304,N_5652,N_5022);
nand U9305 (N_9305,N_7231,N_4893);
and U9306 (N_9306,N_4716,N_6762);
and U9307 (N_9307,N_5880,N_7623);
and U9308 (N_9308,N_4765,N_6328);
nor U9309 (N_9309,N_4975,N_4951);
xnor U9310 (N_9310,N_4667,N_6037);
nor U9311 (N_9311,N_6244,N_7390);
or U9312 (N_9312,N_7931,N_7626);
nand U9313 (N_9313,N_6496,N_7063);
or U9314 (N_9314,N_6708,N_5420);
nor U9315 (N_9315,N_7869,N_5544);
and U9316 (N_9316,N_6691,N_5948);
nand U9317 (N_9317,N_6221,N_6711);
nand U9318 (N_9318,N_6479,N_7449);
xnor U9319 (N_9319,N_5191,N_7858);
and U9320 (N_9320,N_5374,N_5449);
nor U9321 (N_9321,N_4772,N_5716);
and U9322 (N_9322,N_5182,N_7961);
or U9323 (N_9323,N_7884,N_4979);
and U9324 (N_9324,N_4162,N_4356);
and U9325 (N_9325,N_5777,N_6025);
xor U9326 (N_9326,N_5811,N_5983);
and U9327 (N_9327,N_7668,N_7222);
and U9328 (N_9328,N_4623,N_4574);
nor U9329 (N_9329,N_4427,N_6351);
nand U9330 (N_9330,N_7395,N_6821);
and U9331 (N_9331,N_5121,N_6870);
xnor U9332 (N_9332,N_4685,N_5466);
or U9333 (N_9333,N_6231,N_6632);
or U9334 (N_9334,N_6178,N_6209);
or U9335 (N_9335,N_5717,N_6952);
nor U9336 (N_9336,N_4910,N_5007);
nand U9337 (N_9337,N_5024,N_7660);
xnor U9338 (N_9338,N_6070,N_7825);
nand U9339 (N_9339,N_7369,N_5331);
or U9340 (N_9340,N_6092,N_7472);
xnor U9341 (N_9341,N_5912,N_6509);
nand U9342 (N_9342,N_4245,N_5335);
nor U9343 (N_9343,N_5578,N_4596);
nor U9344 (N_9344,N_5707,N_4362);
xnor U9345 (N_9345,N_6683,N_6395);
nand U9346 (N_9346,N_6859,N_6575);
nand U9347 (N_9347,N_4638,N_4806);
or U9348 (N_9348,N_4799,N_5885);
or U9349 (N_9349,N_4751,N_7544);
nor U9350 (N_9350,N_6306,N_7384);
nor U9351 (N_9351,N_5600,N_7612);
or U9352 (N_9352,N_7702,N_6193);
nor U9353 (N_9353,N_4616,N_4437);
nand U9354 (N_9354,N_7550,N_5048);
and U9355 (N_9355,N_4714,N_4506);
nand U9356 (N_9356,N_4156,N_6036);
xnor U9357 (N_9357,N_7212,N_7629);
and U9358 (N_9358,N_5114,N_6059);
xor U9359 (N_9359,N_6802,N_4257);
xnor U9360 (N_9360,N_7600,N_7627);
or U9361 (N_9361,N_4607,N_6484);
nand U9362 (N_9362,N_5865,N_7937);
nor U9363 (N_9363,N_7136,N_6587);
and U9364 (N_9364,N_7062,N_6522);
and U9365 (N_9365,N_7882,N_4187);
and U9366 (N_9366,N_4738,N_7542);
nand U9367 (N_9367,N_4299,N_5644);
or U9368 (N_9368,N_6996,N_6806);
or U9369 (N_9369,N_7488,N_6527);
nor U9370 (N_9370,N_7382,N_5947);
and U9371 (N_9371,N_6718,N_5774);
nand U9372 (N_9372,N_5926,N_6348);
or U9373 (N_9373,N_6115,N_4229);
and U9374 (N_9374,N_6462,N_6139);
or U9375 (N_9375,N_6435,N_5352);
or U9376 (N_9376,N_7838,N_7989);
xor U9377 (N_9377,N_4763,N_7706);
nor U9378 (N_9378,N_5300,N_6048);
nor U9379 (N_9379,N_6106,N_7667);
and U9380 (N_9380,N_4109,N_5396);
and U9381 (N_9381,N_7133,N_4213);
nor U9382 (N_9382,N_6090,N_4999);
or U9383 (N_9383,N_4080,N_4489);
nor U9384 (N_9384,N_5736,N_4298);
or U9385 (N_9385,N_7732,N_5020);
nand U9386 (N_9386,N_6783,N_4291);
nand U9387 (N_9387,N_5719,N_6181);
nand U9388 (N_9388,N_6526,N_5606);
nor U9389 (N_9389,N_7676,N_4647);
xor U9390 (N_9390,N_6245,N_5927);
nand U9391 (N_9391,N_5086,N_6534);
or U9392 (N_9392,N_4309,N_6097);
or U9393 (N_9393,N_4496,N_7169);
nand U9394 (N_9394,N_6559,N_4352);
and U9395 (N_9395,N_4703,N_7052);
or U9396 (N_9396,N_7548,N_4985);
or U9397 (N_9397,N_6322,N_7647);
nor U9398 (N_9398,N_6363,N_5091);
nor U9399 (N_9399,N_7336,N_7473);
and U9400 (N_9400,N_4039,N_6415);
nand U9401 (N_9401,N_6666,N_5339);
nand U9402 (N_9402,N_5357,N_5404);
and U9403 (N_9403,N_4660,N_6050);
or U9404 (N_9404,N_6771,N_4605);
nand U9405 (N_9405,N_5399,N_6332);
nand U9406 (N_9406,N_6259,N_6954);
and U9407 (N_9407,N_5131,N_5400);
or U9408 (N_9408,N_4409,N_4107);
or U9409 (N_9409,N_5835,N_4313);
nor U9410 (N_9410,N_6968,N_6145);
nor U9411 (N_9411,N_4485,N_5209);
xnor U9412 (N_9412,N_7635,N_4849);
and U9413 (N_9413,N_7686,N_6552);
and U9414 (N_9414,N_5798,N_4279);
xor U9415 (N_9415,N_7078,N_7871);
nand U9416 (N_9416,N_5519,N_6608);
nor U9417 (N_9417,N_5955,N_5189);
and U9418 (N_9418,N_7948,N_7446);
and U9419 (N_9419,N_6856,N_4501);
nand U9420 (N_9420,N_4478,N_6301);
or U9421 (N_9421,N_4712,N_6168);
xnor U9422 (N_9422,N_5129,N_4174);
nand U9423 (N_9423,N_7328,N_5635);
or U9424 (N_9424,N_6029,N_4527);
and U9425 (N_9425,N_7239,N_5664);
or U9426 (N_9426,N_5925,N_5233);
or U9427 (N_9427,N_4693,N_7912);
nand U9428 (N_9428,N_6689,N_7796);
or U9429 (N_9429,N_6704,N_5649);
and U9430 (N_9430,N_5171,N_4764);
or U9431 (N_9431,N_5797,N_6343);
nand U9432 (N_9432,N_6692,N_7338);
and U9433 (N_9433,N_5741,N_5207);
nor U9434 (N_9434,N_6201,N_5392);
nand U9435 (N_9435,N_6769,N_6381);
or U9436 (N_9436,N_4097,N_5368);
xor U9437 (N_9437,N_7061,N_7187);
and U9438 (N_9438,N_7643,N_6161);
nor U9439 (N_9439,N_5605,N_7818);
xor U9440 (N_9440,N_6270,N_6942);
xor U9441 (N_9441,N_7300,N_7784);
nand U9442 (N_9442,N_6874,N_5906);
and U9443 (N_9443,N_7528,N_5894);
nor U9444 (N_9444,N_6981,N_7015);
xnor U9445 (N_9445,N_6653,N_5902);
or U9446 (N_9446,N_5708,N_6624);
and U9447 (N_9447,N_5451,N_6474);
and U9448 (N_9448,N_4057,N_4973);
or U9449 (N_9449,N_7185,N_5324);
nor U9450 (N_9450,N_5638,N_4516);
or U9451 (N_9451,N_6472,N_6267);
or U9452 (N_9452,N_5160,N_6705);
nor U9453 (N_9453,N_5197,N_7103);
or U9454 (N_9454,N_4650,N_7833);
or U9455 (N_9455,N_4237,N_7164);
nand U9456 (N_9456,N_7982,N_5252);
nor U9457 (N_9457,N_6588,N_6214);
xor U9458 (N_9458,N_6296,N_6817);
nand U9459 (N_9459,N_5565,N_4221);
and U9460 (N_9460,N_4176,N_7641);
and U9461 (N_9461,N_5759,N_6677);
and U9462 (N_9462,N_5915,N_4116);
nand U9463 (N_9463,N_6317,N_6994);
nor U9464 (N_9464,N_5491,N_5145);
nor U9465 (N_9465,N_4528,N_5437);
nand U9466 (N_9466,N_5415,N_4125);
xor U9467 (N_9467,N_7268,N_4955);
nor U9468 (N_9468,N_5890,N_7889);
nor U9469 (N_9469,N_7748,N_7761);
nor U9470 (N_9470,N_5043,N_6909);
or U9471 (N_9471,N_7843,N_5127);
nor U9472 (N_9472,N_6189,N_4702);
and U9473 (N_9473,N_6816,N_4498);
nand U9474 (N_9474,N_4360,N_6634);
and U9475 (N_9475,N_7960,N_4612);
and U9476 (N_9476,N_4759,N_7083);
or U9477 (N_9477,N_6669,N_6706);
xnor U9478 (N_9478,N_7622,N_6585);
and U9479 (N_9479,N_7204,N_7209);
or U9480 (N_9480,N_7304,N_7337);
nand U9481 (N_9481,N_4774,N_6466);
xnor U9482 (N_9482,N_7953,N_7802);
or U9483 (N_9483,N_7474,N_5395);
nor U9484 (N_9484,N_6668,N_5425);
nor U9485 (N_9485,N_4549,N_5383);
nand U9486 (N_9486,N_6230,N_7370);
and U9487 (N_9487,N_7253,N_5297);
nor U9488 (N_9488,N_6165,N_7428);
nand U9489 (N_9489,N_7689,N_6731);
nor U9490 (N_9490,N_5060,N_5080);
nor U9491 (N_9491,N_4307,N_6887);
nand U9492 (N_9492,N_5487,N_6116);
xor U9493 (N_9493,N_6105,N_6826);
nand U9494 (N_9494,N_7016,N_7445);
and U9495 (N_9495,N_4112,N_7272);
nor U9496 (N_9496,N_4863,N_5873);
and U9497 (N_9497,N_7294,N_7654);
nor U9498 (N_9498,N_5904,N_7656);
nor U9499 (N_9499,N_4636,N_7867);
nand U9500 (N_9500,N_4028,N_5646);
nor U9501 (N_9501,N_5590,N_7902);
and U9502 (N_9502,N_5283,N_5502);
nand U9503 (N_9503,N_7152,N_7410);
nor U9504 (N_9504,N_5276,N_4268);
and U9505 (N_9505,N_5328,N_5409);
and U9506 (N_9506,N_5481,N_4465);
nand U9507 (N_9507,N_4817,N_4239);
nand U9508 (N_9508,N_7778,N_6586);
xnor U9509 (N_9509,N_4025,N_5398);
nor U9510 (N_9510,N_4407,N_7701);
xnor U9511 (N_9511,N_6895,N_7565);
xor U9512 (N_9512,N_5081,N_4874);
nor U9513 (N_9513,N_4583,N_5469);
and U9514 (N_9514,N_6908,N_5677);
and U9515 (N_9515,N_7716,N_6153);
nand U9516 (N_9516,N_7285,N_5843);
nor U9517 (N_9517,N_6009,N_4707);
or U9518 (N_9518,N_7981,N_4466);
and U9519 (N_9519,N_7535,N_5799);
or U9520 (N_9520,N_7484,N_5468);
nor U9521 (N_9521,N_6104,N_7135);
nor U9522 (N_9522,N_5075,N_7605);
or U9523 (N_9523,N_5648,N_7318);
xnor U9524 (N_9524,N_4038,N_4153);
nand U9525 (N_9525,N_5090,N_6837);
and U9526 (N_9526,N_6247,N_4566);
nor U9527 (N_9527,N_7760,N_5718);
nor U9528 (N_9528,N_6208,N_6119);
nand U9529 (N_9529,N_6748,N_5461);
nor U9530 (N_9530,N_5117,N_4890);
or U9531 (N_9531,N_5302,N_7102);
and U9532 (N_9532,N_6277,N_4511);
or U9533 (N_9533,N_6977,N_7547);
and U9534 (N_9534,N_6693,N_7767);
or U9535 (N_9535,N_6792,N_5170);
nor U9536 (N_9536,N_6897,N_7509);
or U9537 (N_9537,N_4499,N_7495);
or U9538 (N_9538,N_5055,N_7974);
or U9539 (N_9539,N_7973,N_7144);
or U9540 (N_9540,N_6356,N_7165);
or U9541 (N_9541,N_4040,N_6482);
nor U9542 (N_9542,N_6606,N_7658);
or U9543 (N_9543,N_5183,N_5995);
or U9544 (N_9544,N_6679,N_5367);
or U9545 (N_9545,N_5930,N_4081);
or U9546 (N_9546,N_5965,N_4065);
or U9547 (N_9547,N_4008,N_5102);
nor U9548 (N_9548,N_7841,N_5992);
nand U9549 (N_9549,N_4341,N_6182);
and U9550 (N_9550,N_4000,N_6709);
or U9551 (N_9551,N_6739,N_5711);
nor U9552 (N_9552,N_5895,N_6154);
nor U9553 (N_9553,N_7860,N_6341);
and U9554 (N_9554,N_7712,N_5295);
nand U9555 (N_9555,N_5032,N_7967);
nor U9556 (N_9556,N_6752,N_6832);
nor U9557 (N_9557,N_6647,N_4788);
nor U9558 (N_9558,N_6061,N_6580);
xor U9559 (N_9559,N_7516,N_4358);
and U9560 (N_9560,N_6233,N_4404);
or U9561 (N_9561,N_6645,N_6095);
or U9562 (N_9562,N_7704,N_6664);
or U9563 (N_9563,N_5924,N_5211);
or U9564 (N_9564,N_4625,N_6584);
nand U9565 (N_9565,N_6336,N_4618);
nor U9566 (N_9566,N_5941,N_4630);
and U9567 (N_9567,N_6524,N_7774);
nor U9568 (N_9568,N_6347,N_7991);
nand U9569 (N_9569,N_7645,N_6700);
xor U9570 (N_9570,N_4856,N_5346);
or U9571 (N_9571,N_4821,N_7377);
or U9572 (N_9572,N_7603,N_6544);
nor U9573 (N_9573,N_4442,N_5515);
nor U9574 (N_9574,N_6186,N_6567);
and U9575 (N_9575,N_6570,N_6133);
or U9576 (N_9576,N_7151,N_6089);
nor U9577 (N_9577,N_7132,N_4537);
xor U9578 (N_9578,N_5951,N_5699);
nand U9579 (N_9579,N_4001,N_7724);
nand U9580 (N_9580,N_7801,N_6982);
and U9581 (N_9581,N_6800,N_7687);
and U9582 (N_9582,N_7800,N_5237);
or U9583 (N_9583,N_7891,N_6236);
or U9584 (N_9584,N_4419,N_7719);
nand U9585 (N_9585,N_6956,N_7717);
xor U9586 (N_9586,N_7980,N_6915);
and U9587 (N_9587,N_7804,N_4248);
nor U9588 (N_9588,N_5200,N_6194);
nand U9589 (N_9589,N_4203,N_4921);
nand U9590 (N_9590,N_5307,N_7546);
and U9591 (N_9591,N_7375,N_7842);
xnor U9592 (N_9592,N_6126,N_6989);
or U9593 (N_9593,N_4481,N_5077);
or U9594 (N_9594,N_6180,N_7652);
nand U9595 (N_9595,N_7696,N_4829);
or U9596 (N_9596,N_5673,N_4931);
and U9597 (N_9597,N_5107,N_4901);
nand U9598 (N_9598,N_4852,N_7478);
or U9599 (N_9599,N_6483,N_6538);
nand U9600 (N_9600,N_5030,N_6756);
nand U9601 (N_9601,N_5268,N_6251);
and U9602 (N_9602,N_7811,N_4440);
or U9603 (N_9603,N_4822,N_6946);
xor U9604 (N_9604,N_5658,N_6834);
nor U9605 (N_9605,N_4066,N_7707);
or U9606 (N_9606,N_7076,N_6644);
and U9607 (N_9607,N_5003,N_7945);
and U9608 (N_9608,N_5866,N_5260);
and U9609 (N_9609,N_6445,N_4970);
xor U9610 (N_9610,N_4800,N_6240);
and U9611 (N_9611,N_4939,N_5172);
and U9612 (N_9612,N_4058,N_4011);
nor U9613 (N_9613,N_7476,N_6255);
nor U9614 (N_9614,N_6250,N_4851);
xor U9615 (N_9615,N_4389,N_7238);
nor U9616 (N_9616,N_4514,N_4331);
or U9617 (N_9617,N_6141,N_7789);
nand U9618 (N_9618,N_4775,N_7271);
or U9619 (N_9619,N_4748,N_4564);
and U9620 (N_9620,N_7043,N_7501);
nand U9621 (N_9621,N_4659,N_7549);
nor U9622 (N_9622,N_7720,N_4960);
or U9623 (N_9623,N_6091,N_6019);
nand U9624 (N_9624,N_5414,N_5737);
and U9625 (N_9625,N_5901,N_5938);
and U9626 (N_9626,N_6819,N_4538);
nor U9627 (N_9627,N_7970,N_7162);
nor U9628 (N_9628,N_7407,N_6755);
or U9629 (N_9629,N_7845,N_5088);
nand U9630 (N_9630,N_6164,N_6437);
or U9631 (N_9631,N_6983,N_6405);
xnor U9632 (N_9632,N_4878,N_4305);
or U9633 (N_9633,N_4853,N_6101);
nand U9634 (N_9634,N_4512,N_5809);
nor U9635 (N_9635,N_4603,N_5004);
and U9636 (N_9636,N_5540,N_4924);
nand U9637 (N_9637,N_6423,N_7023);
xnor U9638 (N_9638,N_7192,N_5998);
or U9639 (N_9639,N_7346,N_7047);
nor U9640 (N_9640,N_6903,N_7996);
and U9641 (N_9641,N_5933,N_5173);
and U9642 (N_9642,N_5615,N_5111);
xnor U9643 (N_9643,N_4833,N_4165);
or U9644 (N_9644,N_6637,N_4114);
nand U9645 (N_9645,N_7573,N_4199);
and U9646 (N_9646,N_7332,N_4425);
and U9647 (N_9647,N_4734,N_4431);
or U9648 (N_9648,N_5639,N_7123);
and U9649 (N_9649,N_6224,N_4393);
nor U9650 (N_9650,N_4254,N_5571);
or U9651 (N_9651,N_4049,N_6428);
and U9652 (N_9652,N_5854,N_4838);
or U9653 (N_9653,N_5558,N_5294);
and U9654 (N_9654,N_7934,N_7759);
and U9655 (N_9655,N_5036,N_5899);
and U9656 (N_9656,N_7245,N_4832);
or U9657 (N_9657,N_5722,N_4982);
or U9658 (N_9658,N_7555,N_5730);
or U9659 (N_9659,N_5701,N_6345);
xnor U9660 (N_9660,N_4390,N_4972);
nand U9661 (N_9661,N_4797,N_6916);
or U9662 (N_9662,N_4015,N_5342);
or U9663 (N_9663,N_7477,N_6672);
nand U9664 (N_9664,N_5097,N_5417);
nand U9665 (N_9665,N_4108,N_6430);
or U9666 (N_9666,N_7522,N_6074);
or U9667 (N_9667,N_6506,N_7633);
nor U9668 (N_9668,N_7303,N_5773);
nand U9669 (N_9669,N_4363,N_7965);
and U9670 (N_9670,N_7404,N_4054);
or U9671 (N_9671,N_7736,N_6213);
or U9672 (N_9672,N_5378,N_6571);
or U9673 (N_9673,N_6658,N_6156);
nor U9674 (N_9674,N_4743,N_4267);
or U9675 (N_9675,N_4067,N_5217);
and U9676 (N_9676,N_5358,N_4455);
and U9677 (N_9677,N_7335,N_6321);
nand U9678 (N_9678,N_5304,N_6851);
and U9679 (N_9679,N_6790,N_7031);
and U9680 (N_9680,N_5178,N_7917);
or U9681 (N_9681,N_6334,N_6449);
nand U9682 (N_9682,N_7233,N_7461);
nor U9683 (N_9683,N_7183,N_4639);
nor U9684 (N_9684,N_7246,N_4280);
nor U9685 (N_9685,N_6146,N_5177);
nor U9686 (N_9686,N_5790,N_4819);
and U9687 (N_9687,N_4414,N_5039);
or U9688 (N_9688,N_7188,N_7288);
nand U9689 (N_9689,N_5279,N_7483);
or U9690 (N_9690,N_6873,N_7296);
nand U9691 (N_9691,N_5641,N_5988);
nand U9692 (N_9692,N_7586,N_5068);
and U9693 (N_9693,N_7085,N_4925);
or U9694 (N_9694,N_5052,N_5010);
nand U9695 (N_9695,N_7491,N_7106);
xnor U9696 (N_9696,N_6674,N_4536);
or U9697 (N_9697,N_6365,N_7630);
or U9698 (N_9698,N_4857,N_4885);
nor U9699 (N_9699,N_6476,N_5393);
or U9700 (N_9700,N_7688,N_6885);
nand U9701 (N_9701,N_6451,N_7916);
nand U9702 (N_9702,N_5286,N_6498);
xnor U9703 (N_9703,N_6135,N_6784);
nor U9704 (N_9704,N_6184,N_5909);
xor U9705 (N_9705,N_6617,N_4330);
nor U9706 (N_9706,N_7462,N_6450);
nand U9707 (N_9707,N_7678,N_6004);
nor U9708 (N_9708,N_7816,N_5479);
nor U9709 (N_9709,N_6598,N_6085);
or U9710 (N_9710,N_4629,N_7456);
xnor U9711 (N_9711,N_7038,N_4184);
nor U9712 (N_9712,N_4190,N_5444);
or U9713 (N_9713,N_4050,N_7709);
nand U9714 (N_9714,N_6572,N_7648);
and U9715 (N_9715,N_7806,N_6997);
nor U9716 (N_9716,N_4719,N_7533);
and U9717 (N_9717,N_5175,N_6582);
nand U9718 (N_9718,N_7266,N_4997);
nand U9719 (N_9719,N_5681,N_4754);
and U9720 (N_9720,N_4847,N_7280);
nor U9721 (N_9721,N_5761,N_5014);
nand U9722 (N_9722,N_5120,N_4875);
xnor U9723 (N_9723,N_5167,N_5019);
nor U9724 (N_9724,N_5472,N_6906);
nor U9725 (N_9725,N_7379,N_5096);
nor U9726 (N_9726,N_7824,N_4500);
xnor U9727 (N_9727,N_7459,N_7554);
and U9728 (N_9728,N_7545,N_4575);
nor U9729 (N_9729,N_6040,N_6505);
and U9730 (N_9730,N_7511,N_4035);
and U9731 (N_9731,N_6350,N_7326);
nor U9732 (N_9732,N_4919,N_7409);
nand U9733 (N_9733,N_6086,N_4060);
and U9734 (N_9734,N_7131,N_7082);
nor U9735 (N_9735,N_6424,N_4316);
or U9736 (N_9736,N_4621,N_6174);
xor U9737 (N_9737,N_6237,N_5802);
nand U9738 (N_9738,N_4472,N_7977);
nor U9739 (N_9739,N_6008,N_4681);
nand U9740 (N_9740,N_5325,N_4091);
and U9741 (N_9741,N_6797,N_7830);
nor U9742 (N_9742,N_5359,N_7032);
and U9743 (N_9743,N_7878,N_6776);
nor U9744 (N_9744,N_6872,N_7562);
nand U9745 (N_9745,N_4606,N_7956);
nor U9746 (N_9746,N_7978,N_5489);
and U9747 (N_9747,N_5148,N_5212);
and U9748 (N_9748,N_5246,N_6383);
or U9749 (N_9749,N_4812,N_4323);
nand U9750 (N_9750,N_5139,N_7127);
nand U9751 (N_9751,N_4675,N_7166);
or U9752 (N_9752,N_5384,N_7413);
xor U9753 (N_9753,N_6489,N_4013);
nand U9754 (N_9754,N_5533,N_6640);
nand U9755 (N_9755,N_5976,N_4044);
nor U9756 (N_9756,N_5538,N_7923);
nor U9757 (N_9757,N_7734,N_6923);
or U9758 (N_9758,N_5421,N_4026);
nand U9759 (N_9759,N_7341,N_7773);
nand U9760 (N_9760,N_4998,N_4377);
or U9761 (N_9761,N_4698,N_6978);
or U9762 (N_9762,N_7907,N_5593);
nand U9763 (N_9763,N_4398,N_7208);
nand U9764 (N_9764,N_6927,N_6014);
nor U9765 (N_9765,N_5660,N_5239);
or U9766 (N_9766,N_4991,N_4926);
or U9767 (N_9767,N_5228,N_7008);
or U9768 (N_9768,N_4666,N_6902);
nand U9769 (N_9769,N_5512,N_4289);
and U9770 (N_9770,N_4007,N_6170);
or U9771 (N_9771,N_4121,N_7080);
nand U9772 (N_9772,N_6442,N_7617);
nor U9773 (N_9773,N_7698,N_7611);
and U9774 (N_9774,N_4808,N_4594);
nand U9775 (N_9775,N_6295,N_7269);
xnor U9776 (N_9776,N_5067,N_4770);
and U9777 (N_9777,N_4366,N_6042);
xnor U9778 (N_9778,N_5299,N_4789);
nand U9779 (N_9779,N_7797,N_6805);
and U9780 (N_9780,N_5263,N_6313);
xor U9781 (N_9781,N_5857,N_4535);
nand U9782 (N_9782,N_6176,N_4430);
or U9783 (N_9783,N_5418,N_6680);
nor U9784 (N_9784,N_4720,N_4099);
xnor U9785 (N_9785,N_5712,N_7439);
or U9786 (N_9786,N_5169,N_6543);
nand U9787 (N_9787,N_5147,N_5397);
nand U9788 (N_9788,N_5366,N_4474);
or U9789 (N_9789,N_7971,N_5957);
or U9790 (N_9790,N_7628,N_4696);
and U9791 (N_9791,N_6881,N_4967);
nand U9792 (N_9792,N_5371,N_7120);
nor U9793 (N_9793,N_5541,N_7769);
and U9794 (N_9794,N_6390,N_6261);
nor U9795 (N_9795,N_6928,N_7744);
or U9796 (N_9796,N_4102,N_5863);
nor U9797 (N_9797,N_4908,N_4104);
or U9798 (N_9798,N_4508,N_6195);
nand U9799 (N_9799,N_7441,N_4375);
nand U9800 (N_9800,N_7220,N_6678);
nand U9801 (N_9801,N_5251,N_4340);
or U9802 (N_9802,N_6812,N_4308);
xor U9803 (N_9803,N_6330,N_6254);
xor U9804 (N_9804,N_6880,N_7396);
nor U9805 (N_9805,N_5534,N_6815);
nand U9806 (N_9806,N_6542,N_5569);
and U9807 (N_9807,N_4648,N_6600);
or U9808 (N_9808,N_7685,N_6300);
and U9809 (N_9809,N_7364,N_5587);
or U9810 (N_9810,N_6204,N_7122);
nor U9811 (N_9811,N_7069,N_6432);
nor U9812 (N_9812,N_5675,N_4421);
and U9813 (N_9813,N_5932,N_7393);
nand U9814 (N_9814,N_6855,N_7093);
nand U9815 (N_9815,N_7249,N_6338);
or U9816 (N_9816,N_6337,N_5918);
nor U9817 (N_9817,N_6131,N_5033);
and U9818 (N_9818,N_7345,N_7564);
nand U9819 (N_9819,N_7017,N_5443);
and U9820 (N_9820,N_7481,N_6055);
nor U9821 (N_9821,N_4620,N_5931);
or U9822 (N_9822,N_4787,N_7149);
xnor U9823 (N_9823,N_5659,N_6073);
or U9824 (N_9824,N_4076,N_6862);
and U9825 (N_9825,N_6458,N_5896);
and U9826 (N_9826,N_6030,N_5124);
nand U9827 (N_9827,N_5158,N_6845);
nor U9828 (N_9828,N_5185,N_5760);
and U9829 (N_9829,N_7178,N_6065);
nor U9830 (N_9830,N_7826,N_7933);
and U9831 (N_9831,N_4403,N_5598);
and U9832 (N_9832,N_5390,N_6079);
nand U9833 (N_9833,N_5261,N_5619);
xnor U9834 (N_9834,N_6223,N_5018);
or U9835 (N_9835,N_5892,N_7557);
or U9836 (N_9836,N_5053,N_5698);
or U9837 (N_9837,N_5792,N_5474);
nor U9838 (N_9838,N_4063,N_6950);
and U9839 (N_9839,N_7084,N_6471);
nand U9840 (N_9840,N_5385,N_4086);
nand U9841 (N_9841,N_7829,N_6454);
or U9842 (N_9842,N_4862,N_4072);
nor U9843 (N_9843,N_4945,N_6431);
xnor U9844 (N_9844,N_5274,N_5198);
nor U9845 (N_9845,N_7115,N_7150);
nand U9846 (N_9846,N_7324,N_7705);
and U9847 (N_9847,N_4391,N_4470);
or U9848 (N_9848,N_6190,N_4644);
nor U9849 (N_9849,N_6713,N_7065);
nor U9850 (N_9850,N_5424,N_5700);
nor U9851 (N_9851,N_7566,N_4785);
and U9852 (N_9852,N_7275,N_6272);
and U9853 (N_9853,N_4029,N_6403);
nor U9854 (N_9854,N_6590,N_7270);
or U9855 (N_9855,N_5377,N_7423);
nor U9856 (N_9856,N_5628,N_6938);
nand U9857 (N_9857,N_6751,N_4683);
nand U9858 (N_9858,N_6759,N_7587);
and U9859 (N_9859,N_4117,N_7598);
nand U9860 (N_9860,N_5093,N_7751);
nand U9861 (N_9861,N_5214,N_7505);
xnor U9862 (N_9862,N_6068,N_6961);
and U9863 (N_9863,N_5387,N_7568);
nand U9864 (N_9864,N_6907,N_7898);
or U9865 (N_9865,N_6191,N_4126);
nand U9866 (N_9866,N_6558,N_4637);
xor U9867 (N_9867,N_4173,N_4211);
xnor U9868 (N_9868,N_5762,N_7429);
or U9869 (N_9869,N_6562,N_5589);
xor U9870 (N_9870,N_5074,N_6599);
nor U9871 (N_9871,N_6248,N_4587);
nor U9872 (N_9872,N_5344,N_4105);
nand U9873 (N_9873,N_7585,N_6212);
nand U9874 (N_9874,N_6636,N_5151);
xor U9875 (N_9875,N_4944,N_4641);
and U9876 (N_9876,N_5744,N_5168);
nand U9877 (N_9877,N_7469,N_4530);
nor U9878 (N_9878,N_6697,N_5671);
and U9879 (N_9879,N_6046,N_4415);
nand U9880 (N_9880,N_5910,N_4152);
nand U9881 (N_9881,N_7862,N_5817);
nand U9882 (N_9882,N_7490,N_4287);
and U9883 (N_9883,N_4463,N_5284);
or U9884 (N_9884,N_5546,N_7217);
xnor U9885 (N_9885,N_6228,N_5432);
nand U9886 (N_9886,N_4668,N_5095);
nor U9887 (N_9887,N_5694,N_6076);
xnor U9888 (N_9888,N_4006,N_6360);
or U9889 (N_9889,N_5679,N_7134);
and U9890 (N_9890,N_4169,N_6864);
xor U9891 (N_9891,N_5517,N_5063);
xor U9892 (N_9892,N_4147,N_5490);
nor U9893 (N_9893,N_5323,N_4487);
nor U9894 (N_9894,N_4198,N_7060);
xnor U9895 (N_9895,N_6919,N_5669);
and U9896 (N_9896,N_6794,N_5321);
nor U9897 (N_9897,N_4236,N_4293);
and U9898 (N_9898,N_6047,N_5758);
or U9899 (N_9899,N_7042,N_5428);
xnor U9900 (N_9900,N_4524,N_7711);
nor U9901 (N_9901,N_4634,N_6545);
or U9902 (N_9902,N_6917,N_6379);
and U9903 (N_9903,N_6732,N_6303);
or U9904 (N_9904,N_6293,N_6256);
or U9905 (N_9905,N_6124,N_7525);
or U9906 (N_9906,N_5740,N_5536);
or U9907 (N_9907,N_5319,N_6926);
nand U9908 (N_9908,N_6616,N_7539);
or U9909 (N_9909,N_7048,N_4534);
and U9910 (N_9910,N_5029,N_4405);
nand U9911 (N_9911,N_7260,N_6093);
or U9912 (N_9912,N_4941,N_5630);
nand U9913 (N_9913,N_7753,N_5099);
nor U9914 (N_9914,N_7835,N_6331);
nor U9915 (N_9915,N_4816,N_7321);
and U9916 (N_9916,N_7176,N_5190);
nand U9917 (N_9917,N_5985,N_4995);
nand U9918 (N_9918,N_4103,N_6464);
nand U9919 (N_9919,N_4845,N_4002);
or U9920 (N_9920,N_4133,N_7881);
xor U9921 (N_9921,N_5503,N_7416);
or U9922 (N_9922,N_6717,N_7936);
nand U9923 (N_9923,N_6108,N_5913);
nor U9924 (N_9924,N_4127,N_7987);
nor U9925 (N_9925,N_6854,N_4980);
xnor U9926 (N_9926,N_6686,N_6399);
or U9927 (N_9927,N_6595,N_5439);
nand U9928 (N_9928,N_6344,N_4938);
nor U9929 (N_9929,N_5257,N_4795);
nand U9930 (N_9930,N_4604,N_6714);
xnor U9931 (N_9931,N_4410,N_4835);
nand U9932 (N_9932,N_4034,N_4753);
and U9933 (N_9933,N_6985,N_5793);
nor U9934 (N_9934,N_5847,N_5192);
or U9935 (N_9935,N_5584,N_4074);
nor U9936 (N_9936,N_5822,N_4697);
nor U9937 (N_9937,N_6052,N_4796);
nor U9938 (N_9938,N_6302,N_4892);
or U9939 (N_9939,N_6993,N_4750);
nor U9940 (N_9940,N_7356,N_4225);
or U9941 (N_9941,N_7485,N_6882);
xnor U9942 (N_9942,N_4729,N_6563);
and U9943 (N_9943,N_7854,N_7515);
and U9944 (N_9944,N_4469,N_4679);
and U9945 (N_9945,N_5999,N_4226);
or U9946 (N_9946,N_7655,N_5878);
or U9947 (N_9947,N_7747,N_5776);
and U9948 (N_9948,N_7765,N_7358);
nand U9949 (N_9949,N_6444,N_6809);
or U9950 (N_9950,N_6967,N_5369);
and U9951 (N_9951,N_7172,N_5746);
nand U9952 (N_9952,N_7095,N_5464);
or U9953 (N_9953,N_6589,N_4122);
or U9954 (N_9954,N_6122,N_5388);
and U9955 (N_9955,N_7412,N_4525);
xor U9956 (N_9956,N_7684,N_7097);
nand U9957 (N_9957,N_5898,N_5620);
and U9958 (N_9958,N_4790,N_6452);
and U9959 (N_9959,N_6966,N_5568);
and U9960 (N_9960,N_7029,N_6467);
or U9961 (N_9961,N_4075,N_6229);
and U9962 (N_9962,N_7559,N_4601);
and U9963 (N_9963,N_4260,N_6389);
or U9964 (N_9964,N_5800,N_6955);
or U9965 (N_9965,N_6529,N_6532);
nand U9966 (N_9966,N_5853,N_7030);
nor U9967 (N_9967,N_6659,N_6160);
xnor U9968 (N_9968,N_7234,N_6210);
and U9969 (N_9969,N_7531,N_7110);
nand U9970 (N_9970,N_6187,N_6426);
or U9971 (N_9971,N_4947,N_4311);
nor U9972 (N_9972,N_7750,N_5508);
nor U9973 (N_9973,N_4568,N_6865);
and U9974 (N_9974,N_4059,N_7922);
nand U9975 (N_9975,N_6561,N_5038);
nor U9976 (N_9976,N_7785,N_6396);
nand U9977 (N_9977,N_7694,N_6280);
nor U9978 (N_9978,N_4294,N_4959);
xnor U9979 (N_9979,N_5518,N_7053);
and U9980 (N_9980,N_4382,N_5275);
or U9981 (N_9981,N_5796,N_7033);
nor U9982 (N_9982,N_5435,N_7002);
or U9983 (N_9983,N_4047,N_6687);
nor U9984 (N_9984,N_6747,N_5273);
nor U9985 (N_9985,N_6556,N_7954);
or U9986 (N_9986,N_5689,N_4447);
or U9987 (N_9987,N_4095,N_6609);
or U9988 (N_9988,N_6026,N_6286);
nor U9989 (N_9989,N_5427,N_7457);
nor U9990 (N_9990,N_7494,N_6744);
or U9991 (N_9991,N_7831,N_7815);
nand U9992 (N_9992,N_6354,N_6998);
nand U9993 (N_9993,N_5579,N_4334);
nand U9994 (N_9994,N_5083,N_7855);
and U9995 (N_9995,N_5333,N_7487);
or U9996 (N_9996,N_5657,N_5492);
or U9997 (N_9997,N_4768,N_7787);
xor U9998 (N_9998,N_7117,N_5703);
nor U9999 (N_9999,N_6436,N_7025);
or U10000 (N_10000,N_5577,N_7653);
or U10001 (N_10001,N_6125,N_5533);
nand U10002 (N_10002,N_5354,N_6562);
and U10003 (N_10003,N_7427,N_6969);
nor U10004 (N_10004,N_6510,N_6732);
or U10005 (N_10005,N_5832,N_5547);
nand U10006 (N_10006,N_7072,N_7557);
or U10007 (N_10007,N_5235,N_5047);
and U10008 (N_10008,N_6633,N_6747);
and U10009 (N_10009,N_7786,N_4469);
and U10010 (N_10010,N_7296,N_5808);
or U10011 (N_10011,N_4440,N_4701);
nor U10012 (N_10012,N_7077,N_5651);
and U10013 (N_10013,N_6478,N_5021);
nor U10014 (N_10014,N_7076,N_6693);
xnor U10015 (N_10015,N_6456,N_4198);
nor U10016 (N_10016,N_5265,N_4175);
and U10017 (N_10017,N_6918,N_5678);
or U10018 (N_10018,N_4303,N_5725);
nand U10019 (N_10019,N_7944,N_5827);
nor U10020 (N_10020,N_5192,N_4521);
nand U10021 (N_10021,N_5202,N_5187);
or U10022 (N_10022,N_4373,N_4527);
nor U10023 (N_10023,N_4557,N_5524);
or U10024 (N_10024,N_6190,N_5736);
xnor U10025 (N_10025,N_7350,N_5953);
or U10026 (N_10026,N_7293,N_4134);
nand U10027 (N_10027,N_5778,N_6112);
or U10028 (N_10028,N_5402,N_4272);
or U10029 (N_10029,N_7606,N_5656);
and U10030 (N_10030,N_5806,N_6874);
and U10031 (N_10031,N_7845,N_6326);
or U10032 (N_10032,N_4449,N_5960);
nor U10033 (N_10033,N_7776,N_4383);
nand U10034 (N_10034,N_5896,N_5534);
nand U10035 (N_10035,N_4276,N_7266);
nor U10036 (N_10036,N_7068,N_7145);
nand U10037 (N_10037,N_6677,N_6631);
and U10038 (N_10038,N_5399,N_5319);
nand U10039 (N_10039,N_6845,N_4636);
nor U10040 (N_10040,N_4420,N_6796);
nor U10041 (N_10041,N_6443,N_6812);
nand U10042 (N_10042,N_5693,N_7388);
xnor U10043 (N_10043,N_7245,N_7361);
nand U10044 (N_10044,N_6242,N_7584);
and U10045 (N_10045,N_7739,N_6902);
nor U10046 (N_10046,N_5065,N_7563);
nand U10047 (N_10047,N_7844,N_4698);
or U10048 (N_10048,N_4421,N_5487);
and U10049 (N_10049,N_5607,N_7788);
and U10050 (N_10050,N_5677,N_7254);
nand U10051 (N_10051,N_4664,N_7779);
nand U10052 (N_10052,N_5028,N_7485);
and U10053 (N_10053,N_7945,N_6747);
and U10054 (N_10054,N_5713,N_5027);
or U10055 (N_10055,N_5427,N_7693);
nand U10056 (N_10056,N_4800,N_6282);
or U10057 (N_10057,N_5652,N_7680);
nand U10058 (N_10058,N_7276,N_6429);
nand U10059 (N_10059,N_5704,N_5672);
nand U10060 (N_10060,N_7072,N_5604);
nand U10061 (N_10061,N_5642,N_4920);
xnor U10062 (N_10062,N_4248,N_4859);
or U10063 (N_10063,N_5792,N_6696);
nor U10064 (N_10064,N_6452,N_6964);
nand U10065 (N_10065,N_5638,N_7030);
nor U10066 (N_10066,N_4619,N_7416);
and U10067 (N_10067,N_4246,N_4518);
xnor U10068 (N_10068,N_5966,N_7912);
or U10069 (N_10069,N_7551,N_7961);
or U10070 (N_10070,N_7779,N_7193);
xor U10071 (N_10071,N_7423,N_4493);
and U10072 (N_10072,N_4424,N_5100);
or U10073 (N_10073,N_6199,N_5950);
nor U10074 (N_10074,N_5196,N_6008);
and U10075 (N_10075,N_6167,N_6498);
or U10076 (N_10076,N_5028,N_7866);
nor U10077 (N_10077,N_4758,N_6659);
nand U10078 (N_10078,N_4125,N_4852);
or U10079 (N_10079,N_6830,N_6368);
nand U10080 (N_10080,N_5708,N_7820);
or U10081 (N_10081,N_6572,N_7624);
and U10082 (N_10082,N_4891,N_4527);
or U10083 (N_10083,N_5636,N_5562);
and U10084 (N_10084,N_5675,N_7102);
nor U10085 (N_10085,N_6206,N_7116);
xor U10086 (N_10086,N_6699,N_6737);
nor U10087 (N_10087,N_4323,N_6736);
or U10088 (N_10088,N_6178,N_6691);
xnor U10089 (N_10089,N_6911,N_4415);
or U10090 (N_10090,N_4082,N_5653);
nand U10091 (N_10091,N_6156,N_5639);
xnor U10092 (N_10092,N_6568,N_6132);
and U10093 (N_10093,N_7882,N_5979);
and U10094 (N_10094,N_5080,N_7295);
nand U10095 (N_10095,N_7883,N_6656);
nor U10096 (N_10096,N_6379,N_4746);
nand U10097 (N_10097,N_6841,N_4581);
nor U10098 (N_10098,N_4456,N_7799);
nor U10099 (N_10099,N_6631,N_5597);
nand U10100 (N_10100,N_7429,N_7055);
or U10101 (N_10101,N_4306,N_5031);
or U10102 (N_10102,N_6943,N_7312);
and U10103 (N_10103,N_7533,N_6575);
nand U10104 (N_10104,N_7799,N_5478);
nand U10105 (N_10105,N_6617,N_7377);
nand U10106 (N_10106,N_6323,N_4097);
nand U10107 (N_10107,N_6650,N_4269);
nand U10108 (N_10108,N_6895,N_4245);
nor U10109 (N_10109,N_7579,N_4101);
or U10110 (N_10110,N_5496,N_7403);
and U10111 (N_10111,N_5005,N_6956);
xor U10112 (N_10112,N_7887,N_4146);
or U10113 (N_10113,N_7851,N_5219);
nand U10114 (N_10114,N_4096,N_4462);
or U10115 (N_10115,N_6397,N_7441);
nand U10116 (N_10116,N_5634,N_5172);
nand U10117 (N_10117,N_5112,N_7483);
or U10118 (N_10118,N_7488,N_5412);
nand U10119 (N_10119,N_7170,N_7567);
xor U10120 (N_10120,N_6648,N_6878);
and U10121 (N_10121,N_7296,N_6484);
xor U10122 (N_10122,N_6980,N_4565);
nor U10123 (N_10123,N_4844,N_4460);
xnor U10124 (N_10124,N_5933,N_6560);
or U10125 (N_10125,N_7425,N_7867);
nand U10126 (N_10126,N_7715,N_4582);
and U10127 (N_10127,N_7755,N_6117);
nor U10128 (N_10128,N_7818,N_7047);
nor U10129 (N_10129,N_7326,N_5995);
nor U10130 (N_10130,N_6628,N_4867);
and U10131 (N_10131,N_4690,N_4723);
nor U10132 (N_10132,N_6802,N_7803);
or U10133 (N_10133,N_6550,N_5555);
and U10134 (N_10134,N_7128,N_6944);
or U10135 (N_10135,N_4635,N_7492);
nand U10136 (N_10136,N_5429,N_6263);
nor U10137 (N_10137,N_6206,N_5699);
or U10138 (N_10138,N_5832,N_4385);
xor U10139 (N_10139,N_7002,N_4351);
xnor U10140 (N_10140,N_6857,N_4281);
or U10141 (N_10141,N_5792,N_7546);
or U10142 (N_10142,N_7849,N_5979);
nor U10143 (N_10143,N_4102,N_7826);
nor U10144 (N_10144,N_5140,N_4621);
xnor U10145 (N_10145,N_6787,N_4027);
nor U10146 (N_10146,N_5621,N_7669);
xnor U10147 (N_10147,N_6194,N_4757);
and U10148 (N_10148,N_6693,N_4837);
nand U10149 (N_10149,N_5797,N_5415);
and U10150 (N_10150,N_5012,N_5288);
nor U10151 (N_10151,N_4663,N_4602);
xor U10152 (N_10152,N_4519,N_4112);
nand U10153 (N_10153,N_6359,N_5507);
and U10154 (N_10154,N_5911,N_4881);
nor U10155 (N_10155,N_7782,N_4105);
nor U10156 (N_10156,N_7146,N_6926);
nand U10157 (N_10157,N_7002,N_6915);
nand U10158 (N_10158,N_7177,N_4622);
nor U10159 (N_10159,N_5884,N_6400);
nor U10160 (N_10160,N_6137,N_6599);
nor U10161 (N_10161,N_7752,N_6416);
xnor U10162 (N_10162,N_7221,N_7520);
nand U10163 (N_10163,N_4515,N_7565);
or U10164 (N_10164,N_6283,N_6521);
or U10165 (N_10165,N_5677,N_6427);
and U10166 (N_10166,N_7906,N_7995);
or U10167 (N_10167,N_7698,N_5436);
and U10168 (N_10168,N_5177,N_7142);
nor U10169 (N_10169,N_7228,N_6696);
nand U10170 (N_10170,N_4623,N_4327);
and U10171 (N_10171,N_4347,N_7538);
nand U10172 (N_10172,N_4150,N_4410);
xor U10173 (N_10173,N_7739,N_7122);
nor U10174 (N_10174,N_6638,N_5452);
nand U10175 (N_10175,N_7625,N_4377);
or U10176 (N_10176,N_5212,N_5818);
xnor U10177 (N_10177,N_7022,N_5013);
nand U10178 (N_10178,N_5654,N_4008);
nor U10179 (N_10179,N_5030,N_5333);
or U10180 (N_10180,N_6752,N_6746);
or U10181 (N_10181,N_7657,N_4843);
nand U10182 (N_10182,N_4576,N_6885);
and U10183 (N_10183,N_7443,N_4615);
and U10184 (N_10184,N_7051,N_4065);
or U10185 (N_10185,N_7147,N_5273);
and U10186 (N_10186,N_7115,N_6461);
nand U10187 (N_10187,N_5477,N_6727);
xnor U10188 (N_10188,N_7336,N_4451);
nand U10189 (N_10189,N_5621,N_7576);
xnor U10190 (N_10190,N_5862,N_6103);
and U10191 (N_10191,N_4811,N_4509);
nor U10192 (N_10192,N_6589,N_5829);
nor U10193 (N_10193,N_4336,N_5210);
nor U10194 (N_10194,N_5372,N_4712);
and U10195 (N_10195,N_7345,N_5492);
nor U10196 (N_10196,N_5488,N_5300);
nand U10197 (N_10197,N_4434,N_6174);
nand U10198 (N_10198,N_5834,N_6401);
or U10199 (N_10199,N_7334,N_6924);
and U10200 (N_10200,N_7224,N_7508);
or U10201 (N_10201,N_6978,N_5085);
or U10202 (N_10202,N_5025,N_6578);
nand U10203 (N_10203,N_5967,N_4448);
and U10204 (N_10204,N_4390,N_7513);
and U10205 (N_10205,N_4685,N_7423);
nand U10206 (N_10206,N_5256,N_4780);
or U10207 (N_10207,N_5524,N_6613);
nor U10208 (N_10208,N_5972,N_6214);
and U10209 (N_10209,N_4449,N_7366);
nor U10210 (N_10210,N_7866,N_4717);
and U10211 (N_10211,N_4808,N_6646);
or U10212 (N_10212,N_5960,N_5414);
nand U10213 (N_10213,N_5720,N_5778);
or U10214 (N_10214,N_7568,N_6766);
or U10215 (N_10215,N_7673,N_5715);
and U10216 (N_10216,N_7642,N_6605);
and U10217 (N_10217,N_6111,N_7850);
or U10218 (N_10218,N_6811,N_5528);
nand U10219 (N_10219,N_7680,N_4648);
nor U10220 (N_10220,N_5733,N_4217);
nand U10221 (N_10221,N_4417,N_6568);
nand U10222 (N_10222,N_7552,N_7878);
nor U10223 (N_10223,N_7437,N_4397);
nor U10224 (N_10224,N_7858,N_6155);
and U10225 (N_10225,N_4989,N_5145);
or U10226 (N_10226,N_5751,N_6033);
nand U10227 (N_10227,N_4890,N_5027);
nor U10228 (N_10228,N_7795,N_4194);
nor U10229 (N_10229,N_5582,N_5495);
nor U10230 (N_10230,N_7843,N_6129);
or U10231 (N_10231,N_4992,N_5517);
or U10232 (N_10232,N_7870,N_5856);
nor U10233 (N_10233,N_5709,N_4114);
nand U10234 (N_10234,N_5031,N_6747);
xnor U10235 (N_10235,N_5798,N_6250);
nand U10236 (N_10236,N_7911,N_6900);
nor U10237 (N_10237,N_6639,N_5437);
or U10238 (N_10238,N_7770,N_6099);
nor U10239 (N_10239,N_6644,N_5576);
and U10240 (N_10240,N_4730,N_7260);
and U10241 (N_10241,N_4806,N_5627);
or U10242 (N_10242,N_6036,N_7776);
xor U10243 (N_10243,N_5558,N_7360);
and U10244 (N_10244,N_7821,N_7537);
or U10245 (N_10245,N_7641,N_7225);
and U10246 (N_10246,N_4755,N_7391);
xnor U10247 (N_10247,N_6558,N_4434);
nand U10248 (N_10248,N_6407,N_4565);
xnor U10249 (N_10249,N_6968,N_4062);
nand U10250 (N_10250,N_6232,N_5693);
and U10251 (N_10251,N_6547,N_5841);
xor U10252 (N_10252,N_6047,N_7043);
nor U10253 (N_10253,N_4532,N_6252);
nor U10254 (N_10254,N_6782,N_6254);
and U10255 (N_10255,N_6262,N_5711);
nand U10256 (N_10256,N_6381,N_6627);
xnor U10257 (N_10257,N_6180,N_5307);
and U10258 (N_10258,N_7250,N_7162);
or U10259 (N_10259,N_7555,N_4170);
nor U10260 (N_10260,N_6213,N_6608);
nor U10261 (N_10261,N_7374,N_7363);
nor U10262 (N_10262,N_7475,N_6472);
nor U10263 (N_10263,N_5030,N_6155);
or U10264 (N_10264,N_7010,N_6353);
nor U10265 (N_10265,N_6555,N_6471);
and U10266 (N_10266,N_6475,N_4180);
nor U10267 (N_10267,N_5901,N_6457);
nand U10268 (N_10268,N_7906,N_4986);
or U10269 (N_10269,N_7453,N_5193);
nand U10270 (N_10270,N_7951,N_7131);
nand U10271 (N_10271,N_5209,N_7933);
or U10272 (N_10272,N_5189,N_6358);
nand U10273 (N_10273,N_6770,N_7731);
or U10274 (N_10274,N_4490,N_7737);
xnor U10275 (N_10275,N_6112,N_5598);
or U10276 (N_10276,N_5110,N_4875);
xnor U10277 (N_10277,N_6681,N_6124);
nand U10278 (N_10278,N_7441,N_6857);
nand U10279 (N_10279,N_5438,N_6030);
nand U10280 (N_10280,N_5669,N_6336);
nor U10281 (N_10281,N_5522,N_7545);
and U10282 (N_10282,N_4347,N_6285);
xor U10283 (N_10283,N_5900,N_4633);
or U10284 (N_10284,N_5976,N_5007);
or U10285 (N_10285,N_7680,N_4840);
or U10286 (N_10286,N_4320,N_7879);
or U10287 (N_10287,N_4473,N_7729);
or U10288 (N_10288,N_4970,N_5999);
xor U10289 (N_10289,N_4825,N_6389);
nor U10290 (N_10290,N_4313,N_5909);
or U10291 (N_10291,N_5241,N_6131);
nand U10292 (N_10292,N_5965,N_7354);
nand U10293 (N_10293,N_5229,N_6995);
or U10294 (N_10294,N_7154,N_7062);
nand U10295 (N_10295,N_6523,N_7527);
or U10296 (N_10296,N_5498,N_7645);
nand U10297 (N_10297,N_5637,N_5522);
xnor U10298 (N_10298,N_6956,N_6573);
or U10299 (N_10299,N_5883,N_4988);
nor U10300 (N_10300,N_4193,N_6376);
and U10301 (N_10301,N_5503,N_5469);
and U10302 (N_10302,N_6413,N_6484);
nor U10303 (N_10303,N_5520,N_4227);
nor U10304 (N_10304,N_6359,N_6476);
and U10305 (N_10305,N_4534,N_6989);
and U10306 (N_10306,N_6976,N_4077);
or U10307 (N_10307,N_7595,N_6181);
xor U10308 (N_10308,N_4820,N_5841);
and U10309 (N_10309,N_6169,N_4740);
or U10310 (N_10310,N_5335,N_5079);
and U10311 (N_10311,N_7714,N_4350);
or U10312 (N_10312,N_7515,N_6468);
or U10313 (N_10313,N_7411,N_4189);
nor U10314 (N_10314,N_7794,N_6606);
nor U10315 (N_10315,N_7632,N_5370);
nor U10316 (N_10316,N_4717,N_7828);
or U10317 (N_10317,N_6122,N_7462);
nor U10318 (N_10318,N_6782,N_4000);
and U10319 (N_10319,N_7094,N_7555);
and U10320 (N_10320,N_6590,N_7113);
xnor U10321 (N_10321,N_6442,N_4756);
nor U10322 (N_10322,N_4274,N_4788);
nand U10323 (N_10323,N_4519,N_7401);
or U10324 (N_10324,N_6956,N_5798);
nand U10325 (N_10325,N_7957,N_6008);
and U10326 (N_10326,N_4915,N_6444);
nand U10327 (N_10327,N_6232,N_5899);
and U10328 (N_10328,N_6484,N_7597);
nand U10329 (N_10329,N_4383,N_6952);
nor U10330 (N_10330,N_5841,N_5244);
and U10331 (N_10331,N_4159,N_7034);
or U10332 (N_10332,N_6600,N_7698);
nand U10333 (N_10333,N_7791,N_7314);
and U10334 (N_10334,N_7718,N_6168);
nand U10335 (N_10335,N_7118,N_7503);
or U10336 (N_10336,N_5589,N_4623);
and U10337 (N_10337,N_7965,N_5372);
nor U10338 (N_10338,N_5745,N_6064);
nand U10339 (N_10339,N_7500,N_4851);
or U10340 (N_10340,N_7590,N_7221);
nand U10341 (N_10341,N_5314,N_6856);
and U10342 (N_10342,N_6719,N_5920);
or U10343 (N_10343,N_5237,N_7244);
nor U10344 (N_10344,N_4499,N_5229);
and U10345 (N_10345,N_6504,N_5716);
nor U10346 (N_10346,N_6889,N_7671);
and U10347 (N_10347,N_7105,N_6533);
and U10348 (N_10348,N_6470,N_7338);
nor U10349 (N_10349,N_6038,N_5999);
nand U10350 (N_10350,N_7193,N_5592);
or U10351 (N_10351,N_5304,N_5484);
and U10352 (N_10352,N_5094,N_5588);
nor U10353 (N_10353,N_5404,N_4495);
and U10354 (N_10354,N_4203,N_6468);
nor U10355 (N_10355,N_5259,N_6831);
and U10356 (N_10356,N_4088,N_5596);
and U10357 (N_10357,N_6294,N_4117);
nand U10358 (N_10358,N_7135,N_6354);
or U10359 (N_10359,N_5567,N_5488);
nand U10360 (N_10360,N_5583,N_6056);
nor U10361 (N_10361,N_7579,N_7009);
and U10362 (N_10362,N_5035,N_4462);
nand U10363 (N_10363,N_6291,N_5833);
nor U10364 (N_10364,N_4249,N_7601);
or U10365 (N_10365,N_6273,N_7114);
nand U10366 (N_10366,N_5482,N_6086);
nand U10367 (N_10367,N_6410,N_6714);
nand U10368 (N_10368,N_7289,N_6437);
nand U10369 (N_10369,N_6010,N_7190);
nand U10370 (N_10370,N_7872,N_5936);
and U10371 (N_10371,N_6960,N_6306);
or U10372 (N_10372,N_7603,N_6551);
and U10373 (N_10373,N_6519,N_6344);
or U10374 (N_10374,N_6406,N_5066);
or U10375 (N_10375,N_7841,N_6349);
nor U10376 (N_10376,N_7401,N_4531);
or U10377 (N_10377,N_5297,N_4082);
and U10378 (N_10378,N_4950,N_4550);
nor U10379 (N_10379,N_6428,N_4118);
nor U10380 (N_10380,N_7865,N_6700);
and U10381 (N_10381,N_7836,N_7845);
nor U10382 (N_10382,N_5459,N_6005);
nor U10383 (N_10383,N_4540,N_4160);
or U10384 (N_10384,N_4038,N_7875);
xor U10385 (N_10385,N_5421,N_6810);
nand U10386 (N_10386,N_5567,N_7408);
nor U10387 (N_10387,N_6951,N_4248);
and U10388 (N_10388,N_6543,N_4532);
nor U10389 (N_10389,N_7322,N_7950);
nand U10390 (N_10390,N_7330,N_4727);
nor U10391 (N_10391,N_6803,N_6041);
nand U10392 (N_10392,N_7011,N_4472);
nor U10393 (N_10393,N_6686,N_4263);
nor U10394 (N_10394,N_6618,N_6100);
and U10395 (N_10395,N_7693,N_5577);
nand U10396 (N_10396,N_6112,N_4402);
and U10397 (N_10397,N_6447,N_6975);
nand U10398 (N_10398,N_6047,N_7527);
or U10399 (N_10399,N_7213,N_7665);
and U10400 (N_10400,N_5143,N_7096);
nand U10401 (N_10401,N_4564,N_7711);
and U10402 (N_10402,N_4524,N_6668);
xnor U10403 (N_10403,N_7148,N_7237);
xor U10404 (N_10404,N_6584,N_5577);
and U10405 (N_10405,N_6798,N_7120);
and U10406 (N_10406,N_5283,N_6511);
and U10407 (N_10407,N_5517,N_5909);
or U10408 (N_10408,N_5487,N_4235);
or U10409 (N_10409,N_4647,N_4199);
and U10410 (N_10410,N_6521,N_6495);
nor U10411 (N_10411,N_5637,N_6616);
xnor U10412 (N_10412,N_4734,N_7174);
and U10413 (N_10413,N_7191,N_7484);
nand U10414 (N_10414,N_5163,N_7069);
and U10415 (N_10415,N_6999,N_4965);
and U10416 (N_10416,N_5645,N_7195);
and U10417 (N_10417,N_5388,N_6861);
nor U10418 (N_10418,N_4719,N_5962);
and U10419 (N_10419,N_6051,N_5827);
or U10420 (N_10420,N_5168,N_6692);
nor U10421 (N_10421,N_7507,N_7780);
nor U10422 (N_10422,N_6323,N_7521);
nor U10423 (N_10423,N_6157,N_6850);
nor U10424 (N_10424,N_4444,N_5690);
or U10425 (N_10425,N_4017,N_5883);
and U10426 (N_10426,N_6772,N_4345);
nand U10427 (N_10427,N_5621,N_7197);
nor U10428 (N_10428,N_6442,N_7332);
nand U10429 (N_10429,N_6465,N_4069);
nand U10430 (N_10430,N_6262,N_6081);
or U10431 (N_10431,N_4637,N_6545);
nor U10432 (N_10432,N_4503,N_5596);
nor U10433 (N_10433,N_5751,N_7886);
and U10434 (N_10434,N_5101,N_5972);
or U10435 (N_10435,N_4706,N_4097);
and U10436 (N_10436,N_5950,N_5649);
nand U10437 (N_10437,N_7177,N_5482);
nor U10438 (N_10438,N_7305,N_5053);
nand U10439 (N_10439,N_5183,N_6899);
or U10440 (N_10440,N_7116,N_7311);
or U10441 (N_10441,N_7331,N_6624);
and U10442 (N_10442,N_6112,N_5502);
nand U10443 (N_10443,N_7120,N_5214);
nor U10444 (N_10444,N_7598,N_4387);
and U10445 (N_10445,N_4138,N_7954);
and U10446 (N_10446,N_7990,N_6343);
xor U10447 (N_10447,N_6881,N_5373);
nand U10448 (N_10448,N_6282,N_7939);
nand U10449 (N_10449,N_4554,N_7769);
and U10450 (N_10450,N_4421,N_4140);
and U10451 (N_10451,N_5532,N_4385);
and U10452 (N_10452,N_5629,N_6279);
and U10453 (N_10453,N_4995,N_5503);
xor U10454 (N_10454,N_7824,N_5594);
nand U10455 (N_10455,N_4080,N_5464);
or U10456 (N_10456,N_5801,N_5363);
and U10457 (N_10457,N_5280,N_5709);
nor U10458 (N_10458,N_6642,N_5743);
nand U10459 (N_10459,N_6142,N_5922);
or U10460 (N_10460,N_5174,N_4846);
xor U10461 (N_10461,N_5880,N_4021);
nor U10462 (N_10462,N_7151,N_4695);
nor U10463 (N_10463,N_4973,N_4872);
or U10464 (N_10464,N_7382,N_4858);
nand U10465 (N_10465,N_6610,N_7634);
or U10466 (N_10466,N_6997,N_6745);
nand U10467 (N_10467,N_5721,N_5718);
nor U10468 (N_10468,N_5888,N_5330);
nor U10469 (N_10469,N_6783,N_5171);
nor U10470 (N_10470,N_5186,N_7807);
and U10471 (N_10471,N_5539,N_4751);
or U10472 (N_10472,N_5962,N_7828);
or U10473 (N_10473,N_6609,N_5645);
and U10474 (N_10474,N_5315,N_5936);
nand U10475 (N_10475,N_4386,N_6613);
nand U10476 (N_10476,N_6771,N_4103);
or U10477 (N_10477,N_5425,N_6430);
and U10478 (N_10478,N_4010,N_7434);
nor U10479 (N_10479,N_4181,N_4157);
xnor U10480 (N_10480,N_4406,N_7172);
and U10481 (N_10481,N_4333,N_7938);
nor U10482 (N_10482,N_5386,N_4828);
nor U10483 (N_10483,N_5425,N_7813);
and U10484 (N_10484,N_7892,N_4786);
and U10485 (N_10485,N_6942,N_7701);
nand U10486 (N_10486,N_5713,N_6410);
xnor U10487 (N_10487,N_7100,N_6267);
nand U10488 (N_10488,N_6457,N_4696);
and U10489 (N_10489,N_5107,N_4886);
nor U10490 (N_10490,N_5478,N_6088);
nor U10491 (N_10491,N_4371,N_7391);
nor U10492 (N_10492,N_5446,N_6373);
nand U10493 (N_10493,N_6525,N_7300);
and U10494 (N_10494,N_4719,N_7149);
nor U10495 (N_10495,N_5893,N_7166);
nor U10496 (N_10496,N_5011,N_4392);
and U10497 (N_10497,N_4362,N_5488);
xor U10498 (N_10498,N_4947,N_7068);
xnor U10499 (N_10499,N_4435,N_6661);
or U10500 (N_10500,N_7170,N_4675);
nand U10501 (N_10501,N_7491,N_7173);
nand U10502 (N_10502,N_5041,N_4915);
nand U10503 (N_10503,N_7714,N_4469);
xor U10504 (N_10504,N_5386,N_6847);
and U10505 (N_10505,N_4190,N_7205);
nand U10506 (N_10506,N_4557,N_7010);
and U10507 (N_10507,N_7350,N_6122);
or U10508 (N_10508,N_5699,N_4444);
and U10509 (N_10509,N_4601,N_6380);
nor U10510 (N_10510,N_4325,N_6369);
nor U10511 (N_10511,N_4438,N_5113);
xnor U10512 (N_10512,N_6065,N_7714);
or U10513 (N_10513,N_5804,N_7736);
nor U10514 (N_10514,N_4712,N_5155);
nor U10515 (N_10515,N_6723,N_6852);
nand U10516 (N_10516,N_7539,N_5152);
nand U10517 (N_10517,N_5200,N_4097);
nand U10518 (N_10518,N_6050,N_5917);
nor U10519 (N_10519,N_4479,N_4287);
or U10520 (N_10520,N_5507,N_5685);
xnor U10521 (N_10521,N_5443,N_4779);
or U10522 (N_10522,N_6144,N_4907);
and U10523 (N_10523,N_6171,N_4491);
nor U10524 (N_10524,N_4290,N_7725);
nand U10525 (N_10525,N_7327,N_5285);
and U10526 (N_10526,N_4793,N_5468);
and U10527 (N_10527,N_6541,N_7568);
or U10528 (N_10528,N_7333,N_5803);
and U10529 (N_10529,N_5895,N_5985);
nor U10530 (N_10530,N_5424,N_7978);
nand U10531 (N_10531,N_7507,N_7215);
xnor U10532 (N_10532,N_5411,N_4267);
nand U10533 (N_10533,N_5035,N_4224);
or U10534 (N_10534,N_4961,N_5124);
or U10535 (N_10535,N_7154,N_5856);
nor U10536 (N_10536,N_4220,N_6811);
or U10537 (N_10537,N_7909,N_6779);
nor U10538 (N_10538,N_4542,N_5395);
nand U10539 (N_10539,N_4095,N_6087);
and U10540 (N_10540,N_7679,N_7117);
or U10541 (N_10541,N_4515,N_7198);
nand U10542 (N_10542,N_4799,N_4318);
nand U10543 (N_10543,N_7109,N_4612);
nor U10544 (N_10544,N_6539,N_6204);
and U10545 (N_10545,N_6462,N_5819);
nand U10546 (N_10546,N_7807,N_6443);
or U10547 (N_10547,N_4508,N_7524);
nor U10548 (N_10548,N_4896,N_6391);
and U10549 (N_10549,N_6186,N_4430);
nand U10550 (N_10550,N_6336,N_6734);
or U10551 (N_10551,N_4523,N_6771);
nand U10552 (N_10552,N_7660,N_6067);
and U10553 (N_10553,N_5445,N_5222);
xor U10554 (N_10554,N_6305,N_7253);
xor U10555 (N_10555,N_7140,N_7695);
and U10556 (N_10556,N_4017,N_7873);
and U10557 (N_10557,N_6214,N_6394);
or U10558 (N_10558,N_4182,N_5771);
and U10559 (N_10559,N_7654,N_7207);
and U10560 (N_10560,N_5476,N_4666);
or U10561 (N_10561,N_4659,N_4914);
and U10562 (N_10562,N_4295,N_5201);
or U10563 (N_10563,N_7146,N_4621);
or U10564 (N_10564,N_5742,N_4432);
or U10565 (N_10565,N_4163,N_4646);
nor U10566 (N_10566,N_4111,N_7557);
nand U10567 (N_10567,N_7221,N_6271);
or U10568 (N_10568,N_7576,N_5832);
or U10569 (N_10569,N_7728,N_7636);
xor U10570 (N_10570,N_5145,N_4032);
nor U10571 (N_10571,N_4989,N_7660);
and U10572 (N_10572,N_7902,N_6191);
nand U10573 (N_10573,N_5872,N_7885);
xnor U10574 (N_10574,N_5758,N_6202);
nand U10575 (N_10575,N_6839,N_4198);
nand U10576 (N_10576,N_4344,N_5234);
and U10577 (N_10577,N_5790,N_7382);
nor U10578 (N_10578,N_4051,N_6020);
nand U10579 (N_10579,N_7992,N_6646);
xor U10580 (N_10580,N_6531,N_4461);
nand U10581 (N_10581,N_7777,N_5755);
xor U10582 (N_10582,N_7912,N_6653);
or U10583 (N_10583,N_4471,N_4341);
nand U10584 (N_10584,N_4089,N_4762);
and U10585 (N_10585,N_4882,N_6892);
nor U10586 (N_10586,N_7321,N_7682);
or U10587 (N_10587,N_4565,N_6816);
and U10588 (N_10588,N_7191,N_6357);
nor U10589 (N_10589,N_6506,N_5806);
nand U10590 (N_10590,N_6402,N_7591);
or U10591 (N_10591,N_7026,N_6355);
xnor U10592 (N_10592,N_4246,N_6987);
nand U10593 (N_10593,N_5265,N_7452);
and U10594 (N_10594,N_6257,N_4177);
or U10595 (N_10595,N_7413,N_5733);
nand U10596 (N_10596,N_7033,N_4240);
or U10597 (N_10597,N_7162,N_5179);
or U10598 (N_10598,N_7702,N_6109);
xor U10599 (N_10599,N_5299,N_4035);
nand U10600 (N_10600,N_5724,N_5815);
nand U10601 (N_10601,N_4420,N_4439);
or U10602 (N_10602,N_4870,N_4411);
or U10603 (N_10603,N_6879,N_6794);
and U10604 (N_10604,N_6367,N_5359);
or U10605 (N_10605,N_7674,N_5331);
nor U10606 (N_10606,N_7868,N_7269);
nor U10607 (N_10607,N_7580,N_4323);
and U10608 (N_10608,N_4705,N_4189);
nand U10609 (N_10609,N_6687,N_5651);
xor U10610 (N_10610,N_7049,N_4508);
and U10611 (N_10611,N_6237,N_7066);
or U10612 (N_10612,N_7306,N_4777);
nor U10613 (N_10613,N_7981,N_5874);
and U10614 (N_10614,N_6594,N_5967);
nor U10615 (N_10615,N_5379,N_5460);
nor U10616 (N_10616,N_7218,N_5610);
nor U10617 (N_10617,N_4346,N_6372);
nor U10618 (N_10618,N_4381,N_6854);
or U10619 (N_10619,N_5166,N_5874);
nor U10620 (N_10620,N_4102,N_6166);
nor U10621 (N_10621,N_4964,N_7386);
nand U10622 (N_10622,N_5660,N_6359);
nor U10623 (N_10623,N_6584,N_7138);
nor U10624 (N_10624,N_7414,N_7315);
nor U10625 (N_10625,N_7272,N_4470);
nor U10626 (N_10626,N_5697,N_5286);
nand U10627 (N_10627,N_6863,N_7775);
nor U10628 (N_10628,N_6304,N_7933);
nand U10629 (N_10629,N_5118,N_6492);
nand U10630 (N_10630,N_7053,N_7840);
xor U10631 (N_10631,N_7453,N_5933);
nand U10632 (N_10632,N_4760,N_4987);
nand U10633 (N_10633,N_5445,N_4184);
or U10634 (N_10634,N_5020,N_5720);
xnor U10635 (N_10635,N_4783,N_5207);
nand U10636 (N_10636,N_5097,N_5135);
and U10637 (N_10637,N_7469,N_7574);
nand U10638 (N_10638,N_7594,N_7652);
nor U10639 (N_10639,N_4505,N_4797);
xor U10640 (N_10640,N_4926,N_4340);
or U10641 (N_10641,N_6602,N_5586);
xnor U10642 (N_10642,N_5718,N_7202);
or U10643 (N_10643,N_6390,N_5956);
or U10644 (N_10644,N_5489,N_7330);
and U10645 (N_10645,N_6585,N_5097);
nor U10646 (N_10646,N_5320,N_7213);
or U10647 (N_10647,N_4660,N_7099);
and U10648 (N_10648,N_5575,N_7774);
and U10649 (N_10649,N_7652,N_7753);
or U10650 (N_10650,N_5889,N_5062);
nand U10651 (N_10651,N_5871,N_5435);
nor U10652 (N_10652,N_4384,N_4500);
xor U10653 (N_10653,N_4223,N_6422);
nor U10654 (N_10654,N_5110,N_5361);
nand U10655 (N_10655,N_6704,N_4279);
or U10656 (N_10656,N_7943,N_4450);
nor U10657 (N_10657,N_6278,N_7920);
or U10658 (N_10658,N_7407,N_6435);
and U10659 (N_10659,N_6590,N_6827);
nand U10660 (N_10660,N_4961,N_7942);
or U10661 (N_10661,N_6063,N_6346);
and U10662 (N_10662,N_6961,N_7711);
nand U10663 (N_10663,N_4687,N_7189);
and U10664 (N_10664,N_7572,N_6245);
nand U10665 (N_10665,N_4496,N_7389);
nor U10666 (N_10666,N_7278,N_4909);
nor U10667 (N_10667,N_4120,N_5450);
and U10668 (N_10668,N_5510,N_7385);
xor U10669 (N_10669,N_7237,N_5105);
or U10670 (N_10670,N_5913,N_7058);
or U10671 (N_10671,N_6562,N_7297);
nand U10672 (N_10672,N_6154,N_7838);
and U10673 (N_10673,N_6238,N_5832);
or U10674 (N_10674,N_5053,N_6791);
nor U10675 (N_10675,N_5338,N_4960);
nor U10676 (N_10676,N_5090,N_4492);
and U10677 (N_10677,N_4130,N_7851);
nor U10678 (N_10678,N_7888,N_6501);
and U10679 (N_10679,N_5327,N_6105);
or U10680 (N_10680,N_4058,N_4002);
and U10681 (N_10681,N_4859,N_6582);
nor U10682 (N_10682,N_7289,N_5234);
and U10683 (N_10683,N_6719,N_5334);
nor U10684 (N_10684,N_4183,N_5098);
xor U10685 (N_10685,N_4780,N_5693);
nand U10686 (N_10686,N_7779,N_5019);
nor U10687 (N_10687,N_4936,N_7405);
nand U10688 (N_10688,N_5920,N_6090);
or U10689 (N_10689,N_4813,N_7388);
nor U10690 (N_10690,N_4748,N_6016);
and U10691 (N_10691,N_4632,N_4388);
nand U10692 (N_10692,N_4776,N_5572);
xnor U10693 (N_10693,N_5795,N_5687);
nor U10694 (N_10694,N_7307,N_7943);
or U10695 (N_10695,N_7859,N_5327);
or U10696 (N_10696,N_7081,N_6449);
or U10697 (N_10697,N_6921,N_5825);
nor U10698 (N_10698,N_4816,N_7893);
nor U10699 (N_10699,N_7411,N_6107);
nand U10700 (N_10700,N_7316,N_5637);
or U10701 (N_10701,N_5976,N_4606);
and U10702 (N_10702,N_4361,N_7173);
nand U10703 (N_10703,N_4236,N_4941);
xor U10704 (N_10704,N_7934,N_4144);
nor U10705 (N_10705,N_7980,N_6205);
or U10706 (N_10706,N_7830,N_4931);
or U10707 (N_10707,N_7368,N_4771);
nand U10708 (N_10708,N_5500,N_4056);
and U10709 (N_10709,N_7982,N_7274);
nand U10710 (N_10710,N_6270,N_7495);
or U10711 (N_10711,N_6113,N_4824);
nor U10712 (N_10712,N_7795,N_5356);
and U10713 (N_10713,N_5180,N_5072);
and U10714 (N_10714,N_6902,N_6323);
nor U10715 (N_10715,N_6700,N_6105);
nor U10716 (N_10716,N_5823,N_5915);
nor U10717 (N_10717,N_7335,N_5281);
or U10718 (N_10718,N_5324,N_4682);
nor U10719 (N_10719,N_7934,N_4470);
nor U10720 (N_10720,N_5917,N_7839);
and U10721 (N_10721,N_4643,N_5307);
and U10722 (N_10722,N_5636,N_4567);
xor U10723 (N_10723,N_6302,N_4392);
nor U10724 (N_10724,N_4942,N_5880);
or U10725 (N_10725,N_5294,N_6043);
nand U10726 (N_10726,N_6593,N_4873);
or U10727 (N_10727,N_5050,N_4465);
or U10728 (N_10728,N_4622,N_5577);
nor U10729 (N_10729,N_6266,N_5737);
nand U10730 (N_10730,N_5204,N_7051);
nand U10731 (N_10731,N_5360,N_7802);
nand U10732 (N_10732,N_5780,N_4232);
nor U10733 (N_10733,N_7758,N_4270);
nor U10734 (N_10734,N_7607,N_5517);
nor U10735 (N_10735,N_4768,N_5763);
xor U10736 (N_10736,N_4609,N_5602);
or U10737 (N_10737,N_4227,N_4592);
and U10738 (N_10738,N_5826,N_4182);
or U10739 (N_10739,N_4139,N_6296);
and U10740 (N_10740,N_7005,N_7589);
and U10741 (N_10741,N_4251,N_5575);
nand U10742 (N_10742,N_6768,N_7733);
and U10743 (N_10743,N_6506,N_5804);
nor U10744 (N_10744,N_6441,N_4714);
and U10745 (N_10745,N_5562,N_6785);
xor U10746 (N_10746,N_6353,N_5913);
nor U10747 (N_10747,N_4996,N_5941);
nor U10748 (N_10748,N_7468,N_4909);
nor U10749 (N_10749,N_4486,N_7983);
and U10750 (N_10750,N_7942,N_5076);
or U10751 (N_10751,N_5533,N_4725);
nand U10752 (N_10752,N_5961,N_5930);
nor U10753 (N_10753,N_6414,N_4370);
or U10754 (N_10754,N_5695,N_5751);
nand U10755 (N_10755,N_4210,N_5606);
or U10756 (N_10756,N_7769,N_7549);
nor U10757 (N_10757,N_6581,N_6217);
nand U10758 (N_10758,N_6700,N_6607);
and U10759 (N_10759,N_6505,N_4410);
and U10760 (N_10760,N_7286,N_7726);
and U10761 (N_10761,N_6251,N_6148);
or U10762 (N_10762,N_5309,N_6614);
and U10763 (N_10763,N_5257,N_6384);
or U10764 (N_10764,N_5255,N_6179);
and U10765 (N_10765,N_7852,N_6559);
or U10766 (N_10766,N_6628,N_7600);
or U10767 (N_10767,N_7697,N_6671);
or U10768 (N_10768,N_6432,N_4546);
nand U10769 (N_10769,N_5759,N_5231);
nor U10770 (N_10770,N_5148,N_5582);
nand U10771 (N_10771,N_5543,N_6979);
nor U10772 (N_10772,N_6924,N_5746);
nor U10773 (N_10773,N_6890,N_6500);
xnor U10774 (N_10774,N_7395,N_4805);
nor U10775 (N_10775,N_5562,N_4518);
nor U10776 (N_10776,N_7785,N_5291);
nor U10777 (N_10777,N_7805,N_6544);
and U10778 (N_10778,N_4362,N_4857);
or U10779 (N_10779,N_7058,N_5063);
nor U10780 (N_10780,N_6110,N_4628);
or U10781 (N_10781,N_6249,N_5492);
and U10782 (N_10782,N_6688,N_6126);
nand U10783 (N_10783,N_7760,N_7439);
nor U10784 (N_10784,N_6903,N_4356);
xor U10785 (N_10785,N_6526,N_6118);
nor U10786 (N_10786,N_6258,N_7980);
nor U10787 (N_10787,N_5904,N_6727);
or U10788 (N_10788,N_7879,N_4312);
and U10789 (N_10789,N_7648,N_6432);
nand U10790 (N_10790,N_6052,N_7710);
or U10791 (N_10791,N_5455,N_6105);
nand U10792 (N_10792,N_5540,N_4680);
and U10793 (N_10793,N_7352,N_5410);
nor U10794 (N_10794,N_5246,N_7396);
nand U10795 (N_10795,N_6343,N_6820);
nand U10796 (N_10796,N_7018,N_4492);
and U10797 (N_10797,N_6869,N_7357);
and U10798 (N_10798,N_7173,N_5723);
xnor U10799 (N_10799,N_5916,N_7347);
nor U10800 (N_10800,N_4918,N_7843);
nand U10801 (N_10801,N_6910,N_6374);
and U10802 (N_10802,N_7997,N_5607);
nand U10803 (N_10803,N_6604,N_4933);
nand U10804 (N_10804,N_6618,N_4091);
or U10805 (N_10805,N_6029,N_4540);
nor U10806 (N_10806,N_4076,N_6678);
nand U10807 (N_10807,N_4166,N_5878);
nand U10808 (N_10808,N_5922,N_4846);
nand U10809 (N_10809,N_5253,N_7123);
nand U10810 (N_10810,N_4469,N_7481);
nor U10811 (N_10811,N_5749,N_7238);
or U10812 (N_10812,N_6677,N_7155);
nand U10813 (N_10813,N_6881,N_4630);
or U10814 (N_10814,N_7678,N_4613);
nand U10815 (N_10815,N_5969,N_5483);
and U10816 (N_10816,N_5766,N_5251);
nor U10817 (N_10817,N_5109,N_6064);
and U10818 (N_10818,N_5821,N_5830);
or U10819 (N_10819,N_7167,N_4268);
or U10820 (N_10820,N_4800,N_7554);
nor U10821 (N_10821,N_5728,N_6130);
or U10822 (N_10822,N_7401,N_7645);
nand U10823 (N_10823,N_4361,N_6480);
and U10824 (N_10824,N_4581,N_7605);
or U10825 (N_10825,N_7523,N_7924);
and U10826 (N_10826,N_4067,N_6952);
nand U10827 (N_10827,N_5055,N_7319);
and U10828 (N_10828,N_7267,N_5819);
nand U10829 (N_10829,N_4526,N_5775);
and U10830 (N_10830,N_6788,N_6092);
nor U10831 (N_10831,N_7292,N_4852);
xnor U10832 (N_10832,N_4815,N_6254);
or U10833 (N_10833,N_7408,N_5283);
nand U10834 (N_10834,N_4927,N_7966);
nor U10835 (N_10835,N_6865,N_6224);
and U10836 (N_10836,N_5641,N_6466);
nand U10837 (N_10837,N_6700,N_6377);
xor U10838 (N_10838,N_6008,N_6839);
nand U10839 (N_10839,N_4341,N_7823);
or U10840 (N_10840,N_6558,N_6643);
nor U10841 (N_10841,N_4287,N_4585);
and U10842 (N_10842,N_6024,N_7527);
nor U10843 (N_10843,N_7492,N_5502);
and U10844 (N_10844,N_4497,N_4699);
xor U10845 (N_10845,N_4471,N_5113);
and U10846 (N_10846,N_5925,N_5354);
nand U10847 (N_10847,N_4541,N_5446);
and U10848 (N_10848,N_6926,N_4063);
and U10849 (N_10849,N_6456,N_7157);
nand U10850 (N_10850,N_5403,N_6149);
and U10851 (N_10851,N_5799,N_7050);
nor U10852 (N_10852,N_5235,N_7664);
xnor U10853 (N_10853,N_7313,N_5894);
nor U10854 (N_10854,N_5344,N_4908);
nor U10855 (N_10855,N_4893,N_4201);
xor U10856 (N_10856,N_7124,N_6308);
nand U10857 (N_10857,N_4981,N_6911);
and U10858 (N_10858,N_6717,N_4535);
and U10859 (N_10859,N_4875,N_4252);
nor U10860 (N_10860,N_4840,N_6005);
nor U10861 (N_10861,N_4552,N_4362);
or U10862 (N_10862,N_5335,N_4220);
nor U10863 (N_10863,N_4039,N_4497);
nor U10864 (N_10864,N_4109,N_6694);
or U10865 (N_10865,N_6359,N_5501);
nand U10866 (N_10866,N_5945,N_7661);
xnor U10867 (N_10867,N_6599,N_7882);
xor U10868 (N_10868,N_5292,N_7948);
and U10869 (N_10869,N_4620,N_7588);
nor U10870 (N_10870,N_4303,N_5053);
nor U10871 (N_10871,N_7940,N_7795);
and U10872 (N_10872,N_5779,N_4072);
or U10873 (N_10873,N_6116,N_7197);
nand U10874 (N_10874,N_6340,N_5285);
nor U10875 (N_10875,N_4117,N_6622);
and U10876 (N_10876,N_4007,N_7057);
and U10877 (N_10877,N_5416,N_4513);
nor U10878 (N_10878,N_7127,N_7581);
nor U10879 (N_10879,N_5916,N_7465);
nor U10880 (N_10880,N_7662,N_6967);
xor U10881 (N_10881,N_7513,N_6763);
nor U10882 (N_10882,N_5458,N_4512);
or U10883 (N_10883,N_5805,N_6751);
or U10884 (N_10884,N_4948,N_4385);
nand U10885 (N_10885,N_5764,N_6582);
or U10886 (N_10886,N_6811,N_6271);
and U10887 (N_10887,N_6551,N_4466);
or U10888 (N_10888,N_7031,N_4081);
nor U10889 (N_10889,N_7722,N_4579);
or U10890 (N_10890,N_4822,N_6328);
nand U10891 (N_10891,N_4907,N_5506);
nand U10892 (N_10892,N_4848,N_4373);
and U10893 (N_10893,N_5836,N_7924);
and U10894 (N_10894,N_6260,N_4378);
nor U10895 (N_10895,N_6298,N_5084);
or U10896 (N_10896,N_5709,N_7059);
xor U10897 (N_10897,N_7216,N_5053);
or U10898 (N_10898,N_7257,N_5062);
or U10899 (N_10899,N_6968,N_7752);
and U10900 (N_10900,N_5345,N_6547);
xor U10901 (N_10901,N_7413,N_6308);
nand U10902 (N_10902,N_4627,N_7617);
or U10903 (N_10903,N_4805,N_6538);
or U10904 (N_10904,N_5802,N_7599);
and U10905 (N_10905,N_5478,N_4323);
xor U10906 (N_10906,N_7122,N_4104);
and U10907 (N_10907,N_7662,N_4862);
nor U10908 (N_10908,N_5297,N_4961);
nand U10909 (N_10909,N_5273,N_6780);
xor U10910 (N_10910,N_7601,N_5314);
and U10911 (N_10911,N_6935,N_4203);
or U10912 (N_10912,N_5481,N_6248);
or U10913 (N_10913,N_7205,N_5615);
nor U10914 (N_10914,N_6108,N_5446);
or U10915 (N_10915,N_5593,N_7084);
and U10916 (N_10916,N_7938,N_6275);
and U10917 (N_10917,N_6137,N_4663);
or U10918 (N_10918,N_6560,N_5343);
and U10919 (N_10919,N_7227,N_4048);
nor U10920 (N_10920,N_6458,N_4637);
xnor U10921 (N_10921,N_7339,N_5794);
nor U10922 (N_10922,N_5121,N_5418);
nand U10923 (N_10923,N_6836,N_7327);
nand U10924 (N_10924,N_6081,N_6659);
nand U10925 (N_10925,N_5293,N_5986);
nand U10926 (N_10926,N_6540,N_6413);
nor U10927 (N_10927,N_7245,N_7032);
or U10928 (N_10928,N_5621,N_7948);
nand U10929 (N_10929,N_5609,N_5098);
or U10930 (N_10930,N_5399,N_5121);
nor U10931 (N_10931,N_5603,N_4887);
or U10932 (N_10932,N_7270,N_5589);
nor U10933 (N_10933,N_5757,N_7779);
xor U10934 (N_10934,N_6689,N_7578);
xnor U10935 (N_10935,N_5265,N_6952);
nor U10936 (N_10936,N_5992,N_6175);
xnor U10937 (N_10937,N_6008,N_6718);
or U10938 (N_10938,N_7897,N_7444);
nor U10939 (N_10939,N_4031,N_7772);
and U10940 (N_10940,N_6183,N_5943);
xor U10941 (N_10941,N_6884,N_4892);
nor U10942 (N_10942,N_5602,N_6836);
nor U10943 (N_10943,N_4037,N_4130);
nand U10944 (N_10944,N_5865,N_6846);
or U10945 (N_10945,N_6143,N_5501);
nand U10946 (N_10946,N_6857,N_5354);
or U10947 (N_10947,N_7039,N_7508);
and U10948 (N_10948,N_7607,N_4617);
nand U10949 (N_10949,N_7414,N_4829);
and U10950 (N_10950,N_5716,N_7112);
and U10951 (N_10951,N_5881,N_5221);
or U10952 (N_10952,N_7175,N_5743);
nor U10953 (N_10953,N_7294,N_5714);
nand U10954 (N_10954,N_7048,N_4382);
and U10955 (N_10955,N_5278,N_5980);
nand U10956 (N_10956,N_6649,N_5210);
nor U10957 (N_10957,N_7772,N_4502);
nor U10958 (N_10958,N_7767,N_7105);
or U10959 (N_10959,N_7618,N_5847);
nand U10960 (N_10960,N_4124,N_6883);
or U10961 (N_10961,N_6829,N_7568);
nor U10962 (N_10962,N_5284,N_7209);
nor U10963 (N_10963,N_4462,N_7621);
xor U10964 (N_10964,N_4537,N_7059);
and U10965 (N_10965,N_7148,N_6158);
or U10966 (N_10966,N_6485,N_4878);
and U10967 (N_10967,N_5082,N_4673);
or U10968 (N_10968,N_5286,N_7314);
xnor U10969 (N_10969,N_6003,N_4476);
and U10970 (N_10970,N_7675,N_5883);
and U10971 (N_10971,N_6355,N_5310);
xnor U10972 (N_10972,N_5891,N_6161);
xnor U10973 (N_10973,N_7565,N_4185);
nor U10974 (N_10974,N_4270,N_6681);
nand U10975 (N_10975,N_4284,N_5285);
nor U10976 (N_10976,N_5907,N_4051);
nand U10977 (N_10977,N_7438,N_4691);
and U10978 (N_10978,N_4903,N_7202);
xor U10979 (N_10979,N_5114,N_5108);
or U10980 (N_10980,N_4808,N_7396);
nand U10981 (N_10981,N_5643,N_4500);
nand U10982 (N_10982,N_7350,N_5615);
and U10983 (N_10983,N_6022,N_7788);
or U10984 (N_10984,N_5355,N_6414);
or U10985 (N_10985,N_4290,N_4577);
or U10986 (N_10986,N_7487,N_5453);
nand U10987 (N_10987,N_7754,N_4338);
nand U10988 (N_10988,N_5258,N_4725);
nand U10989 (N_10989,N_4222,N_4169);
and U10990 (N_10990,N_5472,N_4862);
nor U10991 (N_10991,N_6511,N_6100);
xnor U10992 (N_10992,N_5339,N_6665);
nand U10993 (N_10993,N_4495,N_7957);
nand U10994 (N_10994,N_7452,N_6278);
or U10995 (N_10995,N_6921,N_4098);
nor U10996 (N_10996,N_5235,N_5951);
nand U10997 (N_10997,N_5567,N_5036);
and U10998 (N_10998,N_5217,N_6940);
nor U10999 (N_10999,N_4587,N_5361);
nor U11000 (N_11000,N_5498,N_6009);
nor U11001 (N_11001,N_5569,N_4064);
nand U11002 (N_11002,N_4671,N_5794);
nand U11003 (N_11003,N_4275,N_5563);
nor U11004 (N_11004,N_7666,N_5615);
nor U11005 (N_11005,N_7288,N_7815);
or U11006 (N_11006,N_5977,N_4309);
or U11007 (N_11007,N_5978,N_6727);
nand U11008 (N_11008,N_5971,N_6939);
and U11009 (N_11009,N_4653,N_6068);
nand U11010 (N_11010,N_7747,N_4436);
nand U11011 (N_11011,N_5688,N_5831);
or U11012 (N_11012,N_7944,N_6147);
nand U11013 (N_11013,N_4877,N_5777);
nor U11014 (N_11014,N_7983,N_7291);
xor U11015 (N_11015,N_4656,N_7214);
nor U11016 (N_11016,N_5413,N_7441);
or U11017 (N_11017,N_6390,N_6252);
and U11018 (N_11018,N_7149,N_4289);
nand U11019 (N_11019,N_7411,N_5728);
nand U11020 (N_11020,N_7545,N_7992);
nand U11021 (N_11021,N_7498,N_7231);
or U11022 (N_11022,N_6802,N_7927);
nand U11023 (N_11023,N_5466,N_7586);
and U11024 (N_11024,N_7677,N_5730);
or U11025 (N_11025,N_4847,N_5753);
nand U11026 (N_11026,N_5929,N_5964);
or U11027 (N_11027,N_7041,N_7289);
nor U11028 (N_11028,N_6168,N_6539);
xnor U11029 (N_11029,N_7156,N_5703);
nor U11030 (N_11030,N_5948,N_5277);
and U11031 (N_11031,N_6606,N_5726);
nor U11032 (N_11032,N_4514,N_6763);
or U11033 (N_11033,N_5440,N_6201);
nor U11034 (N_11034,N_7660,N_4678);
nand U11035 (N_11035,N_7255,N_5474);
nor U11036 (N_11036,N_4041,N_4651);
nor U11037 (N_11037,N_5580,N_6197);
nor U11038 (N_11038,N_4791,N_7718);
nor U11039 (N_11039,N_7805,N_7789);
nor U11040 (N_11040,N_6333,N_7365);
nand U11041 (N_11041,N_4777,N_6000);
nor U11042 (N_11042,N_5313,N_7258);
or U11043 (N_11043,N_7296,N_6938);
or U11044 (N_11044,N_5243,N_7181);
nand U11045 (N_11045,N_7421,N_4864);
nand U11046 (N_11046,N_7506,N_7741);
nand U11047 (N_11047,N_7405,N_7246);
nor U11048 (N_11048,N_7740,N_6062);
nor U11049 (N_11049,N_5040,N_7754);
nand U11050 (N_11050,N_6278,N_4499);
nor U11051 (N_11051,N_4642,N_6529);
or U11052 (N_11052,N_6775,N_5517);
nand U11053 (N_11053,N_7560,N_4227);
or U11054 (N_11054,N_6455,N_4746);
xnor U11055 (N_11055,N_5473,N_6119);
or U11056 (N_11056,N_5359,N_7713);
and U11057 (N_11057,N_4465,N_4488);
nand U11058 (N_11058,N_4891,N_5327);
nand U11059 (N_11059,N_5109,N_6528);
xnor U11060 (N_11060,N_5275,N_6129);
and U11061 (N_11061,N_5259,N_5985);
or U11062 (N_11062,N_4832,N_4528);
or U11063 (N_11063,N_6976,N_7703);
nand U11064 (N_11064,N_7952,N_6348);
nor U11065 (N_11065,N_7083,N_7078);
nor U11066 (N_11066,N_5579,N_7440);
nor U11067 (N_11067,N_6949,N_6464);
nor U11068 (N_11068,N_4538,N_4147);
nand U11069 (N_11069,N_7299,N_4742);
nand U11070 (N_11070,N_7961,N_7695);
or U11071 (N_11071,N_7891,N_4287);
nand U11072 (N_11072,N_4205,N_7217);
and U11073 (N_11073,N_6773,N_5191);
and U11074 (N_11074,N_7371,N_4379);
and U11075 (N_11075,N_7673,N_7912);
xnor U11076 (N_11076,N_6744,N_7292);
xor U11077 (N_11077,N_5014,N_6706);
or U11078 (N_11078,N_5079,N_7099);
or U11079 (N_11079,N_7043,N_7764);
or U11080 (N_11080,N_7648,N_6288);
nor U11081 (N_11081,N_7179,N_7916);
nor U11082 (N_11082,N_6947,N_5243);
or U11083 (N_11083,N_4978,N_6260);
or U11084 (N_11084,N_6129,N_6357);
and U11085 (N_11085,N_4638,N_5751);
or U11086 (N_11086,N_6537,N_5620);
or U11087 (N_11087,N_5008,N_4061);
nor U11088 (N_11088,N_5300,N_6873);
and U11089 (N_11089,N_6611,N_5865);
nand U11090 (N_11090,N_6986,N_6214);
and U11091 (N_11091,N_4345,N_6761);
and U11092 (N_11092,N_7475,N_5926);
nor U11093 (N_11093,N_6143,N_6239);
or U11094 (N_11094,N_7657,N_5694);
or U11095 (N_11095,N_6440,N_5050);
and U11096 (N_11096,N_6504,N_7479);
nor U11097 (N_11097,N_7221,N_6238);
nand U11098 (N_11098,N_6670,N_7468);
nand U11099 (N_11099,N_6991,N_5669);
and U11100 (N_11100,N_6556,N_6202);
nand U11101 (N_11101,N_6239,N_5501);
xnor U11102 (N_11102,N_7594,N_5204);
and U11103 (N_11103,N_4046,N_6377);
or U11104 (N_11104,N_4197,N_5663);
xnor U11105 (N_11105,N_6849,N_4730);
nand U11106 (N_11106,N_5229,N_6531);
nand U11107 (N_11107,N_5245,N_7588);
and U11108 (N_11108,N_6747,N_5013);
and U11109 (N_11109,N_7679,N_6795);
nand U11110 (N_11110,N_4487,N_4056);
or U11111 (N_11111,N_5866,N_4359);
and U11112 (N_11112,N_6812,N_6656);
nor U11113 (N_11113,N_6584,N_5437);
or U11114 (N_11114,N_6373,N_6277);
nand U11115 (N_11115,N_7233,N_7129);
and U11116 (N_11116,N_7924,N_5011);
or U11117 (N_11117,N_4981,N_5823);
nand U11118 (N_11118,N_4470,N_5255);
nor U11119 (N_11119,N_6725,N_5212);
or U11120 (N_11120,N_4686,N_4994);
or U11121 (N_11121,N_6129,N_7828);
nor U11122 (N_11122,N_4167,N_4236);
or U11123 (N_11123,N_4905,N_5341);
or U11124 (N_11124,N_7187,N_7992);
xnor U11125 (N_11125,N_4910,N_4334);
nor U11126 (N_11126,N_7254,N_7826);
nor U11127 (N_11127,N_5534,N_7833);
and U11128 (N_11128,N_4714,N_4694);
or U11129 (N_11129,N_5322,N_7829);
xor U11130 (N_11130,N_6330,N_6152);
and U11131 (N_11131,N_7190,N_4302);
nor U11132 (N_11132,N_6771,N_7060);
nand U11133 (N_11133,N_7933,N_6216);
nor U11134 (N_11134,N_6007,N_5042);
nor U11135 (N_11135,N_7531,N_6476);
nand U11136 (N_11136,N_6779,N_5314);
xnor U11137 (N_11137,N_6815,N_4849);
nor U11138 (N_11138,N_7575,N_4120);
and U11139 (N_11139,N_6480,N_5446);
and U11140 (N_11140,N_4523,N_6079);
and U11141 (N_11141,N_7829,N_4500);
xnor U11142 (N_11142,N_7816,N_7911);
xnor U11143 (N_11143,N_4854,N_7727);
nor U11144 (N_11144,N_7554,N_6187);
and U11145 (N_11145,N_5418,N_4748);
nor U11146 (N_11146,N_6652,N_6756);
and U11147 (N_11147,N_4641,N_6766);
nor U11148 (N_11148,N_6746,N_5567);
nand U11149 (N_11149,N_5321,N_7642);
nor U11150 (N_11150,N_5949,N_7934);
nor U11151 (N_11151,N_7879,N_6135);
and U11152 (N_11152,N_5603,N_4097);
xnor U11153 (N_11153,N_5969,N_4786);
or U11154 (N_11154,N_5288,N_5987);
xor U11155 (N_11155,N_7753,N_4788);
nand U11156 (N_11156,N_5209,N_5936);
nor U11157 (N_11157,N_6748,N_6453);
nand U11158 (N_11158,N_4200,N_6674);
or U11159 (N_11159,N_7986,N_5350);
or U11160 (N_11160,N_5229,N_6123);
nor U11161 (N_11161,N_5435,N_6888);
xor U11162 (N_11162,N_4514,N_4327);
or U11163 (N_11163,N_7254,N_4884);
nor U11164 (N_11164,N_6029,N_6970);
xnor U11165 (N_11165,N_5353,N_6261);
or U11166 (N_11166,N_7463,N_5521);
nor U11167 (N_11167,N_6776,N_6323);
or U11168 (N_11168,N_4618,N_7194);
or U11169 (N_11169,N_6253,N_4463);
or U11170 (N_11170,N_5163,N_7112);
and U11171 (N_11171,N_5517,N_4472);
nor U11172 (N_11172,N_7757,N_5618);
or U11173 (N_11173,N_5600,N_5568);
xnor U11174 (N_11174,N_4276,N_4699);
xor U11175 (N_11175,N_7224,N_6411);
and U11176 (N_11176,N_5389,N_7184);
xnor U11177 (N_11177,N_7621,N_7856);
or U11178 (N_11178,N_6389,N_5661);
and U11179 (N_11179,N_7332,N_6302);
and U11180 (N_11180,N_6998,N_5189);
and U11181 (N_11181,N_7790,N_7935);
or U11182 (N_11182,N_6148,N_7511);
nor U11183 (N_11183,N_6035,N_7607);
or U11184 (N_11184,N_7612,N_6318);
or U11185 (N_11185,N_5204,N_4178);
or U11186 (N_11186,N_4790,N_7029);
nand U11187 (N_11187,N_6237,N_6739);
nand U11188 (N_11188,N_5574,N_7729);
and U11189 (N_11189,N_4021,N_6244);
and U11190 (N_11190,N_5924,N_4450);
xor U11191 (N_11191,N_4684,N_4840);
nand U11192 (N_11192,N_7755,N_4131);
or U11193 (N_11193,N_5070,N_4311);
and U11194 (N_11194,N_5076,N_5594);
nand U11195 (N_11195,N_4927,N_7317);
xnor U11196 (N_11196,N_4371,N_5378);
nand U11197 (N_11197,N_5592,N_7251);
and U11198 (N_11198,N_5221,N_7298);
and U11199 (N_11199,N_5358,N_4698);
nand U11200 (N_11200,N_7333,N_6636);
or U11201 (N_11201,N_5584,N_4758);
and U11202 (N_11202,N_6252,N_4919);
or U11203 (N_11203,N_7831,N_6033);
nor U11204 (N_11204,N_6810,N_6929);
and U11205 (N_11205,N_7539,N_7253);
nor U11206 (N_11206,N_5893,N_6020);
and U11207 (N_11207,N_6434,N_4137);
and U11208 (N_11208,N_4718,N_6740);
and U11209 (N_11209,N_6099,N_5977);
nand U11210 (N_11210,N_5947,N_4826);
and U11211 (N_11211,N_5289,N_5166);
and U11212 (N_11212,N_5622,N_4059);
nor U11213 (N_11213,N_5510,N_5975);
nor U11214 (N_11214,N_5995,N_4806);
or U11215 (N_11215,N_4516,N_4703);
xnor U11216 (N_11216,N_7038,N_4159);
nand U11217 (N_11217,N_7253,N_6818);
or U11218 (N_11218,N_6624,N_7807);
or U11219 (N_11219,N_5096,N_7991);
nand U11220 (N_11220,N_5097,N_4015);
nand U11221 (N_11221,N_6164,N_6089);
and U11222 (N_11222,N_7946,N_4396);
nand U11223 (N_11223,N_5512,N_4103);
nor U11224 (N_11224,N_6877,N_4596);
xor U11225 (N_11225,N_6654,N_5504);
nor U11226 (N_11226,N_5147,N_7230);
nand U11227 (N_11227,N_5105,N_4510);
xnor U11228 (N_11228,N_5218,N_7969);
and U11229 (N_11229,N_7269,N_4726);
and U11230 (N_11230,N_5651,N_7072);
or U11231 (N_11231,N_4516,N_6766);
nand U11232 (N_11232,N_6233,N_4145);
nand U11233 (N_11233,N_4444,N_5628);
or U11234 (N_11234,N_5922,N_4663);
nand U11235 (N_11235,N_7882,N_7707);
and U11236 (N_11236,N_7503,N_5269);
or U11237 (N_11237,N_5043,N_4209);
or U11238 (N_11238,N_6443,N_7266);
and U11239 (N_11239,N_4179,N_5276);
nand U11240 (N_11240,N_5007,N_4578);
nand U11241 (N_11241,N_7604,N_4095);
nor U11242 (N_11242,N_6372,N_5839);
and U11243 (N_11243,N_5683,N_5206);
or U11244 (N_11244,N_6943,N_7848);
nor U11245 (N_11245,N_4968,N_6528);
nor U11246 (N_11246,N_4004,N_5392);
nand U11247 (N_11247,N_7031,N_4163);
xor U11248 (N_11248,N_4682,N_4772);
nor U11249 (N_11249,N_6449,N_5529);
or U11250 (N_11250,N_5496,N_4051);
xnor U11251 (N_11251,N_4237,N_7218);
xor U11252 (N_11252,N_6977,N_4423);
and U11253 (N_11253,N_5206,N_4688);
or U11254 (N_11254,N_7667,N_6391);
nand U11255 (N_11255,N_7020,N_6735);
and U11256 (N_11256,N_4823,N_5800);
or U11257 (N_11257,N_6170,N_5637);
nor U11258 (N_11258,N_7609,N_4137);
nor U11259 (N_11259,N_4968,N_7289);
or U11260 (N_11260,N_7058,N_6180);
nor U11261 (N_11261,N_5823,N_4836);
nor U11262 (N_11262,N_6923,N_5644);
xnor U11263 (N_11263,N_7947,N_4439);
and U11264 (N_11264,N_6749,N_5883);
nand U11265 (N_11265,N_5638,N_7680);
nand U11266 (N_11266,N_6922,N_7501);
and U11267 (N_11267,N_7073,N_5151);
xnor U11268 (N_11268,N_7966,N_7386);
and U11269 (N_11269,N_4867,N_7803);
xnor U11270 (N_11270,N_4650,N_5766);
nand U11271 (N_11271,N_4006,N_5094);
and U11272 (N_11272,N_6547,N_6289);
nor U11273 (N_11273,N_6483,N_4382);
or U11274 (N_11274,N_4521,N_4148);
nor U11275 (N_11275,N_4086,N_4827);
and U11276 (N_11276,N_6283,N_4913);
nand U11277 (N_11277,N_4793,N_7747);
and U11278 (N_11278,N_5616,N_4081);
nor U11279 (N_11279,N_4102,N_5399);
nor U11280 (N_11280,N_5961,N_6448);
nor U11281 (N_11281,N_6587,N_7281);
and U11282 (N_11282,N_6564,N_7249);
and U11283 (N_11283,N_4129,N_7294);
and U11284 (N_11284,N_4946,N_7862);
nand U11285 (N_11285,N_6037,N_7988);
or U11286 (N_11286,N_6226,N_5757);
and U11287 (N_11287,N_7263,N_5823);
nand U11288 (N_11288,N_5629,N_7214);
nand U11289 (N_11289,N_6437,N_5634);
or U11290 (N_11290,N_6770,N_5537);
nor U11291 (N_11291,N_6237,N_7797);
and U11292 (N_11292,N_5224,N_7120);
nand U11293 (N_11293,N_7842,N_5051);
or U11294 (N_11294,N_6148,N_5220);
nand U11295 (N_11295,N_6887,N_6760);
and U11296 (N_11296,N_5794,N_5537);
xnor U11297 (N_11297,N_7868,N_6040);
or U11298 (N_11298,N_5266,N_5612);
or U11299 (N_11299,N_7056,N_6848);
or U11300 (N_11300,N_6403,N_4146);
nand U11301 (N_11301,N_7599,N_5201);
and U11302 (N_11302,N_7021,N_4128);
and U11303 (N_11303,N_5831,N_7399);
nand U11304 (N_11304,N_5135,N_5843);
and U11305 (N_11305,N_4422,N_6035);
xor U11306 (N_11306,N_5746,N_4180);
xor U11307 (N_11307,N_5744,N_7003);
nand U11308 (N_11308,N_6590,N_4399);
nand U11309 (N_11309,N_7134,N_6241);
xnor U11310 (N_11310,N_4377,N_4337);
nand U11311 (N_11311,N_5532,N_5704);
nor U11312 (N_11312,N_6552,N_5617);
nor U11313 (N_11313,N_5646,N_5952);
xnor U11314 (N_11314,N_4193,N_7388);
or U11315 (N_11315,N_7155,N_6100);
and U11316 (N_11316,N_6792,N_5684);
or U11317 (N_11317,N_4016,N_4362);
xnor U11318 (N_11318,N_7508,N_4373);
xnor U11319 (N_11319,N_4282,N_5567);
nor U11320 (N_11320,N_6633,N_6282);
or U11321 (N_11321,N_7859,N_7820);
xor U11322 (N_11322,N_6690,N_4859);
nand U11323 (N_11323,N_5304,N_5609);
and U11324 (N_11324,N_4641,N_4560);
or U11325 (N_11325,N_5493,N_5164);
or U11326 (N_11326,N_7433,N_7283);
or U11327 (N_11327,N_6101,N_4456);
or U11328 (N_11328,N_4410,N_5568);
nor U11329 (N_11329,N_7175,N_7778);
or U11330 (N_11330,N_5648,N_5965);
or U11331 (N_11331,N_6302,N_4004);
and U11332 (N_11332,N_7200,N_4516);
and U11333 (N_11333,N_6678,N_7253);
nand U11334 (N_11334,N_5340,N_7109);
or U11335 (N_11335,N_6736,N_5784);
and U11336 (N_11336,N_7121,N_6123);
xor U11337 (N_11337,N_4117,N_6940);
and U11338 (N_11338,N_7144,N_5244);
or U11339 (N_11339,N_6334,N_5972);
xnor U11340 (N_11340,N_6016,N_4819);
nor U11341 (N_11341,N_6435,N_5920);
and U11342 (N_11342,N_5242,N_6762);
and U11343 (N_11343,N_5686,N_5215);
or U11344 (N_11344,N_5086,N_5581);
nand U11345 (N_11345,N_4165,N_7837);
xnor U11346 (N_11346,N_6689,N_5654);
nor U11347 (N_11347,N_5261,N_5998);
nand U11348 (N_11348,N_5568,N_5478);
nor U11349 (N_11349,N_4847,N_7622);
and U11350 (N_11350,N_6175,N_5007);
or U11351 (N_11351,N_4436,N_7693);
and U11352 (N_11352,N_7123,N_5900);
and U11353 (N_11353,N_5465,N_6669);
nand U11354 (N_11354,N_5207,N_5316);
nand U11355 (N_11355,N_4244,N_6923);
and U11356 (N_11356,N_4307,N_7150);
or U11357 (N_11357,N_7952,N_5051);
xnor U11358 (N_11358,N_7553,N_4375);
or U11359 (N_11359,N_5574,N_4337);
and U11360 (N_11360,N_5486,N_4075);
nand U11361 (N_11361,N_7689,N_7593);
nand U11362 (N_11362,N_4874,N_6082);
nand U11363 (N_11363,N_7147,N_4379);
nand U11364 (N_11364,N_5764,N_6216);
nand U11365 (N_11365,N_5761,N_6359);
and U11366 (N_11366,N_4799,N_6987);
nand U11367 (N_11367,N_5708,N_7592);
and U11368 (N_11368,N_4614,N_7082);
nand U11369 (N_11369,N_5776,N_7949);
or U11370 (N_11370,N_7504,N_5281);
or U11371 (N_11371,N_7558,N_7204);
nand U11372 (N_11372,N_5377,N_5915);
and U11373 (N_11373,N_6613,N_5495);
and U11374 (N_11374,N_4385,N_6333);
and U11375 (N_11375,N_7609,N_7441);
xor U11376 (N_11376,N_7682,N_7794);
nand U11377 (N_11377,N_4135,N_5372);
and U11378 (N_11378,N_5810,N_4206);
nand U11379 (N_11379,N_5651,N_4671);
nor U11380 (N_11380,N_7808,N_6246);
nand U11381 (N_11381,N_7085,N_4751);
nor U11382 (N_11382,N_5243,N_4478);
or U11383 (N_11383,N_5849,N_6156);
or U11384 (N_11384,N_5228,N_4728);
and U11385 (N_11385,N_5802,N_7631);
and U11386 (N_11386,N_4158,N_7686);
and U11387 (N_11387,N_4449,N_5450);
nand U11388 (N_11388,N_7301,N_4677);
and U11389 (N_11389,N_4049,N_6064);
nand U11390 (N_11390,N_5642,N_7694);
nor U11391 (N_11391,N_5379,N_5323);
nand U11392 (N_11392,N_4163,N_4254);
and U11393 (N_11393,N_7150,N_6004);
nand U11394 (N_11394,N_5264,N_7752);
and U11395 (N_11395,N_6277,N_7051);
or U11396 (N_11396,N_4111,N_7439);
nand U11397 (N_11397,N_6513,N_7793);
or U11398 (N_11398,N_4938,N_6844);
or U11399 (N_11399,N_7552,N_6072);
nor U11400 (N_11400,N_7956,N_5491);
nor U11401 (N_11401,N_4012,N_4226);
nor U11402 (N_11402,N_6823,N_5484);
nand U11403 (N_11403,N_4715,N_4747);
nand U11404 (N_11404,N_4574,N_4405);
nor U11405 (N_11405,N_7628,N_4295);
or U11406 (N_11406,N_5259,N_4628);
nor U11407 (N_11407,N_7166,N_4185);
and U11408 (N_11408,N_7412,N_7834);
nor U11409 (N_11409,N_5279,N_7464);
xnor U11410 (N_11410,N_4052,N_5571);
or U11411 (N_11411,N_5083,N_6515);
nand U11412 (N_11412,N_7549,N_7533);
nand U11413 (N_11413,N_7473,N_6564);
nand U11414 (N_11414,N_4772,N_4307);
nor U11415 (N_11415,N_7143,N_6186);
and U11416 (N_11416,N_5799,N_6388);
and U11417 (N_11417,N_5456,N_4248);
nor U11418 (N_11418,N_6055,N_5901);
or U11419 (N_11419,N_4385,N_6926);
and U11420 (N_11420,N_4213,N_7114);
nor U11421 (N_11421,N_4290,N_5837);
nor U11422 (N_11422,N_7318,N_5589);
nand U11423 (N_11423,N_5665,N_7929);
nor U11424 (N_11424,N_6177,N_7193);
nand U11425 (N_11425,N_6762,N_6898);
xnor U11426 (N_11426,N_5574,N_4776);
xor U11427 (N_11427,N_4572,N_7433);
nor U11428 (N_11428,N_7423,N_6957);
nor U11429 (N_11429,N_6569,N_7689);
nand U11430 (N_11430,N_4422,N_6719);
nor U11431 (N_11431,N_4886,N_5069);
or U11432 (N_11432,N_4207,N_5463);
xor U11433 (N_11433,N_4441,N_7987);
and U11434 (N_11434,N_6786,N_7076);
nand U11435 (N_11435,N_6006,N_5869);
nor U11436 (N_11436,N_5440,N_5435);
nand U11437 (N_11437,N_6366,N_5816);
nor U11438 (N_11438,N_7188,N_7226);
nand U11439 (N_11439,N_7945,N_5206);
xor U11440 (N_11440,N_5062,N_6166);
nand U11441 (N_11441,N_5470,N_4118);
nand U11442 (N_11442,N_4370,N_6198);
nor U11443 (N_11443,N_5658,N_4447);
nor U11444 (N_11444,N_4330,N_7191);
and U11445 (N_11445,N_7208,N_7740);
xnor U11446 (N_11446,N_5490,N_4021);
and U11447 (N_11447,N_6654,N_5298);
or U11448 (N_11448,N_7463,N_6528);
and U11449 (N_11449,N_7477,N_4414);
or U11450 (N_11450,N_5673,N_7693);
nand U11451 (N_11451,N_7513,N_5902);
or U11452 (N_11452,N_4849,N_4731);
nor U11453 (N_11453,N_5495,N_7887);
xnor U11454 (N_11454,N_5376,N_5207);
and U11455 (N_11455,N_4298,N_6358);
or U11456 (N_11456,N_5339,N_6107);
or U11457 (N_11457,N_7090,N_6085);
nand U11458 (N_11458,N_5819,N_6808);
nand U11459 (N_11459,N_7045,N_7601);
or U11460 (N_11460,N_5938,N_6611);
xor U11461 (N_11461,N_7338,N_5362);
nand U11462 (N_11462,N_6642,N_7586);
xor U11463 (N_11463,N_6300,N_6898);
and U11464 (N_11464,N_6369,N_7109);
nor U11465 (N_11465,N_5611,N_7521);
or U11466 (N_11466,N_7819,N_7264);
nor U11467 (N_11467,N_4101,N_6965);
nor U11468 (N_11468,N_6251,N_4042);
nand U11469 (N_11469,N_6435,N_5068);
or U11470 (N_11470,N_5803,N_6722);
nand U11471 (N_11471,N_4775,N_4539);
nand U11472 (N_11472,N_5756,N_7548);
xor U11473 (N_11473,N_6294,N_4833);
or U11474 (N_11474,N_4084,N_7021);
or U11475 (N_11475,N_5316,N_7611);
nor U11476 (N_11476,N_6311,N_4840);
and U11477 (N_11477,N_4165,N_7799);
and U11478 (N_11478,N_6480,N_4094);
and U11479 (N_11479,N_7896,N_4907);
xor U11480 (N_11480,N_5543,N_4669);
xnor U11481 (N_11481,N_5752,N_5741);
nor U11482 (N_11482,N_7910,N_7224);
xor U11483 (N_11483,N_6326,N_6028);
and U11484 (N_11484,N_7699,N_6159);
and U11485 (N_11485,N_4418,N_5265);
xnor U11486 (N_11486,N_7427,N_6758);
nand U11487 (N_11487,N_6950,N_7737);
nor U11488 (N_11488,N_5586,N_6173);
and U11489 (N_11489,N_4945,N_6040);
or U11490 (N_11490,N_4894,N_4399);
and U11491 (N_11491,N_4023,N_4657);
nand U11492 (N_11492,N_5963,N_6398);
or U11493 (N_11493,N_4266,N_6658);
or U11494 (N_11494,N_7922,N_6295);
or U11495 (N_11495,N_5496,N_7310);
and U11496 (N_11496,N_7110,N_6935);
nand U11497 (N_11497,N_6359,N_7545);
and U11498 (N_11498,N_6062,N_6206);
nand U11499 (N_11499,N_5598,N_7864);
nand U11500 (N_11500,N_4408,N_6836);
nor U11501 (N_11501,N_7084,N_5302);
and U11502 (N_11502,N_4139,N_4932);
and U11503 (N_11503,N_7768,N_6669);
and U11504 (N_11504,N_5405,N_4744);
or U11505 (N_11505,N_7796,N_5994);
nand U11506 (N_11506,N_6730,N_7795);
and U11507 (N_11507,N_6409,N_5763);
nor U11508 (N_11508,N_7933,N_4835);
xor U11509 (N_11509,N_4423,N_7941);
and U11510 (N_11510,N_4230,N_5475);
or U11511 (N_11511,N_5402,N_5978);
and U11512 (N_11512,N_4990,N_6623);
xnor U11513 (N_11513,N_7821,N_6271);
and U11514 (N_11514,N_6954,N_6689);
and U11515 (N_11515,N_6386,N_5834);
xor U11516 (N_11516,N_4067,N_7460);
or U11517 (N_11517,N_5900,N_7188);
and U11518 (N_11518,N_7469,N_7046);
or U11519 (N_11519,N_7939,N_6367);
nand U11520 (N_11520,N_5575,N_4135);
nand U11521 (N_11521,N_6868,N_4242);
and U11522 (N_11522,N_4429,N_7444);
or U11523 (N_11523,N_5846,N_4032);
nand U11524 (N_11524,N_7768,N_7307);
and U11525 (N_11525,N_5909,N_7814);
and U11526 (N_11526,N_7393,N_4467);
nor U11527 (N_11527,N_4860,N_6232);
nor U11528 (N_11528,N_6410,N_6292);
and U11529 (N_11529,N_5186,N_7069);
nand U11530 (N_11530,N_6843,N_4598);
nor U11531 (N_11531,N_4507,N_5088);
or U11532 (N_11532,N_4750,N_5676);
xnor U11533 (N_11533,N_7597,N_6016);
nand U11534 (N_11534,N_5419,N_4172);
nor U11535 (N_11535,N_4348,N_7495);
or U11536 (N_11536,N_5919,N_6354);
or U11537 (N_11537,N_6909,N_4231);
nor U11538 (N_11538,N_5104,N_5031);
nand U11539 (N_11539,N_7937,N_5703);
and U11540 (N_11540,N_7575,N_5662);
or U11541 (N_11541,N_7423,N_6058);
and U11542 (N_11542,N_7490,N_4222);
nor U11543 (N_11543,N_5587,N_4652);
nand U11544 (N_11544,N_4056,N_5438);
nand U11545 (N_11545,N_6235,N_4277);
or U11546 (N_11546,N_7165,N_6280);
nand U11547 (N_11547,N_7504,N_6075);
and U11548 (N_11548,N_7648,N_5500);
and U11549 (N_11549,N_4477,N_5869);
or U11550 (N_11550,N_6632,N_5131);
and U11551 (N_11551,N_7467,N_4771);
nand U11552 (N_11552,N_6761,N_7274);
xor U11553 (N_11553,N_7131,N_7061);
nor U11554 (N_11554,N_7047,N_4187);
or U11555 (N_11555,N_5344,N_6561);
nand U11556 (N_11556,N_4070,N_4004);
nand U11557 (N_11557,N_5893,N_6151);
or U11558 (N_11558,N_4348,N_6128);
nor U11559 (N_11559,N_4824,N_7542);
nand U11560 (N_11560,N_4886,N_6740);
nand U11561 (N_11561,N_6498,N_7718);
and U11562 (N_11562,N_6695,N_4387);
and U11563 (N_11563,N_7813,N_6491);
or U11564 (N_11564,N_6418,N_5512);
or U11565 (N_11565,N_5656,N_7106);
and U11566 (N_11566,N_4520,N_4289);
and U11567 (N_11567,N_4045,N_6479);
and U11568 (N_11568,N_4501,N_6604);
and U11569 (N_11569,N_5287,N_4027);
nor U11570 (N_11570,N_5583,N_6949);
nor U11571 (N_11571,N_5287,N_6666);
nor U11572 (N_11572,N_6582,N_6168);
nand U11573 (N_11573,N_7888,N_6388);
xnor U11574 (N_11574,N_5232,N_5788);
and U11575 (N_11575,N_5685,N_4281);
or U11576 (N_11576,N_6760,N_7280);
and U11577 (N_11577,N_4553,N_7045);
nor U11578 (N_11578,N_5681,N_6315);
nand U11579 (N_11579,N_6422,N_7744);
nor U11580 (N_11580,N_4689,N_5341);
nand U11581 (N_11581,N_4498,N_6824);
nor U11582 (N_11582,N_7260,N_4442);
nor U11583 (N_11583,N_4371,N_4274);
xnor U11584 (N_11584,N_5871,N_7604);
and U11585 (N_11585,N_7128,N_5476);
xnor U11586 (N_11586,N_5921,N_6152);
nand U11587 (N_11587,N_7941,N_4935);
nor U11588 (N_11588,N_7814,N_5754);
or U11589 (N_11589,N_5602,N_7670);
nand U11590 (N_11590,N_6740,N_6657);
or U11591 (N_11591,N_4181,N_4979);
and U11592 (N_11592,N_5781,N_5228);
nand U11593 (N_11593,N_6575,N_7427);
nor U11594 (N_11594,N_4872,N_7592);
nor U11595 (N_11595,N_6522,N_6971);
nand U11596 (N_11596,N_6979,N_7566);
nand U11597 (N_11597,N_6329,N_6656);
xnor U11598 (N_11598,N_6296,N_4415);
nor U11599 (N_11599,N_7009,N_5872);
nor U11600 (N_11600,N_4557,N_7121);
nand U11601 (N_11601,N_4641,N_5877);
and U11602 (N_11602,N_7155,N_4788);
nand U11603 (N_11603,N_4558,N_4073);
or U11604 (N_11604,N_7878,N_5272);
nand U11605 (N_11605,N_5016,N_5487);
nand U11606 (N_11606,N_7249,N_4727);
or U11607 (N_11607,N_6482,N_4697);
and U11608 (N_11608,N_6692,N_5732);
and U11609 (N_11609,N_5344,N_5819);
and U11610 (N_11610,N_6293,N_7356);
and U11611 (N_11611,N_4428,N_4773);
nor U11612 (N_11612,N_6772,N_6328);
and U11613 (N_11613,N_5506,N_7573);
xor U11614 (N_11614,N_6510,N_4788);
or U11615 (N_11615,N_5709,N_7757);
nor U11616 (N_11616,N_5402,N_5298);
xor U11617 (N_11617,N_6860,N_6688);
and U11618 (N_11618,N_7058,N_4354);
or U11619 (N_11619,N_4958,N_4072);
nand U11620 (N_11620,N_5963,N_6294);
xor U11621 (N_11621,N_4954,N_7362);
xnor U11622 (N_11622,N_5571,N_6125);
nor U11623 (N_11623,N_6872,N_6290);
and U11624 (N_11624,N_6708,N_5449);
nor U11625 (N_11625,N_7378,N_5173);
and U11626 (N_11626,N_7187,N_4633);
and U11627 (N_11627,N_4310,N_6526);
nor U11628 (N_11628,N_6353,N_4207);
nand U11629 (N_11629,N_7582,N_6756);
and U11630 (N_11630,N_6007,N_5365);
or U11631 (N_11631,N_4996,N_7389);
and U11632 (N_11632,N_7832,N_7671);
or U11633 (N_11633,N_4520,N_6152);
or U11634 (N_11634,N_7982,N_7777);
and U11635 (N_11635,N_5376,N_5640);
nand U11636 (N_11636,N_7753,N_7938);
or U11637 (N_11637,N_4894,N_5551);
or U11638 (N_11638,N_6097,N_5200);
and U11639 (N_11639,N_4077,N_7834);
and U11640 (N_11640,N_6941,N_7011);
nand U11641 (N_11641,N_6726,N_4699);
and U11642 (N_11642,N_5030,N_4497);
nand U11643 (N_11643,N_5255,N_7653);
nand U11644 (N_11644,N_6864,N_4455);
nand U11645 (N_11645,N_4804,N_4385);
nand U11646 (N_11646,N_7680,N_5479);
nor U11647 (N_11647,N_4958,N_5644);
or U11648 (N_11648,N_5610,N_6697);
xor U11649 (N_11649,N_5710,N_4047);
xor U11650 (N_11650,N_6307,N_7349);
and U11651 (N_11651,N_4189,N_4424);
or U11652 (N_11652,N_7831,N_7826);
or U11653 (N_11653,N_7312,N_5692);
nand U11654 (N_11654,N_6428,N_7592);
or U11655 (N_11655,N_5119,N_5157);
and U11656 (N_11656,N_5892,N_7187);
and U11657 (N_11657,N_6814,N_4872);
and U11658 (N_11658,N_5511,N_7542);
nor U11659 (N_11659,N_7208,N_5168);
nor U11660 (N_11660,N_7474,N_6238);
or U11661 (N_11661,N_4456,N_6053);
and U11662 (N_11662,N_4099,N_4687);
or U11663 (N_11663,N_7769,N_4888);
nor U11664 (N_11664,N_4985,N_4475);
nor U11665 (N_11665,N_6313,N_4528);
or U11666 (N_11666,N_7350,N_4387);
and U11667 (N_11667,N_6097,N_4414);
nor U11668 (N_11668,N_5409,N_7329);
nor U11669 (N_11669,N_5005,N_4988);
nand U11670 (N_11670,N_6184,N_6978);
and U11671 (N_11671,N_6973,N_5705);
nor U11672 (N_11672,N_7485,N_5940);
and U11673 (N_11673,N_7924,N_4094);
xor U11674 (N_11674,N_6299,N_7457);
nor U11675 (N_11675,N_5041,N_7151);
or U11676 (N_11676,N_4214,N_6164);
and U11677 (N_11677,N_4001,N_4065);
nor U11678 (N_11678,N_4734,N_7565);
or U11679 (N_11679,N_4031,N_4676);
and U11680 (N_11680,N_6459,N_4148);
nor U11681 (N_11681,N_7904,N_7830);
and U11682 (N_11682,N_6287,N_5596);
nor U11683 (N_11683,N_6280,N_6004);
nor U11684 (N_11684,N_6438,N_4696);
and U11685 (N_11685,N_4898,N_6408);
nor U11686 (N_11686,N_7924,N_4879);
or U11687 (N_11687,N_4834,N_7913);
or U11688 (N_11688,N_6649,N_6803);
nand U11689 (N_11689,N_6883,N_4806);
or U11690 (N_11690,N_6668,N_4827);
and U11691 (N_11691,N_7632,N_4458);
nand U11692 (N_11692,N_4813,N_7778);
nand U11693 (N_11693,N_4044,N_7615);
nand U11694 (N_11694,N_7280,N_5306);
nand U11695 (N_11695,N_6607,N_4276);
nand U11696 (N_11696,N_6759,N_4268);
or U11697 (N_11697,N_6846,N_5214);
nor U11698 (N_11698,N_6137,N_5134);
and U11699 (N_11699,N_7940,N_5334);
nand U11700 (N_11700,N_4868,N_6491);
xor U11701 (N_11701,N_5199,N_4075);
and U11702 (N_11702,N_7255,N_7977);
or U11703 (N_11703,N_7263,N_5054);
nor U11704 (N_11704,N_5705,N_7667);
nor U11705 (N_11705,N_6364,N_5134);
nor U11706 (N_11706,N_7839,N_7549);
nand U11707 (N_11707,N_7792,N_6014);
nor U11708 (N_11708,N_7888,N_7924);
nand U11709 (N_11709,N_4044,N_6249);
and U11710 (N_11710,N_4385,N_4082);
nor U11711 (N_11711,N_7894,N_7478);
or U11712 (N_11712,N_4543,N_7126);
nand U11713 (N_11713,N_4385,N_5760);
nand U11714 (N_11714,N_7782,N_7094);
nor U11715 (N_11715,N_6269,N_7471);
and U11716 (N_11716,N_6491,N_6807);
nand U11717 (N_11717,N_6952,N_5656);
nor U11718 (N_11718,N_5373,N_4580);
nand U11719 (N_11719,N_4114,N_6031);
and U11720 (N_11720,N_7006,N_5084);
and U11721 (N_11721,N_7380,N_4302);
nor U11722 (N_11722,N_5088,N_7309);
or U11723 (N_11723,N_5820,N_6039);
xnor U11724 (N_11724,N_5717,N_5995);
or U11725 (N_11725,N_6490,N_7695);
nand U11726 (N_11726,N_5332,N_4771);
xnor U11727 (N_11727,N_5700,N_5605);
nor U11728 (N_11728,N_7065,N_6294);
and U11729 (N_11729,N_4679,N_6096);
nand U11730 (N_11730,N_5338,N_5883);
or U11731 (N_11731,N_7460,N_7887);
or U11732 (N_11732,N_5225,N_7884);
nand U11733 (N_11733,N_5370,N_5925);
and U11734 (N_11734,N_4068,N_4846);
xnor U11735 (N_11735,N_4416,N_6068);
nand U11736 (N_11736,N_7316,N_4138);
or U11737 (N_11737,N_4222,N_6815);
nor U11738 (N_11738,N_6393,N_4137);
nor U11739 (N_11739,N_6087,N_6263);
or U11740 (N_11740,N_7744,N_5895);
xor U11741 (N_11741,N_5161,N_4543);
and U11742 (N_11742,N_6804,N_5626);
nand U11743 (N_11743,N_7059,N_7215);
nand U11744 (N_11744,N_7438,N_4287);
nand U11745 (N_11745,N_4262,N_6596);
and U11746 (N_11746,N_5601,N_6877);
and U11747 (N_11747,N_7104,N_6030);
and U11748 (N_11748,N_7394,N_6669);
nand U11749 (N_11749,N_6442,N_7931);
nand U11750 (N_11750,N_6299,N_6832);
and U11751 (N_11751,N_7029,N_4358);
xor U11752 (N_11752,N_7758,N_7879);
and U11753 (N_11753,N_6892,N_6083);
nand U11754 (N_11754,N_4472,N_7936);
and U11755 (N_11755,N_4705,N_5324);
nand U11756 (N_11756,N_5414,N_7664);
or U11757 (N_11757,N_5218,N_5721);
nand U11758 (N_11758,N_7348,N_5595);
nor U11759 (N_11759,N_5962,N_5530);
nand U11760 (N_11760,N_5196,N_7359);
nor U11761 (N_11761,N_4469,N_5627);
xnor U11762 (N_11762,N_4279,N_4902);
and U11763 (N_11763,N_6366,N_7674);
nor U11764 (N_11764,N_6563,N_5572);
nor U11765 (N_11765,N_7450,N_5957);
nor U11766 (N_11766,N_6693,N_6123);
or U11767 (N_11767,N_5419,N_5389);
nor U11768 (N_11768,N_6568,N_7918);
or U11769 (N_11769,N_4066,N_5317);
nor U11770 (N_11770,N_4459,N_4856);
nor U11771 (N_11771,N_7189,N_4694);
nor U11772 (N_11772,N_7827,N_6441);
nor U11773 (N_11773,N_4724,N_4294);
xnor U11774 (N_11774,N_7319,N_6978);
and U11775 (N_11775,N_6196,N_5523);
and U11776 (N_11776,N_4118,N_5193);
xnor U11777 (N_11777,N_7826,N_7081);
and U11778 (N_11778,N_7826,N_6657);
or U11779 (N_11779,N_6869,N_6980);
nand U11780 (N_11780,N_7328,N_7039);
and U11781 (N_11781,N_6078,N_6302);
or U11782 (N_11782,N_6444,N_4610);
or U11783 (N_11783,N_4615,N_7322);
xor U11784 (N_11784,N_6586,N_5881);
and U11785 (N_11785,N_7618,N_5798);
or U11786 (N_11786,N_4273,N_6394);
and U11787 (N_11787,N_7008,N_7877);
or U11788 (N_11788,N_7955,N_7226);
nor U11789 (N_11789,N_7204,N_6020);
or U11790 (N_11790,N_6780,N_5237);
and U11791 (N_11791,N_7613,N_6832);
nor U11792 (N_11792,N_7210,N_4616);
xnor U11793 (N_11793,N_7900,N_7870);
and U11794 (N_11794,N_4171,N_6088);
or U11795 (N_11795,N_7092,N_5479);
and U11796 (N_11796,N_6090,N_7139);
and U11797 (N_11797,N_4328,N_7824);
nor U11798 (N_11798,N_7109,N_7318);
nor U11799 (N_11799,N_5488,N_7299);
nand U11800 (N_11800,N_6585,N_4477);
nand U11801 (N_11801,N_5530,N_5713);
nand U11802 (N_11802,N_4451,N_4009);
or U11803 (N_11803,N_6501,N_7333);
or U11804 (N_11804,N_7305,N_5634);
xor U11805 (N_11805,N_6467,N_7062);
nand U11806 (N_11806,N_4303,N_7567);
or U11807 (N_11807,N_7738,N_5412);
nand U11808 (N_11808,N_7175,N_7602);
nand U11809 (N_11809,N_6381,N_5829);
and U11810 (N_11810,N_5668,N_6650);
and U11811 (N_11811,N_5061,N_6386);
xor U11812 (N_11812,N_7229,N_6917);
and U11813 (N_11813,N_6407,N_4632);
and U11814 (N_11814,N_4420,N_5566);
nor U11815 (N_11815,N_7276,N_5209);
nor U11816 (N_11816,N_6569,N_6493);
or U11817 (N_11817,N_7455,N_6949);
and U11818 (N_11818,N_5770,N_6540);
nor U11819 (N_11819,N_7658,N_5688);
nor U11820 (N_11820,N_7244,N_4668);
and U11821 (N_11821,N_6584,N_7359);
nand U11822 (N_11822,N_6028,N_5439);
nor U11823 (N_11823,N_4619,N_6401);
and U11824 (N_11824,N_7398,N_6470);
and U11825 (N_11825,N_6346,N_5541);
and U11826 (N_11826,N_4394,N_4577);
and U11827 (N_11827,N_6021,N_6659);
or U11828 (N_11828,N_7357,N_7798);
nand U11829 (N_11829,N_4570,N_7184);
nand U11830 (N_11830,N_5344,N_5370);
nand U11831 (N_11831,N_5743,N_6629);
or U11832 (N_11832,N_6140,N_6506);
nor U11833 (N_11833,N_4674,N_6142);
nand U11834 (N_11834,N_4768,N_6660);
and U11835 (N_11835,N_7556,N_4474);
xnor U11836 (N_11836,N_6387,N_6677);
nand U11837 (N_11837,N_5331,N_4562);
nor U11838 (N_11838,N_7733,N_5674);
and U11839 (N_11839,N_7221,N_6129);
nand U11840 (N_11840,N_6930,N_5252);
or U11841 (N_11841,N_6656,N_7169);
nand U11842 (N_11842,N_4830,N_5478);
nand U11843 (N_11843,N_6413,N_5342);
or U11844 (N_11844,N_6921,N_6485);
nand U11845 (N_11845,N_4514,N_6705);
xor U11846 (N_11846,N_6175,N_5127);
and U11847 (N_11847,N_5907,N_4056);
and U11848 (N_11848,N_4297,N_5322);
and U11849 (N_11849,N_4826,N_4263);
or U11850 (N_11850,N_4362,N_6643);
and U11851 (N_11851,N_7460,N_5239);
or U11852 (N_11852,N_6340,N_7883);
or U11853 (N_11853,N_6118,N_6668);
or U11854 (N_11854,N_4949,N_7223);
nor U11855 (N_11855,N_7224,N_4377);
and U11856 (N_11856,N_6167,N_4813);
nor U11857 (N_11857,N_5028,N_4565);
nor U11858 (N_11858,N_6063,N_4418);
nand U11859 (N_11859,N_6602,N_5208);
nand U11860 (N_11860,N_5909,N_4387);
xor U11861 (N_11861,N_4974,N_4457);
and U11862 (N_11862,N_5689,N_5324);
nor U11863 (N_11863,N_6690,N_6459);
nor U11864 (N_11864,N_6210,N_7764);
and U11865 (N_11865,N_7632,N_7344);
or U11866 (N_11866,N_5796,N_5328);
and U11867 (N_11867,N_7495,N_7583);
nand U11868 (N_11868,N_5870,N_5142);
nor U11869 (N_11869,N_5455,N_7810);
nand U11870 (N_11870,N_5241,N_4077);
nand U11871 (N_11871,N_4434,N_4838);
and U11872 (N_11872,N_4412,N_5857);
nand U11873 (N_11873,N_6993,N_4636);
nand U11874 (N_11874,N_5627,N_5316);
or U11875 (N_11875,N_4736,N_7736);
nand U11876 (N_11876,N_5043,N_4007);
or U11877 (N_11877,N_7451,N_7031);
nand U11878 (N_11878,N_4521,N_5507);
and U11879 (N_11879,N_7556,N_4402);
and U11880 (N_11880,N_7786,N_4096);
and U11881 (N_11881,N_4319,N_6599);
nor U11882 (N_11882,N_5421,N_5635);
nor U11883 (N_11883,N_7416,N_4214);
xor U11884 (N_11884,N_5345,N_6717);
and U11885 (N_11885,N_6152,N_4055);
xnor U11886 (N_11886,N_4340,N_4920);
and U11887 (N_11887,N_4558,N_6915);
nand U11888 (N_11888,N_4101,N_7186);
or U11889 (N_11889,N_6845,N_6673);
nand U11890 (N_11890,N_7070,N_7673);
nor U11891 (N_11891,N_5264,N_6863);
xor U11892 (N_11892,N_5652,N_4530);
nor U11893 (N_11893,N_7187,N_6331);
and U11894 (N_11894,N_7685,N_6626);
and U11895 (N_11895,N_5872,N_6149);
and U11896 (N_11896,N_6352,N_6565);
nand U11897 (N_11897,N_4267,N_5351);
xor U11898 (N_11898,N_7411,N_7441);
and U11899 (N_11899,N_7706,N_6145);
or U11900 (N_11900,N_6606,N_5319);
and U11901 (N_11901,N_7299,N_4095);
and U11902 (N_11902,N_6109,N_4220);
and U11903 (N_11903,N_5946,N_5893);
or U11904 (N_11904,N_7516,N_5349);
nor U11905 (N_11905,N_7190,N_7441);
nand U11906 (N_11906,N_5306,N_4284);
nand U11907 (N_11907,N_5435,N_7769);
nand U11908 (N_11908,N_4155,N_5493);
nand U11909 (N_11909,N_4855,N_6915);
nor U11910 (N_11910,N_4431,N_7912);
and U11911 (N_11911,N_5150,N_4989);
or U11912 (N_11912,N_6661,N_6677);
nor U11913 (N_11913,N_5786,N_5672);
and U11914 (N_11914,N_5157,N_5242);
and U11915 (N_11915,N_6530,N_7930);
nor U11916 (N_11916,N_7327,N_5707);
and U11917 (N_11917,N_6798,N_7130);
nor U11918 (N_11918,N_6612,N_6411);
nor U11919 (N_11919,N_7544,N_5615);
nand U11920 (N_11920,N_4785,N_7731);
or U11921 (N_11921,N_4756,N_6426);
nand U11922 (N_11922,N_6061,N_5998);
and U11923 (N_11923,N_5630,N_7106);
nand U11924 (N_11924,N_7677,N_6020);
or U11925 (N_11925,N_7284,N_6125);
nor U11926 (N_11926,N_7879,N_6985);
nor U11927 (N_11927,N_4432,N_7445);
and U11928 (N_11928,N_6979,N_4662);
or U11929 (N_11929,N_5909,N_4960);
and U11930 (N_11930,N_5991,N_4659);
and U11931 (N_11931,N_4051,N_5970);
nor U11932 (N_11932,N_4662,N_5216);
nand U11933 (N_11933,N_4247,N_6082);
and U11934 (N_11934,N_6831,N_6310);
xor U11935 (N_11935,N_7093,N_7741);
nor U11936 (N_11936,N_5744,N_6814);
and U11937 (N_11937,N_5954,N_4685);
nand U11938 (N_11938,N_6268,N_4760);
or U11939 (N_11939,N_6111,N_7998);
nand U11940 (N_11940,N_4983,N_4215);
nand U11941 (N_11941,N_5728,N_7980);
or U11942 (N_11942,N_7481,N_7894);
and U11943 (N_11943,N_5209,N_5437);
or U11944 (N_11944,N_4299,N_4533);
nand U11945 (N_11945,N_6982,N_5056);
nor U11946 (N_11946,N_7361,N_4952);
and U11947 (N_11947,N_6752,N_7093);
and U11948 (N_11948,N_4421,N_5997);
or U11949 (N_11949,N_5993,N_4942);
and U11950 (N_11950,N_5110,N_5470);
and U11951 (N_11951,N_4529,N_6738);
nand U11952 (N_11952,N_5926,N_6787);
nor U11953 (N_11953,N_7796,N_5329);
or U11954 (N_11954,N_5330,N_7808);
and U11955 (N_11955,N_5103,N_4050);
xor U11956 (N_11956,N_5752,N_4631);
nand U11957 (N_11957,N_5877,N_5992);
or U11958 (N_11958,N_6585,N_6029);
and U11959 (N_11959,N_6794,N_5219);
and U11960 (N_11960,N_4892,N_5273);
nand U11961 (N_11961,N_7526,N_6463);
or U11962 (N_11962,N_6810,N_5828);
nand U11963 (N_11963,N_7093,N_7577);
xor U11964 (N_11964,N_7606,N_4539);
nand U11965 (N_11965,N_6215,N_4516);
nand U11966 (N_11966,N_6962,N_4209);
or U11967 (N_11967,N_7148,N_6380);
nand U11968 (N_11968,N_5504,N_6464);
nand U11969 (N_11969,N_5844,N_4077);
or U11970 (N_11970,N_7906,N_4654);
and U11971 (N_11971,N_6197,N_7176);
nor U11972 (N_11972,N_7182,N_5692);
nor U11973 (N_11973,N_5769,N_7791);
or U11974 (N_11974,N_5856,N_6680);
xnor U11975 (N_11975,N_4653,N_7596);
or U11976 (N_11976,N_7876,N_6109);
and U11977 (N_11977,N_4217,N_7905);
xor U11978 (N_11978,N_4749,N_6827);
nand U11979 (N_11979,N_6758,N_4397);
nand U11980 (N_11980,N_4502,N_5094);
nand U11981 (N_11981,N_6107,N_6980);
and U11982 (N_11982,N_5270,N_7774);
or U11983 (N_11983,N_7665,N_6286);
nand U11984 (N_11984,N_5850,N_5238);
or U11985 (N_11985,N_4168,N_4542);
and U11986 (N_11986,N_6667,N_5759);
xor U11987 (N_11987,N_6861,N_6028);
nand U11988 (N_11988,N_6504,N_6698);
and U11989 (N_11989,N_6612,N_7426);
nand U11990 (N_11990,N_5262,N_7081);
or U11991 (N_11991,N_4347,N_4587);
and U11992 (N_11992,N_5277,N_5177);
or U11993 (N_11993,N_7654,N_4727);
and U11994 (N_11994,N_7744,N_5542);
or U11995 (N_11995,N_4240,N_6810);
and U11996 (N_11996,N_4064,N_5646);
nor U11997 (N_11997,N_7458,N_7361);
nor U11998 (N_11998,N_6848,N_4775);
nand U11999 (N_11999,N_4808,N_6969);
nand U12000 (N_12000,N_9465,N_10846);
nand U12001 (N_12001,N_9998,N_9288);
or U12002 (N_12002,N_10763,N_8375);
and U12003 (N_12003,N_8793,N_9663);
or U12004 (N_12004,N_9383,N_9179);
or U12005 (N_12005,N_8177,N_9181);
and U12006 (N_12006,N_11419,N_10696);
nand U12007 (N_12007,N_9357,N_8234);
xnor U12008 (N_12008,N_9840,N_8500);
or U12009 (N_12009,N_8784,N_9162);
or U12010 (N_12010,N_11644,N_9964);
nand U12011 (N_12011,N_9106,N_8045);
and U12012 (N_12012,N_9767,N_11766);
or U12013 (N_12013,N_9248,N_11093);
nand U12014 (N_12014,N_9361,N_10707);
or U12015 (N_12015,N_9716,N_8438);
and U12016 (N_12016,N_10237,N_11333);
or U12017 (N_12017,N_9947,N_11487);
nor U12018 (N_12018,N_11116,N_9300);
and U12019 (N_12019,N_10184,N_8389);
nand U12020 (N_12020,N_9538,N_9630);
nor U12021 (N_12021,N_8964,N_10308);
nand U12022 (N_12022,N_11041,N_9305);
nand U12023 (N_12023,N_11143,N_9139);
or U12024 (N_12024,N_11294,N_9675);
and U12025 (N_12025,N_9384,N_9527);
or U12026 (N_12026,N_8312,N_9202);
nand U12027 (N_12027,N_9402,N_10716);
or U12028 (N_12028,N_9635,N_10810);
or U12029 (N_12029,N_10396,N_10080);
and U12030 (N_12030,N_8497,N_8086);
and U12031 (N_12031,N_9578,N_9397);
or U12032 (N_12032,N_10619,N_8037);
nand U12033 (N_12033,N_8049,N_8927);
or U12034 (N_12034,N_9223,N_11592);
xnor U12035 (N_12035,N_11400,N_10127);
or U12036 (N_12036,N_8236,N_8881);
and U12037 (N_12037,N_11296,N_11313);
nand U12038 (N_12038,N_10444,N_10056);
and U12039 (N_12039,N_8851,N_10286);
nand U12040 (N_12040,N_9283,N_11035);
or U12041 (N_12041,N_9647,N_8485);
nand U12042 (N_12042,N_9913,N_9270);
and U12043 (N_12043,N_11544,N_10424);
nor U12044 (N_12044,N_10465,N_11861);
nor U12045 (N_12045,N_10365,N_8939);
xor U12046 (N_12046,N_9791,N_10381);
nor U12047 (N_12047,N_11027,N_10828);
nor U12048 (N_12048,N_9793,N_9129);
nor U12049 (N_12049,N_11744,N_9028);
nor U12050 (N_12050,N_11841,N_9780);
nand U12051 (N_12051,N_9299,N_10743);
and U12052 (N_12052,N_9885,N_11546);
nand U12053 (N_12053,N_9001,N_10714);
or U12054 (N_12054,N_11600,N_11240);
or U12055 (N_12055,N_10000,N_8025);
nand U12056 (N_12056,N_10276,N_9726);
nor U12057 (N_12057,N_11016,N_9719);
nand U12058 (N_12058,N_8433,N_11922);
and U12059 (N_12059,N_8777,N_10524);
nand U12060 (N_12060,N_8783,N_10998);
nor U12061 (N_12061,N_9347,N_10339);
or U12062 (N_12062,N_10493,N_9467);
nand U12063 (N_12063,N_11479,N_8039);
xor U12064 (N_12064,N_10871,N_10126);
and U12065 (N_12065,N_8863,N_8709);
nor U12066 (N_12066,N_8085,N_11950);
or U12067 (N_12067,N_11739,N_9188);
nor U12068 (N_12068,N_11297,N_11439);
nor U12069 (N_12069,N_10712,N_8016);
nor U12070 (N_12070,N_8405,N_11295);
and U12071 (N_12071,N_8904,N_8144);
nor U12072 (N_12072,N_11945,N_9956);
and U12073 (N_12073,N_10477,N_11451);
and U12074 (N_12074,N_11475,N_9280);
or U12075 (N_12075,N_9441,N_10075);
nor U12076 (N_12076,N_8490,N_11241);
and U12077 (N_12077,N_8638,N_10136);
nand U12078 (N_12078,N_9433,N_10019);
nand U12079 (N_12079,N_8203,N_10672);
xnor U12080 (N_12080,N_11010,N_9083);
or U12081 (N_12081,N_11593,N_8183);
nor U12082 (N_12082,N_11008,N_9275);
or U12083 (N_12083,N_8191,N_11071);
xnor U12084 (N_12084,N_11534,N_8410);
nand U12085 (N_12085,N_10976,N_8316);
and U12086 (N_12086,N_9459,N_10020);
or U12087 (N_12087,N_10663,N_9134);
and U12088 (N_12088,N_11696,N_11166);
and U12089 (N_12089,N_11024,N_9651);
nand U12090 (N_12090,N_8298,N_10840);
nand U12091 (N_12091,N_8214,N_9395);
or U12092 (N_12092,N_10336,N_8816);
nor U12093 (N_12093,N_11216,N_10618);
and U12094 (N_12094,N_9566,N_10590);
or U12095 (N_12095,N_8984,N_9387);
nand U12096 (N_12096,N_8978,N_8237);
and U12097 (N_12097,N_11787,N_9727);
nand U12098 (N_12098,N_11520,N_9250);
nor U12099 (N_12099,N_11213,N_9611);
nor U12100 (N_12100,N_9479,N_9285);
or U12101 (N_12101,N_10287,N_11595);
nand U12102 (N_12102,N_11773,N_11290);
nor U12103 (N_12103,N_10397,N_9989);
nor U12104 (N_12104,N_11959,N_11690);
or U12105 (N_12105,N_9853,N_8598);
xnor U12106 (N_12106,N_11127,N_11536);
xor U12107 (N_12107,N_10166,N_8604);
or U12108 (N_12108,N_9512,N_8969);
nor U12109 (N_12109,N_9564,N_10596);
xor U12110 (N_12110,N_11459,N_8326);
or U12111 (N_12111,N_9468,N_9205);
nand U12112 (N_12112,N_11780,N_8911);
and U12113 (N_12113,N_9375,N_8390);
and U12114 (N_12114,N_9101,N_10503);
and U12115 (N_12115,N_8530,N_8213);
and U12116 (N_12116,N_8993,N_11556);
nand U12117 (N_12117,N_10558,N_9811);
or U12118 (N_12118,N_8593,N_8082);
xnor U12119 (N_12119,N_10082,N_11302);
nand U12120 (N_12120,N_10621,N_10173);
or U12121 (N_12121,N_11233,N_8714);
and U12122 (N_12122,N_8163,N_8317);
and U12123 (N_12123,N_8459,N_8658);
and U12124 (N_12124,N_8003,N_10710);
nand U12125 (N_12125,N_11303,N_10749);
or U12126 (N_12126,N_11506,N_11801);
or U12127 (N_12127,N_9581,N_9539);
nor U12128 (N_12128,N_8853,N_9152);
and U12129 (N_12129,N_9546,N_8131);
xor U12130 (N_12130,N_11443,N_11731);
nand U12131 (N_12131,N_10818,N_8865);
nor U12132 (N_12132,N_8648,N_11412);
or U12133 (N_12133,N_8513,N_11949);
nand U12134 (N_12134,N_9007,N_9355);
nor U12135 (N_12135,N_11114,N_11692);
and U12136 (N_12136,N_10108,N_8813);
and U12137 (N_12137,N_10335,N_9554);
nand U12138 (N_12138,N_10599,N_11624);
and U12139 (N_12139,N_10474,N_11620);
nor U12140 (N_12140,N_9379,N_9458);
and U12141 (N_12141,N_9303,N_11069);
or U12142 (N_12142,N_8992,N_10652);
and U12143 (N_12143,N_11853,N_11594);
or U12144 (N_12144,N_11613,N_8745);
and U12145 (N_12145,N_11401,N_11433);
nor U12146 (N_12146,N_10378,N_10701);
and U12147 (N_12147,N_8129,N_10057);
and U12148 (N_12148,N_8474,N_8948);
nor U12149 (N_12149,N_8182,N_11157);
nor U12150 (N_12150,N_8726,N_10333);
nor U12151 (N_12151,N_9960,N_10016);
nor U12152 (N_12152,N_10345,N_10757);
and U12153 (N_12153,N_10782,N_10122);
xor U12154 (N_12154,N_8636,N_10670);
nor U12155 (N_12155,N_11445,N_8437);
or U12156 (N_12156,N_10900,N_9660);
xnor U12157 (N_12157,N_8737,N_11524);
or U12158 (N_12158,N_9551,N_9757);
nand U12159 (N_12159,N_9605,N_8599);
xor U12160 (N_12160,N_10482,N_11695);
xnor U12161 (N_12161,N_10758,N_10880);
and U12162 (N_12162,N_11342,N_9157);
nand U12163 (N_12163,N_8041,N_9901);
xor U12164 (N_12164,N_8871,N_10984);
nand U12165 (N_12165,N_8616,N_10206);
and U12166 (N_12166,N_10901,N_11080);
or U12167 (N_12167,N_9213,N_10483);
or U12168 (N_12168,N_9484,N_11647);
and U12169 (N_12169,N_11628,N_8534);
nor U12170 (N_12170,N_8850,N_9813);
xor U12171 (N_12171,N_9431,N_8884);
or U12172 (N_12172,N_8882,N_10580);
nand U12173 (N_12173,N_9472,N_10198);
and U12174 (N_12174,N_11703,N_11381);
and U12175 (N_12175,N_8834,N_10827);
nor U12176 (N_12176,N_11153,N_10756);
nor U12177 (N_12177,N_11428,N_9087);
and U12178 (N_12178,N_9585,N_10935);
nand U12179 (N_12179,N_10191,N_8046);
nor U12180 (N_12180,N_11623,N_8702);
nand U12181 (N_12181,N_8098,N_11854);
or U12182 (N_12182,N_9600,N_9449);
nand U12183 (N_12183,N_11011,N_9615);
nand U12184 (N_12184,N_8220,N_9573);
nand U12185 (N_12185,N_10711,N_9323);
and U12186 (N_12186,N_8304,N_10594);
nand U12187 (N_12187,N_8968,N_10211);
nand U12188 (N_12188,N_9511,N_10414);
nand U12189 (N_12189,N_9750,N_8828);
nor U12190 (N_12190,N_9498,N_11037);
and U12191 (N_12191,N_9020,N_8716);
nor U12192 (N_12192,N_9473,N_8125);
nand U12193 (N_12193,N_9483,N_9827);
nand U12194 (N_12194,N_8914,N_10575);
nor U12195 (N_12195,N_10052,N_8178);
or U12196 (N_12196,N_9272,N_10263);
nor U12197 (N_12197,N_8071,N_9787);
nand U12198 (N_12198,N_10450,N_11305);
or U12199 (N_12199,N_8331,N_11847);
or U12200 (N_12200,N_11023,N_11700);
nand U12201 (N_12201,N_11872,N_8509);
xnor U12202 (N_12202,N_9273,N_8977);
and U12203 (N_12203,N_11043,N_8947);
and U12204 (N_12204,N_9343,N_10802);
and U12205 (N_12205,N_11179,N_8647);
nand U12206 (N_12206,N_10642,N_9783);
nor U12207 (N_12207,N_11525,N_8473);
nand U12208 (N_12208,N_8681,N_11065);
nor U12209 (N_12209,N_8337,N_10403);
and U12210 (N_12210,N_9871,N_8728);
xnor U12211 (N_12211,N_10447,N_8406);
or U12212 (N_12212,N_8276,N_9888);
nand U12213 (N_12213,N_8527,N_8376);
or U12214 (N_12214,N_8397,N_9359);
nor U12215 (N_12215,N_8916,N_10864);
and U12216 (N_12216,N_9426,N_11691);
and U12217 (N_12217,N_8357,N_8102);
xnor U12218 (N_12218,N_10819,N_11880);
or U12219 (N_12219,N_9768,N_8209);
or U12220 (N_12220,N_11809,N_11667);
nor U12221 (N_12221,N_10309,N_11927);
and U12222 (N_12222,N_9525,N_8832);
and U12223 (N_12223,N_9632,N_9386);
nand U12224 (N_12224,N_10844,N_9576);
nor U12225 (N_12225,N_8999,N_11588);
or U12226 (N_12226,N_8570,N_9860);
nand U12227 (N_12227,N_10167,N_9709);
nor U12228 (N_12228,N_9971,N_9494);
nand U12229 (N_12229,N_9341,N_8201);
and U12230 (N_12230,N_11911,N_9419);
and U12231 (N_12231,N_8836,N_8306);
nor U12232 (N_12232,N_11357,N_11490);
and U12233 (N_12233,N_10713,N_9666);
nand U12234 (N_12234,N_9688,N_8730);
nand U12235 (N_12235,N_11150,N_10692);
nand U12236 (N_12236,N_9646,N_8718);
nor U12237 (N_12237,N_8305,N_10364);
and U12238 (N_12238,N_9741,N_10165);
and U12239 (N_12239,N_9061,N_9259);
nand U12240 (N_12240,N_8496,N_11225);
nor U12241 (N_12241,N_9798,N_10574);
and U12242 (N_12242,N_8738,N_8552);
or U12243 (N_12243,N_11929,N_9540);
and U12244 (N_12244,N_11991,N_9580);
and U12245 (N_12245,N_10585,N_9126);
or U12246 (N_12246,N_9364,N_9905);
and U12247 (N_12247,N_10839,N_8385);
nand U12248 (N_12248,N_11317,N_11722);
xnor U12249 (N_12249,N_10028,N_10369);
and U12250 (N_12250,N_11109,N_9837);
nand U12251 (N_12251,N_9481,N_9969);
and U12252 (N_12252,N_10281,N_8244);
nand U12253 (N_12253,N_11148,N_11952);
or U12254 (N_12254,N_11259,N_9992);
nand U12255 (N_12255,N_11204,N_9194);
and U12256 (N_12256,N_10552,N_9808);
and U12257 (N_12257,N_9316,N_10491);
or U12258 (N_12258,N_11542,N_9409);
nor U12259 (N_12259,N_10650,N_9867);
and U12260 (N_12260,N_10374,N_10046);
or U12261 (N_12261,N_10469,N_8601);
nand U12262 (N_12262,N_10232,N_11777);
and U12263 (N_12263,N_8266,N_11115);
nand U12264 (N_12264,N_9346,N_11341);
nand U12265 (N_12265,N_10533,N_9211);
nor U12266 (N_12266,N_9477,N_9220);
and U12267 (N_12267,N_9993,N_10944);
and U12268 (N_12268,N_9671,N_9593);
nand U12269 (N_12269,N_11059,N_11774);
nand U12270 (N_12270,N_9046,N_8769);
nand U12271 (N_12271,N_10008,N_11319);
or U12272 (N_12272,N_10514,N_9940);
nor U12273 (N_12273,N_11382,N_8290);
or U12274 (N_12274,N_10736,N_11615);
or U12275 (N_12275,N_11423,N_11395);
or U12276 (N_12276,N_9936,N_10975);
or U12277 (N_12277,N_10139,N_9256);
nand U12278 (N_12278,N_8581,N_11481);
or U12279 (N_12279,N_9943,N_10578);
nor U12280 (N_12280,N_11285,N_10836);
and U12281 (N_12281,N_10732,N_11102);
or U12282 (N_12282,N_11476,N_11852);
nand U12283 (N_12283,N_9035,N_9064);
nor U12284 (N_12284,N_10305,N_10625);
nor U12285 (N_12285,N_9510,N_11310);
nand U12286 (N_12286,N_9985,N_8370);
nor U12287 (N_12287,N_10092,N_9369);
nor U12288 (N_12288,N_9542,N_8151);
or U12289 (N_12289,N_8380,N_9060);
xnor U12290 (N_12290,N_9980,N_8377);
or U12291 (N_12291,N_9563,N_9463);
nor U12292 (N_12292,N_10413,N_11374);
nor U12293 (N_12293,N_9487,N_10013);
and U12294 (N_12294,N_8631,N_11222);
and U12295 (N_12295,N_9855,N_8966);
xnor U12296 (N_12296,N_10107,N_10200);
or U12297 (N_12297,N_9655,N_11064);
nor U12298 (N_12298,N_9756,N_11616);
and U12299 (N_12299,N_10831,N_9167);
xor U12300 (N_12300,N_11420,N_11463);
nor U12301 (N_12301,N_8122,N_8486);
and U12302 (N_12302,N_9024,N_8367);
xnor U12303 (N_12303,N_9330,N_11752);
nor U12304 (N_12304,N_8619,N_10860);
and U12305 (N_12305,N_9720,N_8786);
or U12306 (N_12306,N_11768,N_10487);
and U12307 (N_12307,N_11858,N_9899);
nor U12308 (N_12308,N_10292,N_10768);
xnor U12309 (N_12309,N_8143,N_8983);
and U12310 (N_12310,N_8625,N_9521);
nand U12311 (N_12311,N_10683,N_10037);
nand U12312 (N_12312,N_9434,N_9242);
nand U12313 (N_12313,N_10517,N_10382);
nor U12314 (N_12314,N_10467,N_8195);
and U12315 (N_12315,N_11464,N_9037);
nand U12316 (N_12316,N_8760,N_11656);
and U12317 (N_12317,N_8642,N_8362);
or U12318 (N_12318,N_10848,N_8958);
nand U12319 (N_12319,N_8436,N_10176);
and U12320 (N_12320,N_11617,N_10603);
xnor U12321 (N_12321,N_11055,N_8303);
nand U12322 (N_12322,N_9959,N_9785);
and U12323 (N_12323,N_11688,N_10304);
and U12324 (N_12324,N_11005,N_11707);
nor U12325 (N_12325,N_10267,N_11376);
nor U12326 (N_12326,N_11121,N_10679);
nand U12327 (N_12327,N_10761,N_9495);
nor U12328 (N_12328,N_10180,N_8081);
nand U12329 (N_12329,N_10129,N_11640);
nand U12330 (N_12330,N_11020,N_11790);
nand U12331 (N_12331,N_10101,N_11203);
or U12332 (N_12332,N_10573,N_9643);
or U12333 (N_12333,N_11477,N_8259);
or U12334 (N_12334,N_8324,N_9416);
nor U12335 (N_12335,N_10722,N_9258);
or U12336 (N_12336,N_11794,N_10772);
nand U12337 (N_12337,N_8492,N_10079);
and U12338 (N_12338,N_11152,N_11194);
or U12339 (N_12339,N_11170,N_8193);
xor U12340 (N_12340,N_9407,N_11388);
nor U12341 (N_12341,N_9009,N_10589);
or U12342 (N_12342,N_8349,N_9047);
nand U12343 (N_12343,N_8652,N_9432);
nor U12344 (N_12344,N_11942,N_9862);
nand U12345 (N_12345,N_8704,N_10434);
or U12346 (N_12346,N_10560,N_8868);
or U12347 (N_12347,N_10155,N_11493);
and U12348 (N_12348,N_11432,N_9146);
nand U12349 (N_12349,N_10912,N_8336);
nor U12350 (N_12350,N_8613,N_10769);
xor U12351 (N_12351,N_8279,N_9200);
and U12352 (N_12352,N_10576,N_10423);
and U12353 (N_12353,N_10090,N_8132);
and U12354 (N_12354,N_9036,N_9382);
or U12355 (N_12355,N_9108,N_11834);
or U12356 (N_12356,N_9851,N_11648);
or U12357 (N_12357,N_10971,N_11226);
nor U12358 (N_12358,N_10217,N_8960);
xor U12359 (N_12359,N_10693,N_10706);
xnor U12360 (N_12360,N_8668,N_10620);
nand U12361 (N_12361,N_8525,N_10204);
nor U12362 (N_12362,N_9547,N_11119);
nor U12363 (N_12363,N_8764,N_10592);
xor U12364 (N_12364,N_10982,N_9849);
nor U12365 (N_12365,N_8857,N_9872);
and U12366 (N_12366,N_9529,N_11492);
xor U12367 (N_12367,N_9567,N_10432);
nand U12368 (N_12368,N_10197,N_8804);
nand U12369 (N_12369,N_10279,N_10437);
and U12370 (N_12370,N_10641,N_8514);
nand U12371 (N_12371,N_9881,N_11193);
and U12372 (N_12372,N_10032,N_11273);
nand U12373 (N_12373,N_8427,N_9360);
nand U12374 (N_12374,N_9310,N_11097);
nor U12375 (N_12375,N_8000,N_8185);
and U12376 (N_12376,N_9291,N_8054);
nor U12377 (N_12377,N_9640,N_10086);
nand U12378 (N_12378,N_11175,N_8695);
nor U12379 (N_12379,N_9986,N_11100);
xnor U12380 (N_12380,N_11753,N_8061);
nand U12381 (N_12381,N_8150,N_10132);
and U12382 (N_12382,N_11118,N_10402);
and U12383 (N_12383,N_11245,N_9678);
or U12384 (N_12384,N_8121,N_8651);
nand U12385 (N_12385,N_9894,N_9492);
xor U12386 (N_12386,N_11291,N_9889);
nand U12387 (N_12387,N_10087,N_9074);
and U12388 (N_12388,N_9313,N_9136);
or U12389 (N_12389,N_8249,N_11070);
and U12390 (N_12390,N_11304,N_11308);
and U12391 (N_12391,N_9208,N_9085);
nand U12392 (N_12392,N_10917,N_10881);
xor U12393 (N_12393,N_11772,N_8577);
or U12394 (N_12394,N_11047,N_9648);
nor U12395 (N_12395,N_10100,N_11239);
and U12396 (N_12396,N_11249,N_8562);
and U12397 (N_12397,N_9728,N_10440);
nor U12398 (N_12398,N_11701,N_10480);
xnor U12399 (N_12399,N_8284,N_10405);
xnor U12400 (N_12400,N_9760,N_9053);
and U12401 (N_12401,N_10653,N_11255);
or U12402 (N_12402,N_10609,N_10615);
or U12403 (N_12403,N_11084,N_10331);
or U12404 (N_12404,N_9598,N_9437);
and U12405 (N_12405,N_10608,N_10148);
or U12406 (N_12406,N_8140,N_10421);
or U12407 (N_12407,N_11257,N_9244);
nand U12408 (N_12408,N_10239,N_10992);
nand U12409 (N_12409,N_8751,N_10986);
and U12410 (N_12410,N_11403,N_8149);
nand U12411 (N_12411,N_10130,N_10829);
and U12412 (N_12412,N_9089,N_8488);
nor U12413 (N_12413,N_8949,N_11572);
or U12414 (N_12414,N_10376,N_9314);
xnor U12415 (N_12415,N_11545,N_8699);
nand U12416 (N_12416,N_10207,N_10518);
and U12417 (N_12417,N_9224,N_9026);
nand U12418 (N_12418,N_10416,N_8192);
or U12419 (N_12419,N_11456,N_10442);
and U12420 (N_12420,N_9017,N_9696);
and U12421 (N_12421,N_8797,N_11599);
or U12422 (N_12422,N_9027,N_9818);
nor U12423 (N_12423,N_8053,N_11919);
nand U12424 (N_12424,N_11930,N_10932);
or U12425 (N_12425,N_9826,N_8360);
nand U12426 (N_12426,N_10311,N_11651);
nor U12427 (N_12427,N_9311,N_8065);
xnor U12428 (N_12428,N_8088,N_9717);
nor U12429 (N_12429,N_11377,N_11621);
nand U12430 (N_12430,N_9245,N_9592);
or U12431 (N_12431,N_8494,N_8050);
or U12432 (N_12432,N_9486,N_8471);
and U12433 (N_12433,N_11947,N_11817);
or U12434 (N_12434,N_9874,N_9625);
nor U12435 (N_12435,N_9496,N_11888);
xor U12436 (N_12436,N_11349,N_9955);
or U12437 (N_12437,N_11923,N_10938);
nor U12438 (N_12438,N_10577,N_11253);
nand U12439 (N_12439,N_11968,N_10225);
nand U12440 (N_12440,N_10581,N_10337);
xnor U12441 (N_12441,N_10520,N_11737);
or U12442 (N_12442,N_8844,N_9620);
and U12443 (N_12443,N_9264,N_11045);
or U12444 (N_12444,N_8021,N_11778);
and U12445 (N_12445,N_9081,N_10168);
xor U12446 (N_12446,N_8837,N_10522);
nand U12447 (N_12447,N_9044,N_11474);
nor U12448 (N_12448,N_11346,N_10956);
and U12449 (N_12449,N_8168,N_10586);
nand U12450 (N_12450,N_11606,N_10728);
nand U12451 (N_12451,N_11575,N_10216);
nand U12452 (N_12452,N_10505,N_9192);
and U12453 (N_12453,N_8062,N_8624);
nor U12454 (N_12454,N_9105,N_10438);
nand U12455 (N_12455,N_11279,N_11563);
xnor U12456 (N_12456,N_11960,N_10298);
or U12457 (N_12457,N_11073,N_8369);
nand U12458 (N_12458,N_8734,N_8395);
and U12459 (N_12459,N_11026,N_9684);
or U12460 (N_12460,N_8590,N_9110);
and U12461 (N_12461,N_11992,N_9196);
nand U12462 (N_12462,N_8152,N_10024);
nand U12463 (N_12463,N_10564,N_10835);
nor U12464 (N_12464,N_8650,N_9619);
and U12465 (N_12465,N_10435,N_10534);
nand U12466 (N_12466,N_9987,N_9673);
or U12467 (N_12467,N_10041,N_11601);
nand U12468 (N_12468,N_10513,N_9831);
nor U12469 (N_12469,N_10995,N_9095);
and U12470 (N_12470,N_8645,N_10053);
xnor U12471 (N_12471,N_10118,N_10675);
nand U12472 (N_12472,N_10242,N_11495);
nand U12473 (N_12473,N_8399,N_10913);
nor U12474 (N_12474,N_11881,N_8972);
nand U12475 (N_12475,N_11028,N_8394);
or U12476 (N_12476,N_9925,N_11828);
or U12477 (N_12477,N_8603,N_11658);
or U12478 (N_12478,N_9802,N_10955);
nor U12479 (N_12479,N_10735,N_9507);
and U12480 (N_12480,N_9832,N_11709);
or U12481 (N_12481,N_9003,N_8515);
nand U12482 (N_12482,N_8216,N_11404);
or U12483 (N_12483,N_10760,N_10636);
or U12484 (N_12484,N_9518,N_10627);
nor U12485 (N_12485,N_9412,N_9586);
and U12486 (N_12486,N_8678,N_10762);
or U12487 (N_12487,N_9623,N_10770);
nand U12488 (N_12488,N_11725,N_10948);
xor U12489 (N_12489,N_8897,N_11939);
and U12490 (N_12490,N_8371,N_10094);
nor U12491 (N_12491,N_9772,N_9921);
or U12492 (N_12492,N_9506,N_11156);
xnor U12493 (N_12493,N_10822,N_10776);
nor U12494 (N_12494,N_8372,N_9394);
nand U12495 (N_12495,N_9160,N_8923);
xor U12496 (N_12496,N_8103,N_11164);
xnor U12497 (N_12497,N_9180,N_8011);
or U12498 (N_12498,N_11670,N_10326);
nand U12499 (N_12499,N_9251,N_9191);
and U12500 (N_12500,N_8523,N_9902);
nor U12501 (N_12501,N_11887,N_10143);
nand U12502 (N_12502,N_11642,N_11356);
or U12503 (N_12503,N_9637,N_11051);
or U12504 (N_12504,N_9657,N_11176);
and U12505 (N_12505,N_9092,N_10657);
nor U12506 (N_12506,N_10492,N_11824);
nand U12507 (N_12507,N_8456,N_9603);
or U12508 (N_12508,N_8339,N_9005);
or U12509 (N_12509,N_8484,N_9363);
nand U12510 (N_12510,N_11999,N_11315);
xor U12511 (N_12511,N_9173,N_9878);
nor U12512 (N_12512,N_10791,N_11364);
and U12513 (N_12513,N_8556,N_10297);
nand U12514 (N_12514,N_10027,N_9935);
nor U12515 (N_12515,N_10417,N_11147);
nor U12516 (N_12516,N_10865,N_11533);
and U12517 (N_12517,N_10799,N_10395);
nor U12518 (N_12518,N_8020,N_11316);
and U12519 (N_12519,N_11675,N_10549);
nand U12520 (N_12520,N_10060,N_8340);
nand U12521 (N_12521,N_11622,N_8172);
and U12522 (N_12522,N_10315,N_11091);
and U12523 (N_12523,N_9296,N_8166);
or U12524 (N_12524,N_11272,N_11483);
xor U12525 (N_12525,N_10384,N_10571);
nand U12526 (N_12526,N_8073,N_9759);
and U12527 (N_12527,N_11275,N_9252);
nand U12528 (N_12528,N_9743,N_9286);
or U12529 (N_12529,N_8169,N_10222);
xor U12530 (N_12530,N_8611,N_8950);
nor U12531 (N_12531,N_9503,N_11365);
xor U12532 (N_12532,N_9777,N_11212);
nand U12533 (N_12533,N_9910,N_8123);
or U12534 (N_12534,N_9634,N_8566);
nor U12535 (N_12535,N_11025,N_9163);
and U12536 (N_12536,N_8731,N_10527);
nand U12537 (N_12537,N_10502,N_10669);
and U12538 (N_12538,N_8398,N_9983);
nand U12539 (N_12539,N_11618,N_10656);
and U12540 (N_12540,N_8812,N_10039);
nand U12541 (N_12541,N_11396,N_10613);
and U12542 (N_12542,N_10065,N_8956);
or U12543 (N_12543,N_10379,N_8318);
and U12544 (N_12544,N_10733,N_10662);
nand U12545 (N_12545,N_8447,N_10295);
and U12546 (N_12546,N_10346,N_8986);
nand U12547 (N_12547,N_11502,N_8781);
or U12548 (N_12548,N_10241,N_8971);
nand U12549 (N_12549,N_10996,N_8198);
nand U12550 (N_12550,N_9923,N_9471);
nor U12551 (N_12551,N_10389,N_8898);
and U12552 (N_12552,N_9842,N_8133);
or U12553 (N_12553,N_9297,N_10358);
or U12554 (N_12554,N_9282,N_10705);
and U12555 (N_12555,N_9415,N_9099);
nor U12556 (N_12556,N_11230,N_10754);
and U12557 (N_12557,N_10076,N_9672);
nand U12558 (N_12558,N_11450,N_11174);
and U12559 (N_12559,N_10660,N_8481);
nand U12560 (N_12560,N_8040,N_11636);
and U12561 (N_12561,N_10189,N_8479);
nand U12562 (N_12562,N_9774,N_10545);
nor U12563 (N_12563,N_8345,N_8024);
nand U12564 (N_12564,N_10431,N_9833);
nand U12565 (N_12565,N_8811,N_8374);
nand U12566 (N_12566,N_10957,N_11605);
and U12567 (N_12567,N_11775,N_8869);
nor U12568 (N_12568,N_10853,N_9107);
xnor U12569 (N_12569,N_11229,N_11387);
or U12570 (N_12570,N_11271,N_11815);
nor U12571 (N_12571,N_9939,N_8520);
nor U12572 (N_12572,N_8157,N_11111);
nor U12573 (N_12573,N_10813,N_11472);
and U12574 (N_12574,N_10348,N_10426);
and U12575 (N_12575,N_8270,N_8981);
nor U12576 (N_12576,N_11014,N_10746);
nor U12577 (N_12577,N_11705,N_8944);
xnor U12578 (N_12578,N_10209,N_8591);
nor U12579 (N_12579,N_9979,N_8917);
nor U12580 (N_12580,N_8356,N_10099);
nand U12581 (N_12581,N_10473,N_9156);
or U12582 (N_12582,N_9978,N_9873);
or U12583 (N_12583,N_11454,N_10767);
nor U12584 (N_12584,N_8892,N_10805);
or U12585 (N_12585,N_10678,N_11610);
nor U12586 (N_12586,N_9765,N_8124);
or U12587 (N_12587,N_8240,N_8655);
or U12588 (N_12588,N_8014,N_9420);
xnor U12589 (N_12589,N_8779,N_11082);
and U12590 (N_12590,N_8495,N_8221);
or U12591 (N_12591,N_10089,N_11218);
nand U12592 (N_12592,N_8444,N_8013);
nand U12593 (N_12593,N_10734,N_10457);
and U12594 (N_12594,N_8368,N_9941);
nor U12595 (N_12595,N_11154,N_8359);
or U12596 (N_12596,N_11083,N_11738);
or U12597 (N_12597,N_9400,N_8592);
or U12598 (N_12598,N_11321,N_8285);
nand U12599 (N_12599,N_10918,N_11602);
nor U12600 (N_12600,N_8223,N_9924);
nor U12601 (N_12601,N_11711,N_9770);
or U12602 (N_12602,N_9976,N_11567);
nand U12603 (N_12603,N_8239,N_8818);
or U12604 (N_12604,N_11674,N_8864);
nor U12605 (N_12605,N_9870,N_9414);
and U12606 (N_12606,N_8211,N_8557);
xnor U12607 (N_12607,N_8194,N_10147);
and U12608 (N_12608,N_8711,N_10651);
xor U12609 (N_12609,N_8396,N_9591);
nor U12610 (N_12610,N_8788,N_11827);
nand U12611 (N_12611,N_9649,N_10591);
xnor U12612 (N_12612,N_11223,N_8623);
and U12613 (N_12613,N_9689,N_11266);
or U12614 (N_12614,N_11513,N_8031);
or U12615 (N_12615,N_11948,N_10385);
nand U12616 (N_12616,N_8412,N_9218);
nand U12617 (N_12617,N_11105,N_11029);
or U12618 (N_12618,N_11748,N_9307);
nand U12619 (N_12619,N_8036,N_11870);
nand U12620 (N_12620,N_11970,N_9763);
xnor U12621 (N_12621,N_9879,N_9429);
and U12622 (N_12622,N_8549,N_9493);
nand U12623 (N_12623,N_8400,N_11384);
nor U12624 (N_12624,N_11783,N_11391);
and U12625 (N_12625,N_8856,N_11362);
nand U12626 (N_12626,N_10792,N_11301);
or U12627 (N_12627,N_10238,N_10121);
nand U12628 (N_12628,N_8289,N_8895);
nand U12629 (N_12629,N_9175,N_9701);
nor U12630 (N_12630,N_11458,N_11246);
nor U12631 (N_12631,N_10720,N_8142);
nor U12632 (N_12632,N_10464,N_11980);
and U12633 (N_12633,N_11836,N_11438);
xnor U12634 (N_12634,N_8661,N_11771);
nor U12635 (N_12635,N_8894,N_9755);
xnor U12636 (N_12636,N_8536,N_8826);
and U12637 (N_12637,N_9158,N_9775);
nand U12638 (N_12638,N_11838,N_10563);
nand U12639 (N_12639,N_9690,N_10436);
nor U12640 (N_12640,N_11580,N_11159);
nand U12641 (N_12641,N_11351,N_11471);
nand U12642 (N_12642,N_9948,N_10759);
or U12643 (N_12643,N_10507,N_8967);
or U12644 (N_12644,N_9809,N_10624);
nand U12645 (N_12645,N_10610,N_8671);
and U12646 (N_12646,N_8663,N_11633);
or U12647 (N_12647,N_9875,N_10058);
and U12648 (N_12648,N_11724,N_10296);
nand U12649 (N_12649,N_11684,N_8344);
and U12650 (N_12650,N_10872,N_8159);
and U12651 (N_12651,N_10497,N_10318);
xnor U12652 (N_12652,N_10428,N_9219);
nor U12653 (N_12653,N_11925,N_9088);
and U12654 (N_12654,N_11372,N_10149);
or U12655 (N_12655,N_11679,N_10157);
and U12656 (N_12656,N_10902,N_9398);
and U12657 (N_12657,N_8935,N_8775);
nor U12658 (N_12658,N_8245,N_11088);
and U12659 (N_12659,N_8439,N_8342);
and U12660 (N_12660,N_11619,N_9676);
and U12661 (N_12661,N_9221,N_9558);
and U12662 (N_12662,N_9098,N_9408);
nor U12663 (N_12663,N_11900,N_9735);
nand U12664 (N_12664,N_10458,N_9896);
xnor U12665 (N_12665,N_8921,N_11289);
or U12666 (N_12666,N_11375,N_11576);
nor U12667 (N_12667,N_10150,N_10408);
xor U12668 (N_12668,N_10883,N_8996);
nor U12669 (N_12669,N_9844,N_9700);
and U12670 (N_12670,N_11671,N_8130);
or U12671 (N_12671,N_10949,N_10074);
or U12672 (N_12672,N_11205,N_9893);
or U12673 (N_12673,N_9570,N_10934);
nor U12674 (N_12674,N_10821,N_11306);
and U12675 (N_12675,N_9583,N_11369);
nand U12676 (N_12676,N_10877,N_9730);
or U12677 (N_12677,N_8033,N_9550);
nand U12678 (N_12678,N_11762,N_8461);
and U12679 (N_12679,N_11270,N_9002);
xor U12680 (N_12680,N_9410,N_9544);
nor U12681 (N_12681,N_11687,N_11158);
nand U12682 (N_12682,N_11448,N_8888);
or U12683 (N_12683,N_10499,N_11050);
or U12684 (N_12684,N_8468,N_8548);
and U12685 (N_12685,N_8112,N_8723);
and U12686 (N_12686,N_8454,N_9066);
xor U12687 (N_12687,N_9466,N_8970);
nor U12688 (N_12688,N_10271,N_10164);
and U12689 (N_12689,N_8026,N_10034);
xnor U12690 (N_12690,N_9253,N_11200);
and U12691 (N_12691,N_11281,N_10380);
or U12692 (N_12692,N_8134,N_10419);
nand U12693 (N_12693,N_11188,N_9895);
or U12694 (N_12694,N_8629,N_10889);
nor U12695 (N_12695,N_10774,N_9920);
nand U12696 (N_12696,N_8409,N_11017);
or U12697 (N_12697,N_8578,N_8105);
nor U12698 (N_12698,N_8408,N_10059);
nor U12699 (N_12699,N_11682,N_8379);
nand U12700 (N_12700,N_10715,N_8338);
nor U12701 (N_12701,N_10826,N_11574);
or U12702 (N_12702,N_11565,N_10634);
or U12703 (N_12703,N_10302,N_11117);
and U12704 (N_12704,N_9413,N_10231);
nand U12705 (N_12705,N_11747,N_11803);
and U12706 (N_12706,N_10694,N_8429);
nand U12707 (N_12707,N_11087,N_8156);
and U12708 (N_12708,N_8847,N_10373);
nand U12709 (N_12709,N_10366,N_11585);
xor U12710 (N_12710,N_8262,N_10054);
nor U12711 (N_12711,N_11873,N_11857);
and U12712 (N_12712,N_11799,N_11486);
nor U12713 (N_12713,N_11363,N_11081);
nand U12714 (N_12714,N_11373,N_8343);
or U12715 (N_12715,N_11046,N_11631);
nor U12716 (N_12716,N_11664,N_11066);
or U12717 (N_12717,N_9900,N_9556);
nand U12718 (N_12718,N_9277,N_11535);
and U12719 (N_12719,N_9533,N_11800);
or U12720 (N_12720,N_11324,N_11044);
xnor U12721 (N_12721,N_10055,N_11981);
nand U12722 (N_12722,N_10637,N_11899);
and U12723 (N_12723,N_9612,N_10354);
and U12724 (N_12724,N_10192,N_8776);
or U12725 (N_12725,N_11979,N_9997);
or U12726 (N_12726,N_8703,N_10486);
nand U12727 (N_12727,N_10879,N_11425);
or U12728 (N_12728,N_10851,N_11639);
and U12729 (N_12729,N_8720,N_11522);
nand U12730 (N_12730,N_10541,N_11446);
or U12731 (N_12731,N_10855,N_9267);
nor U12732 (N_12732,N_10033,N_8256);
nor U12733 (N_12733,N_8780,N_8038);
and U12734 (N_12734,N_10832,N_10698);
nand U12735 (N_12735,N_8962,N_10867);
nor U12736 (N_12736,N_10868,N_10806);
and U12737 (N_12737,N_8846,N_8043);
nor U12738 (N_12738,N_10042,N_9548);
and U12739 (N_12739,N_10936,N_9736);
or U12740 (N_12740,N_11751,N_10301);
or U12741 (N_12741,N_10259,N_8982);
or U12742 (N_12742,N_11996,N_9012);
or U12743 (N_12743,N_9464,N_11136);
nand U12744 (N_12744,N_9707,N_9589);
xnor U12745 (N_12745,N_10842,N_9949);
nor U12746 (N_12746,N_9794,N_11661);
or U12747 (N_12747,N_9990,N_11819);
and U12748 (N_12748,N_9752,N_10562);
or U12749 (N_12749,N_11498,N_8633);
or U12750 (N_12750,N_8170,N_8874);
or U12751 (N_12751,N_8990,N_11846);
nor U12752 (N_12752,N_10245,N_11267);
and U12753 (N_12753,N_11178,N_8540);
nor U12754 (N_12754,N_10962,N_11839);
nand U12755 (N_12755,N_9662,N_10771);
xnor U12756 (N_12756,N_9519,N_11795);
nand U12757 (N_12757,N_9132,N_10006);
and U12758 (N_12758,N_9151,N_10597);
nor U12759 (N_12759,N_10980,N_10540);
or U12760 (N_12760,N_10249,N_9608);
nand U12761 (N_12761,N_11577,N_9816);
nand U12762 (N_12762,N_9358,N_9193);
nor U12763 (N_12763,N_8586,N_8567);
nor U12764 (N_12764,N_8052,N_11033);
nor U12765 (N_12765,N_8934,N_8539);
nor U12766 (N_12766,N_11672,N_11039);
xor U12767 (N_12767,N_11825,N_10638);
xnor U12768 (N_12768,N_10282,N_10970);
nor U12769 (N_12769,N_10208,N_9169);
nand U12770 (N_12770,N_9999,N_9504);
nor U12771 (N_12771,N_8146,N_10151);
or U12772 (N_12772,N_11263,N_10617);
nor U12773 (N_12773,N_10886,N_11882);
nor U12774 (N_12774,N_10911,N_10113);
nand U12775 (N_12775,N_8354,N_10030);
xnor U12776 (N_12776,N_9056,N_10448);
or U12777 (N_12777,N_8684,N_10285);
or U12778 (N_12778,N_8765,N_8579);
xor U12779 (N_12779,N_9515,N_10789);
nand U12780 (N_12780,N_10943,N_11591);
xnor U12781 (N_12781,N_11860,N_10676);
or U12782 (N_12782,N_9025,N_10223);
and U12783 (N_12783,N_11352,N_8985);
and U12784 (N_12784,N_9930,N_9255);
xnor U12785 (N_12785,N_10884,N_9232);
or U12786 (N_12786,N_8278,N_9929);
nand U12787 (N_12787,N_11826,N_8792);
nand U12788 (N_12788,N_10171,N_10658);
nor U12789 (N_12789,N_10745,N_10390);
xor U12790 (N_12790,N_10025,N_10070);
nor U12791 (N_12791,N_8600,N_10084);
or U12792 (N_12792,N_11300,N_10644);
and U12793 (N_12793,N_10343,N_10510);
or U12794 (N_12794,N_10370,N_11250);
and U12795 (N_12795,N_9238,N_9376);
nand U12796 (N_12796,N_8424,N_9804);
or U12797 (N_12797,N_8622,N_11764);
or U12798 (N_12798,N_10026,N_8012);
or U12799 (N_12799,N_9128,N_9008);
nand U12800 (N_12800,N_8618,N_8452);
nor U12801 (N_12801,N_8323,N_9500);
and U12802 (N_12802,N_8487,N_8363);
and U12803 (N_12803,N_9805,N_11569);
nand U12804 (N_12804,N_9938,N_8758);
nand U12805 (N_12805,N_8582,N_8640);
or U12806 (N_12806,N_8936,N_11074);
nand U12807 (N_12807,N_10233,N_10471);
and U12808 (N_12808,N_10461,N_11151);
nand U12809 (N_12809,N_8348,N_8809);
and U12810 (N_12810,N_11537,N_10063);
nand U12811 (N_12811,N_8924,N_9958);
nor U12812 (N_12812,N_10035,N_9751);
xnor U12813 (N_12813,N_8407,N_9077);
nor U12814 (N_12814,N_8426,N_8091);
nand U12815 (N_12815,N_11413,N_10340);
nand U12816 (N_12816,N_11969,N_10324);
nand U12817 (N_12817,N_9290,N_11864);
nor U12818 (N_12818,N_11370,N_8879);
or U12819 (N_12819,N_8995,N_9182);
xnor U12820 (N_12820,N_11385,N_9829);
or U12821 (N_12821,N_8908,N_8228);
nand U12822 (N_12822,N_9198,N_10102);
and U12823 (N_12823,N_11217,N_9292);
nand U12824 (N_12824,N_10300,N_10188);
nor U12825 (N_12825,N_8997,N_8698);
and U12826 (N_12826,N_11890,N_9071);
nor U12827 (N_12827,N_11729,N_11095);
nand U12828 (N_12828,N_11550,N_9891);
nor U12829 (N_12829,N_8258,N_10538);
xnor U12830 (N_12830,N_11090,N_11519);
xnor U12831 (N_12831,N_11571,N_8807);
xnor U12832 (N_12832,N_11172,N_9337);
and U12833 (N_12833,N_8753,N_11538);
or U12834 (N_12834,N_10319,N_11918);
nand U12835 (N_12835,N_11680,N_10981);
and U12836 (N_12836,N_11926,N_11169);
nor U12837 (N_12837,N_10808,N_10144);
or U12838 (N_12838,N_8218,N_10874);
or U12839 (N_12839,N_9228,N_9462);
nand U12840 (N_12840,N_11763,N_9754);
nand U12841 (N_12841,N_9801,N_8383);
nand U12842 (N_12842,N_10219,N_11211);
or U12843 (N_12843,N_10386,N_8926);
nand U12844 (N_12844,N_9766,N_8878);
or U12845 (N_12845,N_8411,N_9237);
or U12846 (N_12846,N_8332,N_11986);
nand U12847 (N_12847,N_10398,N_9771);
and U12848 (N_12848,N_8190,N_10937);
nand U12849 (N_12849,N_9694,N_10478);
or U12850 (N_12850,N_9240,N_11835);
or U12851 (N_12851,N_9335,N_10077);
or U12852 (N_12852,N_8621,N_11702);
nand U12853 (N_12853,N_10110,N_8801);
and U12854 (N_12854,N_8453,N_9215);
nor U12855 (N_12855,N_8018,N_10002);
and U12856 (N_12856,N_11909,N_9178);
nand U12857 (N_12857,N_9439,N_10556);
or U12858 (N_12858,N_8767,N_10203);
nand U12859 (N_12859,N_10071,N_10293);
or U12860 (N_12860,N_11262,N_10910);
nand U12861 (N_12861,N_9886,N_10530);
and U12862 (N_12862,N_8859,N_11859);
nand U12863 (N_12863,N_9532,N_11532);
nand U12864 (N_12864,N_8875,N_9396);
and U12865 (N_12865,N_10078,N_11447);
nand U12866 (N_12866,N_10958,N_9207);
nand U12867 (N_12867,N_8246,N_10856);
or U12868 (N_12868,N_11440,N_9942);
and U12869 (N_12869,N_11552,N_8007);
nor U12870 (N_12870,N_10048,N_11767);
xnor U12871 (N_12871,N_8605,N_10323);
nor U12872 (N_12872,N_9679,N_10882);
and U12873 (N_12873,N_10727,N_8329);
and U12874 (N_12874,N_11368,N_8754);
nand U12875 (N_12875,N_8055,N_9226);
xor U12876 (N_12876,N_9911,N_9575);
nor U12877 (N_12877,N_8048,N_8051);
xnor U12878 (N_12878,N_8953,N_11231);
nand U12879 (N_12879,N_10229,N_9430);
xnor U12880 (N_12880,N_11134,N_10960);
or U12881 (N_12881,N_8267,N_9524);
or U12882 (N_12882,N_10137,N_10394);
nand U12883 (N_12883,N_8998,N_10228);
xor U12884 (N_12884,N_8717,N_10131);
and U12885 (N_12885,N_10512,N_11484);
nand U12886 (N_12886,N_10142,N_9041);
or U12887 (N_12887,N_9747,N_9738);
nand U12888 (N_12888,N_10400,N_9352);
nand U12889 (N_12889,N_10959,N_8814);
nand U12890 (N_12890,N_10584,N_10258);
nand U12891 (N_12891,N_9366,N_10800);
nor U12892 (N_12892,N_11383,N_9934);
nand U12893 (N_12893,N_9974,N_8042);
or U12894 (N_12894,N_9450,N_11061);
and U12895 (N_12895,N_9456,N_10344);
and U12896 (N_12896,N_10744,N_8646);
nor U12897 (N_12897,N_11712,N_8858);
and U12898 (N_12898,N_11441,N_10363);
nor U12899 (N_12899,N_9365,N_8715);
or U12900 (N_12900,N_11829,N_10012);
nand U12901 (N_12901,N_10334,N_11570);
nor U12902 (N_12902,N_10999,N_8512);
nand U12903 (N_12903,N_9796,N_10342);
nor U12904 (N_12904,N_8706,N_11057);
nor U12905 (N_12905,N_10681,N_8275);
or U12906 (N_12906,N_9266,N_10449);
nor U12907 (N_12907,N_9868,N_11954);
and U12908 (N_12908,N_10947,N_11390);
and U12909 (N_12909,N_10244,N_9317);
and U12910 (N_12910,N_10040,N_8691);
and U12911 (N_12911,N_8587,N_8403);
nand U12912 (N_12912,N_8257,N_11198);
nor U12913 (N_12913,N_8446,N_8819);
or U12914 (N_12914,N_8035,N_8067);
nor U12915 (N_12915,N_11042,N_10067);
nor U12916 (N_12916,N_10635,N_10177);
nor U12917 (N_12917,N_8815,N_8277);
and U12918 (N_12918,N_9225,N_8373);
nor U12919 (N_12919,N_9664,N_10583);
nor U12920 (N_12920,N_11277,N_10796);
nand U12921 (N_12921,N_10045,N_11662);
and U12922 (N_12922,N_10001,N_11485);
or U12923 (N_12923,N_10531,N_10931);
nor U12924 (N_12924,N_11110,N_11104);
nand U12925 (N_12925,N_11358,N_11683);
nor U12926 (N_12926,N_11978,N_9260);
or U12927 (N_12927,N_11378,N_8222);
and U12928 (N_12928,N_9858,N_11353);
and U12929 (N_12929,N_10815,N_10903);
nand U12930 (N_12930,N_11886,N_10160);
nor U12931 (N_12931,N_8596,N_10648);
nand U12932 (N_12932,N_9442,N_9597);
and U12933 (N_12933,N_10907,N_9033);
and U12934 (N_12934,N_8138,N_11254);
and U12935 (N_12935,N_8175,N_9417);
nand U12936 (N_12936,N_11704,N_8108);
nor U12937 (N_12937,N_11288,N_9571);
or U12938 (N_12938,N_11583,N_11242);
nand U12939 (N_12939,N_9897,N_10940);
nor U12940 (N_12940,N_8798,N_8742);
and U12941 (N_12941,N_11944,N_9918);
xnor U12942 (N_12942,N_10372,N_9869);
nor U12943 (N_12943,N_10159,N_8565);
or U12944 (N_12944,N_11504,N_11921);
xnor U12945 (N_12945,N_9887,N_8656);
nand U12946 (N_12946,N_8574,N_10753);
or U12947 (N_12947,N_10686,N_9405);
and U12948 (N_12948,N_8355,N_10083);
or U12949 (N_12949,N_10368,N_9502);
or U12950 (N_12950,N_8679,N_9806);
and U12951 (N_12951,N_11453,N_11019);
and U12952 (N_12952,N_9616,N_11142);
and U12953 (N_12953,N_9594,N_11160);
nor U12954 (N_12954,N_11329,N_11003);
or U12955 (N_12955,N_10411,N_9469);
nand U12956 (N_12956,N_8153,N_9779);
or U12957 (N_12957,N_10310,N_11894);
or U12958 (N_12958,N_8489,N_10993);
or U12959 (N_12959,N_11842,N_9216);
nand U12960 (N_12960,N_8466,N_10489);
nor U12961 (N_12961,N_10227,N_9823);
nor U12962 (N_12962,N_10726,N_8330);
or U12963 (N_12963,N_11598,N_10554);
nand U12964 (N_12964,N_9820,N_10854);
and U12965 (N_12965,N_10633,N_10314);
or U12966 (N_12966,N_9954,N_9204);
and U12967 (N_12967,N_8872,N_11234);
or U12968 (N_12968,N_11982,N_8297);
and U12969 (N_12969,N_8015,N_11086);
nor U12970 (N_12970,N_10330,N_9595);
nand U12971 (N_12971,N_10185,N_9229);
nand U12972 (N_12972,N_9537,N_11966);
xnor U12973 (N_12973,N_9729,N_11228);
nand U12974 (N_12974,N_11098,N_8669);
and U12975 (N_12975,N_10718,N_8919);
or U12976 (N_12976,N_9916,N_11155);
and U12977 (N_12977,N_10044,N_11505);
nand U12978 (N_12978,N_8006,N_11686);
and U12979 (N_12979,N_8458,N_8269);
and U12980 (N_12980,N_8119,N_10290);
nand U12981 (N_12981,N_9118,N_10454);
and U12982 (N_12982,N_8402,N_11343);
nor U12983 (N_12983,N_10500,N_11112);
nand U12984 (N_12984,N_11128,N_8079);
and U12985 (N_12985,N_11810,N_8181);
nand U12986 (N_12986,N_8900,N_10704);
or U12987 (N_12987,N_10506,N_10187);
and U12988 (N_12988,N_9946,N_10923);
and U12989 (N_12989,N_10969,N_9617);
and U12990 (N_12990,N_9276,N_10673);
or U12991 (N_12991,N_11488,N_9000);
nand U12992 (N_12992,N_11394,N_10647);
nor U12993 (N_12993,N_8282,N_8639);
nand U12994 (N_12994,N_10158,N_8682);
nand U12995 (N_12995,N_11759,N_10106);
or U12996 (N_12996,N_11500,N_8662);
nand U12997 (N_12997,N_9803,N_10655);
or U12998 (N_12998,N_8909,N_9372);
nor U12999 (N_12999,N_11379,N_8938);
nand U13000 (N_13000,N_11913,N_8414);
or U13001 (N_13001,N_9517,N_8667);
xnor U13002 (N_13002,N_10925,N_8415);
or U13003 (N_13003,N_10899,N_11320);
nand U13004 (N_13004,N_10250,N_11455);
and U13005 (N_13005,N_11060,N_11733);
nand U13006 (N_13006,N_11496,N_10264);
and U13007 (N_13007,N_8227,N_9476);
nand U13008 (N_13008,N_11626,N_10968);
or U13009 (N_13009,N_11514,N_9509);
or U13010 (N_13010,N_8576,N_10406);
nand U13011 (N_13011,N_11685,N_10214);
and U13012 (N_13012,N_11036,N_8563);
nor U13013 (N_13013,N_8531,N_8829);
xnor U13014 (N_13014,N_9968,N_11614);
nor U13015 (N_13015,N_11501,N_8002);
and U13016 (N_13016,N_8320,N_9454);
nand U13017 (N_13017,N_11587,N_10038);
nor U13018 (N_13018,N_9301,N_8920);
nor U13019 (N_13019,N_11937,N_11818);
or U13020 (N_13020,N_8867,N_10841);
and U13021 (N_13021,N_8058,N_9247);
and U13022 (N_13022,N_8225,N_9665);
and U13023 (N_13023,N_9206,N_9306);
or U13024 (N_13024,N_8551,N_8825);
or U13025 (N_13025,N_8876,N_8806);
or U13026 (N_13026,N_10817,N_11435);
nor U13027 (N_13027,N_8918,N_8388);
nor U13028 (N_13028,N_9569,N_10196);
nor U13029 (N_13029,N_11964,N_11907);
nor U13030 (N_13030,N_8519,N_10654);
or U13031 (N_13031,N_8160,N_8802);
xor U13032 (N_13032,N_10626,N_11511);
and U13033 (N_13033,N_10788,N_9243);
nand U13034 (N_13034,N_8743,N_9115);
and U13035 (N_13035,N_9799,N_10036);
nand U13036 (N_13036,N_11867,N_8381);
xor U13037 (N_13037,N_10909,N_9096);
or U13038 (N_13038,N_9094,N_11655);
or U13039 (N_13039,N_8127,N_9782);
and U13040 (N_13040,N_11889,N_11096);
xor U13041 (N_13041,N_11967,N_9865);
and U13042 (N_13042,N_8094,N_9014);
or U13043 (N_13043,N_11883,N_8762);
nor U13044 (N_13044,N_9201,N_10921);
nor U13045 (N_13045,N_9257,N_9520);
or U13046 (N_13046,N_9543,N_9489);
nand U13047 (N_13047,N_8028,N_11697);
nand U13048 (N_13048,N_11227,N_8741);
nand U13049 (N_13049,N_11287,N_9991);
xor U13050 (N_13050,N_11983,N_8740);
nand U13051 (N_13051,N_11261,N_9199);
and U13052 (N_13052,N_10725,N_9596);
and U13053 (N_13053,N_8782,N_10731);
nand U13054 (N_13054,N_8899,N_9488);
or U13055 (N_13055,N_10415,N_11562);
nor U13056 (N_13056,N_10154,N_8333);
or U13057 (N_13057,N_9706,N_9082);
and U13058 (N_13058,N_11791,N_9577);
xor U13059 (N_13059,N_11742,N_8205);
and U13060 (N_13060,N_11634,N_10724);
nand U13061 (N_13061,N_10125,N_10128);
nand U13062 (N_13062,N_9142,N_11515);
and U13063 (N_13063,N_8009,N_11885);
nor U13064 (N_13064,N_10313,N_11843);
nand U13065 (N_13065,N_8693,N_9042);
nand U13066 (N_13066,N_11268,N_9845);
nor U13067 (N_13067,N_8774,N_11963);
nor U13068 (N_13068,N_8059,N_8521);
or U13069 (N_13069,N_10162,N_10135);
nand U13070 (N_13070,N_11935,N_10823);
and U13071 (N_13071,N_9497,N_10773);
nor U13072 (N_13072,N_8547,N_8202);
nor U13073 (N_13073,N_11543,N_11411);
or U13074 (N_13074,N_10632,N_9737);
or U13075 (N_13075,N_11280,N_9549);
and U13076 (N_13076,N_10268,N_10748);
or U13077 (N_13077,N_11730,N_11723);
and U13078 (N_13078,N_9154,N_8148);
and U13079 (N_13079,N_9528,N_9090);
nor U13080 (N_13080,N_9579,N_10875);
nor U13081 (N_13081,N_8147,N_11699);
xnor U13082 (N_13082,N_10973,N_10787);
nor U13083 (N_13083,N_8905,N_8643);
xnor U13084 (N_13084,N_8773,N_11761);
nor U13085 (N_13085,N_9164,N_8308);
or U13086 (N_13086,N_10022,N_10565);
nand U13087 (N_13087,N_8689,N_10750);
and U13088 (N_13088,N_9781,N_9824);
nand U13089 (N_13089,N_10085,N_10009);
and U13090 (N_13090,N_10509,N_8335);
and U13091 (N_13091,N_9293,N_9601);
nor U13092 (N_13092,N_9327,N_11659);
and U13093 (N_13093,N_11946,N_10684);
nand U13094 (N_13094,N_10081,N_11000);
or U13095 (N_13095,N_11990,N_11427);
nor U13096 (N_13096,N_9638,N_9446);
nand U13097 (N_13097,N_8569,N_10124);
and U13098 (N_13098,N_9553,N_8069);
nand U13099 (N_13099,N_11689,N_11077);
and U13100 (N_13100,N_11746,N_9121);
and U13101 (N_13101,N_8787,N_11736);
nand U13102 (N_13102,N_10401,N_10804);
nor U13103 (N_13103,N_9746,N_10977);
and U13104 (N_13104,N_10383,N_8120);
or U13105 (N_13105,N_10479,N_8187);
and U13106 (N_13106,N_9069,N_8075);
or U13107 (N_13107,N_8008,N_10614);
nand U13108 (N_13108,N_9470,N_9367);
and U13109 (N_13109,N_9695,N_8692);
nor U13110 (N_13110,N_8353,N_8455);
xnor U13111 (N_13111,N_8107,N_9745);
and U13112 (N_13112,N_9084,N_10926);
nand U13113 (N_13113,N_10096,N_10280);
nor U13114 (N_13114,N_8440,N_10014);
or U13115 (N_13115,N_11491,N_11653);
nor U13116 (N_13116,N_11101,N_10870);
or U13117 (N_13117,N_10451,N_11941);
and U13118 (N_13118,N_10161,N_8634);
and U13119 (N_13119,N_11197,N_10890);
and U13120 (N_13120,N_10604,N_8230);
nand U13121 (N_13121,N_11573,N_10929);
xnor U13122 (N_13122,N_10221,N_10537);
or U13123 (N_13123,N_11933,N_8635);
nor U13124 (N_13124,N_11063,N_11260);
and U13125 (N_13125,N_11754,N_10220);
and U13126 (N_13126,N_10526,N_9677);
or U13127 (N_13127,N_11755,N_9970);
and U13128 (N_13128,N_10946,N_10115);
and U13129 (N_13129,N_10961,N_8238);
and U13130 (N_13130,N_11354,N_9120);
and U13131 (N_13131,N_9961,N_10407);
nand U13132 (N_13132,N_9038,N_9734);
nand U13133 (N_13133,N_8293,N_10430);
xnor U13134 (N_13134,N_10003,N_9076);
nor U13135 (N_13135,N_10777,N_11089);
xor U13136 (N_13136,N_8545,N_10795);
or U13137 (N_13137,N_9331,N_8617);
and U13138 (N_13138,N_9861,N_9740);
or U13139 (N_13139,N_11876,N_9059);
nor U13140 (N_13140,N_9797,N_10072);
or U13141 (N_13141,N_10649,N_8165);
nand U13142 (N_13142,N_11004,N_9319);
and U13143 (N_13143,N_8524,N_9086);
nand U13144 (N_13144,N_11936,N_10420);
nand U13145 (N_13145,N_8763,N_9344);
xor U13146 (N_13146,N_11052,N_9246);
or U13147 (N_13147,N_8219,N_11276);
and U13148 (N_13148,N_9123,N_9147);
xor U13149 (N_13149,N_10446,N_10945);
nor U13150 (N_13150,N_9825,N_8942);
nand U13151 (N_13151,N_8179,N_10270);
xnor U13152 (N_13152,N_11814,N_11512);
nor U13153 (N_13153,N_8463,N_10210);
nor U13154 (N_13154,N_11195,N_11541);
nor U13155 (N_13155,N_11566,N_11916);
or U13156 (N_13156,N_10361,N_11779);
or U13157 (N_13157,N_11219,N_10470);
xnor U13158 (N_13158,N_11629,N_10289);
and U13159 (N_13159,N_10004,N_8422);
and U13160 (N_13160,N_8089,N_8955);
nand U13161 (N_13161,N_8886,N_8477);
xor U13162 (N_13162,N_10475,N_11878);
nor U13163 (N_13163,N_11478,N_9909);
or U13164 (N_13164,N_10273,N_10213);
and U13165 (N_13165,N_9011,N_11627);
nand U13166 (N_13166,N_8542,N_11347);
and U13167 (N_13167,N_11564,N_9731);
xor U13168 (N_13168,N_9308,N_9841);
and U13169 (N_13169,N_11582,N_10194);
nor U13170 (N_13170,N_10569,N_9150);
nor U13171 (N_13171,N_11855,N_10062);
or U13172 (N_13172,N_8104,N_9650);
or U13173 (N_13173,N_10234,N_10593);
nand U13174 (N_13174,N_8005,N_8637);
nor U13175 (N_13175,N_8722,N_11034);
xor U13176 (N_13176,N_10941,N_11129);
or U13177 (N_13177,N_8980,N_10021);
and U13178 (N_13178,N_9362,N_11597);
and U13179 (N_13179,N_9687,N_9545);
or U13180 (N_13180,N_10643,N_9535);
xor U13181 (N_13181,N_10201,N_8861);
xor U13182 (N_13182,N_8393,N_10752);
and U13183 (N_13183,N_10906,N_8929);
or U13184 (N_13184,N_8632,N_9328);
or U13185 (N_13185,N_10175,N_11798);
nor U13186 (N_13186,N_8705,N_9661);
or U13187 (N_13187,N_10801,N_8620);
or U13188 (N_13188,N_11716,N_8680);
nor U13189 (N_13189,N_11972,N_10439);
nand U13190 (N_13190,N_9906,N_10328);
or U13191 (N_13191,N_9859,N_9457);
nor U13192 (N_13192,N_9210,N_9764);
nor U13193 (N_13193,N_11130,N_8965);
nand U13194 (N_13194,N_8475,N_10965);
and U13195 (N_13195,N_10332,N_11210);
or U13196 (N_13196,N_8286,N_9668);
and U13197 (N_13197,N_9404,N_9117);
nand U13198 (N_13198,N_9642,N_9863);
nand U13199 (N_13199,N_10579,N_11769);
and U13200 (N_13200,N_11251,N_11844);
and U13201 (N_13201,N_11467,N_9124);
or U13202 (N_13202,N_9022,N_9356);
nor U13203 (N_13203,N_8665,N_10862);
nand U13204 (N_13204,N_8478,N_10677);
nor U13205 (N_13205,N_9015,N_11804);
xnor U13206 (N_13206,N_8940,N_8885);
and U13207 (N_13207,N_11892,N_10111);
or U13208 (N_13208,N_10516,N_8606);
and U13209 (N_13209,N_11189,N_11283);
nand U13210 (N_13210,N_9722,N_8027);
xor U13211 (N_13211,N_11603,N_10138);
xnor U13212 (N_13212,N_9127,N_10697);
and U13213 (N_13213,N_11144,N_8457);
nor U13214 (N_13214,N_8800,N_10043);
or U13215 (N_13215,N_9713,N_11840);
nor U13216 (N_13216,N_8873,N_9880);
nor U13217 (N_13217,N_11557,N_11549);
nand U13218 (N_13218,N_10646,N_11932);
and U13219 (N_13219,N_11958,N_9508);
nand U13220 (N_13220,N_9749,N_9324);
nand U13221 (N_13221,N_9838,N_10939);
xnor U13222 (N_13222,N_8309,N_11167);
and U13223 (N_13223,N_10963,N_8880);
nand U13224 (N_13224,N_10205,N_9641);
nand U13225 (N_13225,N_9944,N_10254);
nor U13226 (N_13226,N_9057,N_9049);
xor U13227 (N_13227,N_10978,N_8830);
and U13228 (N_13228,N_11107,N_10476);
nor U13229 (N_13229,N_8838,N_9340);
nor U13230 (N_13230,N_10668,N_8441);
nor U13231 (N_13231,N_9058,N_8649);
nand U13232 (N_13232,N_8180,N_10252);
nand U13233 (N_13233,N_9890,N_11406);
nand U13234 (N_13234,N_11192,N_8994);
and U13235 (N_13235,N_8795,N_9233);
nand U13236 (N_13236,N_8822,N_10495);
and U13237 (N_13237,N_8912,N_8272);
or U13238 (N_13238,N_10066,N_10181);
nand U13239 (N_13239,N_10018,N_9447);
or U13240 (N_13240,N_8502,N_8664);
xor U13241 (N_13241,N_10916,N_8421);
nor U13242 (N_13242,N_9453,N_10667);
and U13243 (N_13243,N_9111,N_9166);
and U13244 (N_13244,N_9336,N_8750);
nand U13245 (N_13245,N_8361,N_10399);
nor U13246 (N_13246,N_9531,N_11540);
xnor U13247 (N_13247,N_11539,N_8247);
nand U13248 (N_13248,N_11022,N_11424);
nor U13249 (N_13249,N_8378,N_11429);
and U13250 (N_13250,N_11811,N_11635);
xnor U13251 (N_13251,N_11956,N_10404);
nand U13252 (N_13252,N_9318,N_10896);
nor U13253 (N_13253,N_9691,N_9385);
nand U13254 (N_13254,N_10778,N_9866);
nor U13255 (N_13255,N_9807,N_11468);
and U13256 (N_13256,N_8034,N_8736);
nor U13257 (N_13257,N_8827,N_9438);
and U13258 (N_13258,N_10622,N_9177);
nand U13259 (N_13259,N_8493,N_11865);
and U13260 (N_13260,N_11607,N_9176);
and U13261 (N_13261,N_10850,N_8066);
xnor U13262 (N_13262,N_9354,N_9830);
and U13263 (N_13263,N_10224,N_10741);
or U13264 (N_13264,N_9155,N_9065);
or U13265 (N_13265,N_11875,N_10141);
and U13266 (N_13266,N_9977,N_9023);
or U13267 (N_13267,N_8084,N_8173);
nor U13268 (N_13268,N_8959,N_11437);
and U13269 (N_13269,N_10983,N_11187);
nand U13270 (N_13270,N_11398,N_11135);
and U13271 (N_13271,N_9652,N_10320);
or U13272 (N_13272,N_10703,N_8322);
nand U13273 (N_13273,N_11792,N_11499);
or U13274 (N_13274,N_11015,N_9236);
xor U13275 (N_13275,N_11503,N_9792);
and U13276 (N_13276,N_10501,N_8974);
xnor U13277 (N_13277,N_9190,N_10990);
nand U13278 (N_13278,N_11868,N_9790);
nor U13279 (N_13279,N_9698,N_11902);
and U13280 (N_13280,N_9628,N_11106);
or U13281 (N_13281,N_11489,N_11355);
nand U13282 (N_13282,N_9294,N_11528);
nor U13283 (N_13283,N_8261,N_10730);
nand U13284 (N_13284,N_8232,N_10291);
and U13285 (N_13285,N_11898,N_11660);
nand U13286 (N_13286,N_9184,N_11221);
nor U13287 (N_13287,N_10623,N_8264);
nor U13288 (N_13288,N_9705,N_8100);
xnor U13289 (N_13289,N_8243,N_11663);
nand U13290 (N_13290,N_11224,N_10069);
and U13291 (N_13291,N_10357,N_10845);
nand U13292 (N_13292,N_8199,N_11951);
xor U13293 (N_13293,N_11793,N_10690);
nand U13294 (N_13294,N_9075,N_9460);
nand U13295 (N_13295,N_11641,N_8961);
nor U13296 (N_13296,N_11590,N_10887);
or U13297 (N_13297,N_9505,N_10833);
nor U13298 (N_13298,N_9045,N_8690);
and U13299 (N_13299,N_8010,N_11940);
or U13300 (N_13300,N_10550,N_10114);
or U13301 (N_13301,N_11866,N_8660);
and U13302 (N_13302,N_9326,N_8571);
nor U13303 (N_13303,N_11465,N_10322);
nand U13304 (N_13304,N_11910,N_8506);
nand U13305 (N_13305,N_9669,N_10511);
nand U13306 (N_13306,N_11345,N_8840);
nor U13307 (N_13307,N_9451,N_10640);
xnor U13308 (N_13308,N_11407,N_9590);
xor U13309 (N_13309,N_8137,N_8989);
nor U13310 (N_13310,N_9032,N_9010);
nand U13311 (N_13311,N_10628,N_11507);
nand U13312 (N_13312,N_10611,N_10719);
nand U13313 (N_13313,N_10798,N_8641);
or U13314 (N_13314,N_10905,N_9922);
and U13315 (N_13315,N_11998,N_11209);
and U13316 (N_13316,N_9658,N_10109);
and U13317 (N_13317,N_8817,N_10857);
nor U13318 (N_13318,N_11509,N_10967);
nor U13319 (N_13319,N_10519,N_8350);
nor U13320 (N_13320,N_10539,N_9786);
nor U13321 (N_13321,N_11903,N_8467);
and U13322 (N_13322,N_10793,N_10257);
nor U13323 (N_13323,N_10794,N_8080);
or U13324 (N_13324,N_10737,N_8451);
nand U13325 (N_13325,N_10433,N_10607);
or U13326 (N_13326,N_9812,N_9744);
or U13327 (N_13327,N_10341,N_10387);
and U13328 (N_13328,N_11649,N_11431);
nand U13329 (N_13329,N_8325,N_10169);
or U13330 (N_13330,N_8694,N_9670);
nand U13331 (N_13331,N_11326,N_10265);
nor U13332 (N_13332,N_11236,N_10616);
nand U13333 (N_13333,N_10459,N_9230);
nand U13334 (N_13334,N_8476,N_8314);
nand U13335 (N_13335,N_10256,N_9876);
xor U13336 (N_13336,N_10306,N_8845);
and U13337 (N_13337,N_8208,N_9937);
xnor U13338 (N_13338,N_10352,N_8491);
nor U13339 (N_13339,N_11989,N_10659);
and U13340 (N_13340,N_11669,N_9742);
or U13341 (N_13341,N_8352,N_10723);
nor U13342 (N_13342,N_10997,N_10140);
or U13343 (N_13343,N_9289,N_10104);
or U13344 (N_13344,N_11637,N_9917);
nor U13345 (N_13345,N_11392,N_9685);
and U13346 (N_13346,N_8564,N_9116);
xnor U13347 (N_13347,N_10606,N_10595);
and U13348 (N_13348,N_11031,N_10784);
and U13349 (N_13349,N_9915,N_9321);
nor U13350 (N_13350,N_10484,N_11508);
and U13351 (N_13351,N_11806,N_11924);
nand U13352 (N_13352,N_10182,N_10785);
and U13353 (N_13353,N_8188,N_9390);
nand U13354 (N_13354,N_10349,N_9274);
nand U13355 (N_13355,N_9836,N_10535);
nand U13356 (N_13356,N_10742,N_11596);
nand U13357 (N_13357,N_11318,N_10532);
and U13358 (N_13358,N_10103,N_8387);
nand U13359 (N_13359,N_11006,N_8973);
nor U13360 (N_13360,N_9418,N_10029);
nor U13361 (N_13361,N_11630,N_11745);
or U13362 (N_13362,N_10456,N_11845);
nor U13363 (N_13363,N_9114,N_10445);
and U13364 (N_13364,N_8790,N_11099);
nor U13365 (N_13365,N_10212,N_9856);
or U13366 (N_13366,N_8553,N_11145);
nor U13367 (N_13367,N_10803,N_10351);
xor U13368 (N_13368,N_9183,N_10153);
and U13369 (N_13369,N_10236,N_9710);
and U13370 (N_13370,N_10288,N_10455);
or U13371 (N_13371,N_11146,N_8976);
xnor U13372 (N_13372,N_8364,N_10523);
nand U13373 (N_13373,N_9119,N_8794);
nand U13374 (N_13374,N_8933,N_9403);
and U13375 (N_13375,N_11426,N_11149);
and U13376 (N_13376,N_9513,N_9951);
or U13377 (N_13377,N_10721,N_9070);
nand U13378 (N_13378,N_8470,N_10891);
or U13379 (N_13379,N_9271,N_9112);
or U13380 (N_13380,N_9624,N_8113);
nor U13381 (N_13381,N_9654,N_10260);
nand U13382 (N_13382,N_11920,N_10152);
or U13383 (N_13383,N_9234,N_10170);
nor U13384 (N_13384,N_8511,N_11863);
nor U13385 (N_13385,N_8673,N_9898);
nand U13386 (N_13386,N_11124,N_8252);
nor U13387 (N_13387,N_10568,N_9721);
or U13388 (N_13388,N_11274,N_9031);
and U13389 (N_13389,N_8460,N_9399);
xor U13390 (N_13390,N_10566,N_9068);
or U13391 (N_13391,N_11013,N_10866);
nor U13392 (N_13392,N_9030,N_11735);
nor U13393 (N_13393,N_11553,N_11917);
xnor U13394 (N_13394,N_10316,N_9209);
xnor U13395 (N_13395,N_8469,N_11988);
or U13396 (N_13396,N_11643,N_8766);
or U13397 (N_13397,N_8287,N_10546);
nor U13398 (N_13398,N_10355,N_10481);
or U13399 (N_13399,N_8310,N_9161);
xnor U13400 (N_13400,N_8595,N_10543);
nor U13401 (N_13401,N_8670,N_11604);
or U13402 (N_13402,N_11650,N_10255);
and U13403 (N_13403,N_11191,N_11417);
or U13404 (N_13404,N_9148,N_8568);
and U13405 (N_13405,N_8887,N_9189);
nand U13406 (N_13406,N_9686,N_9621);
and U13407 (N_13407,N_11938,N_10095);
nand U13408 (N_13408,N_11001,N_8416);
or U13409 (N_13409,N_8167,N_9636);
nand U13410 (N_13410,N_9485,N_10824);
or U13411 (N_13411,N_8915,N_8657);
nor U13412 (N_13412,N_9693,N_8626);
nor U13413 (N_13413,N_11132,N_9428);
and U13414 (N_13414,N_9988,N_10356);
nand U13415 (N_13415,N_8533,N_11997);
nand U13416 (N_13416,N_10325,N_8095);
or U13417 (N_13417,N_10425,N_9659);
or U13418 (N_13418,N_8609,N_9604);
or U13419 (N_13419,N_11482,N_9618);
and U13420 (N_13420,N_8943,N_9165);
or U13421 (N_13421,N_11652,N_8543);
nand U13422 (N_13422,N_10786,N_9063);
nor U13423 (N_13423,N_10031,N_9153);
or U13424 (N_13424,N_8291,N_11740);
xnor U13425 (N_13425,N_9018,N_10572);
and U13426 (N_13426,N_8430,N_8280);
nand U13427 (N_13427,N_9345,N_11813);
nand U13428 (N_13428,N_9424,N_9882);
or U13429 (N_13429,N_8321,N_10709);
nand U13430 (N_13430,N_9263,N_11531);
nand U13431 (N_13431,N_8273,N_9195);
and U13432 (N_13432,N_9217,N_9261);
and U13433 (N_13433,N_9265,N_10494);
nor U13434 (N_13434,N_11214,N_8311);
nand U13435 (N_13435,N_11589,N_8109);
and U13436 (N_13436,N_8070,N_8833);
nand U13437 (N_13437,N_8883,N_8283);
and U13438 (N_13438,N_11568,N_11708);
nor U13439 (N_13439,N_11830,N_9653);
or U13440 (N_13440,N_11470,N_9287);
or U13441 (N_13441,N_8612,N_10895);
or U13442 (N_13442,N_9295,N_8841);
nand U13443 (N_13443,N_10989,N_10664);
nand U13444 (N_13444,N_9478,N_8017);
and U13445 (N_13445,N_9953,N_10739);
nand U13446 (N_13446,N_11232,N_11327);
nor U13447 (N_13447,N_8445,N_11756);
and U13448 (N_13448,N_11177,N_9392);
or U13449 (N_13449,N_8231,N_9928);
or U13450 (N_13450,N_11410,N_10427);
xor U13451 (N_13451,N_8739,N_9733);
nor U13452 (N_13452,N_8174,N_8849);
xor U13453 (N_13453,N_9109,N_10740);
or U13454 (N_13454,N_9034,N_11749);
or U13455 (N_13455,N_10371,N_11021);
and U13456 (N_13456,N_11137,N_9332);
nand U13457 (N_13457,N_11995,N_8450);
nor U13458 (N_13458,N_8392,N_9144);
and U13459 (N_13459,N_10011,N_10338);
or U13460 (N_13460,N_10797,N_8341);
or U13461 (N_13461,N_11823,N_11258);
or U13462 (N_13462,N_11141,N_11578);
or U13463 (N_13463,N_8295,N_10751);
nand U13464 (N_13464,N_10859,N_8226);
and U13465 (N_13465,N_11962,N_9159);
nor U13466 (N_13466,N_10600,N_11665);
nor U13467 (N_13467,N_10460,N_11314);
xor U13468 (N_13468,N_9278,N_10994);
or U13469 (N_13469,N_8821,N_8093);
or U13470 (N_13470,N_11201,N_10780);
and U13471 (N_13471,N_11168,N_9374);
or U13472 (N_13472,N_8063,N_8386);
nand U13473 (N_13473,N_10375,N_11206);
or U13474 (N_13474,N_8957,N_11473);
and U13475 (N_13475,N_8126,N_11312);
and U13476 (N_13476,N_11361,N_10987);
nor U13477 (N_13477,N_8001,N_8701);
and U13478 (N_13478,N_8327,N_8419);
or U13479 (N_13479,N_9933,N_10097);
xnor U13480 (N_13480,N_8614,N_8890);
nor U13481 (N_13481,N_10561,N_8854);
or U13482 (N_13482,N_9715,N_8823);
nand U13483 (N_13483,N_10953,N_10117);
nor U13484 (N_13484,N_11785,N_11608);
nor U13485 (N_13485,N_10235,N_9079);
nor U13486 (N_13486,N_10061,N_11165);
nand U13487 (N_13487,N_11322,N_8480);
xnor U13488 (N_13488,N_11714,N_11292);
xor U13489 (N_13489,N_9143,N_8791);
or U13490 (N_13490,N_9984,N_11494);
and U13491 (N_13491,N_11559,N_11673);
xnor U13492 (N_13492,N_11350,N_10174);
and U13493 (N_13493,N_10226,N_11943);
or U13494 (N_13494,N_9982,N_10179);
or U13495 (N_13495,N_11516,N_11180);
nor U13496 (N_13496,N_9474,N_9712);
nor U13497 (N_13497,N_9973,N_9950);
nand U13498 (N_13498,N_8560,N_8161);
nor U13499 (N_13499,N_8076,N_9883);
nand U13500 (N_13500,N_11797,N_11957);
nand U13501 (N_13501,N_8507,N_10942);
nor U13502 (N_13502,N_11460,N_10612);
and U13503 (N_13503,N_11584,N_10353);
nand U13504 (N_13504,N_8975,N_11421);
xor U13505 (N_13505,N_11625,N_11196);
xnor U13506 (N_13506,N_10468,N_11269);
nor U13507 (N_13507,N_9262,N_10007);
or U13508 (N_13508,N_8064,N_11405);
or U13509 (N_13509,N_11386,N_8583);
and U13510 (N_13510,N_11698,N_8842);
nor U13511 (N_13511,N_8843,N_9067);
nand U13512 (N_13512,N_9021,N_11955);
or U13513 (N_13513,N_11760,N_11284);
and U13514 (N_13514,N_8260,N_9834);
or U13515 (N_13515,N_8907,N_8532);
or U13516 (N_13516,N_9443,N_8597);
or U13517 (N_13517,N_10893,N_9391);
nand U13518 (N_13518,N_8724,N_11914);
xnor U13519 (N_13519,N_10974,N_8889);
nor U13520 (N_13520,N_8550,N_11461);
nand U13521 (N_13521,N_8659,N_8032);
xnor U13522 (N_13522,N_8505,N_11293);
xnor U13523 (N_13523,N_10347,N_8607);
and U13524 (N_13524,N_9475,N_8083);
nor U13525 (N_13525,N_9683,N_9814);
xnor U13526 (N_13526,N_8068,N_11389);
nand U13527 (N_13527,N_11666,N_11796);
or U13528 (N_13528,N_8382,N_11497);
and U13529 (N_13529,N_8906,N_11323);
nand U13530 (N_13530,N_8630,N_9645);
nor U13531 (N_13531,N_8499,N_10892);
nor U13532 (N_13532,N_9584,N_8072);
and U13533 (N_13533,N_9561,N_8056);
nor U13534 (N_13534,N_9957,N_11517);
or U13535 (N_13535,N_9350,N_9349);
nor U13536 (N_13536,N_8465,N_9568);
nor U13537 (N_13537,N_9480,N_11961);
nor U13538 (N_13538,N_8855,N_9903);
nor U13539 (N_13539,N_8449,N_9848);
nand U13540 (N_13540,N_9013,N_9994);
xnor U13541 (N_13541,N_10954,N_10269);
nand U13542 (N_13542,N_8954,N_9490);
nand U13543 (N_13543,N_10790,N_8115);
or U13544 (N_13544,N_9091,N_10915);
nand U13545 (N_13545,N_9052,N_10218);
nand U13546 (N_13546,N_10277,N_9351);
nor U13547 (N_13547,N_10047,N_8186);
nand U13548 (N_13548,N_8526,N_10775);
xnor U13549 (N_13549,N_10548,N_11247);
xnor U13550 (N_13550,N_11334,N_10779);
nand U13551 (N_13551,N_11480,N_9857);
or U13552 (N_13552,N_9455,N_10687);
or U13553 (N_13553,N_11654,N_11199);
xor U13554 (N_13554,N_9491,N_10878);
nor U13555 (N_13555,N_8963,N_11182);
and U13556 (N_13556,N_8503,N_9140);
or U13557 (N_13557,N_8128,N_9452);
nor U13558 (N_13558,N_8504,N_11208);
nand U13559 (N_13559,N_11523,N_11256);
or U13560 (N_13560,N_9846,N_10146);
xor U13561 (N_13561,N_10567,N_9312);
and U13562 (N_13562,N_10972,N_11348);
nand U13563 (N_13563,N_9239,N_11139);
and U13564 (N_13564,N_11449,N_9708);
and U13565 (N_13565,N_11706,N_8434);
and U13566 (N_13566,N_11007,N_9904);
xor U13567 (N_13567,N_10496,N_8029);
and U13568 (N_13568,N_8700,N_8744);
nand U13569 (N_13569,N_8555,N_10178);
or U13570 (N_13570,N_11638,N_11032);
xnor U13571 (N_13571,N_8300,N_9040);
nand U13572 (N_13572,N_8319,N_8413);
nand U13573 (N_13573,N_10525,N_11393);
nor U13574 (N_13574,N_8749,N_11113);
nor U13575 (N_13575,N_10933,N_11931);
nand U13576 (N_13576,N_9789,N_9704);
or U13577 (N_13577,N_8675,N_8877);
and U13578 (N_13578,N_10781,N_8145);
nor U13579 (N_13579,N_10544,N_8541);
or U13580 (N_13580,N_9373,N_8241);
xor U13581 (N_13581,N_10283,N_8768);
nand U13582 (N_13582,N_11750,N_8988);
and U13583 (N_13583,N_11335,N_8951);
and U13584 (N_13584,N_8483,N_8296);
xor U13585 (N_13585,N_11220,N_11120);
or U13586 (N_13586,N_11657,N_8748);
nor U13587 (N_13587,N_10145,N_10515);
xnor U13588 (N_13588,N_8778,N_8831);
nor U13589 (N_13589,N_11123,N_10666);
or U13590 (N_13590,N_11108,N_10215);
or U13591 (N_13591,N_10068,N_11561);
or U13592 (N_13592,N_10091,N_8559);
and U13593 (N_13593,N_8274,N_10120);
xnor U13594 (N_13594,N_11727,N_9125);
nand U13595 (N_13595,N_10392,N_9436);
and U13596 (N_13596,N_10463,N_10452);
nand U13597 (N_13597,N_11422,N_11344);
nand U13598 (N_13598,N_10508,N_11965);
and U13599 (N_13599,N_8535,N_10631);
or U13600 (N_13600,N_8610,N_8200);
nor U13601 (N_13601,N_8685,N_10838);
nand U13602 (N_13602,N_8092,N_9702);
nand U13603 (N_13603,N_11530,N_11307);
xnor U13604 (N_13604,N_10246,N_10547);
nand U13605 (N_13605,N_8432,N_10274);
nand U13606 (N_13606,N_8746,N_9370);
or U13607 (N_13607,N_9839,N_11896);
nor U13608 (N_13608,N_8210,N_9981);
and U13609 (N_13609,N_10764,N_8030);
and U13610 (N_13610,N_8789,N_9378);
nand U13611 (N_13611,N_8852,N_8602);
nor U13612 (N_13612,N_11190,N_9401);
or U13613 (N_13613,N_8683,N_9975);
nand U13614 (N_13614,N_11976,N_10847);
and U13615 (N_13615,N_11905,N_10551);
nand U13616 (N_13616,N_11243,N_8110);
nor U13617 (N_13617,N_10837,N_10017);
and U13618 (N_13618,N_10816,N_8255);
nand U13619 (N_13619,N_11067,N_10825);
nand U13620 (N_13620,N_8294,N_11237);
and U13621 (N_13621,N_8589,N_11821);
and U13622 (N_13622,N_9565,N_10156);
or U13623 (N_13623,N_8913,N_8019);
xor U13624 (N_13624,N_11973,N_10443);
nor U13625 (N_13625,N_10843,N_8759);
nor U13626 (N_13626,N_11849,N_10964);
or U13627 (N_13627,N_9892,N_8820);
nand U13628 (N_13628,N_11719,N_8528);
or U13629 (N_13629,N_8585,N_8910);
and U13630 (N_13630,N_8677,N_9877);
nor U13631 (N_13631,N_8666,N_9631);
and U13632 (N_13632,N_11820,N_10904);
and U13633 (N_13633,N_8196,N_9445);
and U13634 (N_13634,N_10098,N_9339);
nand U13635 (N_13635,N_10312,N_10588);
and U13636 (N_13636,N_11402,N_11058);
or U13637 (N_13637,N_11054,N_8418);
nand U13638 (N_13638,N_8608,N_10015);
nand U13639 (N_13639,N_9269,N_11122);
xnor U13640 (N_13640,N_11832,N_11874);
or U13641 (N_13641,N_10064,N_11862);
nor U13642 (N_13642,N_8118,N_11646);
nand U13643 (N_13643,N_9029,N_11367);
nand U13644 (N_13644,N_11330,N_11904);
and U13645 (N_13645,N_9054,N_10717);
nand U13646 (N_13646,N_10873,N_9614);
nor U13647 (N_13647,N_9427,N_10393);
nor U13648 (N_13648,N_10689,N_8135);
and U13649 (N_13649,N_11786,N_10183);
nor U13650 (N_13650,N_8803,N_10601);
and U13651 (N_13651,N_11555,N_8707);
nor U13652 (N_13652,N_9187,N_11645);
nand U13653 (N_13653,N_8401,N_9557);
nand U13654 (N_13654,N_8752,N_9062);
and U13655 (N_13655,N_10193,N_11466);
or U13656 (N_13656,N_10367,N_9703);
nor U13657 (N_13657,N_9333,N_9078);
nor U13658 (N_13658,N_11415,N_11728);
and U13659 (N_13659,N_10418,N_9835);
nor U13660 (N_13660,N_11436,N_10602);
nand U13661 (N_13661,N_9599,N_9073);
and U13662 (N_13662,N_8472,N_11278);
nor U13663 (N_13663,N_9602,N_8197);
xor U13664 (N_13664,N_11822,N_8931);
nor U13665 (N_13665,N_11399,N_9972);
and U13666 (N_13666,N_8932,N_11311);
and U13667 (N_13667,N_11678,N_9932);
or U13668 (N_13668,N_10809,N_10674);
nand U13669 (N_13669,N_9644,N_11851);
nor U13670 (N_13670,N_8891,N_11612);
nor U13671 (N_13671,N_8824,N_9298);
or U13672 (N_13672,N_11934,N_8158);
nor U13673 (N_13673,N_9758,N_11974);
xor U13674 (N_13674,N_10307,N_10202);
nand U13675 (N_13675,N_8796,N_8154);
nand U13676 (N_13676,N_9714,N_8233);
nand U13677 (N_13677,N_11848,N_9817);
or U13678 (N_13678,N_8087,N_11072);
or U13679 (N_13679,N_11282,N_10521);
and U13680 (N_13680,N_11802,N_8176);
xnor U13681 (N_13681,N_8301,N_10807);
or U13682 (N_13682,N_9966,N_11328);
or U13683 (N_13683,N_11068,N_9607);
xnor U13684 (N_13684,N_9461,N_11677);
nor U13685 (N_13685,N_9815,N_9680);
and U13686 (N_13686,N_10005,N_8428);
and U13687 (N_13687,N_11518,N_8420);
nand U13688 (N_13688,N_11238,N_8171);
or U13689 (N_13689,N_8945,N_8719);
nor U13690 (N_13690,N_10329,N_11062);
nand U13691 (N_13691,N_10422,N_8101);
xnor U13692 (N_13692,N_9927,N_9784);
nor U13693 (N_13693,N_10988,N_9995);
or U13694 (N_13694,N_11409,N_11789);
and U13695 (N_13695,N_9168,N_9864);
or U13696 (N_13696,N_9145,N_8292);
nor U13697 (N_13697,N_8644,N_10262);
or U13698 (N_13698,N_8464,N_11126);
nor U13699 (N_13699,N_9222,N_10914);
nand U13700 (N_13700,N_10528,N_8448);
nand U13701 (N_13701,N_11092,N_8366);
and U13702 (N_13702,N_8733,N_8987);
and U13703 (N_13703,N_11527,N_11215);
nor U13704 (N_13704,N_11163,N_9674);
and U13705 (N_13705,N_11984,N_9773);
and U13706 (N_13706,N_8004,N_8584);
nor U13707 (N_13707,N_9389,N_10317);
nor U13708 (N_13708,N_11893,N_9131);
or U13709 (N_13709,N_10950,N_8346);
nor U13710 (N_13710,N_9560,N_9574);
or U13711 (N_13711,N_8116,N_8281);
nor U13712 (N_13712,N_8575,N_9967);
or U13713 (N_13713,N_9530,N_10472);
nor U13714 (N_13714,N_9435,N_8937);
nor U13715 (N_13715,N_11430,N_11908);
and U13716 (N_13716,N_8254,N_11131);
or U13717 (N_13717,N_11551,N_11184);
and U13718 (N_13718,N_10834,N_10685);
nor U13719 (N_13719,N_8139,N_11397);
and U13720 (N_13720,N_10952,N_9931);
or U13721 (N_13721,N_10820,N_8756);
nor U13722 (N_13722,N_8044,N_9281);
nand U13723 (N_13723,N_10863,N_8141);
or U13724 (N_13724,N_11741,N_11075);
nand U13725 (N_13725,N_10598,N_10093);
and U13726 (N_13726,N_11103,N_10922);
or U13727 (N_13727,N_8710,N_10928);
or U13728 (N_13728,N_8136,N_8057);
and U13729 (N_13729,N_8351,N_9197);
nand U13730 (N_13730,N_9699,N_11012);
or U13731 (N_13731,N_9149,N_11871);
or U13732 (N_13732,N_11856,N_8074);
or U13733 (N_13733,N_11668,N_8808);
or U13734 (N_13734,N_8893,N_8417);
nand U13735 (N_13735,N_9965,N_11884);
nand U13736 (N_13736,N_9279,N_11788);
nor U13737 (N_13737,N_10700,N_11632);
nand U13738 (N_13738,N_8482,N_10105);
and U13739 (N_13739,N_11586,N_9828);
and U13740 (N_13740,N_8696,N_11906);
and U13741 (N_13741,N_9609,N_11248);
xnor U13742 (N_13742,N_9377,N_11078);
nand U13743 (N_13743,N_8561,N_9050);
or U13744 (N_13744,N_8224,N_11207);
nor U13745 (N_13745,N_10898,N_10362);
and U13746 (N_13746,N_10979,N_9368);
and U13747 (N_13747,N_10133,N_11833);
nor U13748 (N_13748,N_11325,N_9753);
nand U13749 (N_13749,N_11805,N_8251);
nand U13750 (N_13750,N_9227,N_9423);
nor U13751 (N_13751,N_9843,N_10708);
or U13752 (N_13752,N_9141,N_10498);
nor U13753 (N_13753,N_10294,N_9100);
nor U13754 (N_13754,N_10275,N_8217);
nor U13755 (N_13755,N_9411,N_8687);
nor U13756 (N_13756,N_9788,N_10195);
or U13757 (N_13757,N_9329,N_8404);
or U13758 (N_13758,N_10410,N_8235);
nand U13759 (N_13759,N_11079,N_9682);
nand U13760 (N_13760,N_10051,N_8588);
nor U13761 (N_13761,N_11125,N_11710);
nor U13762 (N_13762,N_9448,N_11416);
nand U13763 (N_13763,N_8529,N_9778);
nand U13764 (N_13764,N_11837,N_8672);
and U13765 (N_13765,N_9945,N_11452);
and U13766 (N_13766,N_8979,N_10504);
nor U13767 (N_13767,N_10350,N_11186);
nand U13768 (N_13768,N_8271,N_9723);
nor U13769 (N_13769,N_10639,N_8727);
and U13770 (N_13770,N_8628,N_11994);
or U13771 (N_13771,N_11558,N_9122);
or U13772 (N_13772,N_9315,N_8946);
nor U13773 (N_13773,N_10951,N_11094);
nor U13774 (N_13774,N_9393,N_11469);
nor U13775 (N_13775,N_10991,N_9572);
nand U13776 (N_13776,N_10783,N_8111);
nor U13777 (N_13777,N_10680,N_9613);
nand U13778 (N_13778,N_11879,N_8755);
and U13779 (N_13779,N_11056,N_9952);
and U13780 (N_13780,N_8544,N_8713);
and U13781 (N_13781,N_9097,N_10699);
nor U13782 (N_13782,N_9516,N_10247);
nor U13783 (N_13783,N_9534,N_9627);
and U13784 (N_13784,N_9622,N_10924);
nor U13785 (N_13785,N_11462,N_8517);
nand U13786 (N_13786,N_9138,N_8299);
and U13787 (N_13787,N_9309,N_8263);
or U13788 (N_13788,N_9610,N_9522);
and U13789 (N_13789,N_10605,N_11331);
or U13790 (N_13790,N_11812,N_8315);
nand U13791 (N_13791,N_10766,N_10412);
and U13792 (N_13792,N_11510,N_11869);
and U13793 (N_13793,N_11521,N_10702);
nand U13794 (N_13794,N_8307,N_9810);
nand U13795 (N_13795,N_9697,N_8721);
and U13796 (N_13796,N_8835,N_10240);
nand U13797 (N_13797,N_8558,N_11611);
nand U13798 (N_13798,N_9284,N_9113);
and U13799 (N_13799,N_9656,N_11560);
or U13800 (N_13800,N_9440,N_9582);
and U13801 (N_13801,N_9847,N_11529);
or U13802 (N_13802,N_10248,N_8265);
xor U13803 (N_13803,N_8732,N_9692);
and U13804 (N_13804,N_8288,N_8653);
nand U13805 (N_13805,N_8860,N_10682);
nand U13806 (N_13806,N_11581,N_8546);
and U13807 (N_13807,N_8023,N_9587);
or U13808 (N_13808,N_8810,N_8443);
and U13809 (N_13809,N_8688,N_11049);
nand U13810 (N_13810,N_9231,N_8785);
xnor U13811 (N_13811,N_9541,N_9186);
nor U13812 (N_13812,N_8925,N_8930);
and U13813 (N_13813,N_10894,N_10230);
nand U13814 (N_13814,N_8928,N_8903);
or U13815 (N_13815,N_11140,N_9093);
nand U13816 (N_13816,N_9724,N_8498);
or U13817 (N_13817,N_10920,N_9302);
and U13818 (N_13818,N_9380,N_11018);
nor U13819 (N_13819,N_8654,N_11765);
or U13820 (N_13820,N_8799,N_9055);
nor U13821 (N_13821,N_9536,N_10811);
nor U13822 (N_13822,N_9919,N_9325);
or U13823 (N_13823,N_10388,N_11309);
or U13824 (N_13824,N_8442,N_9137);
or U13825 (N_13825,N_11891,N_8423);
nor U13826 (N_13826,N_9212,N_8757);
xor U13827 (N_13827,N_10243,N_10671);
nor U13828 (N_13828,N_8106,N_8077);
nor U13829 (N_13829,N_11339,N_8431);
nor U13830 (N_13830,N_11901,N_9761);
xnor U13831 (N_13831,N_10088,N_9353);
and U13832 (N_13832,N_10112,N_11183);
xnor U13833 (N_13833,N_9501,N_10299);
nand U13834 (N_13834,N_10251,N_10429);
and U13835 (N_13835,N_9552,N_10861);
nor U13836 (N_13836,N_10278,N_10582);
and U13837 (N_13837,N_8772,N_9555);
nor U13838 (N_13838,N_11971,N_9821);
and U13839 (N_13839,N_8952,N_9776);
and U13840 (N_13840,N_10876,N_8184);
and U13841 (N_13841,N_10261,N_9338);
or U13842 (N_13842,N_8155,N_9800);
nand U13843 (N_13843,N_11726,N_8922);
or U13844 (N_13844,N_8384,N_8771);
nor U13845 (N_13845,N_10134,N_10409);
or U13846 (N_13846,N_8204,N_11252);
nand U13847 (N_13847,N_11975,N_8060);
and U13848 (N_13848,N_10284,N_9388);
nand U13849 (N_13849,N_9254,N_9739);
nor U13850 (N_13850,N_11298,N_10688);
xnor U13851 (N_13851,N_10985,N_11360);
or U13852 (N_13852,N_8358,N_8162);
and U13853 (N_13853,N_9711,N_10199);
and U13854 (N_13854,N_11030,N_9322);
or U13855 (N_13855,N_9235,N_10755);
nor U13856 (N_13856,N_9526,N_10630);
and U13857 (N_13857,N_9732,N_10629);
and U13858 (N_13858,N_10163,N_10266);
nand U13859 (N_13859,N_9718,N_9725);
nor U13860 (N_13860,N_10186,N_9171);
nor U13861 (N_13861,N_11053,N_8839);
xnor U13862 (N_13862,N_9633,N_8554);
nand U13863 (N_13863,N_8097,N_10559);
and U13864 (N_13864,N_10010,N_9130);
and U13865 (N_13865,N_9514,N_10966);
nand U13866 (N_13866,N_8735,N_8117);
nor U13867 (N_13867,N_9926,N_8253);
and U13868 (N_13868,N_8538,N_10321);
nor U13869 (N_13869,N_9072,N_8212);
nor U13870 (N_13870,N_9214,N_9006);
xnor U13871 (N_13871,N_8572,N_8697);
nand U13872 (N_13872,N_8805,N_9249);
nor U13873 (N_13873,N_8206,N_9822);
and U13874 (N_13874,N_11359,N_8207);
xor U13875 (N_13875,N_11076,N_11784);
xor U13876 (N_13876,N_11173,N_8096);
nor U13877 (N_13877,N_10485,N_9626);
xor U13878 (N_13878,N_10536,N_8250);
or U13879 (N_13879,N_8099,N_10665);
or U13880 (N_13880,N_9421,N_11721);
and U13881 (N_13881,N_11713,N_11265);
and U13882 (N_13882,N_11138,N_10858);
nor U13883 (N_13883,N_9482,N_10557);
nand U13884 (N_13884,N_9103,N_11202);
and U13885 (N_13885,N_10661,N_11912);
nand U13886 (N_13886,N_9174,N_10462);
nand U13887 (N_13887,N_11286,N_10529);
or U13888 (N_13888,N_10908,N_8615);
and U13889 (N_13889,N_11676,N_9104);
or U13890 (N_13890,N_9170,N_8725);
and U13891 (N_13891,N_10927,N_10765);
or U13892 (N_13892,N_8516,N_11299);
or U13893 (N_13893,N_9795,N_8761);
nor U13894 (N_13894,N_8594,N_10190);
nand U13895 (N_13895,N_9371,N_10691);
and U13896 (N_13896,N_9016,N_8114);
or U13897 (N_13897,N_9819,N_10919);
nand U13898 (N_13898,N_10123,N_11987);
nand U13899 (N_13899,N_8627,N_9963);
and U13900 (N_13900,N_11717,N_9912);
nand U13901 (N_13901,N_11953,N_11897);
or U13902 (N_13902,N_10490,N_11414);
nor U13903 (N_13903,N_8770,N_11579);
or U13904 (N_13904,N_10488,N_9629);
or U13905 (N_13905,N_10360,N_11002);
and U13906 (N_13906,N_10555,N_10729);
nand U13907 (N_13907,N_8242,N_11718);
or U13908 (N_13908,N_8501,N_10453);
nor U13909 (N_13909,N_9019,N_11694);
or U13910 (N_13910,N_9051,N_11171);
or U13911 (N_13911,N_8522,N_11444);
nor U13912 (N_13912,N_9342,N_11332);
xor U13913 (N_13913,N_9748,N_11340);
nand U13914 (N_13914,N_9854,N_10542);
nor U13915 (N_13915,N_11715,N_8462);
and U13916 (N_13916,N_9268,N_8508);
or U13917 (N_13917,N_9422,N_9320);
nand U13918 (N_13918,N_11442,N_8248);
or U13919 (N_13919,N_10023,N_8334);
and U13920 (N_13920,N_11993,N_8674);
nor U13921 (N_13921,N_8347,N_11808);
and U13922 (N_13922,N_11734,N_9962);
nand U13923 (N_13923,N_11877,N_9559);
or U13924 (N_13924,N_9241,N_9639);
nand U13925 (N_13925,N_11161,N_10852);
nand U13926 (N_13926,N_8580,N_9203);
and U13927 (N_13927,N_8747,N_9348);
or U13928 (N_13928,N_11380,N_9080);
nor U13929 (N_13929,N_11915,N_8215);
nor U13930 (N_13930,N_10830,N_11850);
nor U13931 (N_13931,N_9172,N_9606);
nand U13932 (N_13932,N_11609,N_9004);
or U13933 (N_13933,N_10119,N_8365);
and U13934 (N_13934,N_11048,N_9523);
or U13935 (N_13935,N_11743,N_10553);
nor U13936 (N_13936,N_10814,N_9304);
or U13937 (N_13937,N_8896,N_11816);
xor U13938 (N_13938,N_10869,N_11693);
xor U13939 (N_13939,N_9769,N_10073);
xor U13940 (N_13940,N_11181,N_11185);
xnor U13941 (N_13941,N_8391,N_11133);
nor U13942 (N_13942,N_8902,N_10272);
nand U13943 (N_13943,N_8229,N_10050);
and U13944 (N_13944,N_8328,N_10747);
or U13945 (N_13945,N_11757,N_11408);
or U13946 (N_13946,N_8047,N_9667);
nand U13947 (N_13947,N_9499,N_11554);
and U13948 (N_13948,N_8866,N_10930);
or U13949 (N_13949,N_11681,N_8537);
nor U13950 (N_13950,N_11547,N_10885);
xor U13951 (N_13951,N_9381,N_11548);
nor U13952 (N_13952,N_11782,N_10897);
and U13953 (N_13953,N_8686,N_8189);
nor U13954 (N_13954,N_10377,N_10812);
and U13955 (N_13955,N_9039,N_10466);
and U13956 (N_13956,N_11434,N_10327);
nor U13957 (N_13957,N_11418,N_10441);
nor U13958 (N_13958,N_11831,N_11009);
nor U13959 (N_13959,N_11977,N_8862);
and U13960 (N_13960,N_9444,N_8991);
and U13961 (N_13961,N_11770,N_10116);
or U13962 (N_13962,N_10570,N_8164);
nand U13963 (N_13963,N_11038,N_8901);
xnor U13964 (N_13964,N_9852,N_11457);
or U13965 (N_13965,N_9681,N_9185);
nor U13966 (N_13966,N_10587,N_11371);
or U13967 (N_13967,N_9406,N_11337);
or U13968 (N_13968,N_8573,N_11732);
nor U13969 (N_13969,N_8708,N_10172);
xnor U13970 (N_13970,N_11895,N_10645);
nor U13971 (N_13971,N_11807,N_8435);
nor U13972 (N_13972,N_11085,N_9562);
and U13973 (N_13973,N_9048,N_8302);
nand U13974 (N_13974,N_11336,N_11758);
and U13975 (N_13975,N_8313,N_10049);
and U13976 (N_13976,N_9043,N_8078);
nor U13977 (N_13977,N_11162,N_11985);
or U13978 (N_13978,N_10391,N_8090);
nor U13979 (N_13979,N_11366,N_9425);
xor U13980 (N_13980,N_9102,N_9907);
and U13981 (N_13981,N_9133,N_9135);
nor U13982 (N_13982,N_9884,N_9334);
or U13983 (N_13983,N_10359,N_10695);
or U13984 (N_13984,N_8510,N_9914);
and U13985 (N_13985,N_11720,N_9588);
nor U13986 (N_13986,N_11781,N_9908);
or U13987 (N_13987,N_8712,N_11776);
or U13988 (N_13988,N_11928,N_10888);
nand U13989 (N_13989,N_11264,N_8941);
and U13990 (N_13990,N_11526,N_11040);
nand U13991 (N_13991,N_11244,N_9850);
or U13992 (N_13992,N_8022,N_8848);
nor U13993 (N_13993,N_8676,N_10849);
or U13994 (N_13994,N_10253,N_11235);
and U13995 (N_13995,N_8425,N_10738);
nor U13996 (N_13996,N_9762,N_11338);
and U13997 (N_13997,N_8268,N_8518);
and U13998 (N_13998,N_10303,N_9996);
and U13999 (N_13999,N_8870,N_8729);
nand U14000 (N_14000,N_10940,N_9504);
nand U14001 (N_14001,N_11522,N_11575);
or U14002 (N_14002,N_9010,N_11987);
nor U14003 (N_14003,N_8492,N_8707);
xnor U14004 (N_14004,N_8765,N_9849);
nor U14005 (N_14005,N_9809,N_9254);
and U14006 (N_14006,N_8809,N_9526);
or U14007 (N_14007,N_11209,N_11204);
nand U14008 (N_14008,N_9786,N_10804);
nor U14009 (N_14009,N_8573,N_9662);
nand U14010 (N_14010,N_10167,N_8600);
or U14011 (N_14011,N_11917,N_9798);
nor U14012 (N_14012,N_11483,N_8592);
or U14013 (N_14013,N_10848,N_8135);
nand U14014 (N_14014,N_9331,N_10160);
nor U14015 (N_14015,N_9442,N_10378);
or U14016 (N_14016,N_9573,N_10214);
xor U14017 (N_14017,N_11399,N_10285);
nand U14018 (N_14018,N_11770,N_10190);
nor U14019 (N_14019,N_9677,N_11970);
nand U14020 (N_14020,N_8081,N_8918);
nor U14021 (N_14021,N_8304,N_8831);
nand U14022 (N_14022,N_11451,N_11944);
xor U14023 (N_14023,N_8040,N_8212);
or U14024 (N_14024,N_11947,N_8690);
or U14025 (N_14025,N_8663,N_11763);
nand U14026 (N_14026,N_10590,N_10379);
nand U14027 (N_14027,N_11511,N_11683);
nand U14028 (N_14028,N_10565,N_8791);
nor U14029 (N_14029,N_8462,N_9265);
and U14030 (N_14030,N_10920,N_10688);
nand U14031 (N_14031,N_11566,N_8735);
and U14032 (N_14032,N_9412,N_10987);
and U14033 (N_14033,N_10656,N_10240);
and U14034 (N_14034,N_10791,N_9675);
nand U14035 (N_14035,N_10248,N_9645);
or U14036 (N_14036,N_11359,N_11267);
or U14037 (N_14037,N_8910,N_11145);
nand U14038 (N_14038,N_8866,N_8053);
nor U14039 (N_14039,N_10500,N_9085);
nor U14040 (N_14040,N_11205,N_9942);
and U14041 (N_14041,N_9607,N_10552);
and U14042 (N_14042,N_10979,N_9508);
and U14043 (N_14043,N_10138,N_10706);
xnor U14044 (N_14044,N_8644,N_10657);
nor U14045 (N_14045,N_10294,N_10596);
xnor U14046 (N_14046,N_9759,N_8228);
nand U14047 (N_14047,N_9644,N_8804);
nor U14048 (N_14048,N_10176,N_11211);
nand U14049 (N_14049,N_11747,N_8034);
and U14050 (N_14050,N_11300,N_10696);
nor U14051 (N_14051,N_10869,N_8690);
or U14052 (N_14052,N_10455,N_10989);
or U14053 (N_14053,N_10049,N_11485);
nor U14054 (N_14054,N_9535,N_9667);
nand U14055 (N_14055,N_10326,N_8779);
nand U14056 (N_14056,N_11931,N_11283);
nand U14057 (N_14057,N_8262,N_10449);
nand U14058 (N_14058,N_8649,N_8425);
nor U14059 (N_14059,N_10516,N_11849);
or U14060 (N_14060,N_11919,N_8901);
or U14061 (N_14061,N_8369,N_8601);
nor U14062 (N_14062,N_8796,N_11991);
xor U14063 (N_14063,N_11652,N_8774);
or U14064 (N_14064,N_10652,N_8335);
nand U14065 (N_14065,N_8167,N_10130);
nand U14066 (N_14066,N_11645,N_11288);
or U14067 (N_14067,N_8276,N_9820);
nand U14068 (N_14068,N_8540,N_11066);
and U14069 (N_14069,N_8680,N_10784);
and U14070 (N_14070,N_9268,N_10163);
nand U14071 (N_14071,N_9619,N_8801);
and U14072 (N_14072,N_10936,N_11852);
and U14073 (N_14073,N_9388,N_11149);
and U14074 (N_14074,N_9634,N_10145);
nor U14075 (N_14075,N_11466,N_9970);
or U14076 (N_14076,N_10831,N_8674);
nor U14077 (N_14077,N_8571,N_11546);
or U14078 (N_14078,N_11008,N_10870);
nand U14079 (N_14079,N_8156,N_11038);
nand U14080 (N_14080,N_9123,N_9281);
xnor U14081 (N_14081,N_10330,N_10302);
or U14082 (N_14082,N_9033,N_8008);
nand U14083 (N_14083,N_10397,N_8534);
or U14084 (N_14084,N_9603,N_9718);
nand U14085 (N_14085,N_10117,N_10760);
nand U14086 (N_14086,N_11341,N_9493);
nand U14087 (N_14087,N_11207,N_8792);
xnor U14088 (N_14088,N_10618,N_10601);
nand U14089 (N_14089,N_8804,N_9954);
xnor U14090 (N_14090,N_8000,N_11751);
xnor U14091 (N_14091,N_10122,N_8744);
or U14092 (N_14092,N_9206,N_10809);
or U14093 (N_14093,N_9906,N_11904);
xor U14094 (N_14094,N_8774,N_8549);
nand U14095 (N_14095,N_10881,N_8085);
nand U14096 (N_14096,N_9777,N_8930);
and U14097 (N_14097,N_8872,N_11908);
nand U14098 (N_14098,N_9746,N_11582);
and U14099 (N_14099,N_10099,N_10948);
or U14100 (N_14100,N_8187,N_8209);
nor U14101 (N_14101,N_11867,N_9680);
or U14102 (N_14102,N_10233,N_9867);
nand U14103 (N_14103,N_11746,N_11811);
nand U14104 (N_14104,N_8737,N_10343);
nor U14105 (N_14105,N_9502,N_8993);
and U14106 (N_14106,N_11759,N_11186);
nand U14107 (N_14107,N_9812,N_11725);
xor U14108 (N_14108,N_10096,N_10104);
nor U14109 (N_14109,N_10085,N_10046);
or U14110 (N_14110,N_8519,N_10226);
nand U14111 (N_14111,N_9573,N_11178);
and U14112 (N_14112,N_10207,N_11127);
or U14113 (N_14113,N_9417,N_8759);
xnor U14114 (N_14114,N_9333,N_8542);
or U14115 (N_14115,N_11464,N_10525);
nand U14116 (N_14116,N_11169,N_8787);
nand U14117 (N_14117,N_8443,N_11533);
nor U14118 (N_14118,N_9075,N_9805);
xnor U14119 (N_14119,N_8973,N_9392);
or U14120 (N_14120,N_8453,N_10799);
nor U14121 (N_14121,N_9633,N_10633);
nand U14122 (N_14122,N_11278,N_11346);
nor U14123 (N_14123,N_11984,N_11508);
or U14124 (N_14124,N_9566,N_8339);
or U14125 (N_14125,N_10686,N_8378);
nand U14126 (N_14126,N_11087,N_8717);
or U14127 (N_14127,N_9375,N_11021);
nor U14128 (N_14128,N_8499,N_11629);
nor U14129 (N_14129,N_9228,N_11527);
or U14130 (N_14130,N_10974,N_11628);
nand U14131 (N_14131,N_10190,N_10555);
nor U14132 (N_14132,N_8939,N_10968);
nor U14133 (N_14133,N_11879,N_11421);
xnor U14134 (N_14134,N_8822,N_10244);
and U14135 (N_14135,N_10719,N_8800);
and U14136 (N_14136,N_10359,N_11977);
nand U14137 (N_14137,N_11664,N_8403);
or U14138 (N_14138,N_10986,N_8855);
xor U14139 (N_14139,N_9651,N_8418);
xor U14140 (N_14140,N_10749,N_10347);
or U14141 (N_14141,N_10667,N_9533);
nor U14142 (N_14142,N_8840,N_9520);
nor U14143 (N_14143,N_8454,N_9016);
nor U14144 (N_14144,N_11502,N_9915);
xnor U14145 (N_14145,N_11271,N_10598);
and U14146 (N_14146,N_11936,N_10666);
xor U14147 (N_14147,N_11736,N_10279);
nand U14148 (N_14148,N_8199,N_11305);
nand U14149 (N_14149,N_10947,N_11847);
nor U14150 (N_14150,N_8259,N_11423);
nor U14151 (N_14151,N_8950,N_8351);
xor U14152 (N_14152,N_9305,N_10517);
nor U14153 (N_14153,N_8608,N_10193);
and U14154 (N_14154,N_8050,N_8526);
nand U14155 (N_14155,N_10622,N_8457);
nor U14156 (N_14156,N_8170,N_9078);
nand U14157 (N_14157,N_8906,N_11547);
xor U14158 (N_14158,N_11272,N_10615);
nand U14159 (N_14159,N_9434,N_11294);
and U14160 (N_14160,N_9045,N_8621);
nor U14161 (N_14161,N_10672,N_8873);
nand U14162 (N_14162,N_9028,N_10237);
and U14163 (N_14163,N_9651,N_9021);
nand U14164 (N_14164,N_8850,N_9781);
or U14165 (N_14165,N_10837,N_10264);
nand U14166 (N_14166,N_8566,N_8691);
nor U14167 (N_14167,N_10154,N_8429);
and U14168 (N_14168,N_11906,N_8554);
and U14169 (N_14169,N_9029,N_8354);
nand U14170 (N_14170,N_10060,N_9732);
or U14171 (N_14171,N_11648,N_11066);
xnor U14172 (N_14172,N_8037,N_9977);
nor U14173 (N_14173,N_8678,N_9772);
and U14174 (N_14174,N_10089,N_8680);
xnor U14175 (N_14175,N_11391,N_8244);
nand U14176 (N_14176,N_8090,N_8122);
nand U14177 (N_14177,N_9695,N_8501);
nand U14178 (N_14178,N_11455,N_11809);
or U14179 (N_14179,N_10368,N_11162);
or U14180 (N_14180,N_11281,N_10694);
xnor U14181 (N_14181,N_8102,N_8304);
nand U14182 (N_14182,N_9295,N_10058);
nor U14183 (N_14183,N_9098,N_11910);
and U14184 (N_14184,N_11695,N_10361);
xor U14185 (N_14185,N_9053,N_11392);
or U14186 (N_14186,N_10764,N_9824);
nand U14187 (N_14187,N_9492,N_11799);
nand U14188 (N_14188,N_9734,N_9304);
and U14189 (N_14189,N_10329,N_9601);
nand U14190 (N_14190,N_9451,N_8492);
or U14191 (N_14191,N_10847,N_10054);
or U14192 (N_14192,N_8686,N_8078);
or U14193 (N_14193,N_9790,N_9619);
nor U14194 (N_14194,N_11807,N_11249);
and U14195 (N_14195,N_11232,N_11348);
nor U14196 (N_14196,N_9447,N_9953);
xor U14197 (N_14197,N_11823,N_8244);
xnor U14198 (N_14198,N_10009,N_9709);
nor U14199 (N_14199,N_9285,N_8438);
or U14200 (N_14200,N_9921,N_8729);
nand U14201 (N_14201,N_10801,N_11319);
nor U14202 (N_14202,N_8222,N_8273);
xor U14203 (N_14203,N_11968,N_10839);
xnor U14204 (N_14204,N_8028,N_10728);
or U14205 (N_14205,N_11870,N_9943);
and U14206 (N_14206,N_11240,N_9501);
nor U14207 (N_14207,N_8766,N_9158);
nand U14208 (N_14208,N_11696,N_10486);
nor U14209 (N_14209,N_9294,N_9704);
xnor U14210 (N_14210,N_11431,N_9409);
and U14211 (N_14211,N_8290,N_9489);
nor U14212 (N_14212,N_10630,N_9229);
and U14213 (N_14213,N_9176,N_9729);
or U14214 (N_14214,N_10211,N_11362);
nor U14215 (N_14215,N_8607,N_8964);
or U14216 (N_14216,N_9367,N_10261);
nor U14217 (N_14217,N_10074,N_10867);
or U14218 (N_14218,N_9101,N_11048);
nand U14219 (N_14219,N_9210,N_11365);
and U14220 (N_14220,N_11925,N_11580);
nor U14221 (N_14221,N_11817,N_10973);
and U14222 (N_14222,N_8703,N_11465);
and U14223 (N_14223,N_10963,N_10639);
nor U14224 (N_14224,N_9138,N_11722);
or U14225 (N_14225,N_11253,N_11702);
and U14226 (N_14226,N_11514,N_9506);
xor U14227 (N_14227,N_8147,N_8924);
or U14228 (N_14228,N_11525,N_9637);
nand U14229 (N_14229,N_11018,N_11334);
nand U14230 (N_14230,N_11432,N_10053);
and U14231 (N_14231,N_8468,N_11307);
xnor U14232 (N_14232,N_10349,N_11510);
xor U14233 (N_14233,N_9537,N_11462);
xnor U14234 (N_14234,N_9619,N_9711);
and U14235 (N_14235,N_10816,N_11720);
nand U14236 (N_14236,N_8842,N_11386);
nor U14237 (N_14237,N_8118,N_8999);
and U14238 (N_14238,N_8526,N_11574);
nand U14239 (N_14239,N_8234,N_11695);
and U14240 (N_14240,N_11240,N_11980);
nand U14241 (N_14241,N_10646,N_9520);
and U14242 (N_14242,N_9456,N_10786);
or U14243 (N_14243,N_9738,N_11533);
and U14244 (N_14244,N_10850,N_8065);
or U14245 (N_14245,N_8183,N_9964);
and U14246 (N_14246,N_9075,N_8151);
nand U14247 (N_14247,N_8634,N_8185);
and U14248 (N_14248,N_11051,N_9419);
nand U14249 (N_14249,N_11666,N_11308);
or U14250 (N_14250,N_10507,N_9064);
and U14251 (N_14251,N_8024,N_10363);
or U14252 (N_14252,N_11596,N_10475);
or U14253 (N_14253,N_10085,N_8481);
and U14254 (N_14254,N_8703,N_10157);
and U14255 (N_14255,N_11537,N_10015);
nand U14256 (N_14256,N_10675,N_9724);
nor U14257 (N_14257,N_9988,N_10866);
or U14258 (N_14258,N_11913,N_9405);
and U14259 (N_14259,N_8384,N_10918);
and U14260 (N_14260,N_9110,N_9215);
xnor U14261 (N_14261,N_11367,N_11244);
and U14262 (N_14262,N_10802,N_8963);
or U14263 (N_14263,N_10292,N_11822);
nor U14264 (N_14264,N_9169,N_9775);
or U14265 (N_14265,N_8727,N_8440);
and U14266 (N_14266,N_8459,N_10421);
nor U14267 (N_14267,N_11734,N_10625);
nor U14268 (N_14268,N_11542,N_10585);
nand U14269 (N_14269,N_10339,N_11499);
nand U14270 (N_14270,N_9473,N_11379);
xor U14271 (N_14271,N_11474,N_8779);
nor U14272 (N_14272,N_11216,N_8845);
nor U14273 (N_14273,N_11139,N_9114);
or U14274 (N_14274,N_9894,N_8678);
and U14275 (N_14275,N_10264,N_8089);
nand U14276 (N_14276,N_8044,N_11290);
nor U14277 (N_14277,N_11305,N_10920);
and U14278 (N_14278,N_9024,N_10876);
and U14279 (N_14279,N_10460,N_8033);
nand U14280 (N_14280,N_10448,N_8223);
and U14281 (N_14281,N_8460,N_10111);
nand U14282 (N_14282,N_9560,N_10633);
nand U14283 (N_14283,N_11550,N_9504);
nor U14284 (N_14284,N_11648,N_9367);
or U14285 (N_14285,N_8799,N_9591);
or U14286 (N_14286,N_11801,N_11977);
xor U14287 (N_14287,N_11567,N_8469);
or U14288 (N_14288,N_11306,N_9999);
nor U14289 (N_14289,N_11208,N_11385);
nor U14290 (N_14290,N_8639,N_8308);
nand U14291 (N_14291,N_9414,N_8270);
or U14292 (N_14292,N_8733,N_8574);
nor U14293 (N_14293,N_8918,N_10480);
and U14294 (N_14294,N_8053,N_8434);
nand U14295 (N_14295,N_10168,N_10517);
and U14296 (N_14296,N_10166,N_9106);
nand U14297 (N_14297,N_8285,N_10431);
nand U14298 (N_14298,N_8401,N_10085);
xnor U14299 (N_14299,N_10206,N_11267);
or U14300 (N_14300,N_8119,N_11707);
or U14301 (N_14301,N_8108,N_8300);
or U14302 (N_14302,N_10178,N_11677);
and U14303 (N_14303,N_10637,N_11858);
or U14304 (N_14304,N_8706,N_8947);
nand U14305 (N_14305,N_10964,N_8766);
nor U14306 (N_14306,N_8259,N_8826);
nand U14307 (N_14307,N_9336,N_8759);
xnor U14308 (N_14308,N_11304,N_8404);
and U14309 (N_14309,N_8689,N_11343);
and U14310 (N_14310,N_9218,N_8010);
nand U14311 (N_14311,N_11168,N_9052);
xnor U14312 (N_14312,N_8557,N_9603);
nand U14313 (N_14313,N_10305,N_8493);
and U14314 (N_14314,N_8722,N_10063);
nor U14315 (N_14315,N_9895,N_9243);
and U14316 (N_14316,N_8856,N_9667);
nand U14317 (N_14317,N_10198,N_10137);
or U14318 (N_14318,N_10105,N_8185);
nand U14319 (N_14319,N_8988,N_11996);
and U14320 (N_14320,N_8362,N_9873);
nor U14321 (N_14321,N_9766,N_9346);
nor U14322 (N_14322,N_9921,N_8390);
nand U14323 (N_14323,N_8636,N_8417);
nor U14324 (N_14324,N_8308,N_9061);
xnor U14325 (N_14325,N_11656,N_9719);
or U14326 (N_14326,N_11269,N_9558);
or U14327 (N_14327,N_8359,N_9920);
nor U14328 (N_14328,N_8629,N_9819);
xor U14329 (N_14329,N_11859,N_10746);
and U14330 (N_14330,N_8278,N_9282);
and U14331 (N_14331,N_10985,N_8775);
nor U14332 (N_14332,N_8082,N_8771);
xor U14333 (N_14333,N_8892,N_8485);
nor U14334 (N_14334,N_10045,N_8406);
or U14335 (N_14335,N_10924,N_8689);
and U14336 (N_14336,N_8011,N_8639);
or U14337 (N_14337,N_11534,N_9294);
xor U14338 (N_14338,N_11868,N_10726);
nand U14339 (N_14339,N_10496,N_9199);
xnor U14340 (N_14340,N_11743,N_10851);
or U14341 (N_14341,N_8559,N_11133);
and U14342 (N_14342,N_11701,N_8505);
or U14343 (N_14343,N_9606,N_10380);
xor U14344 (N_14344,N_11022,N_9601);
or U14345 (N_14345,N_11712,N_9410);
nand U14346 (N_14346,N_8347,N_11940);
or U14347 (N_14347,N_11883,N_9385);
nand U14348 (N_14348,N_9554,N_10709);
nor U14349 (N_14349,N_10879,N_10518);
nor U14350 (N_14350,N_11396,N_10184);
or U14351 (N_14351,N_11691,N_10911);
nor U14352 (N_14352,N_8160,N_8283);
nor U14353 (N_14353,N_10362,N_11379);
and U14354 (N_14354,N_8064,N_8362);
and U14355 (N_14355,N_11758,N_10183);
and U14356 (N_14356,N_11360,N_8636);
nor U14357 (N_14357,N_11536,N_8501);
or U14358 (N_14358,N_8719,N_9057);
xor U14359 (N_14359,N_10761,N_11654);
nand U14360 (N_14360,N_9430,N_8238);
nor U14361 (N_14361,N_9534,N_9905);
and U14362 (N_14362,N_8467,N_9135);
nor U14363 (N_14363,N_11754,N_11895);
xnor U14364 (N_14364,N_8865,N_11303);
nor U14365 (N_14365,N_8052,N_10300);
and U14366 (N_14366,N_8550,N_10692);
xnor U14367 (N_14367,N_9438,N_8357);
nand U14368 (N_14368,N_9980,N_10232);
nor U14369 (N_14369,N_9715,N_10903);
or U14370 (N_14370,N_8934,N_9392);
or U14371 (N_14371,N_10976,N_10773);
or U14372 (N_14372,N_8498,N_11104);
nor U14373 (N_14373,N_8764,N_9315);
and U14374 (N_14374,N_10174,N_10862);
and U14375 (N_14375,N_9496,N_11047);
nand U14376 (N_14376,N_10455,N_11569);
or U14377 (N_14377,N_10474,N_11662);
nand U14378 (N_14378,N_11715,N_10164);
nand U14379 (N_14379,N_9112,N_9294);
nor U14380 (N_14380,N_10996,N_11464);
xor U14381 (N_14381,N_10029,N_11897);
nor U14382 (N_14382,N_11448,N_10043);
nand U14383 (N_14383,N_10120,N_10681);
nor U14384 (N_14384,N_8958,N_8562);
nand U14385 (N_14385,N_10948,N_9058);
or U14386 (N_14386,N_11843,N_9789);
and U14387 (N_14387,N_11727,N_8911);
and U14388 (N_14388,N_8925,N_10922);
nor U14389 (N_14389,N_9295,N_8964);
nor U14390 (N_14390,N_10678,N_9869);
and U14391 (N_14391,N_10046,N_11942);
xor U14392 (N_14392,N_11466,N_10105);
nor U14393 (N_14393,N_8795,N_10076);
nor U14394 (N_14394,N_9569,N_9725);
and U14395 (N_14395,N_9735,N_10521);
xnor U14396 (N_14396,N_11633,N_10363);
and U14397 (N_14397,N_10558,N_11072);
nand U14398 (N_14398,N_10393,N_11551);
nor U14399 (N_14399,N_10101,N_10689);
or U14400 (N_14400,N_8524,N_9058);
or U14401 (N_14401,N_9712,N_11616);
nand U14402 (N_14402,N_11503,N_11489);
and U14403 (N_14403,N_10839,N_8967);
and U14404 (N_14404,N_11305,N_11237);
nor U14405 (N_14405,N_10170,N_10777);
nor U14406 (N_14406,N_9186,N_9982);
or U14407 (N_14407,N_10427,N_11077);
and U14408 (N_14408,N_11254,N_8824);
and U14409 (N_14409,N_10566,N_11613);
nand U14410 (N_14410,N_11606,N_9493);
or U14411 (N_14411,N_8607,N_11332);
and U14412 (N_14412,N_10112,N_11271);
or U14413 (N_14413,N_8572,N_9787);
nand U14414 (N_14414,N_10309,N_8558);
nand U14415 (N_14415,N_10061,N_8043);
xor U14416 (N_14416,N_11358,N_8506);
or U14417 (N_14417,N_10483,N_11225);
nand U14418 (N_14418,N_11421,N_10640);
or U14419 (N_14419,N_8546,N_11536);
or U14420 (N_14420,N_8954,N_9555);
or U14421 (N_14421,N_8881,N_9250);
nand U14422 (N_14422,N_10147,N_8286);
nand U14423 (N_14423,N_9439,N_10935);
or U14424 (N_14424,N_8067,N_10427);
or U14425 (N_14425,N_11350,N_11992);
nand U14426 (N_14426,N_11492,N_9388);
nand U14427 (N_14427,N_8027,N_10100);
nor U14428 (N_14428,N_9821,N_10773);
nor U14429 (N_14429,N_9208,N_8405);
nor U14430 (N_14430,N_8911,N_11445);
nor U14431 (N_14431,N_9096,N_8027);
xnor U14432 (N_14432,N_10838,N_10188);
nor U14433 (N_14433,N_8356,N_10497);
and U14434 (N_14434,N_11636,N_11939);
nor U14435 (N_14435,N_10931,N_8256);
and U14436 (N_14436,N_10018,N_8806);
and U14437 (N_14437,N_9647,N_11249);
and U14438 (N_14438,N_8456,N_10952);
or U14439 (N_14439,N_8235,N_9220);
nand U14440 (N_14440,N_10040,N_11939);
or U14441 (N_14441,N_9670,N_8462);
and U14442 (N_14442,N_11941,N_10157);
nand U14443 (N_14443,N_10816,N_10762);
and U14444 (N_14444,N_9639,N_8730);
nor U14445 (N_14445,N_9513,N_9667);
nand U14446 (N_14446,N_8666,N_8550);
and U14447 (N_14447,N_9778,N_8526);
nor U14448 (N_14448,N_10583,N_8769);
and U14449 (N_14449,N_10844,N_9547);
nand U14450 (N_14450,N_9561,N_10256);
xnor U14451 (N_14451,N_11963,N_10268);
nor U14452 (N_14452,N_9676,N_11247);
or U14453 (N_14453,N_9559,N_11570);
nor U14454 (N_14454,N_11870,N_11898);
xnor U14455 (N_14455,N_8588,N_9015);
or U14456 (N_14456,N_10390,N_10555);
nand U14457 (N_14457,N_9884,N_8660);
nand U14458 (N_14458,N_9171,N_8021);
nor U14459 (N_14459,N_9225,N_10064);
and U14460 (N_14460,N_11034,N_10880);
xnor U14461 (N_14461,N_10795,N_8976);
nor U14462 (N_14462,N_10942,N_11776);
or U14463 (N_14463,N_9712,N_10866);
and U14464 (N_14464,N_9576,N_9140);
nor U14465 (N_14465,N_9455,N_10934);
nand U14466 (N_14466,N_8205,N_9149);
and U14467 (N_14467,N_8345,N_9117);
or U14468 (N_14468,N_10353,N_8782);
nand U14469 (N_14469,N_9422,N_9154);
nand U14470 (N_14470,N_10973,N_8285);
or U14471 (N_14471,N_10417,N_9528);
nand U14472 (N_14472,N_9860,N_11726);
nor U14473 (N_14473,N_10004,N_10525);
or U14474 (N_14474,N_10839,N_8503);
xor U14475 (N_14475,N_8223,N_11355);
nor U14476 (N_14476,N_8596,N_9764);
and U14477 (N_14477,N_9026,N_10233);
or U14478 (N_14478,N_10839,N_9940);
nand U14479 (N_14479,N_11553,N_9358);
and U14480 (N_14480,N_10720,N_11773);
and U14481 (N_14481,N_11702,N_9446);
nor U14482 (N_14482,N_8009,N_10385);
or U14483 (N_14483,N_9778,N_11508);
nor U14484 (N_14484,N_8077,N_11138);
xor U14485 (N_14485,N_11852,N_9374);
nand U14486 (N_14486,N_8478,N_10521);
nor U14487 (N_14487,N_9135,N_10151);
or U14488 (N_14488,N_10380,N_8513);
and U14489 (N_14489,N_10877,N_11471);
nand U14490 (N_14490,N_9322,N_8503);
nand U14491 (N_14491,N_9306,N_9210);
nand U14492 (N_14492,N_8038,N_8690);
and U14493 (N_14493,N_9900,N_10419);
and U14494 (N_14494,N_10591,N_11858);
or U14495 (N_14495,N_10958,N_9530);
or U14496 (N_14496,N_10159,N_11163);
nor U14497 (N_14497,N_11256,N_10022);
and U14498 (N_14498,N_10706,N_9652);
or U14499 (N_14499,N_8812,N_10764);
and U14500 (N_14500,N_11476,N_8926);
nand U14501 (N_14501,N_11449,N_8693);
nand U14502 (N_14502,N_9911,N_9332);
xor U14503 (N_14503,N_11332,N_11286);
nor U14504 (N_14504,N_9651,N_11138);
or U14505 (N_14505,N_8960,N_9770);
nand U14506 (N_14506,N_11406,N_9826);
nand U14507 (N_14507,N_9753,N_11982);
nand U14508 (N_14508,N_11406,N_10934);
nand U14509 (N_14509,N_11623,N_10544);
nand U14510 (N_14510,N_9556,N_10802);
and U14511 (N_14511,N_9183,N_9090);
nand U14512 (N_14512,N_9277,N_10424);
and U14513 (N_14513,N_10551,N_11687);
nand U14514 (N_14514,N_11476,N_10901);
nand U14515 (N_14515,N_9798,N_10723);
and U14516 (N_14516,N_9193,N_10267);
xor U14517 (N_14517,N_10928,N_10504);
xor U14518 (N_14518,N_11401,N_9563);
and U14519 (N_14519,N_9193,N_8626);
and U14520 (N_14520,N_8110,N_9159);
nor U14521 (N_14521,N_9176,N_8836);
xor U14522 (N_14522,N_11816,N_8972);
nor U14523 (N_14523,N_10455,N_8032);
or U14524 (N_14524,N_11562,N_9853);
xnor U14525 (N_14525,N_9313,N_8791);
and U14526 (N_14526,N_10460,N_8993);
nand U14527 (N_14527,N_8514,N_11647);
nor U14528 (N_14528,N_10423,N_11700);
nand U14529 (N_14529,N_8149,N_11746);
or U14530 (N_14530,N_8617,N_9828);
and U14531 (N_14531,N_8384,N_10434);
nand U14532 (N_14532,N_8362,N_11022);
nor U14533 (N_14533,N_11824,N_8251);
nand U14534 (N_14534,N_10456,N_9341);
xnor U14535 (N_14535,N_9754,N_9908);
or U14536 (N_14536,N_11923,N_8103);
xor U14537 (N_14537,N_11488,N_9015);
xor U14538 (N_14538,N_8800,N_11056);
or U14539 (N_14539,N_8740,N_11985);
nor U14540 (N_14540,N_9240,N_11297);
nand U14541 (N_14541,N_11253,N_8062);
or U14542 (N_14542,N_8922,N_10248);
nor U14543 (N_14543,N_11478,N_8394);
xnor U14544 (N_14544,N_11070,N_9510);
and U14545 (N_14545,N_9703,N_10536);
nor U14546 (N_14546,N_9544,N_8374);
xnor U14547 (N_14547,N_8892,N_11729);
or U14548 (N_14548,N_9423,N_10559);
and U14549 (N_14549,N_10078,N_11430);
nor U14550 (N_14550,N_10827,N_9771);
nand U14551 (N_14551,N_11187,N_9836);
or U14552 (N_14552,N_10242,N_10775);
xor U14553 (N_14553,N_11315,N_11765);
nor U14554 (N_14554,N_10446,N_8454);
or U14555 (N_14555,N_11503,N_9734);
or U14556 (N_14556,N_10698,N_9896);
and U14557 (N_14557,N_9180,N_10902);
or U14558 (N_14558,N_9060,N_11019);
nor U14559 (N_14559,N_10227,N_9808);
or U14560 (N_14560,N_8177,N_9934);
or U14561 (N_14561,N_10334,N_10548);
or U14562 (N_14562,N_11611,N_8087);
and U14563 (N_14563,N_11673,N_10196);
or U14564 (N_14564,N_10539,N_11246);
xnor U14565 (N_14565,N_8396,N_11379);
or U14566 (N_14566,N_11299,N_11960);
or U14567 (N_14567,N_11322,N_8825);
xor U14568 (N_14568,N_10404,N_11711);
xnor U14569 (N_14569,N_11144,N_11982);
nor U14570 (N_14570,N_11672,N_9867);
and U14571 (N_14571,N_11946,N_10895);
nor U14572 (N_14572,N_9125,N_9787);
nor U14573 (N_14573,N_10342,N_8094);
nor U14574 (N_14574,N_9829,N_8448);
xnor U14575 (N_14575,N_8708,N_10560);
nand U14576 (N_14576,N_10011,N_9280);
nor U14577 (N_14577,N_11555,N_8458);
nor U14578 (N_14578,N_9172,N_8878);
nor U14579 (N_14579,N_9133,N_11575);
nand U14580 (N_14580,N_10763,N_11212);
nand U14581 (N_14581,N_11856,N_10903);
and U14582 (N_14582,N_8865,N_11853);
nand U14583 (N_14583,N_9050,N_11880);
nand U14584 (N_14584,N_11558,N_10407);
nor U14585 (N_14585,N_10951,N_8473);
or U14586 (N_14586,N_11735,N_10747);
nand U14587 (N_14587,N_11340,N_9603);
xnor U14588 (N_14588,N_10352,N_8147);
and U14589 (N_14589,N_9091,N_8140);
and U14590 (N_14590,N_10991,N_8455);
or U14591 (N_14591,N_9358,N_10964);
or U14592 (N_14592,N_8877,N_10352);
or U14593 (N_14593,N_10338,N_8369);
and U14594 (N_14594,N_11232,N_9418);
and U14595 (N_14595,N_9765,N_11041);
nand U14596 (N_14596,N_9134,N_8038);
or U14597 (N_14597,N_9284,N_9883);
and U14598 (N_14598,N_10896,N_8473);
nor U14599 (N_14599,N_11395,N_11068);
nor U14600 (N_14600,N_11312,N_10152);
nor U14601 (N_14601,N_9083,N_8715);
nand U14602 (N_14602,N_9180,N_8438);
and U14603 (N_14603,N_9589,N_11516);
nand U14604 (N_14604,N_8612,N_9736);
nor U14605 (N_14605,N_11118,N_9090);
nand U14606 (N_14606,N_8489,N_10952);
or U14607 (N_14607,N_8847,N_11535);
nand U14608 (N_14608,N_9514,N_9569);
nand U14609 (N_14609,N_9172,N_10582);
nand U14610 (N_14610,N_9644,N_8136);
or U14611 (N_14611,N_8276,N_8065);
or U14612 (N_14612,N_10460,N_11570);
and U14613 (N_14613,N_10357,N_10417);
xor U14614 (N_14614,N_10021,N_11842);
or U14615 (N_14615,N_9492,N_9564);
nand U14616 (N_14616,N_9453,N_10443);
and U14617 (N_14617,N_9972,N_11309);
nor U14618 (N_14618,N_8576,N_8765);
or U14619 (N_14619,N_11197,N_11116);
nand U14620 (N_14620,N_11894,N_9714);
nor U14621 (N_14621,N_11339,N_9246);
nand U14622 (N_14622,N_9979,N_10838);
xnor U14623 (N_14623,N_8990,N_9131);
and U14624 (N_14624,N_9387,N_11114);
nand U14625 (N_14625,N_9037,N_11875);
nand U14626 (N_14626,N_11512,N_9324);
and U14627 (N_14627,N_9593,N_10350);
nand U14628 (N_14628,N_10659,N_11643);
and U14629 (N_14629,N_8142,N_8731);
nor U14630 (N_14630,N_11221,N_10421);
and U14631 (N_14631,N_8568,N_8266);
or U14632 (N_14632,N_10458,N_8643);
nor U14633 (N_14633,N_9652,N_10700);
or U14634 (N_14634,N_9546,N_9414);
and U14635 (N_14635,N_11955,N_10045);
and U14636 (N_14636,N_11343,N_10136);
nor U14637 (N_14637,N_10354,N_11863);
xor U14638 (N_14638,N_10383,N_8999);
nand U14639 (N_14639,N_10924,N_8287);
and U14640 (N_14640,N_9212,N_9772);
or U14641 (N_14641,N_11080,N_10598);
xnor U14642 (N_14642,N_10252,N_11985);
and U14643 (N_14643,N_9871,N_9835);
or U14644 (N_14644,N_9613,N_11339);
nor U14645 (N_14645,N_8739,N_9958);
nor U14646 (N_14646,N_9949,N_8876);
nand U14647 (N_14647,N_11994,N_10227);
nor U14648 (N_14648,N_8181,N_9462);
xnor U14649 (N_14649,N_9973,N_11839);
nand U14650 (N_14650,N_9795,N_9334);
or U14651 (N_14651,N_9451,N_10181);
nor U14652 (N_14652,N_9749,N_10593);
and U14653 (N_14653,N_11133,N_8309);
xor U14654 (N_14654,N_8748,N_10320);
or U14655 (N_14655,N_9990,N_10920);
or U14656 (N_14656,N_11995,N_9156);
nor U14657 (N_14657,N_11524,N_9061);
nand U14658 (N_14658,N_11576,N_9966);
nand U14659 (N_14659,N_11801,N_9531);
nor U14660 (N_14660,N_10357,N_11681);
nand U14661 (N_14661,N_9025,N_10784);
nor U14662 (N_14662,N_9293,N_8196);
or U14663 (N_14663,N_8591,N_8222);
nand U14664 (N_14664,N_10320,N_9984);
and U14665 (N_14665,N_11082,N_11445);
and U14666 (N_14666,N_8372,N_10754);
nand U14667 (N_14667,N_10255,N_8261);
nor U14668 (N_14668,N_10551,N_11070);
or U14669 (N_14669,N_9597,N_11692);
nand U14670 (N_14670,N_8773,N_11607);
xnor U14671 (N_14671,N_11465,N_11801);
nand U14672 (N_14672,N_9060,N_10112);
and U14673 (N_14673,N_9446,N_10029);
or U14674 (N_14674,N_8279,N_10200);
xor U14675 (N_14675,N_8034,N_11534);
nand U14676 (N_14676,N_10805,N_9673);
nor U14677 (N_14677,N_10315,N_8272);
nand U14678 (N_14678,N_11550,N_8800);
and U14679 (N_14679,N_10779,N_9219);
nand U14680 (N_14680,N_8909,N_8636);
and U14681 (N_14681,N_8521,N_11532);
nor U14682 (N_14682,N_11166,N_10561);
or U14683 (N_14683,N_9051,N_10488);
nand U14684 (N_14684,N_11471,N_8877);
or U14685 (N_14685,N_8312,N_8048);
nand U14686 (N_14686,N_9390,N_9467);
xnor U14687 (N_14687,N_9913,N_10317);
nand U14688 (N_14688,N_9680,N_10973);
or U14689 (N_14689,N_10081,N_11049);
or U14690 (N_14690,N_8612,N_10845);
and U14691 (N_14691,N_11992,N_9888);
nand U14692 (N_14692,N_8152,N_10589);
or U14693 (N_14693,N_8210,N_11637);
xor U14694 (N_14694,N_8286,N_11026);
xnor U14695 (N_14695,N_8884,N_8042);
nor U14696 (N_14696,N_10196,N_10359);
or U14697 (N_14697,N_10359,N_9762);
or U14698 (N_14698,N_10974,N_11629);
or U14699 (N_14699,N_11506,N_9781);
and U14700 (N_14700,N_11302,N_11872);
nand U14701 (N_14701,N_10778,N_8441);
xor U14702 (N_14702,N_10786,N_8905);
nand U14703 (N_14703,N_10327,N_8624);
nor U14704 (N_14704,N_8746,N_9661);
or U14705 (N_14705,N_10549,N_9415);
and U14706 (N_14706,N_11719,N_10036);
nor U14707 (N_14707,N_8346,N_10795);
nor U14708 (N_14708,N_9500,N_10055);
xor U14709 (N_14709,N_10900,N_11786);
and U14710 (N_14710,N_9740,N_11502);
nor U14711 (N_14711,N_11869,N_8221);
or U14712 (N_14712,N_10834,N_8204);
nand U14713 (N_14713,N_8278,N_10943);
nand U14714 (N_14714,N_10528,N_8492);
nand U14715 (N_14715,N_10134,N_9649);
or U14716 (N_14716,N_10890,N_10374);
or U14717 (N_14717,N_11667,N_10562);
nand U14718 (N_14718,N_11331,N_10694);
and U14719 (N_14719,N_8374,N_9897);
or U14720 (N_14720,N_8344,N_8357);
xnor U14721 (N_14721,N_10560,N_10244);
and U14722 (N_14722,N_10235,N_11214);
nor U14723 (N_14723,N_11891,N_9853);
nor U14724 (N_14724,N_10661,N_9695);
nor U14725 (N_14725,N_10797,N_10017);
nand U14726 (N_14726,N_8989,N_9532);
or U14727 (N_14727,N_11777,N_10586);
xnor U14728 (N_14728,N_11483,N_9457);
and U14729 (N_14729,N_10534,N_11224);
xnor U14730 (N_14730,N_10494,N_9855);
nor U14731 (N_14731,N_9904,N_10634);
or U14732 (N_14732,N_10106,N_8339);
and U14733 (N_14733,N_8728,N_10507);
nand U14734 (N_14734,N_10019,N_10637);
or U14735 (N_14735,N_10505,N_10338);
nand U14736 (N_14736,N_8196,N_11770);
and U14737 (N_14737,N_10072,N_11957);
and U14738 (N_14738,N_10136,N_8108);
nand U14739 (N_14739,N_11892,N_8202);
and U14740 (N_14740,N_8102,N_11155);
and U14741 (N_14741,N_11947,N_8387);
and U14742 (N_14742,N_11918,N_10523);
nor U14743 (N_14743,N_9272,N_10622);
nor U14744 (N_14744,N_9876,N_9844);
and U14745 (N_14745,N_9499,N_8164);
or U14746 (N_14746,N_11477,N_8891);
nand U14747 (N_14747,N_11150,N_10225);
nand U14748 (N_14748,N_9124,N_9253);
nor U14749 (N_14749,N_10949,N_10971);
nor U14750 (N_14750,N_10441,N_11096);
or U14751 (N_14751,N_8888,N_8519);
or U14752 (N_14752,N_9281,N_10925);
or U14753 (N_14753,N_10473,N_8818);
nor U14754 (N_14754,N_11279,N_9198);
or U14755 (N_14755,N_8906,N_9857);
and U14756 (N_14756,N_9561,N_11423);
or U14757 (N_14757,N_8325,N_11335);
and U14758 (N_14758,N_8896,N_9660);
or U14759 (N_14759,N_8269,N_11481);
or U14760 (N_14760,N_10941,N_10175);
nand U14761 (N_14761,N_10020,N_11946);
or U14762 (N_14762,N_10128,N_10668);
nand U14763 (N_14763,N_8282,N_8202);
or U14764 (N_14764,N_8963,N_9685);
nor U14765 (N_14765,N_10042,N_9688);
nor U14766 (N_14766,N_10387,N_8203);
or U14767 (N_14767,N_9093,N_8833);
nor U14768 (N_14768,N_10201,N_8010);
and U14769 (N_14769,N_9731,N_10376);
xnor U14770 (N_14770,N_9610,N_10389);
nand U14771 (N_14771,N_9113,N_10980);
or U14772 (N_14772,N_9110,N_9152);
and U14773 (N_14773,N_9789,N_9836);
or U14774 (N_14774,N_9438,N_9684);
nor U14775 (N_14775,N_9840,N_10581);
or U14776 (N_14776,N_8113,N_10349);
and U14777 (N_14777,N_9991,N_11645);
nor U14778 (N_14778,N_11454,N_9460);
nor U14779 (N_14779,N_10172,N_11213);
and U14780 (N_14780,N_8651,N_11079);
and U14781 (N_14781,N_11920,N_8360);
nand U14782 (N_14782,N_11506,N_9164);
nand U14783 (N_14783,N_8600,N_8607);
xnor U14784 (N_14784,N_11961,N_11516);
nand U14785 (N_14785,N_8058,N_8837);
or U14786 (N_14786,N_10249,N_8342);
and U14787 (N_14787,N_9236,N_8860);
xor U14788 (N_14788,N_11147,N_11569);
and U14789 (N_14789,N_10398,N_9459);
or U14790 (N_14790,N_9625,N_9861);
nor U14791 (N_14791,N_8812,N_8497);
or U14792 (N_14792,N_9605,N_8664);
and U14793 (N_14793,N_10757,N_11864);
or U14794 (N_14794,N_11882,N_10627);
or U14795 (N_14795,N_10131,N_8429);
and U14796 (N_14796,N_8301,N_9565);
and U14797 (N_14797,N_11034,N_10360);
nand U14798 (N_14798,N_10564,N_9404);
or U14799 (N_14799,N_9139,N_8949);
xnor U14800 (N_14800,N_9097,N_11120);
and U14801 (N_14801,N_10272,N_11223);
nor U14802 (N_14802,N_11798,N_8271);
or U14803 (N_14803,N_8851,N_9265);
and U14804 (N_14804,N_8463,N_11670);
and U14805 (N_14805,N_8005,N_9387);
and U14806 (N_14806,N_10997,N_10575);
or U14807 (N_14807,N_11845,N_8540);
nand U14808 (N_14808,N_9474,N_10901);
nand U14809 (N_14809,N_8470,N_11351);
nor U14810 (N_14810,N_10741,N_10055);
nor U14811 (N_14811,N_9902,N_9882);
nor U14812 (N_14812,N_8925,N_9147);
nand U14813 (N_14813,N_9120,N_9838);
or U14814 (N_14814,N_9418,N_9110);
xnor U14815 (N_14815,N_8365,N_11853);
nor U14816 (N_14816,N_10493,N_10818);
nor U14817 (N_14817,N_11263,N_9415);
and U14818 (N_14818,N_9160,N_8099);
and U14819 (N_14819,N_9983,N_11646);
nand U14820 (N_14820,N_8876,N_8183);
or U14821 (N_14821,N_10294,N_10008);
and U14822 (N_14822,N_9936,N_11953);
or U14823 (N_14823,N_9938,N_11827);
nand U14824 (N_14824,N_9204,N_10292);
nor U14825 (N_14825,N_10534,N_10993);
nand U14826 (N_14826,N_9135,N_11266);
and U14827 (N_14827,N_11257,N_8577);
or U14828 (N_14828,N_11706,N_10400);
nand U14829 (N_14829,N_10044,N_9110);
nand U14830 (N_14830,N_11291,N_9035);
or U14831 (N_14831,N_8519,N_9916);
or U14832 (N_14832,N_10775,N_11947);
nand U14833 (N_14833,N_8586,N_9910);
nor U14834 (N_14834,N_9818,N_8856);
nand U14835 (N_14835,N_11519,N_10010);
nand U14836 (N_14836,N_10431,N_10691);
xnor U14837 (N_14837,N_11421,N_10228);
nand U14838 (N_14838,N_10957,N_11122);
or U14839 (N_14839,N_10282,N_8081);
nand U14840 (N_14840,N_8068,N_8552);
nand U14841 (N_14841,N_10992,N_10971);
or U14842 (N_14842,N_11373,N_11601);
xor U14843 (N_14843,N_11782,N_8253);
nor U14844 (N_14844,N_11169,N_11162);
nand U14845 (N_14845,N_8972,N_10700);
or U14846 (N_14846,N_8451,N_10510);
xnor U14847 (N_14847,N_10291,N_8458);
xnor U14848 (N_14848,N_11343,N_9052);
and U14849 (N_14849,N_8358,N_10899);
or U14850 (N_14850,N_9186,N_11510);
and U14851 (N_14851,N_10909,N_10224);
or U14852 (N_14852,N_10375,N_11976);
nand U14853 (N_14853,N_11499,N_10323);
or U14854 (N_14854,N_9982,N_10609);
xnor U14855 (N_14855,N_8632,N_11776);
and U14856 (N_14856,N_9418,N_11494);
nand U14857 (N_14857,N_11722,N_9509);
or U14858 (N_14858,N_8334,N_8901);
nand U14859 (N_14859,N_9969,N_8757);
nor U14860 (N_14860,N_8230,N_8877);
and U14861 (N_14861,N_11715,N_9452);
nor U14862 (N_14862,N_11604,N_8058);
nand U14863 (N_14863,N_10853,N_8886);
or U14864 (N_14864,N_9133,N_10775);
nand U14865 (N_14865,N_8699,N_10250);
xor U14866 (N_14866,N_9153,N_8245);
or U14867 (N_14867,N_10907,N_11177);
nor U14868 (N_14868,N_9865,N_9176);
nor U14869 (N_14869,N_10308,N_8380);
or U14870 (N_14870,N_10202,N_11953);
or U14871 (N_14871,N_10417,N_8600);
or U14872 (N_14872,N_11582,N_11776);
nand U14873 (N_14873,N_8992,N_11523);
and U14874 (N_14874,N_11861,N_11403);
nand U14875 (N_14875,N_11776,N_11813);
xnor U14876 (N_14876,N_10960,N_9392);
and U14877 (N_14877,N_9659,N_8971);
nor U14878 (N_14878,N_11355,N_11904);
and U14879 (N_14879,N_9617,N_10759);
xor U14880 (N_14880,N_9311,N_10979);
nand U14881 (N_14881,N_11905,N_10935);
nor U14882 (N_14882,N_8514,N_11340);
or U14883 (N_14883,N_10939,N_8795);
or U14884 (N_14884,N_11928,N_9480);
or U14885 (N_14885,N_8977,N_8806);
xnor U14886 (N_14886,N_10394,N_11271);
or U14887 (N_14887,N_10295,N_9766);
nor U14888 (N_14888,N_10528,N_11155);
nor U14889 (N_14889,N_8091,N_11371);
nand U14890 (N_14890,N_11838,N_11104);
or U14891 (N_14891,N_11027,N_11037);
and U14892 (N_14892,N_8443,N_9893);
nand U14893 (N_14893,N_11714,N_11002);
nand U14894 (N_14894,N_11399,N_11467);
and U14895 (N_14895,N_8580,N_10730);
and U14896 (N_14896,N_10189,N_10104);
nor U14897 (N_14897,N_8252,N_10529);
nor U14898 (N_14898,N_9675,N_8242);
and U14899 (N_14899,N_11462,N_9550);
nand U14900 (N_14900,N_11491,N_9940);
nor U14901 (N_14901,N_9761,N_11355);
or U14902 (N_14902,N_11887,N_9599);
nor U14903 (N_14903,N_8198,N_9119);
nor U14904 (N_14904,N_10345,N_8555);
nand U14905 (N_14905,N_9589,N_9082);
and U14906 (N_14906,N_9013,N_9971);
xnor U14907 (N_14907,N_9336,N_8096);
or U14908 (N_14908,N_8158,N_8777);
or U14909 (N_14909,N_10817,N_8833);
or U14910 (N_14910,N_9808,N_8942);
or U14911 (N_14911,N_9517,N_9197);
and U14912 (N_14912,N_8323,N_10471);
nand U14913 (N_14913,N_9508,N_9872);
and U14914 (N_14914,N_8110,N_9157);
nand U14915 (N_14915,N_10451,N_9770);
or U14916 (N_14916,N_9332,N_10429);
and U14917 (N_14917,N_9199,N_11108);
and U14918 (N_14918,N_10108,N_10584);
nor U14919 (N_14919,N_11867,N_11994);
or U14920 (N_14920,N_8419,N_8713);
and U14921 (N_14921,N_11204,N_11023);
and U14922 (N_14922,N_8880,N_8602);
and U14923 (N_14923,N_8296,N_10755);
nand U14924 (N_14924,N_10339,N_8166);
xor U14925 (N_14925,N_9849,N_10443);
nor U14926 (N_14926,N_8988,N_9169);
or U14927 (N_14927,N_10228,N_8469);
and U14928 (N_14928,N_8710,N_9384);
nand U14929 (N_14929,N_10776,N_8979);
and U14930 (N_14930,N_9910,N_9345);
nor U14931 (N_14931,N_8838,N_9843);
xnor U14932 (N_14932,N_10644,N_10916);
and U14933 (N_14933,N_9966,N_10300);
nor U14934 (N_14934,N_10830,N_11937);
or U14935 (N_14935,N_11517,N_10553);
nor U14936 (N_14936,N_11668,N_11075);
nor U14937 (N_14937,N_8344,N_10932);
or U14938 (N_14938,N_8477,N_11592);
nor U14939 (N_14939,N_9407,N_8559);
and U14940 (N_14940,N_9939,N_11288);
or U14941 (N_14941,N_10123,N_10296);
or U14942 (N_14942,N_10272,N_10940);
nor U14943 (N_14943,N_10800,N_11406);
and U14944 (N_14944,N_9494,N_10176);
or U14945 (N_14945,N_10673,N_10552);
nor U14946 (N_14946,N_8036,N_11784);
nand U14947 (N_14947,N_8313,N_11472);
and U14948 (N_14948,N_11387,N_8814);
or U14949 (N_14949,N_8538,N_9305);
and U14950 (N_14950,N_8013,N_10739);
nand U14951 (N_14951,N_10850,N_9853);
nand U14952 (N_14952,N_10298,N_9422);
xnor U14953 (N_14953,N_11161,N_8811);
nor U14954 (N_14954,N_9967,N_11747);
nor U14955 (N_14955,N_10199,N_11817);
nor U14956 (N_14956,N_10764,N_11337);
nor U14957 (N_14957,N_8391,N_8898);
and U14958 (N_14958,N_9749,N_8441);
and U14959 (N_14959,N_11477,N_11168);
nor U14960 (N_14960,N_10085,N_11581);
nand U14961 (N_14961,N_11221,N_9702);
nor U14962 (N_14962,N_11426,N_10281);
or U14963 (N_14963,N_9724,N_9743);
nor U14964 (N_14964,N_11319,N_11281);
or U14965 (N_14965,N_8768,N_8865);
nand U14966 (N_14966,N_11907,N_10071);
nor U14967 (N_14967,N_10938,N_10183);
or U14968 (N_14968,N_8819,N_8329);
and U14969 (N_14969,N_11610,N_11597);
and U14970 (N_14970,N_10008,N_10627);
and U14971 (N_14971,N_8117,N_8193);
and U14972 (N_14972,N_8770,N_9173);
nor U14973 (N_14973,N_8886,N_8606);
and U14974 (N_14974,N_11019,N_9273);
or U14975 (N_14975,N_10580,N_11659);
or U14976 (N_14976,N_9535,N_10812);
nor U14977 (N_14977,N_10215,N_8851);
nor U14978 (N_14978,N_10551,N_10176);
or U14979 (N_14979,N_8553,N_10609);
nor U14980 (N_14980,N_10147,N_8034);
nor U14981 (N_14981,N_8532,N_11522);
nor U14982 (N_14982,N_8417,N_10183);
or U14983 (N_14983,N_11939,N_10522);
or U14984 (N_14984,N_9850,N_8680);
nor U14985 (N_14985,N_11062,N_11688);
and U14986 (N_14986,N_8802,N_10682);
nand U14987 (N_14987,N_9007,N_9730);
or U14988 (N_14988,N_10920,N_9516);
nand U14989 (N_14989,N_9739,N_11513);
nor U14990 (N_14990,N_9381,N_8099);
xor U14991 (N_14991,N_11052,N_10667);
xnor U14992 (N_14992,N_10978,N_11279);
and U14993 (N_14993,N_9494,N_10458);
nor U14994 (N_14994,N_8336,N_11185);
nand U14995 (N_14995,N_10932,N_11083);
or U14996 (N_14996,N_8096,N_11784);
nor U14997 (N_14997,N_10404,N_11074);
nand U14998 (N_14998,N_8578,N_9662);
or U14999 (N_14999,N_9408,N_8993);
or U15000 (N_15000,N_8543,N_8186);
and U15001 (N_15001,N_8857,N_10020);
nor U15002 (N_15002,N_10074,N_8643);
and U15003 (N_15003,N_9920,N_8716);
and U15004 (N_15004,N_9868,N_11739);
and U15005 (N_15005,N_8746,N_9049);
or U15006 (N_15006,N_11716,N_10753);
or U15007 (N_15007,N_9214,N_8512);
nand U15008 (N_15008,N_8463,N_8340);
or U15009 (N_15009,N_8560,N_9818);
xor U15010 (N_15010,N_11059,N_8550);
nand U15011 (N_15011,N_11827,N_11769);
nor U15012 (N_15012,N_9048,N_10427);
or U15013 (N_15013,N_10911,N_11852);
xnor U15014 (N_15014,N_8607,N_11051);
or U15015 (N_15015,N_9798,N_8537);
nor U15016 (N_15016,N_11495,N_8009);
nor U15017 (N_15017,N_11681,N_8217);
nor U15018 (N_15018,N_10400,N_9487);
or U15019 (N_15019,N_9239,N_9300);
and U15020 (N_15020,N_9697,N_8097);
and U15021 (N_15021,N_10097,N_8048);
and U15022 (N_15022,N_8015,N_11507);
and U15023 (N_15023,N_11942,N_9586);
nand U15024 (N_15024,N_10746,N_10335);
and U15025 (N_15025,N_10782,N_10386);
xnor U15026 (N_15026,N_8131,N_11604);
and U15027 (N_15027,N_10336,N_11951);
nor U15028 (N_15028,N_9825,N_11516);
nor U15029 (N_15029,N_11251,N_9224);
and U15030 (N_15030,N_10444,N_11261);
or U15031 (N_15031,N_10357,N_8197);
or U15032 (N_15032,N_10826,N_11668);
nand U15033 (N_15033,N_8339,N_9057);
nor U15034 (N_15034,N_11614,N_9738);
nand U15035 (N_15035,N_10238,N_8579);
and U15036 (N_15036,N_8239,N_8320);
nand U15037 (N_15037,N_11788,N_11171);
nor U15038 (N_15038,N_11787,N_10008);
or U15039 (N_15039,N_8804,N_10666);
xnor U15040 (N_15040,N_9633,N_9088);
nand U15041 (N_15041,N_11722,N_8619);
xnor U15042 (N_15042,N_10334,N_9981);
nor U15043 (N_15043,N_8102,N_9282);
or U15044 (N_15044,N_10266,N_10678);
nor U15045 (N_15045,N_8912,N_10915);
and U15046 (N_15046,N_9142,N_11352);
nor U15047 (N_15047,N_10316,N_8876);
nor U15048 (N_15048,N_11429,N_9288);
and U15049 (N_15049,N_11522,N_11549);
or U15050 (N_15050,N_9965,N_9964);
and U15051 (N_15051,N_8857,N_9306);
and U15052 (N_15052,N_8518,N_11707);
nor U15053 (N_15053,N_11852,N_11611);
nand U15054 (N_15054,N_9024,N_8144);
xnor U15055 (N_15055,N_8770,N_11828);
nor U15056 (N_15056,N_9868,N_8933);
nor U15057 (N_15057,N_10312,N_8467);
or U15058 (N_15058,N_10754,N_8096);
and U15059 (N_15059,N_9670,N_9625);
nor U15060 (N_15060,N_11498,N_10665);
and U15061 (N_15061,N_10741,N_9468);
nor U15062 (N_15062,N_8320,N_8160);
nand U15063 (N_15063,N_11594,N_10256);
nand U15064 (N_15064,N_10277,N_9399);
nand U15065 (N_15065,N_11547,N_9551);
and U15066 (N_15066,N_8354,N_9308);
and U15067 (N_15067,N_8670,N_9027);
nor U15068 (N_15068,N_9511,N_11900);
xor U15069 (N_15069,N_8507,N_8618);
and U15070 (N_15070,N_9102,N_10614);
or U15071 (N_15071,N_9458,N_8953);
and U15072 (N_15072,N_10798,N_11213);
xnor U15073 (N_15073,N_8924,N_9881);
nor U15074 (N_15074,N_8987,N_9679);
and U15075 (N_15075,N_11698,N_10720);
and U15076 (N_15076,N_10808,N_10409);
and U15077 (N_15077,N_10388,N_11019);
nand U15078 (N_15078,N_9513,N_9580);
xnor U15079 (N_15079,N_8833,N_9435);
and U15080 (N_15080,N_9599,N_8472);
nand U15081 (N_15081,N_9406,N_9435);
or U15082 (N_15082,N_9113,N_10286);
nand U15083 (N_15083,N_8052,N_11947);
nor U15084 (N_15084,N_9879,N_11096);
and U15085 (N_15085,N_8439,N_9993);
nor U15086 (N_15086,N_8435,N_9692);
nor U15087 (N_15087,N_11477,N_11195);
nand U15088 (N_15088,N_8216,N_9509);
nor U15089 (N_15089,N_10203,N_8500);
nand U15090 (N_15090,N_10014,N_8657);
nand U15091 (N_15091,N_10745,N_8345);
nor U15092 (N_15092,N_11575,N_10666);
xor U15093 (N_15093,N_10616,N_9626);
or U15094 (N_15094,N_10288,N_9409);
nor U15095 (N_15095,N_8219,N_10081);
and U15096 (N_15096,N_10038,N_9250);
or U15097 (N_15097,N_10969,N_10387);
nor U15098 (N_15098,N_11338,N_8141);
or U15099 (N_15099,N_11656,N_9896);
xnor U15100 (N_15100,N_8232,N_8120);
and U15101 (N_15101,N_9104,N_11380);
and U15102 (N_15102,N_10527,N_8033);
nor U15103 (N_15103,N_9997,N_9769);
or U15104 (N_15104,N_9991,N_9247);
or U15105 (N_15105,N_11172,N_9795);
xor U15106 (N_15106,N_11509,N_9093);
nand U15107 (N_15107,N_11923,N_10828);
nand U15108 (N_15108,N_9824,N_11034);
and U15109 (N_15109,N_10375,N_10158);
or U15110 (N_15110,N_9467,N_8701);
or U15111 (N_15111,N_11429,N_8844);
and U15112 (N_15112,N_11605,N_9113);
nor U15113 (N_15113,N_8399,N_11490);
or U15114 (N_15114,N_8246,N_10991);
or U15115 (N_15115,N_8557,N_11587);
nand U15116 (N_15116,N_9244,N_10531);
and U15117 (N_15117,N_11667,N_11233);
or U15118 (N_15118,N_9170,N_11626);
or U15119 (N_15119,N_8866,N_9352);
nor U15120 (N_15120,N_11231,N_9528);
nand U15121 (N_15121,N_8653,N_10363);
and U15122 (N_15122,N_9529,N_11601);
nand U15123 (N_15123,N_11164,N_8093);
and U15124 (N_15124,N_9587,N_9077);
nor U15125 (N_15125,N_8418,N_9076);
or U15126 (N_15126,N_9639,N_9155);
and U15127 (N_15127,N_11686,N_11933);
nand U15128 (N_15128,N_8186,N_11103);
nand U15129 (N_15129,N_11454,N_9399);
and U15130 (N_15130,N_8842,N_11272);
or U15131 (N_15131,N_8588,N_11233);
or U15132 (N_15132,N_9401,N_9219);
xor U15133 (N_15133,N_8002,N_8721);
and U15134 (N_15134,N_11108,N_11522);
and U15135 (N_15135,N_8794,N_11016);
xor U15136 (N_15136,N_8430,N_9390);
and U15137 (N_15137,N_8505,N_9337);
and U15138 (N_15138,N_11133,N_9800);
nor U15139 (N_15139,N_10904,N_11328);
or U15140 (N_15140,N_9424,N_8158);
nor U15141 (N_15141,N_11421,N_8127);
nand U15142 (N_15142,N_10473,N_11888);
or U15143 (N_15143,N_9223,N_10741);
and U15144 (N_15144,N_9090,N_11535);
and U15145 (N_15145,N_9669,N_10759);
xor U15146 (N_15146,N_8907,N_8458);
nor U15147 (N_15147,N_9076,N_9420);
nand U15148 (N_15148,N_10815,N_11486);
and U15149 (N_15149,N_10849,N_9193);
or U15150 (N_15150,N_9836,N_10445);
nand U15151 (N_15151,N_11344,N_11357);
or U15152 (N_15152,N_11659,N_8846);
nand U15153 (N_15153,N_9720,N_8518);
nor U15154 (N_15154,N_8069,N_10103);
xnor U15155 (N_15155,N_8475,N_10691);
and U15156 (N_15156,N_11259,N_11585);
nand U15157 (N_15157,N_8346,N_8254);
and U15158 (N_15158,N_10094,N_10017);
nand U15159 (N_15159,N_10726,N_9890);
and U15160 (N_15160,N_10704,N_9075);
nand U15161 (N_15161,N_8185,N_8201);
nor U15162 (N_15162,N_11541,N_10989);
nor U15163 (N_15163,N_11542,N_10963);
nor U15164 (N_15164,N_10390,N_11195);
nand U15165 (N_15165,N_11938,N_8986);
or U15166 (N_15166,N_8885,N_8773);
nor U15167 (N_15167,N_11315,N_11075);
or U15168 (N_15168,N_9917,N_9538);
nor U15169 (N_15169,N_9564,N_8713);
and U15170 (N_15170,N_9354,N_11660);
nor U15171 (N_15171,N_8915,N_11905);
xnor U15172 (N_15172,N_10893,N_11157);
or U15173 (N_15173,N_9840,N_9836);
nand U15174 (N_15174,N_9758,N_9771);
nor U15175 (N_15175,N_11893,N_8635);
or U15176 (N_15176,N_11698,N_9054);
nor U15177 (N_15177,N_8108,N_9595);
or U15178 (N_15178,N_8232,N_9057);
or U15179 (N_15179,N_10245,N_10177);
and U15180 (N_15180,N_8941,N_10081);
nand U15181 (N_15181,N_11905,N_9951);
and U15182 (N_15182,N_9523,N_9110);
nand U15183 (N_15183,N_10527,N_9241);
and U15184 (N_15184,N_11481,N_8705);
nand U15185 (N_15185,N_10914,N_11289);
nand U15186 (N_15186,N_10445,N_8788);
xnor U15187 (N_15187,N_11355,N_8091);
xnor U15188 (N_15188,N_10370,N_8009);
nand U15189 (N_15189,N_8532,N_11445);
or U15190 (N_15190,N_10081,N_10082);
nor U15191 (N_15191,N_8563,N_9576);
or U15192 (N_15192,N_10526,N_11822);
nor U15193 (N_15193,N_8116,N_10227);
nor U15194 (N_15194,N_10319,N_8362);
or U15195 (N_15195,N_8734,N_11229);
nand U15196 (N_15196,N_10374,N_11547);
or U15197 (N_15197,N_9931,N_8870);
or U15198 (N_15198,N_11705,N_11814);
and U15199 (N_15199,N_10414,N_8051);
nor U15200 (N_15200,N_11046,N_10117);
nor U15201 (N_15201,N_9782,N_9481);
xor U15202 (N_15202,N_8825,N_11102);
and U15203 (N_15203,N_8181,N_8551);
and U15204 (N_15204,N_11189,N_9162);
nor U15205 (N_15205,N_10512,N_10160);
xor U15206 (N_15206,N_11859,N_11884);
nor U15207 (N_15207,N_8251,N_8477);
or U15208 (N_15208,N_9741,N_11782);
xor U15209 (N_15209,N_8976,N_9074);
nor U15210 (N_15210,N_8836,N_8753);
and U15211 (N_15211,N_9856,N_9018);
and U15212 (N_15212,N_8224,N_8233);
or U15213 (N_15213,N_11375,N_8605);
and U15214 (N_15214,N_8302,N_9085);
nor U15215 (N_15215,N_10272,N_9881);
nand U15216 (N_15216,N_10798,N_11846);
and U15217 (N_15217,N_9507,N_9569);
nand U15218 (N_15218,N_11811,N_11780);
or U15219 (N_15219,N_8356,N_10850);
or U15220 (N_15220,N_8367,N_8005);
nor U15221 (N_15221,N_9990,N_9317);
and U15222 (N_15222,N_11564,N_11218);
and U15223 (N_15223,N_10930,N_9802);
nand U15224 (N_15224,N_10584,N_11763);
and U15225 (N_15225,N_9362,N_8451);
xnor U15226 (N_15226,N_8208,N_9268);
nor U15227 (N_15227,N_9935,N_10746);
nor U15228 (N_15228,N_9311,N_9208);
xor U15229 (N_15229,N_9960,N_9542);
or U15230 (N_15230,N_11631,N_11316);
nand U15231 (N_15231,N_8120,N_10246);
and U15232 (N_15232,N_11641,N_10738);
and U15233 (N_15233,N_8880,N_10538);
or U15234 (N_15234,N_9007,N_8180);
and U15235 (N_15235,N_8308,N_9192);
or U15236 (N_15236,N_11280,N_8473);
nand U15237 (N_15237,N_8826,N_11968);
nand U15238 (N_15238,N_9509,N_11501);
or U15239 (N_15239,N_11378,N_10820);
and U15240 (N_15240,N_8396,N_10366);
nand U15241 (N_15241,N_9168,N_9372);
and U15242 (N_15242,N_11267,N_11587);
nor U15243 (N_15243,N_8108,N_11159);
xnor U15244 (N_15244,N_9644,N_10150);
nand U15245 (N_15245,N_9249,N_8133);
nand U15246 (N_15246,N_9785,N_8761);
and U15247 (N_15247,N_10661,N_10463);
nand U15248 (N_15248,N_8468,N_8755);
nand U15249 (N_15249,N_11600,N_11248);
or U15250 (N_15250,N_10234,N_10295);
and U15251 (N_15251,N_11255,N_9470);
and U15252 (N_15252,N_10304,N_8481);
nand U15253 (N_15253,N_9991,N_11584);
nor U15254 (N_15254,N_8517,N_8374);
and U15255 (N_15255,N_9341,N_11606);
xor U15256 (N_15256,N_9642,N_11972);
nand U15257 (N_15257,N_11223,N_8262);
nor U15258 (N_15258,N_10227,N_10997);
nand U15259 (N_15259,N_8284,N_10241);
and U15260 (N_15260,N_10978,N_10631);
nand U15261 (N_15261,N_10707,N_8880);
nor U15262 (N_15262,N_11400,N_10643);
nand U15263 (N_15263,N_10939,N_10876);
xor U15264 (N_15264,N_11467,N_9391);
nor U15265 (N_15265,N_9300,N_8646);
nor U15266 (N_15266,N_11780,N_8626);
nor U15267 (N_15267,N_8007,N_9462);
nand U15268 (N_15268,N_9803,N_9980);
xor U15269 (N_15269,N_9435,N_8357);
or U15270 (N_15270,N_11920,N_10960);
nand U15271 (N_15271,N_9442,N_10179);
nor U15272 (N_15272,N_11535,N_10332);
nor U15273 (N_15273,N_9557,N_10828);
or U15274 (N_15274,N_10050,N_8640);
or U15275 (N_15275,N_8299,N_11247);
nor U15276 (N_15276,N_10956,N_10842);
nor U15277 (N_15277,N_10808,N_8934);
nand U15278 (N_15278,N_11288,N_9734);
nand U15279 (N_15279,N_8581,N_10447);
nand U15280 (N_15280,N_10988,N_11305);
and U15281 (N_15281,N_8599,N_9797);
or U15282 (N_15282,N_8922,N_10469);
and U15283 (N_15283,N_11822,N_11387);
xor U15284 (N_15284,N_10310,N_11385);
nand U15285 (N_15285,N_10050,N_11782);
nor U15286 (N_15286,N_8193,N_11378);
or U15287 (N_15287,N_11326,N_8732);
and U15288 (N_15288,N_10420,N_11022);
and U15289 (N_15289,N_8328,N_9044);
nor U15290 (N_15290,N_9201,N_9806);
nand U15291 (N_15291,N_8608,N_10599);
nor U15292 (N_15292,N_10375,N_9021);
nand U15293 (N_15293,N_8372,N_8802);
xor U15294 (N_15294,N_9732,N_9607);
nor U15295 (N_15295,N_8981,N_10784);
xnor U15296 (N_15296,N_8401,N_8658);
nand U15297 (N_15297,N_9750,N_8092);
nand U15298 (N_15298,N_9555,N_10263);
nor U15299 (N_15299,N_11684,N_11159);
and U15300 (N_15300,N_11976,N_8486);
nand U15301 (N_15301,N_9977,N_11984);
and U15302 (N_15302,N_8491,N_8028);
xnor U15303 (N_15303,N_11493,N_11066);
and U15304 (N_15304,N_11025,N_10173);
and U15305 (N_15305,N_8031,N_8914);
and U15306 (N_15306,N_8103,N_8378);
nor U15307 (N_15307,N_9521,N_8804);
nand U15308 (N_15308,N_10071,N_11223);
and U15309 (N_15309,N_11997,N_8466);
nor U15310 (N_15310,N_11814,N_8250);
nand U15311 (N_15311,N_9352,N_9268);
or U15312 (N_15312,N_10724,N_8344);
and U15313 (N_15313,N_10983,N_11528);
nor U15314 (N_15314,N_9591,N_9848);
xnor U15315 (N_15315,N_9777,N_11754);
xor U15316 (N_15316,N_11386,N_8759);
nor U15317 (N_15317,N_11714,N_8067);
nand U15318 (N_15318,N_10650,N_10590);
or U15319 (N_15319,N_10640,N_10215);
or U15320 (N_15320,N_9073,N_9103);
nand U15321 (N_15321,N_8224,N_10511);
nand U15322 (N_15322,N_8692,N_11406);
and U15323 (N_15323,N_10517,N_8066);
nor U15324 (N_15324,N_8477,N_10187);
xor U15325 (N_15325,N_11901,N_9092);
or U15326 (N_15326,N_10419,N_11003);
and U15327 (N_15327,N_8082,N_9521);
xnor U15328 (N_15328,N_10353,N_8918);
and U15329 (N_15329,N_10303,N_10185);
and U15330 (N_15330,N_10519,N_9808);
or U15331 (N_15331,N_9169,N_11898);
nand U15332 (N_15332,N_11893,N_8463);
or U15333 (N_15333,N_10512,N_9404);
xnor U15334 (N_15334,N_8140,N_9481);
and U15335 (N_15335,N_11131,N_9606);
nand U15336 (N_15336,N_8158,N_8590);
and U15337 (N_15337,N_9986,N_8702);
or U15338 (N_15338,N_8848,N_10257);
and U15339 (N_15339,N_8442,N_9801);
and U15340 (N_15340,N_9658,N_8409);
and U15341 (N_15341,N_8835,N_10908);
and U15342 (N_15342,N_9604,N_11179);
nand U15343 (N_15343,N_9629,N_8941);
nor U15344 (N_15344,N_9183,N_10849);
or U15345 (N_15345,N_10615,N_11186);
xor U15346 (N_15346,N_11224,N_9283);
xor U15347 (N_15347,N_9978,N_11811);
nand U15348 (N_15348,N_10619,N_9563);
nor U15349 (N_15349,N_9601,N_9807);
xor U15350 (N_15350,N_8218,N_9144);
and U15351 (N_15351,N_9473,N_8584);
nor U15352 (N_15352,N_10137,N_8468);
or U15353 (N_15353,N_9672,N_10119);
or U15354 (N_15354,N_10543,N_9860);
and U15355 (N_15355,N_8576,N_11120);
and U15356 (N_15356,N_11243,N_8274);
and U15357 (N_15357,N_8020,N_8254);
nor U15358 (N_15358,N_10368,N_8235);
nor U15359 (N_15359,N_8858,N_9015);
and U15360 (N_15360,N_10823,N_9471);
nor U15361 (N_15361,N_11080,N_10916);
and U15362 (N_15362,N_11634,N_8668);
nor U15363 (N_15363,N_9632,N_10913);
nor U15364 (N_15364,N_11632,N_11839);
nand U15365 (N_15365,N_9725,N_8060);
nand U15366 (N_15366,N_8079,N_9394);
nor U15367 (N_15367,N_11697,N_11564);
xor U15368 (N_15368,N_11490,N_11451);
xnor U15369 (N_15369,N_10129,N_11877);
xor U15370 (N_15370,N_11429,N_11403);
xnor U15371 (N_15371,N_9487,N_8241);
or U15372 (N_15372,N_11302,N_8778);
or U15373 (N_15373,N_8787,N_9209);
xnor U15374 (N_15374,N_10133,N_11283);
nor U15375 (N_15375,N_10484,N_11465);
and U15376 (N_15376,N_11750,N_10583);
nor U15377 (N_15377,N_8515,N_8627);
nor U15378 (N_15378,N_8555,N_11130);
and U15379 (N_15379,N_11216,N_10890);
xor U15380 (N_15380,N_9965,N_8239);
nor U15381 (N_15381,N_10273,N_9649);
nor U15382 (N_15382,N_8486,N_9736);
nor U15383 (N_15383,N_10875,N_9872);
nor U15384 (N_15384,N_8413,N_10036);
or U15385 (N_15385,N_10310,N_10889);
and U15386 (N_15386,N_9900,N_9478);
nand U15387 (N_15387,N_10560,N_11080);
or U15388 (N_15388,N_8332,N_11537);
nand U15389 (N_15389,N_8933,N_10980);
nand U15390 (N_15390,N_10046,N_11025);
nor U15391 (N_15391,N_11790,N_8659);
or U15392 (N_15392,N_10535,N_11199);
nand U15393 (N_15393,N_8492,N_8870);
or U15394 (N_15394,N_10264,N_8946);
nand U15395 (N_15395,N_10265,N_10719);
xor U15396 (N_15396,N_8476,N_8676);
or U15397 (N_15397,N_8616,N_8482);
xor U15398 (N_15398,N_8557,N_8031);
and U15399 (N_15399,N_11142,N_8637);
and U15400 (N_15400,N_8084,N_8471);
and U15401 (N_15401,N_9384,N_9479);
nand U15402 (N_15402,N_10815,N_11720);
nor U15403 (N_15403,N_9703,N_9772);
nand U15404 (N_15404,N_10411,N_10245);
or U15405 (N_15405,N_11283,N_8875);
and U15406 (N_15406,N_9705,N_10061);
nand U15407 (N_15407,N_8799,N_11471);
or U15408 (N_15408,N_9738,N_9053);
or U15409 (N_15409,N_11259,N_10758);
nor U15410 (N_15410,N_8603,N_8664);
or U15411 (N_15411,N_10396,N_10279);
nor U15412 (N_15412,N_9200,N_11412);
or U15413 (N_15413,N_11867,N_10889);
nand U15414 (N_15414,N_10977,N_9769);
nor U15415 (N_15415,N_9277,N_8200);
or U15416 (N_15416,N_11581,N_9787);
or U15417 (N_15417,N_10426,N_11127);
nand U15418 (N_15418,N_8691,N_9186);
nand U15419 (N_15419,N_8846,N_9953);
or U15420 (N_15420,N_11907,N_9147);
nand U15421 (N_15421,N_9786,N_10107);
nor U15422 (N_15422,N_11760,N_8084);
nor U15423 (N_15423,N_10820,N_10632);
nand U15424 (N_15424,N_11181,N_8055);
xor U15425 (N_15425,N_8367,N_9865);
nor U15426 (N_15426,N_9103,N_10003);
and U15427 (N_15427,N_10665,N_9779);
nor U15428 (N_15428,N_11011,N_8447);
xnor U15429 (N_15429,N_9879,N_10974);
xnor U15430 (N_15430,N_9687,N_9629);
nand U15431 (N_15431,N_10507,N_8841);
and U15432 (N_15432,N_10886,N_8984);
or U15433 (N_15433,N_11810,N_9254);
or U15434 (N_15434,N_10765,N_10279);
and U15435 (N_15435,N_10769,N_8903);
or U15436 (N_15436,N_10093,N_8449);
nor U15437 (N_15437,N_9559,N_11098);
and U15438 (N_15438,N_8124,N_10280);
or U15439 (N_15439,N_11118,N_10213);
nor U15440 (N_15440,N_10630,N_11710);
xor U15441 (N_15441,N_10760,N_9399);
nand U15442 (N_15442,N_9267,N_9740);
and U15443 (N_15443,N_9925,N_10037);
xor U15444 (N_15444,N_10550,N_10962);
nand U15445 (N_15445,N_10705,N_10431);
nor U15446 (N_15446,N_8320,N_9124);
or U15447 (N_15447,N_10336,N_11848);
xor U15448 (N_15448,N_8063,N_11860);
nor U15449 (N_15449,N_10973,N_8806);
or U15450 (N_15450,N_10457,N_11128);
nor U15451 (N_15451,N_9747,N_8135);
and U15452 (N_15452,N_9288,N_8115);
nor U15453 (N_15453,N_11339,N_9656);
or U15454 (N_15454,N_8704,N_11137);
or U15455 (N_15455,N_11428,N_9491);
and U15456 (N_15456,N_9377,N_11561);
or U15457 (N_15457,N_8883,N_11998);
or U15458 (N_15458,N_9994,N_8127);
nand U15459 (N_15459,N_9515,N_8007);
or U15460 (N_15460,N_11812,N_8843);
nor U15461 (N_15461,N_8038,N_8073);
and U15462 (N_15462,N_11287,N_10338);
nor U15463 (N_15463,N_9921,N_11875);
nand U15464 (N_15464,N_8909,N_9199);
xnor U15465 (N_15465,N_10992,N_10069);
nand U15466 (N_15466,N_10765,N_10398);
nor U15467 (N_15467,N_11246,N_8409);
and U15468 (N_15468,N_8190,N_8750);
nand U15469 (N_15469,N_10527,N_8070);
xnor U15470 (N_15470,N_8242,N_9474);
nor U15471 (N_15471,N_9094,N_11745);
and U15472 (N_15472,N_11313,N_10700);
nor U15473 (N_15473,N_8276,N_10758);
or U15474 (N_15474,N_10023,N_8187);
and U15475 (N_15475,N_8911,N_9045);
or U15476 (N_15476,N_9554,N_10940);
or U15477 (N_15477,N_9986,N_10862);
and U15478 (N_15478,N_8600,N_10695);
or U15479 (N_15479,N_9467,N_9572);
nor U15480 (N_15480,N_11130,N_9943);
and U15481 (N_15481,N_10996,N_10456);
nor U15482 (N_15482,N_9258,N_10435);
nand U15483 (N_15483,N_10510,N_9098);
nor U15484 (N_15484,N_11415,N_8659);
nand U15485 (N_15485,N_8658,N_11952);
nor U15486 (N_15486,N_11511,N_11190);
nor U15487 (N_15487,N_10403,N_9977);
and U15488 (N_15488,N_11208,N_11210);
and U15489 (N_15489,N_10818,N_11889);
nor U15490 (N_15490,N_10374,N_11872);
xor U15491 (N_15491,N_11009,N_8610);
nor U15492 (N_15492,N_8031,N_10926);
or U15493 (N_15493,N_9964,N_11665);
xor U15494 (N_15494,N_10861,N_10506);
or U15495 (N_15495,N_11527,N_11282);
and U15496 (N_15496,N_8603,N_10405);
nor U15497 (N_15497,N_11163,N_10736);
or U15498 (N_15498,N_10405,N_11877);
nand U15499 (N_15499,N_11896,N_10662);
nor U15500 (N_15500,N_9303,N_8919);
xnor U15501 (N_15501,N_11742,N_9397);
nor U15502 (N_15502,N_10010,N_8401);
nand U15503 (N_15503,N_10444,N_8786);
or U15504 (N_15504,N_11012,N_8709);
nor U15505 (N_15505,N_11738,N_11564);
or U15506 (N_15506,N_9554,N_9176);
or U15507 (N_15507,N_11069,N_9716);
and U15508 (N_15508,N_9993,N_8730);
or U15509 (N_15509,N_10082,N_8117);
and U15510 (N_15510,N_9075,N_9462);
or U15511 (N_15511,N_11487,N_8109);
and U15512 (N_15512,N_10575,N_10475);
or U15513 (N_15513,N_11766,N_11271);
xnor U15514 (N_15514,N_10993,N_10791);
or U15515 (N_15515,N_11277,N_10897);
or U15516 (N_15516,N_9606,N_10901);
or U15517 (N_15517,N_9925,N_10337);
and U15518 (N_15518,N_10963,N_8917);
xnor U15519 (N_15519,N_9202,N_11021);
nor U15520 (N_15520,N_9865,N_8704);
nand U15521 (N_15521,N_9973,N_11626);
and U15522 (N_15522,N_10424,N_9330);
nand U15523 (N_15523,N_11945,N_9870);
or U15524 (N_15524,N_11810,N_10979);
xnor U15525 (N_15525,N_11153,N_9427);
and U15526 (N_15526,N_8719,N_9217);
nand U15527 (N_15527,N_8975,N_10623);
nand U15528 (N_15528,N_9609,N_8945);
or U15529 (N_15529,N_8597,N_8712);
nand U15530 (N_15530,N_10701,N_11026);
nor U15531 (N_15531,N_8728,N_10110);
or U15532 (N_15532,N_11571,N_9061);
nor U15533 (N_15533,N_9203,N_8604);
or U15534 (N_15534,N_8510,N_9332);
nor U15535 (N_15535,N_11558,N_8251);
nand U15536 (N_15536,N_8572,N_9252);
nor U15537 (N_15537,N_9234,N_10475);
nand U15538 (N_15538,N_8938,N_9778);
nand U15539 (N_15539,N_9678,N_9615);
or U15540 (N_15540,N_11322,N_9173);
nand U15541 (N_15541,N_8727,N_11843);
nand U15542 (N_15542,N_8085,N_8911);
nor U15543 (N_15543,N_10194,N_9501);
xnor U15544 (N_15544,N_11450,N_9698);
nor U15545 (N_15545,N_9677,N_8828);
and U15546 (N_15546,N_11831,N_8564);
nand U15547 (N_15547,N_9690,N_9658);
and U15548 (N_15548,N_11795,N_10752);
nand U15549 (N_15549,N_10102,N_11811);
and U15550 (N_15550,N_8774,N_11934);
nor U15551 (N_15551,N_11840,N_8815);
nand U15552 (N_15552,N_8576,N_9366);
nand U15553 (N_15553,N_11151,N_8696);
or U15554 (N_15554,N_9668,N_10086);
nand U15555 (N_15555,N_11072,N_9987);
and U15556 (N_15556,N_9652,N_11406);
nor U15557 (N_15557,N_8928,N_10176);
or U15558 (N_15558,N_10143,N_8047);
nor U15559 (N_15559,N_9402,N_9958);
nand U15560 (N_15560,N_11642,N_10668);
nor U15561 (N_15561,N_9964,N_9725);
nor U15562 (N_15562,N_10159,N_9107);
nand U15563 (N_15563,N_9132,N_11860);
and U15564 (N_15564,N_8285,N_11515);
or U15565 (N_15565,N_9014,N_11647);
nand U15566 (N_15566,N_9607,N_8372);
or U15567 (N_15567,N_8852,N_8004);
xnor U15568 (N_15568,N_10814,N_8223);
or U15569 (N_15569,N_8854,N_9844);
nor U15570 (N_15570,N_9223,N_8090);
nor U15571 (N_15571,N_10918,N_8958);
nand U15572 (N_15572,N_10842,N_9442);
or U15573 (N_15573,N_11026,N_8280);
xor U15574 (N_15574,N_11769,N_8098);
and U15575 (N_15575,N_9065,N_9499);
or U15576 (N_15576,N_11060,N_11681);
and U15577 (N_15577,N_11861,N_11827);
and U15578 (N_15578,N_8397,N_11213);
and U15579 (N_15579,N_9477,N_9307);
xnor U15580 (N_15580,N_11557,N_8945);
or U15581 (N_15581,N_10537,N_9190);
or U15582 (N_15582,N_8727,N_8792);
and U15583 (N_15583,N_9500,N_10844);
or U15584 (N_15584,N_11272,N_8315);
nand U15585 (N_15585,N_10928,N_10430);
and U15586 (N_15586,N_8557,N_8336);
nand U15587 (N_15587,N_8499,N_11022);
nand U15588 (N_15588,N_11435,N_8493);
and U15589 (N_15589,N_11877,N_9963);
and U15590 (N_15590,N_9185,N_8787);
or U15591 (N_15591,N_9046,N_9570);
or U15592 (N_15592,N_8757,N_9189);
and U15593 (N_15593,N_11505,N_9364);
nor U15594 (N_15594,N_8566,N_9230);
and U15595 (N_15595,N_8592,N_10632);
or U15596 (N_15596,N_9184,N_9921);
xnor U15597 (N_15597,N_9063,N_11958);
or U15598 (N_15598,N_10257,N_10670);
and U15599 (N_15599,N_8699,N_8223);
or U15600 (N_15600,N_8146,N_11021);
nor U15601 (N_15601,N_8439,N_9138);
nor U15602 (N_15602,N_10284,N_10509);
and U15603 (N_15603,N_11083,N_11352);
xnor U15604 (N_15604,N_10787,N_10057);
nand U15605 (N_15605,N_10219,N_10374);
nand U15606 (N_15606,N_9103,N_8299);
xnor U15607 (N_15607,N_11891,N_9946);
and U15608 (N_15608,N_9624,N_9577);
nand U15609 (N_15609,N_8391,N_11305);
nand U15610 (N_15610,N_9493,N_10166);
or U15611 (N_15611,N_11483,N_11341);
xnor U15612 (N_15612,N_11911,N_10842);
nand U15613 (N_15613,N_11691,N_10949);
nor U15614 (N_15614,N_9029,N_11917);
nand U15615 (N_15615,N_9212,N_9613);
and U15616 (N_15616,N_8265,N_8565);
xnor U15617 (N_15617,N_11940,N_9545);
or U15618 (N_15618,N_10010,N_11321);
or U15619 (N_15619,N_9705,N_10058);
or U15620 (N_15620,N_11652,N_10729);
and U15621 (N_15621,N_9565,N_9176);
nand U15622 (N_15622,N_10778,N_10913);
nor U15623 (N_15623,N_10401,N_9003);
and U15624 (N_15624,N_11011,N_11403);
and U15625 (N_15625,N_8773,N_8242);
or U15626 (N_15626,N_9144,N_8144);
nand U15627 (N_15627,N_9236,N_10978);
nand U15628 (N_15628,N_10808,N_10145);
nor U15629 (N_15629,N_8239,N_10925);
or U15630 (N_15630,N_10288,N_8837);
nand U15631 (N_15631,N_10819,N_8563);
or U15632 (N_15632,N_9878,N_11971);
nand U15633 (N_15633,N_8311,N_9664);
nor U15634 (N_15634,N_10932,N_10405);
nand U15635 (N_15635,N_8856,N_8961);
nand U15636 (N_15636,N_8886,N_9125);
or U15637 (N_15637,N_10034,N_10490);
and U15638 (N_15638,N_9996,N_11557);
nor U15639 (N_15639,N_9819,N_11761);
nand U15640 (N_15640,N_8490,N_11521);
nor U15641 (N_15641,N_9983,N_8916);
nand U15642 (N_15642,N_10649,N_9476);
and U15643 (N_15643,N_8284,N_9736);
or U15644 (N_15644,N_8953,N_8745);
nand U15645 (N_15645,N_9873,N_8139);
nand U15646 (N_15646,N_10209,N_8240);
nor U15647 (N_15647,N_8608,N_10842);
nor U15648 (N_15648,N_11612,N_10735);
and U15649 (N_15649,N_8613,N_10886);
nor U15650 (N_15650,N_10290,N_9100);
nand U15651 (N_15651,N_8488,N_10472);
nor U15652 (N_15652,N_10957,N_8727);
nand U15653 (N_15653,N_11787,N_9470);
xnor U15654 (N_15654,N_9585,N_9191);
or U15655 (N_15655,N_8718,N_9152);
and U15656 (N_15656,N_9658,N_11081);
and U15657 (N_15657,N_9624,N_8828);
and U15658 (N_15658,N_11254,N_9248);
nand U15659 (N_15659,N_9790,N_9499);
nand U15660 (N_15660,N_10277,N_10228);
or U15661 (N_15661,N_8090,N_11442);
or U15662 (N_15662,N_9556,N_11861);
nor U15663 (N_15663,N_10508,N_10308);
or U15664 (N_15664,N_11551,N_8473);
and U15665 (N_15665,N_10943,N_10391);
and U15666 (N_15666,N_11323,N_10915);
nand U15667 (N_15667,N_11815,N_8441);
nor U15668 (N_15668,N_10368,N_8718);
or U15669 (N_15669,N_10956,N_9780);
nand U15670 (N_15670,N_11372,N_10566);
and U15671 (N_15671,N_11630,N_11968);
or U15672 (N_15672,N_10472,N_10087);
xor U15673 (N_15673,N_8872,N_10888);
or U15674 (N_15674,N_11814,N_10957);
xnor U15675 (N_15675,N_11998,N_11481);
nor U15676 (N_15676,N_11253,N_11315);
or U15677 (N_15677,N_9676,N_11123);
and U15678 (N_15678,N_10731,N_8882);
nor U15679 (N_15679,N_8948,N_10883);
and U15680 (N_15680,N_8030,N_10619);
or U15681 (N_15681,N_9007,N_11605);
nor U15682 (N_15682,N_11669,N_9502);
nand U15683 (N_15683,N_8959,N_10185);
or U15684 (N_15684,N_9150,N_11897);
nor U15685 (N_15685,N_11906,N_8397);
nor U15686 (N_15686,N_9790,N_10419);
or U15687 (N_15687,N_11027,N_9072);
xnor U15688 (N_15688,N_8104,N_8227);
or U15689 (N_15689,N_11461,N_10925);
nand U15690 (N_15690,N_8159,N_8716);
nor U15691 (N_15691,N_11885,N_11553);
and U15692 (N_15692,N_9548,N_10026);
nand U15693 (N_15693,N_8981,N_10270);
and U15694 (N_15694,N_11572,N_9077);
nor U15695 (N_15695,N_8397,N_8759);
or U15696 (N_15696,N_11217,N_8901);
nand U15697 (N_15697,N_9198,N_9441);
xor U15698 (N_15698,N_10939,N_9606);
nor U15699 (N_15699,N_10545,N_8265);
nand U15700 (N_15700,N_10255,N_8626);
nand U15701 (N_15701,N_11433,N_8413);
nand U15702 (N_15702,N_8392,N_9880);
and U15703 (N_15703,N_8561,N_8671);
xor U15704 (N_15704,N_9149,N_10115);
xor U15705 (N_15705,N_11811,N_8478);
nand U15706 (N_15706,N_10104,N_8195);
or U15707 (N_15707,N_11037,N_9308);
nand U15708 (N_15708,N_9928,N_9839);
xor U15709 (N_15709,N_9708,N_11021);
or U15710 (N_15710,N_11483,N_8679);
or U15711 (N_15711,N_9948,N_11954);
or U15712 (N_15712,N_9548,N_8711);
nor U15713 (N_15713,N_8618,N_9031);
nand U15714 (N_15714,N_10703,N_11308);
nor U15715 (N_15715,N_11195,N_10432);
or U15716 (N_15716,N_8443,N_8766);
and U15717 (N_15717,N_9359,N_10863);
nor U15718 (N_15718,N_8395,N_10820);
and U15719 (N_15719,N_10771,N_11349);
nand U15720 (N_15720,N_10299,N_11452);
or U15721 (N_15721,N_10910,N_11638);
and U15722 (N_15722,N_8161,N_10517);
nor U15723 (N_15723,N_11325,N_10340);
nor U15724 (N_15724,N_8600,N_8659);
and U15725 (N_15725,N_10061,N_10336);
and U15726 (N_15726,N_9197,N_10809);
nor U15727 (N_15727,N_11808,N_8282);
nor U15728 (N_15728,N_8355,N_8417);
and U15729 (N_15729,N_8249,N_11415);
nand U15730 (N_15730,N_10223,N_11218);
and U15731 (N_15731,N_10719,N_11506);
nand U15732 (N_15732,N_10769,N_11210);
or U15733 (N_15733,N_9385,N_8236);
and U15734 (N_15734,N_9849,N_9449);
nand U15735 (N_15735,N_10170,N_10400);
nand U15736 (N_15736,N_11402,N_9807);
or U15737 (N_15737,N_10318,N_10619);
and U15738 (N_15738,N_10216,N_11392);
or U15739 (N_15739,N_11414,N_11094);
xnor U15740 (N_15740,N_10966,N_11595);
or U15741 (N_15741,N_8714,N_10023);
xnor U15742 (N_15742,N_8114,N_9888);
or U15743 (N_15743,N_9721,N_9405);
xnor U15744 (N_15744,N_11090,N_11515);
and U15745 (N_15745,N_8901,N_10674);
and U15746 (N_15746,N_8456,N_11396);
or U15747 (N_15747,N_10016,N_9687);
and U15748 (N_15748,N_9518,N_11832);
xor U15749 (N_15749,N_10614,N_11465);
and U15750 (N_15750,N_11689,N_9102);
and U15751 (N_15751,N_11466,N_9513);
and U15752 (N_15752,N_8904,N_9710);
or U15753 (N_15753,N_11914,N_10374);
nand U15754 (N_15754,N_8503,N_11786);
xor U15755 (N_15755,N_11640,N_8635);
xor U15756 (N_15756,N_11837,N_11956);
nor U15757 (N_15757,N_10696,N_8224);
nand U15758 (N_15758,N_10012,N_10988);
and U15759 (N_15759,N_11539,N_11227);
or U15760 (N_15760,N_11796,N_11137);
and U15761 (N_15761,N_8961,N_8441);
or U15762 (N_15762,N_8471,N_8792);
nor U15763 (N_15763,N_8291,N_10319);
nand U15764 (N_15764,N_11389,N_10695);
nand U15765 (N_15765,N_10880,N_10316);
nand U15766 (N_15766,N_10076,N_8212);
nand U15767 (N_15767,N_11098,N_10315);
and U15768 (N_15768,N_11094,N_10886);
and U15769 (N_15769,N_9723,N_8224);
nand U15770 (N_15770,N_9757,N_9035);
nand U15771 (N_15771,N_10644,N_8637);
xnor U15772 (N_15772,N_10041,N_8410);
and U15773 (N_15773,N_9998,N_10636);
nor U15774 (N_15774,N_9561,N_9805);
and U15775 (N_15775,N_10746,N_10336);
nor U15776 (N_15776,N_11979,N_11074);
xor U15777 (N_15777,N_8543,N_10304);
nand U15778 (N_15778,N_8698,N_10849);
or U15779 (N_15779,N_8197,N_10403);
xor U15780 (N_15780,N_10017,N_10728);
nor U15781 (N_15781,N_8671,N_11702);
nand U15782 (N_15782,N_9543,N_10760);
nor U15783 (N_15783,N_10665,N_10153);
nand U15784 (N_15784,N_9328,N_10902);
and U15785 (N_15785,N_11568,N_11938);
nor U15786 (N_15786,N_8814,N_9717);
nor U15787 (N_15787,N_9644,N_9514);
nand U15788 (N_15788,N_11765,N_8882);
nand U15789 (N_15789,N_9438,N_10956);
and U15790 (N_15790,N_9609,N_11302);
or U15791 (N_15791,N_11687,N_11051);
or U15792 (N_15792,N_9507,N_9695);
nand U15793 (N_15793,N_11485,N_10449);
and U15794 (N_15794,N_11563,N_9661);
and U15795 (N_15795,N_10671,N_8574);
nor U15796 (N_15796,N_11408,N_9173);
nand U15797 (N_15797,N_10878,N_11876);
and U15798 (N_15798,N_9016,N_10655);
nand U15799 (N_15799,N_9861,N_11390);
or U15800 (N_15800,N_10806,N_8020);
nand U15801 (N_15801,N_10702,N_8395);
nand U15802 (N_15802,N_8243,N_8319);
or U15803 (N_15803,N_9752,N_8202);
and U15804 (N_15804,N_10120,N_9242);
nor U15805 (N_15805,N_8280,N_10642);
nor U15806 (N_15806,N_9210,N_10564);
nand U15807 (N_15807,N_11906,N_8727);
nand U15808 (N_15808,N_8019,N_10107);
xnor U15809 (N_15809,N_10014,N_10337);
nor U15810 (N_15810,N_11386,N_11713);
nor U15811 (N_15811,N_9735,N_9444);
nand U15812 (N_15812,N_10024,N_11268);
nor U15813 (N_15813,N_9688,N_10720);
or U15814 (N_15814,N_11192,N_9356);
and U15815 (N_15815,N_9660,N_8091);
nand U15816 (N_15816,N_11567,N_8302);
nand U15817 (N_15817,N_10397,N_8097);
nand U15818 (N_15818,N_10640,N_11200);
or U15819 (N_15819,N_8891,N_9600);
nor U15820 (N_15820,N_9742,N_10084);
or U15821 (N_15821,N_9237,N_9553);
or U15822 (N_15822,N_11174,N_11258);
or U15823 (N_15823,N_8200,N_8877);
nand U15824 (N_15824,N_10239,N_9487);
and U15825 (N_15825,N_11212,N_9497);
nor U15826 (N_15826,N_9111,N_11653);
nand U15827 (N_15827,N_8971,N_9653);
and U15828 (N_15828,N_11330,N_9901);
xnor U15829 (N_15829,N_9520,N_9144);
nand U15830 (N_15830,N_10779,N_10887);
or U15831 (N_15831,N_11613,N_9187);
nand U15832 (N_15832,N_9770,N_8031);
xor U15833 (N_15833,N_10832,N_8893);
nand U15834 (N_15834,N_9684,N_8450);
nand U15835 (N_15835,N_9748,N_10207);
nor U15836 (N_15836,N_11389,N_9457);
and U15837 (N_15837,N_10856,N_11491);
and U15838 (N_15838,N_9512,N_10945);
nand U15839 (N_15839,N_11548,N_10945);
xnor U15840 (N_15840,N_8809,N_10698);
and U15841 (N_15841,N_9076,N_9594);
nand U15842 (N_15842,N_8109,N_10977);
and U15843 (N_15843,N_11089,N_8352);
or U15844 (N_15844,N_11495,N_9534);
nor U15845 (N_15845,N_8279,N_9279);
or U15846 (N_15846,N_10328,N_9545);
and U15847 (N_15847,N_8364,N_11713);
and U15848 (N_15848,N_10155,N_10791);
nor U15849 (N_15849,N_9441,N_11889);
and U15850 (N_15850,N_8112,N_10033);
or U15851 (N_15851,N_9779,N_8735);
and U15852 (N_15852,N_11123,N_9452);
xor U15853 (N_15853,N_9208,N_9275);
xor U15854 (N_15854,N_8515,N_8409);
xor U15855 (N_15855,N_10288,N_8476);
or U15856 (N_15856,N_8712,N_10688);
or U15857 (N_15857,N_9156,N_11110);
nor U15858 (N_15858,N_11557,N_8892);
and U15859 (N_15859,N_8844,N_9054);
or U15860 (N_15860,N_9721,N_8493);
nor U15861 (N_15861,N_8023,N_11872);
nand U15862 (N_15862,N_8867,N_9014);
nand U15863 (N_15863,N_11075,N_10941);
xor U15864 (N_15864,N_9800,N_8608);
nand U15865 (N_15865,N_9549,N_9288);
nor U15866 (N_15866,N_10100,N_11135);
or U15867 (N_15867,N_11245,N_8905);
or U15868 (N_15868,N_11899,N_11731);
or U15869 (N_15869,N_8276,N_10733);
or U15870 (N_15870,N_10150,N_9243);
nor U15871 (N_15871,N_10645,N_8730);
or U15872 (N_15872,N_8816,N_11654);
or U15873 (N_15873,N_8797,N_11270);
nand U15874 (N_15874,N_11491,N_10992);
and U15875 (N_15875,N_10741,N_9174);
nor U15876 (N_15876,N_9281,N_8584);
xnor U15877 (N_15877,N_10074,N_8152);
or U15878 (N_15878,N_8976,N_9077);
nor U15879 (N_15879,N_10923,N_10746);
or U15880 (N_15880,N_11047,N_8801);
nand U15881 (N_15881,N_11778,N_10787);
and U15882 (N_15882,N_11006,N_11587);
nand U15883 (N_15883,N_9703,N_9575);
nor U15884 (N_15884,N_9304,N_11772);
or U15885 (N_15885,N_11342,N_8604);
or U15886 (N_15886,N_11326,N_9903);
xor U15887 (N_15887,N_10686,N_8837);
and U15888 (N_15888,N_11373,N_10289);
and U15889 (N_15889,N_10478,N_11427);
or U15890 (N_15890,N_11805,N_9716);
nand U15891 (N_15891,N_11032,N_9703);
nor U15892 (N_15892,N_9295,N_10342);
nor U15893 (N_15893,N_11488,N_9433);
or U15894 (N_15894,N_8245,N_9488);
xnor U15895 (N_15895,N_8335,N_8272);
xnor U15896 (N_15896,N_9231,N_11786);
and U15897 (N_15897,N_8457,N_10463);
or U15898 (N_15898,N_8808,N_8660);
nor U15899 (N_15899,N_11039,N_11368);
nor U15900 (N_15900,N_8468,N_11071);
nor U15901 (N_15901,N_9198,N_8592);
xnor U15902 (N_15902,N_11110,N_11671);
or U15903 (N_15903,N_11203,N_9574);
nand U15904 (N_15904,N_10959,N_9269);
nand U15905 (N_15905,N_8393,N_9942);
nor U15906 (N_15906,N_10285,N_9075);
or U15907 (N_15907,N_9797,N_9987);
nor U15908 (N_15908,N_9286,N_11588);
and U15909 (N_15909,N_10695,N_11312);
nor U15910 (N_15910,N_11509,N_11294);
nand U15911 (N_15911,N_10754,N_10729);
and U15912 (N_15912,N_8076,N_11384);
nor U15913 (N_15913,N_11774,N_8856);
and U15914 (N_15914,N_8784,N_8474);
nand U15915 (N_15915,N_10699,N_8714);
xnor U15916 (N_15916,N_8455,N_11611);
nor U15917 (N_15917,N_11014,N_8469);
nor U15918 (N_15918,N_10064,N_11706);
or U15919 (N_15919,N_10137,N_11617);
or U15920 (N_15920,N_11267,N_8919);
or U15921 (N_15921,N_10526,N_8197);
and U15922 (N_15922,N_9082,N_9669);
and U15923 (N_15923,N_8009,N_9098);
nand U15924 (N_15924,N_8745,N_8190);
or U15925 (N_15925,N_10699,N_8327);
or U15926 (N_15926,N_11474,N_9672);
nand U15927 (N_15927,N_8190,N_9259);
nor U15928 (N_15928,N_10525,N_10700);
xnor U15929 (N_15929,N_8524,N_10251);
nand U15930 (N_15930,N_11931,N_11570);
or U15931 (N_15931,N_8730,N_9864);
nor U15932 (N_15932,N_10606,N_10579);
xnor U15933 (N_15933,N_10008,N_11729);
nand U15934 (N_15934,N_11923,N_9371);
xnor U15935 (N_15935,N_8294,N_10116);
and U15936 (N_15936,N_11210,N_8674);
nand U15937 (N_15937,N_8900,N_9491);
or U15938 (N_15938,N_11537,N_10193);
xnor U15939 (N_15939,N_10861,N_8765);
and U15940 (N_15940,N_10135,N_8631);
or U15941 (N_15941,N_8349,N_8880);
or U15942 (N_15942,N_10761,N_11997);
or U15943 (N_15943,N_8152,N_10430);
xnor U15944 (N_15944,N_11803,N_10066);
and U15945 (N_15945,N_11523,N_9722);
nor U15946 (N_15946,N_11411,N_8695);
nor U15947 (N_15947,N_8774,N_10797);
nor U15948 (N_15948,N_8688,N_9606);
xnor U15949 (N_15949,N_11635,N_9784);
nor U15950 (N_15950,N_10442,N_10804);
and U15951 (N_15951,N_11677,N_10846);
nand U15952 (N_15952,N_11993,N_9917);
nand U15953 (N_15953,N_9081,N_11307);
nand U15954 (N_15954,N_10311,N_11395);
nand U15955 (N_15955,N_10557,N_8851);
nand U15956 (N_15956,N_11134,N_8449);
nor U15957 (N_15957,N_8083,N_10636);
nand U15958 (N_15958,N_9197,N_9964);
nand U15959 (N_15959,N_8436,N_10686);
nand U15960 (N_15960,N_11467,N_8691);
xor U15961 (N_15961,N_11865,N_8339);
or U15962 (N_15962,N_9616,N_8533);
or U15963 (N_15963,N_9116,N_10574);
and U15964 (N_15964,N_8483,N_10442);
xnor U15965 (N_15965,N_9249,N_8309);
or U15966 (N_15966,N_11350,N_8434);
and U15967 (N_15967,N_11152,N_10822);
nand U15968 (N_15968,N_8462,N_8198);
nor U15969 (N_15969,N_9473,N_10861);
or U15970 (N_15970,N_11863,N_9462);
xor U15971 (N_15971,N_9426,N_8483);
or U15972 (N_15972,N_9770,N_9988);
nand U15973 (N_15973,N_10224,N_10340);
xor U15974 (N_15974,N_11471,N_10493);
and U15975 (N_15975,N_9204,N_10736);
nor U15976 (N_15976,N_10442,N_10058);
nor U15977 (N_15977,N_10293,N_8606);
and U15978 (N_15978,N_11363,N_9386);
or U15979 (N_15979,N_11633,N_9188);
or U15980 (N_15980,N_9611,N_10207);
nand U15981 (N_15981,N_10831,N_10366);
nand U15982 (N_15982,N_10557,N_9484);
nand U15983 (N_15983,N_9091,N_10648);
and U15984 (N_15984,N_9011,N_8822);
or U15985 (N_15985,N_9079,N_10722);
xor U15986 (N_15986,N_11165,N_11670);
and U15987 (N_15987,N_10035,N_9413);
nor U15988 (N_15988,N_10389,N_10375);
nand U15989 (N_15989,N_11009,N_8349);
nor U15990 (N_15990,N_11209,N_10906);
or U15991 (N_15991,N_9270,N_9475);
xnor U15992 (N_15992,N_9398,N_8815);
and U15993 (N_15993,N_8826,N_8709);
nor U15994 (N_15994,N_11710,N_10908);
nor U15995 (N_15995,N_8499,N_11373);
and U15996 (N_15996,N_10158,N_9439);
or U15997 (N_15997,N_8140,N_9304);
and U15998 (N_15998,N_10801,N_9603);
nor U15999 (N_15999,N_10216,N_9524);
nand U16000 (N_16000,N_14362,N_15916);
and U16001 (N_16001,N_15603,N_15817);
nand U16002 (N_16002,N_13293,N_12311);
nor U16003 (N_16003,N_12651,N_12848);
or U16004 (N_16004,N_14083,N_13491);
nand U16005 (N_16005,N_13947,N_12939);
and U16006 (N_16006,N_14770,N_12202);
nor U16007 (N_16007,N_14012,N_12199);
nor U16008 (N_16008,N_14884,N_14729);
or U16009 (N_16009,N_12921,N_12302);
nor U16010 (N_16010,N_15542,N_13239);
xnor U16011 (N_16011,N_13722,N_12523);
nand U16012 (N_16012,N_14368,N_14399);
nor U16013 (N_16013,N_14065,N_15952);
xor U16014 (N_16014,N_15708,N_14206);
nand U16015 (N_16015,N_14375,N_15528);
nand U16016 (N_16016,N_14601,N_13974);
nand U16017 (N_16017,N_12804,N_12639);
xor U16018 (N_16018,N_14158,N_12935);
and U16019 (N_16019,N_14181,N_15811);
xor U16020 (N_16020,N_12173,N_12235);
and U16021 (N_16021,N_13814,N_13210);
xnor U16022 (N_16022,N_13318,N_13826);
nand U16023 (N_16023,N_12405,N_15631);
nor U16024 (N_16024,N_13460,N_13070);
and U16025 (N_16025,N_12113,N_13767);
nor U16026 (N_16026,N_14221,N_12619);
xnor U16027 (N_16027,N_13436,N_13801);
or U16028 (N_16028,N_14632,N_12197);
or U16029 (N_16029,N_14283,N_13909);
or U16030 (N_16030,N_13805,N_15043);
or U16031 (N_16031,N_15187,N_13457);
xor U16032 (N_16032,N_15608,N_14483);
nand U16033 (N_16033,N_12415,N_13168);
and U16034 (N_16034,N_15490,N_13228);
xor U16035 (N_16035,N_15024,N_13453);
nor U16036 (N_16036,N_14517,N_15977);
nor U16037 (N_16037,N_15832,N_15077);
nand U16038 (N_16038,N_15264,N_15706);
nor U16039 (N_16039,N_15434,N_15257);
nand U16040 (N_16040,N_13887,N_13363);
or U16041 (N_16041,N_12857,N_14702);
nor U16042 (N_16042,N_13764,N_14124);
nand U16043 (N_16043,N_15173,N_13047);
nand U16044 (N_16044,N_13308,N_14244);
nand U16045 (N_16045,N_14230,N_15272);
or U16046 (N_16046,N_12563,N_12350);
and U16047 (N_16047,N_15580,N_12386);
nor U16048 (N_16048,N_13594,N_12986);
nor U16049 (N_16049,N_15109,N_15871);
and U16050 (N_16050,N_15049,N_15632);
nand U16051 (N_16051,N_14425,N_14552);
and U16052 (N_16052,N_15932,N_13451);
xnor U16053 (N_16053,N_12275,N_15888);
or U16054 (N_16054,N_13096,N_14280);
nand U16055 (N_16055,N_14306,N_12205);
nand U16056 (N_16056,N_13093,N_13086);
and U16057 (N_16057,N_14711,N_14655);
or U16058 (N_16058,N_12352,N_13470);
xor U16059 (N_16059,N_15305,N_15941);
nand U16060 (N_16060,N_12474,N_14153);
and U16061 (N_16061,N_13265,N_13721);
nor U16062 (N_16062,N_14423,N_15254);
nand U16063 (N_16063,N_12014,N_14037);
or U16064 (N_16064,N_12198,N_14551);
or U16065 (N_16065,N_14363,N_12347);
and U16066 (N_16066,N_12394,N_13654);
or U16067 (N_16067,N_12642,N_12375);
nor U16068 (N_16068,N_13343,N_14851);
nor U16069 (N_16069,N_12504,N_13957);
and U16070 (N_16070,N_12367,N_14698);
or U16071 (N_16071,N_14993,N_12750);
and U16072 (N_16072,N_15799,N_14455);
and U16073 (N_16073,N_13071,N_12254);
and U16074 (N_16074,N_13135,N_13568);
or U16075 (N_16075,N_12952,N_15126);
or U16076 (N_16076,N_14695,N_14835);
xnor U16077 (N_16077,N_14373,N_15050);
nand U16078 (N_16078,N_12053,N_15219);
or U16079 (N_16079,N_13632,N_15802);
xnor U16080 (N_16080,N_15336,N_13283);
nor U16081 (N_16081,N_12412,N_14670);
nor U16082 (N_16082,N_12892,N_13400);
nand U16083 (N_16083,N_15467,N_14262);
xor U16084 (N_16084,N_14001,N_15710);
nor U16085 (N_16085,N_14496,N_13307);
nor U16086 (N_16086,N_15395,N_12627);
xnor U16087 (N_16087,N_14449,N_14417);
nor U16088 (N_16088,N_15124,N_13324);
nor U16089 (N_16089,N_13083,N_14047);
nor U16090 (N_16090,N_15876,N_15172);
nand U16091 (N_16091,N_12353,N_14328);
nor U16092 (N_16092,N_15521,N_15170);
or U16093 (N_16093,N_15056,N_12344);
nand U16094 (N_16094,N_15990,N_15839);
and U16095 (N_16095,N_12381,N_15202);
and U16096 (N_16096,N_15954,N_13510);
nor U16097 (N_16097,N_12324,N_14934);
nor U16098 (N_16098,N_15934,N_12150);
or U16099 (N_16099,N_15252,N_12900);
nand U16100 (N_16100,N_13976,N_12989);
or U16101 (N_16101,N_12182,N_13884);
nor U16102 (N_16102,N_13671,N_15098);
and U16103 (N_16103,N_14808,N_13028);
and U16104 (N_16104,N_13745,N_14218);
nand U16105 (N_16105,N_15984,N_13389);
or U16106 (N_16106,N_13301,N_15999);
xor U16107 (N_16107,N_13736,N_12169);
and U16108 (N_16108,N_12317,N_15074);
or U16109 (N_16109,N_12835,N_14506);
xor U16110 (N_16110,N_14612,N_13647);
nand U16111 (N_16111,N_15496,N_12700);
and U16112 (N_16112,N_14853,N_13998);
or U16113 (N_16113,N_15417,N_15776);
and U16114 (N_16114,N_15825,N_15551);
or U16115 (N_16115,N_12822,N_12458);
or U16116 (N_16116,N_12409,N_12468);
nand U16117 (N_16117,N_12707,N_15891);
and U16118 (N_16118,N_15860,N_15095);
nor U16119 (N_16119,N_15849,N_14329);
or U16120 (N_16120,N_12723,N_15485);
nand U16121 (N_16121,N_12300,N_12692);
nand U16122 (N_16122,N_12897,N_15645);
nor U16123 (N_16123,N_12784,N_15287);
or U16124 (N_16124,N_12508,N_15457);
and U16125 (N_16125,N_14849,N_14560);
or U16126 (N_16126,N_13178,N_14164);
or U16127 (N_16127,N_13375,N_15728);
and U16128 (N_16128,N_15499,N_14769);
nand U16129 (N_16129,N_12288,N_15174);
or U16130 (N_16130,N_14205,N_13452);
or U16131 (N_16131,N_12759,N_12237);
nand U16132 (N_16132,N_15230,N_14875);
nand U16133 (N_16133,N_14666,N_14928);
and U16134 (N_16134,N_14340,N_14510);
and U16135 (N_16135,N_15694,N_12511);
and U16136 (N_16136,N_13734,N_14672);
or U16137 (N_16137,N_12719,N_14296);
and U16138 (N_16138,N_12355,N_12172);
or U16139 (N_16139,N_14781,N_13134);
and U16140 (N_16140,N_12851,N_14173);
nor U16141 (N_16141,N_12956,N_15851);
nand U16142 (N_16142,N_15702,N_14051);
nor U16143 (N_16143,N_15899,N_14997);
xnor U16144 (N_16144,N_15514,N_14028);
nor U16145 (N_16145,N_15415,N_15732);
nor U16146 (N_16146,N_15620,N_14841);
nand U16147 (N_16147,N_14401,N_12282);
or U16148 (N_16148,N_13876,N_12675);
xnor U16149 (N_16149,N_14624,N_13298);
and U16150 (N_16150,N_14380,N_13030);
xor U16151 (N_16151,N_12085,N_13468);
and U16152 (N_16152,N_14342,N_13098);
and U16153 (N_16153,N_15391,N_12534);
and U16154 (N_16154,N_14305,N_15923);
or U16155 (N_16155,N_12180,N_12365);
and U16156 (N_16156,N_14764,N_13089);
or U16157 (N_16157,N_14241,N_13497);
nor U16158 (N_16158,N_12633,N_12335);
nor U16159 (N_16159,N_12208,N_15800);
and U16160 (N_16160,N_15628,N_12343);
nor U16161 (N_16161,N_13760,N_15016);
or U16162 (N_16162,N_14169,N_13675);
or U16163 (N_16163,N_14656,N_14099);
or U16164 (N_16164,N_15078,N_14822);
nand U16165 (N_16165,N_15365,N_12859);
nand U16166 (N_16166,N_15648,N_13322);
nor U16167 (N_16167,N_14383,N_14029);
nand U16168 (N_16168,N_12338,N_13713);
or U16169 (N_16169,N_13459,N_13575);
nor U16170 (N_16170,N_15427,N_15707);
nor U16171 (N_16171,N_15379,N_14319);
nor U16172 (N_16172,N_15213,N_15418);
nor U16173 (N_16173,N_15502,N_13182);
nand U16174 (N_16174,N_15668,N_14093);
and U16175 (N_16175,N_13190,N_15053);
xnor U16176 (N_16176,N_15764,N_13592);
and U16177 (N_16177,N_12366,N_15903);
or U16178 (N_16178,N_13469,N_14662);
or U16179 (N_16179,N_13427,N_12230);
nand U16180 (N_16180,N_13062,N_13603);
xor U16181 (N_16181,N_12506,N_13292);
or U16182 (N_16182,N_13549,N_15150);
nand U16183 (N_16183,N_14497,N_15048);
nand U16184 (N_16184,N_14701,N_15890);
nor U16185 (N_16185,N_14238,N_14035);
or U16186 (N_16186,N_13320,N_14416);
nand U16187 (N_16187,N_13938,N_12397);
and U16188 (N_16188,N_14141,N_14617);
xor U16189 (N_16189,N_13751,N_13091);
or U16190 (N_16190,N_14457,N_12837);
nor U16191 (N_16191,N_13838,N_15996);
and U16192 (N_16192,N_14436,N_12466);
xnor U16193 (N_16193,N_14405,N_15303);
nor U16194 (N_16194,N_15870,N_14864);
nor U16195 (N_16195,N_12874,N_14160);
or U16196 (N_16196,N_13445,N_15279);
and U16197 (N_16197,N_14253,N_12174);
nor U16198 (N_16198,N_15037,N_15138);
nand U16199 (N_16199,N_12864,N_15614);
nor U16200 (N_16200,N_14795,N_15674);
or U16201 (N_16201,N_14117,N_13865);
and U16202 (N_16202,N_13197,N_13414);
nor U16203 (N_16203,N_12153,N_12994);
and U16204 (N_16204,N_14608,N_14650);
xor U16205 (N_16205,N_13153,N_15667);
or U16206 (N_16206,N_14390,N_14096);
nand U16207 (N_16207,N_14235,N_13765);
nor U16208 (N_16208,N_15167,N_12188);
and U16209 (N_16209,N_12801,N_13822);
or U16210 (N_16210,N_12682,N_15258);
and U16211 (N_16211,N_12094,N_13705);
or U16212 (N_16212,N_12330,N_12727);
or U16213 (N_16213,N_13557,N_14988);
nand U16214 (N_16214,N_13063,N_13779);
and U16215 (N_16215,N_14842,N_15306);
and U16216 (N_16216,N_15743,N_12167);
nand U16217 (N_16217,N_13531,N_13581);
nand U16218 (N_16218,N_15002,N_13563);
and U16219 (N_16219,N_15943,N_13064);
or U16220 (N_16220,N_15063,N_12526);
nor U16221 (N_16221,N_12507,N_15778);
nor U16222 (N_16222,N_14881,N_14123);
or U16223 (N_16223,N_12697,N_13276);
nand U16224 (N_16224,N_15406,N_12918);
nor U16225 (N_16225,N_15388,N_15399);
nor U16226 (N_16226,N_14925,N_14703);
nand U16227 (N_16227,N_13836,N_12616);
nand U16228 (N_16228,N_15346,N_13576);
and U16229 (N_16229,N_13201,N_14438);
nor U16230 (N_16230,N_15164,N_14558);
and U16231 (N_16231,N_13430,N_12098);
or U16232 (N_16232,N_12543,N_13862);
nand U16233 (N_16233,N_14897,N_12362);
nand U16234 (N_16234,N_12611,N_13449);
or U16235 (N_16235,N_13516,N_12867);
nor U16236 (N_16236,N_12449,N_14771);
and U16237 (N_16237,N_15746,N_15848);
nand U16238 (N_16238,N_12933,N_14208);
nor U16239 (N_16239,N_15685,N_13198);
nand U16240 (N_16240,N_13382,N_12159);
or U16241 (N_16241,N_13248,N_15135);
nor U16242 (N_16242,N_13519,N_14069);
nor U16243 (N_16243,N_12915,N_15843);
or U16244 (N_16244,N_13044,N_14815);
nor U16245 (N_16245,N_15662,N_12402);
or U16246 (N_16246,N_15171,N_15709);
xor U16247 (N_16247,N_14765,N_14227);
or U16248 (N_16248,N_12834,N_12909);
nor U16249 (N_16249,N_14013,N_13102);
nor U16250 (N_16250,N_15091,N_13368);
or U16251 (N_16251,N_12104,N_14710);
and U16252 (N_16252,N_12763,N_12877);
or U16253 (N_16253,N_13795,N_13856);
nand U16254 (N_16254,N_14282,N_12329);
nand U16255 (N_16255,N_12790,N_12592);
and U16256 (N_16256,N_12512,N_13811);
or U16257 (N_16257,N_12886,N_15299);
xor U16258 (N_16258,N_14615,N_14751);
or U16259 (N_16259,N_14185,N_15148);
and U16260 (N_16260,N_12179,N_13321);
xnor U16261 (N_16261,N_12500,N_15634);
and U16262 (N_16262,N_15791,N_12714);
and U16263 (N_16263,N_13180,N_13274);
or U16264 (N_16264,N_13435,N_14814);
nor U16265 (N_16265,N_15922,N_15821);
nor U16266 (N_16266,N_14437,N_14357);
or U16267 (N_16267,N_12751,N_15731);
nand U16268 (N_16268,N_13746,N_12152);
nor U16269 (N_16269,N_15130,N_15482);
and U16270 (N_16270,N_12146,N_12966);
and U16271 (N_16271,N_14568,N_13335);
nand U16272 (N_16272,N_13599,N_12919);
and U16273 (N_16273,N_13036,N_12090);
xor U16274 (N_16274,N_13257,N_13716);
xor U16275 (N_16275,N_14184,N_13867);
xor U16276 (N_16276,N_12003,N_14189);
and U16277 (N_16277,N_12297,N_14435);
nand U16278 (N_16278,N_12071,N_13069);
nor U16279 (N_16279,N_14345,N_13633);
or U16280 (N_16280,N_15838,N_15412);
and U16281 (N_16281,N_12339,N_15245);
or U16282 (N_16282,N_13571,N_12789);
or U16283 (N_16283,N_13217,N_15655);
and U16284 (N_16284,N_14445,N_15926);
or U16285 (N_16285,N_14343,N_15720);
nor U16286 (N_16286,N_12788,N_13004);
nor U16287 (N_16287,N_12965,N_15924);
or U16288 (N_16288,N_14162,N_12456);
and U16289 (N_16289,N_14247,N_13562);
nand U16290 (N_16290,N_14775,N_15525);
or U16291 (N_16291,N_13117,N_13858);
or U16292 (N_16292,N_13181,N_13680);
or U16293 (N_16293,N_15976,N_12881);
or U16294 (N_16294,N_13328,N_13254);
or U16295 (N_16295,N_15880,N_13275);
and U16296 (N_16296,N_12433,N_15759);
nand U16297 (N_16297,N_12677,N_14646);
or U16298 (N_16298,N_12882,N_13940);
and U16299 (N_16299,N_13235,N_14188);
or U16300 (N_16300,N_12521,N_15535);
nor U16301 (N_16301,N_12970,N_13475);
nand U16302 (N_16302,N_13933,N_14923);
or U16303 (N_16303,N_13530,N_14723);
nor U16304 (N_16304,N_12284,N_13169);
nor U16305 (N_16305,N_13698,N_12184);
or U16306 (N_16306,N_14931,N_12967);
and U16307 (N_16307,N_13524,N_14687);
or U16308 (N_16308,N_12029,N_12513);
nor U16309 (N_16309,N_12624,N_15868);
nor U16310 (N_16310,N_13611,N_15065);
and U16311 (N_16311,N_14613,N_13806);
nand U16312 (N_16312,N_12728,N_14346);
and U16313 (N_16313,N_12483,N_15211);
or U16314 (N_16314,N_14921,N_14545);
nor U16315 (N_16315,N_15593,N_15621);
nand U16316 (N_16316,N_15760,N_14970);
nand U16317 (N_16317,N_14979,N_15275);
xnor U16318 (N_16318,N_13419,N_15330);
or U16319 (N_16319,N_12696,N_13099);
or U16320 (N_16320,N_13750,N_14706);
and U16321 (N_16321,N_14025,N_15221);
or U16322 (N_16322,N_15937,N_12493);
or U16323 (N_16323,N_12062,N_14092);
or U16324 (N_16324,N_14130,N_14216);
or U16325 (N_16325,N_15297,N_15637);
nand U16326 (N_16326,N_15563,N_15179);
and U16327 (N_16327,N_12059,N_14817);
or U16328 (N_16328,N_15315,N_13300);
nor U16329 (N_16329,N_15956,N_13554);
and U16330 (N_16330,N_12811,N_15624);
xnor U16331 (N_16331,N_15483,N_13392);
or U16332 (N_16332,N_14913,N_13537);
nor U16333 (N_16333,N_14571,N_13617);
or U16334 (N_16334,N_14180,N_15332);
xnor U16335 (N_16335,N_13781,N_15501);
xor U16336 (N_16336,N_12555,N_15573);
and U16337 (N_16337,N_12833,N_14107);
nor U16338 (N_16338,N_15653,N_14264);
nand U16339 (N_16339,N_13232,N_13923);
or U16340 (N_16340,N_12139,N_13622);
and U16341 (N_16341,N_12431,N_14178);
nand U16342 (N_16342,N_13586,N_15103);
nor U16343 (N_16343,N_15107,N_12068);
or U16344 (N_16344,N_13643,N_15886);
or U16345 (N_16345,N_13958,N_14067);
or U16346 (N_16346,N_14690,N_15072);
and U16347 (N_16347,N_14048,N_13955);
nand U16348 (N_16348,N_13610,N_14103);
nand U16349 (N_16349,N_13142,N_12705);
and U16350 (N_16350,N_14868,N_15265);
nand U16351 (N_16351,N_12299,N_13725);
or U16352 (N_16352,N_13573,N_14780);
nand U16353 (N_16353,N_13898,N_13708);
xor U16354 (N_16354,N_12914,N_13697);
or U16355 (N_16355,N_15598,N_12536);
nor U16356 (N_16356,N_14316,N_13249);
nor U16357 (N_16357,N_14322,N_12021);
xor U16358 (N_16358,N_14738,N_13986);
and U16359 (N_16359,N_14014,N_13523);
and U16360 (N_16360,N_15664,N_15461);
nor U16361 (N_16361,N_13227,N_12259);
nor U16362 (N_16362,N_15145,N_14137);
and U16363 (N_16363,N_14888,N_14196);
nand U16364 (N_16364,N_13953,N_14356);
or U16365 (N_16365,N_15479,N_15904);
and U16366 (N_16366,N_12088,N_12749);
and U16367 (N_16367,N_13304,N_15547);
or U16368 (N_16368,N_12584,N_12648);
xor U16369 (N_16369,N_12757,N_13390);
or U16370 (N_16370,N_13535,N_12485);
or U16371 (N_16371,N_12849,N_12314);
xnor U16372 (N_16372,N_15131,N_13966);
nand U16373 (N_16373,N_13315,N_15355);
and U16374 (N_16374,N_15527,N_12741);
nand U16375 (N_16375,N_12980,N_13580);
or U16376 (N_16376,N_14501,N_15796);
xor U16377 (N_16377,N_13970,N_14844);
nand U16378 (N_16378,N_15612,N_12583);
or U16379 (N_16379,N_13821,N_12033);
xor U16380 (N_16380,N_13886,N_14284);
or U16381 (N_16381,N_14947,N_14140);
and U16382 (N_16382,N_14724,N_14951);
nand U16383 (N_16383,N_12794,N_15729);
or U16384 (N_16384,N_12709,N_14492);
or U16385 (N_16385,N_15830,N_13917);
nor U16386 (N_16386,N_14395,N_14739);
and U16387 (N_16387,N_14467,N_15007);
or U16388 (N_16388,N_13015,N_12827);
or U16389 (N_16389,N_15044,N_13710);
nor U16390 (N_16390,N_15835,N_13831);
xnor U16391 (N_16391,N_13583,N_13040);
xor U16392 (N_16392,N_15907,N_15576);
nor U16393 (N_16393,N_14430,N_15913);
nand U16394 (N_16394,N_12327,N_15749);
nand U16395 (N_16395,N_15325,N_12002);
xnor U16396 (N_16396,N_14597,N_12040);
xor U16397 (N_16397,N_12129,N_15883);
nor U16398 (N_16398,N_12349,N_13034);
nor U16399 (N_16399,N_12221,N_15021);
and U16400 (N_16400,N_15840,N_15722);
nor U16401 (N_16401,N_14960,N_15734);
nand U16402 (N_16402,N_14179,N_13900);
nor U16403 (N_16403,N_15726,N_13337);
nand U16404 (N_16404,N_15495,N_12434);
or U16405 (N_16405,N_14303,N_12929);
nor U16406 (N_16406,N_14254,N_14422);
nand U16407 (N_16407,N_12030,N_15392);
or U16408 (N_16408,N_12769,N_12137);
or U16409 (N_16409,N_15152,N_12122);
nand U16410 (N_16410,N_13890,N_13553);
and U16411 (N_16411,N_13521,N_14144);
nor U16412 (N_16412,N_15567,N_12678);
nor U16413 (N_16413,N_13560,N_13914);
nand U16414 (N_16414,N_15176,N_12773);
nand U16415 (N_16415,N_15503,N_12662);
nand U16416 (N_16416,N_13003,N_15733);
or U16417 (N_16417,N_14427,N_13798);
nor U16418 (N_16418,N_15777,N_12191);
or U16419 (N_16419,N_15538,N_15426);
or U16420 (N_16420,N_15139,N_13855);
nor U16421 (N_16421,N_15945,N_15288);
and U16422 (N_16422,N_15805,N_14882);
or U16423 (N_16423,N_15912,N_14339);
and U16424 (N_16424,N_13372,N_13029);
or U16425 (N_16425,N_15957,N_14073);
nor U16426 (N_16426,N_12303,N_12177);
nand U16427 (N_16427,N_12008,N_13299);
nor U16428 (N_16428,N_12628,N_15433);
nand U16429 (N_16429,N_12617,N_15545);
or U16430 (N_16430,N_14630,N_14293);
nand U16431 (N_16431,N_13126,N_15396);
or U16432 (N_16432,N_13336,N_12683);
or U16433 (N_16433,N_15562,N_12636);
or U16434 (N_16434,N_12178,N_14653);
nand U16435 (N_16435,N_14861,N_14966);
or U16436 (N_16436,N_12600,N_15615);
or U16437 (N_16437,N_15676,N_14072);
or U16438 (N_16438,N_12136,N_14637);
and U16439 (N_16439,N_13796,N_14940);
or U16440 (N_16440,N_12274,N_13238);
nor U16441 (N_16441,N_14157,N_13157);
nand U16442 (N_16442,N_13832,N_13311);
and U16443 (N_16443,N_13183,N_13339);
or U16444 (N_16444,N_14573,N_15253);
or U16445 (N_16445,N_13833,N_15752);
and U16446 (N_16446,N_14217,N_12666);
xor U16447 (N_16447,N_12452,N_12004);
nor U16448 (N_16448,N_12250,N_13850);
or U16449 (N_16449,N_15313,N_14606);
xnor U16450 (N_16450,N_15289,N_14628);
nor U16451 (N_16451,N_15052,N_15572);
nor U16452 (N_16452,N_13127,N_13442);
nand U16453 (N_16453,N_14251,N_12847);
nand U16454 (N_16454,N_15651,N_14054);
or U16455 (N_16455,N_15524,N_12482);
nand U16456 (N_16456,N_14354,N_13170);
and U16457 (N_16457,N_12845,N_12391);
and U16458 (N_16458,N_13910,N_15029);
nor U16459 (N_16459,N_14252,N_14819);
nor U16460 (N_16460,N_13055,N_14039);
nand U16461 (N_16461,N_14289,N_15023);
nor U16462 (N_16462,N_15407,N_15920);
nand U16463 (N_16463,N_15142,N_13493);
nor U16464 (N_16464,N_15969,N_13724);
nor U16465 (N_16465,N_14478,N_12465);
or U16466 (N_16466,N_14287,N_13569);
nand U16467 (N_16467,N_14465,N_15097);
nand U16468 (N_16468,N_14320,N_14161);
or U16469 (N_16469,N_14636,N_13369);
nand U16470 (N_16470,N_14838,N_12428);
xnor U16471 (N_16471,N_12528,N_14727);
xor U16472 (N_16472,N_15267,N_15909);
or U16473 (N_16473,N_15670,N_13247);
and U16474 (N_16474,N_12450,N_14064);
nor U16475 (N_16475,N_15057,N_13027);
or U16476 (N_16476,N_14379,N_13601);
and U16477 (N_16477,N_15697,N_13810);
nor U16478 (N_16478,N_13207,N_15128);
nor U16479 (N_16479,N_14862,N_14991);
and U16480 (N_16480,N_12893,N_15588);
xnor U16481 (N_16481,N_13447,N_15911);
nor U16482 (N_16482,N_13902,N_15274);
nor U16483 (N_16483,N_12479,N_12517);
or U16484 (N_16484,N_13915,N_12393);
or U16485 (N_16485,N_13066,N_13607);
nor U16486 (N_16486,N_13837,N_12541);
nand U16487 (N_16487,N_13478,N_15177);
xor U16488 (N_16488,N_14136,N_14880);
nor U16489 (N_16489,N_15896,N_14195);
or U16490 (N_16490,N_12830,N_12876);
nor U16491 (N_16491,N_13788,N_14783);
or U16492 (N_16492,N_15410,N_15988);
nand U16493 (N_16493,N_13679,N_14716);
nor U16494 (N_16494,N_15698,N_13686);
and U16495 (N_16495,N_15358,N_12594);
and U16496 (N_16496,N_13965,N_14643);
or U16497 (N_16497,N_13663,N_15225);
nand U16498 (N_16498,N_15682,N_14100);
or U16499 (N_16499,N_13661,N_13682);
and U16500 (N_16500,N_13025,N_15004);
nand U16501 (N_16501,N_15737,N_15693);
nor U16502 (N_16502,N_12175,N_15669);
nor U16503 (N_16503,N_14503,N_15064);
nand U16504 (N_16504,N_15140,N_12440);
xnor U16505 (N_16505,N_13812,N_15822);
nor U16506 (N_16506,N_12200,N_14858);
nand U16507 (N_16507,N_12319,N_12052);
xor U16508 (N_16508,N_14207,N_14779);
nand U16509 (N_16509,N_15966,N_13773);
and U16510 (N_16510,N_14298,N_15214);
nor U16511 (N_16511,N_13808,N_15865);
nand U16512 (N_16512,N_15233,N_13200);
or U16513 (N_16513,N_14790,N_15244);
and U16514 (N_16514,N_15110,N_15032);
or U16515 (N_16515,N_15643,N_12034);
and U16516 (N_16516,N_14150,N_13849);
nor U16517 (N_16517,N_13656,N_15122);
nor U16518 (N_16518,N_15683,N_13809);
nor U16519 (N_16519,N_13060,N_12341);
or U16520 (N_16520,N_14959,N_15897);
nor U16521 (N_16521,N_12716,N_13268);
nor U16522 (N_16522,N_14419,N_15480);
nand U16523 (N_16523,N_14098,N_14257);
or U16524 (N_16524,N_12287,N_15581);
nor U16525 (N_16525,N_15605,N_13199);
and U16526 (N_16526,N_12291,N_12560);
xor U16527 (N_16527,N_12289,N_15350);
nor U16528 (N_16528,N_12561,N_15936);
or U16529 (N_16529,N_12011,N_15440);
nor U16530 (N_16530,N_13800,N_15570);
or U16531 (N_16531,N_14640,N_12404);
nor U16532 (N_16532,N_14762,N_15413);
or U16533 (N_16533,N_15533,N_13906);
and U16534 (N_16534,N_12272,N_14741);
and U16535 (N_16535,N_15857,N_14059);
or U16536 (N_16536,N_13627,N_15012);
nor U16537 (N_16537,N_12006,N_12304);
nand U16538 (N_16538,N_14202,N_14269);
or U16539 (N_16539,N_14519,N_14521);
xnor U16540 (N_16540,N_13108,N_12127);
nand U16541 (N_16541,N_15804,N_12850);
or U16542 (N_16542,N_15280,N_14803);
xnor U16543 (N_16543,N_13694,N_14145);
or U16544 (N_16544,N_15680,N_15675);
nand U16545 (N_16545,N_15120,N_15424);
nor U16546 (N_16546,N_15951,N_14883);
and U16547 (N_16547,N_13234,N_15003);
nand U16548 (N_16548,N_13061,N_15345);
and U16549 (N_16549,N_13279,N_14263);
nand U16550 (N_16550,N_14344,N_15744);
nor U16551 (N_16551,N_15224,N_14155);
nor U16552 (N_16552,N_15270,N_15803);
and U16553 (N_16553,N_12038,N_13319);
nor U16554 (N_16554,N_14945,N_12470);
nand U16555 (N_16555,N_12778,N_13657);
nor U16556 (N_16556,N_15686,N_15557);
or U16557 (N_16557,N_14793,N_12125);
xnor U16558 (N_16558,N_13536,N_15329);
xor U16559 (N_16559,N_15773,N_12661);
and U16560 (N_16560,N_12185,N_14062);
nor U16561 (N_16561,N_12663,N_14045);
or U16562 (N_16562,N_15959,N_14313);
and U16563 (N_16563,N_13489,N_15587);
nand U16564 (N_16564,N_14611,N_14243);
nand U16565 (N_16565,N_15979,N_15046);
nand U16566 (N_16566,N_14429,N_13048);
or U16567 (N_16567,N_12109,N_15222);
and U16568 (N_16568,N_12447,N_12799);
nor U16569 (N_16569,N_13973,N_12753);
nand U16570 (N_16570,N_12761,N_13263);
and U16571 (N_16571,N_13219,N_15905);
or U16572 (N_16572,N_13981,N_15242);
and U16573 (N_16573,N_12791,N_13340);
and U16574 (N_16574,N_12229,N_14975);
and U16575 (N_16575,N_14663,N_13196);
nand U16576 (N_16576,N_14258,N_12704);
and U16577 (N_16577,N_15982,N_14004);
or U16578 (N_16578,N_14872,N_15983);
nor U16579 (N_16579,N_12346,N_15075);
nand U16580 (N_16580,N_14871,N_13899);
and U16581 (N_16581,N_12055,N_14042);
and U16582 (N_16582,N_15558,N_14255);
and U16583 (N_16583,N_14555,N_14992);
nand U16584 (N_16584,N_13709,N_15797);
nor U16585 (N_16585,N_12457,N_13990);
and U16586 (N_16586,N_13415,N_12643);
nand U16587 (N_16587,N_15376,N_13286);
nor U16588 (N_16588,N_12975,N_13748);
nand U16589 (N_16589,N_15657,N_14292);
nand U16590 (N_16590,N_12039,N_14006);
or U16591 (N_16591,N_12887,N_13059);
nor U16592 (N_16592,N_14610,N_14917);
and U16593 (N_16593,N_15882,N_14768);
nand U16594 (N_16594,N_12051,N_14041);
nor U16595 (N_16595,N_12599,N_12234);
or U16596 (N_16596,N_12087,N_13297);
nand U16597 (N_16597,N_14933,N_14210);
xnor U16598 (N_16598,N_13131,N_13589);
xor U16599 (N_16599,N_12253,N_12671);
nand U16600 (N_16600,N_15568,N_13065);
nand U16601 (N_16601,N_12907,N_13889);
and U16602 (N_16602,N_12548,N_14523);
or U16603 (N_16603,N_13250,N_15146);
nor U16604 (N_16604,N_14736,N_12702);
or U16605 (N_16605,N_12313,N_13101);
or U16606 (N_16606,N_12570,N_15595);
and U16607 (N_16607,N_14261,N_13213);
and U16608 (N_16608,N_12490,N_12244);
and U16609 (N_16609,N_14956,N_15561);
nand U16610 (N_16610,N_12101,N_12036);
nor U16611 (N_16611,N_12340,N_12414);
nor U16612 (N_16612,N_12392,N_15460);
or U16613 (N_16613,N_15181,N_14397);
nor U16614 (N_16614,N_12279,N_12774);
nand U16615 (N_16615,N_15281,N_13112);
or U16616 (N_16616,N_15765,N_14910);
nand U16617 (N_16617,N_15509,N_14604);
and U16618 (N_16618,N_14929,N_14609);
xor U16619 (N_16619,N_15199,N_12119);
nand U16620 (N_16620,N_12993,N_13792);
or U16621 (N_16621,N_14452,N_13230);
or U16622 (N_16622,N_12023,N_12061);
and U16623 (N_16623,N_14843,N_12370);
and U16624 (N_16624,N_13528,N_14318);
or U16625 (N_16625,N_12941,N_14514);
or U16626 (N_16626,N_12813,N_13762);
nand U16627 (N_16627,N_14531,N_12816);
or U16628 (N_16628,N_12667,N_14337);
nand U16629 (N_16629,N_15735,N_14616);
and U16630 (N_16630,N_13735,N_12398);
nand U16631 (N_16631,N_15333,N_12780);
nand U16632 (N_16632,N_14224,N_14327);
nand U16633 (N_16633,N_15687,N_13072);
and U16634 (N_16634,N_12710,N_15194);
and U16635 (N_16635,N_13717,N_15921);
and U16636 (N_16636,N_15314,N_15508);
nor U16637 (N_16637,N_15872,N_14660);
nor U16638 (N_16638,N_15955,N_15610);
and U16639 (N_16639,N_12227,N_13929);
and U16640 (N_16640,N_13012,N_12815);
nand U16641 (N_16641,N_12281,N_13194);
nor U16642 (N_16642,N_14954,N_12233);
or U16643 (N_16643,N_12135,N_12484);
nand U16644 (N_16644,N_12609,N_12944);
or U16645 (N_16645,N_12765,N_13024);
or U16646 (N_16646,N_14654,N_14480);
nor U16647 (N_16647,N_12472,N_13094);
nor U16648 (N_16648,N_13780,N_12024);
and U16649 (N_16649,N_14677,N_12186);
nand U16650 (N_16650,N_14985,N_13212);
nand U16651 (N_16651,N_14109,N_13464);
or U16652 (N_16652,N_12664,N_12080);
nand U16653 (N_16653,N_13208,N_13068);
xor U16654 (N_16654,N_13187,N_12800);
and U16655 (N_16655,N_14891,N_14171);
nor U16656 (N_16656,N_14376,N_13141);
xor U16657 (N_16657,N_12640,N_13732);
nor U16658 (N_16658,N_12562,N_15236);
or U16659 (N_16659,N_15318,N_14030);
nand U16660 (N_16660,N_15432,N_15324);
nor U16661 (N_16661,N_14271,N_14546);
nand U16662 (N_16662,N_13737,N_15102);
xnor U16663 (N_16663,N_12357,N_13409);
or U16664 (N_16664,N_15591,N_13114);
nor U16665 (N_16665,N_14007,N_13753);
xnor U16666 (N_16666,N_12931,N_13487);
or U16667 (N_16667,N_12641,N_14213);
nand U16668 (N_16668,N_14002,N_14104);
nor U16669 (N_16669,N_14839,N_13640);
nor U16670 (N_16670,N_15786,N_12565);
nor U16671 (N_16671,N_13723,N_12522);
or U16672 (N_16672,N_15690,N_12672);
and U16673 (N_16673,N_13429,N_13685);
and U16674 (N_16674,N_12831,N_15466);
or U16675 (N_16675,N_14477,N_13163);
or U16676 (N_16676,N_14476,N_14448);
nand U16677 (N_16677,N_14094,N_12768);
nand U16678 (N_16678,N_14746,N_13222);
nor U16679 (N_16679,N_14394,N_15577);
and U16680 (N_16680,N_12937,N_13350);
nand U16681 (N_16681,N_13695,N_12401);
nor U16682 (N_16682,N_13362,N_15665);
nor U16683 (N_16683,N_13472,N_13995);
nand U16684 (N_16684,N_12558,N_12884);
and U16685 (N_16685,N_12708,N_12128);
nand U16686 (N_16686,N_13410,N_13873);
nor U16687 (N_16687,N_13245,N_15134);
and U16688 (N_16688,N_13512,N_13403);
or U16689 (N_16689,N_12295,N_12820);
nor U16690 (N_16690,N_15105,N_15200);
nor U16691 (N_16691,N_14902,N_14498);
nand U16692 (N_16692,N_14219,N_14091);
or U16693 (N_16693,N_14892,N_12574);
xor U16694 (N_16694,N_15186,N_12650);
and U16695 (N_16695,N_13936,N_12502);
or U16696 (N_16696,N_12880,N_13804);
or U16697 (N_16697,N_14441,N_12770);
and U16698 (N_16698,N_13202,N_14347);
or U16699 (N_16699,N_15650,N_13883);
xnor U16700 (N_16700,N_15649,N_13149);
or U16701 (N_16701,N_13755,N_14374);
and U16702 (N_16702,N_15783,N_14018);
and U16703 (N_16703,N_12693,N_12334);
nor U16704 (N_16704,N_14421,N_12764);
or U16705 (N_16705,N_13786,N_15813);
nand U16706 (N_16706,N_12567,N_15845);
nor U16707 (N_16707,N_15974,N_14638);
or U16708 (N_16708,N_12657,N_14308);
and U16709 (N_16709,N_14743,N_14969);
or U16710 (N_16710,N_14777,N_13529);
xnor U16711 (N_16711,N_15944,N_15196);
and U16712 (N_16712,N_13120,N_14056);
nor U16713 (N_16713,N_12096,N_12498);
or U16714 (N_16714,N_14413,N_14631);
nand U16715 (N_16715,N_12945,N_14796);
nor U16716 (N_16716,N_12509,N_12832);
or U16717 (N_16717,N_12435,N_12806);
or U16718 (N_16718,N_15422,N_12852);
xor U16719 (N_16719,N_13303,N_14513);
or U16720 (N_16720,N_12539,N_12622);
nand U16721 (N_16721,N_15606,N_15335);
xor U16722 (N_16722,N_13638,N_12298);
nor U16723 (N_16723,N_14664,N_15592);
nor U16724 (N_16724,N_12432,N_12568);
and U16725 (N_16725,N_13880,N_12307);
and U16726 (N_16726,N_14623,N_13790);
nor U16727 (N_16727,N_14311,N_15755);
and U16728 (N_16728,N_12383,N_13176);
or U16729 (N_16729,N_14453,N_13613);
nor U16730 (N_16730,N_14786,N_15477);
nor U16731 (N_16731,N_15394,N_15464);
nor U16732 (N_16732,N_12015,N_14548);
xnor U16733 (N_16733,N_12267,N_12105);
and U16734 (N_16734,N_12223,N_12990);
nand U16735 (N_16735,N_14290,N_13294);
nor U16736 (N_16736,N_15112,N_13421);
nor U16737 (N_16737,N_13155,N_12825);
and U16738 (N_16738,N_14887,N_13033);
nor U16739 (N_16739,N_12000,N_13963);
nor U16740 (N_16740,N_15991,N_14505);
nand U16741 (N_16741,N_13132,N_15559);
xor U16742 (N_16742,N_14588,N_14138);
xor U16743 (N_16743,N_15864,N_12787);
nor U16744 (N_16744,N_12792,N_12316);
xor U16745 (N_16745,N_13815,N_14528);
nand U16746 (N_16746,N_13467,N_13282);
xnor U16747 (N_16747,N_13195,N_15384);
xor U16748 (N_16748,N_14846,N_13766);
or U16749 (N_16749,N_15011,N_14057);
nand U16750 (N_16750,N_15256,N_13824);
xor U16751 (N_16751,N_14381,N_13629);
xor U16752 (N_16752,N_12629,N_15473);
or U16753 (N_16753,N_13747,N_13660);
or U16754 (N_16754,N_15180,N_14938);
nor U16755 (N_16755,N_12031,N_14806);
nand U16756 (N_16756,N_14798,N_14502);
nor U16757 (N_16757,N_13143,N_15900);
and U16758 (N_16758,N_14489,N_15444);
or U16759 (N_16759,N_14309,N_12533);
nor U16760 (N_16760,N_15962,N_13829);
or U16761 (N_16761,N_15001,N_12901);
or U16762 (N_16762,N_13628,N_13121);
and U16763 (N_16763,N_12537,N_13948);
nand U16764 (N_16764,N_13188,N_13776);
and U16765 (N_16765,N_12999,N_14500);
or U16766 (N_16766,N_12322,N_14222);
nand U16767 (N_16767,N_12913,N_12903);
nand U16768 (N_16768,N_15429,N_12928);
and U16769 (N_16769,N_12812,N_15356);
and U16770 (N_16770,N_13446,N_15484);
xor U16771 (N_16771,N_14634,N_14756);
nor U16772 (N_16772,N_15635,N_12856);
and U16773 (N_16773,N_14245,N_13712);
xnor U16774 (N_16774,N_14299,N_12044);
xnor U16775 (N_16775,N_13720,N_15847);
xor U16776 (N_16776,N_12955,N_14234);
nand U16777 (N_16777,N_13477,N_15877);
nor U16778 (N_16778,N_15311,N_14825);
xor U16779 (N_16779,N_14393,N_15168);
and U16780 (N_16780,N_12043,N_12445);
nand U16781 (N_16781,N_13742,N_13859);
or U16782 (N_16782,N_14125,N_14682);
or U16783 (N_16783,N_13431,N_14068);
or U16784 (N_16784,N_12211,N_13006);
or U16785 (N_16785,N_14719,N_12425);
and U16786 (N_16786,N_15442,N_13996);
nand U16787 (N_16787,N_15554,N_12625);
or U16788 (N_16788,N_13619,N_14256);
and U16789 (N_16789,N_15992,N_13354);
xnor U16790 (N_16790,N_14961,N_14275);
and U16791 (N_16791,N_15677,N_14592);
nand U16792 (N_16792,N_14046,N_15859);
or U16793 (N_16793,N_13352,N_15090);
or U16794 (N_16794,N_12446,N_14128);
xor U16795 (N_16795,N_14367,N_14621);
and U16796 (N_16796,N_12618,N_14070);
or U16797 (N_16797,N_15678,N_14856);
nand U16798 (N_16798,N_12280,N_13864);
nand U16799 (N_16799,N_12905,N_15104);
nand U16800 (N_16800,N_15769,N_15045);
nand U16801 (N_16801,N_13678,N_14763);
or U16802 (N_16802,N_12145,N_13551);
nor U16803 (N_16803,N_15188,N_12608);
nand U16804 (N_16804,N_13402,N_13636);
or U16805 (N_16805,N_14493,N_12271);
nand U16806 (N_16806,N_14456,N_13258);
nand U16807 (N_16807,N_15809,N_14300);
and U16808 (N_16808,N_14008,N_15742);
xor U16809 (N_16809,N_13193,N_12164);
and U16810 (N_16810,N_12766,N_13492);
nor U16811 (N_16811,N_12688,N_15639);
or U16812 (N_16812,N_12217,N_14544);
nor U16813 (N_16813,N_13803,N_12487);
and U16814 (N_16814,N_12958,N_12596);
nor U16815 (N_16815,N_12544,N_12163);
nor U16816 (N_16816,N_14183,N_13295);
nand U16817 (N_16817,N_12531,N_14950);
nor U16818 (N_16818,N_13399,N_15842);
and U16819 (N_16819,N_15569,N_12444);
nor U16820 (N_16820,N_15961,N_12582);
and U16821 (N_16821,N_13018,N_13972);
nor U16822 (N_16822,N_15371,N_12963);
or U16823 (N_16823,N_15282,N_15088);
and U16824 (N_16824,N_13908,N_12860);
and U16825 (N_16825,N_12066,N_14700);
nor U16826 (N_16826,N_14829,N_14159);
and U16827 (N_16827,N_14927,N_12817);
and U16828 (N_16828,N_14944,N_12016);
xnor U16829 (N_16829,N_12454,N_15564);
xnor U16830 (N_16830,N_12406,N_13416);
xor U16831 (N_16831,N_12196,N_13479);
or U16832 (N_16832,N_15958,N_13513);
nor U16833 (N_16833,N_14909,N_14442);
or U16834 (N_16834,N_15642,N_13844);
and U16835 (N_16835,N_12097,N_15918);
nand U16836 (N_16836,N_13151,N_13782);
xnor U16837 (N_16837,N_15512,N_12077);
nand U16838 (N_16838,N_15430,N_14081);
and U16839 (N_16839,N_14142,N_15183);
nor U16840 (N_16840,N_12240,N_14156);
or U16841 (N_16841,N_15774,N_12144);
and U16842 (N_16842,N_15030,N_14766);
nor U16843 (N_16843,N_12891,N_13615);
nand U16844 (N_16844,N_12050,N_15713);
or U16845 (N_16845,N_13438,N_12193);
nand U16846 (N_16846,N_12155,N_12576);
nor U16847 (N_16847,N_14095,N_13758);
or U16848 (N_16848,N_14127,N_13038);
nor U16849 (N_16849,N_14542,N_12610);
nor U16850 (N_16850,N_15475,N_13305);
and U16851 (N_16851,N_14968,N_15017);
nand U16852 (N_16852,N_12118,N_14952);
or U16853 (N_16853,N_14863,N_14387);
and U16854 (N_16854,N_12262,N_15302);
or U16855 (N_16855,N_13246,N_13273);
nor U16856 (N_16856,N_14223,N_15543);
or U16857 (N_16857,N_15641,N_15553);
nand U16858 (N_16858,N_12987,N_15038);
or U16859 (N_16859,N_13313,N_14939);
or U16860 (N_16860,N_14335,N_15986);
nor U16861 (N_16861,N_15447,N_14635);
xor U16862 (N_16862,N_13683,N_15155);
nand U16863 (N_16863,N_12497,N_12252);
nand U16864 (N_16864,N_13049,N_13075);
and U16865 (N_16865,N_15334,N_12579);
nand U16866 (N_16866,N_13546,N_14462);
nor U16867 (N_16867,N_12898,N_14231);
nand U16868 (N_16868,N_15827,N_14330);
xor U16869 (N_16869,N_12360,N_13105);
nand U16870 (N_16870,N_14755,N_15402);
or U16871 (N_16871,N_14237,N_13253);
or U16872 (N_16872,N_13042,N_14444);
nand U16873 (N_16873,N_15950,N_15792);
and U16874 (N_16874,N_15491,N_13356);
xnor U16875 (N_16875,N_13532,N_13330);
nor U16876 (N_16876,N_14259,N_15630);
nand U16877 (N_16877,N_13013,N_15008);
nor U16878 (N_16878,N_13272,N_12598);
or U16879 (N_16879,N_13860,N_12255);
and U16880 (N_16880,N_13424,N_12048);
and U16881 (N_16881,N_13462,N_12843);
nand U16882 (N_16882,N_12838,N_14389);
and U16883 (N_16883,N_13944,N_14038);
and U16884 (N_16884,N_15082,N_13920);
nor U16885 (N_16885,N_13740,N_12418);
nand U16886 (N_16886,N_14277,N_14977);
or U16887 (N_16887,N_12308,N_13624);
xnor U16888 (N_16888,N_14450,N_15465);
nor U16889 (N_16889,N_14304,N_13612);
and U16890 (N_16890,N_15226,N_13262);
nand U16891 (N_16891,N_15266,N_15623);
and U16892 (N_16892,N_14774,N_14584);
or U16893 (N_16893,N_13820,N_15377);
xor U16894 (N_16894,N_12679,N_14794);
xnor U16895 (N_16895,N_13278,N_15714);
nand U16896 (N_16896,N_13509,N_15906);
and U16897 (N_16897,N_14003,N_13655);
nand U16898 (N_16898,N_13139,N_15393);
and U16899 (N_16899,N_15307,N_14577);
nand U16900 (N_16900,N_12862,N_13395);
nor U16901 (N_16901,N_13357,N_12294);
or U16902 (N_16902,N_14633,N_14569);
or U16903 (N_16903,N_13000,N_12046);
xnor U16904 (N_16904,N_13150,N_15087);
nand U16905 (N_16905,N_13882,N_14900);
and U16906 (N_16906,N_14873,N_12613);
nor U16907 (N_16907,N_15312,N_15441);
or U16908 (N_16908,N_15010,N_15080);
xor U16909 (N_16909,N_15820,N_12637);
or U16910 (N_16910,N_15374,N_15448);
nand U16911 (N_16911,N_15454,N_12976);
nor U16912 (N_16912,N_15411,N_14126);
and U16913 (N_16913,N_12861,N_12417);
and U16914 (N_16914,N_13527,N_15060);
nor U16915 (N_16915,N_12413,N_12181);
and U16916 (N_16916,N_15207,N_12732);
nand U16917 (N_16917,N_12489,N_13897);
and U16918 (N_16918,N_13514,N_15340);
or U16919 (N_16919,N_12149,N_15964);
and U16920 (N_16920,N_13444,N_12156);
and U16921 (N_16921,N_14473,N_12203);
xnor U16922 (N_16922,N_15756,N_14015);
xnor U16923 (N_16923,N_13085,N_15818);
and U16924 (N_16924,N_12143,N_15638);
or U16925 (N_16925,N_15552,N_12212);
nand U16926 (N_16926,N_14549,N_14129);
or U16927 (N_16927,N_12997,N_14464);
and U16928 (N_16928,N_13649,N_15887);
or U16929 (N_16929,N_13552,N_14086);
nor U16930 (N_16930,N_12738,N_12828);
and U16931 (N_16931,N_12949,N_14332);
xor U16932 (N_16932,N_12602,N_14722);
nand U16933 (N_16933,N_14267,N_13674);
or U16934 (N_16934,N_13830,N_15205);
or U16935 (N_16935,N_13608,N_14108);
or U16936 (N_16936,N_12220,N_15967);
nor U16937 (N_16937,N_13456,N_14471);
nor U16938 (N_16938,N_15235,N_12699);
or U16939 (N_16939,N_13133,N_15529);
nor U16940 (N_16940,N_12422,N_12243);
or U16941 (N_16941,N_14955,N_15321);
nor U16942 (N_16942,N_14567,N_14973);
nand U16943 (N_16943,N_12872,N_15028);
nand U16944 (N_16944,N_12013,N_12606);
nand U16945 (N_16945,N_15691,N_12380);
and U16946 (N_16946,N_13323,N_12351);
xor U16947 (N_16947,N_13949,N_12668);
or U16948 (N_16948,N_12706,N_15414);
nand U16949 (N_16949,N_14182,N_14914);
nand U16950 (N_16950,N_13848,N_13097);
or U16951 (N_16951,N_13022,N_13138);
or U16952 (N_16952,N_14325,N_12373);
or U16953 (N_16953,N_15980,N_15522);
nor U16954 (N_16954,N_15898,N_14075);
and U16955 (N_16955,N_13379,N_12995);
xnor U16956 (N_16956,N_14893,N_13539);
nand U16957 (N_16957,N_14475,N_12906);
nand U16958 (N_16958,N_13463,N_13302);
nor U16959 (N_16959,N_14433,N_14586);
nor U16960 (N_16960,N_12201,N_15575);
nand U16961 (N_16961,N_12923,N_15425);
or U16962 (N_16962,N_15227,N_15878);
and U16963 (N_16963,N_12908,N_12361);
xor U16964 (N_16964,N_14268,N_15523);
and U16965 (N_16965,N_15815,N_13014);
nor U16966 (N_16966,N_13261,N_14801);
nand U16967 (N_16967,N_15323,N_13146);
and U16968 (N_16968,N_13124,N_14805);
nor U16969 (N_16969,N_13999,N_14816);
nor U16970 (N_16970,N_13621,N_14112);
nand U16971 (N_16971,N_14889,N_12158);
or U16972 (N_16972,N_13501,N_12998);
nor U16973 (N_16973,N_14733,N_14524);
nor U16974 (N_16974,N_13752,N_14369);
nand U16975 (N_16975,N_14472,N_12868);
and U16976 (N_16976,N_14625,N_14668);
xor U16977 (N_16977,N_12585,N_12809);
nand U16978 (N_16978,N_12566,N_12009);
nand U16979 (N_16979,N_13076,N_15566);
nor U16980 (N_16980,N_13688,N_13604);
and U16981 (N_16981,N_15993,N_13540);
nor U16982 (N_16982,N_15248,N_15507);
nor U16983 (N_16983,N_13370,N_13280);
and U16984 (N_16984,N_13398,N_14076);
nor U16985 (N_16985,N_14834,N_13700);
xnor U16986 (N_16986,N_12476,N_12020);
or U16987 (N_16987,N_12591,N_14986);
xor U16988 (N_16988,N_13291,N_12083);
nand U16989 (N_16989,N_12865,N_15452);
or U16990 (N_16990,N_13518,N_14942);
nand U16991 (N_16991,N_14757,N_14341);
or U16992 (N_16992,N_14576,N_13775);
nand U16993 (N_16993,N_15054,N_13658);
nor U16994 (N_16994,N_15548,N_15293);
and U16995 (N_16995,N_14040,N_13852);
and U16996 (N_16996,N_13458,N_14017);
nand U16997 (N_16997,N_12276,N_14132);
nand U16998 (N_16998,N_13704,N_12142);
nand U16999 (N_16999,N_12855,N_14191);
xor U17000 (N_17000,N_12894,N_13652);
nor U17001 (N_17001,N_14333,N_15965);
nor U17002 (N_17002,N_12285,N_13729);
or U17003 (N_17003,N_14704,N_13504);
xnor U17004 (N_17004,N_14833,N_12226);
or U17005 (N_17005,N_14810,N_15055);
xnor U17006 (N_17006,N_14581,N_14823);
nor U17007 (N_17007,N_13107,N_12595);
nor U17008 (N_17008,N_13244,N_15526);
nand U17009 (N_17009,N_15816,N_12273);
xor U17010 (N_17010,N_15239,N_12701);
xor U17011 (N_17011,N_14958,N_14055);
nand U17012 (N_17012,N_13895,N_12378);
nand U17013 (N_17013,N_12577,N_14642);
and U17014 (N_17014,N_12631,N_12925);
and U17015 (N_17015,N_13714,N_14481);
and U17016 (N_17016,N_15215,N_12121);
nor U17017 (N_17017,N_12962,N_12364);
or U17018 (N_17018,N_13797,N_14163);
or U17019 (N_17019,N_15889,N_14543);
nor U17020 (N_17020,N_14370,N_12559);
and U17021 (N_17021,N_12093,N_12501);
and U17022 (N_17022,N_13668,N_14302);
nor U17023 (N_17023,N_15443,N_12518);
nand U17024 (N_17024,N_14044,N_12251);
and U17025 (N_17025,N_13872,N_15879);
nor U17026 (N_17026,N_15459,N_14023);
and U17027 (N_17027,N_13577,N_15320);
or U17028 (N_17028,N_15513,N_14139);
nand U17029 (N_17029,N_13606,N_14683);
nor U17030 (N_17030,N_15910,N_14301);
and U17031 (N_17031,N_13517,N_14582);
nand U17032 (N_17032,N_13125,N_12210);
nor U17033 (N_17033,N_13769,N_14499);
nand U17034 (N_17034,N_12443,N_13229);
or U17035 (N_17035,N_14460,N_15892);
or U17036 (N_17036,N_15468,N_13651);
nand U17037 (N_17037,N_14657,N_14731);
nor U17038 (N_17038,N_14879,N_14818);
or U17039 (N_17039,N_13645,N_15539);
nand U17040 (N_17040,N_15341,N_14461);
nor U17041 (N_17041,N_12377,N_15328);
nor U17042 (N_17042,N_12190,N_14504);
and U17043 (N_17043,N_13461,N_12017);
and U17044 (N_17044,N_13136,N_13835);
nand U17045 (N_17045,N_12363,N_13347);
or U17046 (N_17046,N_15939,N_14855);
or U17047 (N_17047,N_13269,N_12578);
nor U17048 (N_17048,N_13408,N_15451);
nor U17049 (N_17049,N_14593,N_15861);
or U17050 (N_17050,N_12168,N_13158);
and U17051 (N_17051,N_13572,N_15658);
nand U17052 (N_17052,N_12007,N_15544);
or U17053 (N_17053,N_13787,N_14361);
or U17054 (N_17054,N_15076,N_14532);
and U17055 (N_17055,N_15362,N_12310);
nand U17056 (N_17056,N_14326,N_14649);
nand U17057 (N_17057,N_15617,N_12745);
nand U17058 (N_17058,N_15423,N_15361);
nor U17059 (N_17059,N_15846,N_14463);
nand U17060 (N_17060,N_15894,N_15370);
and U17061 (N_17061,N_14937,N_13932);
nand U17062 (N_17062,N_14052,N_12293);
nand U17063 (N_17063,N_12292,N_14876);
and U17064 (N_17064,N_12516,N_15987);
nor U17065 (N_17065,N_12904,N_13166);
or U17066 (N_17066,N_12106,N_12448);
and U17067 (N_17067,N_12183,N_15625);
and U17068 (N_17068,N_15185,N_12134);
or U17069 (N_17069,N_13079,N_13252);
nor U17070 (N_17070,N_12455,N_13407);
nor U17071 (N_17071,N_12231,N_15159);
or U17072 (N_17072,N_12328,N_13823);
and U17073 (N_17073,N_12286,N_12814);
or U17074 (N_17074,N_15971,N_14288);
nand U17075 (N_17075,N_13574,N_12462);
or U17076 (N_17076,N_14186,N_13980);
and U17077 (N_17077,N_13508,N_14285);
nor U17078 (N_17078,N_14671,N_14494);
and U17079 (N_17079,N_13422,N_14744);
and U17080 (N_17080,N_12395,N_13561);
and U17081 (N_17081,N_14151,N_12588);
or U17082 (N_17082,N_12659,N_13962);
or U17083 (N_17083,N_12532,N_15232);
or U17084 (N_17084,N_13991,N_13417);
nor U17085 (N_17085,N_14079,N_15000);
nor U17086 (N_17086,N_14228,N_12797);
nand U17087 (N_17087,N_15854,N_12656);
or U17088 (N_17088,N_15681,N_14976);
and U17089 (N_17089,N_12807,N_13215);
or U17090 (N_17090,N_15753,N_13715);
and U17091 (N_17091,N_14990,N_14033);
or U17092 (N_17092,N_15885,N_14845);
or U17093 (N_17093,N_14759,N_13366);
nor U17094 (N_17094,N_15463,N_13595);
and U17095 (N_17095,N_15850,N_15375);
or U17096 (N_17096,N_12333,N_13349);
and U17097 (N_17097,N_13677,N_14848);
nand U17098 (N_17098,N_15009,N_14382);
nor U17099 (N_17099,N_14175,N_14550);
nor U17100 (N_17100,N_15115,N_15583);
nand U17101 (N_17101,N_12803,N_13544);
and U17102 (N_17102,N_12095,N_12219);
xor U17103 (N_17103,N_13770,N_14418);
or U17104 (N_17104,N_13123,N_14984);
xnor U17105 (N_17105,N_13016,N_15705);
xnor U17106 (N_17106,N_13405,N_14820);
nand U17107 (N_17107,N_15500,N_12166);
nor U17108 (N_17108,N_12369,N_14240);
or U17109 (N_17109,N_15398,N_12037);
nand U17110 (N_17110,N_13376,N_12726);
or U17111 (N_17111,N_13148,N_14885);
or U17112 (N_17112,N_15099,N_15382);
nor U17113 (N_17113,N_13499,N_13984);
and U17114 (N_17114,N_14050,N_13777);
or U17115 (N_17115,N_14260,N_13360);
nand U17116 (N_17116,N_14590,N_15636);
nor U17117 (N_17117,N_14619,N_15478);
and U17118 (N_17118,N_15915,N_13743);
nor U17119 (N_17119,N_14010,N_14557);
xnor U17120 (N_17120,N_12161,N_12634);
or U17121 (N_17121,N_13987,N_15616);
nor U17122 (N_17122,N_13863,N_15640);
nand U17123 (N_17123,N_14458,N_13959);
and U17124 (N_17124,N_15806,N_14404);
nand U17125 (N_17125,N_13918,N_14034);
nor U17126 (N_17126,N_12514,N_13383);
nand U17127 (N_17127,N_15511,N_13943);
nor U17128 (N_17128,N_13570,N_14114);
xor U17129 (N_17129,N_14618,N_12420);
nor U17130 (N_17130,N_15238,N_13807);
nor U17131 (N_17131,N_15339,N_12342);
nand U17132 (N_17132,N_13681,N_13893);
and U17133 (N_17133,N_15929,N_13707);
or U17134 (N_17134,N_13404,N_15497);
or U17135 (N_17135,N_13432,N_15039);
or U17136 (N_17136,N_12073,N_15450);
nor U17137 (N_17137,N_14693,N_15970);
and U17138 (N_17138,N_13388,N_14229);
nand U17139 (N_17139,N_13378,N_13559);
or U17140 (N_17140,N_12653,N_15574);
or U17141 (N_17141,N_13623,N_14907);
xnor U17142 (N_17142,N_15519,N_12524);
or U17143 (N_17143,N_15604,N_12480);
nand U17144 (N_17144,N_13256,N_12960);
xnor U17145 (N_17145,N_15094,N_12684);
or U17146 (N_17146,N_12730,N_14585);
nor U17147 (N_17147,N_15151,N_14085);
and U17148 (N_17148,N_12321,N_13223);
or U17149 (N_17149,N_15163,N_15357);
nor U17150 (N_17150,N_14509,N_13702);
nand U17151 (N_17151,N_12863,N_13871);
or U17152 (N_17152,N_14559,N_12916);
nand U17153 (N_17153,N_15518,N_15342);
nand U17154 (N_17154,N_14000,N_13271);
or U17155 (N_17155,N_14689,N_13160);
nor U17156 (N_17156,N_13056,N_13333);
nor U17157 (N_17157,N_13465,N_15963);
and U17158 (N_17158,N_12407,N_13281);
xnor U17159 (N_17159,N_13005,N_13118);
nor U17160 (N_17160,N_12601,N_12742);
and U17161 (N_17161,N_13401,N_13052);
or U17162 (N_17162,N_14377,N_12160);
or U17163 (N_17163,N_14676,N_14681);
xor U17164 (N_17164,N_13924,N_14084);
and U17165 (N_17165,N_15436,N_15486);
xor U17166 (N_17166,N_13332,N_13754);
and U17167 (N_17167,N_12379,N_12384);
nor U17168 (N_17168,N_15372,N_15101);
nand U17169 (N_17169,N_14336,N_13466);
xnor U17170 (N_17170,N_14575,N_14522);
or U17171 (N_17171,N_12027,N_15960);
xor U17172 (N_17172,N_15123,N_13498);
nand U17173 (N_17173,N_12575,N_15663);
and U17174 (N_17174,N_12290,N_12926);
or U17175 (N_17175,N_13474,N_13935);
or U17176 (N_17176,N_13888,N_14167);
nor U17177 (N_17177,N_13179,N_14995);
nor U17178 (N_17178,N_15327,N_12752);
xor U17179 (N_17179,N_12141,N_13975);
nor U17180 (N_17180,N_12974,N_15858);
nand U17181 (N_17181,N_12552,N_14547);
and U17182 (N_17182,N_15034,N_14579);
or U17183 (N_17183,N_13706,N_14270);
or U17184 (N_17184,N_13596,N_14378);
nand U17185 (N_17185,N_14286,N_12735);
nand U17186 (N_17186,N_12632,N_12388);
nand U17187 (N_17187,N_13939,N_12553);
and U17188 (N_17188,N_15844,N_15079);
or U17189 (N_17189,N_15420,N_12890);
xor U17190 (N_17190,N_15397,N_15873);
and U17191 (N_17191,N_15069,N_12256);
and U17192 (N_17192,N_15416,N_14273);
or U17193 (N_17193,N_15578,N_13175);
and U17194 (N_17194,N_12858,N_14971);
xor U17195 (N_17195,N_14894,N_13626);
and U17196 (N_17196,N_15532,N_13317);
and U17197 (N_17197,N_12471,N_12382);
nand U17198 (N_17198,N_12771,N_14791);
or U17199 (N_17199,N_15251,N_15555);
xor U17200 (N_17200,N_14459,N_12495);
nor U17201 (N_17201,N_15727,N_14936);
nor U17202 (N_17202,N_12486,N_13087);
or U17203 (N_17203,N_15875,N_15829);
xor U17204 (N_17204,N_13978,N_14011);
and U17205 (N_17205,N_12120,N_12777);
xor U17206 (N_17206,N_12326,N_13662);
or U17207 (N_17207,N_13008,N_14411);
or U17208 (N_17208,N_15724,N_15661);
nand U17209 (N_17209,N_12525,N_15717);
xor U17210 (N_17210,N_15741,N_13567);
and U17211 (N_17211,N_14589,N_13009);
and U17212 (N_17212,N_15471,N_15317);
or U17213 (N_17213,N_14174,N_14591);
nor U17214 (N_17214,N_13174,N_15068);
or U17215 (N_17215,N_14314,N_12138);
nand U17216 (N_17216,N_14516,N_13511);
or U17217 (N_17217,N_15337,N_14384);
nor U17218 (N_17218,N_13290,N_12744);
nor U17219 (N_17219,N_15114,N_15981);
and U17220 (N_17220,N_13749,N_14605);
xnor U17221 (N_17221,N_14276,N_13870);
nand U17222 (N_17222,N_14847,N_14199);
nor U17223 (N_17223,N_13566,N_14176);
nand U17224 (N_17224,N_12224,N_13556);
or U17225 (N_17225,N_13609,N_12888);
nand U17226 (N_17226,N_15673,N_13894);
or U17227 (N_17227,N_14680,N_15352);
nand U17228 (N_17228,N_15925,N_12047);
xor U17229 (N_17229,N_12301,N_13503);
nor U17230 (N_17230,N_12356,N_14165);
and U17231 (N_17231,N_15530,N_15647);
xor U17232 (N_17232,N_13359,N_12306);
and U17233 (N_17233,N_13500,N_15041);
nor U17234 (N_17234,N_12424,N_12157);
nand U17235 (N_17235,N_12597,N_12408);
or U17236 (N_17236,N_13768,N_12439);
and U17237 (N_17237,N_13799,N_12959);
and U17238 (N_17238,N_13450,N_13903);
or U17239 (N_17239,N_15571,N_12954);
nor U17240 (N_17240,N_13054,N_15834);
nand U17241 (N_17241,N_14334,N_14998);
or U17242 (N_17242,N_14916,N_14946);
or U17243 (N_17243,N_12189,N_12505);
nand U17244 (N_17244,N_15494,N_15326);
xor U17245 (N_17245,N_14599,N_13639);
nand U17246 (N_17246,N_14203,N_14760);
nor U17247 (N_17247,N_15836,N_15240);
and U17248 (N_17248,N_15489,N_12116);
and U17249 (N_17249,N_12821,N_14895);
xor U17250 (N_17250,N_12551,N_15458);
nor U17251 (N_17251,N_14854,N_12946);
nand U17252 (N_17252,N_12478,N_14016);
nand U17253 (N_17253,N_13763,N_13802);
nand U17254 (N_17254,N_15106,N_14915);
and U17255 (N_17255,N_15020,N_13919);
nand U17256 (N_17256,N_15470,N_12996);
and U17257 (N_17257,N_12841,N_12400);
nor U17258 (N_17258,N_12782,N_12515);
and U17259 (N_17259,N_15309,N_15549);
nand U17260 (N_17260,N_13367,N_14530);
nand U17261 (N_17261,N_15066,N_12315);
or U17262 (N_17262,N_15721,N_14209);
nor U17263 (N_17263,N_15400,N_15206);
or U17264 (N_17264,N_14684,N_12494);
nand U17265 (N_17265,N_13428,N_13744);
or U17266 (N_17266,N_12964,N_14474);
xnor U17267 (N_17267,N_14930,N_12535);
and U17268 (N_17268,N_15298,N_14053);
and U17269 (N_17269,N_14626,N_14912);
and U17270 (N_17270,N_12074,N_15117);
nand U17271 (N_17271,N_13001,N_13701);
or U17272 (N_17272,N_14877,N_14541);
or U17273 (N_17273,N_13448,N_13922);
nand U17274 (N_17274,N_12810,N_15116);
nor U17275 (N_17275,N_13520,N_12054);
nor U17276 (N_17276,N_15300,N_13505);
nand U17277 (N_17277,N_14926,N_13921);
and U17278 (N_17278,N_15292,N_15178);
nand U17279 (N_17279,N_14639,N_14154);
nor U17280 (N_17280,N_12724,N_12325);
or U17281 (N_17281,N_15059,N_15191);
xor U17282 (N_17282,N_15127,N_13266);
and U17283 (N_17283,N_15626,N_15234);
nor U17284 (N_17284,N_15269,N_15855);
or U17285 (N_17285,N_13853,N_12586);
or U17286 (N_17286,N_15819,N_12823);
nand U17287 (N_17287,N_15136,N_13095);
nand U17288 (N_17288,N_12460,N_14021);
xnor U17289 (N_17289,N_12195,N_15537);
or U17290 (N_17290,N_15472,N_12056);
nand U17291 (N_17291,N_12075,N_15599);
nand U17292 (N_17292,N_15428,N_12740);
xnor U17293 (N_17293,N_15607,N_15541);
and U17294 (N_17294,N_14694,N_12260);
and U17295 (N_17295,N_15689,N_14143);
or U17296 (N_17296,N_12572,N_12018);
xor U17297 (N_17297,N_12099,N_13385);
nand U17298 (N_17298,N_12463,N_12660);
nand U17299 (N_17299,N_14748,N_15018);
or U17300 (N_17300,N_15536,N_12442);
nor U17301 (N_17301,N_13406,N_14454);
and U17302 (N_17302,N_13925,N_15086);
and U17303 (N_17303,N_14372,N_13325);
nand U17304 (N_17304,N_12057,N_13164);
and U17305 (N_17305,N_15597,N_12162);
and U17306 (N_17306,N_15033,N_14890);
and U17307 (N_17307,N_15261,N_12070);
or U17308 (N_17308,N_13847,N_13983);
nand U17309 (N_17309,N_12266,N_15736);
nor U17310 (N_17310,N_15492,N_14878);
nand U17311 (N_17311,N_15364,N_14852);
and U17312 (N_17312,N_15684,N_15504);
nor U17313 (N_17313,N_14412,N_12305);
nand U17314 (N_17314,N_14556,N_14242);
nand U17315 (N_17315,N_14728,N_13334);
and U17316 (N_17316,N_14121,N_14274);
nand U17317 (N_17317,N_12419,N_13726);
nand U17318 (N_17318,N_12028,N_13237);
nand U17319 (N_17319,N_15217,N_14999);
nand U17320 (N_17320,N_14972,N_13969);
and U17321 (N_17321,N_14696,N_14146);
xor U17322 (N_17322,N_15938,N_13699);
nand U17323 (N_17323,N_14758,N_12140);
nand U17324 (N_17324,N_13486,N_12895);
nand U17325 (N_17325,N_15790,N_12649);
nor U17326 (N_17326,N_12010,N_15505);
or U17327 (N_17327,N_14198,N_13177);
and U17328 (N_17328,N_13039,N_15273);
or U17329 (N_17329,N_12991,N_15715);
or U17330 (N_17330,N_12589,N_15438);
and U17331 (N_17331,N_14526,N_15935);
nor U17332 (N_17332,N_15852,N_13259);
or U17333 (N_17333,N_14233,N_14031);
or U17334 (N_17334,N_14310,N_12713);
and U17335 (N_17335,N_12529,N_15022);
nor U17336 (N_17336,N_14898,N_12924);
and U17337 (N_17337,N_14726,N_13670);
nor U17338 (N_17338,N_14226,N_12358);
nand U17339 (N_17339,N_13653,N_12779);
and U17340 (N_17340,N_15995,N_13993);
and U17341 (N_17341,N_15488,N_14540);
nor U17342 (N_17342,N_15165,N_14200);
and U17343 (N_17343,N_12604,N_14088);
nor U17344 (N_17344,N_14730,N_13051);
xor U17345 (N_17345,N_14807,N_15071);
nor U17346 (N_17346,N_14250,N_14058);
and U17347 (N_17347,N_14778,N_14426);
xor U17348 (N_17348,N_13533,N_13730);
and U17349 (N_17349,N_13411,N_13687);
and U17350 (N_17350,N_13931,N_14715);
and U17351 (N_17351,N_12836,N_12703);
nor U17352 (N_17352,N_15940,N_14685);
and U17353 (N_17353,N_13672,N_12739);
xnor U17354 (N_17354,N_13412,N_15209);
and U17355 (N_17355,N_12111,N_15419);
nor U17356 (N_17356,N_14622,N_15771);
nor U17357 (N_17357,N_15121,N_14903);
and U17358 (N_17358,N_13785,N_12973);
nor U17359 (N_17359,N_12846,N_14439);
nand U17360 (N_17360,N_13927,N_15700);
nand U17361 (N_17361,N_15143,N_14321);
or U17362 (N_17362,N_12676,N_12246);
and U17363 (N_17363,N_15296,N_12278);
and U17364 (N_17364,N_14800,N_13774);
nand U17365 (N_17365,N_13997,N_12680);
and U17366 (N_17366,N_13579,N_12687);
nor U17367 (N_17367,N_13851,N_12978);
or U17368 (N_17368,N_15711,N_12354);
and U17369 (N_17369,N_13173,N_13437);
or U17370 (N_17370,N_15201,N_14331);
and U17371 (N_17371,N_12371,N_14686);
nor U17372 (N_17372,N_13879,N_12665);
nand U17373 (N_17373,N_12620,N_13502);
and U17374 (N_17374,N_12348,N_15387);
nor U17375 (N_17375,N_13846,N_12236);
or U17376 (N_17376,N_13819,N_13380);
or U17377 (N_17377,N_12520,N_15250);
nand U17378 (N_17378,N_12124,N_15453);
nor U17379 (N_17379,N_13558,N_15241);
nand U17380 (N_17380,N_12547,N_13971);
nor U17381 (N_17381,N_14784,N_15949);
and U17382 (N_17382,N_12712,N_13950);
nand U17383 (N_17383,N_14607,N_13397);
or U17384 (N_17384,N_13728,N_14113);
nor U17385 (N_17385,N_15901,N_15808);
nand U17386 (N_17386,N_13618,N_13346);
nor U17387 (N_17387,N_13693,N_15343);
or U17388 (N_17388,N_13425,N_12942);
or U17389 (N_17389,N_15862,N_15259);
or U17390 (N_17390,N_14574,N_13152);
nand U17391 (N_17391,N_12670,N_14565);
nand U17392 (N_17392,N_14603,N_12110);
and U17393 (N_17393,N_15354,N_12605);
or U17394 (N_17394,N_13147,N_12437);
nor U17395 (N_17395,N_13676,N_12781);
nand U17396 (N_17396,N_12019,N_15347);
nor U17397 (N_17397,N_12427,N_12258);
and U17398 (N_17398,N_14679,N_13203);
or U17399 (N_17399,N_14749,N_13122);
nand U17400 (N_17400,N_13192,N_14515);
and U17401 (N_17401,N_14932,N_14266);
and U17402 (N_17402,N_12123,N_12131);
xor U17403 (N_17403,N_13896,N_13994);
or U17404 (N_17404,N_13226,N_15703);
nand U17405 (N_17405,N_15534,N_13582);
nand U17406 (N_17406,N_12065,N_13496);
or U17407 (N_17407,N_15609,N_14077);
xor U17408 (N_17408,N_15619,N_12950);
and U17409 (N_17409,N_12721,N_15255);
or U17410 (N_17410,N_12718,N_13941);
nand U17411 (N_17411,N_14911,N_13074);
nand U17412 (N_17412,N_12345,N_13046);
xnor U17413 (N_17413,N_13365,N_15019);
nand U17414 (N_17414,N_14352,N_15754);
nand U17415 (N_17415,N_12854,N_15161);
nor U17416 (N_17416,N_15409,N_12879);
or U17417 (N_17417,N_13371,N_12695);
nand U17418 (N_17418,N_15005,N_12982);
nor U17419 (N_17419,N_12264,N_14828);
nor U17420 (N_17420,N_14720,N_12654);
and U17421 (N_17421,N_14761,N_12387);
nand U17422 (N_17422,N_15439,N_12103);
and U17423 (N_17423,N_14918,N_13032);
xnor U17424 (N_17424,N_13041,N_15978);
or U17425 (N_17425,N_12492,N_14566);
and U17426 (N_17426,N_14974,N_13587);
nand U17427 (N_17427,N_14678,N_13162);
nand U17428 (N_17428,N_15748,N_12438);
and U17429 (N_17429,N_13067,N_15190);
nor U17430 (N_17430,N_14060,N_14994);
and U17431 (N_17431,N_15718,N_12154);
xor U17432 (N_17432,N_13620,N_12840);
nor U17433 (N_17433,N_15828,N_12948);
and U17434 (N_17434,N_13209,N_13907);
nor U17435 (N_17435,N_14922,N_15035);
or U17436 (N_17436,N_13002,N_15144);
xor U17437 (N_17437,N_15975,N_15763);
nand U17438 (N_17438,N_15798,N_14168);
nand U17439 (N_17439,N_13696,N_14537);
and U17440 (N_17440,N_15192,N_14082);
and U17441 (N_17441,N_13934,N_12268);
or U17442 (N_17442,N_14595,N_13538);
nor U17443 (N_17443,N_15767,N_12429);
or U17444 (N_17444,N_13326,N_12239);
xor U17445 (N_17445,N_12187,N_15216);
or U17446 (N_17446,N_12421,N_12911);
and U17447 (N_17447,N_13355,N_14249);
xnor U17448 (N_17448,N_14194,N_12530);
and U17449 (N_17449,N_14967,N_12165);
xnor U17450 (N_17450,N_13129,N_12910);
nand U17451 (N_17451,N_12844,N_15286);
nand U17452 (N_17452,N_15100,N_14572);
and U17453 (N_17453,N_14414,N_14466);
nor U17454 (N_17454,N_14063,N_12557);
xor U17455 (N_17455,N_12527,N_12743);
nor U17456 (N_17456,N_13992,N_15841);
and U17457 (N_17457,N_12368,N_15363);
nor U17458 (N_17458,N_13264,N_14674);
nor U17459 (N_17459,N_13605,N_12883);
and U17460 (N_17460,N_13167,N_13240);
or U17461 (N_17461,N_13593,N_14410);
or U17462 (N_17462,N_12323,N_13641);
or U17463 (N_17463,N_13243,N_13216);
nor U17464 (N_17464,N_15716,N_15596);
xor U17465 (N_17465,N_13082,N_13031);
and U17466 (N_17466,N_14246,N_12758);
nand U17467 (N_17467,N_12416,N_14752);
or U17468 (N_17468,N_12932,N_15582);
and U17469 (N_17469,N_14978,N_12228);
and U17470 (N_17470,N_15316,N_14061);
or U17471 (N_17471,N_13945,N_14767);
nand U17472 (N_17472,N_13224,N_14518);
and U17473 (N_17473,N_15359,N_14281);
nand U17474 (N_17474,N_12151,N_13719);
nand U17475 (N_17475,N_14953,N_15158);
nor U17476 (N_17476,N_14049,N_12538);
nand U17477 (N_17477,N_12947,N_14920);
nor U17478 (N_17478,N_13771,N_15195);
or U17479 (N_17479,N_12510,N_14627);
nor U17480 (N_17480,N_14115,N_14440);
nand U17481 (N_17481,N_15319,N_15948);
nand U17482 (N_17482,N_12968,N_12725);
nor U17483 (N_17483,N_15204,N_13912);
nand U17484 (N_17484,N_13364,N_14133);
and U17485 (N_17485,N_15092,N_12969);
and U17486 (N_17486,N_15455,N_14651);
nor U17487 (N_17487,N_14193,N_12580);
nor U17488 (N_17488,N_13818,N_14753);
nor U17489 (N_17489,N_14824,N_13784);
nand U17490 (N_17490,N_14177,N_12072);
nor U17491 (N_17491,N_14870,N_13021);
nand U17492 (N_17492,N_12920,N_14102);
and U17493 (N_17493,N_14750,N_13081);
nand U17494 (N_17494,N_13391,N_13473);
nand U17495 (N_17495,N_14534,N_15953);
nand U17496 (N_17496,N_15782,N_12902);
nand U17497 (N_17497,N_13597,N_15745);
nor U17498 (N_17498,N_13555,N_15153);
and U17499 (N_17499,N_14553,N_14398);
and U17500 (N_17500,N_15560,N_13703);
nand U17501 (N_17501,N_12079,N_14707);
nand U17502 (N_17502,N_14773,N_13309);
or U17503 (N_17503,N_15946,N_13840);
and U17504 (N_17504,N_13650,N_15197);
nor U17505 (N_17505,N_13866,N_14166);
or U17506 (N_17506,N_14149,N_12587);
nor U17507 (N_17507,N_12148,N_13526);
nand U17508 (N_17508,N_14665,N_12748);
or U17509 (N_17509,N_13154,N_14486);
nor U17510 (N_17510,N_15093,N_14220);
nor U17511 (N_17511,N_15157,N_12385);
nand U17512 (N_17512,N_15184,N_15083);
or U17513 (N_17513,N_13058,N_15389);
nand U17514 (N_17514,N_13396,N_14826);
nand U17515 (N_17515,N_15627,N_12238);
or U17516 (N_17516,N_15015,N_13184);
xor U17517 (N_17517,N_12491,N_15404);
or U17518 (N_17518,N_12222,N_13023);
or U17519 (N_17519,N_14350,N_12084);
or U17520 (N_17520,N_15431,N_13035);
or U17521 (N_17521,N_14529,N_12107);
and U17522 (N_17522,N_13930,N_13358);
xor U17523 (N_17523,N_15218,N_14594);
nor U17524 (N_17524,N_14578,N_15565);
xor U17525 (N_17525,N_12426,N_12938);
and U17526 (N_17526,N_13741,N_12698);
nand U17527 (N_17527,N_14447,N_13377);
nor U17528 (N_17528,N_12078,N_14596);
xnor U17529 (N_17529,N_14563,N_12934);
and U17530 (N_17530,N_14831,N_15042);
nand U17531 (N_17531,N_14620,N_12795);
nor U17532 (N_17532,N_13084,N_13961);
nand U17533 (N_17533,N_14036,N_13731);
nor U17534 (N_17534,N_13443,N_15147);
xnor U17535 (N_17535,N_12265,N_13793);
nor U17536 (N_17536,N_12658,N_12496);
nor U17537 (N_17537,N_12001,N_14026);
xnor U17538 (N_17538,N_15445,N_12819);
xnor U17539 (N_17539,N_13960,N_15119);
nand U17540 (N_17540,N_14239,N_15853);
or U17541 (N_17541,N_12032,N_15919);
nand U17542 (N_17542,N_14420,N_14469);
and U17543 (N_17543,N_13869,N_12331);
nand U17544 (N_17544,N_12459,N_14641);
nand U17545 (N_17545,N_15629,N_12988);
and U17546 (N_17546,N_13659,N_12499);
nand U17547 (N_17547,N_13050,N_13221);
nor U17548 (N_17548,N_14120,N_13171);
and U17549 (N_17549,N_13361,N_13759);
nand U17550 (N_17550,N_12540,N_13861);
nand U17551 (N_17551,N_15688,N_15276);
or U17552 (N_17552,N_14349,N_13964);
nand U17553 (N_17553,N_13310,N_15449);
nand U17554 (N_17554,N_12681,N_14850);
xnor U17555 (N_17555,N_12793,N_15812);
or U17556 (N_17556,N_14122,N_12423);
and U17557 (N_17557,N_15435,N_12783);
nand U17558 (N_17558,N_13951,N_15166);
nor U17559 (N_17559,N_13841,N_15210);
xor U17560 (N_17560,N_12296,N_13854);
xnor U17561 (N_17561,N_14943,N_13426);
and U17562 (N_17562,N_13080,N_12669);
or U17563 (N_17563,N_13077,N_14297);
and U17564 (N_17564,N_14152,N_15212);
and U17565 (N_17565,N_15933,N_14562);
or U17566 (N_17566,N_14734,N_12644);
xnor U17567 (N_17567,N_14272,N_12117);
and U17568 (N_17568,N_13791,N_13384);
nor U17569 (N_17569,N_14647,N_13545);
or U17570 (N_17570,N_12571,N_14089);
nand U17571 (N_17571,N_13584,N_15546);
and U17572 (N_17572,N_14982,N_15795);
nor U17573 (N_17573,N_14119,N_14131);
nand U17574 (N_17574,N_13946,N_13270);
or U17575 (N_17575,N_15633,N_14388);
and U17576 (N_17576,N_14919,N_15644);
nand U17577 (N_17577,N_14533,N_14172);
nand U17578 (N_17578,N_14400,N_12086);
or U17579 (N_17579,N_14192,N_13296);
nor U17580 (N_17580,N_13692,N_14491);
xnor U17581 (N_17581,N_15930,N_13251);
or U17582 (N_17582,N_15338,N_15719);
nor U17583 (N_17583,N_12026,N_13137);
nor U17584 (N_17584,N_12829,N_13942);
and U17585 (N_17585,N_12269,N_13434);
nand U17586 (N_17586,N_14479,N_14747);
nor U17587 (N_17587,N_12058,N_13007);
nor U17588 (N_17588,N_13485,N_12556);
xor U17589 (N_17589,N_14386,N_15474);
or U17590 (N_17590,N_15757,N_15520);
nor U17591 (N_17591,N_13494,N_14201);
and U17592 (N_17592,N_13691,N_14204);
xor U17593 (N_17593,N_13130,N_15263);
nand U17594 (N_17594,N_15223,N_13441);
and U17595 (N_17595,N_14836,N_13140);
and U17596 (N_17596,N_14965,N_12473);
and U17597 (N_17597,N_12207,N_12100);
and U17598 (N_17598,N_13189,N_13739);
and U17599 (N_17599,N_14074,N_15208);
nand U17600 (N_17600,N_13738,N_14236);
nor U17601 (N_17601,N_15837,N_13225);
nand U17602 (N_17602,N_13110,N_12569);
nand U17603 (N_17603,N_12866,N_14996);
nand U17604 (N_17604,N_12746,N_12081);
and U17605 (N_17605,N_14737,N_15118);
xnor U17606 (N_17606,N_13161,N_12689);
or U17607 (N_17607,N_13578,N_13817);
nand U17608 (N_17608,N_12312,N_14078);
nand U17609 (N_17609,N_12971,N_15456);
nand U17610 (N_17610,N_15874,N_15968);
nand U17611 (N_17611,N_13967,N_12102);
and U17612 (N_17612,N_13891,N_13644);
or U17613 (N_17613,N_12694,N_12612);
or U17614 (N_17614,N_12573,N_14317);
nand U17615 (N_17615,N_13666,N_15160);
nor U17616 (N_17616,N_14987,N_12076);
xnor U17617 (N_17617,N_13351,N_13928);
and U17618 (N_17618,N_14717,N_13648);
nand U17619 (N_17619,N_13353,N_14866);
xnor U17620 (N_17620,N_15437,N_13338);
nor U17621 (N_17621,N_15770,N_14403);
nand U17622 (N_17622,N_14580,N_14813);
nand U17623 (N_17623,N_14214,N_15895);
nand U17624 (N_17624,N_14886,N_13522);
xnor U17625 (N_17625,N_13690,N_13646);
and U17626 (N_17626,N_13843,N_15793);
and U17627 (N_17627,N_14351,N_13017);
nand U17628 (N_17628,N_14406,N_15203);
or U17629 (N_17629,N_15154,N_12206);
or U17630 (N_17630,N_12005,N_15073);
or U17631 (N_17631,N_15162,N_13111);
or U17632 (N_17632,N_15304,N_13954);
or U17633 (N_17633,N_14962,N_14468);
nor U17634 (N_17634,N_14600,N_12734);
or U17635 (N_17635,N_15169,N_15740);
nand U17636 (N_17636,N_12012,N_13073);
nor U17637 (N_17637,N_13165,N_14667);
and U17638 (N_17638,N_15931,N_15866);
xor U17639 (N_17639,N_12147,N_13664);
and U17640 (N_17640,N_15973,N_13542);
nand U17641 (N_17641,N_15831,N_15730);
and U17642 (N_17642,N_13314,N_13255);
nand U17643 (N_17643,N_12630,N_13602);
or U17644 (N_17644,N_13794,N_13374);
nand U17645 (N_17645,N_15125,N_12092);
nor U17646 (N_17646,N_14508,N_14348);
and U17647 (N_17647,N_13090,N_14554);
nand U17648 (N_17648,N_15469,N_12645);
nand U17649 (N_17649,N_14338,N_14725);
and U17650 (N_17650,N_13634,N_15516);
or U17651 (N_17651,N_15220,N_13541);
and U17652 (N_17652,N_14772,N_14983);
nand U17653 (N_17653,N_15051,N_15998);
nor U17654 (N_17654,N_15881,N_12940);
nand U17655 (N_17655,N_15367,N_14396);
nor U17656 (N_17656,N_15385,N_14294);
or U17657 (N_17657,N_14147,N_12722);
nand U17658 (N_17658,N_12623,N_15927);
or U17659 (N_17659,N_12899,N_14090);
nand U17660 (N_17660,N_14659,N_13393);
and U17661 (N_17661,N_12132,N_14101);
nor U17662 (N_17662,N_15613,N_12674);
and U17663 (N_17663,N_14106,N_14941);
xor U17664 (N_17664,N_14488,N_14520);
or U17665 (N_17665,N_15540,N_15283);
or U17666 (N_17666,N_13506,N_14797);
and U17667 (N_17667,N_15243,N_12232);
nand U17668 (N_17668,N_14714,N_12564);
nand U17669 (N_17669,N_12957,N_12464);
and U17670 (N_17670,N_12686,N_15515);
nor U17671 (N_17671,N_12922,N_12756);
or U17672 (N_17672,N_15025,N_14358);
or U17673 (N_17673,N_15646,N_12826);
or U17674 (N_17674,N_14776,N_13439);
xor U17675 (N_17675,N_12320,N_15738);
or U17676 (N_17676,N_14443,N_13956);
nand U17677 (N_17677,N_12992,N_13892);
and U17678 (N_17678,N_12214,N_12818);
or U17679 (N_17679,N_15351,N_13989);
and U17680 (N_17680,N_12225,N_15290);
xor U17681 (N_17681,N_15994,N_12372);
nand U17682 (N_17682,N_12277,N_12115);
nand U17683 (N_17683,N_14721,N_13834);
nand U17684 (N_17684,N_14535,N_14360);
or U17685 (N_17685,N_13106,N_15781);
nor U17686 (N_17686,N_13839,N_15833);
or U17687 (N_17687,N_15137,N_12082);
nor U17688 (N_17688,N_12133,N_12871);
nand U17689 (N_17689,N_15656,N_13454);
nor U17690 (N_17690,N_15408,N_13342);
nor U17691 (N_17691,N_12045,N_13825);
or U17692 (N_17692,N_14279,N_14809);
xnor U17693 (N_17693,N_15246,N_14484);
or U17694 (N_17694,N_13913,N_13488);
nand U17695 (N_17695,N_13968,N_15390);
or U17696 (N_17696,N_13037,N_15366);
nand U17697 (N_17697,N_12720,N_12762);
xnor U17698 (N_17698,N_15129,N_12870);
nor U17699 (N_17699,N_13673,N_15291);
nand U17700 (N_17700,N_15788,N_15824);
nand U17701 (N_17701,N_14652,N_12614);
nor U17702 (N_17702,N_15602,N_14905);
or U17703 (N_17703,N_13344,N_13345);
and U17704 (N_17704,N_13206,N_14248);
nand U17705 (N_17705,N_13550,N_15751);
or U17706 (N_17706,N_15369,N_14392);
nand U17707 (N_17707,N_15446,N_12546);
nor U17708 (N_17708,N_15348,N_12025);
xor U17709 (N_17709,N_13490,N_12691);
xor U17710 (N_17710,N_14673,N_13525);
nor U17711 (N_17711,N_15696,N_15723);
xor U17712 (N_17712,N_15268,N_13214);
and U17713 (N_17713,N_13267,N_15622);
nand U17714 (N_17714,N_15590,N_14365);
and U17715 (N_17715,N_14527,N_15403);
nor U17716 (N_17716,N_14669,N_14538);
or U17717 (N_17717,N_15589,N_15807);
and U17718 (N_17718,N_12842,N_12554);
nand U17719 (N_17719,N_14190,N_15133);
nand U17720 (N_17720,N_13220,N_14906);
or U17721 (N_17721,N_13159,N_15766);
nor U17722 (N_17722,N_14110,N_13420);
nor U17723 (N_17723,N_15556,N_14215);
nand U17724 (N_17724,N_14867,N_14212);
nand U17725 (N_17725,N_12390,N_12760);
and U17726 (N_17726,N_12241,N_15869);
or U17727 (N_17727,N_15378,N_15014);
xnor U17728 (N_17728,N_15062,N_14371);
or U17729 (N_17729,N_13440,N_14583);
and U17730 (N_17730,N_13191,N_15260);
nand U17731 (N_17731,N_14291,N_14470);
and U17732 (N_17732,N_15481,N_13875);
and U17733 (N_17733,N_15611,N_15322);
nor U17734 (N_17734,N_13211,N_14043);
nor U17735 (N_17735,N_13543,N_14904);
nor U17736 (N_17736,N_15660,N_12673);
nor U17737 (N_17737,N_14525,N_13642);
and U17738 (N_17738,N_14602,N_13078);
and U17739 (N_17739,N_14135,N_13010);
xor U17740 (N_17740,N_14648,N_12802);
and U17741 (N_17741,N_13053,N_13625);
and U17742 (N_17742,N_13828,N_12607);
nor U17743 (N_17743,N_12912,N_12621);
nand U17744 (N_17744,N_13481,N_12824);
and U17745 (N_17745,N_13631,N_13614);
nor U17746 (N_17746,N_14869,N_15671);
nor U17747 (N_17747,N_14512,N_14699);
and U17748 (N_17748,N_12638,N_14507);
nor U17749 (N_17749,N_15814,N_15510);
or U17750 (N_17750,N_13684,N_13635);
or U17751 (N_17751,N_14415,N_12796);
nand U17752 (N_17752,N_14307,N_13316);
or U17753 (N_17753,N_12581,N_15863);
xnor U17754 (N_17754,N_12927,N_12108);
nand U17755 (N_17755,N_15084,N_13116);
nor U17756 (N_17756,N_14111,N_14860);
and U17757 (N_17757,N_12209,N_13877);
and U17758 (N_17758,N_14799,N_13476);
and U17759 (N_17759,N_12772,N_14432);
nor U17760 (N_17760,N_14366,N_13113);
and U17761 (N_17761,N_14027,N_12089);
xor U17762 (N_17762,N_15654,N_13711);
or U17763 (N_17763,N_12374,N_14837);
or U17764 (N_17764,N_12248,N_14645);
nand U17765 (N_17765,N_13904,N_14949);
nor U17766 (N_17766,N_13394,N_14788);
and U17767 (N_17767,N_14712,N_12069);
or U17768 (N_17768,N_13598,N_12972);
xnor U17769 (N_17769,N_14924,N_13916);
xor U17770 (N_17770,N_14832,N_15006);
and U17771 (N_17771,N_13483,N_13104);
xnor U17772 (N_17772,N_12091,N_14785);
nor U17773 (N_17773,N_15349,N_15972);
and U17774 (N_17774,N_14232,N_14118);
or U17775 (N_17775,N_14804,N_15618);
and U17776 (N_17776,N_15725,N_14211);
xor U17777 (N_17777,N_12318,N_13218);
and U17778 (N_17778,N_12270,N_15278);
xor U17779 (N_17779,N_15089,N_12453);
and U17780 (N_17780,N_14446,N_12981);
and U17781 (N_17781,N_15789,N_15893);
or U17782 (N_17782,N_13761,N_13115);
nand U17783 (N_17783,N_13418,N_14865);
and U17784 (N_17784,N_12451,N_12798);
nand U17785 (N_17785,N_13952,N_12467);
or U17786 (N_17786,N_14874,N_12853);
nor U17787 (N_17787,N_14901,N_15381);
nand U17788 (N_17788,N_15902,N_13534);
and U17789 (N_17789,N_12519,N_12112);
and U17790 (N_17790,N_12717,N_14811);
nor U17791 (N_17791,N_12176,N_13144);
nand U17792 (N_17792,N_12441,N_15193);
or U17793 (N_17793,N_14782,N_14812);
nand U17794 (N_17794,N_14827,N_12192);
and U17795 (N_17795,N_15908,N_12542);
xnor U17796 (N_17796,N_15772,N_14278);
nor U17797 (N_17797,N_15031,N_13306);
or U17798 (N_17798,N_12715,N_13288);
or U17799 (N_17799,N_12403,N_14688);
or U17800 (N_17800,N_12461,N_15989);
or U17801 (N_17801,N_14539,N_12477);
and U17802 (N_17802,N_14353,N_15768);
and U17803 (N_17803,N_13233,N_13756);
nor U17804 (N_17804,N_13088,N_12063);
nor U17805 (N_17805,N_12283,N_12690);
and U17806 (N_17806,N_13778,N_13733);
or U17807 (N_17807,N_12984,N_13284);
or U17808 (N_17808,N_15701,N_14424);
nand U17809 (N_17809,N_15081,N_13977);
nor U17810 (N_17810,N_15156,N_14705);
nand U17811 (N_17811,N_13590,N_12336);
or U17812 (N_17812,N_12961,N_14735);
and U17813 (N_17813,N_14071,N_14859);
xor U17814 (N_17814,N_15229,N_15113);
nor U17815 (N_17815,N_15794,N_15586);
and U17816 (N_17816,N_13433,N_14697);
nand U17817 (N_17817,N_12481,N_14265);
nand U17818 (N_17818,N_15928,N_14644);
and U17819 (N_17819,N_15985,N_15331);
or U17820 (N_17820,N_12549,N_13019);
and U17821 (N_17821,N_15383,N_15067);
and U17822 (N_17822,N_14324,N_15652);
xor U17823 (N_17823,N_13718,N_13515);
nor U17824 (N_17824,N_15801,N_13236);
nand U17825 (N_17825,N_13988,N_12733);
nor U17826 (N_17826,N_15247,N_12337);
or U17827 (N_17827,N_15917,N_13868);
or U17828 (N_17828,N_15692,N_15198);
or U17829 (N_17829,N_12550,N_13484);
and U17830 (N_17830,N_14355,N_15784);
nor U17831 (N_17831,N_12754,N_12839);
nand U17832 (N_17832,N_12711,N_13185);
and U17833 (N_17833,N_14148,N_12126);
nor U17834 (N_17834,N_13881,N_15672);
nor U17835 (N_17835,N_12216,N_12399);
nand U17836 (N_17836,N_14087,N_13242);
nor U17837 (N_17837,N_12635,N_14409);
and U17838 (N_17838,N_14957,N_15353);
nor U17839 (N_17839,N_13287,N_15061);
nor U17840 (N_17840,N_13172,N_12869);
or U17841 (N_17841,N_12503,N_13471);
nor U17842 (N_17842,N_13482,N_15584);
nand U17843 (N_17843,N_13156,N_12049);
xnor U17844 (N_17844,N_14732,N_15579);
nand U17845 (N_17845,N_13331,N_14009);
or U17846 (N_17846,N_14170,N_14451);
and U17847 (N_17847,N_15739,N_15175);
and U17848 (N_17848,N_12309,N_13413);
or U17849 (N_17849,N_12410,N_12767);
and U17850 (N_17850,N_15373,N_12590);
nor U17851 (N_17851,N_14197,N_14066);
and U17852 (N_17852,N_14487,N_15704);
or U17853 (N_17853,N_13507,N_15047);
and U17854 (N_17854,N_15108,N_15040);
or U17855 (N_17855,N_12475,N_12469);
and U17856 (N_17856,N_12430,N_14570);
xnor U17857 (N_17857,N_12647,N_12785);
and U17858 (N_17858,N_13480,N_15386);
and U17859 (N_17859,N_12257,N_12261);
or U17860 (N_17860,N_13011,N_14981);
nand U17861 (N_17861,N_14080,N_12215);
or U17862 (N_17862,N_13186,N_14598);
nand U17863 (N_17863,N_14295,N_12035);
or U17864 (N_17864,N_15884,N_12376);
xor U17865 (N_17865,N_14980,N_15070);
xnor U17866 (N_17866,N_13128,N_14935);
nor U17867 (N_17867,N_13827,N_14391);
and U17868 (N_17868,N_14908,N_15301);
or U17869 (N_17869,N_15585,N_14187);
nand U17870 (N_17870,N_15421,N_14116);
nor U17871 (N_17871,N_15228,N_12067);
and U17872 (N_17872,N_14428,N_14561);
nor U17873 (N_17873,N_15111,N_12396);
nor U17874 (N_17874,N_14312,N_12436);
xor U17875 (N_17875,N_15531,N_13341);
and U17876 (N_17876,N_15750,N_12603);
or U17877 (N_17877,N_15498,N_13979);
and U17878 (N_17878,N_13260,N_13109);
or U17879 (N_17879,N_13327,N_14434);
nor U17880 (N_17880,N_12114,N_14840);
and U17881 (N_17881,N_15310,N_12194);
or U17882 (N_17882,N_13387,N_14020);
nand U17883 (N_17883,N_13874,N_12064);
and U17884 (N_17884,N_14708,N_14364);
and U17885 (N_17885,N_15550,N_13911);
nor U17886 (N_17886,N_15761,N_13789);
or U17887 (N_17887,N_12943,N_15308);
xor U17888 (N_17888,N_14323,N_13145);
nor U17889 (N_17889,N_15779,N_13591);
or U17890 (N_17890,N_13092,N_13857);
nor U17891 (N_17891,N_15368,N_12130);
xor U17892 (N_17892,N_12685,N_15036);
and U17893 (N_17893,N_15594,N_13565);
nand U17894 (N_17894,N_15476,N_12213);
or U17895 (N_17895,N_13630,N_13845);
nand U17896 (N_17896,N_12889,N_12930);
nor U17897 (N_17897,N_15947,N_12808);
nor U17898 (N_17898,N_14709,N_12042);
and U17899 (N_17899,N_15026,N_13103);
or U17900 (N_17900,N_12805,N_12731);
xor U17901 (N_17901,N_13241,N_15679);
nand U17902 (N_17902,N_12747,N_15189);
and U17903 (N_17903,N_14024,N_15856);
nand U17904 (N_17904,N_12218,N_15284);
nand U17905 (N_17905,N_14408,N_15600);
or U17906 (N_17906,N_15277,N_13772);
xor U17907 (N_17907,N_13386,N_12263);
nor U17908 (N_17908,N_15182,N_12729);
and U17909 (N_17909,N_15085,N_15775);
nand U17910 (N_17910,N_12979,N_13423);
nand U17911 (N_17911,N_15013,N_13757);
nand U17912 (N_17912,N_12332,N_13689);
and U17913 (N_17913,N_14490,N_15747);
or U17914 (N_17914,N_12545,N_15659);
nand U17915 (N_17915,N_15487,N_12249);
or U17916 (N_17916,N_13783,N_14792);
nor U17917 (N_17917,N_14989,N_12775);
nor U17918 (N_17918,N_14742,N_14614);
or U17919 (N_17919,N_13043,N_13665);
and U17920 (N_17920,N_15601,N_13637);
nor U17921 (N_17921,N_15295,N_15294);
nor U17922 (N_17922,N_14692,N_12983);
nor U17923 (N_17923,N_12875,N_12022);
and U17924 (N_17924,N_13381,N_13020);
and U17925 (N_17925,N_13616,N_14661);
or U17926 (N_17926,N_15785,N_12936);
nand U17927 (N_17927,N_14032,N_12985);
nor U17928 (N_17928,N_12878,N_12247);
nor U17929 (N_17929,N_14745,N_15810);
and U17930 (N_17930,N_13348,N_15149);
xor U17931 (N_17931,N_13901,N_15823);
nor U17932 (N_17932,N_14899,N_14431);
and U17933 (N_17933,N_12917,N_12977);
or U17934 (N_17934,N_14485,N_12626);
and U17935 (N_17935,N_14948,N_15096);
nand U17936 (N_17936,N_14830,N_12060);
or U17937 (N_17937,N_13100,N_15666);
and U17938 (N_17938,N_14482,N_13231);
nand U17939 (N_17939,N_14005,N_13669);
nand U17940 (N_17940,N_15231,N_13588);
and U17941 (N_17941,N_12655,N_15027);
nand U17942 (N_17942,N_14564,N_15780);
nand U17943 (N_17943,N_13905,N_13547);
xnor U17944 (N_17944,N_12041,N_13277);
nand U17945 (N_17945,N_13455,N_12411);
or U17946 (N_17946,N_12755,N_13045);
nand U17947 (N_17947,N_15401,N_14787);
nand U17948 (N_17948,N_12389,N_14385);
and U17949 (N_17949,N_14407,N_12242);
and U17950 (N_17950,N_15141,N_14789);
nand U17951 (N_17951,N_12170,N_14587);
and U17952 (N_17952,N_14821,N_14019);
nand U17953 (N_17953,N_15132,N_12245);
nor U17954 (N_17954,N_14225,N_15787);
nand U17955 (N_17955,N_12171,N_15271);
nor U17956 (N_17956,N_12776,N_12736);
nor U17957 (N_17957,N_13878,N_12873);
xor U17958 (N_17958,N_14134,N_12488);
and U17959 (N_17959,N_14658,N_15405);
nor U17960 (N_17960,N_15285,N_13285);
nor U17961 (N_17961,N_13937,N_12885);
or U17962 (N_17962,N_15826,N_15237);
and U17963 (N_17963,N_12593,N_14691);
or U17964 (N_17964,N_14675,N_12359);
nand U17965 (N_17965,N_13564,N_14359);
xnor U17966 (N_17966,N_13057,N_14896);
or U17967 (N_17967,N_12951,N_12953);
and U17968 (N_17968,N_14105,N_13885);
nand U17969 (N_17969,N_15380,N_14315);
nand U17970 (N_17970,N_14713,N_14536);
or U17971 (N_17971,N_12786,N_14629);
nand U17972 (N_17972,N_15867,N_13204);
or U17973 (N_17973,N_15695,N_12652);
nor U17974 (N_17974,N_14754,N_15360);
or U17975 (N_17975,N_12737,N_13667);
and U17976 (N_17976,N_13926,N_15914);
and U17977 (N_17977,N_13312,N_13600);
xor U17978 (N_17978,N_12646,N_14495);
nand U17979 (N_17979,N_14740,N_13289);
or U17980 (N_17980,N_15344,N_14402);
or U17981 (N_17981,N_13985,N_15762);
xor U17982 (N_17982,N_13813,N_15249);
and U17983 (N_17983,N_13585,N_15506);
and U17984 (N_17984,N_14511,N_13548);
or U17985 (N_17985,N_13119,N_15997);
nor U17986 (N_17986,N_14964,N_15462);
nor U17987 (N_17987,N_15058,N_12204);
nor U17988 (N_17988,N_13842,N_13205);
nor U17989 (N_17989,N_13816,N_15262);
or U17990 (N_17990,N_13373,N_14802);
or U17991 (N_17991,N_14857,N_14963);
nor U17992 (N_17992,N_13727,N_15493);
xor U17993 (N_17993,N_15942,N_15758);
and U17994 (N_17994,N_13329,N_15699);
nand U17995 (N_17995,N_13495,N_14022);
and U17996 (N_17996,N_15517,N_14718);
nor U17997 (N_17997,N_14097,N_15712);
nor U17998 (N_17998,N_13026,N_12896);
nand U17999 (N_17999,N_12615,N_13982);
or U18000 (N_18000,N_12833,N_15201);
and U18001 (N_18001,N_12161,N_14269);
and U18002 (N_18002,N_13557,N_12222);
nand U18003 (N_18003,N_14934,N_15816);
or U18004 (N_18004,N_13197,N_13155);
and U18005 (N_18005,N_15792,N_15398);
nor U18006 (N_18006,N_15831,N_15023);
nor U18007 (N_18007,N_13529,N_12149);
nor U18008 (N_18008,N_12306,N_15735);
nand U18009 (N_18009,N_15910,N_15069);
and U18010 (N_18010,N_14130,N_13918);
and U18011 (N_18011,N_15343,N_12665);
xor U18012 (N_18012,N_14448,N_15061);
nor U18013 (N_18013,N_13269,N_15449);
nand U18014 (N_18014,N_14136,N_13114);
and U18015 (N_18015,N_13131,N_15927);
nor U18016 (N_18016,N_15371,N_13799);
and U18017 (N_18017,N_13672,N_15178);
or U18018 (N_18018,N_12684,N_13412);
and U18019 (N_18019,N_13321,N_12401);
and U18020 (N_18020,N_14193,N_13547);
xnor U18021 (N_18021,N_13304,N_15937);
nor U18022 (N_18022,N_14255,N_14031);
nand U18023 (N_18023,N_14622,N_12692);
nand U18024 (N_18024,N_13198,N_13105);
nand U18025 (N_18025,N_13953,N_12362);
nand U18026 (N_18026,N_13550,N_14326);
nor U18027 (N_18027,N_12406,N_13750);
nand U18028 (N_18028,N_13535,N_15119);
nand U18029 (N_18029,N_13039,N_14678);
nand U18030 (N_18030,N_15872,N_13374);
xor U18031 (N_18031,N_15741,N_14423);
and U18032 (N_18032,N_12428,N_12579);
nor U18033 (N_18033,N_13458,N_12053);
or U18034 (N_18034,N_14403,N_15148);
xnor U18035 (N_18035,N_12799,N_15141);
or U18036 (N_18036,N_13157,N_14954);
and U18037 (N_18037,N_14650,N_15011);
and U18038 (N_18038,N_12698,N_14458);
nand U18039 (N_18039,N_14536,N_12814);
nand U18040 (N_18040,N_12025,N_14350);
or U18041 (N_18041,N_14247,N_13861);
nand U18042 (N_18042,N_12803,N_13877);
nor U18043 (N_18043,N_13602,N_13450);
nand U18044 (N_18044,N_15551,N_13569);
nor U18045 (N_18045,N_13655,N_14717);
and U18046 (N_18046,N_12184,N_15629);
nor U18047 (N_18047,N_12104,N_13120);
and U18048 (N_18048,N_14594,N_13861);
nand U18049 (N_18049,N_13605,N_14166);
and U18050 (N_18050,N_12246,N_14766);
nand U18051 (N_18051,N_14627,N_14813);
nor U18052 (N_18052,N_12676,N_12163);
nand U18053 (N_18053,N_13647,N_14912);
xnor U18054 (N_18054,N_12732,N_15396);
or U18055 (N_18055,N_14279,N_13373);
nand U18056 (N_18056,N_14459,N_14106);
and U18057 (N_18057,N_12107,N_15905);
and U18058 (N_18058,N_15879,N_12649);
nor U18059 (N_18059,N_13849,N_12073);
nor U18060 (N_18060,N_12038,N_13059);
nand U18061 (N_18061,N_14991,N_13107);
nor U18062 (N_18062,N_13007,N_13123);
or U18063 (N_18063,N_13570,N_12050);
nand U18064 (N_18064,N_15070,N_12944);
or U18065 (N_18065,N_12458,N_15587);
or U18066 (N_18066,N_14814,N_15040);
nand U18067 (N_18067,N_14070,N_13650);
xnor U18068 (N_18068,N_15292,N_15583);
and U18069 (N_18069,N_14877,N_14279);
or U18070 (N_18070,N_15119,N_15352);
and U18071 (N_18071,N_12484,N_15461);
or U18072 (N_18072,N_12728,N_15948);
and U18073 (N_18073,N_12899,N_14518);
nand U18074 (N_18074,N_13626,N_15502);
nand U18075 (N_18075,N_15791,N_12894);
nand U18076 (N_18076,N_13792,N_13646);
nand U18077 (N_18077,N_13347,N_12115);
nand U18078 (N_18078,N_15083,N_12001);
nand U18079 (N_18079,N_12364,N_15670);
or U18080 (N_18080,N_12929,N_14232);
nand U18081 (N_18081,N_14653,N_12340);
or U18082 (N_18082,N_12956,N_14546);
xnor U18083 (N_18083,N_13090,N_15692);
or U18084 (N_18084,N_13782,N_12479);
nand U18085 (N_18085,N_14047,N_12847);
and U18086 (N_18086,N_14167,N_15900);
and U18087 (N_18087,N_13229,N_13147);
nor U18088 (N_18088,N_15955,N_14618);
xnor U18089 (N_18089,N_12870,N_13588);
nor U18090 (N_18090,N_15964,N_14674);
or U18091 (N_18091,N_12051,N_12918);
and U18092 (N_18092,N_15378,N_15478);
nand U18093 (N_18093,N_15173,N_14326);
nor U18094 (N_18094,N_12634,N_12530);
nand U18095 (N_18095,N_12171,N_13583);
or U18096 (N_18096,N_15539,N_15530);
nor U18097 (N_18097,N_14302,N_14432);
nor U18098 (N_18098,N_13093,N_15864);
or U18099 (N_18099,N_13421,N_13182);
or U18100 (N_18100,N_12376,N_13535);
or U18101 (N_18101,N_12674,N_12213);
nand U18102 (N_18102,N_15458,N_15304);
and U18103 (N_18103,N_13459,N_12100);
xor U18104 (N_18104,N_12900,N_12053);
xnor U18105 (N_18105,N_15377,N_12820);
nand U18106 (N_18106,N_13871,N_14373);
or U18107 (N_18107,N_12997,N_15426);
nand U18108 (N_18108,N_15834,N_13446);
nand U18109 (N_18109,N_12532,N_15307);
nand U18110 (N_18110,N_12257,N_15953);
and U18111 (N_18111,N_12403,N_15114);
nand U18112 (N_18112,N_12693,N_12234);
nand U18113 (N_18113,N_12268,N_15195);
or U18114 (N_18114,N_14982,N_13300);
nand U18115 (N_18115,N_12702,N_15227);
and U18116 (N_18116,N_15691,N_14996);
nand U18117 (N_18117,N_12921,N_14959);
nand U18118 (N_18118,N_12642,N_15091);
or U18119 (N_18119,N_13831,N_12828);
nand U18120 (N_18120,N_15208,N_12304);
nor U18121 (N_18121,N_13676,N_15479);
nor U18122 (N_18122,N_13606,N_13153);
and U18123 (N_18123,N_12266,N_14537);
or U18124 (N_18124,N_12878,N_15416);
nor U18125 (N_18125,N_12114,N_12388);
nor U18126 (N_18126,N_12577,N_15797);
nor U18127 (N_18127,N_13018,N_12396);
xor U18128 (N_18128,N_15010,N_14449);
xor U18129 (N_18129,N_13158,N_15765);
nor U18130 (N_18130,N_13098,N_14232);
nor U18131 (N_18131,N_12653,N_14643);
nor U18132 (N_18132,N_15083,N_14185);
and U18133 (N_18133,N_14964,N_13643);
nor U18134 (N_18134,N_12514,N_13287);
nand U18135 (N_18135,N_12913,N_15452);
nor U18136 (N_18136,N_15002,N_12258);
xnor U18137 (N_18137,N_13551,N_15160);
nor U18138 (N_18138,N_15663,N_12840);
nand U18139 (N_18139,N_12348,N_13079);
or U18140 (N_18140,N_12483,N_14272);
and U18141 (N_18141,N_15022,N_14630);
nor U18142 (N_18142,N_13023,N_14980);
nand U18143 (N_18143,N_14600,N_12128);
and U18144 (N_18144,N_13403,N_14911);
and U18145 (N_18145,N_13075,N_12171);
nor U18146 (N_18146,N_14215,N_14625);
nand U18147 (N_18147,N_15457,N_12385);
nand U18148 (N_18148,N_15324,N_15667);
nand U18149 (N_18149,N_15128,N_12803);
xnor U18150 (N_18150,N_14066,N_15785);
and U18151 (N_18151,N_15856,N_12141);
and U18152 (N_18152,N_15907,N_14304);
and U18153 (N_18153,N_15599,N_14952);
or U18154 (N_18154,N_12254,N_13695);
nor U18155 (N_18155,N_12599,N_15382);
nor U18156 (N_18156,N_13468,N_13534);
nand U18157 (N_18157,N_15413,N_12132);
and U18158 (N_18158,N_12937,N_14737);
or U18159 (N_18159,N_13254,N_12017);
and U18160 (N_18160,N_15304,N_15003);
or U18161 (N_18161,N_12006,N_13609);
nand U18162 (N_18162,N_12085,N_15630);
and U18163 (N_18163,N_15352,N_12425);
nor U18164 (N_18164,N_14603,N_13614);
nand U18165 (N_18165,N_12487,N_12576);
nor U18166 (N_18166,N_15071,N_15298);
nor U18167 (N_18167,N_13346,N_13979);
nor U18168 (N_18168,N_12297,N_15285);
or U18169 (N_18169,N_13822,N_13048);
or U18170 (N_18170,N_12494,N_13568);
nor U18171 (N_18171,N_13549,N_15444);
nand U18172 (N_18172,N_12793,N_15978);
and U18173 (N_18173,N_12069,N_13517);
nor U18174 (N_18174,N_13620,N_12919);
xor U18175 (N_18175,N_13252,N_12769);
or U18176 (N_18176,N_15293,N_12638);
or U18177 (N_18177,N_12227,N_12594);
nor U18178 (N_18178,N_12727,N_15244);
and U18179 (N_18179,N_12958,N_15794);
and U18180 (N_18180,N_13730,N_12475);
and U18181 (N_18181,N_15407,N_14663);
nor U18182 (N_18182,N_13323,N_15390);
and U18183 (N_18183,N_15010,N_13583);
nand U18184 (N_18184,N_12651,N_15370);
and U18185 (N_18185,N_13917,N_13878);
nor U18186 (N_18186,N_12925,N_12167);
and U18187 (N_18187,N_15929,N_15890);
nor U18188 (N_18188,N_12312,N_13628);
or U18189 (N_18189,N_15713,N_12464);
nor U18190 (N_18190,N_14816,N_13481);
and U18191 (N_18191,N_13476,N_12951);
or U18192 (N_18192,N_14787,N_15774);
nand U18193 (N_18193,N_13029,N_13671);
nor U18194 (N_18194,N_12630,N_13751);
nand U18195 (N_18195,N_15206,N_12052);
or U18196 (N_18196,N_15262,N_12892);
and U18197 (N_18197,N_15389,N_12265);
or U18198 (N_18198,N_12709,N_14771);
nor U18199 (N_18199,N_12180,N_14170);
nand U18200 (N_18200,N_14157,N_15894);
nor U18201 (N_18201,N_13868,N_13006);
nor U18202 (N_18202,N_13111,N_12216);
and U18203 (N_18203,N_12092,N_14288);
nor U18204 (N_18204,N_14569,N_13786);
or U18205 (N_18205,N_13175,N_12678);
and U18206 (N_18206,N_13809,N_15157);
or U18207 (N_18207,N_12933,N_13656);
nand U18208 (N_18208,N_14532,N_12047);
or U18209 (N_18209,N_12768,N_12153);
xor U18210 (N_18210,N_14948,N_12239);
nand U18211 (N_18211,N_15721,N_12220);
or U18212 (N_18212,N_15298,N_13945);
or U18213 (N_18213,N_12108,N_14071);
nand U18214 (N_18214,N_13410,N_12025);
nand U18215 (N_18215,N_13952,N_15350);
and U18216 (N_18216,N_14161,N_15099);
or U18217 (N_18217,N_12864,N_15346);
and U18218 (N_18218,N_15270,N_14356);
nor U18219 (N_18219,N_14178,N_13043);
nand U18220 (N_18220,N_14386,N_12398);
or U18221 (N_18221,N_13132,N_12382);
nor U18222 (N_18222,N_15312,N_12641);
and U18223 (N_18223,N_13376,N_12838);
nand U18224 (N_18224,N_15053,N_14938);
or U18225 (N_18225,N_14272,N_15805);
nand U18226 (N_18226,N_13244,N_12036);
nand U18227 (N_18227,N_15903,N_15945);
xnor U18228 (N_18228,N_14766,N_15765);
or U18229 (N_18229,N_13178,N_12335);
xor U18230 (N_18230,N_12701,N_12869);
nand U18231 (N_18231,N_13254,N_14630);
and U18232 (N_18232,N_15122,N_15558);
and U18233 (N_18233,N_15582,N_15401);
or U18234 (N_18234,N_14891,N_13585);
nand U18235 (N_18235,N_15075,N_15291);
and U18236 (N_18236,N_13445,N_13950);
nor U18237 (N_18237,N_12145,N_15923);
or U18238 (N_18238,N_15301,N_15604);
and U18239 (N_18239,N_13139,N_14749);
nand U18240 (N_18240,N_13862,N_12847);
and U18241 (N_18241,N_14971,N_12345);
nand U18242 (N_18242,N_13507,N_12109);
and U18243 (N_18243,N_14714,N_13763);
xnor U18244 (N_18244,N_15384,N_12069);
or U18245 (N_18245,N_15151,N_15723);
and U18246 (N_18246,N_14884,N_14534);
or U18247 (N_18247,N_12163,N_12232);
xor U18248 (N_18248,N_15213,N_15798);
and U18249 (N_18249,N_14408,N_14944);
or U18250 (N_18250,N_12282,N_14895);
nand U18251 (N_18251,N_14899,N_13008);
nand U18252 (N_18252,N_13329,N_15890);
or U18253 (N_18253,N_12752,N_15867);
nor U18254 (N_18254,N_15199,N_12794);
or U18255 (N_18255,N_15316,N_12610);
nor U18256 (N_18256,N_12021,N_12339);
and U18257 (N_18257,N_13808,N_13261);
or U18258 (N_18258,N_12469,N_12509);
nand U18259 (N_18259,N_15520,N_14252);
nand U18260 (N_18260,N_14935,N_13131);
and U18261 (N_18261,N_15083,N_14080);
xnor U18262 (N_18262,N_15366,N_13152);
nand U18263 (N_18263,N_14789,N_12838);
or U18264 (N_18264,N_15937,N_12999);
and U18265 (N_18265,N_13982,N_14699);
and U18266 (N_18266,N_14616,N_12592);
nor U18267 (N_18267,N_13676,N_14778);
or U18268 (N_18268,N_15195,N_14685);
or U18269 (N_18269,N_14384,N_14655);
or U18270 (N_18270,N_14566,N_15530);
nor U18271 (N_18271,N_14361,N_14702);
and U18272 (N_18272,N_13914,N_15980);
and U18273 (N_18273,N_15881,N_15765);
or U18274 (N_18274,N_14948,N_14871);
nand U18275 (N_18275,N_15197,N_14384);
nor U18276 (N_18276,N_14483,N_15833);
and U18277 (N_18277,N_12065,N_12276);
or U18278 (N_18278,N_15398,N_14832);
or U18279 (N_18279,N_12312,N_15740);
and U18280 (N_18280,N_12320,N_14927);
nor U18281 (N_18281,N_12653,N_13866);
xor U18282 (N_18282,N_15201,N_14558);
nor U18283 (N_18283,N_14689,N_14475);
and U18284 (N_18284,N_14480,N_13330);
or U18285 (N_18285,N_13848,N_13231);
nand U18286 (N_18286,N_14378,N_14833);
and U18287 (N_18287,N_14166,N_13701);
xnor U18288 (N_18288,N_14654,N_15730);
or U18289 (N_18289,N_12228,N_14705);
and U18290 (N_18290,N_13704,N_14089);
nor U18291 (N_18291,N_13272,N_14311);
nor U18292 (N_18292,N_15546,N_15963);
xnor U18293 (N_18293,N_13803,N_13031);
xnor U18294 (N_18294,N_15298,N_12058);
nor U18295 (N_18295,N_13537,N_13969);
nor U18296 (N_18296,N_13057,N_13572);
or U18297 (N_18297,N_13766,N_12403);
nand U18298 (N_18298,N_14721,N_14867);
or U18299 (N_18299,N_14806,N_15282);
nor U18300 (N_18300,N_13199,N_15592);
xnor U18301 (N_18301,N_13510,N_14661);
nand U18302 (N_18302,N_15830,N_14926);
and U18303 (N_18303,N_14264,N_13810);
nor U18304 (N_18304,N_12151,N_12698);
nand U18305 (N_18305,N_13215,N_13678);
nor U18306 (N_18306,N_13403,N_12760);
and U18307 (N_18307,N_14454,N_12299);
nor U18308 (N_18308,N_15090,N_12053);
xor U18309 (N_18309,N_13784,N_12894);
or U18310 (N_18310,N_15433,N_13471);
or U18311 (N_18311,N_15032,N_14872);
and U18312 (N_18312,N_15058,N_12250);
xor U18313 (N_18313,N_13416,N_13788);
or U18314 (N_18314,N_15627,N_12524);
nor U18315 (N_18315,N_13286,N_13082);
and U18316 (N_18316,N_14798,N_15994);
nand U18317 (N_18317,N_12461,N_14506);
nand U18318 (N_18318,N_15708,N_14479);
nand U18319 (N_18319,N_15147,N_15993);
and U18320 (N_18320,N_12868,N_12561);
xnor U18321 (N_18321,N_14077,N_13030);
or U18322 (N_18322,N_13601,N_12317);
nand U18323 (N_18323,N_13798,N_14638);
xor U18324 (N_18324,N_12784,N_15484);
and U18325 (N_18325,N_12972,N_12047);
nand U18326 (N_18326,N_15670,N_15392);
nand U18327 (N_18327,N_15964,N_13124);
nor U18328 (N_18328,N_14217,N_15981);
and U18329 (N_18329,N_12565,N_14358);
nand U18330 (N_18330,N_15607,N_15784);
nand U18331 (N_18331,N_15926,N_15549);
or U18332 (N_18332,N_13348,N_15202);
nand U18333 (N_18333,N_15719,N_12925);
or U18334 (N_18334,N_12466,N_14097);
nor U18335 (N_18335,N_15697,N_12452);
nor U18336 (N_18336,N_14506,N_15087);
and U18337 (N_18337,N_13565,N_13488);
nand U18338 (N_18338,N_12496,N_14435);
or U18339 (N_18339,N_14681,N_13580);
nand U18340 (N_18340,N_12877,N_14104);
xnor U18341 (N_18341,N_15107,N_15650);
nand U18342 (N_18342,N_13366,N_12562);
or U18343 (N_18343,N_12629,N_13093);
xor U18344 (N_18344,N_12666,N_14252);
or U18345 (N_18345,N_15607,N_12109);
nand U18346 (N_18346,N_12607,N_14603);
and U18347 (N_18347,N_12659,N_15608);
or U18348 (N_18348,N_14039,N_12907);
or U18349 (N_18349,N_14925,N_14527);
nor U18350 (N_18350,N_13902,N_15966);
nand U18351 (N_18351,N_15883,N_14801);
and U18352 (N_18352,N_15901,N_15612);
and U18353 (N_18353,N_14662,N_14824);
nor U18354 (N_18354,N_14256,N_12452);
xnor U18355 (N_18355,N_13308,N_12004);
nand U18356 (N_18356,N_12419,N_13352);
nor U18357 (N_18357,N_15855,N_14175);
and U18358 (N_18358,N_15348,N_12072);
or U18359 (N_18359,N_14261,N_13980);
or U18360 (N_18360,N_14609,N_13321);
or U18361 (N_18361,N_12848,N_12835);
and U18362 (N_18362,N_15641,N_12297);
and U18363 (N_18363,N_15083,N_14112);
and U18364 (N_18364,N_15508,N_13730);
xor U18365 (N_18365,N_14404,N_14553);
and U18366 (N_18366,N_15445,N_13897);
or U18367 (N_18367,N_14722,N_13032);
nand U18368 (N_18368,N_15492,N_12873);
nand U18369 (N_18369,N_14907,N_14098);
or U18370 (N_18370,N_13551,N_12833);
and U18371 (N_18371,N_15115,N_12495);
nand U18372 (N_18372,N_14440,N_14796);
and U18373 (N_18373,N_14883,N_12710);
nand U18374 (N_18374,N_13717,N_12943);
or U18375 (N_18375,N_14348,N_15331);
or U18376 (N_18376,N_14251,N_15715);
or U18377 (N_18377,N_14860,N_13958);
and U18378 (N_18378,N_13066,N_12810);
or U18379 (N_18379,N_13217,N_15574);
or U18380 (N_18380,N_13065,N_13294);
and U18381 (N_18381,N_12584,N_13810);
nor U18382 (N_18382,N_12648,N_15396);
nand U18383 (N_18383,N_12921,N_15305);
nor U18384 (N_18384,N_12369,N_12230);
or U18385 (N_18385,N_12425,N_15722);
and U18386 (N_18386,N_13123,N_14409);
nor U18387 (N_18387,N_14754,N_15212);
and U18388 (N_18388,N_12371,N_15962);
or U18389 (N_18389,N_14431,N_15323);
nand U18390 (N_18390,N_13968,N_15548);
and U18391 (N_18391,N_12775,N_14217);
and U18392 (N_18392,N_13427,N_15350);
and U18393 (N_18393,N_12552,N_12240);
nor U18394 (N_18394,N_14417,N_14494);
or U18395 (N_18395,N_15588,N_12192);
nand U18396 (N_18396,N_13567,N_14207);
and U18397 (N_18397,N_15926,N_12657);
xor U18398 (N_18398,N_14217,N_15214);
xor U18399 (N_18399,N_12971,N_13383);
nor U18400 (N_18400,N_15385,N_13002);
xor U18401 (N_18401,N_12596,N_12343);
or U18402 (N_18402,N_12323,N_13888);
or U18403 (N_18403,N_12860,N_14635);
and U18404 (N_18404,N_14229,N_12052);
and U18405 (N_18405,N_12293,N_15671);
nand U18406 (N_18406,N_13143,N_13041);
and U18407 (N_18407,N_13338,N_12958);
and U18408 (N_18408,N_12774,N_14750);
nand U18409 (N_18409,N_14985,N_13609);
or U18410 (N_18410,N_14430,N_13241);
or U18411 (N_18411,N_15343,N_13991);
nor U18412 (N_18412,N_14422,N_14832);
nor U18413 (N_18413,N_15404,N_14526);
nand U18414 (N_18414,N_13609,N_15930);
nor U18415 (N_18415,N_12156,N_13180);
and U18416 (N_18416,N_12251,N_14282);
nor U18417 (N_18417,N_15216,N_14492);
nor U18418 (N_18418,N_14611,N_12030);
nand U18419 (N_18419,N_15810,N_13376);
nor U18420 (N_18420,N_15665,N_14654);
nor U18421 (N_18421,N_13265,N_15729);
and U18422 (N_18422,N_13129,N_14101);
nor U18423 (N_18423,N_15840,N_15663);
or U18424 (N_18424,N_13137,N_14226);
and U18425 (N_18425,N_14291,N_12601);
nor U18426 (N_18426,N_13527,N_13638);
nand U18427 (N_18427,N_12773,N_12636);
and U18428 (N_18428,N_14112,N_14512);
nand U18429 (N_18429,N_15729,N_15508);
xnor U18430 (N_18430,N_14443,N_13671);
nor U18431 (N_18431,N_15379,N_12802);
nor U18432 (N_18432,N_13219,N_12095);
and U18433 (N_18433,N_15578,N_13608);
and U18434 (N_18434,N_14417,N_14265);
nor U18435 (N_18435,N_15189,N_15319);
or U18436 (N_18436,N_13131,N_14471);
or U18437 (N_18437,N_14950,N_13821);
nor U18438 (N_18438,N_12456,N_14065);
nand U18439 (N_18439,N_12835,N_14637);
xor U18440 (N_18440,N_12085,N_15982);
nor U18441 (N_18441,N_12873,N_15516);
nor U18442 (N_18442,N_12333,N_14954);
and U18443 (N_18443,N_13730,N_14588);
and U18444 (N_18444,N_12052,N_13011);
or U18445 (N_18445,N_13784,N_15446);
nand U18446 (N_18446,N_14879,N_13667);
nor U18447 (N_18447,N_15134,N_15132);
or U18448 (N_18448,N_14038,N_14699);
nor U18449 (N_18449,N_15427,N_12294);
nor U18450 (N_18450,N_13669,N_15446);
or U18451 (N_18451,N_15611,N_13033);
nand U18452 (N_18452,N_15103,N_12288);
nor U18453 (N_18453,N_15003,N_14211);
nor U18454 (N_18454,N_15650,N_14533);
or U18455 (N_18455,N_13463,N_12452);
and U18456 (N_18456,N_15313,N_13814);
xnor U18457 (N_18457,N_14419,N_12461);
and U18458 (N_18458,N_15863,N_12774);
and U18459 (N_18459,N_15723,N_12156);
or U18460 (N_18460,N_13667,N_13544);
and U18461 (N_18461,N_14596,N_12735);
or U18462 (N_18462,N_14604,N_14612);
or U18463 (N_18463,N_13299,N_14938);
nor U18464 (N_18464,N_13824,N_12756);
xor U18465 (N_18465,N_12676,N_13770);
nor U18466 (N_18466,N_12474,N_15373);
xnor U18467 (N_18467,N_14338,N_14064);
or U18468 (N_18468,N_14093,N_14957);
or U18469 (N_18469,N_13609,N_12219);
and U18470 (N_18470,N_13795,N_12748);
and U18471 (N_18471,N_12013,N_15146);
and U18472 (N_18472,N_14527,N_13554);
or U18473 (N_18473,N_14365,N_12506);
xor U18474 (N_18474,N_13136,N_13223);
and U18475 (N_18475,N_14131,N_12385);
or U18476 (N_18476,N_14736,N_13504);
and U18477 (N_18477,N_13518,N_14783);
nand U18478 (N_18478,N_13735,N_13658);
nand U18479 (N_18479,N_12820,N_15059);
nand U18480 (N_18480,N_15803,N_15335);
nor U18481 (N_18481,N_12877,N_14416);
nor U18482 (N_18482,N_13496,N_12267);
nand U18483 (N_18483,N_12289,N_12699);
or U18484 (N_18484,N_13449,N_15107);
and U18485 (N_18485,N_13754,N_13813);
nand U18486 (N_18486,N_13712,N_14254);
nand U18487 (N_18487,N_12166,N_13498);
nand U18488 (N_18488,N_15597,N_14033);
or U18489 (N_18489,N_12933,N_14119);
nand U18490 (N_18490,N_15000,N_15922);
and U18491 (N_18491,N_15701,N_15488);
nand U18492 (N_18492,N_15013,N_12275);
nor U18493 (N_18493,N_15541,N_12473);
or U18494 (N_18494,N_12579,N_13338);
and U18495 (N_18495,N_12749,N_12055);
nand U18496 (N_18496,N_15682,N_12771);
or U18497 (N_18497,N_15362,N_14547);
and U18498 (N_18498,N_13622,N_14475);
or U18499 (N_18499,N_14235,N_13784);
and U18500 (N_18500,N_12953,N_14305);
and U18501 (N_18501,N_13413,N_14465);
xnor U18502 (N_18502,N_14108,N_12826);
or U18503 (N_18503,N_12659,N_13560);
or U18504 (N_18504,N_14287,N_15251);
and U18505 (N_18505,N_14581,N_12569);
nor U18506 (N_18506,N_15176,N_12972);
nand U18507 (N_18507,N_14550,N_12630);
nand U18508 (N_18508,N_13194,N_14734);
or U18509 (N_18509,N_13458,N_14861);
and U18510 (N_18510,N_12734,N_13103);
nand U18511 (N_18511,N_14716,N_15990);
or U18512 (N_18512,N_12858,N_14899);
and U18513 (N_18513,N_12312,N_15258);
nand U18514 (N_18514,N_13318,N_12710);
nor U18515 (N_18515,N_14878,N_14950);
nor U18516 (N_18516,N_14118,N_15694);
or U18517 (N_18517,N_15417,N_13396);
or U18518 (N_18518,N_15910,N_15432);
nand U18519 (N_18519,N_15824,N_15206);
and U18520 (N_18520,N_14596,N_14591);
and U18521 (N_18521,N_14836,N_13495);
nand U18522 (N_18522,N_14000,N_12186);
nor U18523 (N_18523,N_15448,N_12093);
and U18524 (N_18524,N_15305,N_14960);
or U18525 (N_18525,N_14752,N_14244);
nor U18526 (N_18526,N_15324,N_13665);
nor U18527 (N_18527,N_13408,N_12692);
nand U18528 (N_18528,N_15806,N_14624);
nand U18529 (N_18529,N_14351,N_12554);
and U18530 (N_18530,N_12261,N_12930);
and U18531 (N_18531,N_13879,N_15580);
nand U18532 (N_18532,N_14302,N_14310);
nand U18533 (N_18533,N_15997,N_12235);
nor U18534 (N_18534,N_13696,N_14382);
or U18535 (N_18535,N_13372,N_15008);
nand U18536 (N_18536,N_15941,N_13890);
nand U18537 (N_18537,N_13908,N_14780);
or U18538 (N_18538,N_12371,N_15687);
and U18539 (N_18539,N_13504,N_14389);
and U18540 (N_18540,N_14428,N_15374);
nand U18541 (N_18541,N_13857,N_12324);
nor U18542 (N_18542,N_12765,N_13437);
nand U18543 (N_18543,N_14969,N_14771);
and U18544 (N_18544,N_13898,N_13126);
or U18545 (N_18545,N_15891,N_15890);
nand U18546 (N_18546,N_15206,N_13768);
or U18547 (N_18547,N_13580,N_13543);
or U18548 (N_18548,N_12417,N_13829);
nor U18549 (N_18549,N_15019,N_12046);
nand U18550 (N_18550,N_13615,N_13128);
and U18551 (N_18551,N_12078,N_12961);
and U18552 (N_18552,N_14344,N_14925);
and U18553 (N_18553,N_12572,N_12472);
nand U18554 (N_18554,N_15061,N_12120);
or U18555 (N_18555,N_12784,N_15135);
nor U18556 (N_18556,N_12041,N_15193);
xnor U18557 (N_18557,N_12755,N_14056);
nand U18558 (N_18558,N_14902,N_15853);
or U18559 (N_18559,N_14492,N_14512);
xnor U18560 (N_18560,N_13836,N_13596);
and U18561 (N_18561,N_13643,N_12524);
or U18562 (N_18562,N_13047,N_14672);
and U18563 (N_18563,N_14959,N_15720);
nand U18564 (N_18564,N_13648,N_13263);
xor U18565 (N_18565,N_13566,N_15684);
or U18566 (N_18566,N_12702,N_12765);
nor U18567 (N_18567,N_13439,N_12581);
or U18568 (N_18568,N_12493,N_15027);
and U18569 (N_18569,N_14818,N_13044);
or U18570 (N_18570,N_12444,N_15640);
or U18571 (N_18571,N_12197,N_15578);
nor U18572 (N_18572,N_15247,N_15294);
and U18573 (N_18573,N_15321,N_12695);
xnor U18574 (N_18574,N_12133,N_14065);
and U18575 (N_18575,N_12337,N_14607);
and U18576 (N_18576,N_12289,N_12065);
xor U18577 (N_18577,N_13274,N_14071);
nand U18578 (N_18578,N_15690,N_12348);
nand U18579 (N_18579,N_12216,N_14057);
nor U18580 (N_18580,N_13932,N_14462);
and U18581 (N_18581,N_14335,N_14647);
or U18582 (N_18582,N_13745,N_14844);
xor U18583 (N_18583,N_12055,N_15434);
or U18584 (N_18584,N_15995,N_15158);
and U18585 (N_18585,N_14375,N_13131);
and U18586 (N_18586,N_13466,N_13328);
nor U18587 (N_18587,N_13822,N_12648);
or U18588 (N_18588,N_13371,N_12233);
or U18589 (N_18589,N_13819,N_12128);
or U18590 (N_18590,N_13121,N_15094);
xnor U18591 (N_18591,N_14358,N_14782);
nand U18592 (N_18592,N_14240,N_15782);
and U18593 (N_18593,N_13808,N_14393);
and U18594 (N_18594,N_15548,N_14354);
xnor U18595 (N_18595,N_15725,N_12700);
or U18596 (N_18596,N_14844,N_15473);
or U18597 (N_18597,N_15393,N_15686);
and U18598 (N_18598,N_15381,N_13506);
nor U18599 (N_18599,N_14694,N_13372);
or U18600 (N_18600,N_12412,N_15975);
or U18601 (N_18601,N_15821,N_14051);
and U18602 (N_18602,N_14613,N_13460);
and U18603 (N_18603,N_13486,N_14686);
and U18604 (N_18604,N_13475,N_15701);
nor U18605 (N_18605,N_14313,N_12453);
and U18606 (N_18606,N_13078,N_13003);
nand U18607 (N_18607,N_13926,N_12170);
nor U18608 (N_18608,N_12124,N_12238);
and U18609 (N_18609,N_15671,N_13433);
and U18610 (N_18610,N_14400,N_14512);
and U18611 (N_18611,N_15292,N_13877);
nand U18612 (N_18612,N_12771,N_14344);
nand U18613 (N_18613,N_12188,N_15355);
nand U18614 (N_18614,N_14659,N_12956);
or U18615 (N_18615,N_15863,N_13540);
or U18616 (N_18616,N_15032,N_13983);
nand U18617 (N_18617,N_12201,N_15113);
or U18618 (N_18618,N_14310,N_13658);
nand U18619 (N_18619,N_12392,N_14841);
or U18620 (N_18620,N_12077,N_12494);
nand U18621 (N_18621,N_15922,N_13134);
nor U18622 (N_18622,N_14274,N_13444);
nand U18623 (N_18623,N_12601,N_15132);
xor U18624 (N_18624,N_14394,N_14189);
nor U18625 (N_18625,N_13458,N_13473);
nor U18626 (N_18626,N_12339,N_14160);
and U18627 (N_18627,N_13962,N_15959);
nand U18628 (N_18628,N_15862,N_13015);
nor U18629 (N_18629,N_13798,N_13121);
or U18630 (N_18630,N_14204,N_15047);
or U18631 (N_18631,N_13172,N_14204);
or U18632 (N_18632,N_15499,N_12038);
or U18633 (N_18633,N_15163,N_15676);
and U18634 (N_18634,N_13372,N_15979);
nor U18635 (N_18635,N_14026,N_12398);
and U18636 (N_18636,N_15536,N_15016);
or U18637 (N_18637,N_15387,N_15886);
nor U18638 (N_18638,N_15186,N_13329);
or U18639 (N_18639,N_14019,N_13249);
nor U18640 (N_18640,N_12877,N_13737);
xor U18641 (N_18641,N_14640,N_12330);
nand U18642 (N_18642,N_14756,N_15344);
and U18643 (N_18643,N_13004,N_14627);
and U18644 (N_18644,N_13250,N_12320);
or U18645 (N_18645,N_15374,N_14407);
nor U18646 (N_18646,N_13451,N_13032);
nand U18647 (N_18647,N_12716,N_15880);
nor U18648 (N_18648,N_14403,N_13176);
or U18649 (N_18649,N_13162,N_12222);
nand U18650 (N_18650,N_15243,N_12217);
nand U18651 (N_18651,N_14336,N_12515);
xnor U18652 (N_18652,N_15288,N_12386);
nand U18653 (N_18653,N_14681,N_13934);
xnor U18654 (N_18654,N_13695,N_14353);
nand U18655 (N_18655,N_13897,N_15043);
nor U18656 (N_18656,N_14727,N_13493);
or U18657 (N_18657,N_14829,N_15407);
nor U18658 (N_18658,N_14622,N_12725);
xnor U18659 (N_18659,N_14441,N_15970);
or U18660 (N_18660,N_15675,N_14860);
or U18661 (N_18661,N_14818,N_13091);
nor U18662 (N_18662,N_14001,N_15084);
nand U18663 (N_18663,N_13995,N_14484);
nand U18664 (N_18664,N_15927,N_14083);
and U18665 (N_18665,N_14852,N_15995);
or U18666 (N_18666,N_12384,N_15583);
and U18667 (N_18667,N_12401,N_12448);
nand U18668 (N_18668,N_13738,N_13783);
or U18669 (N_18669,N_14203,N_12272);
or U18670 (N_18670,N_13181,N_13532);
nor U18671 (N_18671,N_15357,N_13360);
and U18672 (N_18672,N_12811,N_13716);
xnor U18673 (N_18673,N_12648,N_14210);
xor U18674 (N_18674,N_15679,N_12280);
or U18675 (N_18675,N_14162,N_13304);
and U18676 (N_18676,N_12421,N_14185);
and U18677 (N_18677,N_12727,N_12774);
or U18678 (N_18678,N_15651,N_13065);
and U18679 (N_18679,N_14467,N_15286);
nor U18680 (N_18680,N_15006,N_15012);
and U18681 (N_18681,N_14780,N_14644);
or U18682 (N_18682,N_13061,N_14735);
nor U18683 (N_18683,N_15585,N_14521);
nor U18684 (N_18684,N_14296,N_12828);
or U18685 (N_18685,N_15081,N_14647);
nand U18686 (N_18686,N_15108,N_14141);
and U18687 (N_18687,N_15090,N_15354);
or U18688 (N_18688,N_13014,N_12719);
nor U18689 (N_18689,N_15927,N_12265);
nor U18690 (N_18690,N_12641,N_15753);
xnor U18691 (N_18691,N_13014,N_13296);
and U18692 (N_18692,N_15359,N_13067);
or U18693 (N_18693,N_14311,N_13388);
and U18694 (N_18694,N_13056,N_13722);
or U18695 (N_18695,N_14619,N_13897);
and U18696 (N_18696,N_13287,N_13339);
xnor U18697 (N_18697,N_14917,N_14310);
and U18698 (N_18698,N_15096,N_14145);
nor U18699 (N_18699,N_14571,N_14206);
nand U18700 (N_18700,N_12442,N_15267);
nor U18701 (N_18701,N_13276,N_12270);
and U18702 (N_18702,N_13837,N_13029);
nor U18703 (N_18703,N_13268,N_15740);
nor U18704 (N_18704,N_14009,N_12750);
and U18705 (N_18705,N_14998,N_15601);
and U18706 (N_18706,N_14542,N_15737);
nor U18707 (N_18707,N_12566,N_13181);
and U18708 (N_18708,N_14708,N_13745);
and U18709 (N_18709,N_13313,N_15549);
nor U18710 (N_18710,N_12305,N_15363);
or U18711 (N_18711,N_13423,N_15878);
nand U18712 (N_18712,N_14454,N_13489);
or U18713 (N_18713,N_13218,N_13550);
and U18714 (N_18714,N_15933,N_15713);
nand U18715 (N_18715,N_15434,N_12111);
nand U18716 (N_18716,N_13208,N_14163);
nor U18717 (N_18717,N_12201,N_15845);
nand U18718 (N_18718,N_15806,N_13298);
and U18719 (N_18719,N_13441,N_15211);
and U18720 (N_18720,N_12764,N_12412);
or U18721 (N_18721,N_15895,N_15465);
nor U18722 (N_18722,N_12527,N_14021);
nor U18723 (N_18723,N_15932,N_12726);
and U18724 (N_18724,N_14228,N_13267);
or U18725 (N_18725,N_14358,N_14606);
xnor U18726 (N_18726,N_15660,N_12713);
or U18727 (N_18727,N_14260,N_14128);
or U18728 (N_18728,N_13262,N_14007);
and U18729 (N_18729,N_14403,N_14974);
and U18730 (N_18730,N_14456,N_13049);
xnor U18731 (N_18731,N_12574,N_14535);
nand U18732 (N_18732,N_15820,N_13341);
and U18733 (N_18733,N_13981,N_14107);
nor U18734 (N_18734,N_15010,N_14267);
and U18735 (N_18735,N_15796,N_15299);
xnor U18736 (N_18736,N_14468,N_12995);
nand U18737 (N_18737,N_12076,N_12908);
or U18738 (N_18738,N_13286,N_15622);
nand U18739 (N_18739,N_15844,N_14234);
nand U18740 (N_18740,N_15714,N_13566);
nand U18741 (N_18741,N_14968,N_15817);
or U18742 (N_18742,N_14829,N_13507);
nor U18743 (N_18743,N_15692,N_15793);
and U18744 (N_18744,N_14623,N_13956);
and U18745 (N_18745,N_13402,N_13109);
xnor U18746 (N_18746,N_12035,N_14465);
nand U18747 (N_18747,N_14709,N_13480);
or U18748 (N_18748,N_13988,N_15269);
or U18749 (N_18749,N_15956,N_13400);
nor U18750 (N_18750,N_12527,N_13770);
nor U18751 (N_18751,N_15404,N_14112);
or U18752 (N_18752,N_15202,N_14395);
nor U18753 (N_18753,N_12345,N_13936);
or U18754 (N_18754,N_15141,N_12211);
and U18755 (N_18755,N_14254,N_15534);
and U18756 (N_18756,N_13984,N_14918);
or U18757 (N_18757,N_12656,N_14343);
xor U18758 (N_18758,N_14446,N_15813);
and U18759 (N_18759,N_12510,N_12210);
nand U18760 (N_18760,N_14048,N_13364);
nand U18761 (N_18761,N_13308,N_12793);
nor U18762 (N_18762,N_12356,N_15256);
or U18763 (N_18763,N_13084,N_15175);
and U18764 (N_18764,N_14626,N_15512);
or U18765 (N_18765,N_15916,N_15808);
and U18766 (N_18766,N_15060,N_15155);
nand U18767 (N_18767,N_15634,N_12515);
xor U18768 (N_18768,N_14096,N_12929);
nor U18769 (N_18769,N_14962,N_13183);
or U18770 (N_18770,N_14568,N_12399);
nand U18771 (N_18771,N_14923,N_12057);
or U18772 (N_18772,N_14642,N_15362);
nor U18773 (N_18773,N_14223,N_12422);
nor U18774 (N_18774,N_14123,N_15466);
and U18775 (N_18775,N_12422,N_13065);
nand U18776 (N_18776,N_12726,N_13955);
and U18777 (N_18777,N_14855,N_15080);
and U18778 (N_18778,N_12042,N_12704);
nand U18779 (N_18779,N_13930,N_14085);
nand U18780 (N_18780,N_14247,N_13648);
or U18781 (N_18781,N_12606,N_15647);
xor U18782 (N_18782,N_12982,N_13710);
and U18783 (N_18783,N_14952,N_12637);
xnor U18784 (N_18784,N_12546,N_14713);
nor U18785 (N_18785,N_12039,N_14102);
nand U18786 (N_18786,N_12314,N_14881);
nand U18787 (N_18787,N_12409,N_15208);
xnor U18788 (N_18788,N_15770,N_14251);
nor U18789 (N_18789,N_13026,N_13318);
nand U18790 (N_18790,N_14971,N_13519);
or U18791 (N_18791,N_13124,N_12818);
nand U18792 (N_18792,N_13289,N_13130);
xnor U18793 (N_18793,N_15394,N_15374);
nor U18794 (N_18794,N_15557,N_14265);
nand U18795 (N_18795,N_15166,N_12288);
or U18796 (N_18796,N_15343,N_12945);
nor U18797 (N_18797,N_13365,N_15120);
and U18798 (N_18798,N_15219,N_14591);
nand U18799 (N_18799,N_14613,N_14341);
xnor U18800 (N_18800,N_12556,N_13290);
and U18801 (N_18801,N_15370,N_12545);
or U18802 (N_18802,N_14468,N_12021);
nand U18803 (N_18803,N_12360,N_12823);
nand U18804 (N_18804,N_15578,N_15990);
nand U18805 (N_18805,N_12744,N_12380);
or U18806 (N_18806,N_12245,N_13951);
nor U18807 (N_18807,N_14152,N_15637);
and U18808 (N_18808,N_12928,N_15433);
xor U18809 (N_18809,N_12700,N_14322);
nor U18810 (N_18810,N_15521,N_12686);
and U18811 (N_18811,N_13037,N_12017);
and U18812 (N_18812,N_14357,N_15843);
xor U18813 (N_18813,N_15810,N_15075);
nand U18814 (N_18814,N_12303,N_13805);
nor U18815 (N_18815,N_15814,N_14474);
nand U18816 (N_18816,N_15136,N_13418);
and U18817 (N_18817,N_13227,N_13665);
nor U18818 (N_18818,N_12642,N_13066);
nor U18819 (N_18819,N_13213,N_13670);
or U18820 (N_18820,N_15041,N_12388);
and U18821 (N_18821,N_14210,N_12769);
nand U18822 (N_18822,N_12697,N_14512);
or U18823 (N_18823,N_14449,N_13656);
or U18824 (N_18824,N_14479,N_15054);
xnor U18825 (N_18825,N_12364,N_12774);
nand U18826 (N_18826,N_15529,N_13022);
or U18827 (N_18827,N_13264,N_13374);
nand U18828 (N_18828,N_14121,N_14368);
nor U18829 (N_18829,N_15206,N_13476);
nor U18830 (N_18830,N_12416,N_12957);
and U18831 (N_18831,N_13914,N_15925);
or U18832 (N_18832,N_15695,N_12850);
nand U18833 (N_18833,N_15273,N_12729);
and U18834 (N_18834,N_15612,N_15864);
nand U18835 (N_18835,N_14128,N_15675);
xnor U18836 (N_18836,N_15640,N_14544);
or U18837 (N_18837,N_13948,N_13453);
nor U18838 (N_18838,N_14906,N_14303);
or U18839 (N_18839,N_15787,N_12634);
nand U18840 (N_18840,N_12622,N_13356);
and U18841 (N_18841,N_15097,N_12929);
or U18842 (N_18842,N_12095,N_15507);
xnor U18843 (N_18843,N_12161,N_14813);
xor U18844 (N_18844,N_12028,N_15536);
nor U18845 (N_18845,N_14111,N_15706);
nor U18846 (N_18846,N_14300,N_13124);
nor U18847 (N_18847,N_12292,N_15404);
or U18848 (N_18848,N_15806,N_14299);
and U18849 (N_18849,N_13099,N_13647);
or U18850 (N_18850,N_14846,N_12153);
or U18851 (N_18851,N_14690,N_14086);
or U18852 (N_18852,N_12859,N_15292);
nand U18853 (N_18853,N_12131,N_14076);
or U18854 (N_18854,N_13907,N_15979);
and U18855 (N_18855,N_12837,N_13434);
and U18856 (N_18856,N_15790,N_15839);
nor U18857 (N_18857,N_14372,N_13373);
and U18858 (N_18858,N_12509,N_13207);
xnor U18859 (N_18859,N_14258,N_15681);
and U18860 (N_18860,N_12679,N_12593);
xnor U18861 (N_18861,N_13303,N_13210);
nand U18862 (N_18862,N_14889,N_14456);
and U18863 (N_18863,N_15192,N_15556);
and U18864 (N_18864,N_12336,N_13807);
nand U18865 (N_18865,N_15840,N_14674);
nor U18866 (N_18866,N_13693,N_15834);
or U18867 (N_18867,N_15648,N_15508);
nand U18868 (N_18868,N_15811,N_13945);
nor U18869 (N_18869,N_15774,N_12081);
and U18870 (N_18870,N_14913,N_14801);
nand U18871 (N_18871,N_12361,N_15692);
nand U18872 (N_18872,N_12002,N_12615);
and U18873 (N_18873,N_13589,N_15915);
or U18874 (N_18874,N_14724,N_15613);
nand U18875 (N_18875,N_13500,N_14748);
nand U18876 (N_18876,N_12333,N_12257);
nand U18877 (N_18877,N_14008,N_14742);
nand U18878 (N_18878,N_15259,N_14673);
nor U18879 (N_18879,N_13673,N_12214);
nand U18880 (N_18880,N_15168,N_14289);
or U18881 (N_18881,N_13932,N_12706);
or U18882 (N_18882,N_12765,N_13219);
or U18883 (N_18883,N_12273,N_15753);
or U18884 (N_18884,N_12401,N_14254);
nand U18885 (N_18885,N_15382,N_15940);
nor U18886 (N_18886,N_13705,N_12196);
nand U18887 (N_18887,N_14377,N_12545);
nand U18888 (N_18888,N_13386,N_13402);
nor U18889 (N_18889,N_12602,N_15136);
or U18890 (N_18890,N_14959,N_13404);
xor U18891 (N_18891,N_12482,N_13836);
nor U18892 (N_18892,N_14455,N_13388);
and U18893 (N_18893,N_13072,N_13192);
nand U18894 (N_18894,N_14266,N_15123);
and U18895 (N_18895,N_12408,N_14025);
or U18896 (N_18896,N_14694,N_14140);
and U18897 (N_18897,N_12219,N_14836);
and U18898 (N_18898,N_14623,N_15365);
xor U18899 (N_18899,N_15343,N_15154);
nand U18900 (N_18900,N_13520,N_14173);
nand U18901 (N_18901,N_13758,N_12425);
nor U18902 (N_18902,N_14386,N_12002);
or U18903 (N_18903,N_12540,N_13177);
and U18904 (N_18904,N_15491,N_15714);
nor U18905 (N_18905,N_15422,N_14397);
nand U18906 (N_18906,N_12170,N_12977);
nand U18907 (N_18907,N_12885,N_13411);
nor U18908 (N_18908,N_13783,N_14062);
and U18909 (N_18909,N_15940,N_15082);
and U18910 (N_18910,N_15626,N_14053);
or U18911 (N_18911,N_13743,N_15489);
and U18912 (N_18912,N_12614,N_14217);
nand U18913 (N_18913,N_14664,N_14168);
and U18914 (N_18914,N_12323,N_13725);
xnor U18915 (N_18915,N_12233,N_14194);
nand U18916 (N_18916,N_13214,N_13393);
and U18917 (N_18917,N_15764,N_13750);
and U18918 (N_18918,N_14874,N_13973);
nand U18919 (N_18919,N_14926,N_14690);
nand U18920 (N_18920,N_12705,N_12507);
or U18921 (N_18921,N_15984,N_15802);
or U18922 (N_18922,N_12415,N_13655);
xor U18923 (N_18923,N_12785,N_15776);
or U18924 (N_18924,N_12802,N_15538);
nand U18925 (N_18925,N_15346,N_13796);
or U18926 (N_18926,N_12000,N_13403);
and U18927 (N_18927,N_15027,N_15625);
or U18928 (N_18928,N_12741,N_12580);
nand U18929 (N_18929,N_15557,N_15751);
and U18930 (N_18930,N_14266,N_12312);
nand U18931 (N_18931,N_12667,N_14273);
nor U18932 (N_18932,N_12829,N_12901);
and U18933 (N_18933,N_15889,N_13412);
nor U18934 (N_18934,N_13757,N_12376);
or U18935 (N_18935,N_15639,N_15505);
or U18936 (N_18936,N_13363,N_12075);
xor U18937 (N_18937,N_15997,N_14303);
nand U18938 (N_18938,N_15932,N_12975);
nor U18939 (N_18939,N_14349,N_13457);
nor U18940 (N_18940,N_15415,N_12590);
nor U18941 (N_18941,N_13391,N_14503);
xor U18942 (N_18942,N_12784,N_13144);
nand U18943 (N_18943,N_15505,N_13562);
nand U18944 (N_18944,N_14941,N_12896);
or U18945 (N_18945,N_13528,N_12524);
nand U18946 (N_18946,N_13729,N_13510);
nor U18947 (N_18947,N_15213,N_15763);
and U18948 (N_18948,N_13900,N_15203);
and U18949 (N_18949,N_13956,N_13500);
nor U18950 (N_18950,N_15461,N_15670);
nand U18951 (N_18951,N_15362,N_15330);
nor U18952 (N_18952,N_13806,N_13474);
and U18953 (N_18953,N_14139,N_12345);
nand U18954 (N_18954,N_12042,N_12481);
nor U18955 (N_18955,N_12871,N_12927);
or U18956 (N_18956,N_12454,N_12978);
nand U18957 (N_18957,N_12604,N_12508);
nand U18958 (N_18958,N_12752,N_15425);
nand U18959 (N_18959,N_12898,N_14753);
and U18960 (N_18960,N_13209,N_12625);
or U18961 (N_18961,N_14766,N_13769);
or U18962 (N_18962,N_14056,N_14360);
nand U18963 (N_18963,N_14930,N_15007);
nand U18964 (N_18964,N_14368,N_12547);
or U18965 (N_18965,N_14931,N_15807);
nand U18966 (N_18966,N_15168,N_12094);
nor U18967 (N_18967,N_14347,N_12309);
or U18968 (N_18968,N_12466,N_14440);
nor U18969 (N_18969,N_12193,N_13001);
and U18970 (N_18970,N_12283,N_14974);
or U18971 (N_18971,N_13496,N_14453);
xor U18972 (N_18972,N_13480,N_15125);
or U18973 (N_18973,N_13981,N_15827);
xnor U18974 (N_18974,N_12859,N_15772);
nand U18975 (N_18975,N_15223,N_14857);
xor U18976 (N_18976,N_14728,N_14092);
and U18977 (N_18977,N_13705,N_12962);
nor U18978 (N_18978,N_14785,N_13125);
nand U18979 (N_18979,N_14290,N_14774);
nor U18980 (N_18980,N_13475,N_15844);
or U18981 (N_18981,N_14519,N_12324);
or U18982 (N_18982,N_12800,N_14762);
or U18983 (N_18983,N_12510,N_12981);
or U18984 (N_18984,N_15320,N_13170);
nor U18985 (N_18985,N_13796,N_13119);
or U18986 (N_18986,N_14510,N_15267);
nand U18987 (N_18987,N_12421,N_14746);
and U18988 (N_18988,N_12565,N_15639);
nand U18989 (N_18989,N_12959,N_15948);
and U18990 (N_18990,N_13572,N_12976);
nor U18991 (N_18991,N_12693,N_13478);
and U18992 (N_18992,N_15489,N_15020);
or U18993 (N_18993,N_12767,N_12174);
nor U18994 (N_18994,N_14290,N_13591);
nand U18995 (N_18995,N_12201,N_12649);
nand U18996 (N_18996,N_12086,N_12371);
and U18997 (N_18997,N_15204,N_12829);
nor U18998 (N_18998,N_12956,N_12630);
or U18999 (N_18999,N_14698,N_13346);
nor U19000 (N_19000,N_12601,N_14080);
nand U19001 (N_19001,N_14599,N_14832);
xor U19002 (N_19002,N_12512,N_14288);
nand U19003 (N_19003,N_14435,N_12722);
and U19004 (N_19004,N_12100,N_15458);
nand U19005 (N_19005,N_14132,N_12849);
and U19006 (N_19006,N_15846,N_13787);
or U19007 (N_19007,N_12268,N_14763);
and U19008 (N_19008,N_13152,N_12402);
or U19009 (N_19009,N_15310,N_15378);
nand U19010 (N_19010,N_12291,N_15806);
nand U19011 (N_19011,N_14799,N_15830);
or U19012 (N_19012,N_14727,N_12335);
nand U19013 (N_19013,N_14480,N_15906);
and U19014 (N_19014,N_14721,N_13841);
nor U19015 (N_19015,N_12352,N_15232);
and U19016 (N_19016,N_13611,N_15928);
and U19017 (N_19017,N_12811,N_15723);
and U19018 (N_19018,N_15750,N_15276);
nand U19019 (N_19019,N_15783,N_15071);
or U19020 (N_19020,N_13246,N_13723);
and U19021 (N_19021,N_14648,N_15557);
nor U19022 (N_19022,N_14154,N_12906);
or U19023 (N_19023,N_12254,N_14791);
or U19024 (N_19024,N_14859,N_15430);
xnor U19025 (N_19025,N_14524,N_15660);
or U19026 (N_19026,N_14518,N_15505);
nor U19027 (N_19027,N_14548,N_12875);
and U19028 (N_19028,N_12249,N_15640);
and U19029 (N_19029,N_14689,N_15464);
nor U19030 (N_19030,N_15684,N_15762);
or U19031 (N_19031,N_12399,N_12667);
or U19032 (N_19032,N_14091,N_14742);
nor U19033 (N_19033,N_13536,N_12470);
xnor U19034 (N_19034,N_12252,N_14116);
xnor U19035 (N_19035,N_13028,N_12781);
or U19036 (N_19036,N_15730,N_14075);
and U19037 (N_19037,N_12340,N_13487);
and U19038 (N_19038,N_12880,N_14429);
nand U19039 (N_19039,N_12547,N_12109);
or U19040 (N_19040,N_14082,N_15944);
nor U19041 (N_19041,N_13700,N_14269);
and U19042 (N_19042,N_12359,N_14938);
nor U19043 (N_19043,N_15554,N_14970);
and U19044 (N_19044,N_15488,N_13737);
nor U19045 (N_19045,N_13939,N_12855);
nand U19046 (N_19046,N_15603,N_15437);
xor U19047 (N_19047,N_14188,N_13722);
nand U19048 (N_19048,N_13125,N_15446);
nand U19049 (N_19049,N_12424,N_15943);
nor U19050 (N_19050,N_15782,N_15742);
or U19051 (N_19051,N_14926,N_13534);
nand U19052 (N_19052,N_13922,N_14971);
or U19053 (N_19053,N_12105,N_12453);
and U19054 (N_19054,N_14736,N_15018);
xor U19055 (N_19055,N_13327,N_13611);
or U19056 (N_19056,N_14243,N_15475);
nor U19057 (N_19057,N_13809,N_13778);
or U19058 (N_19058,N_14596,N_14351);
nor U19059 (N_19059,N_12973,N_12801);
or U19060 (N_19060,N_12895,N_15097);
or U19061 (N_19061,N_13559,N_15123);
nand U19062 (N_19062,N_13424,N_12945);
xor U19063 (N_19063,N_15033,N_12215);
nor U19064 (N_19064,N_13332,N_13222);
nand U19065 (N_19065,N_12580,N_13546);
nand U19066 (N_19066,N_13436,N_14879);
nand U19067 (N_19067,N_13436,N_13111);
or U19068 (N_19068,N_14535,N_12030);
and U19069 (N_19069,N_15294,N_12976);
nor U19070 (N_19070,N_14512,N_13053);
xnor U19071 (N_19071,N_15432,N_14165);
nor U19072 (N_19072,N_15573,N_12804);
xnor U19073 (N_19073,N_12574,N_13506);
nor U19074 (N_19074,N_14211,N_13846);
or U19075 (N_19075,N_12257,N_12177);
nand U19076 (N_19076,N_15121,N_14319);
nand U19077 (N_19077,N_15493,N_14528);
and U19078 (N_19078,N_15441,N_14892);
nand U19079 (N_19079,N_12445,N_13100);
nor U19080 (N_19080,N_12420,N_14175);
nor U19081 (N_19081,N_12892,N_15482);
nand U19082 (N_19082,N_15188,N_14891);
and U19083 (N_19083,N_15298,N_15772);
nand U19084 (N_19084,N_13836,N_12172);
xor U19085 (N_19085,N_14808,N_13759);
nor U19086 (N_19086,N_14371,N_12823);
and U19087 (N_19087,N_14752,N_12887);
or U19088 (N_19088,N_15550,N_13820);
xnor U19089 (N_19089,N_14083,N_13621);
or U19090 (N_19090,N_14090,N_15665);
or U19091 (N_19091,N_12801,N_12270);
nor U19092 (N_19092,N_14638,N_15084);
nor U19093 (N_19093,N_14080,N_13601);
and U19094 (N_19094,N_15070,N_15382);
and U19095 (N_19095,N_13333,N_14086);
or U19096 (N_19096,N_13533,N_12639);
or U19097 (N_19097,N_15982,N_12386);
nor U19098 (N_19098,N_14930,N_13490);
or U19099 (N_19099,N_14078,N_13174);
or U19100 (N_19100,N_12050,N_15354);
and U19101 (N_19101,N_15134,N_14562);
and U19102 (N_19102,N_15733,N_13664);
or U19103 (N_19103,N_12979,N_12781);
and U19104 (N_19104,N_14908,N_15823);
or U19105 (N_19105,N_13882,N_15565);
and U19106 (N_19106,N_12245,N_12120);
and U19107 (N_19107,N_14971,N_14009);
nor U19108 (N_19108,N_15332,N_15965);
nor U19109 (N_19109,N_14042,N_13814);
and U19110 (N_19110,N_12290,N_13864);
or U19111 (N_19111,N_14015,N_14816);
nand U19112 (N_19112,N_14841,N_14892);
nand U19113 (N_19113,N_14131,N_15135);
nor U19114 (N_19114,N_12066,N_14201);
and U19115 (N_19115,N_12575,N_15857);
and U19116 (N_19116,N_14140,N_13014);
and U19117 (N_19117,N_15602,N_12886);
or U19118 (N_19118,N_13321,N_13859);
or U19119 (N_19119,N_14546,N_13333);
xor U19120 (N_19120,N_13694,N_15856);
or U19121 (N_19121,N_14967,N_14158);
or U19122 (N_19122,N_14442,N_15700);
nand U19123 (N_19123,N_12337,N_14472);
nor U19124 (N_19124,N_12334,N_13581);
or U19125 (N_19125,N_13687,N_15266);
or U19126 (N_19126,N_12789,N_15795);
xor U19127 (N_19127,N_14032,N_15158);
or U19128 (N_19128,N_13716,N_15819);
or U19129 (N_19129,N_14419,N_12239);
or U19130 (N_19130,N_12913,N_15063);
and U19131 (N_19131,N_12954,N_14854);
or U19132 (N_19132,N_12174,N_12944);
and U19133 (N_19133,N_12958,N_13722);
and U19134 (N_19134,N_15600,N_14458);
nor U19135 (N_19135,N_13156,N_14393);
and U19136 (N_19136,N_12471,N_12582);
xor U19137 (N_19137,N_15825,N_12306);
or U19138 (N_19138,N_12435,N_13579);
nor U19139 (N_19139,N_12631,N_12826);
or U19140 (N_19140,N_14192,N_12879);
or U19141 (N_19141,N_14618,N_13963);
or U19142 (N_19142,N_12616,N_15418);
or U19143 (N_19143,N_12021,N_15493);
nor U19144 (N_19144,N_14281,N_13301);
nand U19145 (N_19145,N_14015,N_12692);
nand U19146 (N_19146,N_14465,N_14629);
or U19147 (N_19147,N_14028,N_13983);
and U19148 (N_19148,N_14432,N_15152);
or U19149 (N_19149,N_14371,N_12866);
and U19150 (N_19150,N_13172,N_12589);
and U19151 (N_19151,N_14612,N_15525);
nand U19152 (N_19152,N_13663,N_14792);
nor U19153 (N_19153,N_12141,N_15715);
xor U19154 (N_19154,N_14871,N_14145);
xor U19155 (N_19155,N_12281,N_13221);
and U19156 (N_19156,N_13505,N_14552);
and U19157 (N_19157,N_14241,N_13683);
nor U19158 (N_19158,N_15878,N_14690);
and U19159 (N_19159,N_14447,N_13904);
nor U19160 (N_19160,N_13405,N_15094);
nand U19161 (N_19161,N_13638,N_12535);
or U19162 (N_19162,N_13599,N_13285);
or U19163 (N_19163,N_14352,N_14663);
or U19164 (N_19164,N_12363,N_15347);
nand U19165 (N_19165,N_12621,N_15612);
and U19166 (N_19166,N_14803,N_13166);
or U19167 (N_19167,N_12697,N_14954);
xnor U19168 (N_19168,N_12129,N_13513);
or U19169 (N_19169,N_14906,N_13763);
nor U19170 (N_19170,N_15723,N_14021);
or U19171 (N_19171,N_15423,N_12463);
nand U19172 (N_19172,N_14888,N_13392);
or U19173 (N_19173,N_13664,N_14794);
or U19174 (N_19174,N_15765,N_14092);
nor U19175 (N_19175,N_13276,N_12659);
xor U19176 (N_19176,N_15697,N_14314);
xor U19177 (N_19177,N_14532,N_13383);
and U19178 (N_19178,N_14748,N_14547);
or U19179 (N_19179,N_14038,N_15541);
nand U19180 (N_19180,N_14255,N_13233);
and U19181 (N_19181,N_12332,N_15511);
or U19182 (N_19182,N_15367,N_15565);
xor U19183 (N_19183,N_12070,N_12433);
nand U19184 (N_19184,N_12622,N_13552);
and U19185 (N_19185,N_12603,N_15968);
nand U19186 (N_19186,N_14573,N_13312);
nor U19187 (N_19187,N_14865,N_15044);
or U19188 (N_19188,N_13936,N_13897);
nand U19189 (N_19189,N_12692,N_14204);
or U19190 (N_19190,N_15851,N_12368);
or U19191 (N_19191,N_14599,N_13477);
or U19192 (N_19192,N_14734,N_12276);
or U19193 (N_19193,N_12103,N_14509);
nor U19194 (N_19194,N_12999,N_14367);
nand U19195 (N_19195,N_12962,N_13316);
nand U19196 (N_19196,N_13425,N_14957);
and U19197 (N_19197,N_15759,N_14808);
nor U19198 (N_19198,N_12618,N_12793);
and U19199 (N_19199,N_12514,N_15304);
nand U19200 (N_19200,N_12730,N_15379);
or U19201 (N_19201,N_13910,N_13030);
or U19202 (N_19202,N_15849,N_14865);
nor U19203 (N_19203,N_14079,N_12977);
and U19204 (N_19204,N_13663,N_14159);
and U19205 (N_19205,N_14708,N_12801);
and U19206 (N_19206,N_15557,N_13443);
and U19207 (N_19207,N_12869,N_12646);
nor U19208 (N_19208,N_13987,N_12316);
nor U19209 (N_19209,N_14893,N_13676);
or U19210 (N_19210,N_14617,N_15081);
and U19211 (N_19211,N_15391,N_13691);
or U19212 (N_19212,N_13525,N_12678);
and U19213 (N_19213,N_13046,N_14987);
nand U19214 (N_19214,N_14628,N_13004);
or U19215 (N_19215,N_12392,N_13905);
and U19216 (N_19216,N_12088,N_15348);
nand U19217 (N_19217,N_13288,N_12988);
or U19218 (N_19218,N_12789,N_14479);
nand U19219 (N_19219,N_13106,N_14207);
or U19220 (N_19220,N_12271,N_14600);
nor U19221 (N_19221,N_15213,N_13976);
or U19222 (N_19222,N_12607,N_15923);
nor U19223 (N_19223,N_15212,N_13704);
and U19224 (N_19224,N_15079,N_13825);
and U19225 (N_19225,N_12353,N_13873);
and U19226 (N_19226,N_14188,N_14056);
or U19227 (N_19227,N_15886,N_13669);
xnor U19228 (N_19228,N_12937,N_13502);
xnor U19229 (N_19229,N_12738,N_13410);
or U19230 (N_19230,N_15871,N_15683);
or U19231 (N_19231,N_12188,N_14367);
nand U19232 (N_19232,N_14669,N_14428);
nor U19233 (N_19233,N_14183,N_12834);
nor U19234 (N_19234,N_15768,N_12997);
nor U19235 (N_19235,N_14462,N_15992);
or U19236 (N_19236,N_12496,N_14976);
nand U19237 (N_19237,N_14638,N_13008);
and U19238 (N_19238,N_14934,N_12318);
nor U19239 (N_19239,N_12115,N_13806);
or U19240 (N_19240,N_14641,N_12123);
and U19241 (N_19241,N_14210,N_12080);
nor U19242 (N_19242,N_14802,N_15143);
nor U19243 (N_19243,N_12072,N_14825);
or U19244 (N_19244,N_12572,N_15928);
and U19245 (N_19245,N_15871,N_13198);
or U19246 (N_19246,N_15563,N_14664);
and U19247 (N_19247,N_13457,N_14454);
nand U19248 (N_19248,N_15743,N_15581);
nand U19249 (N_19249,N_12317,N_13840);
and U19250 (N_19250,N_13209,N_14196);
nand U19251 (N_19251,N_14613,N_12382);
nand U19252 (N_19252,N_15616,N_13120);
nand U19253 (N_19253,N_15096,N_13397);
nand U19254 (N_19254,N_15627,N_12436);
or U19255 (N_19255,N_13449,N_14514);
or U19256 (N_19256,N_14679,N_14623);
and U19257 (N_19257,N_14017,N_12681);
xor U19258 (N_19258,N_14732,N_15534);
nor U19259 (N_19259,N_14885,N_13164);
or U19260 (N_19260,N_14969,N_13617);
xor U19261 (N_19261,N_13768,N_13820);
or U19262 (N_19262,N_15414,N_12468);
or U19263 (N_19263,N_13711,N_13159);
and U19264 (N_19264,N_13552,N_15440);
nor U19265 (N_19265,N_13000,N_13812);
nand U19266 (N_19266,N_13517,N_13694);
nor U19267 (N_19267,N_14652,N_15802);
nor U19268 (N_19268,N_12188,N_12170);
or U19269 (N_19269,N_13055,N_12704);
and U19270 (N_19270,N_14298,N_13105);
xor U19271 (N_19271,N_14519,N_12572);
or U19272 (N_19272,N_13908,N_14992);
nand U19273 (N_19273,N_13381,N_12720);
or U19274 (N_19274,N_14191,N_14904);
nor U19275 (N_19275,N_14352,N_15237);
or U19276 (N_19276,N_13422,N_14216);
or U19277 (N_19277,N_14242,N_14096);
nand U19278 (N_19278,N_12262,N_15924);
and U19279 (N_19279,N_15679,N_15753);
or U19280 (N_19280,N_13773,N_13560);
nand U19281 (N_19281,N_13014,N_14606);
xnor U19282 (N_19282,N_13113,N_15311);
nand U19283 (N_19283,N_12656,N_14862);
xor U19284 (N_19284,N_14359,N_12680);
nor U19285 (N_19285,N_12390,N_15329);
and U19286 (N_19286,N_15100,N_13537);
nand U19287 (N_19287,N_13665,N_15621);
nand U19288 (N_19288,N_12590,N_13121);
nand U19289 (N_19289,N_12462,N_13922);
nor U19290 (N_19290,N_13550,N_13893);
nor U19291 (N_19291,N_15734,N_12476);
nor U19292 (N_19292,N_12343,N_14289);
nand U19293 (N_19293,N_14318,N_13865);
nand U19294 (N_19294,N_12565,N_14987);
and U19295 (N_19295,N_13411,N_13434);
nand U19296 (N_19296,N_15283,N_13551);
nor U19297 (N_19297,N_13062,N_13868);
nand U19298 (N_19298,N_15368,N_13197);
nand U19299 (N_19299,N_14649,N_15754);
or U19300 (N_19300,N_14551,N_13740);
or U19301 (N_19301,N_12829,N_15426);
and U19302 (N_19302,N_13673,N_12223);
or U19303 (N_19303,N_15886,N_14518);
nor U19304 (N_19304,N_12242,N_13676);
nor U19305 (N_19305,N_15534,N_15122);
and U19306 (N_19306,N_12135,N_13485);
nor U19307 (N_19307,N_12114,N_15126);
xor U19308 (N_19308,N_15152,N_12352);
and U19309 (N_19309,N_12116,N_12268);
and U19310 (N_19310,N_12472,N_12058);
nor U19311 (N_19311,N_15711,N_13976);
nor U19312 (N_19312,N_15692,N_12945);
nand U19313 (N_19313,N_13080,N_15376);
xnor U19314 (N_19314,N_13310,N_12309);
nand U19315 (N_19315,N_12559,N_15831);
or U19316 (N_19316,N_15780,N_14461);
or U19317 (N_19317,N_13638,N_14071);
nand U19318 (N_19318,N_12457,N_12586);
or U19319 (N_19319,N_12738,N_15149);
nor U19320 (N_19320,N_14745,N_14143);
and U19321 (N_19321,N_12811,N_14726);
and U19322 (N_19322,N_13167,N_15272);
nand U19323 (N_19323,N_14102,N_12027);
nor U19324 (N_19324,N_13792,N_12440);
nor U19325 (N_19325,N_12594,N_12009);
nor U19326 (N_19326,N_14983,N_14782);
nand U19327 (N_19327,N_13821,N_15756);
nor U19328 (N_19328,N_12180,N_13396);
nor U19329 (N_19329,N_15818,N_12238);
or U19330 (N_19330,N_14955,N_12258);
nand U19331 (N_19331,N_13926,N_15816);
nand U19332 (N_19332,N_12887,N_14663);
nand U19333 (N_19333,N_12558,N_13782);
nor U19334 (N_19334,N_15244,N_13697);
nor U19335 (N_19335,N_14403,N_13690);
nand U19336 (N_19336,N_15610,N_12802);
nand U19337 (N_19337,N_15494,N_14330);
nand U19338 (N_19338,N_15232,N_15513);
nand U19339 (N_19339,N_13567,N_15515);
and U19340 (N_19340,N_14661,N_13827);
nand U19341 (N_19341,N_15997,N_12431);
or U19342 (N_19342,N_12699,N_12304);
nor U19343 (N_19343,N_14068,N_12029);
and U19344 (N_19344,N_15678,N_15644);
nor U19345 (N_19345,N_12946,N_14692);
nor U19346 (N_19346,N_12296,N_15842);
xor U19347 (N_19347,N_15286,N_12916);
and U19348 (N_19348,N_12478,N_12391);
nor U19349 (N_19349,N_15515,N_15455);
nand U19350 (N_19350,N_15583,N_15049);
nor U19351 (N_19351,N_15997,N_13994);
nor U19352 (N_19352,N_15711,N_14144);
and U19353 (N_19353,N_14290,N_14197);
nor U19354 (N_19354,N_15512,N_14985);
nor U19355 (N_19355,N_14593,N_14312);
or U19356 (N_19356,N_13328,N_15577);
xnor U19357 (N_19357,N_13256,N_12030);
nand U19358 (N_19358,N_13104,N_15907);
nor U19359 (N_19359,N_13951,N_15378);
xnor U19360 (N_19360,N_13717,N_12329);
or U19361 (N_19361,N_15508,N_15562);
or U19362 (N_19362,N_13020,N_12437);
nand U19363 (N_19363,N_15225,N_13082);
xor U19364 (N_19364,N_15090,N_15112);
nor U19365 (N_19365,N_15066,N_12441);
xor U19366 (N_19366,N_13684,N_13186);
nor U19367 (N_19367,N_15110,N_15375);
or U19368 (N_19368,N_14775,N_14640);
and U19369 (N_19369,N_12430,N_15463);
or U19370 (N_19370,N_15369,N_15813);
xor U19371 (N_19371,N_13209,N_15458);
nor U19372 (N_19372,N_13246,N_15522);
nand U19373 (N_19373,N_13459,N_12469);
and U19374 (N_19374,N_14870,N_12274);
nand U19375 (N_19375,N_14935,N_13980);
and U19376 (N_19376,N_14021,N_12474);
nand U19377 (N_19377,N_15344,N_14573);
nand U19378 (N_19378,N_12202,N_13248);
and U19379 (N_19379,N_13039,N_14783);
nand U19380 (N_19380,N_13369,N_12356);
nand U19381 (N_19381,N_12241,N_15806);
or U19382 (N_19382,N_15441,N_15349);
and U19383 (N_19383,N_13217,N_12809);
nor U19384 (N_19384,N_13813,N_12725);
nand U19385 (N_19385,N_14160,N_13548);
or U19386 (N_19386,N_12930,N_14645);
xor U19387 (N_19387,N_15233,N_13714);
and U19388 (N_19388,N_12168,N_14761);
and U19389 (N_19389,N_14805,N_14065);
or U19390 (N_19390,N_14744,N_15150);
nand U19391 (N_19391,N_14284,N_12682);
nor U19392 (N_19392,N_13839,N_13118);
and U19393 (N_19393,N_14728,N_15674);
nand U19394 (N_19394,N_15867,N_15931);
nor U19395 (N_19395,N_15803,N_13788);
nand U19396 (N_19396,N_15052,N_15164);
and U19397 (N_19397,N_15293,N_13633);
or U19398 (N_19398,N_12653,N_14555);
nor U19399 (N_19399,N_14580,N_15366);
and U19400 (N_19400,N_15121,N_14954);
xnor U19401 (N_19401,N_14410,N_12322);
nand U19402 (N_19402,N_14172,N_13062);
xor U19403 (N_19403,N_14894,N_14592);
nand U19404 (N_19404,N_13596,N_13566);
or U19405 (N_19405,N_12303,N_13383);
xor U19406 (N_19406,N_12704,N_12514);
nand U19407 (N_19407,N_15745,N_15670);
nor U19408 (N_19408,N_15500,N_14544);
and U19409 (N_19409,N_14891,N_15437);
nand U19410 (N_19410,N_12109,N_15487);
xnor U19411 (N_19411,N_14934,N_14120);
or U19412 (N_19412,N_14558,N_13430);
xnor U19413 (N_19413,N_15027,N_15201);
nand U19414 (N_19414,N_15632,N_13354);
or U19415 (N_19415,N_14543,N_13616);
nand U19416 (N_19416,N_14063,N_12441);
and U19417 (N_19417,N_15255,N_14479);
and U19418 (N_19418,N_14639,N_15761);
nand U19419 (N_19419,N_15056,N_12081);
and U19420 (N_19420,N_13174,N_15610);
or U19421 (N_19421,N_14225,N_13364);
or U19422 (N_19422,N_15817,N_14140);
nand U19423 (N_19423,N_12388,N_13616);
or U19424 (N_19424,N_15381,N_13910);
nand U19425 (N_19425,N_14196,N_13387);
or U19426 (N_19426,N_12660,N_13884);
nand U19427 (N_19427,N_14831,N_13406);
nand U19428 (N_19428,N_13069,N_15691);
nand U19429 (N_19429,N_15204,N_12424);
or U19430 (N_19430,N_13535,N_12112);
or U19431 (N_19431,N_14798,N_12935);
and U19432 (N_19432,N_15335,N_13473);
nand U19433 (N_19433,N_12777,N_15064);
or U19434 (N_19434,N_13490,N_13670);
and U19435 (N_19435,N_14072,N_14750);
or U19436 (N_19436,N_15168,N_13251);
nor U19437 (N_19437,N_14472,N_14972);
nand U19438 (N_19438,N_15551,N_13142);
nor U19439 (N_19439,N_14970,N_14414);
and U19440 (N_19440,N_15293,N_13062);
nor U19441 (N_19441,N_14290,N_13901);
xor U19442 (N_19442,N_14308,N_12834);
nor U19443 (N_19443,N_12047,N_15671);
or U19444 (N_19444,N_15490,N_14563);
or U19445 (N_19445,N_15747,N_13938);
or U19446 (N_19446,N_13026,N_13908);
nand U19447 (N_19447,N_14034,N_14140);
nor U19448 (N_19448,N_15202,N_15221);
and U19449 (N_19449,N_13480,N_12812);
nand U19450 (N_19450,N_14803,N_13068);
xnor U19451 (N_19451,N_15953,N_15647);
nand U19452 (N_19452,N_14339,N_15010);
nand U19453 (N_19453,N_12923,N_12963);
or U19454 (N_19454,N_12402,N_12415);
and U19455 (N_19455,N_12159,N_12613);
nor U19456 (N_19456,N_13147,N_14828);
nor U19457 (N_19457,N_13284,N_14329);
nor U19458 (N_19458,N_15540,N_14417);
or U19459 (N_19459,N_12635,N_13931);
or U19460 (N_19460,N_14063,N_13329);
nand U19461 (N_19461,N_14590,N_13966);
or U19462 (N_19462,N_14449,N_12489);
nor U19463 (N_19463,N_14050,N_15495);
and U19464 (N_19464,N_14380,N_14586);
nor U19465 (N_19465,N_13696,N_14082);
xnor U19466 (N_19466,N_12852,N_15325);
or U19467 (N_19467,N_12428,N_13541);
nand U19468 (N_19468,N_13647,N_13490);
nand U19469 (N_19469,N_12194,N_12262);
or U19470 (N_19470,N_13766,N_13632);
or U19471 (N_19471,N_13096,N_14581);
or U19472 (N_19472,N_13948,N_12332);
and U19473 (N_19473,N_14742,N_12460);
or U19474 (N_19474,N_15679,N_12786);
and U19475 (N_19475,N_14328,N_13127);
nand U19476 (N_19476,N_14760,N_14045);
or U19477 (N_19477,N_12959,N_12388);
nand U19478 (N_19478,N_13621,N_15845);
and U19479 (N_19479,N_12671,N_14868);
nor U19480 (N_19480,N_14619,N_13278);
nor U19481 (N_19481,N_12952,N_13683);
xor U19482 (N_19482,N_14515,N_12885);
nand U19483 (N_19483,N_14639,N_12978);
nor U19484 (N_19484,N_15335,N_14128);
nor U19485 (N_19485,N_12610,N_15672);
and U19486 (N_19486,N_13628,N_13033);
xor U19487 (N_19487,N_14006,N_14913);
nand U19488 (N_19488,N_13878,N_12798);
nor U19489 (N_19489,N_12959,N_12063);
nor U19490 (N_19490,N_12916,N_13451);
nand U19491 (N_19491,N_15103,N_12813);
xnor U19492 (N_19492,N_13669,N_13212);
or U19493 (N_19493,N_12639,N_12047);
or U19494 (N_19494,N_12659,N_14332);
xor U19495 (N_19495,N_12575,N_13521);
and U19496 (N_19496,N_13788,N_15048);
and U19497 (N_19497,N_15471,N_14331);
nor U19498 (N_19498,N_12300,N_14642);
and U19499 (N_19499,N_15748,N_14753);
and U19500 (N_19500,N_15010,N_15804);
and U19501 (N_19501,N_15133,N_15454);
and U19502 (N_19502,N_15649,N_13711);
nor U19503 (N_19503,N_13936,N_12217);
and U19504 (N_19504,N_12583,N_13721);
nor U19505 (N_19505,N_14138,N_13319);
and U19506 (N_19506,N_14774,N_14020);
or U19507 (N_19507,N_12215,N_14250);
xor U19508 (N_19508,N_12468,N_12072);
or U19509 (N_19509,N_15075,N_12913);
nor U19510 (N_19510,N_13831,N_15774);
xor U19511 (N_19511,N_13765,N_12778);
and U19512 (N_19512,N_13524,N_14774);
and U19513 (N_19513,N_14127,N_12780);
and U19514 (N_19514,N_12168,N_12553);
nor U19515 (N_19515,N_14239,N_13045);
nand U19516 (N_19516,N_14158,N_14589);
nand U19517 (N_19517,N_15524,N_13904);
or U19518 (N_19518,N_15378,N_14923);
or U19519 (N_19519,N_15743,N_14650);
nor U19520 (N_19520,N_13981,N_13703);
or U19521 (N_19521,N_12785,N_15503);
nor U19522 (N_19522,N_15333,N_13231);
and U19523 (N_19523,N_13397,N_15755);
nor U19524 (N_19524,N_13018,N_14316);
or U19525 (N_19525,N_15810,N_12419);
and U19526 (N_19526,N_12466,N_15042);
nor U19527 (N_19527,N_14917,N_12343);
xor U19528 (N_19528,N_13658,N_15576);
and U19529 (N_19529,N_15242,N_15452);
or U19530 (N_19530,N_14888,N_15825);
and U19531 (N_19531,N_15810,N_14719);
or U19532 (N_19532,N_12156,N_15477);
or U19533 (N_19533,N_12384,N_15702);
or U19534 (N_19534,N_13426,N_15505);
or U19535 (N_19535,N_12319,N_12906);
nor U19536 (N_19536,N_12564,N_12134);
nand U19537 (N_19537,N_13806,N_12407);
or U19538 (N_19538,N_13994,N_15424);
and U19539 (N_19539,N_13544,N_14443);
nand U19540 (N_19540,N_12852,N_13357);
nand U19541 (N_19541,N_13912,N_14935);
xor U19542 (N_19542,N_13869,N_15537);
xnor U19543 (N_19543,N_12424,N_15215);
nor U19544 (N_19544,N_14421,N_15844);
nand U19545 (N_19545,N_15175,N_14358);
and U19546 (N_19546,N_15682,N_13588);
nor U19547 (N_19547,N_13889,N_15066);
or U19548 (N_19548,N_14741,N_15441);
nand U19549 (N_19549,N_13868,N_12386);
nand U19550 (N_19550,N_14770,N_15943);
nor U19551 (N_19551,N_14192,N_12769);
nor U19552 (N_19552,N_12395,N_12747);
nor U19553 (N_19553,N_15855,N_14030);
nor U19554 (N_19554,N_12936,N_14870);
nand U19555 (N_19555,N_14300,N_15977);
nand U19556 (N_19556,N_12498,N_15607);
or U19557 (N_19557,N_12378,N_14632);
or U19558 (N_19558,N_12174,N_13253);
or U19559 (N_19559,N_13366,N_14976);
nor U19560 (N_19560,N_15469,N_12622);
and U19561 (N_19561,N_12336,N_12196);
or U19562 (N_19562,N_14146,N_14753);
and U19563 (N_19563,N_15194,N_14736);
and U19564 (N_19564,N_14111,N_15284);
or U19565 (N_19565,N_13674,N_12010);
and U19566 (N_19566,N_14720,N_12289);
and U19567 (N_19567,N_12553,N_13741);
nor U19568 (N_19568,N_15112,N_15307);
or U19569 (N_19569,N_15225,N_13699);
nand U19570 (N_19570,N_15118,N_14066);
xor U19571 (N_19571,N_12574,N_12357);
nor U19572 (N_19572,N_13024,N_13015);
and U19573 (N_19573,N_15001,N_15850);
and U19574 (N_19574,N_13934,N_14737);
nand U19575 (N_19575,N_13413,N_13014);
or U19576 (N_19576,N_14391,N_15396);
and U19577 (N_19577,N_12368,N_12592);
or U19578 (N_19578,N_15521,N_14333);
nand U19579 (N_19579,N_15068,N_12971);
xor U19580 (N_19580,N_13713,N_14843);
and U19581 (N_19581,N_14172,N_15328);
or U19582 (N_19582,N_13527,N_15671);
and U19583 (N_19583,N_14453,N_12796);
nor U19584 (N_19584,N_13575,N_12446);
or U19585 (N_19585,N_13053,N_15303);
and U19586 (N_19586,N_12004,N_14349);
or U19587 (N_19587,N_15195,N_15469);
xnor U19588 (N_19588,N_14695,N_14854);
or U19589 (N_19589,N_15200,N_12560);
nand U19590 (N_19590,N_15804,N_15921);
nor U19591 (N_19591,N_14456,N_14229);
and U19592 (N_19592,N_15833,N_15031);
and U19593 (N_19593,N_15359,N_14570);
and U19594 (N_19594,N_12588,N_15593);
xor U19595 (N_19595,N_15547,N_14701);
nand U19596 (N_19596,N_13836,N_15718);
and U19597 (N_19597,N_15105,N_15145);
xnor U19598 (N_19598,N_13389,N_15952);
nor U19599 (N_19599,N_13837,N_14336);
or U19600 (N_19600,N_12792,N_12208);
or U19601 (N_19601,N_13676,N_12799);
and U19602 (N_19602,N_15720,N_15590);
nor U19603 (N_19603,N_13972,N_14980);
nor U19604 (N_19604,N_13800,N_12623);
and U19605 (N_19605,N_14174,N_12912);
nand U19606 (N_19606,N_14514,N_13370);
or U19607 (N_19607,N_14704,N_15760);
nand U19608 (N_19608,N_13125,N_15966);
nand U19609 (N_19609,N_13841,N_15670);
and U19610 (N_19610,N_15113,N_15281);
nor U19611 (N_19611,N_14212,N_15502);
and U19612 (N_19612,N_15989,N_15723);
nand U19613 (N_19613,N_12120,N_13981);
or U19614 (N_19614,N_13763,N_13951);
nand U19615 (N_19615,N_15899,N_14076);
nand U19616 (N_19616,N_12878,N_13988);
nand U19617 (N_19617,N_15291,N_15063);
or U19618 (N_19618,N_12721,N_15902);
or U19619 (N_19619,N_12813,N_13070);
and U19620 (N_19620,N_12394,N_14397);
and U19621 (N_19621,N_12855,N_12197);
and U19622 (N_19622,N_15846,N_14906);
xor U19623 (N_19623,N_13282,N_12722);
xor U19624 (N_19624,N_12646,N_14780);
and U19625 (N_19625,N_13229,N_12395);
nand U19626 (N_19626,N_14660,N_13981);
nand U19627 (N_19627,N_15095,N_13222);
and U19628 (N_19628,N_12524,N_14413);
nor U19629 (N_19629,N_14082,N_12197);
xor U19630 (N_19630,N_13392,N_14776);
and U19631 (N_19631,N_13060,N_12248);
and U19632 (N_19632,N_14951,N_13597);
nor U19633 (N_19633,N_15297,N_15741);
nor U19634 (N_19634,N_13288,N_12270);
nand U19635 (N_19635,N_14262,N_15134);
nand U19636 (N_19636,N_14632,N_14559);
and U19637 (N_19637,N_12585,N_13532);
nand U19638 (N_19638,N_13627,N_12597);
nand U19639 (N_19639,N_15304,N_15227);
and U19640 (N_19640,N_14172,N_13849);
xnor U19641 (N_19641,N_12419,N_15966);
nor U19642 (N_19642,N_13648,N_15670);
or U19643 (N_19643,N_15399,N_14123);
and U19644 (N_19644,N_12647,N_15615);
nand U19645 (N_19645,N_14210,N_15873);
nor U19646 (N_19646,N_13590,N_12072);
or U19647 (N_19647,N_13507,N_13136);
nand U19648 (N_19648,N_12731,N_14415);
xnor U19649 (N_19649,N_15631,N_12489);
and U19650 (N_19650,N_14179,N_15972);
and U19651 (N_19651,N_13437,N_14732);
or U19652 (N_19652,N_15923,N_14019);
or U19653 (N_19653,N_12642,N_13829);
nand U19654 (N_19654,N_14904,N_15980);
nand U19655 (N_19655,N_12929,N_12666);
nor U19656 (N_19656,N_13385,N_15864);
nor U19657 (N_19657,N_14268,N_12106);
or U19658 (N_19658,N_13722,N_14091);
and U19659 (N_19659,N_15176,N_15429);
nor U19660 (N_19660,N_12948,N_13231);
or U19661 (N_19661,N_12874,N_12270);
nand U19662 (N_19662,N_14315,N_14916);
or U19663 (N_19663,N_15356,N_13072);
or U19664 (N_19664,N_15911,N_12874);
nor U19665 (N_19665,N_15448,N_13234);
nor U19666 (N_19666,N_13027,N_13192);
and U19667 (N_19667,N_14453,N_14050);
and U19668 (N_19668,N_15766,N_15369);
nor U19669 (N_19669,N_12916,N_14013);
nor U19670 (N_19670,N_15821,N_12662);
nand U19671 (N_19671,N_15696,N_13686);
xnor U19672 (N_19672,N_15557,N_14123);
or U19673 (N_19673,N_14797,N_12270);
and U19674 (N_19674,N_15267,N_15452);
nor U19675 (N_19675,N_13190,N_14038);
nor U19676 (N_19676,N_13282,N_12852);
nor U19677 (N_19677,N_14110,N_13281);
or U19678 (N_19678,N_15001,N_15496);
and U19679 (N_19679,N_14934,N_15242);
xor U19680 (N_19680,N_13892,N_15128);
nor U19681 (N_19681,N_13541,N_13374);
or U19682 (N_19682,N_13114,N_14404);
or U19683 (N_19683,N_12951,N_12186);
or U19684 (N_19684,N_15548,N_14748);
nand U19685 (N_19685,N_13260,N_15561);
nor U19686 (N_19686,N_14128,N_13169);
nor U19687 (N_19687,N_14377,N_14990);
nand U19688 (N_19688,N_12439,N_15078);
and U19689 (N_19689,N_15323,N_12632);
and U19690 (N_19690,N_14391,N_13412);
nand U19691 (N_19691,N_15099,N_12418);
nand U19692 (N_19692,N_12835,N_14990);
xnor U19693 (N_19693,N_13796,N_14275);
xor U19694 (N_19694,N_13784,N_13421);
or U19695 (N_19695,N_14901,N_13066);
nor U19696 (N_19696,N_13611,N_14991);
xnor U19697 (N_19697,N_12675,N_13344);
nor U19698 (N_19698,N_15930,N_12911);
nand U19699 (N_19699,N_14203,N_13034);
xor U19700 (N_19700,N_15285,N_15992);
or U19701 (N_19701,N_12455,N_12799);
nand U19702 (N_19702,N_12852,N_12381);
nand U19703 (N_19703,N_14649,N_15056);
or U19704 (N_19704,N_13302,N_15176);
or U19705 (N_19705,N_15793,N_15357);
nor U19706 (N_19706,N_15566,N_12153);
or U19707 (N_19707,N_15304,N_13101);
or U19708 (N_19708,N_12715,N_14346);
or U19709 (N_19709,N_15869,N_13583);
nand U19710 (N_19710,N_13279,N_14111);
and U19711 (N_19711,N_14117,N_14498);
nor U19712 (N_19712,N_13137,N_15374);
nand U19713 (N_19713,N_14265,N_13431);
or U19714 (N_19714,N_14027,N_14700);
nor U19715 (N_19715,N_14521,N_14349);
or U19716 (N_19716,N_13648,N_13034);
nor U19717 (N_19717,N_13670,N_14531);
and U19718 (N_19718,N_14614,N_13807);
or U19719 (N_19719,N_13220,N_12559);
nand U19720 (N_19720,N_14130,N_12605);
and U19721 (N_19721,N_15893,N_14290);
nand U19722 (N_19722,N_13905,N_12472);
nand U19723 (N_19723,N_12410,N_15748);
nand U19724 (N_19724,N_12100,N_14056);
or U19725 (N_19725,N_12699,N_12665);
or U19726 (N_19726,N_13623,N_14100);
or U19727 (N_19727,N_15398,N_14248);
nor U19728 (N_19728,N_12282,N_12118);
or U19729 (N_19729,N_13293,N_12277);
or U19730 (N_19730,N_15200,N_13468);
nand U19731 (N_19731,N_14050,N_13215);
nand U19732 (N_19732,N_15386,N_14694);
xnor U19733 (N_19733,N_13492,N_14907);
nor U19734 (N_19734,N_12065,N_15467);
or U19735 (N_19735,N_15770,N_15284);
and U19736 (N_19736,N_13545,N_12879);
and U19737 (N_19737,N_14244,N_14697);
nor U19738 (N_19738,N_15690,N_13303);
or U19739 (N_19739,N_15942,N_12892);
and U19740 (N_19740,N_12798,N_13386);
or U19741 (N_19741,N_12332,N_13136);
nor U19742 (N_19742,N_12400,N_12300);
and U19743 (N_19743,N_13869,N_13151);
and U19744 (N_19744,N_14142,N_14306);
and U19745 (N_19745,N_14429,N_15146);
nor U19746 (N_19746,N_13508,N_14160);
nor U19747 (N_19747,N_15924,N_12387);
xor U19748 (N_19748,N_14191,N_13093);
and U19749 (N_19749,N_14026,N_14755);
or U19750 (N_19750,N_12607,N_12641);
nand U19751 (N_19751,N_14187,N_14383);
or U19752 (N_19752,N_12494,N_15241);
nand U19753 (N_19753,N_12750,N_12709);
nand U19754 (N_19754,N_14160,N_14820);
nor U19755 (N_19755,N_13383,N_14425);
nand U19756 (N_19756,N_15818,N_13131);
nand U19757 (N_19757,N_14815,N_13496);
nand U19758 (N_19758,N_12676,N_13269);
or U19759 (N_19759,N_13718,N_14336);
and U19760 (N_19760,N_13419,N_14065);
nor U19761 (N_19761,N_15591,N_12410);
nor U19762 (N_19762,N_15873,N_14515);
xor U19763 (N_19763,N_15093,N_14165);
and U19764 (N_19764,N_13790,N_14178);
nand U19765 (N_19765,N_13713,N_12259);
or U19766 (N_19766,N_15233,N_13638);
or U19767 (N_19767,N_14427,N_13283);
or U19768 (N_19768,N_13232,N_12144);
nand U19769 (N_19769,N_15044,N_14169);
nor U19770 (N_19770,N_15391,N_12030);
or U19771 (N_19771,N_14498,N_14847);
or U19772 (N_19772,N_13705,N_14092);
nand U19773 (N_19773,N_13096,N_12015);
and U19774 (N_19774,N_13394,N_12178);
xor U19775 (N_19775,N_12643,N_13741);
or U19776 (N_19776,N_13525,N_15820);
nor U19777 (N_19777,N_13993,N_12344);
or U19778 (N_19778,N_14556,N_13364);
and U19779 (N_19779,N_15549,N_12873);
nand U19780 (N_19780,N_15586,N_12849);
nand U19781 (N_19781,N_13889,N_14278);
or U19782 (N_19782,N_12743,N_14955);
or U19783 (N_19783,N_12391,N_14057);
nor U19784 (N_19784,N_12863,N_15534);
nor U19785 (N_19785,N_13373,N_13237);
nand U19786 (N_19786,N_13875,N_13873);
and U19787 (N_19787,N_13195,N_13702);
nor U19788 (N_19788,N_12716,N_15875);
xor U19789 (N_19789,N_12930,N_13688);
nor U19790 (N_19790,N_14677,N_12265);
or U19791 (N_19791,N_13925,N_13673);
or U19792 (N_19792,N_12079,N_12174);
and U19793 (N_19793,N_12228,N_15174);
and U19794 (N_19794,N_13530,N_14118);
or U19795 (N_19795,N_13506,N_12366);
nor U19796 (N_19796,N_13785,N_13307);
and U19797 (N_19797,N_15082,N_12302);
and U19798 (N_19798,N_13875,N_15645);
or U19799 (N_19799,N_12187,N_13013);
and U19800 (N_19800,N_14364,N_12132);
nor U19801 (N_19801,N_14477,N_13923);
and U19802 (N_19802,N_12745,N_15141);
and U19803 (N_19803,N_14385,N_14397);
and U19804 (N_19804,N_13746,N_13556);
nand U19805 (N_19805,N_13242,N_15148);
or U19806 (N_19806,N_13171,N_15855);
xor U19807 (N_19807,N_15425,N_15151);
nor U19808 (N_19808,N_12892,N_14693);
xor U19809 (N_19809,N_12082,N_12941);
nor U19810 (N_19810,N_15399,N_15044);
and U19811 (N_19811,N_13418,N_12067);
nor U19812 (N_19812,N_14436,N_14983);
and U19813 (N_19813,N_14127,N_12325);
or U19814 (N_19814,N_13584,N_13443);
nor U19815 (N_19815,N_12495,N_15606);
nand U19816 (N_19816,N_12477,N_13797);
nor U19817 (N_19817,N_12696,N_13479);
nor U19818 (N_19818,N_14834,N_13570);
xor U19819 (N_19819,N_14450,N_15292);
nor U19820 (N_19820,N_13647,N_13587);
nor U19821 (N_19821,N_13977,N_12650);
nand U19822 (N_19822,N_14971,N_15015);
xor U19823 (N_19823,N_15266,N_12838);
nor U19824 (N_19824,N_15116,N_13648);
nor U19825 (N_19825,N_14376,N_12162);
nor U19826 (N_19826,N_14572,N_12131);
nor U19827 (N_19827,N_15648,N_13768);
and U19828 (N_19828,N_14449,N_13439);
nor U19829 (N_19829,N_15907,N_15333);
or U19830 (N_19830,N_13740,N_13586);
and U19831 (N_19831,N_14133,N_15559);
or U19832 (N_19832,N_12731,N_15683);
nor U19833 (N_19833,N_15450,N_14956);
or U19834 (N_19834,N_12458,N_14132);
nor U19835 (N_19835,N_12634,N_15547);
or U19836 (N_19836,N_15350,N_13824);
nand U19837 (N_19837,N_15073,N_12084);
or U19838 (N_19838,N_15109,N_15736);
or U19839 (N_19839,N_14191,N_12410);
or U19840 (N_19840,N_15688,N_14555);
nand U19841 (N_19841,N_13102,N_12764);
and U19842 (N_19842,N_12273,N_13353);
and U19843 (N_19843,N_13430,N_15337);
or U19844 (N_19844,N_13121,N_12139);
nand U19845 (N_19845,N_12909,N_12432);
and U19846 (N_19846,N_13002,N_14240);
and U19847 (N_19847,N_14446,N_13148);
nand U19848 (N_19848,N_14911,N_12794);
and U19849 (N_19849,N_13758,N_15700);
xor U19850 (N_19850,N_12375,N_13546);
or U19851 (N_19851,N_13105,N_13276);
and U19852 (N_19852,N_15743,N_15848);
or U19853 (N_19853,N_12954,N_15200);
or U19854 (N_19854,N_15593,N_12433);
nand U19855 (N_19855,N_14431,N_14584);
nor U19856 (N_19856,N_12663,N_15214);
and U19857 (N_19857,N_13347,N_12091);
nor U19858 (N_19858,N_14453,N_12356);
nand U19859 (N_19859,N_14103,N_13616);
or U19860 (N_19860,N_13917,N_15836);
and U19861 (N_19861,N_13363,N_13010);
nor U19862 (N_19862,N_15549,N_14923);
nand U19863 (N_19863,N_12261,N_12474);
xor U19864 (N_19864,N_12467,N_14464);
nand U19865 (N_19865,N_12932,N_14352);
nor U19866 (N_19866,N_13495,N_12615);
nand U19867 (N_19867,N_15727,N_12076);
nand U19868 (N_19868,N_12298,N_15631);
nor U19869 (N_19869,N_15825,N_14774);
or U19870 (N_19870,N_14115,N_15081);
or U19871 (N_19871,N_14909,N_14841);
nor U19872 (N_19872,N_14529,N_12621);
nand U19873 (N_19873,N_13929,N_15340);
nand U19874 (N_19874,N_15245,N_12008);
or U19875 (N_19875,N_14027,N_14758);
and U19876 (N_19876,N_12985,N_12031);
xor U19877 (N_19877,N_15497,N_15878);
nor U19878 (N_19878,N_15217,N_12208);
nor U19879 (N_19879,N_14044,N_13623);
or U19880 (N_19880,N_13758,N_14283);
and U19881 (N_19881,N_14618,N_12247);
nor U19882 (N_19882,N_12563,N_13405);
or U19883 (N_19883,N_12623,N_14403);
nor U19884 (N_19884,N_15172,N_13479);
and U19885 (N_19885,N_14594,N_12127);
nand U19886 (N_19886,N_14316,N_14619);
nor U19887 (N_19887,N_15058,N_14955);
nor U19888 (N_19888,N_14269,N_12992);
nand U19889 (N_19889,N_12764,N_14835);
nand U19890 (N_19890,N_13347,N_14840);
nor U19891 (N_19891,N_15424,N_13078);
or U19892 (N_19892,N_14298,N_15427);
nor U19893 (N_19893,N_15564,N_14338);
nand U19894 (N_19894,N_12214,N_14633);
xnor U19895 (N_19895,N_14340,N_15329);
or U19896 (N_19896,N_15598,N_13261);
nor U19897 (N_19897,N_14846,N_14709);
nor U19898 (N_19898,N_13705,N_14636);
or U19899 (N_19899,N_14919,N_13650);
nand U19900 (N_19900,N_13087,N_12618);
nor U19901 (N_19901,N_12674,N_13053);
and U19902 (N_19902,N_15931,N_13859);
nand U19903 (N_19903,N_15640,N_15031);
nand U19904 (N_19904,N_13752,N_14514);
nor U19905 (N_19905,N_12772,N_13828);
nor U19906 (N_19906,N_15175,N_15193);
or U19907 (N_19907,N_12858,N_15192);
nand U19908 (N_19908,N_12373,N_15599);
and U19909 (N_19909,N_13581,N_12762);
or U19910 (N_19910,N_14170,N_14900);
or U19911 (N_19911,N_15250,N_14199);
or U19912 (N_19912,N_13134,N_15146);
nor U19913 (N_19913,N_15450,N_14463);
nor U19914 (N_19914,N_15494,N_13832);
nor U19915 (N_19915,N_13479,N_14339);
nor U19916 (N_19916,N_13395,N_13011);
or U19917 (N_19917,N_12624,N_13171);
nor U19918 (N_19918,N_15735,N_12351);
or U19919 (N_19919,N_12692,N_14831);
xnor U19920 (N_19920,N_15857,N_13442);
xor U19921 (N_19921,N_14179,N_13985);
nand U19922 (N_19922,N_14877,N_12946);
nand U19923 (N_19923,N_14879,N_14962);
or U19924 (N_19924,N_14714,N_13932);
nor U19925 (N_19925,N_14470,N_12771);
nand U19926 (N_19926,N_14353,N_14556);
and U19927 (N_19927,N_12567,N_13108);
nor U19928 (N_19928,N_13425,N_14297);
and U19929 (N_19929,N_13581,N_14652);
or U19930 (N_19930,N_14895,N_14143);
nand U19931 (N_19931,N_14918,N_12213);
and U19932 (N_19932,N_14777,N_13313);
and U19933 (N_19933,N_15985,N_14500);
or U19934 (N_19934,N_14400,N_12008);
xnor U19935 (N_19935,N_14771,N_14095);
nor U19936 (N_19936,N_12122,N_15049);
and U19937 (N_19937,N_15522,N_13140);
nor U19938 (N_19938,N_15772,N_13136);
xor U19939 (N_19939,N_15183,N_14296);
xor U19940 (N_19940,N_14727,N_15120);
nor U19941 (N_19941,N_12212,N_14751);
nand U19942 (N_19942,N_14629,N_12491);
and U19943 (N_19943,N_14693,N_12268);
nand U19944 (N_19944,N_12403,N_15980);
nand U19945 (N_19945,N_14526,N_15967);
nand U19946 (N_19946,N_15643,N_12229);
or U19947 (N_19947,N_12504,N_15378);
nor U19948 (N_19948,N_14610,N_13158);
nand U19949 (N_19949,N_15959,N_15767);
nor U19950 (N_19950,N_14364,N_13096);
and U19951 (N_19951,N_12149,N_13151);
and U19952 (N_19952,N_13263,N_13836);
nor U19953 (N_19953,N_15224,N_15978);
or U19954 (N_19954,N_12103,N_15075);
or U19955 (N_19955,N_12674,N_13407);
nor U19956 (N_19956,N_13301,N_15248);
and U19957 (N_19957,N_15185,N_12047);
nor U19958 (N_19958,N_13154,N_15061);
nor U19959 (N_19959,N_12642,N_15478);
or U19960 (N_19960,N_12822,N_12077);
nor U19961 (N_19961,N_13911,N_14829);
and U19962 (N_19962,N_14777,N_12438);
nand U19963 (N_19963,N_14505,N_14408);
nand U19964 (N_19964,N_13308,N_14044);
or U19965 (N_19965,N_12132,N_12652);
nor U19966 (N_19966,N_15906,N_12162);
or U19967 (N_19967,N_12610,N_15103);
or U19968 (N_19968,N_15400,N_14210);
xor U19969 (N_19969,N_12270,N_13407);
xnor U19970 (N_19970,N_13641,N_15556);
or U19971 (N_19971,N_14321,N_15514);
xnor U19972 (N_19972,N_13807,N_12006);
nor U19973 (N_19973,N_15739,N_12350);
nand U19974 (N_19974,N_14185,N_13996);
nand U19975 (N_19975,N_13787,N_13895);
and U19976 (N_19976,N_12173,N_15410);
xor U19977 (N_19977,N_12291,N_13186);
xnor U19978 (N_19978,N_12650,N_12213);
nor U19979 (N_19979,N_14968,N_13214);
xor U19980 (N_19980,N_15106,N_13958);
and U19981 (N_19981,N_14442,N_14489);
nor U19982 (N_19982,N_15827,N_14282);
or U19983 (N_19983,N_15935,N_12033);
and U19984 (N_19984,N_14377,N_12856);
and U19985 (N_19985,N_12602,N_15111);
nor U19986 (N_19986,N_12781,N_14796);
nand U19987 (N_19987,N_14802,N_13956);
or U19988 (N_19988,N_12803,N_14687);
and U19989 (N_19989,N_13045,N_14097);
nor U19990 (N_19990,N_14050,N_15013);
or U19991 (N_19991,N_13860,N_12539);
and U19992 (N_19992,N_14260,N_14828);
and U19993 (N_19993,N_15309,N_13127);
nor U19994 (N_19994,N_15107,N_13145);
or U19995 (N_19995,N_12784,N_13258);
xor U19996 (N_19996,N_12012,N_13847);
nand U19997 (N_19997,N_15687,N_13168);
nor U19998 (N_19998,N_12664,N_13800);
xnor U19999 (N_19999,N_14497,N_15355);
nor UO_0 (O_0,N_16173,N_16930);
xnor UO_1 (O_1,N_19271,N_18713);
or UO_2 (O_2,N_18269,N_16517);
and UO_3 (O_3,N_16544,N_17339);
and UO_4 (O_4,N_16105,N_17030);
nand UO_5 (O_5,N_18824,N_16264);
nor UO_6 (O_6,N_16942,N_16803);
or UO_7 (O_7,N_19021,N_18700);
nand UO_8 (O_8,N_18232,N_18237);
nor UO_9 (O_9,N_18772,N_19093);
nor UO_10 (O_10,N_16807,N_18317);
or UO_11 (O_11,N_19162,N_16669);
or UO_12 (O_12,N_18021,N_16156);
nand UO_13 (O_13,N_19932,N_16553);
and UO_14 (O_14,N_17883,N_18123);
nand UO_15 (O_15,N_19365,N_19290);
or UO_16 (O_16,N_17548,N_18478);
or UO_17 (O_17,N_18922,N_19265);
and UO_18 (O_18,N_19600,N_16664);
nand UO_19 (O_19,N_17923,N_19546);
or UO_20 (O_20,N_18231,N_18835);
xnor UO_21 (O_21,N_18813,N_19660);
nor UO_22 (O_22,N_18593,N_16355);
nand UO_23 (O_23,N_16232,N_17155);
nor UO_24 (O_24,N_19917,N_17097);
nand UO_25 (O_25,N_17704,N_18843);
xor UO_26 (O_26,N_17696,N_18572);
nor UO_27 (O_27,N_17552,N_16768);
and UO_28 (O_28,N_17145,N_19124);
or UO_29 (O_29,N_19533,N_19159);
nor UO_30 (O_30,N_19618,N_17723);
xor UO_31 (O_31,N_18646,N_16988);
nand UO_32 (O_32,N_17921,N_19389);
nand UO_33 (O_33,N_16361,N_19341);
and UO_34 (O_34,N_18815,N_16075);
nand UO_35 (O_35,N_19530,N_17002);
xnor UO_36 (O_36,N_16437,N_16837);
nor UO_37 (O_37,N_19853,N_16009);
nor UO_38 (O_38,N_19218,N_17112);
or UO_39 (O_39,N_18740,N_17639);
and UO_40 (O_40,N_18717,N_19592);
xnor UO_41 (O_41,N_18250,N_19339);
nand UO_42 (O_42,N_18156,N_19992);
and UO_43 (O_43,N_16711,N_16178);
xnor UO_44 (O_44,N_17091,N_19032);
or UO_45 (O_45,N_18629,N_17175);
or UO_46 (O_46,N_19013,N_19805);
nor UO_47 (O_47,N_17266,N_17806);
nand UO_48 (O_48,N_17858,N_18540);
or UO_49 (O_49,N_18457,N_17259);
and UO_50 (O_50,N_18497,N_17865);
or UO_51 (O_51,N_17746,N_19971);
nor UO_52 (O_52,N_16744,N_18805);
or UO_53 (O_53,N_17184,N_16545);
or UO_54 (O_54,N_16184,N_17942);
nor UO_55 (O_55,N_19369,N_18295);
nand UO_56 (O_56,N_18588,N_19423);
or UO_57 (O_57,N_19869,N_18053);
nand UO_58 (O_58,N_18175,N_19641);
and UO_59 (O_59,N_16706,N_19145);
or UO_60 (O_60,N_18761,N_17785);
and UO_61 (O_61,N_19611,N_18468);
and UO_62 (O_62,N_19567,N_18149);
nor UO_63 (O_63,N_16190,N_18146);
nand UO_64 (O_64,N_18388,N_17692);
nor UO_65 (O_65,N_18715,N_16720);
nand UO_66 (O_66,N_17514,N_18755);
xor UO_67 (O_67,N_18638,N_19571);
nor UO_68 (O_68,N_16113,N_18222);
or UO_69 (O_69,N_16533,N_17345);
or UO_70 (O_70,N_19380,N_16030);
nand UO_71 (O_71,N_17509,N_19368);
nand UO_72 (O_72,N_18644,N_18698);
or UO_73 (O_73,N_16712,N_18329);
xor UO_74 (O_74,N_17636,N_16295);
and UO_75 (O_75,N_17436,N_18863);
or UO_76 (O_76,N_19422,N_18686);
xnor UO_77 (O_77,N_19373,N_19163);
and UO_78 (O_78,N_19781,N_17740);
and UO_79 (O_79,N_18613,N_18058);
and UO_80 (O_80,N_19460,N_17732);
xor UO_81 (O_81,N_18716,N_16569);
and UO_82 (O_82,N_16996,N_18256);
nand UO_83 (O_83,N_18406,N_19889);
nor UO_84 (O_84,N_16230,N_18547);
and UO_85 (O_85,N_16261,N_16426);
nor UO_86 (O_86,N_18080,N_19718);
and UO_87 (O_87,N_17773,N_19830);
nand UO_88 (O_88,N_18958,N_17721);
nor UO_89 (O_89,N_17620,N_16035);
xnor UO_90 (O_90,N_18465,N_18886);
nor UO_91 (O_91,N_19065,N_16096);
and UO_92 (O_92,N_18748,N_17432);
or UO_93 (O_93,N_17497,N_16299);
or UO_94 (O_94,N_17842,N_19721);
nor UO_95 (O_95,N_17351,N_19736);
xor UO_96 (O_96,N_17530,N_17465);
and UO_97 (O_97,N_19578,N_17458);
xnor UO_98 (O_98,N_19964,N_16459);
or UO_99 (O_99,N_18214,N_18801);
or UO_100 (O_100,N_18535,N_17000);
xnor UO_101 (O_101,N_16871,N_16463);
xor UO_102 (O_102,N_18703,N_18320);
nand UO_103 (O_103,N_18020,N_18305);
or UO_104 (O_104,N_19114,N_18890);
or UO_105 (O_105,N_17838,N_19305);
and UO_106 (O_106,N_18879,N_19059);
nand UO_107 (O_107,N_17657,N_17242);
or UO_108 (O_108,N_16448,N_17742);
nor UO_109 (O_109,N_17217,N_18304);
or UO_110 (O_110,N_18009,N_17783);
nand UO_111 (O_111,N_17064,N_17853);
and UO_112 (O_112,N_19906,N_18692);
and UO_113 (O_113,N_16772,N_19088);
nor UO_114 (O_114,N_18432,N_19837);
and UO_115 (O_115,N_19794,N_17529);
nor UO_116 (O_116,N_17974,N_18678);
or UO_117 (O_117,N_16470,N_17847);
and UO_118 (O_118,N_16745,N_16222);
nand UO_119 (O_119,N_18069,N_16131);
nor UO_120 (O_120,N_16610,N_17265);
and UO_121 (O_121,N_18590,N_19832);
or UO_122 (O_122,N_16039,N_19228);
nand UO_123 (O_123,N_16197,N_17161);
or UO_124 (O_124,N_19346,N_16345);
nor UO_125 (O_125,N_17936,N_18695);
nand UO_126 (O_126,N_19040,N_19187);
and UO_127 (O_127,N_17269,N_17132);
xnor UO_128 (O_128,N_16433,N_17755);
nand UO_129 (O_129,N_19690,N_17230);
nand UO_130 (O_130,N_19201,N_17363);
and UO_131 (O_131,N_18733,N_16898);
nand UO_132 (O_132,N_17778,N_17556);
and UO_133 (O_133,N_16163,N_19405);
or UO_134 (O_134,N_19316,N_17210);
or UO_135 (O_135,N_19273,N_19401);
and UO_136 (O_136,N_16976,N_17768);
and UO_137 (O_137,N_16155,N_16319);
and UO_138 (O_138,N_18180,N_18276);
or UO_139 (O_139,N_17357,N_16323);
or UO_140 (O_140,N_19809,N_16028);
nor UO_141 (O_141,N_16481,N_18413);
and UO_142 (O_142,N_19575,N_17261);
nand UO_143 (O_143,N_16682,N_19803);
nor UO_144 (O_144,N_17218,N_17972);
or UO_145 (O_145,N_16093,N_18836);
nand UO_146 (O_146,N_16938,N_18151);
xnor UO_147 (O_147,N_19067,N_16903);
and UO_148 (O_148,N_18431,N_18513);
nor UO_149 (O_149,N_17978,N_19311);
nand UO_150 (O_150,N_18681,N_16736);
or UO_151 (O_151,N_18938,N_18182);
and UO_152 (O_152,N_17807,N_17677);
or UO_153 (O_153,N_19131,N_18929);
and UO_154 (O_154,N_18857,N_16452);
or UO_155 (O_155,N_19982,N_18738);
or UO_156 (O_156,N_16187,N_17549);
xor UO_157 (O_157,N_16383,N_19628);
or UO_158 (O_158,N_16656,N_16825);
and UO_159 (O_159,N_19070,N_18330);
nor UO_160 (O_160,N_16298,N_19119);
nor UO_161 (O_161,N_16074,N_16089);
and UO_162 (O_162,N_18603,N_18035);
nand UO_163 (O_163,N_17307,N_16820);
nor UO_164 (O_164,N_18920,N_16365);
xor UO_165 (O_165,N_19288,N_19955);
nand UO_166 (O_166,N_19846,N_19890);
nand UO_167 (O_167,N_16344,N_16387);
and UO_168 (O_168,N_16786,N_17181);
and UO_169 (O_169,N_16162,N_16106);
nor UO_170 (O_170,N_18280,N_17128);
and UO_171 (O_171,N_19104,N_19604);
nand UO_172 (O_172,N_18694,N_19647);
and UO_173 (O_173,N_19750,N_16715);
or UO_174 (O_174,N_16125,N_19961);
xor UO_175 (O_175,N_19940,N_18293);
nor UO_176 (O_176,N_19709,N_18988);
nand UO_177 (O_177,N_18242,N_17080);
nor UO_178 (O_178,N_17390,N_17444);
and UO_179 (O_179,N_19214,N_19215);
nand UO_180 (O_180,N_18436,N_16116);
nand UO_181 (O_181,N_18865,N_18766);
nand UO_182 (O_182,N_19402,N_18179);
nor UO_183 (O_183,N_19635,N_17365);
nand UO_184 (O_184,N_17037,N_16998);
and UO_185 (O_185,N_16516,N_18561);
nand UO_186 (O_186,N_17087,N_19748);
and UO_187 (O_187,N_16814,N_18341);
or UO_188 (O_188,N_16505,N_19182);
xnor UO_189 (O_189,N_18479,N_18369);
or UO_190 (O_190,N_19160,N_19544);
nor UO_191 (O_191,N_17483,N_18127);
nand UO_192 (O_192,N_16571,N_19893);
nand UO_193 (O_193,N_16047,N_18624);
or UO_194 (O_194,N_18120,N_17739);
or UO_195 (O_195,N_19390,N_17457);
nand UO_196 (O_196,N_19774,N_18187);
and UO_197 (O_197,N_18290,N_17885);
and UO_198 (O_198,N_18441,N_16301);
or UO_199 (O_199,N_17888,N_18043);
or UO_200 (O_200,N_18523,N_17107);
and UO_201 (O_201,N_17477,N_19609);
and UO_202 (O_202,N_16952,N_16062);
nand UO_203 (O_203,N_19195,N_16774);
nor UO_204 (O_204,N_19287,N_18456);
and UO_205 (O_205,N_16221,N_19330);
xor UO_206 (O_206,N_17103,N_19693);
nor UO_207 (O_207,N_19734,N_18852);
or UO_208 (O_208,N_17428,N_17117);
nor UO_209 (O_209,N_17889,N_16243);
nor UO_210 (O_210,N_16010,N_18223);
or UO_211 (O_211,N_16455,N_18707);
or UO_212 (O_212,N_16209,N_19652);
and UO_213 (O_213,N_19474,N_18206);
and UO_214 (O_214,N_18908,N_19644);
or UO_215 (O_215,N_16398,N_17131);
nand UO_216 (O_216,N_17851,N_19134);
nand UO_217 (O_217,N_19226,N_16502);
and UO_218 (O_218,N_18993,N_19520);
nor UO_219 (O_219,N_16286,N_16145);
nand UO_220 (O_220,N_18937,N_17472);
nor UO_221 (O_221,N_19356,N_16204);
and UO_222 (O_222,N_17661,N_17196);
xnor UO_223 (O_223,N_16400,N_18734);
nor UO_224 (O_224,N_17869,N_19199);
and UO_225 (O_225,N_18121,N_19241);
and UO_226 (O_226,N_19801,N_19995);
or UO_227 (O_227,N_17126,N_17570);
nand UO_228 (O_228,N_19101,N_19720);
xor UO_229 (O_229,N_16226,N_19333);
nand UO_230 (O_230,N_18829,N_17038);
or UO_231 (O_231,N_18401,N_18430);
nand UO_232 (O_232,N_17278,N_17756);
nand UO_233 (O_233,N_18022,N_18787);
and UO_234 (O_234,N_18637,N_18794);
or UO_235 (O_235,N_19827,N_17697);
xnor UO_236 (O_236,N_17152,N_17744);
or UO_237 (O_237,N_18181,N_18859);
nor UO_238 (O_238,N_18711,N_18263);
nor UO_239 (O_239,N_19547,N_16979);
xor UO_240 (O_240,N_16646,N_17527);
xnor UO_241 (O_241,N_16064,N_16850);
nor UO_242 (O_242,N_18797,N_16835);
or UO_243 (O_243,N_18289,N_17500);
and UO_244 (O_244,N_19063,N_19825);
or UO_245 (O_245,N_19976,N_18241);
nor UO_246 (O_246,N_16325,N_18054);
or UO_247 (O_247,N_18914,N_16025);
nor UO_248 (O_248,N_16208,N_18571);
nor UO_249 (O_249,N_18537,N_18435);
nand UO_250 (O_250,N_17671,N_19886);
and UO_251 (O_251,N_18439,N_16274);
nand UO_252 (O_252,N_19624,N_17710);
and UO_253 (O_253,N_16154,N_19555);
nand UO_254 (O_254,N_17252,N_17414);
xnor UO_255 (O_255,N_18373,N_19643);
nor UO_256 (O_256,N_19558,N_18191);
nand UO_257 (O_257,N_17380,N_18335);
and UO_258 (O_258,N_18005,N_18301);
or UO_259 (O_259,N_19428,N_17384);
nor UO_260 (O_260,N_19735,N_19417);
or UO_261 (O_261,N_17120,N_16021);
and UO_262 (O_262,N_17068,N_16941);
xor UO_263 (O_263,N_19408,N_16186);
nor UO_264 (O_264,N_19130,N_18531);
nand UO_265 (O_265,N_17860,N_17272);
or UO_266 (O_266,N_17001,N_17029);
xnor UO_267 (O_267,N_17011,N_17163);
and UO_268 (O_268,N_18504,N_19171);
nor UO_269 (O_269,N_17993,N_18783);
and UO_270 (O_270,N_19004,N_19991);
or UO_271 (O_271,N_19458,N_16716);
and UO_272 (O_272,N_19570,N_16273);
nor UO_273 (O_273,N_16024,N_16635);
nand UO_274 (O_274,N_18606,N_19595);
nand UO_275 (O_275,N_18862,N_17224);
and UO_276 (O_276,N_18382,N_17938);
nor UO_277 (O_277,N_18404,N_16633);
or UO_278 (O_278,N_16069,N_16032);
nor UO_279 (O_279,N_19194,N_16218);
nand UO_280 (O_280,N_19106,N_19948);
nor UO_281 (O_281,N_18093,N_18460);
and UO_282 (O_282,N_16411,N_19954);
nor UO_283 (O_283,N_19178,N_17017);
xnor UO_284 (O_284,N_18587,N_19260);
and UO_285 (O_285,N_18583,N_19329);
xnor UO_286 (O_286,N_17931,N_17031);
or UO_287 (O_287,N_16929,N_16622);
and UO_288 (O_288,N_18721,N_17540);
nand UO_289 (O_289,N_18553,N_17244);
or UO_290 (O_290,N_19551,N_18500);
nor UO_291 (O_291,N_19706,N_18362);
and UO_292 (O_292,N_18586,N_17360);
nor UO_293 (O_293,N_17965,N_18024);
or UO_294 (O_294,N_16351,N_17874);
nor UO_295 (O_295,N_16620,N_17738);
nand UO_296 (O_296,N_19248,N_19303);
nand UO_297 (O_297,N_18782,N_17354);
nor UO_298 (O_298,N_16629,N_17944);
nand UO_299 (O_299,N_19023,N_16581);
nand UO_300 (O_300,N_19035,N_19237);
and UO_301 (O_301,N_19623,N_18878);
or UO_302 (O_302,N_19760,N_19648);
nor UO_303 (O_303,N_18639,N_17784);
or UO_304 (O_304,N_19871,N_16504);
nand UO_305 (O_305,N_17822,N_19905);
nor UO_306 (O_306,N_16055,N_16198);
and UO_307 (O_307,N_18853,N_16738);
nor UO_308 (O_308,N_19675,N_16598);
or UO_309 (O_309,N_16991,N_17986);
xnor UO_310 (O_310,N_19470,N_17425);
nand UO_311 (O_311,N_19580,N_17464);
nor UO_312 (O_312,N_18851,N_18913);
xnor UO_313 (O_313,N_16532,N_18450);
and UO_314 (O_314,N_16216,N_17649);
or UO_315 (O_315,N_16844,N_18636);
or UO_316 (O_316,N_19883,N_17624);
and UO_317 (O_317,N_17495,N_18912);
nor UO_318 (O_318,N_16382,N_19859);
nand UO_319 (O_319,N_17857,N_19382);
nand UO_320 (O_320,N_16830,N_16246);
xnor UO_321 (O_321,N_16692,N_19454);
nand UO_322 (O_322,N_16680,N_18243);
nor UO_323 (O_323,N_17338,N_16368);
xnor UO_324 (O_324,N_17769,N_19862);
nand UO_325 (O_325,N_16966,N_16171);
nor UO_326 (O_326,N_16776,N_19348);
nand UO_327 (O_327,N_17182,N_19054);
and UO_328 (O_328,N_16659,N_17115);
or UO_329 (O_329,N_16220,N_18778);
or UO_330 (O_330,N_17321,N_18390);
xnor UO_331 (O_331,N_18148,N_16939);
xor UO_332 (O_332,N_17348,N_17678);
or UO_333 (O_333,N_17485,N_17648);
and UO_334 (O_334,N_17423,N_16217);
nand UO_335 (O_335,N_18960,N_17610);
and UO_336 (O_336,N_19980,N_16493);
nand UO_337 (O_337,N_16780,N_18056);
and UO_338 (O_338,N_19399,N_16657);
and UO_339 (O_339,N_19534,N_18484);
or UO_340 (O_340,N_16613,N_18600);
nor UO_341 (O_341,N_17083,N_18229);
nand UO_342 (O_342,N_17059,N_19005);
and UO_343 (O_343,N_17019,N_17452);
nor UO_344 (O_344,N_19581,N_19150);
and UO_345 (O_345,N_19268,N_18900);
and UO_346 (O_346,N_17534,N_18663);
or UO_347 (O_347,N_18086,N_18454);
nor UO_348 (O_348,N_18059,N_18389);
nor UO_349 (O_349,N_17979,N_17988);
nor UO_350 (O_350,N_18233,N_16636);
xor UO_351 (O_351,N_17735,N_19501);
or UO_352 (O_352,N_18532,N_16135);
nor UO_353 (O_353,N_18732,N_16339);
nand UO_354 (O_354,N_19562,N_19727);
nand UO_355 (O_355,N_17046,N_17194);
or UO_356 (O_356,N_16153,N_19203);
or UO_357 (O_357,N_19996,N_18727);
and UO_358 (O_358,N_19253,N_17295);
nand UO_359 (O_359,N_17111,N_18102);
xor UO_360 (O_360,N_18795,N_16841);
nor UO_361 (O_361,N_16192,N_18252);
nor UO_362 (O_362,N_18495,N_18100);
and UO_363 (O_363,N_16963,N_16641);
nor UO_364 (O_364,N_16707,N_18512);
nand UO_365 (O_365,N_18141,N_16630);
or UO_366 (O_366,N_18568,N_19525);
xor UO_367 (O_367,N_17582,N_16108);
nor UO_368 (O_368,N_18811,N_16290);
or UO_369 (O_369,N_17670,N_16441);
nor UO_370 (O_370,N_17937,N_16360);
nor UO_371 (O_371,N_17439,N_18786);
or UO_372 (O_372,N_19561,N_16372);
and UO_373 (O_373,N_19415,N_19079);
or UO_374 (O_374,N_17257,N_17034);
nand UO_375 (O_375,N_17958,N_16310);
nand UO_376 (O_376,N_18492,N_18403);
and UO_377 (O_377,N_16887,N_18832);
nor UO_378 (O_378,N_16052,N_18816);
nor UO_379 (O_379,N_16847,N_18378);
and UO_380 (O_380,N_18932,N_16619);
and UO_381 (O_381,N_17039,N_17559);
or UO_382 (O_382,N_19563,N_18273);
or UO_383 (O_383,N_18625,N_19489);
nand UO_384 (O_384,N_19385,N_18333);
or UO_385 (O_385,N_17154,N_18933);
nand UO_386 (O_386,N_18701,N_18393);
nand UO_387 (O_387,N_16922,N_19042);
nor UO_388 (O_388,N_16279,N_18463);
and UO_389 (O_389,N_18798,N_18458);
or UO_390 (O_390,N_19753,N_19453);
nor UO_391 (O_391,N_16726,N_18138);
or UO_392 (O_392,N_16765,N_19338);
and UO_393 (O_393,N_16671,N_16110);
and UO_394 (O_394,N_19238,N_19398);
xor UO_395 (O_395,N_16326,N_18567);
and UO_396 (O_396,N_16842,N_17247);
nand UO_397 (O_397,N_17419,N_16698);
nor UO_398 (O_398,N_19321,N_16320);
and UO_399 (O_399,N_17852,N_19684);
nor UO_400 (O_400,N_18291,N_16937);
nor UO_401 (O_401,N_19921,N_18124);
and UO_402 (O_402,N_18380,N_18286);
or UO_403 (O_403,N_17222,N_17854);
nand UO_404 (O_404,N_17725,N_19758);
and UO_405 (O_405,N_19782,N_19866);
xnor UO_406 (O_406,N_19020,N_17947);
and UO_407 (O_407,N_18808,N_19899);
and UO_408 (O_408,N_19127,N_19358);
and UO_409 (O_409,N_17129,N_16067);
nand UO_410 (O_410,N_18780,N_17943);
or UO_411 (O_411,N_17201,N_19936);
nor UO_412 (O_412,N_16138,N_18945);
nand UO_413 (O_413,N_16527,N_16943);
or UO_414 (O_414,N_17764,N_16267);
nand UO_415 (O_415,N_17466,N_16495);
nor UO_416 (O_416,N_19464,N_19442);
xor UO_417 (O_417,N_16119,N_16792);
xnor UO_418 (O_418,N_18855,N_18643);
nand UO_419 (O_419,N_19923,N_17656);
nor UO_420 (O_420,N_18877,N_18521);
or UO_421 (O_421,N_17311,N_19556);
nand UO_422 (O_422,N_19002,N_19989);
and UO_423 (O_423,N_18079,N_16115);
nor UO_424 (O_424,N_19424,N_18381);
nand UO_425 (O_425,N_17082,N_18983);
nand UO_426 (O_426,N_17929,N_19451);
nor UO_427 (O_427,N_18046,N_19632);
nand UO_428 (O_428,N_18641,N_17589);
or UO_429 (O_429,N_19186,N_19788);
and UO_430 (O_430,N_19538,N_19157);
nand UO_431 (O_431,N_18208,N_16925);
or UO_432 (O_432,N_19739,N_19950);
xor UO_433 (O_433,N_19468,N_19509);
nand UO_434 (O_434,N_17253,N_18088);
and UO_435 (O_435,N_16562,N_19816);
nand UO_436 (O_436,N_16755,N_18962);
and UO_437 (O_437,N_18743,N_17192);
nor UO_438 (O_438,N_17282,N_19297);
nor UO_439 (O_439,N_16027,N_19614);
xor UO_440 (O_440,N_17303,N_17199);
nor UO_441 (O_441,N_16843,N_16928);
nand UO_442 (O_442,N_17248,N_17625);
nand UO_443 (O_443,N_16098,N_16017);
xnor UO_444 (O_444,N_18530,N_19123);
nor UO_445 (O_445,N_18055,N_16317);
or UO_446 (O_446,N_16670,N_17366);
or UO_447 (O_447,N_18310,N_19941);
and UO_448 (O_448,N_18582,N_17081);
nor UO_449 (O_449,N_17185,N_19650);
nor UO_450 (O_450,N_17319,N_16330);
and UO_451 (O_451,N_17896,N_17268);
nor UO_452 (O_452,N_19137,N_18105);
nand UO_453 (O_453,N_19713,N_17051);
nand UO_454 (O_454,N_19554,N_16181);
nand UO_455 (O_455,N_19669,N_17007);
nand UO_456 (O_456,N_18515,N_18619);
xor UO_457 (O_457,N_18628,N_17198);
nand UO_458 (O_458,N_16761,N_19599);
nor UO_459 (O_459,N_19550,N_17881);
nand UO_460 (O_460,N_17086,N_17290);
and UO_461 (O_461,N_19642,N_17484);
nor UO_462 (O_462,N_18464,N_18957);
xor UO_463 (O_463,N_16088,N_19662);
nor UO_464 (O_464,N_18528,N_17963);
nor UO_465 (O_465,N_17171,N_19685);
nand UO_466 (O_466,N_16916,N_18031);
nand UO_467 (O_467,N_16833,N_17759);
and UO_468 (O_468,N_19061,N_17167);
nand UO_469 (O_469,N_19045,N_17442);
nand UO_470 (O_470,N_18405,N_16587);
and UO_471 (O_471,N_19416,N_17585);
nor UO_472 (O_472,N_19970,N_18438);
nand UO_473 (O_473,N_18061,N_18419);
and UO_474 (O_474,N_16769,N_17371);
and UO_475 (O_475,N_16696,N_19990);
or UO_476 (O_476,N_18387,N_17151);
nor UO_477 (O_477,N_19053,N_17124);
nand UO_478 (O_478,N_16229,N_16540);
or UO_479 (O_479,N_19603,N_16490);
and UO_480 (O_480,N_16764,N_16611);
or UO_481 (O_481,N_16195,N_18248);
and UO_482 (O_482,N_16424,N_19164);
nand UO_483 (O_483,N_16975,N_19496);
nor UO_484 (O_484,N_18239,N_17026);
and UO_485 (O_485,N_17099,N_18731);
nor UO_486 (O_486,N_16808,N_19136);
xor UO_487 (O_487,N_18475,N_17286);
nand UO_488 (O_488,N_17373,N_16356);
nor UO_489 (O_489,N_19155,N_18095);
nor UO_490 (O_490,N_17309,N_19209);
and UO_491 (O_491,N_18224,N_18128);
or UO_492 (O_492,N_16404,N_18339);
nand UO_493 (O_493,N_17239,N_18397);
nor UO_494 (O_494,N_19027,N_18134);
nor UO_495 (O_495,N_18491,N_18771);
or UO_496 (O_496,N_17962,N_16589);
xor UO_497 (O_497,N_16775,N_19557);
and UO_498 (O_498,N_17310,N_19360);
and UO_499 (O_499,N_17855,N_18259);
or UO_500 (O_500,N_19666,N_19267);
nand UO_501 (O_501,N_16134,N_19780);
nand UO_502 (O_502,N_16787,N_16340);
or UO_503 (O_503,N_16911,N_18842);
xnor UO_504 (O_504,N_19357,N_16564);
nor UO_505 (O_505,N_16308,N_19870);
and UO_506 (O_506,N_16234,N_17004);
and UO_507 (O_507,N_19000,N_18931);
and UO_508 (O_508,N_16281,N_18010);
nand UO_509 (O_509,N_19994,N_16623);
and UO_510 (O_510,N_17119,N_18892);
and UO_511 (O_511,N_17208,N_17950);
nand UO_512 (O_512,N_16227,N_19672);
nand UO_513 (O_513,N_18592,N_17873);
and UO_514 (O_514,N_16704,N_18219);
nor UO_515 (O_515,N_17219,N_17564);
nor UO_516 (O_516,N_19731,N_16260);
nand UO_517 (O_517,N_16268,N_17283);
or UO_518 (O_518,N_18347,N_17596);
and UO_519 (O_519,N_19569,N_16838);
and UO_520 (O_520,N_19011,N_17815);
or UO_521 (O_521,N_18514,N_18887);
and UO_522 (O_522,N_19698,N_17005);
nand UO_523 (O_523,N_18476,N_18621);
nand UO_524 (O_524,N_19472,N_17153);
and UO_525 (O_525,N_16853,N_16215);
xor UO_526 (O_526,N_17737,N_18411);
and UO_527 (O_527,N_19688,N_18420);
and UO_528 (O_528,N_18220,N_16997);
nand UO_529 (O_529,N_18546,N_17177);
nand UO_530 (O_530,N_17511,N_18225);
or UO_531 (O_531,N_18412,N_19847);
or UO_532 (O_532,N_19191,N_16276);
and UO_533 (O_533,N_17623,N_17398);
or UO_534 (O_534,N_19121,N_19469);
or UO_535 (O_535,N_19630,N_19937);
nand UO_536 (O_536,N_17227,N_19953);
nor UO_537 (O_537,N_17651,N_17665);
nand UO_538 (O_538,N_19740,N_19776);
and UO_539 (O_539,N_19174,N_18710);
or UO_540 (O_540,N_19649,N_19345);
and UO_541 (O_541,N_18116,N_17445);
xnor UO_542 (O_542,N_18904,N_19711);
or UO_543 (O_543,N_17687,N_19262);
nor UO_544 (O_544,N_17804,N_18399);
and UO_545 (O_545,N_16640,N_16166);
and UO_546 (O_546,N_18823,N_16759);
or UO_547 (O_547,N_17329,N_17280);
nand UO_548 (O_548,N_17003,N_19340);
nand UO_549 (O_549,N_18007,N_18357);
nor UO_550 (O_550,N_19519,N_17780);
nand UO_551 (O_551,N_17886,N_18204);
nand UO_552 (O_552,N_19466,N_17597);
nor UO_553 (O_553,N_18049,N_16284);
nor UO_554 (O_554,N_19773,N_19754);
and UO_555 (O_555,N_18104,N_16910);
xor UO_556 (O_556,N_17834,N_17264);
or UO_557 (O_557,N_17186,N_16851);
nand UO_558 (O_558,N_16013,N_17925);
nand UO_559 (O_559,N_19456,N_19185);
nand UO_560 (O_560,N_16124,N_16491);
nor UO_561 (O_561,N_19729,N_18089);
or UO_562 (O_562,N_16520,N_17394);
and UO_563 (O_563,N_17959,N_19352);
and UO_564 (O_564,N_18720,N_17109);
xnor UO_565 (O_565,N_19149,N_16120);
nand UO_566 (O_566,N_16019,N_17516);
nand UO_567 (O_567,N_19473,N_16560);
nand UO_568 (O_568,N_19527,N_17376);
or UO_569 (O_569,N_16791,N_19014);
nor UO_570 (O_570,N_18557,N_18323);
or UO_571 (O_571,N_17826,N_19804);
or UO_572 (O_572,N_18246,N_19087);
and UO_573 (O_573,N_16476,N_17492);
nor UO_574 (O_574,N_16626,N_18254);
and UO_575 (O_575,N_18416,N_18640);
or UO_576 (O_576,N_19007,N_16645);
or UO_577 (O_577,N_19486,N_17251);
or UO_578 (O_578,N_19574,N_17116);
nor UO_579 (O_579,N_16129,N_17043);
and UO_580 (O_580,N_16877,N_16492);
nor UO_581 (O_581,N_17320,N_17720);
nand UO_582 (O_582,N_17928,N_18200);
nor UO_583 (O_583,N_17062,N_16824);
or UO_584 (O_584,N_18066,N_17734);
nand UO_585 (O_585,N_17463,N_17254);
or UO_586 (O_586,N_17557,N_17814);
xnor UO_587 (O_587,N_19440,N_19335);
nor UO_588 (O_588,N_18807,N_16957);
nor UO_589 (O_589,N_18833,N_19167);
nor UO_590 (O_590,N_18870,N_19860);
or UO_591 (O_591,N_16416,N_18542);
nor UO_592 (O_592,N_19768,N_18300);
or UO_593 (O_593,N_16354,N_17061);
or UO_594 (O_594,N_16978,N_16812);
nor UO_595 (O_595,N_17799,N_16029);
or UO_596 (O_596,N_19497,N_19141);
nand UO_597 (O_597,N_19103,N_16909);
and UO_598 (O_598,N_19144,N_17825);
or UO_599 (O_599,N_18968,N_18063);
and UO_600 (O_600,N_18257,N_17076);
or UO_601 (O_601,N_18230,N_16758);
nand UO_602 (O_602,N_16603,N_17574);
nand UO_603 (O_603,N_17277,N_17953);
xor UO_604 (O_604,N_19901,N_17545);
nor UO_605 (O_605,N_18605,N_16060);
or UO_606 (O_606,N_18735,N_18402);
nand UO_607 (O_607,N_16384,N_17141);
or UO_608 (O_608,N_16297,N_17907);
and UO_609 (O_609,N_16926,N_18652);
nor UO_610 (O_610,N_18424,N_16888);
and UO_611 (O_611,N_17718,N_18110);
nor UO_612 (O_612,N_16519,N_16172);
and UO_613 (O_613,N_16303,N_18038);
nor UO_614 (O_614,N_18856,N_18171);
nand UO_615 (O_615,N_17933,N_18919);
nand UO_616 (O_616,N_19095,N_18924);
and UO_617 (O_617,N_19500,N_19151);
nand UO_618 (O_618,N_16590,N_19168);
or UO_619 (O_619,N_17147,N_17349);
and UO_620 (O_620,N_19665,N_19105);
or UO_621 (O_621,N_19573,N_19064);
or UO_622 (O_622,N_18996,N_17985);
nand UO_623 (O_623,N_17100,N_18367);
nor UO_624 (O_624,N_16582,N_19397);
and UO_625 (O_625,N_18410,N_18918);
nor UO_626 (O_626,N_17220,N_18944);
xnor UO_627 (O_627,N_16395,N_16484);
nand UO_628 (O_628,N_18576,N_16214);
xor UO_629 (O_629,N_19505,N_19312);
or UO_630 (O_630,N_18068,N_16725);
xor UO_631 (O_631,N_16695,N_18361);
nand UO_632 (O_632,N_19183,N_18327);
nor UO_633 (O_633,N_18334,N_16350);
and UO_634 (O_634,N_19410,N_17588);
nand UO_635 (O_635,N_19560,N_17226);
nand UO_636 (O_636,N_19882,N_16760);
or UO_637 (O_637,N_17956,N_17041);
nor UO_638 (O_638,N_18655,N_19047);
nor UO_639 (O_639,N_17843,N_18213);
and UO_640 (O_640,N_16004,N_17358);
or UO_641 (O_641,N_19579,N_19213);
nand UO_642 (O_642,N_18658,N_19484);
or UO_643 (O_643,N_17638,N_16709);
nor UO_644 (O_644,N_19487,N_19043);
nor UO_645 (O_645,N_16016,N_18839);
nor UO_646 (O_646,N_19792,N_17650);
or UO_647 (O_647,N_16643,N_19715);
or UO_648 (O_648,N_17714,N_18490);
or UO_649 (O_649,N_18489,N_16454);
nand UO_650 (O_650,N_19523,N_17707);
and UO_651 (O_651,N_16907,N_18299);
xor UO_652 (O_652,N_19098,N_16434);
and UO_653 (O_653,N_19717,N_17123);
and UO_654 (O_654,N_18999,N_18076);
xor UO_655 (O_655,N_18326,N_17023);
and UO_656 (O_656,N_17315,N_18363);
nor UO_657 (O_657,N_19283,N_17571);
or UO_658 (O_658,N_18130,N_19317);
and UO_659 (O_659,N_19975,N_16152);
nor UO_660 (O_660,N_17146,N_16628);
nor UO_661 (O_661,N_17058,N_16509);
and UO_662 (O_662,N_19752,N_17203);
and UO_663 (O_663,N_17008,N_18973);
and UO_664 (O_664,N_17158,N_18751);
nand UO_665 (O_665,N_18483,N_19716);
nand UO_666 (O_666,N_16936,N_17518);
nor UO_667 (O_667,N_19694,N_16701);
and UO_668 (O_668,N_16377,N_16415);
nand UO_669 (O_669,N_16348,N_16684);
and UO_670 (O_670,N_17808,N_16256);
nand UO_671 (O_671,N_16955,N_17654);
nor UO_672 (O_672,N_16555,N_17427);
or UO_673 (O_673,N_16456,N_16806);
nor UO_674 (O_674,N_18616,N_19657);
or UO_675 (O_675,N_19799,N_18040);
xor UO_676 (O_676,N_17334,N_17327);
or UO_677 (O_677,N_16444,N_17413);
nor UO_678 (O_678,N_18951,N_18077);
nor UO_679 (O_679,N_17343,N_19420);
or UO_680 (O_680,N_16457,N_19691);
or UO_681 (O_681,N_16231,N_18969);
or UO_682 (O_682,N_16193,N_16225);
nor UO_683 (O_683,N_17350,N_17054);
xor UO_684 (O_684,N_19227,N_18867);
and UO_685 (O_685,N_16447,N_18469);
and UO_686 (O_686,N_16228,N_18013);
nor UO_687 (O_687,N_19277,N_19915);
and UO_688 (O_688,N_19537,N_19077);
or UO_689 (O_689,N_18418,N_17999);
and UO_690 (O_690,N_18757,N_18015);
nor UO_691 (O_691,N_19206,N_18471);
or UO_692 (O_692,N_17359,N_17798);
or UO_693 (O_693,N_17102,N_17903);
and UO_694 (O_694,N_16465,N_17724);
nor UO_695 (O_695,N_18264,N_19229);
nor UO_696 (O_696,N_16427,N_16513);
or UO_697 (O_697,N_18758,N_17235);
or UO_698 (O_698,N_19835,N_18664);
nand UO_699 (O_699,N_17089,N_17871);
nand UO_700 (O_700,N_16046,N_16983);
and UO_701 (O_701,N_19586,N_16041);
nor UO_702 (O_702,N_16794,N_19738);
and UO_703 (O_703,N_19597,N_16521);
or UO_704 (O_704,N_16700,N_19910);
or UO_705 (O_705,N_17992,N_17716);
nand UO_706 (O_706,N_19842,N_18221);
xnor UO_707 (O_707,N_18162,N_16307);
or UO_708 (O_708,N_16065,N_16466);
or UO_709 (O_709,N_16159,N_18173);
xnor UO_710 (O_710,N_17276,N_18365);
and UO_711 (O_711,N_18374,N_18584);
and UO_712 (O_712,N_17353,N_18793);
and UO_713 (O_713,N_17794,N_18910);
or UO_714 (O_714,N_16574,N_19831);
or UO_715 (O_715,N_16935,N_19972);
nor UO_716 (O_716,N_17892,N_19607);
and UO_717 (O_717,N_16994,N_17468);
and UO_718 (O_718,N_19359,N_18342);
and UO_719 (O_719,N_16547,N_16813);
or UO_720 (O_720,N_18085,N_19962);
xor UO_721 (O_721,N_16366,N_18814);
xnor UO_722 (O_722,N_19510,N_18356);
and UO_723 (O_723,N_18895,N_19166);
nor UO_724 (O_724,N_19377,N_18002);
and UO_725 (O_725,N_18610,N_17395);
and UO_726 (O_726,N_19240,N_19018);
nor UO_727 (O_727,N_18360,N_18745);
xor UO_728 (O_728,N_19224,N_19001);
and UO_729 (O_729,N_18891,N_16313);
nand UO_730 (O_730,N_16799,N_18279);
and UO_731 (O_731,N_16327,N_18099);
nor UO_732 (O_732,N_18319,N_18133);
nor UO_733 (O_733,N_16886,N_18661);
and UO_734 (O_734,N_19755,N_18526);
or UO_735 (O_735,N_17281,N_18421);
or UO_736 (O_736,N_17454,N_19412);
xnor UO_737 (O_737,N_16182,N_19111);
or UO_738 (O_738,N_19969,N_17809);
nand UO_739 (O_739,N_16528,N_19848);
and UO_740 (O_740,N_19834,N_17531);
and UO_741 (O_741,N_19289,N_19865);
nor UO_742 (O_742,N_19022,N_16439);
nor UO_743 (O_743,N_18942,N_16538);
nand UO_744 (O_744,N_19880,N_17162);
nand UO_745 (O_745,N_19394,N_17487);
nand UO_746 (O_746,N_19177,N_18529);
nor UO_747 (O_747,N_17053,N_17063);
nand UO_748 (O_748,N_17344,N_16508);
or UO_749 (O_749,N_19493,N_18211);
and UO_750 (O_750,N_19060,N_19565);
or UO_751 (O_751,N_18271,N_19764);
and UO_752 (O_752,N_18524,N_17471);
nor UO_753 (O_753,N_16654,N_17779);
or UO_754 (O_754,N_18792,N_16045);
xnor UO_755 (O_755,N_16379,N_16821);
nor UO_756 (O_756,N_19812,N_19110);
or UO_757 (O_757,N_18218,N_17682);
nor UO_758 (O_758,N_17844,N_19710);
nor UO_759 (O_759,N_17312,N_17749);
xor UO_760 (O_760,N_17601,N_19304);
and UO_761 (O_761,N_18313,N_17954);
xnor UO_762 (O_762,N_17474,N_18984);
or UO_763 (O_763,N_16438,N_19894);
and UO_764 (O_764,N_17998,N_17690);
and UO_765 (O_765,N_18296,N_18118);
nor UO_766 (O_766,N_19967,N_18719);
nand UO_767 (O_767,N_17347,N_19678);
or UO_768 (O_768,N_17482,N_19266);
nor UO_769 (O_769,N_16146,N_17562);
nand UO_770 (O_770,N_17681,N_19908);
xor UO_771 (O_771,N_17407,N_16693);
xor UO_772 (O_772,N_19598,N_19483);
or UO_773 (O_773,N_19122,N_16477);
and UO_774 (O_774,N_19353,N_19270);
or UO_775 (O_775,N_17607,N_17968);
and UO_776 (O_776,N_18725,N_17298);
nand UO_777 (O_777,N_19726,N_18667);
and UO_778 (O_778,N_16189,N_19987);
nand UO_779 (O_779,N_16987,N_17961);
nor UO_780 (O_780,N_17891,N_19478);
nor UO_781 (O_781,N_17872,N_19172);
or UO_782 (O_782,N_19285,N_18470);
nand UO_783 (O_783,N_17662,N_16891);
nor UO_784 (O_784,N_19366,N_16094);
nor UO_785 (O_785,N_19236,N_19524);
and UO_786 (O_786,N_16239,N_17836);
nand UO_787 (O_787,N_16099,N_16717);
nor UO_788 (O_788,N_18712,N_16778);
or UO_789 (O_789,N_17355,N_16127);
nand UO_790 (O_790,N_16752,N_19993);
nor UO_791 (O_791,N_18803,N_17050);
xnor UO_792 (O_792,N_19467,N_18212);
nor UO_793 (O_793,N_19230,N_18275);
and UO_794 (O_794,N_18425,N_18372);
nand UO_795 (O_795,N_19450,N_17595);
xnor UO_796 (O_796,N_18001,N_18650);
xnor UO_797 (O_797,N_18657,N_18087);
and UO_798 (O_798,N_19771,N_18270);
and UO_799 (O_799,N_18287,N_16259);
and UO_800 (O_800,N_18684,N_16449);
or UO_801 (O_801,N_16376,N_19152);
nand UO_802 (O_802,N_18083,N_18488);
nand UO_803 (O_803,N_17326,N_19539);
nand UO_804 (O_804,N_19935,N_17494);
or UO_805 (O_805,N_18776,N_18872);
and UO_806 (O_806,N_16753,N_18144);
and UO_807 (O_807,N_19261,N_19073);
and UO_808 (O_808,N_17684,N_16270);
or UO_809 (O_809,N_17434,N_19637);
nand UO_810 (O_810,N_16254,N_19438);
and UO_811 (O_811,N_17818,N_17489);
and UO_812 (O_812,N_19143,N_19572);
nor UO_813 (O_813,N_19888,N_18699);
and UO_814 (O_814,N_16422,N_17713);
nor UO_815 (O_815,N_17459,N_18169);
nor UO_816 (O_816,N_18481,N_18343);
nand UO_817 (O_817,N_19142,N_19037);
nand UO_818 (O_818,N_18377,N_18680);
nor UO_819 (O_819,N_18979,N_16757);
nor UO_820 (O_820,N_18741,N_18216);
xor UO_821 (O_821,N_16185,N_17021);
nand UO_822 (O_822,N_18107,N_19999);
and UO_823 (O_823,N_16510,N_17473);
nand UO_824 (O_824,N_19084,N_17386);
or UO_825 (O_825,N_18395,N_16867);
and UO_826 (O_826,N_17612,N_16158);
and UO_827 (O_827,N_16906,N_17498);
nor UO_828 (O_828,N_19730,N_17479);
nand UO_829 (O_829,N_18366,N_19234);
nand UO_830 (O_830,N_17300,N_17461);
nor UO_831 (O_831,N_19851,N_16511);
and UO_832 (O_832,N_16722,N_18998);
nand UO_833 (O_833,N_16793,N_19494);
nor UO_834 (O_834,N_17148,N_18551);
and UO_835 (O_835,N_17499,N_19331);
nand UO_836 (O_836,N_17206,N_16782);
nand UO_837 (O_837,N_17635,N_19361);
nor UO_838 (O_838,N_19039,N_16248);
nand UO_839 (O_839,N_19350,N_17827);
nor UO_840 (O_840,N_18519,N_16087);
or UO_841 (O_841,N_16255,N_16381);
and UO_842 (O_842,N_19918,N_17673);
nor UO_843 (O_843,N_18949,N_19849);
and UO_844 (O_844,N_17795,N_18137);
nand UO_845 (O_845,N_17522,N_16801);
nand UO_846 (O_846,N_18718,N_19457);
nand UO_847 (O_847,N_19670,N_18000);
or UO_848 (O_848,N_18074,N_17608);
nand UO_849 (O_849,N_19181,N_17316);
nor UO_850 (O_850,N_16728,N_19324);
nor UO_851 (O_851,N_19388,N_17262);
or UO_852 (O_852,N_19945,N_16714);
or UO_853 (O_853,N_19075,N_18841);
nor UO_854 (O_854,N_18672,N_16421);
nand UO_855 (O_855,N_19725,N_19448);
and UO_856 (O_856,N_16861,N_18422);
nor UO_857 (O_857,N_17400,N_17578);
nor UO_858 (O_858,N_19947,N_18346);
nand UO_859 (O_859,N_18730,N_17774);
and UO_860 (O_860,N_17951,N_16770);
nor UO_861 (O_861,N_18796,N_19190);
and UO_862 (O_862,N_17862,N_17006);
nand UO_863 (O_863,N_19502,N_16293);
nand UO_864 (O_864,N_16450,N_19944);
or UO_865 (O_865,N_17314,N_16205);
nand UO_866 (O_866,N_16332,N_17411);
or UO_867 (O_867,N_16601,N_17644);
or UO_868 (O_868,N_19336,N_16002);
or UO_869 (O_869,N_18186,N_17788);
nor UO_870 (O_870,N_17073,N_19585);
and UO_871 (O_871,N_18119,N_16908);
nand UO_872 (O_872,N_18821,N_18332);
nand UO_873 (O_873,N_16494,N_17946);
or UO_874 (O_874,N_19115,N_16018);
nor UO_875 (O_875,N_16079,N_17817);
xor UO_876 (O_876,N_18834,N_17060);
and UO_877 (O_877,N_18923,N_17417);
and UO_878 (O_878,N_17626,N_19078);
nor UO_879 (O_879,N_16315,N_16213);
or UO_880 (O_880,N_18527,N_18574);
or UO_881 (O_881,N_16179,N_18147);
xor UO_882 (O_882,N_17911,N_16576);
nor UO_883 (O_883,N_18791,N_18467);
or UO_884 (O_884,N_16954,N_17193);
or UO_885 (O_885,N_19627,N_19355);
nand UO_886 (O_886,N_19016,N_17374);
and UO_887 (O_887,N_17913,N_17727);
nor UO_888 (O_888,N_17967,N_19852);
or UO_889 (O_889,N_18423,N_16762);
and UO_890 (O_890,N_19651,N_16335);
nand UO_891 (O_891,N_19049,N_19354);
nand UO_892 (O_892,N_17706,N_16464);
nand UO_893 (O_893,N_19414,N_18981);
nor UO_894 (O_894,N_18520,N_16949);
nor UO_895 (O_895,N_17095,N_16923);
and UO_896 (O_896,N_19522,N_19813);
xor UO_897 (O_897,N_17577,N_18994);
nand UO_898 (O_898,N_18651,N_19833);
nor UO_899 (O_899,N_16418,N_18560);
or UO_900 (O_900,N_17761,N_16201);
nand UO_901 (O_901,N_17402,N_18384);
or UO_902 (O_902,N_16953,N_18507);
nand UO_903 (O_903,N_16734,N_19806);
and UO_904 (O_904,N_16176,N_17187);
xnor UO_905 (O_905,N_17130,N_17437);
nor UO_906 (O_906,N_18648,N_19117);
and UO_907 (O_907,N_19490,N_19272);
nor UO_908 (O_908,N_17521,N_16944);
and UO_909 (O_909,N_16723,N_16848);
nand UO_910 (O_910,N_17621,N_19896);
nor UO_911 (O_911,N_16551,N_18930);
and UO_912 (O_912,N_19819,N_19161);
nor UO_913 (O_913,N_17378,N_17875);
nor UO_914 (O_914,N_16751,N_17032);
nand UO_915 (O_915,N_18548,N_16388);
nor UO_916 (O_916,N_16244,N_17614);
and UO_917 (O_917,N_19003,N_16743);
or UO_918 (O_918,N_19158,N_16524);
or UO_919 (O_919,N_17015,N_17069);
or UO_920 (O_920,N_16423,N_18936);
nand UO_921 (O_921,N_17856,N_17462);
nand UO_922 (O_922,N_17912,N_18809);
xor UO_923 (O_923,N_19582,N_19319);
or UO_924 (O_924,N_16403,N_19913);
nand UO_925 (O_925,N_18452,N_19655);
nor UO_926 (O_926,N_16271,N_17730);
nand UO_927 (O_927,N_18677,N_19540);
nor UO_928 (O_928,N_17204,N_16285);
and UO_929 (O_929,N_19197,N_17787);
or UO_930 (O_930,N_17191,N_18990);
or UO_931 (O_931,N_16058,N_19148);
nand UO_932 (O_932,N_17792,N_19433);
xnor UO_933 (O_933,N_16117,N_19723);
and UO_934 (O_934,N_16073,N_17195);
nor UO_935 (O_935,N_16056,N_17748);
nand UO_936 (O_936,N_17616,N_16443);
xnor UO_937 (O_937,N_16436,N_18398);
xnor UO_938 (O_938,N_16599,N_17028);
nor UO_939 (O_939,N_17969,N_18143);
or UO_940 (O_940,N_19916,N_16037);
or UO_941 (O_941,N_16771,N_16364);
or UO_942 (O_942,N_18352,N_19513);
nand UO_943 (O_943,N_18563,N_16556);
or UO_944 (O_944,N_18746,N_19323);
or UO_945 (O_945,N_18916,N_16101);
nor UO_946 (O_946,N_19634,N_17305);
xor UO_947 (O_947,N_16773,N_18023);
or UO_948 (O_948,N_17387,N_17284);
or UO_949 (O_949,N_19707,N_17634);
and UO_950 (O_950,N_16625,N_18190);
and UO_951 (O_951,N_16914,N_16658);
nor UO_952 (O_952,N_16136,N_17553);
nand UO_953 (O_953,N_19985,N_16174);
or UO_954 (O_954,N_17821,N_18312);
nor UO_955 (O_955,N_18153,N_16374);
or UO_956 (O_956,N_19176,N_19426);
nand UO_957 (O_957,N_17745,N_17405);
and UO_958 (O_958,N_17372,N_19810);
nand UO_959 (O_959,N_16919,N_16014);
or UO_960 (O_960,N_18954,N_16034);
nor UO_961 (O_961,N_19275,N_16503);
nand UO_962 (O_962,N_18072,N_17044);
nand UO_963 (O_963,N_17679,N_16112);
xnor UO_964 (O_964,N_18597,N_17504);
nor UO_965 (O_965,N_18170,N_17125);
or UO_966 (O_966,N_18174,N_19404);
nand UO_967 (O_967,N_18784,N_16139);
xnor UO_968 (O_968,N_19479,N_16137);
and UO_969 (O_969,N_18965,N_16440);
and UO_970 (O_970,N_18907,N_19192);
or UO_971 (O_971,N_19867,N_16985);
and UO_972 (O_972,N_19413,N_17318);
nor UO_973 (O_973,N_19344,N_18084);
and UO_974 (O_974,N_16973,N_18261);
and UO_975 (O_975,N_17563,N_16602);
or UO_976 (O_976,N_18122,N_16177);
or UO_977 (O_977,N_16990,N_19934);
nor UO_978 (O_978,N_16566,N_17065);
nand UO_979 (O_979,N_19041,N_18328);
and UO_980 (O_980,N_16072,N_18714);
nand UO_981 (O_981,N_16219,N_16363);
nand UO_982 (O_982,N_18927,N_18884);
nor UO_983 (O_983,N_18417,N_18306);
or UO_984 (O_984,N_16616,N_17971);
or UO_985 (O_985,N_18285,N_19391);
nand UO_986 (O_986,N_18209,N_17643);
nor UO_987 (O_987,N_19282,N_19300);
and UO_988 (O_988,N_18316,N_18217);
and UO_989 (O_989,N_18627,N_18883);
nand UO_990 (O_990,N_19129,N_18371);
and UO_991 (O_991,N_16653,N_18364);
nor UO_992 (O_992,N_18736,N_19671);
nand UO_993 (O_993,N_19371,N_16885);
and UO_994 (O_994,N_19872,N_16634);
nor UO_995 (O_995,N_16076,N_16277);
or UO_996 (O_996,N_17166,N_19920);
nand UO_997 (O_997,N_17249,N_17127);
nand UO_998 (O_998,N_16870,N_18653);
and UO_999 (O_999,N_18939,N_18846);
or UO_1000 (O_1000,N_17786,N_17642);
nand UO_1001 (O_1001,N_17579,N_17863);
xor UO_1002 (O_1002,N_17441,N_19946);
or UO_1003 (O_1003,N_16586,N_16114);
and UO_1004 (O_1004,N_16282,N_17868);
nor UO_1005 (O_1005,N_17583,N_19400);
xor UO_1006 (O_1006,N_16878,N_18555);
nor UO_1007 (O_1007,N_18028,N_19318);
nor UO_1008 (O_1008,N_19564,N_18917);
and UO_1009 (O_1009,N_18008,N_16600);
nor UO_1010 (O_1010,N_16453,N_16741);
xor UO_1011 (O_1011,N_18349,N_17443);
and UO_1012 (O_1012,N_19411,N_17989);
nor UO_1013 (O_1013,N_16337,N_19793);
nand UO_1014 (O_1014,N_18963,N_16660);
or UO_1015 (O_1015,N_16359,N_17241);
or UO_1016 (O_1016,N_17093,N_19639);
nand UO_1017 (O_1017,N_18820,N_17012);
or UO_1018 (O_1018,N_17293,N_18594);
and UO_1019 (O_1019,N_17702,N_19313);
nor UO_1020 (O_1020,N_17711,N_18057);
and UO_1021 (O_1021,N_18251,N_17144);
nand UO_1022 (O_1022,N_16970,N_19147);
nand UO_1023 (O_1023,N_17389,N_19836);
and UO_1024 (O_1024,N_17020,N_16699);
xor UO_1025 (O_1025,N_16431,N_17149);
and UO_1026 (O_1026,N_17908,N_18959);
nand UO_1027 (O_1027,N_16224,N_17726);
or UO_1028 (O_1028,N_16385,N_17047);
nand UO_1029 (O_1029,N_18184,N_18192);
or UO_1030 (O_1030,N_19892,N_16719);
and UO_1031 (O_1031,N_18687,N_17313);
and UO_1032 (O_1032,N_18697,N_18591);
nand UO_1033 (O_1033,N_19791,N_16302);
or UO_1034 (O_1034,N_19476,N_16604);
nand UO_1035 (O_1035,N_16739,N_16945);
nor UO_1036 (O_1036,N_16927,N_18159);
and UO_1037 (O_1037,N_19284,N_18509);
nand UO_1038 (O_1038,N_19295,N_17758);
nand UO_1039 (O_1039,N_19778,N_17902);
nor UO_1040 (O_1040,N_19767,N_17490);
or UO_1041 (O_1041,N_16668,N_17110);
nand UO_1042 (O_1042,N_17211,N_17743);
and UO_1043 (O_1043,N_19511,N_18508);
nor UO_1044 (O_1044,N_16188,N_18818);
nand UO_1045 (O_1045,N_16249,N_19855);
and UO_1046 (O_1046,N_18307,N_17285);
or UO_1047 (O_1047,N_16638,N_17431);
or UO_1048 (O_1048,N_17832,N_18449);
or UO_1049 (O_1049,N_16357,N_17317);
nand UO_1050 (O_1050,N_17898,N_17114);
and UO_1051 (O_1051,N_16412,N_19973);
nand UO_1052 (O_1052,N_18487,N_17876);
nor UO_1053 (O_1053,N_18739,N_16269);
nand UO_1054 (O_1054,N_16038,N_19974);
or UO_1055 (O_1055,N_19507,N_19258);
and UO_1056 (O_1056,N_18426,N_17750);
nand UO_1057 (O_1057,N_18888,N_17406);
nor UO_1058 (O_1058,N_18129,N_17754);
or UO_1059 (O_1059,N_19843,N_17368);
and UO_1060 (O_1060,N_18656,N_18750);
nand UO_1061 (O_1061,N_17016,N_18502);
nand UO_1062 (O_1062,N_17555,N_17689);
nand UO_1063 (O_1063,N_16904,N_19210);
or UO_1064 (O_1064,N_17523,N_19682);
or UO_1065 (O_1065,N_16683,N_16805);
xnor UO_1066 (O_1066,N_19219,N_16568);
nor UO_1067 (O_1067,N_16413,N_16784);
nor UO_1068 (O_1068,N_16082,N_16829);
nor UO_1069 (O_1069,N_16968,N_18428);
and UO_1070 (O_1070,N_17271,N_18510);
and UO_1071 (O_1071,N_16296,N_17631);
or UO_1072 (O_1072,N_19263,N_17618);
nand UO_1073 (O_1073,N_18747,N_18541);
xnor UO_1074 (O_1074,N_18125,N_19094);
nor UO_1075 (O_1075,N_19712,N_18737);
xor UO_1076 (O_1076,N_16175,N_19817);
or UO_1077 (O_1077,N_18668,N_18749);
or UO_1078 (O_1078,N_17983,N_17895);
and UO_1079 (O_1079,N_17340,N_19783);
or UO_1080 (O_1080,N_19700,N_16535);
nand UO_1081 (O_1081,N_16144,N_18016);
or UO_1082 (O_1082,N_17622,N_16606);
xnor UO_1083 (O_1083,N_19545,N_19396);
nor UO_1084 (O_1084,N_18078,N_18669);
nor UO_1085 (O_1085,N_16984,N_17615);
nor UO_1086 (O_1086,N_17810,N_19326);
nor UO_1087 (O_1087,N_17878,N_18775);
and UO_1088 (O_1088,N_19942,N_17829);
nand UO_1089 (O_1089,N_16899,N_18379);
and UO_1090 (O_1090,N_18762,N_16417);
xor UO_1091 (O_1091,N_17279,N_19968);
nor UO_1092 (O_1092,N_19638,N_19977);
and UO_1093 (O_1093,N_16827,N_16982);
nand UO_1094 (O_1094,N_16920,N_19108);
and UO_1095 (O_1095,N_18966,N_17088);
or UO_1096 (O_1096,N_18683,N_17049);
nor UO_1097 (O_1097,N_19689,N_18763);
or UO_1098 (O_1098,N_17501,N_17572);
or UO_1099 (O_1099,N_16559,N_16334);
and UO_1100 (O_1100,N_19719,N_19620);
nand UO_1101 (O_1101,N_16378,N_17528);
nand UO_1102 (O_1102,N_17113,N_18827);
or UO_1103 (O_1103,N_17587,N_17776);
and UO_1104 (O_1104,N_17772,N_17503);
xnor UO_1105 (O_1105,N_18194,N_16781);
nor UO_1106 (O_1106,N_18967,N_19239);
nor UO_1107 (O_1107,N_16819,N_16446);
nand UO_1108 (O_1108,N_16565,N_19347);
nor UO_1109 (O_1109,N_17712,N_19938);
nor UO_1110 (O_1110,N_18455,N_19528);
nand UO_1111 (O_1111,N_19017,N_19154);
or UO_1112 (O_1112,N_16742,N_19465);
nand UO_1113 (O_1113,N_19212,N_16202);
nand UO_1114 (O_1114,N_17859,N_18722);
or UO_1115 (O_1115,N_19654,N_16593);
and UO_1116 (O_1116,N_18247,N_17491);
nor UO_1117 (O_1117,N_16211,N_16321);
nor UO_1118 (O_1118,N_16070,N_17438);
or UO_1119 (O_1119,N_16501,N_19102);
or UO_1120 (O_1120,N_18448,N_17604);
and UO_1121 (O_1121,N_17507,N_18538);
nor UO_1122 (O_1122,N_17995,N_16042);
and UO_1123 (O_1123,N_19656,N_19309);
and UO_1124 (O_1124,N_18517,N_18953);
nand UO_1125 (O_1125,N_16199,N_18977);
nand UO_1126 (O_1126,N_19252,N_16840);
and UO_1127 (O_1127,N_17245,N_18210);
nand UO_1128 (O_1128,N_17397,N_17502);
nand UO_1129 (O_1129,N_19815,N_18896);
nand UO_1130 (O_1130,N_16609,N_16005);
xor UO_1131 (O_1131,N_17940,N_17105);
xnor UO_1132 (O_1132,N_16872,N_19441);
or UO_1133 (O_1133,N_17143,N_16420);
or UO_1134 (O_1134,N_18847,N_18579);
nor UO_1135 (O_1135,N_17180,N_16648);
nand UO_1136 (O_1136,N_18282,N_19983);
nor UO_1137 (O_1137,N_18274,N_17980);
nor UO_1138 (O_1138,N_18601,N_18685);
xor UO_1139 (O_1139,N_16614,N_16479);
nor UO_1140 (O_1140,N_16817,N_17270);
and UO_1141 (O_1141,N_16409,N_18075);
nor UO_1142 (O_1142,N_18407,N_16522);
and UO_1143 (O_1143,N_17747,N_19128);
or UO_1144 (O_1144,N_17136,N_17379);
nand UO_1145 (O_1145,N_16948,N_17897);
or UO_1146 (O_1146,N_16458,N_17565);
and UO_1147 (O_1147,N_16092,N_18645);
and UO_1148 (O_1148,N_16678,N_18215);
nor UO_1149 (O_1149,N_19364,N_18462);
nand UO_1150 (O_1150,N_18324,N_16068);
or UO_1151 (O_1151,N_16900,N_19626);
nor UO_1152 (O_1152,N_17991,N_19897);
and UO_1153 (O_1153,N_17330,N_16386);
nor UO_1154 (O_1154,N_19135,N_16373);
and UO_1155 (O_1155,N_19747,N_18368);
nor UO_1156 (O_1156,N_17385,N_17361);
nand UO_1157 (O_1157,N_16889,N_19370);
nand UO_1158 (O_1158,N_16567,N_18975);
xnor UO_1159 (O_1159,N_19491,N_19170);
and UO_1160 (O_1160,N_16512,N_16977);
and UO_1161 (O_1161,N_17476,N_18205);
or UO_1162 (O_1162,N_18709,N_17887);
and UO_1163 (O_1163,N_16649,N_19327);
and UO_1164 (O_1164,N_17909,N_17970);
or UO_1165 (O_1165,N_17708,N_19296);
xnor UO_1166 (O_1166,N_19139,N_16394);
nand UO_1167 (O_1167,N_18812,N_17802);
nor UO_1168 (O_1168,N_16257,N_16785);
nor UO_1169 (O_1169,N_19532,N_18544);
nor UO_1170 (O_1170,N_19951,N_16809);
and UO_1171 (O_1171,N_19978,N_16627);
nor UO_1172 (O_1172,N_17517,N_16880);
and UO_1173 (O_1173,N_17569,N_19909);
or UO_1174 (O_1174,N_17010,N_17429);
nor UO_1175 (O_1175,N_16884,N_17346);
and UO_1176 (O_1176,N_18902,N_16389);
or UO_1177 (O_1177,N_17515,N_17237);
nand UO_1178 (O_1178,N_16822,N_19529);
xor UO_1179 (O_1179,N_18898,N_19733);
nor UO_1180 (O_1180,N_19777,N_17835);
nand UO_1181 (O_1181,N_18585,N_18193);
nor UO_1182 (O_1182,N_18160,N_19902);
nand UO_1183 (O_1183,N_16570,N_19986);
and UO_1184 (O_1184,N_17790,N_17106);
xor UO_1185 (O_1185,N_17573,N_17228);
or UO_1186 (O_1186,N_19929,N_17207);
xnor UO_1187 (O_1187,N_19802,N_18268);
nor UO_1188 (O_1188,N_19770,N_17160);
xnor UO_1189 (O_1189,N_19204,N_17435);
xnor UO_1190 (O_1190,N_19257,N_19090);
and UO_1191 (O_1191,N_19868,N_17456);
and UO_1192 (O_1192,N_16486,N_16541);
nand UO_1193 (O_1193,N_18774,N_19891);
xnor UO_1194 (O_1194,N_17633,N_16655);
and UO_1195 (O_1195,N_17652,N_19742);
or UO_1196 (O_1196,N_19153,N_18266);
or UO_1197 (O_1197,N_19030,N_16992);
or UO_1198 (O_1198,N_18781,N_19138);
nand UO_1199 (O_1199,N_19403,N_19387);
and UO_1200 (O_1200,N_19807,N_16583);
and UO_1201 (O_1201,N_18864,N_18704);
and UO_1202 (O_1202,N_16621,N_16691);
xor UO_1203 (O_1203,N_17273,N_16855);
and UO_1204 (O_1204,N_16160,N_18696);
xnor UO_1205 (O_1205,N_19036,N_19988);
xor UO_1206 (O_1206,N_18868,N_18196);
and UO_1207 (O_1207,N_18925,N_19299);
nand UO_1208 (O_1208,N_18501,N_19584);
or UO_1209 (O_1209,N_16913,N_17820);
nand UO_1210 (O_1210,N_16143,N_18940);
nor UO_1211 (O_1211,N_18873,N_18472);
nand UO_1212 (O_1212,N_18348,N_19301);
nand UO_1213 (O_1213,N_18414,N_17955);
or UO_1214 (O_1214,N_19099,N_17609);
or UO_1215 (O_1215,N_17382,N_16475);
nor UO_1216 (O_1216,N_16430,N_19679);
nand UO_1217 (O_1217,N_17409,N_16686);
or UO_1218 (O_1218,N_16091,N_19590);
or UO_1219 (O_1219,N_17302,N_19612);
or UO_1220 (O_1220,N_18682,N_18394);
or UO_1221 (O_1221,N_17846,N_17475);
or UO_1222 (O_1222,N_19841,N_18822);
and UO_1223 (O_1223,N_17766,N_18552);
xnor UO_1224 (O_1224,N_18569,N_18602);
or UO_1225 (O_1225,N_19949,N_19418);
nand UO_1226 (O_1226,N_18064,N_19596);
and UO_1227 (O_1227,N_19858,N_17189);
nor UO_1228 (O_1228,N_18536,N_18612);
and UO_1229 (O_1229,N_16233,N_18321);
xnor UO_1230 (O_1230,N_18011,N_19080);
and UO_1231 (O_1231,N_19066,N_19256);
or UO_1232 (O_1232,N_16892,N_18453);
or UO_1233 (O_1233,N_18135,N_18486);
or UO_1234 (O_1234,N_18671,N_18630);
or UO_1235 (O_1235,N_16735,N_16729);
nor UO_1236 (O_1236,N_17575,N_16250);
and UO_1237 (O_1237,N_18702,N_16341);
and UO_1238 (O_1238,N_19189,N_18189);
nor UO_1239 (O_1239,N_18708,N_18860);
nor UO_1240 (O_1240,N_18350,N_17547);
and UO_1241 (O_1241,N_17924,N_19724);
xor UO_1242 (O_1242,N_18666,N_16247);
or UO_1243 (O_1243,N_17168,N_16932);
or UO_1244 (O_1244,N_17719,N_19499);
xnor UO_1245 (O_1245,N_19658,N_16934);
nand UO_1246 (O_1246,N_18578,N_18875);
nand UO_1247 (O_1247,N_18580,N_16962);
nor UO_1248 (O_1248,N_18336,N_19616);
or UO_1249 (O_1249,N_19482,N_17256);
or UO_1250 (O_1250,N_18496,N_16679);
nor UO_1251 (O_1251,N_16673,N_17118);
or UO_1252 (O_1252,N_19861,N_18802);
nor UO_1253 (O_1253,N_19741,N_18799);
nor UO_1254 (O_1254,N_18253,N_19775);
nor UO_1255 (O_1255,N_19956,N_19765);
xor UO_1256 (O_1256,N_19031,N_18030);
or UO_1257 (O_1257,N_18025,N_19055);
nor UO_1258 (O_1258,N_17663,N_19488);
nand UO_1259 (O_1259,N_17641,N_16428);
nor UO_1260 (O_1260,N_19981,N_18596);
nand UO_1261 (O_1261,N_17840,N_19461);
and UO_1262 (O_1262,N_18019,N_19225);
or UO_1263 (O_1263,N_19033,N_19659);
xnor UO_1264 (O_1264,N_19096,N_17304);
xnor UO_1265 (O_1265,N_18167,N_19292);
nand UO_1266 (O_1266,N_16300,N_18344);
nor UO_1267 (O_1267,N_19048,N_16960);
nor UO_1268 (O_1268,N_18614,N_16258);
nor UO_1269 (O_1269,N_16961,N_17653);
and UO_1270 (O_1270,N_19211,N_16132);
nor UO_1271 (O_1271,N_16488,N_19432);
and UO_1272 (O_1272,N_18202,N_19175);
nand UO_1273 (O_1273,N_19844,N_17488);
and UO_1274 (O_1274,N_19334,N_18765);
nand UO_1275 (O_1275,N_19548,N_17668);
nand UO_1276 (O_1276,N_18152,N_19395);
and UO_1277 (O_1277,N_17092,N_18752);
nor UO_1278 (O_1278,N_16003,N_17637);
xnor UO_1279 (O_1279,N_16875,N_17213);
nand UO_1280 (O_1280,N_17926,N_17598);
nand UO_1281 (O_1281,N_16558,N_19332);
nand UO_1282 (O_1282,N_19086,N_17837);
nand UO_1283 (O_1283,N_16262,N_17341);
xnor UO_1284 (O_1284,N_18779,N_16718);
nand UO_1285 (O_1285,N_18039,N_16868);
xnor UO_1286 (O_1286,N_18197,N_19038);
or UO_1287 (O_1287,N_18178,N_16362);
or UO_1288 (O_1288,N_16917,N_17703);
or UO_1289 (O_1289,N_19351,N_17156);
nand UO_1290 (O_1290,N_17274,N_18042);
nor UO_1291 (O_1291,N_16632,N_18565);
and UO_1292 (O_1292,N_17133,N_19294);
nand UO_1293 (O_1293,N_18831,N_18113);
nand UO_1294 (O_1294,N_18961,N_18992);
nand UO_1295 (O_1295,N_18383,N_17698);
nor UO_1296 (O_1296,N_18037,N_17375);
nor UO_1297 (O_1297,N_17733,N_16080);
nor UO_1298 (O_1298,N_18845,N_18132);
and UO_1299 (O_1299,N_17949,N_18974);
nor UO_1300 (O_1300,N_16157,N_16140);
and UO_1301 (O_1301,N_16036,N_17055);
nor UO_1302 (O_1302,N_17322,N_19701);
and UO_1303 (O_1303,N_16180,N_16167);
and UO_1304 (O_1304,N_19959,N_17801);
nand UO_1305 (O_1305,N_18726,N_18195);
or UO_1306 (O_1306,N_17904,N_19009);
nand UO_1307 (O_1307,N_17561,N_17683);
nand UO_1308 (O_1308,N_16081,N_17426);
nand UO_1309 (O_1309,N_18767,N_17789);
and UO_1310 (O_1310,N_19568,N_18034);
or UO_1311 (O_1311,N_16238,N_18070);
nor UO_1312 (O_1312,N_17688,N_19113);
nor UO_1313 (O_1313,N_18777,N_19591);
nand UO_1314 (O_1314,N_16797,N_19244);
and UO_1315 (O_1315,N_17627,N_17510);
nor UO_1316 (O_1316,N_18899,N_19449);
and UO_1317 (O_1317,N_19826,N_16543);
or UO_1318 (O_1318,N_19372,N_18604);
and UO_1319 (O_1319,N_18635,N_16194);
nor UO_1320 (O_1320,N_19471,N_17765);
nand UO_1321 (O_1321,N_19132,N_16406);
or UO_1322 (O_1322,N_18893,N_17536);
nand UO_1323 (O_1323,N_19251,N_19082);
xnor UO_1324 (O_1324,N_16575,N_17977);
nand UO_1325 (O_1325,N_18459,N_17170);
and UO_1326 (O_1326,N_16461,N_18081);
or UO_1327 (O_1327,N_16507,N_16142);
nand UO_1328 (O_1328,N_19443,N_18956);
nor UO_1329 (O_1329,N_19242,N_19680);
nor UO_1330 (O_1330,N_16894,N_18139);
or UO_1331 (O_1331,N_17918,N_17975);
and UO_1332 (O_1332,N_18370,N_17982);
and UO_1333 (O_1333,N_18598,N_16591);
nor UO_1334 (O_1334,N_17250,N_17691);
nor UO_1335 (O_1335,N_16915,N_16536);
or UO_1336 (O_1336,N_17685,N_19028);
nand UO_1337 (O_1337,N_17263,N_18690);
nor UO_1338 (O_1338,N_18322,N_19126);
or UO_1339 (O_1339,N_16557,N_17576);
and UO_1340 (O_1340,N_19728,N_16305);
and UO_1341 (O_1341,N_19911,N_17451);
and UO_1342 (O_1342,N_17159,N_16107);
or UO_1343 (O_1343,N_16554,N_19481);
nand UO_1344 (O_1344,N_17513,N_18103);
nand UO_1345 (O_1345,N_16288,N_17544);
nor UO_1346 (O_1346,N_16647,N_17420);
nand UO_1347 (O_1347,N_18249,N_19169);
and UO_1348 (O_1348,N_19645,N_17404);
and UO_1349 (O_1349,N_19495,N_16054);
or UO_1350 (O_1350,N_16740,N_17014);
nor UO_1351 (O_1351,N_19477,N_19083);
or UO_1352 (O_1352,N_19091,N_16497);
and UO_1353 (O_1353,N_18539,N_18267);
nand UO_1354 (O_1354,N_19743,N_18742);
nand UO_1355 (O_1355,N_18759,N_19431);
and UO_1356 (O_1356,N_17383,N_19887);
xnor UO_1357 (O_1357,N_18948,N_16165);
and UO_1358 (O_1358,N_18634,N_19746);
or UO_1359 (O_1359,N_16401,N_18554);
and UO_1360 (O_1360,N_17757,N_18609);
nand UO_1361 (O_1361,N_16462,N_18172);
or UO_1362 (O_1362,N_19202,N_16169);
xor UO_1363 (O_1363,N_18817,N_19010);
nor UO_1364 (O_1364,N_19521,N_18434);
nand UO_1365 (O_1365,N_18955,N_19857);
and UO_1366 (O_1366,N_17424,N_18921);
nor UO_1367 (O_1367,N_18876,N_17328);
nand UO_1368 (O_1368,N_17628,N_18850);
xor UO_1369 (O_1369,N_16086,N_18556);
or UO_1370 (O_1370,N_16790,N_18679);
or UO_1371 (O_1371,N_18608,N_16346);
or UO_1372 (O_1372,N_18558,N_16552);
nor UO_1373 (O_1373,N_17717,N_17045);
or UO_1374 (O_1374,N_17401,N_19337);
nor UO_1375 (O_1375,N_16561,N_18026);
and UO_1376 (O_1376,N_16104,N_19704);
nand UO_1377 (O_1377,N_16663,N_19216);
nor UO_1378 (O_1378,N_16639,N_19379);
nor UO_1379 (O_1379,N_16000,N_17709);
and UO_1380 (O_1380,N_19325,N_18228);
nand UO_1381 (O_1381,N_17324,N_16090);
xor UO_1382 (O_1382,N_16749,N_16727);
or UO_1383 (O_1383,N_16972,N_19100);
nand UO_1384 (O_1384,N_19751,N_18589);
and UO_1385 (O_1385,N_18503,N_16314);
or UO_1386 (O_1386,N_18112,N_17731);
and UO_1387 (O_1387,N_18297,N_19549);
or UO_1388 (O_1388,N_19492,N_17864);
or UO_1389 (O_1389,N_19057,N_17433);
or UO_1390 (O_1390,N_16451,N_19307);
or UO_1391 (O_1391,N_16168,N_16651);
and UO_1392 (O_1392,N_19259,N_17966);
xnor UO_1393 (O_1393,N_16306,N_19173);
nor UO_1394 (O_1394,N_19681,N_19421);
and UO_1395 (O_1395,N_16836,N_18573);
or UO_1396 (O_1396,N_19761,N_17370);
nand UO_1397 (O_1397,N_19676,N_19512);
nor UO_1398 (O_1398,N_19593,N_17916);
xor UO_1399 (O_1399,N_17770,N_16322);
or UO_1400 (O_1400,N_17525,N_17632);
nand UO_1401 (O_1401,N_16369,N_18158);
or UO_1402 (O_1402,N_17033,N_18073);
and UO_1403 (O_1403,N_19298,N_17246);
or UO_1404 (O_1404,N_17421,N_16396);
and UO_1405 (O_1405,N_16754,N_16405);
or UO_1406 (O_1406,N_17567,N_16333);
or UO_1407 (O_1407,N_17981,N_17150);
or UO_1408 (O_1408,N_16672,N_18288);
xor UO_1409 (O_1409,N_19245,N_19808);
nand UO_1410 (O_1410,N_17905,N_17542);
nor UO_1411 (O_1411,N_16788,N_19459);
and UO_1412 (O_1412,N_16661,N_17096);
nand UO_1413 (O_1413,N_16650,N_19943);
nor UO_1414 (O_1414,N_19829,N_16548);
or UO_1415 (O_1415,N_16733,N_18240);
nor UO_1416 (O_1416,N_17052,N_18676);
nand UO_1417 (O_1417,N_17056,N_18647);
xnor UO_1418 (O_1418,N_19508,N_18278);
or UO_1419 (O_1419,N_16981,N_16103);
and UO_1420 (O_1420,N_18724,N_16580);
and UO_1421 (O_1421,N_19392,N_19895);
or UO_1422 (O_1422,N_16343,N_17367);
nor UO_1423 (O_1423,N_18284,N_16596);
or UO_1424 (O_1424,N_18115,N_19979);
and UO_1425 (O_1425,N_19960,N_18654);
and UO_1426 (O_1426,N_18109,N_18830);
or UO_1427 (O_1427,N_16881,N_18903);
and UO_1428 (O_1428,N_17591,N_17901);
or UO_1429 (O_1429,N_18071,N_16071);
or UO_1430 (O_1430,N_18894,N_16040);
nand UO_1431 (O_1431,N_18869,N_18429);
nand UO_1432 (O_1432,N_19926,N_18768);
or UO_1433 (O_1433,N_18385,N_19235);
nand UO_1434 (O_1434,N_16578,N_17453);
and UO_1435 (O_1435,N_19850,N_18770);
or UO_1436 (O_1436,N_16478,N_16063);
or UO_1437 (O_1437,N_17782,N_17701);
or UO_1438 (O_1438,N_19898,N_17927);
or UO_1439 (O_1439,N_16266,N_17139);
xor UO_1440 (O_1440,N_19531,N_19046);
and UO_1441 (O_1441,N_19907,N_18978);
nand UO_1442 (O_1442,N_16746,N_16608);
and UO_1443 (O_1443,N_16414,N_16681);
nand UO_1444 (O_1444,N_17369,N_17505);
nand UO_1445 (O_1445,N_17722,N_18800);
nand UO_1446 (O_1446,N_18840,N_17917);
nor UO_1447 (O_1447,N_19594,N_18595);
and UO_1448 (O_1448,N_17024,N_17469);
nor UO_1449 (O_1449,N_18905,N_17035);
or UO_1450 (O_1450,N_18318,N_18131);
nor UO_1451 (O_1451,N_16397,N_17333);
nand UO_1452 (O_1452,N_17075,N_19378);
xor UO_1453 (O_1453,N_16967,N_17108);
xnor UO_1454 (O_1454,N_16612,N_19310);
and UO_1455 (O_1455,N_19601,N_19274);
xnor UO_1456 (O_1456,N_19673,N_18111);
nand UO_1457 (O_1457,N_17694,N_16572);
nand UO_1458 (O_1458,N_16974,N_16804);
or UO_1459 (O_1459,N_18533,N_17669);
nand UO_1460 (O_1460,N_17524,N_16710);
nand UO_1461 (O_1461,N_19342,N_18633);
or UO_1462 (O_1462,N_18415,N_17700);
and UO_1463 (O_1463,N_16563,N_17539);
nor UO_1464 (O_1464,N_19254,N_17558);
or UO_1465 (O_1465,N_19784,N_17816);
nand UO_1466 (O_1466,N_17342,N_16498);
nand UO_1467 (O_1467,N_16026,N_17275);
and UO_1468 (O_1468,N_17101,N_18114);
nand UO_1469 (O_1469,N_19349,N_17695);
and UO_1470 (O_1470,N_16969,N_16534);
or UO_1471 (O_1471,N_16347,N_18534);
nand UO_1472 (O_1472,N_16689,N_18012);
or UO_1473 (O_1473,N_16676,N_16857);
nand UO_1474 (O_1474,N_19553,N_17267);
and UO_1475 (O_1475,N_19587,N_18881);
and UO_1476 (O_1476,N_18117,N_18176);
nand UO_1477 (O_1477,N_17675,N_17094);
nor UO_1478 (O_1478,N_17752,N_17408);
xor UO_1479 (O_1479,N_17813,N_16429);
and UO_1480 (O_1480,N_19044,N_16882);
nor UO_1481 (O_1481,N_17412,N_19452);
nor UO_1482 (O_1482,N_19506,N_17236);
nand UO_1483 (O_1483,N_19208,N_17541);
xor UO_1484 (O_1484,N_17137,N_17403);
nor UO_1485 (O_1485,N_16031,N_19463);
or UO_1486 (O_1486,N_18097,N_16489);
or UO_1487 (O_1487,N_18788,N_16866);
nand UO_1488 (O_1488,N_18941,N_18166);
xor UO_1489 (O_1489,N_19019,N_16241);
xor UO_1490 (O_1490,N_17287,N_19409);
nand UO_1491 (O_1491,N_17948,N_18498);
nor UO_1492 (O_1492,N_16873,N_18355);
nor UO_1493 (O_1493,N_17532,N_17952);
nand UO_1494 (O_1494,N_18506,N_18926);
or UO_1495 (O_1495,N_19631,N_17292);
or UO_1496 (O_1496,N_19264,N_16637);
nor UO_1497 (O_1497,N_18674,N_17930);
nand UO_1498 (O_1498,N_17990,N_19608);
nand UO_1499 (O_1499,N_18014,N_17470);
or UO_1500 (O_1500,N_16164,N_18157);
xor UO_1501 (O_1501,N_16499,N_18036);
and UO_1502 (O_1502,N_19732,N_19762);
xnor UO_1503 (O_1503,N_19661,N_17984);
or UO_1504 (O_1504,N_16795,N_16931);
nor UO_1505 (O_1505,N_16097,N_18032);
and UO_1506 (O_1506,N_18150,N_17255);
nor UO_1507 (O_1507,N_17173,N_17296);
nand UO_1508 (O_1508,N_19744,N_18550);
and UO_1509 (O_1509,N_18691,N_16594);
or UO_1510 (O_1510,N_18660,N_19444);
and UO_1511 (O_1511,N_19179,N_19439);
or UO_1512 (O_1512,N_16644,N_16380);
or UO_1513 (O_1513,N_17554,N_16057);
nor UO_1514 (O_1514,N_17560,N_16328);
nand UO_1515 (O_1515,N_19606,N_16896);
nand UO_1516 (O_1516,N_16747,N_19362);
nor UO_1517 (O_1517,N_18659,N_18806);
nand UO_1518 (O_1518,N_19705,N_17551);
nand UO_1519 (O_1519,N_17960,N_17590);
and UO_1520 (O_1520,N_16485,N_18062);
or UO_1521 (O_1521,N_19692,N_17899);
and UO_1522 (O_1522,N_18262,N_16469);
nor UO_1523 (O_1523,N_19646,N_19965);
nand UO_1524 (O_1524,N_16128,N_19714);
nor UO_1525 (O_1525,N_16049,N_19480);
or UO_1526 (O_1526,N_17613,N_18559);
or UO_1527 (O_1527,N_16283,N_18003);
and UO_1528 (O_1528,N_16818,N_16624);
and UO_1529 (O_1529,N_19952,N_18760);
xnor UO_1530 (O_1530,N_18337,N_18359);
or UO_1531 (O_1531,N_18482,N_16530);
and UO_1532 (O_1532,N_16329,N_16435);
or UO_1533 (O_1533,N_19514,N_18353);
xnor UO_1534 (O_1534,N_18564,N_19109);
or UO_1535 (O_1535,N_16826,N_18283);
nand UO_1536 (O_1536,N_19393,N_19566);
nand UO_1537 (O_1537,N_16312,N_19504);
nand UO_1538 (O_1538,N_16690,N_17331);
and UO_1539 (O_1539,N_19602,N_19576);
and UO_1540 (O_1540,N_17009,N_17478);
xor UO_1541 (O_1541,N_16721,N_18673);
nand UO_1542 (O_1542,N_16595,N_19012);
nand UO_1543 (O_1543,N_16358,N_17915);
nand UO_1544 (O_1544,N_16531,N_16012);
and UO_1545 (O_1545,N_19386,N_18314);
and UO_1546 (O_1546,N_17906,N_19118);
nor UO_1547 (O_1547,N_19779,N_17467);
or UO_1548 (O_1548,N_17996,N_17072);
xnor UO_1549 (O_1549,N_16399,N_18982);
and UO_1550 (O_1550,N_19559,N_19200);
nand UO_1551 (O_1551,N_16902,N_18773);
nand UO_1552 (O_1552,N_17922,N_16811);
or UO_1553 (O_1553,N_17603,N_17215);
nor UO_1554 (O_1554,N_19291,N_18485);
nor UO_1555 (O_1555,N_19933,N_19966);
xor UO_1556 (O_1556,N_18785,N_19667);
nor UO_1557 (O_1557,N_16275,N_17760);
nand UO_1558 (O_1558,N_17025,N_19269);
or UO_1559 (O_1559,N_17460,N_17630);
or UO_1560 (O_1560,N_19363,N_19517);
or UO_1561 (O_1561,N_18442,N_16783);
nor UO_1562 (O_1562,N_17336,N_16059);
or UO_1563 (O_1563,N_18611,N_17850);
nor UO_1564 (O_1564,N_19425,N_18308);
nand UO_1565 (O_1565,N_18244,N_18294);
nor UO_1566 (O_1566,N_18298,N_16500);
nand UO_1567 (O_1567,N_18566,N_18642);
or UO_1568 (O_1568,N_18409,N_16860);
nor UO_1569 (O_1569,N_18090,N_17646);
xnor UO_1570 (O_1570,N_18227,N_16338);
nand UO_1571 (O_1571,N_17332,N_19615);
and UO_1572 (O_1572,N_16506,N_17381);
nand UO_1573 (O_1573,N_16677,N_17231);
and UO_1574 (O_1574,N_16236,N_18292);
nor UO_1575 (O_1575,N_18161,N_16210);
nor UO_1576 (O_1576,N_17455,N_17606);
or UO_1577 (O_1577,N_18309,N_19315);
nand UO_1578 (O_1578,N_19922,N_19029);
nand UO_1579 (O_1579,N_17867,N_17994);
or UO_1580 (O_1580,N_17580,N_16237);
and UO_1581 (O_1581,N_18688,N_17027);
nand UO_1582 (O_1582,N_18408,N_19925);
or UO_1583 (O_1583,N_18826,N_16523);
and UO_1584 (O_1584,N_19795,N_16748);
nor UO_1585 (O_1585,N_16874,N_19140);
or UO_1586 (O_1586,N_19674,N_18203);
nor UO_1587 (O_1587,N_16133,N_19455);
nor UO_1588 (O_1588,N_19314,N_19958);
or UO_1589 (O_1589,N_17833,N_17728);
nand UO_1590 (O_1590,N_18838,N_19745);
or UO_1591 (O_1591,N_16161,N_18828);
and UO_1592 (O_1592,N_16393,N_17593);
and UO_1593 (O_1593,N_18226,N_16391);
nor UO_1594 (O_1594,N_17396,N_18277);
nand UO_1595 (O_1595,N_16777,N_17987);
and UO_1596 (O_1596,N_16905,N_19196);
and UO_1597 (O_1597,N_16816,N_16834);
or UO_1598 (O_1598,N_19281,N_19058);
nor UO_1599 (O_1599,N_16001,N_16078);
nor UO_1600 (O_1600,N_18033,N_17841);
nand UO_1601 (O_1601,N_19184,N_16483);
or UO_1602 (O_1602,N_17288,N_16859);
nand UO_1603 (O_1603,N_17797,N_19050);
xnor UO_1604 (O_1604,N_16750,N_16864);
nand UO_1605 (O_1605,N_19877,N_16597);
nand UO_1606 (O_1606,N_18255,N_19246);
nor UO_1607 (O_1607,N_17519,N_19697);
nor UO_1608 (O_1608,N_16796,N_17699);
and UO_1609 (O_1609,N_16986,N_18943);
nor UO_1610 (O_1610,N_19822,N_16665);
nor UO_1611 (O_1611,N_17077,N_17617);
and UO_1612 (O_1612,N_18623,N_19663);
nand UO_1613 (O_1613,N_16852,N_18338);
and UO_1614 (O_1614,N_18810,N_19824);
nor UO_1615 (O_1615,N_17388,N_17176);
or UO_1616 (O_1616,N_17605,N_18207);
nand UO_1617 (O_1617,N_19787,N_17619);
xor UO_1618 (O_1618,N_16766,N_19052);
and UO_1619 (O_1619,N_19526,N_16100);
nand UO_1620 (O_1620,N_18620,N_17071);
nor UO_1621 (O_1621,N_19749,N_19633);
nand UO_1622 (O_1622,N_19447,N_17828);
or UO_1623 (O_1623,N_16015,N_18575);
or UO_1624 (O_1624,N_17090,N_17805);
and UO_1625 (O_1625,N_18376,N_19435);
or UO_1626 (O_1626,N_16529,N_17520);
xor UO_1627 (O_1627,N_18400,N_19796);
or UO_1628 (O_1628,N_17715,N_16212);
or UO_1629 (O_1629,N_18165,N_18861);
or UO_1630 (O_1630,N_18154,N_17674);
and UO_1631 (O_1631,N_18607,N_17169);
nor UO_1632 (O_1632,N_16349,N_18516);
nand UO_1633 (O_1633,N_19243,N_18880);
nor UO_1634 (O_1634,N_19984,N_18705);
xor UO_1635 (O_1635,N_19687,N_17440);
or UO_1636 (O_1636,N_17599,N_17084);
nand UO_1637 (O_1637,N_18051,N_16123);
nor UO_1638 (O_1638,N_19427,N_17767);
nor UO_1639 (O_1639,N_19085,N_16066);
and UO_1640 (O_1640,N_17221,N_16407);
nor UO_1641 (O_1641,N_18473,N_16370);
or UO_1642 (O_1642,N_19998,N_16947);
nor UO_1643 (O_1643,N_16515,N_19320);
nor UO_1644 (O_1644,N_18649,N_16309);
nand UO_1645 (O_1645,N_16618,N_19375);
nand UO_1646 (O_1646,N_16950,N_17658);
nand UO_1647 (O_1647,N_16666,N_16084);
and UO_1648 (O_1648,N_16223,N_17449);
nand UO_1649 (O_1649,N_16940,N_18354);
or UO_1650 (O_1650,N_19884,N_18911);
and UO_1651 (O_1651,N_18518,N_18615);
nand UO_1652 (O_1652,N_17900,N_18433);
nor UO_1653 (O_1653,N_18934,N_17074);
and UO_1654 (O_1654,N_18577,N_17811);
and UO_1655 (O_1655,N_19437,N_17450);
or UO_1656 (O_1656,N_19879,N_18041);
nor UO_1657 (O_1657,N_16294,N_19006);
nand UO_1658 (O_1658,N_16375,N_18511);
or UO_1659 (O_1659,N_19217,N_17932);
xor UO_1660 (O_1660,N_16607,N_16537);
and UO_1661 (O_1661,N_18581,N_16965);
nand UO_1662 (O_1662,N_19927,N_17416);
nor UO_1663 (O_1663,N_18091,N_16474);
or UO_1664 (O_1664,N_16702,N_16053);
and UO_1665 (O_1665,N_18897,N_16111);
and UO_1666 (O_1666,N_17048,N_17535);
or UO_1667 (O_1667,N_18670,N_17538);
xnor UO_1668 (O_1668,N_17040,N_19015);
or UO_1669 (O_1669,N_17666,N_17910);
nand UO_1670 (O_1670,N_17957,N_17301);
or UO_1671 (O_1671,N_17291,N_18445);
nand UO_1672 (O_1672,N_17997,N_16148);
nand UO_1673 (O_1673,N_17781,N_17212);
nand UO_1674 (O_1674,N_19430,N_16311);
and UO_1675 (O_1675,N_16724,N_18837);
and UO_1676 (O_1676,N_17306,N_17165);
or UO_1677 (O_1677,N_17629,N_19873);
and UO_1678 (O_1678,N_18756,N_19120);
and UO_1679 (O_1679,N_17660,N_19863);
nand UO_1680 (O_1680,N_19249,N_19097);
nor UO_1681 (O_1681,N_16823,N_18915);
and UO_1682 (O_1682,N_16525,N_16895);
nor UO_1683 (O_1683,N_19757,N_16539);
and UO_1684 (O_1684,N_16667,N_17667);
xor UO_1685 (O_1685,N_19051,N_17496);
nor UO_1686 (O_1686,N_18662,N_16410);
and UO_1687 (O_1687,N_17190,N_19376);
and UO_1688 (O_1688,N_16402,N_17209);
nand UO_1689 (O_1689,N_18952,N_18045);
xnor UO_1690 (O_1690,N_17602,N_17581);
nor UO_1691 (O_1691,N_16577,N_18311);
nor UO_1692 (O_1692,N_16518,N_16849);
and UO_1693 (O_1693,N_17238,N_16196);
and UO_1694 (O_1694,N_17771,N_16687);
nand UO_1695 (O_1695,N_18622,N_17939);
nor UO_1696 (O_1696,N_18392,N_19699);
or UO_1697 (O_1697,N_17121,N_17600);
and UO_1698 (O_1698,N_16304,N_18006);
nand UO_1699 (O_1699,N_19436,N_19232);
or UO_1700 (O_1700,N_16473,N_16445);
nand UO_1701 (O_1701,N_18447,N_19856);
or UO_1702 (O_1702,N_16737,N_19766);
and UO_1703 (O_1703,N_19583,N_19683);
nor UO_1704 (O_1704,N_16043,N_18972);
nor UO_1705 (O_1705,N_19384,N_17078);
nand UO_1706 (O_1706,N_16008,N_16011);
xnor UO_1707 (O_1707,N_18082,N_17751);
or UO_1708 (O_1708,N_18980,N_19062);
or UO_1709 (O_1709,N_19875,N_19071);
nor UO_1710 (O_1710,N_18789,N_17297);
or UO_1711 (O_1711,N_16708,N_18351);
and UO_1712 (O_1712,N_17594,N_19503);
nand UO_1713 (O_1713,N_18375,N_19302);
or UO_1714 (O_1714,N_17294,N_19838);
or UO_1715 (O_1715,N_18769,N_16044);
xnor UO_1716 (O_1716,N_18396,N_17036);
nor UO_1717 (O_1717,N_17299,N_18201);
nor UO_1718 (O_1718,N_19133,N_17512);
or UO_1719 (O_1719,N_19769,N_18027);
or UO_1720 (O_1720,N_18901,N_19081);
nor UO_1721 (O_1721,N_18142,N_19188);
and UO_1722 (O_1722,N_16674,N_19840);
nand UO_1723 (O_1723,N_17205,N_16688);
and UO_1724 (O_1724,N_19931,N_16856);
nor UO_1725 (O_1725,N_18728,N_16007);
or UO_1726 (O_1726,N_19930,N_16240);
xnor UO_1727 (O_1727,N_18947,N_19664);
xor UO_1728 (O_1728,N_17640,N_19328);
and UO_1729 (O_1729,N_17831,N_18437);
nor UO_1730 (O_1730,N_19406,N_17839);
nand UO_1731 (O_1731,N_18848,N_17676);
and UO_1732 (O_1732,N_17800,N_17135);
and UO_1733 (O_1733,N_18096,N_18693);
nand UO_1734 (O_1734,N_16526,N_16713);
nor UO_1735 (O_1735,N_18427,N_17481);
or UO_1736 (O_1736,N_18199,N_19903);
xor UO_1737 (O_1737,N_18065,N_19381);
nand UO_1738 (O_1738,N_16342,N_16989);
nor UO_1739 (O_1739,N_18632,N_19900);
and UO_1740 (O_1740,N_17085,N_18493);
or UO_1741 (O_1741,N_17225,N_19367);
nor UO_1742 (O_1742,N_19231,N_16584);
and UO_1743 (O_1743,N_16779,N_16471);
nand UO_1744 (O_1744,N_16546,N_16756);
nand UO_1745 (O_1745,N_19617,N_17399);
and UO_1746 (O_1746,N_17506,N_19963);
or UO_1747 (O_1747,N_17178,N_16077);
nor UO_1748 (O_1748,N_16995,N_19165);
nor UO_1749 (O_1749,N_19885,N_16662);
nor UO_1750 (O_1750,N_18340,N_19076);
and UO_1751 (O_1751,N_19276,N_17845);
nor UO_1752 (O_1752,N_17122,N_17586);
nand UO_1753 (O_1753,N_18029,N_16442);
or UO_1754 (O_1754,N_17775,N_16588);
nand UO_1755 (O_1755,N_16652,N_18885);
nand UO_1756 (O_1756,N_16675,N_16480);
and UO_1757 (O_1757,N_16141,N_18265);
nor UO_1758 (O_1758,N_19912,N_16048);
nor UO_1759 (O_1759,N_19814,N_16006);
nand UO_1760 (O_1760,N_19703,N_19220);
nor UO_1761 (O_1761,N_18804,N_19089);
and UO_1762 (O_1762,N_17174,N_19034);
or UO_1763 (O_1763,N_19407,N_17223);
and UO_1764 (O_1764,N_17592,N_19619);
xnor UO_1765 (O_1765,N_17533,N_19223);
xor UO_1766 (O_1766,N_19205,N_18991);
nand UO_1767 (O_1767,N_19255,N_18964);
and UO_1768 (O_1768,N_19818,N_16730);
xor UO_1769 (O_1769,N_19056,N_19322);
nor UO_1770 (O_1770,N_19419,N_18004);
or UO_1771 (O_1771,N_19696,N_19180);
and UO_1772 (O_1772,N_16901,N_18281);
or UO_1773 (O_1773,N_19839,N_16802);
xnor UO_1774 (O_1774,N_17877,N_16956);
or UO_1775 (O_1775,N_17232,N_19198);
and UO_1776 (O_1776,N_16980,N_19914);
nor UO_1777 (O_1777,N_17179,N_18108);
nor UO_1778 (O_1778,N_16272,N_19072);
and UO_1779 (O_1779,N_16289,N_19535);
nor UO_1780 (O_1780,N_19904,N_17584);
nand UO_1781 (O_1781,N_19286,N_19613);
or UO_1782 (O_1782,N_19024,N_18849);
or UO_1783 (O_1783,N_18744,N_16022);
or UO_1784 (O_1784,N_19112,N_18950);
and UO_1785 (O_1785,N_18386,N_17200);
or UO_1786 (O_1786,N_19756,N_17260);
nand UO_1787 (O_1787,N_19247,N_16767);
xnor UO_1788 (O_1788,N_17935,N_19772);
and UO_1789 (O_1789,N_16893,N_17337);
or UO_1790 (O_1790,N_16122,N_17763);
and UO_1791 (O_1791,N_18477,N_16912);
or UO_1792 (O_1792,N_19785,N_17098);
nor UO_1793 (O_1793,N_16993,N_19498);
and UO_1794 (O_1794,N_17866,N_19222);
or UO_1795 (O_1795,N_19306,N_19919);
or UO_1796 (O_1796,N_19876,N_17070);
nand UO_1797 (O_1797,N_18987,N_16336);
nand UO_1798 (O_1798,N_18505,N_19636);
or UO_1799 (O_1799,N_18094,N_19874);
and UO_1800 (O_1800,N_17364,N_16876);
and UO_1801 (O_1801,N_17645,N_16408);
and UO_1802 (O_1802,N_16472,N_18494);
nand UO_1803 (O_1803,N_17258,N_16924);
xnor UO_1804 (O_1804,N_16798,N_19069);
nor UO_1805 (O_1805,N_18971,N_17647);
nand UO_1806 (O_1806,N_16467,N_17672);
nand UO_1807 (O_1807,N_18136,N_16897);
and UO_1808 (O_1808,N_18302,N_18145);
and UO_1809 (O_1809,N_18325,N_16207);
xor UO_1810 (O_1810,N_18825,N_16353);
or UO_1811 (O_1811,N_18140,N_16573);
and UO_1812 (O_1812,N_18236,N_19854);
nor UO_1813 (O_1813,N_19125,N_16579);
and UO_1814 (O_1814,N_16331,N_16050);
or UO_1815 (O_1815,N_17879,N_16592);
nand UO_1816 (O_1816,N_16951,N_17884);
nand UO_1817 (O_1817,N_19383,N_19542);
and UO_1818 (O_1818,N_19092,N_16318);
or UO_1819 (O_1819,N_18906,N_18060);
nand UO_1820 (O_1820,N_18631,N_19640);
nor UO_1821 (O_1821,N_16367,N_17796);
or UO_1822 (O_1822,N_17240,N_18543);
nand UO_1823 (O_1823,N_17890,N_16846);
nor UO_1824 (O_1824,N_18675,N_18052);
nor UO_1825 (O_1825,N_17233,N_19485);
nand UO_1826 (O_1826,N_18044,N_16971);
nor UO_1827 (O_1827,N_17791,N_17138);
nand UO_1828 (O_1828,N_17188,N_17480);
nand UO_1829 (O_1829,N_16815,N_19605);
nand UO_1830 (O_1830,N_17919,N_16252);
or UO_1831 (O_1831,N_18101,N_16020);
nand UO_1832 (O_1832,N_18461,N_19429);
nand UO_1833 (O_1833,N_16280,N_18155);
or UO_1834 (O_1834,N_17018,N_19446);
nand UO_1835 (O_1835,N_17172,N_16845);
and UO_1836 (O_1836,N_16109,N_17418);
nor UO_1837 (O_1837,N_16200,N_19622);
nand UO_1838 (O_1838,N_18525,N_18995);
or UO_1839 (O_1839,N_17013,N_16496);
and UO_1840 (O_1840,N_18889,N_19343);
nor UO_1841 (O_1841,N_17022,N_19864);
nor UO_1842 (O_1842,N_16235,N_16959);
or UO_1843 (O_1843,N_16831,N_18238);
nand UO_1844 (O_1844,N_17762,N_19686);
or UO_1845 (O_1845,N_16324,N_16839);
nor UO_1846 (O_1846,N_16800,N_16918);
and UO_1847 (O_1847,N_18188,N_17392);
or UO_1848 (O_1848,N_19221,N_17964);
nor UO_1849 (O_1849,N_17566,N_17848);
nor UO_1850 (O_1850,N_17849,N_18185);
xnor UO_1851 (O_1851,N_17934,N_18882);
or UO_1852 (O_1852,N_17377,N_18446);
xor UO_1853 (O_1853,N_18183,N_17819);
and UO_1854 (O_1854,N_16789,N_17705);
nand UO_1855 (O_1855,N_19008,N_19789);
nand UO_1856 (O_1856,N_17753,N_16051);
and UO_1857 (O_1857,N_17216,N_19552);
nand UO_1858 (O_1858,N_18986,N_19924);
nor UO_1859 (O_1859,N_16697,N_17920);
or UO_1860 (O_1860,N_19722,N_19515);
nand UO_1861 (O_1861,N_16023,N_18997);
nand UO_1862 (O_1862,N_18092,N_17693);
nand UO_1863 (O_1863,N_18970,N_17486);
and UO_1864 (O_1864,N_19939,N_19068);
nor UO_1865 (O_1865,N_16854,N_16862);
nand UO_1866 (O_1866,N_19233,N_18764);
and UO_1867 (O_1867,N_17214,N_16964);
nor UO_1868 (O_1868,N_17655,N_16033);
nor UO_1869 (O_1869,N_16316,N_19928);
or UO_1870 (O_1870,N_16482,N_18522);
and UO_1871 (O_1871,N_18617,N_19797);
nand UO_1872 (O_1872,N_18599,N_19653);
nand UO_1873 (O_1873,N_16460,N_17508);
and UO_1874 (O_1874,N_19589,N_18315);
nand UO_1875 (O_1875,N_18790,N_17430);
or UO_1876 (O_1876,N_18331,N_16121);
and UO_1877 (O_1877,N_16352,N_18303);
and UO_1878 (O_1878,N_19536,N_19881);
and UO_1879 (O_1879,N_18706,N_16150);
and UO_1880 (O_1880,N_19828,N_16170);
nor UO_1881 (O_1881,N_19878,N_18871);
nand UO_1882 (O_1882,N_18050,N_19759);
nor UO_1883 (O_1883,N_16390,N_16130);
and UO_1884 (O_1884,N_18391,N_18272);
nand UO_1885 (O_1885,N_17323,N_18177);
and UO_1886 (O_1886,N_18440,N_16253);
nand UO_1887 (O_1887,N_18260,N_19278);
and UO_1888 (O_1888,N_18164,N_16206);
or UO_1889 (O_1889,N_19708,N_17391);
or UO_1890 (O_1890,N_16542,N_16883);
and UO_1891 (O_1891,N_19116,N_16371);
nand UO_1892 (O_1892,N_18989,N_17446);
nand UO_1893 (O_1893,N_19434,N_18444);
nand UO_1894 (O_1894,N_19518,N_17893);
xnor UO_1895 (O_1895,N_18689,N_17197);
xor UO_1896 (O_1896,N_17976,N_17393);
and UO_1897 (O_1897,N_19823,N_19786);
nand UO_1898 (O_1898,N_17680,N_16631);
xor UO_1899 (O_1899,N_18618,N_18570);
nand UO_1900 (O_1900,N_16287,N_19074);
and UO_1901 (O_1901,N_16203,N_16278);
nor UO_1902 (O_1902,N_16685,N_17325);
and UO_1903 (O_1903,N_17042,N_16549);
or UO_1904 (O_1904,N_17537,N_17164);
nand UO_1905 (O_1905,N_18126,N_18928);
nand UO_1906 (O_1906,N_19374,N_16245);
nor UO_1907 (O_1907,N_18258,N_18499);
nor UO_1908 (O_1908,N_16605,N_19026);
nor UO_1909 (O_1909,N_18665,N_16432);
xor UO_1910 (O_1910,N_17308,N_19702);
nor UO_1911 (O_1911,N_19250,N_16083);
and UO_1912 (O_1912,N_17079,N_18018);
and UO_1913 (O_1913,N_16890,N_16392);
nand UO_1914 (O_1914,N_18235,N_16149);
or UO_1915 (O_1915,N_17140,N_17729);
nor UO_1916 (O_1916,N_17861,N_16292);
and UO_1917 (O_1917,N_16095,N_19293);
nor UO_1918 (O_1918,N_17057,N_16731);
or UO_1919 (O_1919,N_17134,N_18067);
nor UO_1920 (O_1920,N_17243,N_19820);
or UO_1921 (O_1921,N_18163,N_19677);
xor UO_1922 (O_1922,N_18549,N_18466);
nand UO_1923 (O_1923,N_16863,N_16183);
xor UO_1924 (O_1924,N_16118,N_17941);
nand UO_1925 (O_1925,N_19811,N_17362);
and UO_1926 (O_1926,N_19462,N_17894);
and UO_1927 (O_1927,N_17803,N_18358);
and UO_1928 (O_1928,N_16869,N_17289);
xor UO_1929 (O_1929,N_19156,N_16642);
or UO_1930 (O_1930,N_19790,N_19193);
nor UO_1931 (O_1931,N_16487,N_17104);
and UO_1932 (O_1932,N_18819,N_18106);
nor UO_1933 (O_1933,N_17335,N_17202);
or UO_1934 (O_1934,N_16958,N_18562);
nor UO_1935 (O_1935,N_19997,N_17066);
xor UO_1936 (O_1936,N_19737,N_16242);
nand UO_1937 (O_1937,N_19763,N_16921);
nand UO_1938 (O_1938,N_18168,N_17067);
or UO_1939 (O_1939,N_16615,N_17526);
and UO_1940 (O_1940,N_16946,N_19625);
xnor UO_1941 (O_1941,N_19821,N_16085);
and UO_1942 (O_1942,N_17157,N_16061);
and UO_1943 (O_1943,N_16810,N_18474);
nor UO_1944 (O_1944,N_17664,N_19798);
or UO_1945 (O_1945,N_17880,N_19207);
nor UO_1946 (O_1946,N_18245,N_17142);
and UO_1947 (O_1947,N_16732,N_17870);
and UO_1948 (O_1948,N_17546,N_16425);
nor UO_1949 (O_1949,N_16550,N_17568);
nor UO_1950 (O_1950,N_16265,N_18909);
xnor UO_1951 (O_1951,N_19543,N_19695);
or UO_1952 (O_1952,N_18874,N_16151);
nand UO_1953 (O_1953,N_17415,N_19475);
xnor UO_1954 (O_1954,N_16832,N_18976);
or UO_1955 (O_1955,N_19516,N_18754);
or UO_1956 (O_1956,N_16291,N_17823);
and UO_1957 (O_1957,N_19025,N_17410);
or UO_1958 (O_1958,N_19146,N_17945);
and UO_1959 (O_1959,N_17422,N_17659);
nor UO_1960 (O_1960,N_19629,N_19800);
nor UO_1961 (O_1961,N_18198,N_16999);
nor UO_1962 (O_1962,N_18098,N_16191);
nor UO_1963 (O_1963,N_16147,N_19588);
nand UO_1964 (O_1964,N_17812,N_17352);
and UO_1965 (O_1965,N_17611,N_18854);
or UO_1966 (O_1966,N_17493,N_16865);
nor UO_1967 (O_1967,N_19957,N_17356);
xnor UO_1968 (O_1968,N_18451,N_18723);
or UO_1969 (O_1969,N_19610,N_19308);
or UO_1970 (O_1970,N_19668,N_16126);
nor UO_1971 (O_1971,N_18985,N_18729);
nor UO_1972 (O_1972,N_16828,N_16419);
nand UO_1973 (O_1973,N_18866,N_16933);
xnor UO_1974 (O_1974,N_17973,N_17550);
or UO_1975 (O_1975,N_18946,N_18048);
or UO_1976 (O_1976,N_18443,N_18047);
xnor UO_1977 (O_1977,N_17741,N_16858);
nor UO_1978 (O_1978,N_17229,N_17882);
or UO_1979 (O_1979,N_16617,N_19541);
or UO_1980 (O_1980,N_16705,N_18844);
xor UO_1981 (O_1981,N_18858,N_19621);
nand UO_1982 (O_1982,N_18017,N_19445);
xor UO_1983 (O_1983,N_17447,N_17777);
xnor UO_1984 (O_1984,N_18234,N_17914);
nand UO_1985 (O_1985,N_18753,N_17824);
nand UO_1986 (O_1986,N_16514,N_19845);
and UO_1987 (O_1987,N_16468,N_16263);
nand UO_1988 (O_1988,N_17543,N_18545);
nand UO_1989 (O_1989,N_19107,N_19577);
xnor UO_1990 (O_1990,N_19280,N_18345);
xor UO_1991 (O_1991,N_16694,N_16585);
xnor UO_1992 (O_1992,N_17830,N_16251);
or UO_1993 (O_1993,N_19279,N_17736);
nor UO_1994 (O_1994,N_16703,N_18626);
nand UO_1995 (O_1995,N_16879,N_18480);
or UO_1996 (O_1996,N_17686,N_17234);
and UO_1997 (O_1997,N_16102,N_17448);
and UO_1998 (O_1998,N_18935,N_16763);
and UO_1999 (O_1999,N_17793,N_17183);
or UO_2000 (O_2000,N_17823,N_18342);
and UO_2001 (O_2001,N_17701,N_17259);
and UO_2002 (O_2002,N_18031,N_19435);
or UO_2003 (O_2003,N_17448,N_18676);
nor UO_2004 (O_2004,N_17835,N_19908);
xor UO_2005 (O_2005,N_19514,N_18432);
xor UO_2006 (O_2006,N_18744,N_17741);
or UO_2007 (O_2007,N_17043,N_18784);
nor UO_2008 (O_2008,N_19648,N_18876);
xor UO_2009 (O_2009,N_19806,N_17627);
nor UO_2010 (O_2010,N_17623,N_18971);
or UO_2011 (O_2011,N_17793,N_19968);
nand UO_2012 (O_2012,N_19217,N_16347);
nor UO_2013 (O_2013,N_18866,N_17087);
and UO_2014 (O_2014,N_16561,N_18502);
or UO_2015 (O_2015,N_16357,N_19755);
nand UO_2016 (O_2016,N_19070,N_18971);
nand UO_2017 (O_2017,N_18406,N_16481);
xnor UO_2018 (O_2018,N_19225,N_18346);
or UO_2019 (O_2019,N_17828,N_16485);
nor UO_2020 (O_2020,N_17589,N_17468);
and UO_2021 (O_2021,N_17483,N_19157);
nand UO_2022 (O_2022,N_17000,N_18396);
or UO_2023 (O_2023,N_18544,N_16710);
nand UO_2024 (O_2024,N_16838,N_19111);
and UO_2025 (O_2025,N_18596,N_16702);
and UO_2026 (O_2026,N_18213,N_19968);
nand UO_2027 (O_2027,N_19445,N_18385);
nand UO_2028 (O_2028,N_17241,N_16244);
or UO_2029 (O_2029,N_19884,N_16890);
nor UO_2030 (O_2030,N_19671,N_19405);
or UO_2031 (O_2031,N_16216,N_19365);
nand UO_2032 (O_2032,N_16520,N_18424);
and UO_2033 (O_2033,N_18833,N_16775);
xor UO_2034 (O_2034,N_19440,N_18399);
nand UO_2035 (O_2035,N_17189,N_19764);
nand UO_2036 (O_2036,N_17354,N_18564);
and UO_2037 (O_2037,N_19746,N_19429);
nor UO_2038 (O_2038,N_18013,N_17958);
or UO_2039 (O_2039,N_19857,N_19985);
nand UO_2040 (O_2040,N_17935,N_18522);
nor UO_2041 (O_2041,N_19980,N_18562);
and UO_2042 (O_2042,N_16290,N_19341);
and UO_2043 (O_2043,N_19168,N_18675);
or UO_2044 (O_2044,N_16002,N_17624);
nor UO_2045 (O_2045,N_19783,N_16805);
or UO_2046 (O_2046,N_17851,N_16894);
nand UO_2047 (O_2047,N_18154,N_17692);
or UO_2048 (O_2048,N_18735,N_16011);
nor UO_2049 (O_2049,N_16277,N_17435);
and UO_2050 (O_2050,N_19677,N_17677);
and UO_2051 (O_2051,N_18622,N_19289);
nor UO_2052 (O_2052,N_16923,N_19018);
nor UO_2053 (O_2053,N_19016,N_18194);
nand UO_2054 (O_2054,N_17585,N_18710);
nor UO_2055 (O_2055,N_16154,N_18143);
nand UO_2056 (O_2056,N_19817,N_19788);
and UO_2057 (O_2057,N_19104,N_19624);
or UO_2058 (O_2058,N_19081,N_19477);
xor UO_2059 (O_2059,N_17453,N_18400);
or UO_2060 (O_2060,N_18313,N_19834);
nor UO_2061 (O_2061,N_18853,N_17081);
or UO_2062 (O_2062,N_17591,N_18707);
or UO_2063 (O_2063,N_18566,N_16203);
nor UO_2064 (O_2064,N_18662,N_16831);
nor UO_2065 (O_2065,N_17234,N_19618);
or UO_2066 (O_2066,N_16300,N_16281);
xnor UO_2067 (O_2067,N_16369,N_16750);
xor UO_2068 (O_2068,N_17891,N_18503);
nor UO_2069 (O_2069,N_16052,N_19741);
or UO_2070 (O_2070,N_16161,N_18899);
nand UO_2071 (O_2071,N_19436,N_16911);
nand UO_2072 (O_2072,N_19170,N_17720);
nand UO_2073 (O_2073,N_17459,N_19609);
or UO_2074 (O_2074,N_18151,N_16150);
or UO_2075 (O_2075,N_19754,N_18464);
or UO_2076 (O_2076,N_18171,N_18122);
or UO_2077 (O_2077,N_16547,N_19667);
nand UO_2078 (O_2078,N_17642,N_17187);
xor UO_2079 (O_2079,N_16011,N_19451);
nand UO_2080 (O_2080,N_19364,N_17368);
or UO_2081 (O_2081,N_18109,N_18938);
nand UO_2082 (O_2082,N_19128,N_17297);
and UO_2083 (O_2083,N_19136,N_18956);
nor UO_2084 (O_2084,N_17847,N_17665);
nor UO_2085 (O_2085,N_16421,N_18132);
nand UO_2086 (O_2086,N_17007,N_17061);
nor UO_2087 (O_2087,N_19763,N_16758);
nand UO_2088 (O_2088,N_16217,N_19575);
nand UO_2089 (O_2089,N_16422,N_16647);
xor UO_2090 (O_2090,N_19397,N_16175);
or UO_2091 (O_2091,N_18502,N_19315);
and UO_2092 (O_2092,N_16859,N_17055);
or UO_2093 (O_2093,N_19699,N_17951);
nand UO_2094 (O_2094,N_16897,N_16755);
xor UO_2095 (O_2095,N_16626,N_17806);
nor UO_2096 (O_2096,N_18144,N_19878);
nand UO_2097 (O_2097,N_17385,N_17524);
nand UO_2098 (O_2098,N_16748,N_16283);
or UO_2099 (O_2099,N_17138,N_17599);
or UO_2100 (O_2100,N_17304,N_19727);
nor UO_2101 (O_2101,N_16946,N_17341);
and UO_2102 (O_2102,N_16818,N_18757);
xor UO_2103 (O_2103,N_18934,N_16820);
nor UO_2104 (O_2104,N_16151,N_16786);
and UO_2105 (O_2105,N_16204,N_19988);
or UO_2106 (O_2106,N_19216,N_17917);
or UO_2107 (O_2107,N_16501,N_19571);
xor UO_2108 (O_2108,N_19063,N_16696);
nor UO_2109 (O_2109,N_18386,N_17792);
and UO_2110 (O_2110,N_19185,N_18323);
and UO_2111 (O_2111,N_17931,N_19682);
and UO_2112 (O_2112,N_17077,N_17699);
nor UO_2113 (O_2113,N_17167,N_18455);
nor UO_2114 (O_2114,N_16657,N_19056);
and UO_2115 (O_2115,N_19329,N_19911);
nand UO_2116 (O_2116,N_19594,N_18306);
or UO_2117 (O_2117,N_17172,N_16912);
nor UO_2118 (O_2118,N_16158,N_16921);
nand UO_2119 (O_2119,N_18692,N_16950);
or UO_2120 (O_2120,N_18778,N_19416);
or UO_2121 (O_2121,N_16141,N_18490);
or UO_2122 (O_2122,N_16658,N_19277);
xnor UO_2123 (O_2123,N_16005,N_17496);
nand UO_2124 (O_2124,N_19634,N_19627);
and UO_2125 (O_2125,N_18890,N_18320);
nand UO_2126 (O_2126,N_16357,N_19124);
nand UO_2127 (O_2127,N_19657,N_17001);
or UO_2128 (O_2128,N_19642,N_17101);
nor UO_2129 (O_2129,N_17377,N_17857);
nor UO_2130 (O_2130,N_19116,N_19224);
and UO_2131 (O_2131,N_17468,N_18682);
or UO_2132 (O_2132,N_18392,N_19272);
and UO_2133 (O_2133,N_16616,N_17984);
xnor UO_2134 (O_2134,N_18868,N_17357);
or UO_2135 (O_2135,N_19109,N_16745);
or UO_2136 (O_2136,N_19630,N_19194);
and UO_2137 (O_2137,N_18811,N_17716);
or UO_2138 (O_2138,N_17501,N_16126);
nand UO_2139 (O_2139,N_18216,N_16462);
or UO_2140 (O_2140,N_16731,N_19322);
nor UO_2141 (O_2141,N_18182,N_18579);
xnor UO_2142 (O_2142,N_18214,N_16833);
and UO_2143 (O_2143,N_18678,N_18498);
nor UO_2144 (O_2144,N_19140,N_16753);
nand UO_2145 (O_2145,N_19070,N_17856);
nand UO_2146 (O_2146,N_18309,N_18948);
nand UO_2147 (O_2147,N_16709,N_17611);
nand UO_2148 (O_2148,N_17985,N_18700);
or UO_2149 (O_2149,N_17358,N_17117);
and UO_2150 (O_2150,N_16860,N_18413);
nand UO_2151 (O_2151,N_18954,N_17902);
and UO_2152 (O_2152,N_18925,N_18448);
and UO_2153 (O_2153,N_16595,N_16713);
and UO_2154 (O_2154,N_18812,N_18749);
or UO_2155 (O_2155,N_17704,N_16520);
nand UO_2156 (O_2156,N_17957,N_19980);
xnor UO_2157 (O_2157,N_16545,N_17432);
nor UO_2158 (O_2158,N_19727,N_16444);
or UO_2159 (O_2159,N_19529,N_18815);
or UO_2160 (O_2160,N_17966,N_16693);
or UO_2161 (O_2161,N_19758,N_19149);
xor UO_2162 (O_2162,N_19302,N_16101);
nor UO_2163 (O_2163,N_18150,N_17207);
nand UO_2164 (O_2164,N_16640,N_17022);
nor UO_2165 (O_2165,N_19495,N_17880);
or UO_2166 (O_2166,N_18397,N_19657);
or UO_2167 (O_2167,N_17499,N_17172);
and UO_2168 (O_2168,N_17490,N_17200);
and UO_2169 (O_2169,N_17852,N_19569);
and UO_2170 (O_2170,N_17660,N_16817);
or UO_2171 (O_2171,N_19747,N_18727);
and UO_2172 (O_2172,N_19741,N_18388);
or UO_2173 (O_2173,N_16097,N_17367);
nor UO_2174 (O_2174,N_19252,N_16062);
or UO_2175 (O_2175,N_17115,N_17783);
nand UO_2176 (O_2176,N_19251,N_19524);
nor UO_2177 (O_2177,N_19622,N_17305);
or UO_2178 (O_2178,N_19834,N_17026);
xnor UO_2179 (O_2179,N_17634,N_16639);
and UO_2180 (O_2180,N_19840,N_16489);
or UO_2181 (O_2181,N_17866,N_18271);
xor UO_2182 (O_2182,N_17984,N_18476);
or UO_2183 (O_2183,N_16685,N_17805);
xnor UO_2184 (O_2184,N_16609,N_17562);
or UO_2185 (O_2185,N_17809,N_19410);
and UO_2186 (O_2186,N_19252,N_16918);
nor UO_2187 (O_2187,N_16177,N_17776);
and UO_2188 (O_2188,N_19387,N_18231);
or UO_2189 (O_2189,N_17837,N_17066);
or UO_2190 (O_2190,N_18526,N_19358);
nand UO_2191 (O_2191,N_16021,N_18880);
nor UO_2192 (O_2192,N_19517,N_17679);
and UO_2193 (O_2193,N_17835,N_16750);
nor UO_2194 (O_2194,N_16043,N_16513);
and UO_2195 (O_2195,N_19038,N_16347);
or UO_2196 (O_2196,N_16744,N_16481);
or UO_2197 (O_2197,N_18687,N_17336);
or UO_2198 (O_2198,N_17322,N_16992);
nand UO_2199 (O_2199,N_18238,N_17647);
nor UO_2200 (O_2200,N_19689,N_18447);
or UO_2201 (O_2201,N_16224,N_19281);
nor UO_2202 (O_2202,N_18309,N_18881);
or UO_2203 (O_2203,N_17792,N_16434);
nor UO_2204 (O_2204,N_16980,N_19704);
nor UO_2205 (O_2205,N_19168,N_16304);
or UO_2206 (O_2206,N_17845,N_17851);
nand UO_2207 (O_2207,N_19143,N_19430);
nor UO_2208 (O_2208,N_19349,N_17049);
and UO_2209 (O_2209,N_18883,N_18903);
nand UO_2210 (O_2210,N_19147,N_16416);
nor UO_2211 (O_2211,N_19421,N_19826);
and UO_2212 (O_2212,N_17999,N_19506);
nor UO_2213 (O_2213,N_18992,N_19144);
and UO_2214 (O_2214,N_17368,N_18407);
or UO_2215 (O_2215,N_18138,N_17780);
nand UO_2216 (O_2216,N_16247,N_19711);
nor UO_2217 (O_2217,N_16860,N_19187);
and UO_2218 (O_2218,N_18990,N_19025);
and UO_2219 (O_2219,N_16150,N_16473);
or UO_2220 (O_2220,N_19445,N_18329);
and UO_2221 (O_2221,N_18547,N_16547);
xor UO_2222 (O_2222,N_17583,N_19011);
xor UO_2223 (O_2223,N_16001,N_19728);
or UO_2224 (O_2224,N_17560,N_17361);
or UO_2225 (O_2225,N_16953,N_19517);
or UO_2226 (O_2226,N_17841,N_19613);
or UO_2227 (O_2227,N_18849,N_18553);
or UO_2228 (O_2228,N_17754,N_19520);
nand UO_2229 (O_2229,N_17948,N_18092);
or UO_2230 (O_2230,N_17392,N_18618);
nand UO_2231 (O_2231,N_18405,N_16619);
and UO_2232 (O_2232,N_16239,N_18123);
nor UO_2233 (O_2233,N_16165,N_18735);
xnor UO_2234 (O_2234,N_19067,N_19243);
and UO_2235 (O_2235,N_17188,N_17031);
nor UO_2236 (O_2236,N_19393,N_17313);
nand UO_2237 (O_2237,N_16564,N_19886);
or UO_2238 (O_2238,N_16515,N_19359);
or UO_2239 (O_2239,N_18952,N_18685);
or UO_2240 (O_2240,N_19275,N_19935);
nor UO_2241 (O_2241,N_16099,N_16010);
and UO_2242 (O_2242,N_17720,N_17016);
nand UO_2243 (O_2243,N_17905,N_16797);
or UO_2244 (O_2244,N_17177,N_16429);
nand UO_2245 (O_2245,N_17457,N_18152);
xnor UO_2246 (O_2246,N_19854,N_16324);
or UO_2247 (O_2247,N_16459,N_16580);
or UO_2248 (O_2248,N_18508,N_19233);
nor UO_2249 (O_2249,N_17149,N_17666);
nand UO_2250 (O_2250,N_19895,N_17584);
or UO_2251 (O_2251,N_17550,N_16853);
nand UO_2252 (O_2252,N_16762,N_19331);
and UO_2253 (O_2253,N_17286,N_16031);
and UO_2254 (O_2254,N_18646,N_16491);
nand UO_2255 (O_2255,N_18442,N_17008);
nand UO_2256 (O_2256,N_19273,N_16870);
nand UO_2257 (O_2257,N_16756,N_18463);
and UO_2258 (O_2258,N_19397,N_17316);
nand UO_2259 (O_2259,N_16576,N_19470);
xor UO_2260 (O_2260,N_16519,N_19389);
or UO_2261 (O_2261,N_17379,N_19803);
and UO_2262 (O_2262,N_19604,N_16042);
nor UO_2263 (O_2263,N_16915,N_16179);
xor UO_2264 (O_2264,N_17033,N_18036);
nand UO_2265 (O_2265,N_17191,N_18274);
xor UO_2266 (O_2266,N_17224,N_17803);
or UO_2267 (O_2267,N_16324,N_17027);
nor UO_2268 (O_2268,N_17681,N_18695);
nor UO_2269 (O_2269,N_16392,N_18244);
xor UO_2270 (O_2270,N_17189,N_17952);
nor UO_2271 (O_2271,N_18481,N_18429);
and UO_2272 (O_2272,N_19424,N_18012);
nor UO_2273 (O_2273,N_19102,N_16024);
nand UO_2274 (O_2274,N_16950,N_19328);
nand UO_2275 (O_2275,N_18575,N_18847);
nor UO_2276 (O_2276,N_19702,N_18139);
nor UO_2277 (O_2277,N_17023,N_19262);
or UO_2278 (O_2278,N_17200,N_16752);
and UO_2279 (O_2279,N_16599,N_19818);
and UO_2280 (O_2280,N_18615,N_16772);
nand UO_2281 (O_2281,N_18830,N_17447);
nand UO_2282 (O_2282,N_16295,N_16305);
and UO_2283 (O_2283,N_16364,N_18347);
xnor UO_2284 (O_2284,N_19759,N_18691);
nor UO_2285 (O_2285,N_18058,N_19452);
and UO_2286 (O_2286,N_18739,N_17956);
or UO_2287 (O_2287,N_19510,N_18264);
or UO_2288 (O_2288,N_19015,N_17777);
and UO_2289 (O_2289,N_17700,N_16559);
nor UO_2290 (O_2290,N_17362,N_19377);
or UO_2291 (O_2291,N_19296,N_19942);
or UO_2292 (O_2292,N_17982,N_16216);
or UO_2293 (O_2293,N_16492,N_17723);
and UO_2294 (O_2294,N_16286,N_19879);
or UO_2295 (O_2295,N_19572,N_16739);
nor UO_2296 (O_2296,N_17226,N_17474);
and UO_2297 (O_2297,N_17981,N_16735);
or UO_2298 (O_2298,N_17770,N_16818);
nand UO_2299 (O_2299,N_19055,N_19824);
nand UO_2300 (O_2300,N_17071,N_18636);
and UO_2301 (O_2301,N_18658,N_19400);
and UO_2302 (O_2302,N_17239,N_16734);
and UO_2303 (O_2303,N_17780,N_17383);
nor UO_2304 (O_2304,N_19385,N_17895);
nand UO_2305 (O_2305,N_19222,N_19823);
and UO_2306 (O_2306,N_19754,N_18340);
and UO_2307 (O_2307,N_17935,N_16202);
and UO_2308 (O_2308,N_19046,N_17415);
and UO_2309 (O_2309,N_19241,N_19944);
or UO_2310 (O_2310,N_17275,N_19155);
nor UO_2311 (O_2311,N_19549,N_17525);
nand UO_2312 (O_2312,N_18526,N_19612);
xnor UO_2313 (O_2313,N_19650,N_17282);
xor UO_2314 (O_2314,N_17705,N_18544);
xor UO_2315 (O_2315,N_17017,N_17426);
or UO_2316 (O_2316,N_19235,N_18824);
nor UO_2317 (O_2317,N_18399,N_19694);
and UO_2318 (O_2318,N_19135,N_18249);
or UO_2319 (O_2319,N_19290,N_16884);
nor UO_2320 (O_2320,N_17942,N_19434);
nand UO_2321 (O_2321,N_18010,N_16252);
nand UO_2322 (O_2322,N_18428,N_17904);
or UO_2323 (O_2323,N_17688,N_17935);
and UO_2324 (O_2324,N_18640,N_19233);
and UO_2325 (O_2325,N_17620,N_18693);
and UO_2326 (O_2326,N_16726,N_16496);
or UO_2327 (O_2327,N_19899,N_19993);
nor UO_2328 (O_2328,N_19178,N_19071);
nand UO_2329 (O_2329,N_16436,N_19046);
nor UO_2330 (O_2330,N_17513,N_18387);
and UO_2331 (O_2331,N_19322,N_16263);
xnor UO_2332 (O_2332,N_18833,N_17489);
nor UO_2333 (O_2333,N_16943,N_18456);
nand UO_2334 (O_2334,N_16196,N_18483);
or UO_2335 (O_2335,N_19227,N_18588);
nor UO_2336 (O_2336,N_18244,N_16790);
or UO_2337 (O_2337,N_16014,N_18435);
nand UO_2338 (O_2338,N_19228,N_16666);
or UO_2339 (O_2339,N_17029,N_17503);
nor UO_2340 (O_2340,N_17017,N_18285);
nor UO_2341 (O_2341,N_17258,N_19767);
xor UO_2342 (O_2342,N_16663,N_18895);
nor UO_2343 (O_2343,N_16288,N_16548);
nand UO_2344 (O_2344,N_18803,N_18072);
nor UO_2345 (O_2345,N_18147,N_18626);
or UO_2346 (O_2346,N_17889,N_17298);
nor UO_2347 (O_2347,N_18190,N_17163);
nand UO_2348 (O_2348,N_18430,N_16984);
nand UO_2349 (O_2349,N_17794,N_19226);
or UO_2350 (O_2350,N_16174,N_18893);
nor UO_2351 (O_2351,N_16431,N_19547);
and UO_2352 (O_2352,N_18276,N_17339);
nand UO_2353 (O_2353,N_17192,N_18057);
nand UO_2354 (O_2354,N_19963,N_16178);
nor UO_2355 (O_2355,N_16431,N_19916);
nor UO_2356 (O_2356,N_16742,N_17500);
or UO_2357 (O_2357,N_17251,N_17470);
xor UO_2358 (O_2358,N_16784,N_16555);
and UO_2359 (O_2359,N_16469,N_17887);
nor UO_2360 (O_2360,N_19665,N_17500);
nor UO_2361 (O_2361,N_17015,N_17027);
xor UO_2362 (O_2362,N_19292,N_18593);
nand UO_2363 (O_2363,N_19046,N_16467);
nor UO_2364 (O_2364,N_19266,N_16809);
and UO_2365 (O_2365,N_19412,N_17604);
or UO_2366 (O_2366,N_16800,N_16665);
or UO_2367 (O_2367,N_19158,N_18046);
xor UO_2368 (O_2368,N_18709,N_18785);
nor UO_2369 (O_2369,N_18843,N_17015);
xor UO_2370 (O_2370,N_18211,N_19371);
or UO_2371 (O_2371,N_19011,N_18641);
nor UO_2372 (O_2372,N_19646,N_18172);
or UO_2373 (O_2373,N_19536,N_16372);
or UO_2374 (O_2374,N_19048,N_16905);
nand UO_2375 (O_2375,N_19266,N_16400);
nor UO_2376 (O_2376,N_18103,N_19714);
nor UO_2377 (O_2377,N_19642,N_18746);
and UO_2378 (O_2378,N_16754,N_17532);
and UO_2379 (O_2379,N_17935,N_19390);
and UO_2380 (O_2380,N_17089,N_18834);
nor UO_2381 (O_2381,N_19706,N_19913);
xnor UO_2382 (O_2382,N_17959,N_19954);
or UO_2383 (O_2383,N_19388,N_16169);
and UO_2384 (O_2384,N_16511,N_18932);
or UO_2385 (O_2385,N_18113,N_17961);
nor UO_2386 (O_2386,N_19647,N_17872);
nor UO_2387 (O_2387,N_16163,N_17762);
nand UO_2388 (O_2388,N_19074,N_18454);
xnor UO_2389 (O_2389,N_17761,N_17630);
and UO_2390 (O_2390,N_19772,N_18387);
and UO_2391 (O_2391,N_19615,N_17082);
nand UO_2392 (O_2392,N_18691,N_19838);
or UO_2393 (O_2393,N_16645,N_17440);
and UO_2394 (O_2394,N_19710,N_19852);
xor UO_2395 (O_2395,N_16181,N_18313);
nand UO_2396 (O_2396,N_16897,N_18169);
nor UO_2397 (O_2397,N_16761,N_17563);
nand UO_2398 (O_2398,N_17258,N_18631);
nand UO_2399 (O_2399,N_18931,N_16580);
nor UO_2400 (O_2400,N_19936,N_19496);
nand UO_2401 (O_2401,N_19415,N_18245);
nor UO_2402 (O_2402,N_18456,N_18569);
nor UO_2403 (O_2403,N_18543,N_18797);
nand UO_2404 (O_2404,N_19353,N_17834);
or UO_2405 (O_2405,N_18404,N_17488);
and UO_2406 (O_2406,N_17689,N_18198);
and UO_2407 (O_2407,N_19273,N_17485);
or UO_2408 (O_2408,N_17773,N_19282);
nor UO_2409 (O_2409,N_17636,N_18017);
xnor UO_2410 (O_2410,N_17381,N_18819);
nor UO_2411 (O_2411,N_16748,N_19465);
nand UO_2412 (O_2412,N_16850,N_18276);
or UO_2413 (O_2413,N_16514,N_19174);
and UO_2414 (O_2414,N_17578,N_18042);
nand UO_2415 (O_2415,N_19016,N_16598);
nand UO_2416 (O_2416,N_17339,N_17638);
nor UO_2417 (O_2417,N_19490,N_17714);
and UO_2418 (O_2418,N_17394,N_18002);
xor UO_2419 (O_2419,N_16189,N_18860);
nor UO_2420 (O_2420,N_16749,N_19047);
nor UO_2421 (O_2421,N_18507,N_18098);
nand UO_2422 (O_2422,N_19427,N_18037);
nand UO_2423 (O_2423,N_17322,N_19187);
nand UO_2424 (O_2424,N_16665,N_19044);
nor UO_2425 (O_2425,N_17190,N_17743);
nand UO_2426 (O_2426,N_17198,N_19985);
and UO_2427 (O_2427,N_18804,N_16597);
nand UO_2428 (O_2428,N_16893,N_18725);
and UO_2429 (O_2429,N_19422,N_18754);
nor UO_2430 (O_2430,N_17300,N_16969);
and UO_2431 (O_2431,N_17088,N_16535);
or UO_2432 (O_2432,N_18191,N_19263);
and UO_2433 (O_2433,N_18359,N_19220);
nor UO_2434 (O_2434,N_17335,N_19521);
or UO_2435 (O_2435,N_19434,N_16521);
nand UO_2436 (O_2436,N_18148,N_17619);
or UO_2437 (O_2437,N_17060,N_16846);
nand UO_2438 (O_2438,N_18199,N_17740);
nand UO_2439 (O_2439,N_18497,N_19284);
and UO_2440 (O_2440,N_18990,N_16508);
or UO_2441 (O_2441,N_17340,N_18751);
or UO_2442 (O_2442,N_16397,N_16944);
nand UO_2443 (O_2443,N_16725,N_18931);
nor UO_2444 (O_2444,N_16917,N_17179);
nand UO_2445 (O_2445,N_19916,N_17872);
nor UO_2446 (O_2446,N_18286,N_17043);
and UO_2447 (O_2447,N_19995,N_19314);
nor UO_2448 (O_2448,N_18015,N_18922);
and UO_2449 (O_2449,N_18273,N_19481);
xnor UO_2450 (O_2450,N_18318,N_16287);
or UO_2451 (O_2451,N_18958,N_18811);
nand UO_2452 (O_2452,N_19863,N_17343);
nor UO_2453 (O_2453,N_18189,N_19964);
nand UO_2454 (O_2454,N_17863,N_18107);
and UO_2455 (O_2455,N_16040,N_17493);
nand UO_2456 (O_2456,N_18683,N_17823);
nand UO_2457 (O_2457,N_17878,N_18221);
nor UO_2458 (O_2458,N_18172,N_16924);
and UO_2459 (O_2459,N_16567,N_18994);
nor UO_2460 (O_2460,N_18254,N_19666);
nor UO_2461 (O_2461,N_19145,N_16248);
or UO_2462 (O_2462,N_16806,N_18389);
nor UO_2463 (O_2463,N_19030,N_19736);
xor UO_2464 (O_2464,N_16404,N_18907);
or UO_2465 (O_2465,N_19106,N_17061);
nand UO_2466 (O_2466,N_16043,N_19331);
and UO_2467 (O_2467,N_19162,N_19694);
nand UO_2468 (O_2468,N_17196,N_19007);
nand UO_2469 (O_2469,N_18682,N_16029);
nor UO_2470 (O_2470,N_18705,N_18708);
nand UO_2471 (O_2471,N_19453,N_16411);
and UO_2472 (O_2472,N_19041,N_18038);
xnor UO_2473 (O_2473,N_18881,N_17899);
nand UO_2474 (O_2474,N_19200,N_18035);
nand UO_2475 (O_2475,N_17878,N_17501);
and UO_2476 (O_2476,N_19388,N_18343);
nor UO_2477 (O_2477,N_18117,N_19080);
and UO_2478 (O_2478,N_18639,N_18801);
or UO_2479 (O_2479,N_16334,N_18294);
or UO_2480 (O_2480,N_17455,N_17913);
and UO_2481 (O_2481,N_16952,N_18323);
nand UO_2482 (O_2482,N_18774,N_17804);
or UO_2483 (O_2483,N_16179,N_19224);
nand UO_2484 (O_2484,N_17233,N_18773);
nor UO_2485 (O_2485,N_18974,N_19293);
and UO_2486 (O_2486,N_17139,N_16889);
or UO_2487 (O_2487,N_17502,N_17875);
nand UO_2488 (O_2488,N_17414,N_18013);
and UO_2489 (O_2489,N_17500,N_17428);
xnor UO_2490 (O_2490,N_18911,N_19398);
xor UO_2491 (O_2491,N_17201,N_16374);
nand UO_2492 (O_2492,N_16214,N_16206);
or UO_2493 (O_2493,N_17900,N_18547);
and UO_2494 (O_2494,N_18488,N_16056);
nand UO_2495 (O_2495,N_16393,N_17781);
nor UO_2496 (O_2496,N_16903,N_19515);
or UO_2497 (O_2497,N_17729,N_17471);
and UO_2498 (O_2498,N_18912,N_19514);
xor UO_2499 (O_2499,N_18576,N_19726);
endmodule