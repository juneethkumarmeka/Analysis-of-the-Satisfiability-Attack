module basic_500_3000_500_3_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_494,In_308);
and U1 (N_1,In_323,In_418);
nor U2 (N_2,In_103,In_100);
nor U3 (N_3,In_208,In_422);
xnor U4 (N_4,In_282,In_120);
or U5 (N_5,In_371,In_463);
nor U6 (N_6,In_246,In_217);
nor U7 (N_7,In_393,In_264);
xnor U8 (N_8,In_295,In_115);
nor U9 (N_9,In_209,In_78);
nor U10 (N_10,In_236,In_343);
and U11 (N_11,In_234,In_222);
and U12 (N_12,In_257,In_170);
nor U13 (N_13,In_486,In_2);
nor U14 (N_14,In_16,In_70);
or U15 (N_15,In_98,In_336);
nor U16 (N_16,In_376,In_91);
nand U17 (N_17,In_347,In_90);
nor U18 (N_18,In_411,In_454);
or U19 (N_19,In_262,In_298);
or U20 (N_20,In_95,In_297);
and U21 (N_21,In_477,In_232);
or U22 (N_22,In_395,In_3);
nand U23 (N_23,In_390,In_263);
and U24 (N_24,In_27,In_169);
nand U25 (N_25,In_230,In_333);
or U26 (N_26,In_14,In_215);
or U27 (N_27,In_438,In_324);
or U28 (N_28,In_174,In_203);
nor U29 (N_29,In_200,In_121);
and U30 (N_30,In_434,In_315);
or U31 (N_31,In_465,In_116);
nor U32 (N_32,In_55,In_173);
or U33 (N_33,In_400,In_41);
nand U34 (N_34,In_410,In_417);
and U35 (N_35,In_310,In_199);
nor U36 (N_36,In_387,In_1);
nand U37 (N_37,In_483,In_441);
nor U38 (N_38,In_216,In_34);
nor U39 (N_39,In_412,In_272);
and U40 (N_40,In_277,In_357);
nand U41 (N_41,In_498,In_339);
nand U42 (N_42,In_276,In_171);
nor U43 (N_43,In_131,In_109);
nand U44 (N_44,In_351,In_221);
and U45 (N_45,In_348,In_142);
nand U46 (N_46,In_460,In_129);
and U47 (N_47,In_374,In_488);
and U48 (N_48,In_327,In_83);
and U49 (N_49,In_338,In_96);
nand U50 (N_50,In_123,In_102);
or U51 (N_51,In_243,In_449);
and U52 (N_52,In_63,In_231);
nand U53 (N_53,In_163,In_9);
and U54 (N_54,In_487,In_185);
and U55 (N_55,In_349,In_495);
or U56 (N_56,In_139,In_396);
nand U57 (N_57,In_341,In_304);
or U58 (N_58,In_320,In_290);
and U59 (N_59,In_401,In_17);
and U60 (N_60,In_162,In_244);
and U61 (N_61,In_255,In_453);
nor U62 (N_62,In_447,In_152);
or U63 (N_63,In_223,In_193);
or U64 (N_64,In_452,In_285);
or U65 (N_65,In_134,In_114);
nand U66 (N_66,In_398,In_358);
and U67 (N_67,In_72,In_479);
nor U68 (N_68,In_287,In_172);
or U69 (N_69,In_226,In_268);
and U70 (N_70,In_196,In_256);
nor U71 (N_71,In_135,In_427);
xnor U72 (N_72,In_367,In_275);
or U73 (N_73,In_490,In_423);
or U74 (N_74,In_77,In_79);
or U75 (N_75,In_24,In_270);
or U76 (N_76,In_286,In_457);
nand U77 (N_77,In_408,In_180);
nor U78 (N_78,In_388,In_312);
nand U79 (N_79,In_440,In_4);
nor U80 (N_80,In_106,In_66);
or U81 (N_81,In_154,In_157);
xnor U82 (N_82,In_303,In_480);
nor U83 (N_83,In_86,In_12);
nand U84 (N_84,In_190,In_380);
and U85 (N_85,In_161,In_273);
nand U86 (N_86,In_108,In_294);
and U87 (N_87,In_326,In_187);
and U88 (N_88,In_489,In_296);
and U89 (N_89,In_325,In_425);
and U90 (N_90,In_68,In_237);
nor U91 (N_91,In_322,In_93);
nand U92 (N_92,In_458,In_317);
and U93 (N_93,In_119,In_168);
nand U94 (N_94,In_403,In_240);
nor U95 (N_95,In_469,In_151);
or U96 (N_96,In_213,In_355);
nand U97 (N_97,In_112,In_318);
or U98 (N_98,In_113,In_197);
nor U99 (N_99,In_379,In_342);
nand U100 (N_100,In_56,In_145);
nor U101 (N_101,In_136,In_265);
nor U102 (N_102,In_143,In_73);
or U103 (N_103,In_468,In_130);
and U104 (N_104,In_58,In_241);
nor U105 (N_105,In_62,In_385);
nor U106 (N_106,In_291,In_155);
and U107 (N_107,In_133,In_110);
or U108 (N_108,In_225,In_175);
nor U109 (N_109,In_330,In_84);
nor U110 (N_110,In_314,In_178);
and U111 (N_111,In_316,In_309);
or U112 (N_112,In_179,In_210);
nor U113 (N_113,In_445,In_75);
nand U114 (N_114,In_87,In_111);
or U115 (N_115,In_7,In_181);
nand U116 (N_116,In_271,In_331);
nand U117 (N_117,In_370,In_212);
and U118 (N_118,In_364,In_424);
nand U119 (N_119,In_25,In_127);
nor U120 (N_120,In_26,In_462);
nor U121 (N_121,In_67,In_284);
nor U122 (N_122,In_207,In_426);
or U123 (N_123,In_356,In_476);
or U124 (N_124,In_220,In_433);
nand U125 (N_125,In_269,In_206);
nor U126 (N_126,In_321,In_247);
or U127 (N_127,In_436,In_101);
nand U128 (N_128,In_383,In_253);
nand U129 (N_129,In_20,In_354);
and U130 (N_130,In_267,In_499);
nand U131 (N_131,In_332,In_429);
nand U132 (N_132,In_82,In_36);
nand U133 (N_133,In_205,In_259);
nor U134 (N_134,In_250,In_340);
nand U135 (N_135,In_252,In_183);
nand U136 (N_136,In_360,In_328);
nand U137 (N_137,In_392,In_335);
and U138 (N_138,In_368,In_413);
or U139 (N_139,In_382,In_283);
nor U140 (N_140,In_496,In_431);
nor U141 (N_141,In_53,In_52);
nor U142 (N_142,In_165,In_45);
nand U143 (N_143,In_38,In_43);
and U144 (N_144,In_153,In_470);
and U145 (N_145,In_279,In_474);
nand U146 (N_146,In_61,In_245);
nor U147 (N_147,In_194,In_88);
nor U148 (N_148,In_435,In_482);
nor U149 (N_149,In_473,In_137);
or U150 (N_150,In_99,In_258);
and U151 (N_151,In_409,In_365);
nand U152 (N_152,In_81,In_92);
nand U153 (N_153,In_233,In_132);
nor U154 (N_154,In_42,In_192);
nand U155 (N_155,In_307,In_299);
or U156 (N_156,In_421,In_359);
and U157 (N_157,In_419,In_144);
nor U158 (N_158,In_344,In_471);
nor U159 (N_159,In_118,In_147);
and U160 (N_160,In_140,In_198);
nand U161 (N_161,In_195,In_74);
nand U162 (N_162,In_158,In_439);
and U163 (N_163,In_218,In_202);
or U164 (N_164,In_302,In_117);
and U165 (N_165,In_229,In_47);
or U166 (N_166,In_278,In_451);
and U167 (N_167,In_107,In_39);
nand U168 (N_168,In_345,In_94);
nor U169 (N_169,In_21,In_289);
nand U170 (N_170,In_46,In_346);
nand U171 (N_171,In_22,In_405);
and U172 (N_172,In_455,In_64);
nor U173 (N_173,In_397,In_149);
or U174 (N_174,In_8,In_399);
or U175 (N_175,In_352,In_50);
or U176 (N_176,In_432,In_485);
nand U177 (N_177,In_76,In_366);
nor U178 (N_178,In_160,In_394);
nor U179 (N_179,In_146,In_159);
or U180 (N_180,In_15,In_0);
nand U181 (N_181,In_211,In_334);
nand U182 (N_182,In_481,In_126);
nand U183 (N_183,In_249,In_238);
or U184 (N_184,In_386,In_260);
nand U185 (N_185,In_49,In_402);
or U186 (N_186,In_391,In_493);
nor U187 (N_187,In_11,In_235);
or U188 (N_188,In_300,In_35);
nor U189 (N_189,In_497,In_51);
nor U190 (N_190,In_228,In_167);
and U191 (N_191,In_375,In_60);
nor U192 (N_192,In_442,In_362);
nand U193 (N_193,In_464,In_23);
nand U194 (N_194,In_448,In_239);
and U195 (N_195,In_122,In_329);
nand U196 (N_196,In_71,In_124);
nor U197 (N_197,In_176,In_384);
nand U198 (N_198,In_188,In_150);
nand U199 (N_199,In_6,In_475);
nor U200 (N_200,In_242,In_361);
nor U201 (N_201,In_189,In_373);
nand U202 (N_202,In_80,In_104);
and U203 (N_203,In_443,In_166);
nor U204 (N_204,In_311,In_288);
or U205 (N_205,In_404,In_461);
nand U206 (N_206,In_491,In_372);
nand U207 (N_207,In_29,In_301);
and U208 (N_208,In_456,In_156);
or U209 (N_209,In_19,In_292);
and U210 (N_210,In_57,In_416);
nand U211 (N_211,In_459,In_184);
nor U212 (N_212,In_13,In_444);
nor U213 (N_213,In_428,In_261);
and U214 (N_214,In_227,In_37);
xor U215 (N_215,In_201,In_97);
and U216 (N_216,In_420,In_138);
or U217 (N_217,In_65,In_484);
nand U218 (N_218,In_467,In_105);
nor U219 (N_219,In_389,In_28);
nor U220 (N_220,In_251,In_378);
or U221 (N_221,In_472,In_492);
nand U222 (N_222,In_319,In_350);
xor U223 (N_223,In_48,In_437);
nor U224 (N_224,In_40,In_182);
and U225 (N_225,In_44,In_280);
nand U226 (N_226,In_415,In_450);
nand U227 (N_227,In_148,In_377);
nor U228 (N_228,In_125,In_306);
or U229 (N_229,In_363,In_224);
nand U230 (N_230,In_337,In_381);
or U231 (N_231,In_266,In_219);
nand U232 (N_232,In_54,In_18);
nand U233 (N_233,In_478,In_281);
and U234 (N_234,In_31,In_274);
nand U235 (N_235,In_33,In_5);
and U236 (N_236,In_69,In_186);
nor U237 (N_237,In_466,In_10);
or U238 (N_238,In_164,In_191);
nor U239 (N_239,In_177,In_89);
xor U240 (N_240,In_369,In_214);
or U241 (N_241,In_305,In_248);
and U242 (N_242,In_430,In_254);
nor U243 (N_243,In_59,In_204);
nand U244 (N_244,In_293,In_32);
and U245 (N_245,In_128,In_85);
or U246 (N_246,In_407,In_141);
and U247 (N_247,In_30,In_353);
or U248 (N_248,In_414,In_446);
or U249 (N_249,In_406,In_313);
and U250 (N_250,In_103,In_468);
and U251 (N_251,In_409,In_277);
or U252 (N_252,In_408,In_403);
nor U253 (N_253,In_386,In_70);
and U254 (N_254,In_335,In_83);
or U255 (N_255,In_144,In_121);
nor U256 (N_256,In_478,In_163);
or U257 (N_257,In_279,In_81);
nor U258 (N_258,In_263,In_3);
nor U259 (N_259,In_434,In_424);
and U260 (N_260,In_75,In_470);
or U261 (N_261,In_253,In_310);
nor U262 (N_262,In_394,In_219);
and U263 (N_263,In_456,In_449);
nor U264 (N_264,In_216,In_120);
nand U265 (N_265,In_83,In_417);
and U266 (N_266,In_473,In_277);
and U267 (N_267,In_321,In_242);
or U268 (N_268,In_226,In_319);
nor U269 (N_269,In_315,In_341);
nor U270 (N_270,In_13,In_22);
or U271 (N_271,In_488,In_137);
nand U272 (N_272,In_405,In_147);
nand U273 (N_273,In_336,In_466);
nor U274 (N_274,In_450,In_492);
nand U275 (N_275,In_441,In_103);
nand U276 (N_276,In_191,In_412);
and U277 (N_277,In_53,In_66);
or U278 (N_278,In_414,In_226);
and U279 (N_279,In_197,In_449);
nand U280 (N_280,In_379,In_158);
xor U281 (N_281,In_97,In_124);
or U282 (N_282,In_101,In_480);
nor U283 (N_283,In_399,In_27);
and U284 (N_284,In_475,In_467);
nand U285 (N_285,In_237,In_174);
and U286 (N_286,In_385,In_96);
xnor U287 (N_287,In_215,In_115);
or U288 (N_288,In_306,In_492);
or U289 (N_289,In_153,In_2);
or U290 (N_290,In_8,In_34);
nand U291 (N_291,In_29,In_102);
and U292 (N_292,In_449,In_193);
nand U293 (N_293,In_310,In_18);
nand U294 (N_294,In_492,In_114);
nand U295 (N_295,In_222,In_120);
nand U296 (N_296,In_356,In_330);
or U297 (N_297,In_16,In_113);
or U298 (N_298,In_408,In_213);
or U299 (N_299,In_93,In_463);
and U300 (N_300,In_373,In_23);
xnor U301 (N_301,In_328,In_467);
nand U302 (N_302,In_181,In_146);
or U303 (N_303,In_216,In_237);
or U304 (N_304,In_138,In_374);
nor U305 (N_305,In_137,In_397);
xor U306 (N_306,In_297,In_211);
or U307 (N_307,In_61,In_264);
and U308 (N_308,In_343,In_331);
nor U309 (N_309,In_333,In_189);
and U310 (N_310,In_70,In_472);
nand U311 (N_311,In_67,In_386);
or U312 (N_312,In_80,In_166);
nor U313 (N_313,In_81,In_273);
nor U314 (N_314,In_370,In_83);
nand U315 (N_315,In_54,In_9);
nor U316 (N_316,In_304,In_185);
nand U317 (N_317,In_285,In_278);
xnor U318 (N_318,In_220,In_79);
nor U319 (N_319,In_222,In_327);
and U320 (N_320,In_428,In_349);
nand U321 (N_321,In_64,In_49);
or U322 (N_322,In_413,In_319);
nand U323 (N_323,In_499,In_95);
nor U324 (N_324,In_82,In_154);
or U325 (N_325,In_185,In_269);
nand U326 (N_326,In_83,In_251);
and U327 (N_327,In_242,In_107);
and U328 (N_328,In_73,In_289);
or U329 (N_329,In_289,In_74);
nor U330 (N_330,In_246,In_363);
nor U331 (N_331,In_246,In_424);
nor U332 (N_332,In_274,In_427);
nand U333 (N_333,In_160,In_460);
or U334 (N_334,In_309,In_326);
nand U335 (N_335,In_78,In_205);
nand U336 (N_336,In_57,In_350);
nor U337 (N_337,In_304,In_357);
nand U338 (N_338,In_106,In_397);
nor U339 (N_339,In_227,In_109);
or U340 (N_340,In_75,In_215);
or U341 (N_341,In_213,In_237);
nand U342 (N_342,In_316,In_144);
xor U343 (N_343,In_408,In_189);
or U344 (N_344,In_30,In_202);
or U345 (N_345,In_461,In_399);
nor U346 (N_346,In_175,In_452);
xor U347 (N_347,In_423,In_494);
or U348 (N_348,In_343,In_317);
xor U349 (N_349,In_265,In_350);
and U350 (N_350,In_156,In_442);
nor U351 (N_351,In_138,In_287);
nand U352 (N_352,In_225,In_21);
or U353 (N_353,In_284,In_237);
and U354 (N_354,In_75,In_43);
nor U355 (N_355,In_314,In_341);
and U356 (N_356,In_334,In_356);
nand U357 (N_357,In_179,In_467);
or U358 (N_358,In_315,In_218);
nand U359 (N_359,In_35,In_416);
nor U360 (N_360,In_215,In_341);
nand U361 (N_361,In_117,In_337);
nor U362 (N_362,In_402,In_112);
or U363 (N_363,In_142,In_21);
nor U364 (N_364,In_322,In_36);
or U365 (N_365,In_493,In_80);
and U366 (N_366,In_259,In_151);
and U367 (N_367,In_85,In_339);
or U368 (N_368,In_92,In_223);
nand U369 (N_369,In_176,In_91);
or U370 (N_370,In_148,In_169);
nor U371 (N_371,In_89,In_203);
nand U372 (N_372,In_211,In_292);
or U373 (N_373,In_437,In_321);
nor U374 (N_374,In_368,In_259);
and U375 (N_375,In_164,In_171);
nand U376 (N_376,In_159,In_194);
nor U377 (N_377,In_148,In_274);
and U378 (N_378,In_16,In_267);
nor U379 (N_379,In_354,In_421);
or U380 (N_380,In_152,In_58);
or U381 (N_381,In_221,In_227);
nor U382 (N_382,In_326,In_51);
and U383 (N_383,In_107,In_450);
nor U384 (N_384,In_448,In_90);
and U385 (N_385,In_369,In_152);
nand U386 (N_386,In_376,In_136);
nand U387 (N_387,In_67,In_306);
or U388 (N_388,In_464,In_54);
nor U389 (N_389,In_484,In_155);
nor U390 (N_390,In_302,In_138);
nor U391 (N_391,In_163,In_224);
nand U392 (N_392,In_163,In_214);
nor U393 (N_393,In_395,In_12);
or U394 (N_394,In_325,In_62);
nand U395 (N_395,In_228,In_400);
nand U396 (N_396,In_357,In_128);
or U397 (N_397,In_230,In_51);
or U398 (N_398,In_122,In_406);
and U399 (N_399,In_370,In_452);
and U400 (N_400,In_29,In_359);
nor U401 (N_401,In_359,In_317);
nand U402 (N_402,In_414,In_388);
and U403 (N_403,In_341,In_482);
xnor U404 (N_404,In_238,In_45);
nand U405 (N_405,In_433,In_438);
or U406 (N_406,In_486,In_209);
or U407 (N_407,In_477,In_189);
nand U408 (N_408,In_230,In_98);
or U409 (N_409,In_58,In_134);
nand U410 (N_410,In_396,In_91);
nand U411 (N_411,In_173,In_117);
or U412 (N_412,In_22,In_324);
or U413 (N_413,In_195,In_24);
or U414 (N_414,In_428,In_398);
nand U415 (N_415,In_408,In_467);
nand U416 (N_416,In_222,In_376);
nor U417 (N_417,In_288,In_464);
nand U418 (N_418,In_314,In_148);
and U419 (N_419,In_99,In_211);
nor U420 (N_420,In_358,In_260);
nor U421 (N_421,In_160,In_105);
or U422 (N_422,In_235,In_261);
or U423 (N_423,In_482,In_406);
nand U424 (N_424,In_77,In_434);
and U425 (N_425,In_299,In_167);
nand U426 (N_426,In_346,In_52);
nor U427 (N_427,In_478,In_378);
nor U428 (N_428,In_248,In_122);
nand U429 (N_429,In_233,In_247);
or U430 (N_430,In_229,In_64);
nor U431 (N_431,In_464,In_330);
nand U432 (N_432,In_490,In_300);
nand U433 (N_433,In_462,In_492);
nand U434 (N_434,In_238,In_161);
nor U435 (N_435,In_39,In_210);
xnor U436 (N_436,In_364,In_175);
and U437 (N_437,In_422,In_73);
or U438 (N_438,In_167,In_206);
nand U439 (N_439,In_266,In_272);
nand U440 (N_440,In_59,In_78);
or U441 (N_441,In_35,In_144);
nor U442 (N_442,In_338,In_335);
and U443 (N_443,In_303,In_202);
nand U444 (N_444,In_495,In_301);
or U445 (N_445,In_484,In_172);
xor U446 (N_446,In_141,In_96);
nand U447 (N_447,In_321,In_187);
xor U448 (N_448,In_104,In_398);
nand U449 (N_449,In_341,In_84);
and U450 (N_450,In_268,In_374);
and U451 (N_451,In_181,In_456);
and U452 (N_452,In_364,In_323);
or U453 (N_453,In_196,In_381);
and U454 (N_454,In_0,In_135);
or U455 (N_455,In_437,In_399);
nand U456 (N_456,In_30,In_219);
nand U457 (N_457,In_56,In_491);
and U458 (N_458,In_408,In_333);
nand U459 (N_459,In_165,In_334);
nand U460 (N_460,In_203,In_464);
xnor U461 (N_461,In_154,In_290);
nand U462 (N_462,In_241,In_30);
nand U463 (N_463,In_155,In_251);
nand U464 (N_464,In_150,In_83);
nor U465 (N_465,In_192,In_476);
nor U466 (N_466,In_345,In_342);
nor U467 (N_467,In_197,In_458);
and U468 (N_468,In_202,In_82);
nand U469 (N_469,In_185,In_442);
and U470 (N_470,In_116,In_319);
or U471 (N_471,In_220,In_209);
and U472 (N_472,In_23,In_105);
and U473 (N_473,In_360,In_48);
nor U474 (N_474,In_176,In_178);
or U475 (N_475,In_201,In_381);
or U476 (N_476,In_306,In_390);
nand U477 (N_477,In_272,In_27);
nor U478 (N_478,In_280,In_428);
nand U479 (N_479,In_289,In_17);
or U480 (N_480,In_239,In_272);
or U481 (N_481,In_202,In_446);
and U482 (N_482,In_440,In_269);
or U483 (N_483,In_183,In_498);
and U484 (N_484,In_294,In_107);
nor U485 (N_485,In_390,In_63);
nand U486 (N_486,In_184,In_316);
or U487 (N_487,In_340,In_202);
or U488 (N_488,In_207,In_203);
or U489 (N_489,In_242,In_5);
and U490 (N_490,In_59,In_357);
nor U491 (N_491,In_83,In_390);
or U492 (N_492,In_197,In_444);
nand U493 (N_493,In_378,In_40);
nand U494 (N_494,In_257,In_198);
nor U495 (N_495,In_158,In_441);
nand U496 (N_496,In_275,In_155);
or U497 (N_497,In_423,In_147);
and U498 (N_498,In_20,In_144);
or U499 (N_499,In_275,In_91);
nor U500 (N_500,In_46,In_267);
nor U501 (N_501,In_395,In_294);
or U502 (N_502,In_344,In_189);
nor U503 (N_503,In_430,In_355);
or U504 (N_504,In_420,In_213);
nand U505 (N_505,In_27,In_215);
and U506 (N_506,In_108,In_207);
and U507 (N_507,In_270,In_126);
nor U508 (N_508,In_493,In_115);
nand U509 (N_509,In_151,In_294);
or U510 (N_510,In_406,In_109);
or U511 (N_511,In_126,In_408);
nand U512 (N_512,In_292,In_90);
and U513 (N_513,In_295,In_251);
nand U514 (N_514,In_20,In_186);
and U515 (N_515,In_188,In_298);
or U516 (N_516,In_200,In_237);
nor U517 (N_517,In_246,In_30);
or U518 (N_518,In_258,In_300);
nor U519 (N_519,In_343,In_387);
nand U520 (N_520,In_348,In_3);
and U521 (N_521,In_175,In_65);
nor U522 (N_522,In_376,In_287);
and U523 (N_523,In_15,In_80);
nand U524 (N_524,In_98,In_278);
and U525 (N_525,In_415,In_189);
or U526 (N_526,In_299,In_187);
nand U527 (N_527,In_133,In_307);
nor U528 (N_528,In_342,In_265);
nand U529 (N_529,In_14,In_113);
and U530 (N_530,In_273,In_309);
and U531 (N_531,In_153,In_381);
or U532 (N_532,In_206,In_338);
or U533 (N_533,In_122,In_432);
nand U534 (N_534,In_305,In_350);
and U535 (N_535,In_280,In_346);
nand U536 (N_536,In_226,In_76);
nand U537 (N_537,In_434,In_71);
nand U538 (N_538,In_294,In_306);
nand U539 (N_539,In_246,In_283);
nor U540 (N_540,In_104,In_57);
or U541 (N_541,In_252,In_120);
and U542 (N_542,In_0,In_45);
nor U543 (N_543,In_113,In_231);
nor U544 (N_544,In_50,In_104);
nor U545 (N_545,In_137,In_264);
nor U546 (N_546,In_473,In_64);
xnor U547 (N_547,In_174,In_289);
and U548 (N_548,In_267,In_88);
nor U549 (N_549,In_26,In_441);
nor U550 (N_550,In_198,In_364);
nand U551 (N_551,In_87,In_410);
nand U552 (N_552,In_199,In_466);
or U553 (N_553,In_376,In_135);
and U554 (N_554,In_365,In_205);
nor U555 (N_555,In_7,In_175);
or U556 (N_556,In_175,In_211);
or U557 (N_557,In_140,In_401);
and U558 (N_558,In_381,In_23);
and U559 (N_559,In_176,In_453);
or U560 (N_560,In_491,In_476);
and U561 (N_561,In_207,In_370);
nand U562 (N_562,In_132,In_119);
nor U563 (N_563,In_48,In_410);
nor U564 (N_564,In_32,In_280);
nand U565 (N_565,In_152,In_243);
or U566 (N_566,In_377,In_124);
nand U567 (N_567,In_324,In_49);
nor U568 (N_568,In_343,In_335);
nand U569 (N_569,In_310,In_210);
nor U570 (N_570,In_492,In_135);
and U571 (N_571,In_181,In_399);
nor U572 (N_572,In_468,In_53);
nor U573 (N_573,In_254,In_26);
and U574 (N_574,In_276,In_399);
and U575 (N_575,In_251,In_491);
or U576 (N_576,In_41,In_247);
or U577 (N_577,In_359,In_7);
or U578 (N_578,In_65,In_207);
nand U579 (N_579,In_320,In_379);
or U580 (N_580,In_223,In_67);
nor U581 (N_581,In_278,In_159);
nand U582 (N_582,In_318,In_116);
and U583 (N_583,In_243,In_332);
or U584 (N_584,In_428,In_492);
nand U585 (N_585,In_38,In_422);
and U586 (N_586,In_451,In_488);
and U587 (N_587,In_325,In_195);
and U588 (N_588,In_207,In_201);
or U589 (N_589,In_191,In_445);
and U590 (N_590,In_176,In_366);
nand U591 (N_591,In_279,In_455);
nor U592 (N_592,In_398,In_337);
and U593 (N_593,In_179,In_482);
and U594 (N_594,In_150,In_130);
or U595 (N_595,In_73,In_107);
and U596 (N_596,In_81,In_314);
and U597 (N_597,In_179,In_19);
and U598 (N_598,In_218,In_233);
nor U599 (N_599,In_475,In_438);
and U600 (N_600,In_232,In_228);
nor U601 (N_601,In_330,In_9);
and U602 (N_602,In_124,In_413);
or U603 (N_603,In_423,In_127);
or U604 (N_604,In_292,In_380);
and U605 (N_605,In_450,In_260);
nand U606 (N_606,In_109,In_474);
nand U607 (N_607,In_192,In_285);
nor U608 (N_608,In_5,In_364);
nor U609 (N_609,In_453,In_216);
and U610 (N_610,In_59,In_91);
and U611 (N_611,In_413,In_37);
and U612 (N_612,In_10,In_173);
nand U613 (N_613,In_76,In_86);
or U614 (N_614,In_385,In_167);
nor U615 (N_615,In_194,In_151);
nand U616 (N_616,In_92,In_203);
nand U617 (N_617,In_437,In_74);
nand U618 (N_618,In_292,In_149);
and U619 (N_619,In_390,In_184);
nand U620 (N_620,In_200,In_246);
or U621 (N_621,In_25,In_394);
nand U622 (N_622,In_175,In_230);
or U623 (N_623,In_247,In_168);
and U624 (N_624,In_477,In_102);
nand U625 (N_625,In_109,In_324);
or U626 (N_626,In_147,In_106);
and U627 (N_627,In_166,In_302);
nor U628 (N_628,In_102,In_414);
and U629 (N_629,In_200,In_447);
and U630 (N_630,In_427,In_371);
and U631 (N_631,In_110,In_218);
or U632 (N_632,In_22,In_425);
or U633 (N_633,In_310,In_409);
or U634 (N_634,In_258,In_243);
nor U635 (N_635,In_258,In_440);
nand U636 (N_636,In_160,In_181);
nand U637 (N_637,In_325,In_115);
nand U638 (N_638,In_446,In_274);
and U639 (N_639,In_409,In_62);
nor U640 (N_640,In_131,In_160);
xor U641 (N_641,In_196,In_467);
and U642 (N_642,In_232,In_346);
nand U643 (N_643,In_8,In_291);
or U644 (N_644,In_113,In_11);
nor U645 (N_645,In_379,In_392);
nand U646 (N_646,In_8,In_191);
and U647 (N_647,In_46,In_180);
nand U648 (N_648,In_247,In_481);
nor U649 (N_649,In_468,In_206);
nand U650 (N_650,In_223,In_54);
nand U651 (N_651,In_110,In_33);
or U652 (N_652,In_227,In_273);
and U653 (N_653,In_117,In_413);
nor U654 (N_654,In_405,In_264);
nor U655 (N_655,In_401,In_405);
nor U656 (N_656,In_373,In_411);
nor U657 (N_657,In_320,In_498);
xor U658 (N_658,In_168,In_409);
nand U659 (N_659,In_468,In_254);
nor U660 (N_660,In_102,In_315);
or U661 (N_661,In_423,In_214);
nor U662 (N_662,In_239,In_48);
or U663 (N_663,In_293,In_79);
nand U664 (N_664,In_42,In_410);
nand U665 (N_665,In_269,In_270);
nor U666 (N_666,In_32,In_447);
and U667 (N_667,In_285,In_459);
or U668 (N_668,In_274,In_312);
nand U669 (N_669,In_354,In_144);
or U670 (N_670,In_165,In_283);
and U671 (N_671,In_77,In_473);
or U672 (N_672,In_313,In_241);
or U673 (N_673,In_432,In_196);
and U674 (N_674,In_371,In_294);
or U675 (N_675,In_346,In_279);
or U676 (N_676,In_207,In_19);
nor U677 (N_677,In_272,In_414);
or U678 (N_678,In_79,In_402);
and U679 (N_679,In_344,In_374);
nand U680 (N_680,In_54,In_122);
and U681 (N_681,In_218,In_24);
nor U682 (N_682,In_313,In_154);
nand U683 (N_683,In_378,In_44);
nor U684 (N_684,In_171,In_478);
nand U685 (N_685,In_73,In_433);
nand U686 (N_686,In_55,In_382);
nor U687 (N_687,In_315,In_58);
or U688 (N_688,In_241,In_447);
nor U689 (N_689,In_255,In_187);
nor U690 (N_690,In_334,In_273);
or U691 (N_691,In_289,In_109);
or U692 (N_692,In_352,In_54);
and U693 (N_693,In_332,In_173);
nor U694 (N_694,In_158,In_260);
nor U695 (N_695,In_495,In_94);
nor U696 (N_696,In_426,In_356);
nand U697 (N_697,In_66,In_459);
or U698 (N_698,In_102,In_290);
or U699 (N_699,In_241,In_119);
or U700 (N_700,In_492,In_11);
or U701 (N_701,In_365,In_312);
and U702 (N_702,In_151,In_176);
or U703 (N_703,In_344,In_399);
nor U704 (N_704,In_145,In_269);
nor U705 (N_705,In_204,In_338);
nor U706 (N_706,In_50,In_60);
and U707 (N_707,In_161,In_486);
and U708 (N_708,In_134,In_449);
nand U709 (N_709,In_139,In_72);
and U710 (N_710,In_346,In_65);
nand U711 (N_711,In_468,In_257);
nand U712 (N_712,In_336,In_224);
nor U713 (N_713,In_489,In_233);
or U714 (N_714,In_242,In_239);
or U715 (N_715,In_97,In_61);
and U716 (N_716,In_494,In_460);
nand U717 (N_717,In_320,In_22);
or U718 (N_718,In_403,In_162);
nand U719 (N_719,In_72,In_119);
nand U720 (N_720,In_411,In_61);
or U721 (N_721,In_44,In_445);
or U722 (N_722,In_106,In_23);
nand U723 (N_723,In_403,In_317);
or U724 (N_724,In_308,In_368);
and U725 (N_725,In_234,In_389);
or U726 (N_726,In_415,In_101);
or U727 (N_727,In_19,In_55);
and U728 (N_728,In_487,In_398);
nor U729 (N_729,In_437,In_232);
nor U730 (N_730,In_253,In_244);
nor U731 (N_731,In_442,In_452);
or U732 (N_732,In_491,In_438);
nor U733 (N_733,In_25,In_442);
nor U734 (N_734,In_392,In_282);
nor U735 (N_735,In_276,In_217);
nor U736 (N_736,In_436,In_379);
or U737 (N_737,In_330,In_410);
nor U738 (N_738,In_151,In_75);
nand U739 (N_739,In_209,In_92);
and U740 (N_740,In_8,In_123);
nand U741 (N_741,In_162,In_116);
nand U742 (N_742,In_242,In_266);
or U743 (N_743,In_110,In_1);
or U744 (N_744,In_468,In_270);
nor U745 (N_745,In_459,In_312);
nand U746 (N_746,In_11,In_79);
nand U747 (N_747,In_238,In_151);
and U748 (N_748,In_431,In_463);
nor U749 (N_749,In_172,In_392);
or U750 (N_750,In_460,In_210);
nor U751 (N_751,In_249,In_23);
and U752 (N_752,In_485,In_417);
or U753 (N_753,In_245,In_170);
or U754 (N_754,In_447,In_235);
nand U755 (N_755,In_56,In_98);
or U756 (N_756,In_153,In_75);
nor U757 (N_757,In_167,In_10);
or U758 (N_758,In_241,In_433);
nor U759 (N_759,In_80,In_421);
and U760 (N_760,In_272,In_235);
and U761 (N_761,In_385,In_28);
nor U762 (N_762,In_379,In_318);
and U763 (N_763,In_444,In_364);
nand U764 (N_764,In_300,In_175);
or U765 (N_765,In_220,In_370);
or U766 (N_766,In_370,In_15);
nand U767 (N_767,In_142,In_298);
nand U768 (N_768,In_134,In_69);
nand U769 (N_769,In_477,In_435);
and U770 (N_770,In_385,In_380);
or U771 (N_771,In_264,In_389);
or U772 (N_772,In_372,In_205);
nand U773 (N_773,In_280,In_112);
nor U774 (N_774,In_489,In_466);
nor U775 (N_775,In_262,In_135);
or U776 (N_776,In_149,In_5);
nor U777 (N_777,In_299,In_413);
and U778 (N_778,In_43,In_368);
and U779 (N_779,In_280,In_34);
xnor U780 (N_780,In_94,In_42);
xor U781 (N_781,In_497,In_495);
or U782 (N_782,In_113,In_413);
and U783 (N_783,In_478,In_304);
nor U784 (N_784,In_396,In_333);
or U785 (N_785,In_225,In_490);
nand U786 (N_786,In_432,In_158);
or U787 (N_787,In_71,In_134);
and U788 (N_788,In_266,In_305);
or U789 (N_789,In_486,In_164);
or U790 (N_790,In_198,In_356);
nor U791 (N_791,In_28,In_205);
nand U792 (N_792,In_18,In_163);
nand U793 (N_793,In_173,In_475);
and U794 (N_794,In_169,In_396);
and U795 (N_795,In_362,In_379);
nor U796 (N_796,In_23,In_253);
nor U797 (N_797,In_407,In_428);
and U798 (N_798,In_143,In_447);
and U799 (N_799,In_417,In_260);
nor U800 (N_800,In_487,In_112);
or U801 (N_801,In_437,In_477);
nor U802 (N_802,In_477,In_155);
nor U803 (N_803,In_147,In_28);
and U804 (N_804,In_52,In_288);
nor U805 (N_805,In_479,In_486);
nor U806 (N_806,In_232,In_446);
nor U807 (N_807,In_496,In_56);
nor U808 (N_808,In_383,In_289);
and U809 (N_809,In_346,In_243);
nand U810 (N_810,In_26,In_310);
or U811 (N_811,In_466,In_122);
or U812 (N_812,In_11,In_213);
nor U813 (N_813,In_245,In_376);
or U814 (N_814,In_471,In_382);
nand U815 (N_815,In_109,In_369);
and U816 (N_816,In_104,In_261);
nor U817 (N_817,In_309,In_104);
nand U818 (N_818,In_391,In_97);
nor U819 (N_819,In_130,In_159);
nand U820 (N_820,In_347,In_401);
xor U821 (N_821,In_230,In_233);
or U822 (N_822,In_159,In_227);
or U823 (N_823,In_237,In_46);
nor U824 (N_824,In_220,In_253);
and U825 (N_825,In_293,In_75);
nor U826 (N_826,In_428,In_19);
nand U827 (N_827,In_236,In_404);
and U828 (N_828,In_49,In_437);
and U829 (N_829,In_243,In_456);
xor U830 (N_830,In_496,In_109);
and U831 (N_831,In_206,In_112);
or U832 (N_832,In_288,In_386);
or U833 (N_833,In_342,In_283);
nand U834 (N_834,In_355,In_278);
nor U835 (N_835,In_92,In_213);
or U836 (N_836,In_288,In_221);
or U837 (N_837,In_354,In_251);
xor U838 (N_838,In_103,In_179);
nand U839 (N_839,In_284,In_219);
or U840 (N_840,In_473,In_51);
nand U841 (N_841,In_113,In_313);
nor U842 (N_842,In_65,In_45);
or U843 (N_843,In_27,In_167);
nor U844 (N_844,In_168,In_388);
or U845 (N_845,In_362,In_370);
nand U846 (N_846,In_14,In_18);
nand U847 (N_847,In_392,In_245);
nand U848 (N_848,In_428,In_467);
nand U849 (N_849,In_268,In_396);
and U850 (N_850,In_361,In_458);
and U851 (N_851,In_46,In_124);
nor U852 (N_852,In_89,In_393);
or U853 (N_853,In_90,In_4);
nand U854 (N_854,In_37,In_245);
or U855 (N_855,In_141,In_351);
and U856 (N_856,In_456,In_455);
nor U857 (N_857,In_42,In_429);
nand U858 (N_858,In_69,In_445);
or U859 (N_859,In_390,In_120);
and U860 (N_860,In_248,In_265);
or U861 (N_861,In_169,In_250);
or U862 (N_862,In_432,In_490);
nor U863 (N_863,In_423,In_335);
nand U864 (N_864,In_24,In_361);
nand U865 (N_865,In_244,In_35);
and U866 (N_866,In_290,In_8);
nand U867 (N_867,In_458,In_164);
or U868 (N_868,In_165,In_322);
xnor U869 (N_869,In_250,In_156);
nor U870 (N_870,In_334,In_406);
nor U871 (N_871,In_319,In_483);
nor U872 (N_872,In_429,In_196);
nand U873 (N_873,In_338,In_487);
or U874 (N_874,In_247,In_14);
nor U875 (N_875,In_48,In_499);
or U876 (N_876,In_387,In_266);
or U877 (N_877,In_499,In_112);
and U878 (N_878,In_141,In_497);
nor U879 (N_879,In_490,In_13);
and U880 (N_880,In_14,In_448);
nand U881 (N_881,In_3,In_356);
or U882 (N_882,In_282,In_455);
nand U883 (N_883,In_455,In_62);
and U884 (N_884,In_69,In_442);
or U885 (N_885,In_190,In_92);
nand U886 (N_886,In_359,In_276);
nor U887 (N_887,In_162,In_318);
and U888 (N_888,In_124,In_213);
and U889 (N_889,In_99,In_207);
and U890 (N_890,In_66,In_366);
nand U891 (N_891,In_194,In_244);
nand U892 (N_892,In_381,In_260);
nor U893 (N_893,In_48,In_403);
nor U894 (N_894,In_218,In_14);
nand U895 (N_895,In_496,In_95);
nor U896 (N_896,In_124,In_318);
nand U897 (N_897,In_50,In_97);
and U898 (N_898,In_330,In_192);
nor U899 (N_899,In_419,In_14);
and U900 (N_900,In_307,In_135);
nand U901 (N_901,In_253,In_432);
nand U902 (N_902,In_178,In_35);
nor U903 (N_903,In_200,In_319);
nor U904 (N_904,In_464,In_181);
and U905 (N_905,In_462,In_483);
nor U906 (N_906,In_451,In_443);
or U907 (N_907,In_352,In_333);
nand U908 (N_908,In_477,In_26);
nand U909 (N_909,In_350,In_215);
nand U910 (N_910,In_142,In_344);
nand U911 (N_911,In_82,In_298);
nand U912 (N_912,In_478,In_24);
and U913 (N_913,In_398,In_64);
and U914 (N_914,In_141,In_165);
and U915 (N_915,In_274,In_362);
nor U916 (N_916,In_297,In_346);
or U917 (N_917,In_368,In_154);
nor U918 (N_918,In_457,In_368);
nor U919 (N_919,In_367,In_238);
nand U920 (N_920,In_72,In_144);
nand U921 (N_921,In_51,In_115);
or U922 (N_922,In_397,In_105);
nand U923 (N_923,In_124,In_339);
nor U924 (N_924,In_380,In_71);
and U925 (N_925,In_258,In_92);
and U926 (N_926,In_128,In_69);
nor U927 (N_927,In_307,In_461);
and U928 (N_928,In_7,In_197);
nand U929 (N_929,In_450,In_195);
nand U930 (N_930,In_464,In_223);
and U931 (N_931,In_272,In_108);
nor U932 (N_932,In_258,In_152);
nand U933 (N_933,In_46,In_349);
nand U934 (N_934,In_388,In_189);
or U935 (N_935,In_443,In_384);
and U936 (N_936,In_63,In_349);
nand U937 (N_937,In_76,In_128);
nor U938 (N_938,In_351,In_113);
nand U939 (N_939,In_335,In_260);
nand U940 (N_940,In_11,In_130);
nand U941 (N_941,In_303,In_433);
or U942 (N_942,In_150,In_423);
or U943 (N_943,In_272,In_428);
nand U944 (N_944,In_266,In_29);
or U945 (N_945,In_221,In_287);
nor U946 (N_946,In_490,In_221);
nand U947 (N_947,In_91,In_331);
nor U948 (N_948,In_424,In_331);
nand U949 (N_949,In_302,In_136);
and U950 (N_950,In_253,In_391);
nor U951 (N_951,In_486,In_70);
or U952 (N_952,In_233,In_329);
nand U953 (N_953,In_481,In_215);
nand U954 (N_954,In_272,In_129);
nor U955 (N_955,In_327,In_144);
nor U956 (N_956,In_324,In_134);
nand U957 (N_957,In_140,In_122);
or U958 (N_958,In_235,In_190);
and U959 (N_959,In_329,In_453);
and U960 (N_960,In_378,In_180);
nor U961 (N_961,In_343,In_10);
nand U962 (N_962,In_442,In_313);
nor U963 (N_963,In_465,In_257);
and U964 (N_964,In_17,In_470);
nand U965 (N_965,In_61,In_64);
or U966 (N_966,In_45,In_194);
or U967 (N_967,In_443,In_79);
or U968 (N_968,In_131,In_11);
nand U969 (N_969,In_189,In_306);
or U970 (N_970,In_51,In_16);
or U971 (N_971,In_362,In_494);
nand U972 (N_972,In_100,In_275);
and U973 (N_973,In_130,In_399);
nor U974 (N_974,In_355,In_379);
nand U975 (N_975,In_383,In_493);
nor U976 (N_976,In_196,In_485);
nor U977 (N_977,In_454,In_481);
nor U978 (N_978,In_378,In_155);
and U979 (N_979,In_376,In_73);
nand U980 (N_980,In_455,In_344);
nand U981 (N_981,In_114,In_81);
nor U982 (N_982,In_34,In_148);
or U983 (N_983,In_280,In_259);
and U984 (N_984,In_86,In_36);
and U985 (N_985,In_333,In_170);
nand U986 (N_986,In_188,In_343);
nor U987 (N_987,In_243,In_182);
xnor U988 (N_988,In_398,In_298);
or U989 (N_989,In_105,In_408);
or U990 (N_990,In_120,In_361);
nand U991 (N_991,In_6,In_204);
or U992 (N_992,In_357,In_328);
xnor U993 (N_993,In_493,In_186);
nor U994 (N_994,In_14,In_181);
xor U995 (N_995,In_294,In_209);
or U996 (N_996,In_318,In_302);
nor U997 (N_997,In_67,In_31);
nor U998 (N_998,In_208,In_260);
and U999 (N_999,In_256,In_143);
or U1000 (N_1000,N_626,N_966);
or U1001 (N_1001,N_373,N_474);
or U1002 (N_1002,N_978,N_446);
nand U1003 (N_1003,N_28,N_103);
xor U1004 (N_1004,N_976,N_150);
xnor U1005 (N_1005,N_17,N_79);
and U1006 (N_1006,N_868,N_266);
nand U1007 (N_1007,N_121,N_859);
nor U1008 (N_1008,N_669,N_956);
or U1009 (N_1009,N_393,N_276);
nand U1010 (N_1010,N_720,N_9);
and U1011 (N_1011,N_597,N_456);
and U1012 (N_1012,N_149,N_361);
nor U1013 (N_1013,N_256,N_858);
nor U1014 (N_1014,N_535,N_621);
or U1015 (N_1015,N_118,N_277);
and U1016 (N_1016,N_551,N_719);
and U1017 (N_1017,N_717,N_916);
nand U1018 (N_1018,N_769,N_680);
nand U1019 (N_1019,N_245,N_210);
nand U1020 (N_1020,N_145,N_421);
or U1021 (N_1021,N_754,N_107);
nand U1022 (N_1022,N_102,N_968);
nor U1023 (N_1023,N_357,N_255);
nor U1024 (N_1024,N_13,N_42);
nand U1025 (N_1025,N_206,N_439);
nor U1026 (N_1026,N_967,N_812);
or U1027 (N_1027,N_142,N_243);
nor U1028 (N_1028,N_908,N_317);
nor U1029 (N_1029,N_259,N_852);
and U1030 (N_1030,N_606,N_557);
and U1031 (N_1031,N_157,N_499);
xnor U1032 (N_1032,N_774,N_485);
and U1033 (N_1033,N_242,N_162);
nor U1034 (N_1034,N_324,N_73);
or U1035 (N_1035,N_82,N_566);
xnor U1036 (N_1036,N_50,N_906);
or U1037 (N_1037,N_971,N_146);
and U1038 (N_1038,N_35,N_211);
and U1039 (N_1039,N_447,N_413);
nor U1040 (N_1040,N_133,N_716);
and U1041 (N_1041,N_166,N_625);
or U1042 (N_1042,N_470,N_177);
xnor U1043 (N_1043,N_386,N_296);
or U1044 (N_1044,N_780,N_476);
nand U1045 (N_1045,N_552,N_466);
and U1046 (N_1046,N_953,N_665);
nand U1047 (N_1047,N_152,N_471);
nor U1048 (N_1048,N_16,N_27);
and U1049 (N_1049,N_500,N_940);
or U1050 (N_1050,N_299,N_718);
and U1051 (N_1051,N_526,N_885);
or U1052 (N_1052,N_705,N_756);
nand U1053 (N_1053,N_935,N_725);
nand U1054 (N_1054,N_742,N_892);
and U1055 (N_1055,N_19,N_676);
nand U1056 (N_1056,N_737,N_576);
nand U1057 (N_1057,N_414,N_382);
nor U1058 (N_1058,N_850,N_931);
nand U1059 (N_1059,N_110,N_498);
nand U1060 (N_1060,N_528,N_723);
and U1061 (N_1061,N_587,N_563);
and U1062 (N_1062,N_882,N_332);
xnor U1063 (N_1063,N_970,N_825);
nand U1064 (N_1064,N_573,N_207);
and U1065 (N_1065,N_543,N_564);
or U1066 (N_1066,N_734,N_410);
xor U1067 (N_1067,N_348,N_538);
nand U1068 (N_1068,N_877,N_38);
nand U1069 (N_1069,N_699,N_448);
nand U1070 (N_1070,N_307,N_738);
or U1071 (N_1071,N_199,N_334);
and U1072 (N_1072,N_48,N_486);
nand U1073 (N_1073,N_463,N_219);
or U1074 (N_1074,N_689,N_525);
nor U1075 (N_1075,N_560,N_104);
nand U1076 (N_1076,N_865,N_338);
nand U1077 (N_1077,N_98,N_411);
or U1078 (N_1078,N_5,N_746);
nor U1079 (N_1079,N_811,N_53);
and U1080 (N_1080,N_436,N_261);
or U1081 (N_1081,N_612,N_640);
nor U1082 (N_1082,N_437,N_202);
and U1083 (N_1083,N_703,N_221);
or U1084 (N_1084,N_356,N_143);
or U1085 (N_1085,N_744,N_764);
nor U1086 (N_1086,N_36,N_325);
nor U1087 (N_1087,N_804,N_92);
and U1088 (N_1088,N_648,N_160);
or U1089 (N_1089,N_187,N_320);
nor U1090 (N_1090,N_955,N_26);
and U1091 (N_1091,N_319,N_924);
xor U1092 (N_1092,N_205,N_828);
or U1093 (N_1093,N_685,N_380);
and U1094 (N_1094,N_736,N_10);
nor U1095 (N_1095,N_113,N_22);
nor U1096 (N_1096,N_313,N_347);
and U1097 (N_1097,N_707,N_438);
and U1098 (N_1098,N_796,N_484);
nand U1099 (N_1099,N_403,N_71);
or U1100 (N_1100,N_252,N_427);
and U1101 (N_1101,N_937,N_189);
xor U1102 (N_1102,N_604,N_875);
and U1103 (N_1103,N_776,N_106);
nand U1104 (N_1104,N_747,N_661);
or U1105 (N_1105,N_568,N_947);
nor U1106 (N_1106,N_330,N_8);
or U1107 (N_1107,N_672,N_362);
nor U1108 (N_1108,N_743,N_925);
nand U1109 (N_1109,N_69,N_377);
nand U1110 (N_1110,N_819,N_312);
nand U1111 (N_1111,N_666,N_643);
or U1112 (N_1112,N_273,N_547);
nor U1113 (N_1113,N_602,N_588);
and U1114 (N_1114,N_579,N_695);
or U1115 (N_1115,N_749,N_425);
or U1116 (N_1116,N_833,N_853);
or U1117 (N_1117,N_141,N_546);
and U1118 (N_1118,N_954,N_548);
nor U1119 (N_1119,N_292,N_264);
or U1120 (N_1120,N_21,N_370);
nand U1121 (N_1121,N_772,N_235);
nand U1122 (N_1122,N_961,N_298);
nor U1123 (N_1123,N_383,N_37);
or U1124 (N_1124,N_511,N_387);
or U1125 (N_1125,N_675,N_980);
and U1126 (N_1126,N_706,N_810);
nand U1127 (N_1127,N_407,N_536);
nor U1128 (N_1128,N_558,N_899);
nor U1129 (N_1129,N_887,N_84);
nor U1130 (N_1130,N_663,N_763);
nor U1131 (N_1131,N_140,N_135);
and U1132 (N_1132,N_957,N_449);
or U1133 (N_1133,N_249,N_131);
nand U1134 (N_1134,N_432,N_992);
or U1135 (N_1135,N_275,N_314);
or U1136 (N_1136,N_807,N_731);
nor U1137 (N_1137,N_550,N_286);
nor U1138 (N_1138,N_979,N_326);
nor U1139 (N_1139,N_213,N_365);
xor U1140 (N_1140,N_590,N_431);
or U1141 (N_1141,N_866,N_180);
and U1142 (N_1142,N_842,N_801);
nand U1143 (N_1143,N_771,N_301);
or U1144 (N_1144,N_884,N_90);
nor U1145 (N_1145,N_698,N_185);
nand U1146 (N_1146,N_230,N_759);
or U1147 (N_1147,N_822,N_417);
nand U1148 (N_1148,N_328,N_70);
nand U1149 (N_1149,N_516,N_170);
xnor U1150 (N_1150,N_4,N_156);
and U1151 (N_1151,N_192,N_805);
or U1152 (N_1152,N_100,N_761);
and U1153 (N_1153,N_798,N_454);
nand U1154 (N_1154,N_639,N_635);
nand U1155 (N_1155,N_302,N_721);
and U1156 (N_1156,N_930,N_477);
or U1157 (N_1157,N_346,N_753);
nand U1158 (N_1158,N_297,N_901);
nand U1159 (N_1159,N_647,N_826);
nor U1160 (N_1160,N_782,N_41);
or U1161 (N_1161,N_862,N_946);
nand U1162 (N_1162,N_422,N_691);
nand U1163 (N_1163,N_282,N_111);
nor U1164 (N_1164,N_654,N_874);
and U1165 (N_1165,N_190,N_949);
nor U1166 (N_1166,N_818,N_915);
or U1167 (N_1167,N_455,N_932);
nand U1168 (N_1168,N_836,N_848);
nor U1169 (N_1169,N_129,N_800);
and U1170 (N_1170,N_784,N_503);
or U1171 (N_1171,N_351,N_684);
nor U1172 (N_1172,N_553,N_231);
nand U1173 (N_1173,N_770,N_23);
or U1174 (N_1174,N_274,N_914);
and U1175 (N_1175,N_857,N_603);
or U1176 (N_1176,N_331,N_589);
nand U1177 (N_1177,N_517,N_785);
nand U1178 (N_1178,N_962,N_618);
and U1179 (N_1179,N_944,N_504);
nand U1180 (N_1180,N_870,N_336);
nor U1181 (N_1181,N_806,N_729);
nor U1182 (N_1182,N_917,N_168);
and U1183 (N_1183,N_938,N_174);
nor U1184 (N_1184,N_963,N_339);
and U1185 (N_1185,N_983,N_136);
or U1186 (N_1186,N_869,N_234);
xnor U1187 (N_1187,N_952,N_343);
or U1188 (N_1188,N_673,N_767);
or U1189 (N_1189,N_327,N_309);
and U1190 (N_1190,N_775,N_555);
or U1191 (N_1191,N_667,N_502);
or U1192 (N_1192,N_481,N_873);
nor U1193 (N_1193,N_352,N_236);
nand U1194 (N_1194,N_722,N_164);
nand U1195 (N_1195,N_284,N_964);
or U1196 (N_1196,N_569,N_795);
or U1197 (N_1197,N_93,N_115);
or U1198 (N_1198,N_495,N_610);
or U1199 (N_1199,N_433,N_56);
and U1200 (N_1200,N_61,N_399);
or U1201 (N_1201,N_209,N_172);
nor U1202 (N_1202,N_493,N_829);
nand U1203 (N_1203,N_613,N_459);
nand U1204 (N_1204,N_167,N_677);
nand U1205 (N_1205,N_549,N_188);
nor U1206 (N_1206,N_122,N_60);
and U1207 (N_1207,N_175,N_396);
or U1208 (N_1208,N_641,N_64);
nand U1209 (N_1209,N_316,N_183);
and U1210 (N_1210,N_794,N_285);
and U1211 (N_1211,N_186,N_375);
nand U1212 (N_1212,N_492,N_994);
and U1213 (N_1213,N_398,N_817);
nand U1214 (N_1214,N_366,N_631);
nor U1215 (N_1215,N_374,N_305);
or U1216 (N_1216,N_620,N_47);
xnor U1217 (N_1217,N_600,N_598);
and U1218 (N_1218,N_44,N_975);
nor U1219 (N_1219,N_861,N_138);
and U1220 (N_1220,N_294,N_488);
and U1221 (N_1221,N_125,N_176);
and U1222 (N_1222,N_395,N_659);
or U1223 (N_1223,N_554,N_559);
or U1224 (N_1224,N_595,N_408);
nand U1225 (N_1225,N_350,N_792);
nand U1226 (N_1226,N_271,N_308);
nand U1227 (N_1227,N_419,N_445);
nand U1228 (N_1228,N_905,N_216);
nand U1229 (N_1229,N_834,N_575);
nor U1230 (N_1230,N_239,N_799);
nor U1231 (N_1231,N_389,N_902);
nor U1232 (N_1232,N_995,N_948);
and U1233 (N_1233,N_11,N_6);
nand U1234 (N_1234,N_123,N_519);
nor U1235 (N_1235,N_991,N_637);
and U1236 (N_1236,N_630,N_132);
nand U1237 (N_1237,N_268,N_39);
and U1238 (N_1238,N_478,N_533);
nand U1239 (N_1239,N_222,N_934);
or U1240 (N_1240,N_982,N_696);
nand U1241 (N_1241,N_959,N_435);
xnor U1242 (N_1242,N_751,N_986);
and U1243 (N_1243,N_879,N_593);
nor U1244 (N_1244,N_632,N_289);
or U1245 (N_1245,N_740,N_368);
nand U1246 (N_1246,N_318,N_75);
nor U1247 (N_1247,N_732,N_591);
and U1248 (N_1248,N_827,N_655);
and U1249 (N_1249,N_950,N_467);
and U1250 (N_1250,N_364,N_184);
or U1251 (N_1251,N_124,N_196);
or U1252 (N_1252,N_928,N_269);
or U1253 (N_1253,N_856,N_367);
nor U1254 (N_1254,N_712,N_824);
nor U1255 (N_1255,N_907,N_97);
and U1256 (N_1256,N_951,N_714);
nand U1257 (N_1257,N_67,N_945);
and U1258 (N_1258,N_522,N_910);
nand U1259 (N_1259,N_662,N_322);
or U1260 (N_1260,N_851,N_768);
nand U1261 (N_1261,N_808,N_708);
or U1262 (N_1262,N_674,N_741);
and U1263 (N_1263,N_344,N_497);
and U1264 (N_1264,N_406,N_614);
or U1265 (N_1265,N_227,N_394);
and U1266 (N_1266,N_473,N_974);
nand U1267 (N_1267,N_159,N_63);
or U1268 (N_1268,N_601,N_570);
nand U1269 (N_1269,N_893,N_173);
nand U1270 (N_1270,N_539,N_617);
and U1271 (N_1271,N_913,N_628);
or U1272 (N_1272,N_154,N_921);
nor U1273 (N_1273,N_897,N_83);
nor U1274 (N_1274,N_163,N_91);
or U1275 (N_1275,N_841,N_545);
and U1276 (N_1276,N_390,N_2);
or U1277 (N_1277,N_845,N_353);
xor U1278 (N_1278,N_624,N_127);
nand U1279 (N_1279,N_594,N_577);
and U1280 (N_1280,N_816,N_81);
nand U1281 (N_1281,N_909,N_397);
and U1282 (N_1282,N_629,N_889);
nor U1283 (N_1283,N_791,N_468);
nor U1284 (N_1284,N_311,N_670);
and U1285 (N_1285,N_74,N_181);
nand U1286 (N_1286,N_355,N_415);
and U1287 (N_1287,N_583,N_57);
nand U1288 (N_1288,N_537,N_730);
nor U1289 (N_1289,N_461,N_671);
or U1290 (N_1290,N_939,N_839);
or U1291 (N_1291,N_534,N_442);
and U1292 (N_1292,N_400,N_918);
or U1293 (N_1293,N_876,N_31);
or U1294 (N_1294,N_820,N_369);
or U1295 (N_1295,N_653,N_43);
nor U1296 (N_1296,N_993,N_489);
nand U1297 (N_1297,N_530,N_750);
nor U1298 (N_1298,N_809,N_457);
or U1299 (N_1299,N_426,N_960);
or U1300 (N_1300,N_409,N_863);
nor U1301 (N_1301,N_68,N_888);
and U1302 (N_1302,N_514,N_258);
or U1303 (N_1303,N_582,N_520);
and U1304 (N_1304,N_288,N_29);
nand U1305 (N_1305,N_996,N_223);
or U1306 (N_1306,N_927,N_1);
nor U1307 (N_1307,N_660,N_650);
nor U1308 (N_1308,N_844,N_658);
or U1309 (N_1309,N_765,N_611);
nand U1310 (N_1310,N_783,N_385);
or U1311 (N_1311,N_479,N_265);
and U1312 (N_1312,N_981,N_883);
or U1313 (N_1313,N_89,N_483);
nand U1314 (N_1314,N_758,N_838);
xor U1315 (N_1315,N_942,N_130);
or U1316 (N_1316,N_441,N_656);
or U1317 (N_1317,N_903,N_896);
and U1318 (N_1318,N_638,N_88);
and U1319 (N_1319,N_12,N_465);
nand U1320 (N_1320,N_835,N_608);
nand U1321 (N_1321,N_193,N_65);
nor U1322 (N_1322,N_253,N_134);
and U1323 (N_1323,N_704,N_444);
or U1324 (N_1324,N_846,N_116);
or U1325 (N_1325,N_321,N_973);
or U1326 (N_1326,N_33,N_283);
and U1327 (N_1327,N_713,N_919);
or U1328 (N_1328,N_496,N_371);
nor U1329 (N_1329,N_451,N_943);
and U1330 (N_1330,N_505,N_657);
nor U1331 (N_1331,N_464,N_507);
or U1332 (N_1332,N_423,N_25);
or U1333 (N_1333,N_105,N_0);
or U1334 (N_1334,N_652,N_803);
nand U1335 (N_1335,N_359,N_198);
and U1336 (N_1336,N_773,N_85);
nand U1337 (N_1337,N_244,N_755);
nor U1338 (N_1338,N_333,N_458);
or U1339 (N_1339,N_787,N_80);
nor U1340 (N_1340,N_257,N_609);
or U1341 (N_1341,N_306,N_237);
or U1342 (N_1342,N_649,N_849);
and U1343 (N_1343,N_599,N_240);
nand U1344 (N_1344,N_335,N_752);
nor U1345 (N_1345,N_891,N_238);
nand U1346 (N_1346,N_220,N_936);
or U1347 (N_1347,N_565,N_315);
or U1348 (N_1348,N_664,N_418);
nand U1349 (N_1349,N_912,N_762);
or U1350 (N_1350,N_941,N_831);
nand U1351 (N_1351,N_358,N_293);
nand U1352 (N_1352,N_596,N_527);
or U1353 (N_1353,N_208,N_521);
nand U1354 (N_1354,N_232,N_692);
xor U1355 (N_1355,N_518,N_329);
or U1356 (N_1356,N_161,N_687);
or U1357 (N_1357,N_900,N_120);
nand U1358 (N_1358,N_529,N_49);
or U1359 (N_1359,N_194,N_94);
or U1360 (N_1360,N_781,N_404);
nand U1361 (N_1361,N_52,N_420);
xor U1362 (N_1362,N_894,N_855);
and U1363 (N_1363,N_790,N_40);
nand U1364 (N_1364,N_508,N_636);
or U1365 (N_1365,N_644,N_179);
or U1366 (N_1366,N_544,N_54);
and U1367 (N_1367,N_586,N_735);
or U1368 (N_1368,N_633,N_679);
or U1369 (N_1369,N_615,N_360);
nand U1370 (N_1370,N_745,N_384);
nor U1371 (N_1371,N_475,N_797);
or U1372 (N_1372,N_815,N_726);
and U1373 (N_1373,N_201,N_472);
nand U1374 (N_1374,N_605,N_542);
xnor U1375 (N_1375,N_3,N_789);
or U1376 (N_1376,N_66,N_204);
nor U1377 (N_1377,N_101,N_86);
and U1378 (N_1378,N_779,N_18);
nor U1379 (N_1379,N_700,N_270);
and U1380 (N_1380,N_279,N_114);
or U1381 (N_1381,N_895,N_645);
and U1382 (N_1382,N_651,N_119);
and U1383 (N_1383,N_233,N_195);
or U1384 (N_1384,N_337,N_760);
nor U1385 (N_1385,N_58,N_191);
nand U1386 (N_1386,N_681,N_592);
and U1387 (N_1387,N_15,N_512);
nand U1388 (N_1388,N_830,N_148);
and U1389 (N_1389,N_709,N_215);
or U1390 (N_1390,N_290,N_151);
nor U1391 (N_1391,N_51,N_376);
nand U1392 (N_1392,N_697,N_251);
xnor U1393 (N_1393,N_254,N_158);
and U1394 (N_1394,N_832,N_777);
or U1395 (N_1395,N_540,N_619);
nand U1396 (N_1396,N_304,N_515);
or U1397 (N_1397,N_574,N_490);
xor U1398 (N_1398,N_686,N_280);
or U1399 (N_1399,N_668,N_989);
nand U1400 (N_1400,N_372,N_491);
nor U1401 (N_1401,N_379,N_990);
and U1402 (N_1402,N_965,N_354);
nand U1403 (N_1403,N_878,N_627);
or U1404 (N_1404,N_724,N_711);
and U1405 (N_1405,N_506,N_572);
and U1406 (N_1406,N_87,N_646);
nor U1407 (N_1407,N_126,N_440);
and U1408 (N_1408,N_388,N_128);
and U1409 (N_1409,N_823,N_217);
nor U1410 (N_1410,N_20,N_690);
nand U1411 (N_1411,N_890,N_847);
nand U1412 (N_1412,N_814,N_112);
nand U1413 (N_1413,N_416,N_212);
and U1414 (N_1414,N_171,N_165);
and U1415 (N_1415,N_402,N_567);
nor U1416 (N_1416,N_920,N_571);
nor U1417 (N_1417,N_923,N_513);
nand U1418 (N_1418,N_250,N_452);
or U1419 (N_1419,N_688,N_933);
and U1420 (N_1420,N_793,N_281);
or U1421 (N_1421,N_622,N_867);
xnor U1422 (N_1422,N_109,N_453);
and U1423 (N_1423,N_340,N_581);
nor U1424 (N_1424,N_634,N_898);
and U1425 (N_1425,N_341,N_821);
nand U1426 (N_1426,N_682,N_607);
nor U1427 (N_1427,N_226,N_363);
or U1428 (N_1428,N_584,N_303);
nor U1429 (N_1429,N_95,N_860);
nand U1430 (N_1430,N_412,N_999);
nor U1431 (N_1431,N_524,N_580);
and U1432 (N_1432,N_778,N_578);
and U1433 (N_1433,N_998,N_241);
nor U1434 (N_1434,N_278,N_144);
nor U1435 (N_1435,N_424,N_267);
nor U1436 (N_1436,N_532,N_287);
or U1437 (N_1437,N_480,N_556);
or U1438 (N_1438,N_462,N_147);
or U1439 (N_1439,N_96,N_541);
xor U1440 (N_1440,N_985,N_34);
or U1441 (N_1441,N_263,N_77);
nand U1442 (N_1442,N_531,N_788);
or U1443 (N_1443,N_323,N_378);
nand U1444 (N_1444,N_272,N_623);
nor U1445 (N_1445,N_487,N_757);
nand U1446 (N_1446,N_510,N_813);
nand U1447 (N_1447,N_494,N_349);
or U1448 (N_1448,N_295,N_76);
and U1449 (N_1449,N_169,N_733);
and U1450 (N_1450,N_561,N_182);
nor U1451 (N_1451,N_300,N_247);
nor U1452 (N_1452,N_702,N_694);
nand U1453 (N_1453,N_926,N_155);
or U1454 (N_1454,N_678,N_401);
or U1455 (N_1455,N_616,N_997);
or U1456 (N_1456,N_291,N_871);
nand U1457 (N_1457,N_642,N_482);
and U1458 (N_1458,N_24,N_59);
and U1459 (N_1459,N_969,N_840);
and U1460 (N_1460,N_443,N_802);
or U1461 (N_1461,N_693,N_701);
and U1462 (N_1462,N_523,N_229);
and U1463 (N_1463,N_585,N_218);
or U1464 (N_1464,N_99,N_7);
and U1465 (N_1465,N_46,N_429);
nand U1466 (N_1466,N_766,N_434);
nor U1467 (N_1467,N_55,N_260);
nand U1468 (N_1468,N_117,N_710);
or U1469 (N_1469,N_72,N_78);
and U1470 (N_1470,N_342,N_562);
and U1471 (N_1471,N_987,N_854);
or U1472 (N_1472,N_224,N_988);
nand U1473 (N_1473,N_837,N_32);
nand U1474 (N_1474,N_197,N_977);
xor U1475 (N_1475,N_345,N_428);
nor U1476 (N_1476,N_248,N_739);
nand U1477 (N_1477,N_728,N_139);
nor U1478 (N_1478,N_178,N_430);
nand U1479 (N_1479,N_391,N_137);
nand U1480 (N_1480,N_911,N_225);
nand U1481 (N_1481,N_14,N_904);
and U1482 (N_1482,N_864,N_727);
nand U1483 (N_1483,N_786,N_30);
or U1484 (N_1484,N_958,N_501);
nor U1485 (N_1485,N_984,N_203);
nand U1486 (N_1486,N_108,N_153);
or U1487 (N_1487,N_262,N_310);
xor U1488 (N_1488,N_392,N_509);
nor U1489 (N_1489,N_469,N_62);
and U1490 (N_1490,N_45,N_381);
nor U1491 (N_1491,N_881,N_715);
nand U1492 (N_1492,N_929,N_228);
nor U1493 (N_1493,N_880,N_214);
or U1494 (N_1494,N_972,N_872);
or U1495 (N_1495,N_200,N_450);
nand U1496 (N_1496,N_405,N_922);
or U1497 (N_1497,N_748,N_886);
nor U1498 (N_1498,N_843,N_460);
and U1499 (N_1499,N_246,N_683);
nor U1500 (N_1500,N_714,N_673);
and U1501 (N_1501,N_87,N_924);
nand U1502 (N_1502,N_836,N_954);
and U1503 (N_1503,N_963,N_858);
and U1504 (N_1504,N_466,N_514);
nand U1505 (N_1505,N_67,N_322);
and U1506 (N_1506,N_989,N_672);
nor U1507 (N_1507,N_210,N_650);
or U1508 (N_1508,N_512,N_975);
and U1509 (N_1509,N_306,N_808);
and U1510 (N_1510,N_256,N_420);
and U1511 (N_1511,N_359,N_439);
and U1512 (N_1512,N_6,N_92);
and U1513 (N_1513,N_819,N_1);
or U1514 (N_1514,N_877,N_758);
nor U1515 (N_1515,N_58,N_296);
nor U1516 (N_1516,N_200,N_615);
nor U1517 (N_1517,N_175,N_922);
and U1518 (N_1518,N_23,N_705);
nor U1519 (N_1519,N_857,N_69);
and U1520 (N_1520,N_31,N_550);
nor U1521 (N_1521,N_159,N_517);
xor U1522 (N_1522,N_81,N_862);
nor U1523 (N_1523,N_412,N_260);
and U1524 (N_1524,N_807,N_872);
or U1525 (N_1525,N_933,N_833);
or U1526 (N_1526,N_330,N_248);
nor U1527 (N_1527,N_138,N_800);
nand U1528 (N_1528,N_28,N_375);
nor U1529 (N_1529,N_546,N_640);
and U1530 (N_1530,N_481,N_173);
nand U1531 (N_1531,N_878,N_102);
and U1532 (N_1532,N_354,N_727);
and U1533 (N_1533,N_958,N_557);
nor U1534 (N_1534,N_323,N_288);
and U1535 (N_1535,N_100,N_338);
nand U1536 (N_1536,N_292,N_855);
nor U1537 (N_1537,N_409,N_814);
and U1538 (N_1538,N_237,N_36);
or U1539 (N_1539,N_490,N_332);
or U1540 (N_1540,N_18,N_144);
or U1541 (N_1541,N_189,N_66);
nand U1542 (N_1542,N_252,N_528);
and U1543 (N_1543,N_470,N_214);
and U1544 (N_1544,N_878,N_937);
and U1545 (N_1545,N_495,N_333);
nor U1546 (N_1546,N_124,N_549);
nor U1547 (N_1547,N_823,N_29);
and U1548 (N_1548,N_594,N_98);
nor U1549 (N_1549,N_699,N_226);
or U1550 (N_1550,N_138,N_574);
nor U1551 (N_1551,N_666,N_833);
or U1552 (N_1552,N_68,N_794);
and U1553 (N_1553,N_357,N_55);
or U1554 (N_1554,N_498,N_108);
and U1555 (N_1555,N_434,N_390);
nor U1556 (N_1556,N_442,N_209);
or U1557 (N_1557,N_440,N_296);
and U1558 (N_1558,N_45,N_37);
and U1559 (N_1559,N_718,N_435);
nand U1560 (N_1560,N_827,N_124);
and U1561 (N_1561,N_81,N_380);
nor U1562 (N_1562,N_212,N_626);
or U1563 (N_1563,N_393,N_277);
nor U1564 (N_1564,N_422,N_137);
nand U1565 (N_1565,N_803,N_934);
nand U1566 (N_1566,N_279,N_430);
or U1567 (N_1567,N_959,N_807);
nand U1568 (N_1568,N_452,N_71);
and U1569 (N_1569,N_405,N_432);
and U1570 (N_1570,N_196,N_754);
xor U1571 (N_1571,N_764,N_611);
nor U1572 (N_1572,N_270,N_903);
nor U1573 (N_1573,N_347,N_659);
xor U1574 (N_1574,N_144,N_564);
and U1575 (N_1575,N_364,N_713);
nand U1576 (N_1576,N_182,N_495);
nand U1577 (N_1577,N_696,N_590);
nand U1578 (N_1578,N_976,N_578);
nor U1579 (N_1579,N_113,N_571);
and U1580 (N_1580,N_787,N_127);
nand U1581 (N_1581,N_285,N_929);
nand U1582 (N_1582,N_406,N_3);
or U1583 (N_1583,N_470,N_366);
nand U1584 (N_1584,N_424,N_648);
or U1585 (N_1585,N_571,N_694);
nor U1586 (N_1586,N_199,N_541);
nand U1587 (N_1587,N_28,N_411);
nor U1588 (N_1588,N_709,N_736);
nor U1589 (N_1589,N_933,N_422);
nor U1590 (N_1590,N_639,N_700);
or U1591 (N_1591,N_941,N_715);
or U1592 (N_1592,N_908,N_198);
nand U1593 (N_1593,N_913,N_34);
or U1594 (N_1594,N_363,N_753);
or U1595 (N_1595,N_845,N_401);
or U1596 (N_1596,N_61,N_761);
or U1597 (N_1597,N_573,N_334);
or U1598 (N_1598,N_188,N_631);
nor U1599 (N_1599,N_623,N_891);
nor U1600 (N_1600,N_332,N_833);
and U1601 (N_1601,N_214,N_751);
nand U1602 (N_1602,N_448,N_366);
and U1603 (N_1603,N_736,N_176);
nor U1604 (N_1604,N_105,N_135);
and U1605 (N_1605,N_858,N_483);
nand U1606 (N_1606,N_885,N_775);
nor U1607 (N_1607,N_162,N_56);
or U1608 (N_1608,N_174,N_190);
xnor U1609 (N_1609,N_184,N_829);
xor U1610 (N_1610,N_650,N_106);
nor U1611 (N_1611,N_157,N_281);
or U1612 (N_1612,N_640,N_779);
and U1613 (N_1613,N_395,N_25);
nor U1614 (N_1614,N_858,N_491);
nand U1615 (N_1615,N_456,N_104);
nand U1616 (N_1616,N_378,N_212);
nand U1617 (N_1617,N_458,N_474);
and U1618 (N_1618,N_898,N_528);
nand U1619 (N_1619,N_45,N_503);
nand U1620 (N_1620,N_47,N_911);
and U1621 (N_1621,N_800,N_483);
nand U1622 (N_1622,N_85,N_675);
nor U1623 (N_1623,N_724,N_933);
or U1624 (N_1624,N_857,N_992);
nand U1625 (N_1625,N_711,N_654);
or U1626 (N_1626,N_642,N_418);
nor U1627 (N_1627,N_977,N_430);
or U1628 (N_1628,N_500,N_318);
nand U1629 (N_1629,N_843,N_487);
xor U1630 (N_1630,N_946,N_5);
nand U1631 (N_1631,N_340,N_733);
nor U1632 (N_1632,N_425,N_340);
and U1633 (N_1633,N_940,N_704);
nor U1634 (N_1634,N_736,N_158);
nor U1635 (N_1635,N_722,N_476);
and U1636 (N_1636,N_854,N_812);
nand U1637 (N_1637,N_955,N_424);
xor U1638 (N_1638,N_144,N_34);
or U1639 (N_1639,N_89,N_894);
and U1640 (N_1640,N_768,N_806);
nand U1641 (N_1641,N_485,N_539);
nand U1642 (N_1642,N_632,N_352);
nor U1643 (N_1643,N_280,N_616);
nand U1644 (N_1644,N_585,N_848);
nand U1645 (N_1645,N_673,N_556);
or U1646 (N_1646,N_52,N_151);
or U1647 (N_1647,N_467,N_431);
nor U1648 (N_1648,N_366,N_865);
and U1649 (N_1649,N_321,N_732);
nor U1650 (N_1650,N_148,N_39);
or U1651 (N_1651,N_197,N_474);
nor U1652 (N_1652,N_147,N_635);
xnor U1653 (N_1653,N_206,N_565);
or U1654 (N_1654,N_994,N_296);
nor U1655 (N_1655,N_232,N_121);
nand U1656 (N_1656,N_357,N_399);
and U1657 (N_1657,N_996,N_310);
nor U1658 (N_1658,N_871,N_832);
nand U1659 (N_1659,N_465,N_391);
nor U1660 (N_1660,N_234,N_630);
and U1661 (N_1661,N_968,N_570);
nor U1662 (N_1662,N_85,N_77);
and U1663 (N_1663,N_901,N_436);
nor U1664 (N_1664,N_983,N_637);
nor U1665 (N_1665,N_261,N_382);
nor U1666 (N_1666,N_622,N_795);
and U1667 (N_1667,N_259,N_266);
nand U1668 (N_1668,N_212,N_827);
nand U1669 (N_1669,N_747,N_622);
nand U1670 (N_1670,N_974,N_956);
xor U1671 (N_1671,N_713,N_635);
or U1672 (N_1672,N_524,N_238);
nand U1673 (N_1673,N_344,N_573);
nor U1674 (N_1674,N_512,N_634);
and U1675 (N_1675,N_805,N_460);
and U1676 (N_1676,N_357,N_836);
or U1677 (N_1677,N_487,N_734);
nor U1678 (N_1678,N_425,N_48);
and U1679 (N_1679,N_752,N_548);
or U1680 (N_1680,N_833,N_787);
nor U1681 (N_1681,N_91,N_996);
nor U1682 (N_1682,N_978,N_484);
or U1683 (N_1683,N_476,N_213);
or U1684 (N_1684,N_919,N_694);
or U1685 (N_1685,N_872,N_588);
or U1686 (N_1686,N_814,N_192);
nand U1687 (N_1687,N_63,N_389);
nand U1688 (N_1688,N_197,N_985);
nand U1689 (N_1689,N_772,N_455);
and U1690 (N_1690,N_659,N_881);
xor U1691 (N_1691,N_194,N_372);
or U1692 (N_1692,N_781,N_100);
and U1693 (N_1693,N_313,N_781);
and U1694 (N_1694,N_583,N_781);
or U1695 (N_1695,N_640,N_167);
or U1696 (N_1696,N_364,N_1);
or U1697 (N_1697,N_631,N_342);
and U1698 (N_1698,N_182,N_932);
and U1699 (N_1699,N_414,N_268);
and U1700 (N_1700,N_258,N_869);
nor U1701 (N_1701,N_49,N_200);
nand U1702 (N_1702,N_636,N_728);
and U1703 (N_1703,N_578,N_255);
or U1704 (N_1704,N_129,N_789);
or U1705 (N_1705,N_795,N_894);
nand U1706 (N_1706,N_335,N_990);
or U1707 (N_1707,N_707,N_166);
nor U1708 (N_1708,N_180,N_389);
xor U1709 (N_1709,N_77,N_286);
nand U1710 (N_1710,N_941,N_945);
nor U1711 (N_1711,N_31,N_703);
nand U1712 (N_1712,N_594,N_617);
nor U1713 (N_1713,N_512,N_254);
xor U1714 (N_1714,N_145,N_277);
nand U1715 (N_1715,N_365,N_806);
or U1716 (N_1716,N_617,N_581);
nand U1717 (N_1717,N_128,N_439);
nor U1718 (N_1718,N_691,N_805);
nand U1719 (N_1719,N_479,N_610);
nand U1720 (N_1720,N_159,N_242);
nand U1721 (N_1721,N_785,N_252);
nand U1722 (N_1722,N_94,N_834);
nor U1723 (N_1723,N_236,N_336);
nor U1724 (N_1724,N_901,N_76);
nor U1725 (N_1725,N_803,N_660);
and U1726 (N_1726,N_321,N_70);
or U1727 (N_1727,N_89,N_216);
or U1728 (N_1728,N_217,N_443);
or U1729 (N_1729,N_735,N_62);
or U1730 (N_1730,N_621,N_188);
nor U1731 (N_1731,N_493,N_486);
nand U1732 (N_1732,N_924,N_955);
nand U1733 (N_1733,N_846,N_408);
or U1734 (N_1734,N_969,N_550);
nor U1735 (N_1735,N_892,N_497);
or U1736 (N_1736,N_274,N_0);
nand U1737 (N_1737,N_729,N_762);
nor U1738 (N_1738,N_631,N_175);
nand U1739 (N_1739,N_327,N_734);
nor U1740 (N_1740,N_689,N_763);
nor U1741 (N_1741,N_692,N_454);
and U1742 (N_1742,N_625,N_546);
or U1743 (N_1743,N_463,N_883);
and U1744 (N_1744,N_614,N_500);
nand U1745 (N_1745,N_724,N_857);
nor U1746 (N_1746,N_678,N_488);
and U1747 (N_1747,N_920,N_108);
nand U1748 (N_1748,N_92,N_862);
and U1749 (N_1749,N_229,N_461);
nor U1750 (N_1750,N_573,N_385);
and U1751 (N_1751,N_236,N_324);
or U1752 (N_1752,N_10,N_441);
nand U1753 (N_1753,N_578,N_336);
and U1754 (N_1754,N_885,N_500);
or U1755 (N_1755,N_32,N_728);
nor U1756 (N_1756,N_966,N_887);
nor U1757 (N_1757,N_176,N_529);
and U1758 (N_1758,N_973,N_661);
or U1759 (N_1759,N_785,N_494);
or U1760 (N_1760,N_55,N_296);
or U1761 (N_1761,N_156,N_128);
nand U1762 (N_1762,N_869,N_844);
nand U1763 (N_1763,N_713,N_339);
and U1764 (N_1764,N_247,N_647);
or U1765 (N_1765,N_496,N_75);
or U1766 (N_1766,N_964,N_617);
and U1767 (N_1767,N_205,N_519);
and U1768 (N_1768,N_907,N_545);
and U1769 (N_1769,N_322,N_336);
nand U1770 (N_1770,N_237,N_12);
and U1771 (N_1771,N_684,N_151);
nand U1772 (N_1772,N_241,N_79);
or U1773 (N_1773,N_611,N_984);
nor U1774 (N_1774,N_54,N_773);
or U1775 (N_1775,N_961,N_162);
or U1776 (N_1776,N_816,N_629);
xor U1777 (N_1777,N_870,N_468);
and U1778 (N_1778,N_394,N_447);
nor U1779 (N_1779,N_565,N_120);
or U1780 (N_1780,N_244,N_745);
and U1781 (N_1781,N_574,N_720);
and U1782 (N_1782,N_50,N_753);
nor U1783 (N_1783,N_378,N_466);
nand U1784 (N_1784,N_208,N_75);
nand U1785 (N_1785,N_267,N_569);
nor U1786 (N_1786,N_137,N_225);
and U1787 (N_1787,N_831,N_114);
or U1788 (N_1788,N_4,N_758);
or U1789 (N_1789,N_358,N_703);
nor U1790 (N_1790,N_322,N_413);
xnor U1791 (N_1791,N_398,N_338);
nand U1792 (N_1792,N_672,N_10);
or U1793 (N_1793,N_200,N_156);
nor U1794 (N_1794,N_130,N_426);
or U1795 (N_1795,N_481,N_558);
or U1796 (N_1796,N_439,N_658);
nand U1797 (N_1797,N_764,N_35);
xor U1798 (N_1798,N_399,N_490);
or U1799 (N_1799,N_186,N_741);
nor U1800 (N_1800,N_967,N_49);
or U1801 (N_1801,N_894,N_762);
and U1802 (N_1802,N_272,N_854);
nor U1803 (N_1803,N_907,N_198);
xor U1804 (N_1804,N_131,N_11);
nor U1805 (N_1805,N_841,N_176);
nand U1806 (N_1806,N_252,N_651);
nor U1807 (N_1807,N_29,N_291);
or U1808 (N_1808,N_298,N_708);
nand U1809 (N_1809,N_72,N_115);
and U1810 (N_1810,N_442,N_32);
nor U1811 (N_1811,N_757,N_528);
nand U1812 (N_1812,N_363,N_27);
and U1813 (N_1813,N_358,N_295);
and U1814 (N_1814,N_151,N_827);
nor U1815 (N_1815,N_626,N_607);
or U1816 (N_1816,N_718,N_514);
nand U1817 (N_1817,N_344,N_513);
or U1818 (N_1818,N_154,N_755);
nand U1819 (N_1819,N_546,N_179);
and U1820 (N_1820,N_606,N_162);
or U1821 (N_1821,N_779,N_698);
or U1822 (N_1822,N_550,N_288);
nand U1823 (N_1823,N_268,N_138);
nor U1824 (N_1824,N_376,N_728);
nor U1825 (N_1825,N_25,N_324);
nor U1826 (N_1826,N_899,N_404);
or U1827 (N_1827,N_978,N_551);
xnor U1828 (N_1828,N_881,N_703);
nor U1829 (N_1829,N_734,N_265);
nand U1830 (N_1830,N_115,N_615);
and U1831 (N_1831,N_424,N_488);
nor U1832 (N_1832,N_733,N_468);
nor U1833 (N_1833,N_242,N_18);
or U1834 (N_1834,N_698,N_709);
nor U1835 (N_1835,N_750,N_614);
nand U1836 (N_1836,N_350,N_700);
nor U1837 (N_1837,N_719,N_153);
or U1838 (N_1838,N_836,N_414);
or U1839 (N_1839,N_567,N_513);
or U1840 (N_1840,N_598,N_450);
or U1841 (N_1841,N_956,N_882);
nor U1842 (N_1842,N_171,N_872);
nand U1843 (N_1843,N_785,N_653);
nor U1844 (N_1844,N_172,N_3);
nand U1845 (N_1845,N_365,N_855);
nand U1846 (N_1846,N_65,N_912);
or U1847 (N_1847,N_917,N_340);
nand U1848 (N_1848,N_456,N_331);
or U1849 (N_1849,N_330,N_723);
nor U1850 (N_1850,N_278,N_281);
nand U1851 (N_1851,N_208,N_722);
or U1852 (N_1852,N_468,N_485);
nor U1853 (N_1853,N_54,N_403);
or U1854 (N_1854,N_695,N_703);
nand U1855 (N_1855,N_129,N_741);
nor U1856 (N_1856,N_529,N_920);
nor U1857 (N_1857,N_310,N_789);
nor U1858 (N_1858,N_757,N_611);
nand U1859 (N_1859,N_975,N_372);
nor U1860 (N_1860,N_577,N_273);
nor U1861 (N_1861,N_761,N_377);
and U1862 (N_1862,N_634,N_811);
and U1863 (N_1863,N_418,N_500);
or U1864 (N_1864,N_765,N_421);
and U1865 (N_1865,N_479,N_831);
nand U1866 (N_1866,N_469,N_916);
or U1867 (N_1867,N_642,N_562);
nand U1868 (N_1868,N_585,N_770);
nand U1869 (N_1869,N_883,N_859);
nand U1870 (N_1870,N_887,N_335);
nor U1871 (N_1871,N_916,N_606);
or U1872 (N_1872,N_714,N_882);
nand U1873 (N_1873,N_739,N_383);
nor U1874 (N_1874,N_401,N_600);
and U1875 (N_1875,N_39,N_196);
nand U1876 (N_1876,N_627,N_753);
nor U1877 (N_1877,N_759,N_465);
nor U1878 (N_1878,N_113,N_939);
and U1879 (N_1879,N_31,N_197);
nor U1880 (N_1880,N_119,N_516);
or U1881 (N_1881,N_794,N_74);
or U1882 (N_1882,N_61,N_402);
nor U1883 (N_1883,N_734,N_288);
or U1884 (N_1884,N_912,N_721);
and U1885 (N_1885,N_201,N_489);
or U1886 (N_1886,N_844,N_551);
and U1887 (N_1887,N_24,N_872);
or U1888 (N_1888,N_595,N_494);
nand U1889 (N_1889,N_265,N_498);
and U1890 (N_1890,N_904,N_470);
nand U1891 (N_1891,N_351,N_660);
or U1892 (N_1892,N_168,N_100);
and U1893 (N_1893,N_786,N_274);
or U1894 (N_1894,N_321,N_968);
nand U1895 (N_1895,N_108,N_500);
nor U1896 (N_1896,N_181,N_752);
nor U1897 (N_1897,N_441,N_223);
nor U1898 (N_1898,N_631,N_964);
and U1899 (N_1899,N_20,N_850);
or U1900 (N_1900,N_120,N_598);
nor U1901 (N_1901,N_350,N_939);
nand U1902 (N_1902,N_256,N_489);
and U1903 (N_1903,N_462,N_443);
and U1904 (N_1904,N_178,N_391);
nor U1905 (N_1905,N_100,N_297);
nand U1906 (N_1906,N_451,N_223);
nand U1907 (N_1907,N_87,N_793);
and U1908 (N_1908,N_487,N_111);
and U1909 (N_1909,N_881,N_98);
nor U1910 (N_1910,N_973,N_550);
nor U1911 (N_1911,N_31,N_45);
nand U1912 (N_1912,N_186,N_386);
nor U1913 (N_1913,N_720,N_338);
or U1914 (N_1914,N_530,N_620);
xnor U1915 (N_1915,N_893,N_227);
nor U1916 (N_1916,N_375,N_689);
nor U1917 (N_1917,N_67,N_86);
or U1918 (N_1918,N_456,N_130);
nor U1919 (N_1919,N_3,N_931);
nand U1920 (N_1920,N_903,N_82);
nor U1921 (N_1921,N_270,N_383);
nor U1922 (N_1922,N_5,N_246);
or U1923 (N_1923,N_347,N_960);
and U1924 (N_1924,N_98,N_217);
nor U1925 (N_1925,N_156,N_410);
and U1926 (N_1926,N_458,N_890);
and U1927 (N_1927,N_784,N_848);
nor U1928 (N_1928,N_730,N_15);
nor U1929 (N_1929,N_765,N_785);
nor U1930 (N_1930,N_289,N_676);
and U1931 (N_1931,N_455,N_921);
nand U1932 (N_1932,N_7,N_845);
or U1933 (N_1933,N_535,N_516);
and U1934 (N_1934,N_6,N_880);
and U1935 (N_1935,N_529,N_827);
nand U1936 (N_1936,N_275,N_63);
and U1937 (N_1937,N_179,N_405);
nor U1938 (N_1938,N_977,N_320);
nand U1939 (N_1939,N_946,N_381);
or U1940 (N_1940,N_398,N_385);
or U1941 (N_1941,N_752,N_720);
and U1942 (N_1942,N_550,N_783);
and U1943 (N_1943,N_770,N_192);
xor U1944 (N_1944,N_300,N_905);
or U1945 (N_1945,N_870,N_163);
xor U1946 (N_1946,N_412,N_294);
and U1947 (N_1947,N_328,N_157);
nor U1948 (N_1948,N_615,N_62);
and U1949 (N_1949,N_908,N_210);
and U1950 (N_1950,N_538,N_422);
or U1951 (N_1951,N_93,N_886);
or U1952 (N_1952,N_730,N_695);
and U1953 (N_1953,N_785,N_423);
nand U1954 (N_1954,N_603,N_343);
or U1955 (N_1955,N_510,N_424);
and U1956 (N_1956,N_616,N_259);
and U1957 (N_1957,N_852,N_862);
or U1958 (N_1958,N_132,N_33);
and U1959 (N_1959,N_979,N_814);
nand U1960 (N_1960,N_86,N_688);
nor U1961 (N_1961,N_55,N_397);
nor U1962 (N_1962,N_972,N_579);
nand U1963 (N_1963,N_631,N_123);
nor U1964 (N_1964,N_829,N_598);
nor U1965 (N_1965,N_213,N_736);
nand U1966 (N_1966,N_295,N_639);
nand U1967 (N_1967,N_680,N_914);
nand U1968 (N_1968,N_974,N_749);
nand U1969 (N_1969,N_524,N_640);
and U1970 (N_1970,N_763,N_829);
or U1971 (N_1971,N_445,N_596);
nor U1972 (N_1972,N_842,N_897);
nor U1973 (N_1973,N_730,N_64);
or U1974 (N_1974,N_446,N_807);
or U1975 (N_1975,N_764,N_614);
and U1976 (N_1976,N_602,N_485);
nor U1977 (N_1977,N_345,N_538);
and U1978 (N_1978,N_714,N_104);
or U1979 (N_1979,N_904,N_207);
nand U1980 (N_1980,N_176,N_744);
xnor U1981 (N_1981,N_400,N_646);
or U1982 (N_1982,N_732,N_90);
nor U1983 (N_1983,N_276,N_853);
or U1984 (N_1984,N_624,N_798);
xnor U1985 (N_1985,N_189,N_492);
or U1986 (N_1986,N_175,N_303);
and U1987 (N_1987,N_216,N_717);
or U1988 (N_1988,N_735,N_423);
and U1989 (N_1989,N_858,N_198);
nor U1990 (N_1990,N_781,N_978);
nor U1991 (N_1991,N_833,N_86);
nor U1992 (N_1992,N_639,N_745);
or U1993 (N_1993,N_993,N_850);
nor U1994 (N_1994,N_964,N_794);
and U1995 (N_1995,N_848,N_202);
or U1996 (N_1996,N_322,N_147);
nand U1997 (N_1997,N_40,N_755);
nand U1998 (N_1998,N_928,N_629);
nor U1999 (N_1999,N_548,N_321);
nand U2000 (N_2000,N_1010,N_1141);
and U2001 (N_2001,N_1035,N_1799);
or U2002 (N_2002,N_1507,N_1774);
nand U2003 (N_2003,N_1629,N_1715);
and U2004 (N_2004,N_1592,N_1265);
or U2005 (N_2005,N_1742,N_1990);
nand U2006 (N_2006,N_1546,N_1946);
or U2007 (N_2007,N_1430,N_1133);
nor U2008 (N_2008,N_1739,N_1608);
nor U2009 (N_2009,N_1471,N_1517);
and U2010 (N_2010,N_1692,N_1709);
and U2011 (N_2011,N_1037,N_1444);
nand U2012 (N_2012,N_1938,N_1842);
nand U2013 (N_2013,N_1802,N_1058);
nand U2014 (N_2014,N_1260,N_1482);
nor U2015 (N_2015,N_1122,N_1636);
nand U2016 (N_2016,N_1441,N_1987);
and U2017 (N_2017,N_1603,N_1902);
nor U2018 (N_2018,N_1660,N_1810);
nand U2019 (N_2019,N_1247,N_1601);
nand U2020 (N_2020,N_1648,N_1250);
or U2021 (N_2021,N_1824,N_1169);
or U2022 (N_2022,N_1940,N_1955);
nor U2023 (N_2023,N_1489,N_1433);
or U2024 (N_2024,N_1099,N_1459);
nand U2025 (N_2025,N_1670,N_1594);
or U2026 (N_2026,N_1664,N_1532);
and U2027 (N_2027,N_1080,N_1869);
or U2028 (N_2028,N_1610,N_1981);
and U2029 (N_2029,N_1148,N_1278);
or U2030 (N_2030,N_1182,N_1368);
nor U2031 (N_2031,N_1666,N_1496);
nor U2032 (N_2032,N_1092,N_1720);
nor U2033 (N_2033,N_1284,N_1324);
or U2034 (N_2034,N_1781,N_1402);
nor U2035 (N_2035,N_1397,N_1046);
nand U2036 (N_2036,N_1014,N_1374);
nor U2037 (N_2037,N_1944,N_1702);
nor U2038 (N_2038,N_1187,N_1057);
and U2039 (N_2039,N_1039,N_1779);
nand U2040 (N_2040,N_1053,N_1719);
and U2041 (N_2041,N_1729,N_1921);
nand U2042 (N_2042,N_1913,N_1185);
nand U2043 (N_2043,N_1992,N_1412);
nor U2044 (N_2044,N_1645,N_1336);
and U2045 (N_2045,N_1510,N_1366);
or U2046 (N_2046,N_1383,N_1677);
nor U2047 (N_2047,N_1996,N_1595);
nor U2048 (N_2048,N_1661,N_1707);
nor U2049 (N_2049,N_1385,N_1438);
nand U2050 (N_2050,N_1085,N_1375);
nor U2051 (N_2051,N_1146,N_1172);
and U2052 (N_2052,N_1222,N_1686);
nor U2053 (N_2053,N_1695,N_1432);
nor U2054 (N_2054,N_1193,N_1543);
nand U2055 (N_2055,N_1089,N_1463);
nor U2056 (N_2056,N_1223,N_1287);
and U2057 (N_2057,N_1128,N_1115);
and U2058 (N_2058,N_1462,N_1040);
and U2059 (N_2059,N_1490,N_1285);
nand U2060 (N_2060,N_1117,N_1593);
or U2061 (N_2061,N_1120,N_1332);
nand U2062 (N_2062,N_1155,N_1359);
and U2063 (N_2063,N_1018,N_1054);
or U2064 (N_2064,N_1473,N_1088);
nand U2065 (N_2065,N_1371,N_1079);
nor U2066 (N_2066,N_1078,N_1031);
and U2067 (N_2067,N_1678,N_1963);
and U2068 (N_2068,N_1897,N_1620);
and U2069 (N_2069,N_1416,N_1536);
nand U2070 (N_2070,N_1521,N_1047);
and U2071 (N_2071,N_1922,N_1019);
nand U2072 (N_2072,N_1693,N_1884);
nor U2073 (N_2073,N_1920,N_1377);
nor U2074 (N_2074,N_1485,N_1060);
xnor U2075 (N_2075,N_1637,N_1998);
nand U2076 (N_2076,N_1767,N_1007);
nand U2077 (N_2077,N_1290,N_1248);
xnor U2078 (N_2078,N_1134,N_1283);
or U2079 (N_2079,N_1597,N_1343);
nor U2080 (N_2080,N_1043,N_1421);
or U2081 (N_2081,N_1738,N_1221);
nand U2082 (N_2082,N_1795,N_1558);
and U2083 (N_2083,N_1835,N_1952);
and U2084 (N_2084,N_1682,N_1789);
or U2085 (N_2085,N_1360,N_1635);
and U2086 (N_2086,N_1309,N_1062);
nor U2087 (N_2087,N_1737,N_1191);
or U2088 (N_2088,N_1755,N_1964);
and U2089 (N_2089,N_1764,N_1158);
and U2090 (N_2090,N_1991,N_1958);
or U2091 (N_2091,N_1604,N_1560);
or U2092 (N_2092,N_1883,N_1818);
and U2093 (N_2093,N_1206,N_1689);
or U2094 (N_2094,N_1451,N_1492);
nand U2095 (N_2095,N_1863,N_1281);
and U2096 (N_2096,N_1841,N_1184);
and U2097 (N_2097,N_1167,N_1896);
nor U2098 (N_2098,N_1968,N_1082);
or U2099 (N_2099,N_1820,N_1656);
nand U2100 (N_2100,N_1429,N_1937);
or U2101 (N_2101,N_1202,N_1606);
nand U2102 (N_2102,N_1465,N_1044);
nand U2103 (N_2103,N_1993,N_1393);
nand U2104 (N_2104,N_1721,N_1333);
nand U2105 (N_2105,N_1237,N_1026);
xnor U2106 (N_2106,N_1151,N_1346);
and U2107 (N_2107,N_1394,N_1508);
nand U2108 (N_2108,N_1427,N_1551);
nand U2109 (N_2109,N_1400,N_1164);
and U2110 (N_2110,N_1947,N_1272);
and U2111 (N_2111,N_1064,N_1953);
and U2112 (N_2112,N_1559,N_1819);
or U2113 (N_2113,N_1130,N_1114);
nor U2114 (N_2114,N_1590,N_1032);
nor U2115 (N_2115,N_1297,N_1581);
nor U2116 (N_2116,N_1639,N_1143);
nand U2117 (N_2117,N_1973,N_1893);
nor U2118 (N_2118,N_1803,N_1524);
and U2119 (N_2119,N_1984,N_1684);
nor U2120 (N_2120,N_1516,N_1561);
and U2121 (N_2121,N_1618,N_1362);
nor U2122 (N_2122,N_1214,N_1194);
nor U2123 (N_2123,N_1499,N_1912);
nand U2124 (N_2124,N_1527,N_1198);
or U2125 (N_2125,N_1140,N_1259);
and U2126 (N_2126,N_1966,N_1340);
xnor U2127 (N_2127,N_1596,N_1012);
or U2128 (N_2128,N_1780,N_1071);
or U2129 (N_2129,N_1347,N_1887);
or U2130 (N_2130,N_1025,N_1668);
and U2131 (N_2131,N_1541,N_1573);
nand U2132 (N_2132,N_1929,N_1391);
or U2133 (N_2133,N_1305,N_1274);
or U2134 (N_2134,N_1061,N_1915);
nor U2135 (N_2135,N_1483,N_1434);
nand U2136 (N_2136,N_1458,N_1553);
nor U2137 (N_2137,N_1974,N_1049);
or U2138 (N_2138,N_1877,N_1410);
and U2139 (N_2139,N_1226,N_1848);
or U2140 (N_2140,N_1825,N_1150);
and U2141 (N_2141,N_1962,N_1838);
xor U2142 (N_2142,N_1855,N_1584);
nor U2143 (N_2143,N_1399,N_1765);
nand U2144 (N_2144,N_1621,N_1322);
or U2145 (N_2145,N_1854,N_1569);
nor U2146 (N_2146,N_1542,N_1550);
and U2147 (N_2147,N_1022,N_1063);
and U2148 (N_2148,N_1171,N_1997);
or U2149 (N_2149,N_1891,N_1195);
nor U2150 (N_2150,N_1506,N_1667);
nand U2151 (N_2151,N_1116,N_1583);
and U2152 (N_2152,N_1292,N_1706);
nor U2153 (N_2153,N_1724,N_1875);
nand U2154 (N_2154,N_1907,N_1788);
and U2155 (N_2155,N_1228,N_1276);
nand U2156 (N_2156,N_1379,N_1760);
nand U2157 (N_2157,N_1725,N_1727);
or U2158 (N_2158,N_1697,N_1293);
or U2159 (N_2159,N_1833,N_1238);
and U2160 (N_2160,N_1815,N_1509);
or U2161 (N_2161,N_1135,N_1857);
and U2162 (N_2162,N_1520,N_1582);
or U2163 (N_2163,N_1843,N_1055);
or U2164 (N_2164,N_1289,N_1717);
nand U2165 (N_2165,N_1523,N_1578);
and U2166 (N_2166,N_1972,N_1229);
nor U2167 (N_2167,N_1967,N_1005);
nor U2168 (N_2168,N_1392,N_1642);
and U2169 (N_2169,N_1232,N_1980);
nor U2170 (N_2170,N_1793,N_1001);
and U2171 (N_2171,N_1242,N_1933);
nand U2172 (N_2172,N_1943,N_1419);
and U2173 (N_2173,N_1077,N_1251);
or U2174 (N_2174,N_1986,N_1999);
nor U2175 (N_2175,N_1703,N_1280);
nand U2176 (N_2176,N_1249,N_1121);
nand U2177 (N_2177,N_1059,N_1413);
nand U2178 (N_2178,N_1323,N_1839);
nor U2179 (N_2179,N_1207,N_1255);
and U2180 (N_2180,N_1575,N_1978);
or U2181 (N_2181,N_1443,N_1267);
xor U2182 (N_2182,N_1435,N_1196);
and U2183 (N_2183,N_1168,N_1806);
nand U2184 (N_2184,N_1932,N_1052);
nand U2185 (N_2185,N_1270,N_1477);
nor U2186 (N_2186,N_1294,N_1840);
or U2187 (N_2187,N_1562,N_1273);
nand U2188 (N_2188,N_1302,N_1404);
nand U2189 (N_2189,N_1136,N_1622);
nor U2190 (N_2190,N_1812,N_1480);
or U2191 (N_2191,N_1809,N_1328);
nand U2192 (N_2192,N_1565,N_1030);
nor U2193 (N_2193,N_1352,N_1364);
and U2194 (N_2194,N_1740,N_1612);
nand U2195 (N_2195,N_1189,N_1431);
nor U2196 (N_2196,N_1638,N_1256);
nor U2197 (N_2197,N_1448,N_1942);
or U2198 (N_2198,N_1540,N_1488);
and U2199 (N_2199,N_1662,N_1361);
nand U2200 (N_2200,N_1469,N_1501);
or U2201 (N_2201,N_1254,N_1567);
or U2202 (N_2202,N_1500,N_1885);
nor U2203 (N_2203,N_1066,N_1445);
xnor U2204 (N_2204,N_1908,N_1570);
or U2205 (N_2205,N_1036,N_1317);
and U2206 (N_2206,N_1407,N_1977);
nor U2207 (N_2207,N_1801,N_1879);
nand U2208 (N_2208,N_1644,N_1716);
and U2209 (N_2209,N_1205,N_1609);
nand U2210 (N_2210,N_1917,N_1858);
or U2211 (N_2211,N_1827,N_1081);
or U2212 (N_2212,N_1589,N_1425);
nor U2213 (N_2213,N_1466,N_1013);
xor U2214 (N_2214,N_1474,N_1341);
and U2215 (N_2215,N_1663,N_1017);
or U2216 (N_2216,N_1671,N_1950);
and U2217 (N_2217,N_1449,N_1954);
and U2218 (N_2218,N_1310,N_1161);
nor U2219 (N_2219,N_1651,N_1873);
nor U2220 (N_2220,N_1033,N_1023);
nor U2221 (N_2221,N_1188,N_1805);
nand U2222 (N_2222,N_1699,N_1497);
or U2223 (N_2223,N_1514,N_1461);
nand U2224 (N_2224,N_1396,N_1300);
and U2225 (N_2225,N_1734,N_1647);
nor U2226 (N_2226,N_1994,N_1144);
nand U2227 (N_2227,N_1747,N_1787);
and U2228 (N_2228,N_1828,N_1796);
or U2229 (N_2229,N_1041,N_1640);
nand U2230 (N_2230,N_1390,N_1090);
or U2231 (N_2231,N_1102,N_1777);
xor U2232 (N_2232,N_1939,N_1453);
and U2233 (N_2233,N_1487,N_1373);
nand U2234 (N_2234,N_1658,N_1277);
and U2235 (N_2235,N_1166,N_1522);
and U2236 (N_2236,N_1750,N_1535);
nand U2237 (N_2237,N_1288,N_1405);
and U2238 (N_2238,N_1437,N_1985);
and U2239 (N_2239,N_1766,N_1870);
and U2240 (N_2240,N_1100,N_1384);
nand U2241 (N_2241,N_1961,N_1723);
xor U2242 (N_2242,N_1091,N_1547);
or U2243 (N_2243,N_1104,N_1784);
or U2244 (N_2244,N_1528,N_1006);
or U2245 (N_2245,N_1472,N_1674);
nand U2246 (N_2246,N_1587,N_1446);
nor U2247 (N_2247,N_1634,N_1414);
or U2248 (N_2248,N_1538,N_1331);
and U2249 (N_2249,N_1861,N_1586);
and U2250 (N_2250,N_1641,N_1736);
nand U2251 (N_2251,N_1212,N_1756);
or U2252 (N_2252,N_1307,N_1685);
nand U2253 (N_2253,N_1529,N_1512);
or U2254 (N_2254,N_1263,N_1369);
or U2255 (N_2255,N_1452,N_1976);
and U2256 (N_2256,N_1179,N_1983);
or U2257 (N_2257,N_1928,N_1675);
nand U2258 (N_2258,N_1957,N_1086);
and U2259 (N_2259,N_1655,N_1173);
or U2260 (N_2260,N_1710,N_1554);
and U2261 (N_2261,N_1613,N_1113);
nor U2262 (N_2262,N_1890,N_1665);
nand U2263 (N_2263,N_1178,N_1301);
or U2264 (N_2264,N_1881,N_1988);
nor U2265 (N_2265,N_1203,N_1003);
and U2266 (N_2266,N_1852,N_1945);
and U2267 (N_2267,N_1152,N_1252);
nor U2268 (N_2268,N_1856,N_1180);
and U2269 (N_2269,N_1753,N_1979);
nand U2270 (N_2270,N_1970,N_1450);
xnor U2271 (N_2271,N_1577,N_1599);
nand U2272 (N_2272,N_1428,N_1021);
and U2273 (N_2273,N_1325,N_1949);
nand U2274 (N_2274,N_1845,N_1889);
and U2275 (N_2275,N_1770,N_1619);
and U2276 (N_2276,N_1320,N_1817);
nor U2277 (N_2277,N_1365,N_1096);
nor U2278 (N_2278,N_1632,N_1345);
and U2279 (N_2279,N_1264,N_1282);
or U2280 (N_2280,N_1087,N_1681);
and U2281 (N_2281,N_1872,N_1751);
nor U2282 (N_2282,N_1157,N_1775);
nor U2283 (N_2283,N_1306,N_1261);
nor U2284 (N_2284,N_1312,N_1746);
and U2285 (N_2285,N_1935,N_1070);
nand U2286 (N_2286,N_1024,N_1837);
and U2287 (N_2287,N_1145,N_1864);
nand U2288 (N_2288,N_1478,N_1109);
or U2289 (N_2289,N_1515,N_1420);
nand U2290 (N_2290,N_1813,N_1162);
and U2291 (N_2291,N_1201,N_1579);
or U2292 (N_2292,N_1627,N_1042);
nor U2293 (N_2293,N_1778,N_1899);
nand U2294 (N_2294,N_1564,N_1225);
nor U2295 (N_2295,N_1625,N_1349);
nor U2296 (N_2296,N_1235,N_1296);
nor U2297 (N_2297,N_1126,N_1257);
and U2298 (N_2298,N_1726,N_1479);
or U2299 (N_2299,N_1572,N_1163);
nand U2300 (N_2300,N_1909,N_1353);
nor U2301 (N_2301,N_1588,N_1129);
nor U2302 (N_2302,N_1457,N_1672);
and U2303 (N_2303,N_1190,N_1020);
nand U2304 (N_2304,N_1127,N_1916);
or U2305 (N_2305,N_1291,N_1108);
and U2306 (N_2306,N_1823,N_1011);
or U2307 (N_2307,N_1700,N_1050);
nand U2308 (N_2308,N_1519,N_1215);
nand U2309 (N_2309,N_1749,N_1266);
nor U2310 (N_2310,N_1183,N_1069);
or U2311 (N_2311,N_1892,N_1794);
or U2312 (N_2312,N_1376,N_1696);
or U2313 (N_2313,N_1544,N_1904);
nor U2314 (N_2314,N_1722,N_1790);
and U2315 (N_2315,N_1969,N_1243);
nand U2316 (N_2316,N_1192,N_1210);
or U2317 (N_2317,N_1556,N_1357);
and U2318 (N_2318,N_1847,N_1204);
and U2319 (N_2319,N_1800,N_1253);
nand U2320 (N_2320,N_1534,N_1829);
nor U2321 (N_2321,N_1147,N_1028);
nand U2322 (N_2322,N_1244,N_1174);
and U2323 (N_2323,N_1363,N_1093);
nand U2324 (N_2324,N_1084,N_1216);
nand U2325 (N_2325,N_1372,N_1426);
nor U2326 (N_2326,N_1298,N_1111);
nand U2327 (N_2327,N_1866,N_1931);
and U2328 (N_2328,N_1773,N_1918);
nor U2329 (N_2329,N_1549,N_1771);
nand U2330 (N_2330,N_1286,N_1342);
xnor U2331 (N_2331,N_1076,N_1311);
and U2332 (N_2332,N_1768,N_1389);
nand U2333 (N_2333,N_1125,N_1424);
or U2334 (N_2334,N_1808,N_1526);
xor U2335 (N_2335,N_1763,N_1051);
or U2336 (N_2336,N_1844,N_1905);
or U2337 (N_2337,N_1792,N_1495);
and U2338 (N_2338,N_1511,N_1744);
or U2339 (N_2339,N_1350,N_1475);
nand U2340 (N_2340,N_1786,N_1275);
nand U2341 (N_2341,N_1160,N_1387);
or U2342 (N_2342,N_1531,N_1959);
and U2343 (N_2343,N_1901,N_1759);
or U2344 (N_2344,N_1814,N_1073);
nor U2345 (N_2345,N_1447,N_1630);
nor U2346 (N_2346,N_1591,N_1382);
nand U2347 (N_2347,N_1211,N_1505);
nand U2348 (N_2348,N_1851,N_1335);
and U2349 (N_2349,N_1139,N_1075);
nor U2350 (N_2350,N_1712,N_1654);
and U2351 (N_2351,N_1846,N_1914);
and U2352 (N_2352,N_1853,N_1816);
nand U2353 (N_2353,N_1910,N_1611);
nand U2354 (N_2354,N_1628,N_1107);
nand U2355 (N_2355,N_1319,N_1585);
nand U2356 (N_2356,N_1776,N_1791);
nor U2357 (N_2357,N_1455,N_1769);
or U2358 (N_2358,N_1871,N_1924);
or U2359 (N_2359,N_1850,N_1348);
or U2360 (N_2360,N_1308,N_1034);
nand U2361 (N_2361,N_1009,N_1730);
nand U2362 (N_2362,N_1713,N_1690);
nand U2363 (N_2363,N_1548,N_1927);
or U2364 (N_2364,N_1154,N_1874);
and U2365 (N_2365,N_1626,N_1101);
nor U2366 (N_2366,N_1923,N_1498);
nand U2367 (N_2367,N_1315,N_1337);
or U2368 (N_2368,N_1367,N_1240);
nand U2369 (N_2369,N_1209,N_1925);
nand U2370 (N_2370,N_1072,N_1728);
and U2371 (N_2371,N_1423,N_1388);
or U2372 (N_2372,N_1159,N_1200);
or U2373 (N_2373,N_1440,N_1785);
nor U2374 (N_2374,N_1600,N_1068);
and U2375 (N_2375,N_1219,N_1456);
nand U2376 (N_2376,N_1074,N_1408);
nand U2377 (N_2377,N_1934,N_1008);
nor U2378 (N_2378,N_1258,N_1574);
or U2379 (N_2379,N_1502,N_1177);
nand U2380 (N_2380,N_1691,N_1380);
nand U2381 (N_2381,N_1132,N_1355);
nand U2382 (N_2382,N_1330,N_1304);
nor U2383 (N_2383,N_1633,N_1605);
and U2384 (N_2384,N_1381,N_1327);
or U2385 (N_2385,N_1811,N_1580);
nand U2386 (N_2386,N_1227,N_1038);
xnor U2387 (N_2387,N_1454,N_1398);
nand U2388 (N_2388,N_1880,N_1338);
or U2389 (N_2389,N_1643,N_1213);
nor U2390 (N_2390,N_1439,N_1493);
and U2391 (N_2391,N_1231,N_1867);
and U2392 (N_2392,N_1175,N_1862);
or U2393 (N_2393,N_1733,N_1395);
nor U2394 (N_2394,N_1752,N_1262);
or U2395 (N_2395,N_1859,N_1982);
and U2396 (N_2396,N_1906,N_1418);
and U2397 (N_2397,N_1894,N_1743);
nor U2398 (N_2398,N_1926,N_1616);
nor U2399 (N_2399,N_1131,N_1876);
nand U2400 (N_2400,N_1602,N_1110);
or U2401 (N_2401,N_1329,N_1965);
or U2402 (N_2402,N_1002,N_1631);
nor U2403 (N_2403,N_1919,N_1903);
xor U2404 (N_2404,N_1208,N_1732);
nand U2405 (N_2405,N_1748,N_1153);
or U2406 (N_2406,N_1246,N_1659);
nand U2407 (N_2407,N_1941,N_1239);
xor U2408 (N_2408,N_1403,N_1563);
nand U2409 (N_2409,N_1705,N_1236);
nand U2410 (N_2410,N_1518,N_1295);
and U2411 (N_2411,N_1615,N_1783);
or U2412 (N_2412,N_1245,N_1334);
nor U2413 (N_2413,N_1772,N_1411);
and U2414 (N_2414,N_1406,N_1197);
nand U2415 (N_2415,N_1481,N_1149);
nor U2416 (N_2416,N_1165,N_1886);
or U2417 (N_2417,N_1975,N_1545);
and U2418 (N_2418,N_1798,N_1356);
nand U2419 (N_2419,N_1614,N_1936);
or U2420 (N_2420,N_1494,N_1484);
nand U2421 (N_2421,N_1868,N_1989);
and U2422 (N_2422,N_1224,N_1491);
or U2423 (N_2423,N_1436,N_1673);
or U2424 (N_2424,N_1860,N_1401);
nor U2425 (N_2425,N_1220,N_1537);
and U2426 (N_2426,N_1513,N_1878);
or U2427 (N_2427,N_1468,N_1470);
nor U2428 (N_2428,N_1711,N_1676);
and U2429 (N_2429,N_1735,N_1118);
and U2430 (N_2430,N_1797,N_1995);
nor U2431 (N_2431,N_1123,N_1083);
nand U2432 (N_2432,N_1378,N_1679);
and U2433 (N_2433,N_1268,N_1097);
nor U2434 (N_2434,N_1415,N_1714);
or U2435 (N_2435,N_1279,N_1234);
nand U2436 (N_2436,N_1552,N_1318);
or U2437 (N_2437,N_1598,N_1617);
or U2438 (N_2438,N_1299,N_1103);
or U2439 (N_2439,N_1351,N_1176);
nand U2440 (N_2440,N_1657,N_1016);
nor U2441 (N_2441,N_1218,N_1533);
nand U2442 (N_2442,N_1027,N_1186);
nor U2443 (N_2443,N_1741,N_1708);
nand U2444 (N_2444,N_1849,N_1680);
nor U2445 (N_2445,N_1888,N_1822);
or U2446 (N_2446,N_1683,N_1065);
nand U2447 (N_2447,N_1758,N_1386);
and U2448 (N_2448,N_1865,N_1525);
or U2449 (N_2449,N_1313,N_1045);
nand U2450 (N_2450,N_1269,N_1555);
or U2451 (N_2451,N_1095,N_1138);
nand U2452 (N_2452,N_1181,N_1015);
or U2453 (N_2453,N_1836,N_1694);
or U2454 (N_2454,N_1504,N_1048);
or U2455 (N_2455,N_1688,N_1650);
and U2456 (N_2456,N_1757,N_1900);
or U2457 (N_2457,N_1000,N_1067);
or U2458 (N_2458,N_1137,N_1230);
or U2459 (N_2459,N_1119,N_1762);
nor U2460 (N_2460,N_1105,N_1971);
or U2461 (N_2461,N_1124,N_1745);
nor U2462 (N_2462,N_1701,N_1156);
nor U2463 (N_2463,N_1911,N_1142);
nor U2464 (N_2464,N_1882,N_1460);
or U2465 (N_2465,N_1530,N_1503);
or U2466 (N_2466,N_1409,N_1669);
nand U2467 (N_2467,N_1056,N_1539);
nor U2468 (N_2468,N_1170,N_1761);
nor U2469 (N_2469,N_1718,N_1653);
and U2470 (N_2470,N_1467,N_1417);
nor U2471 (N_2471,N_1807,N_1370);
and U2472 (N_2472,N_1316,N_1687);
and U2473 (N_2473,N_1831,N_1754);
or U2474 (N_2474,N_1321,N_1476);
and U2475 (N_2475,N_1623,N_1646);
nor U2476 (N_2476,N_1960,N_1948);
nand U2477 (N_2477,N_1830,N_1098);
or U2478 (N_2478,N_1442,N_1576);
or U2479 (N_2479,N_1112,N_1354);
nand U2480 (N_2480,N_1271,N_1951);
nand U2481 (N_2481,N_1698,N_1344);
and U2482 (N_2482,N_1557,N_1422);
or U2483 (N_2483,N_1571,N_1029);
nand U2484 (N_2484,N_1956,N_1649);
nor U2485 (N_2485,N_1731,N_1004);
and U2486 (N_2486,N_1566,N_1826);
nor U2487 (N_2487,N_1464,N_1326);
nand U2488 (N_2488,N_1834,N_1094);
nand U2489 (N_2489,N_1782,N_1895);
nor U2490 (N_2490,N_1358,N_1314);
nand U2491 (N_2491,N_1339,N_1804);
or U2492 (N_2492,N_1652,N_1217);
nor U2493 (N_2493,N_1821,N_1898);
and U2494 (N_2494,N_1241,N_1303);
nand U2495 (N_2495,N_1486,N_1832);
and U2496 (N_2496,N_1106,N_1568);
and U2497 (N_2497,N_1930,N_1233);
nand U2498 (N_2498,N_1704,N_1607);
and U2499 (N_2499,N_1624,N_1199);
nor U2500 (N_2500,N_1838,N_1814);
and U2501 (N_2501,N_1840,N_1063);
or U2502 (N_2502,N_1757,N_1015);
or U2503 (N_2503,N_1563,N_1477);
nand U2504 (N_2504,N_1462,N_1769);
nor U2505 (N_2505,N_1208,N_1414);
and U2506 (N_2506,N_1836,N_1844);
and U2507 (N_2507,N_1519,N_1807);
nand U2508 (N_2508,N_1569,N_1472);
and U2509 (N_2509,N_1669,N_1618);
nor U2510 (N_2510,N_1349,N_1946);
nor U2511 (N_2511,N_1161,N_1524);
and U2512 (N_2512,N_1596,N_1940);
nor U2513 (N_2513,N_1238,N_1583);
nor U2514 (N_2514,N_1340,N_1582);
or U2515 (N_2515,N_1281,N_1661);
or U2516 (N_2516,N_1020,N_1586);
nand U2517 (N_2517,N_1411,N_1510);
nand U2518 (N_2518,N_1808,N_1697);
xor U2519 (N_2519,N_1057,N_1279);
or U2520 (N_2520,N_1636,N_1273);
nor U2521 (N_2521,N_1282,N_1404);
and U2522 (N_2522,N_1727,N_1136);
or U2523 (N_2523,N_1193,N_1744);
and U2524 (N_2524,N_1457,N_1753);
and U2525 (N_2525,N_1239,N_1543);
nor U2526 (N_2526,N_1116,N_1759);
nand U2527 (N_2527,N_1655,N_1991);
or U2528 (N_2528,N_1336,N_1526);
or U2529 (N_2529,N_1726,N_1075);
nand U2530 (N_2530,N_1990,N_1607);
xnor U2531 (N_2531,N_1856,N_1129);
nor U2532 (N_2532,N_1185,N_1525);
and U2533 (N_2533,N_1878,N_1142);
nand U2534 (N_2534,N_1773,N_1062);
and U2535 (N_2535,N_1753,N_1175);
or U2536 (N_2536,N_1713,N_1759);
nand U2537 (N_2537,N_1100,N_1796);
nand U2538 (N_2538,N_1818,N_1584);
or U2539 (N_2539,N_1724,N_1259);
and U2540 (N_2540,N_1080,N_1170);
and U2541 (N_2541,N_1931,N_1176);
nor U2542 (N_2542,N_1782,N_1468);
and U2543 (N_2543,N_1604,N_1114);
nand U2544 (N_2544,N_1292,N_1159);
nor U2545 (N_2545,N_1853,N_1090);
nand U2546 (N_2546,N_1160,N_1908);
or U2547 (N_2547,N_1582,N_1165);
nor U2548 (N_2548,N_1188,N_1350);
and U2549 (N_2549,N_1074,N_1493);
nor U2550 (N_2550,N_1168,N_1175);
nand U2551 (N_2551,N_1247,N_1558);
nand U2552 (N_2552,N_1189,N_1361);
and U2553 (N_2553,N_1707,N_1884);
or U2554 (N_2554,N_1392,N_1801);
nor U2555 (N_2555,N_1864,N_1666);
nand U2556 (N_2556,N_1131,N_1679);
or U2557 (N_2557,N_1844,N_1017);
nor U2558 (N_2558,N_1012,N_1680);
and U2559 (N_2559,N_1289,N_1460);
nand U2560 (N_2560,N_1743,N_1761);
nand U2561 (N_2561,N_1913,N_1993);
and U2562 (N_2562,N_1302,N_1678);
and U2563 (N_2563,N_1544,N_1346);
nand U2564 (N_2564,N_1721,N_1075);
or U2565 (N_2565,N_1136,N_1354);
or U2566 (N_2566,N_1292,N_1704);
and U2567 (N_2567,N_1317,N_1910);
or U2568 (N_2568,N_1370,N_1761);
nor U2569 (N_2569,N_1982,N_1309);
and U2570 (N_2570,N_1462,N_1536);
or U2571 (N_2571,N_1140,N_1110);
nand U2572 (N_2572,N_1935,N_1439);
nand U2573 (N_2573,N_1542,N_1867);
nand U2574 (N_2574,N_1683,N_1637);
and U2575 (N_2575,N_1686,N_1156);
or U2576 (N_2576,N_1720,N_1380);
and U2577 (N_2577,N_1633,N_1308);
or U2578 (N_2578,N_1730,N_1593);
nand U2579 (N_2579,N_1652,N_1129);
or U2580 (N_2580,N_1638,N_1667);
nor U2581 (N_2581,N_1798,N_1308);
or U2582 (N_2582,N_1359,N_1706);
or U2583 (N_2583,N_1163,N_1929);
or U2584 (N_2584,N_1068,N_1773);
and U2585 (N_2585,N_1029,N_1568);
nand U2586 (N_2586,N_1752,N_1508);
or U2587 (N_2587,N_1777,N_1553);
nand U2588 (N_2588,N_1023,N_1685);
nand U2589 (N_2589,N_1616,N_1043);
nor U2590 (N_2590,N_1472,N_1182);
nor U2591 (N_2591,N_1972,N_1827);
nand U2592 (N_2592,N_1946,N_1635);
and U2593 (N_2593,N_1239,N_1947);
and U2594 (N_2594,N_1766,N_1464);
nand U2595 (N_2595,N_1897,N_1975);
nand U2596 (N_2596,N_1227,N_1602);
and U2597 (N_2597,N_1158,N_1710);
nor U2598 (N_2598,N_1480,N_1436);
or U2599 (N_2599,N_1978,N_1687);
and U2600 (N_2600,N_1054,N_1667);
nand U2601 (N_2601,N_1646,N_1294);
nand U2602 (N_2602,N_1070,N_1306);
and U2603 (N_2603,N_1818,N_1321);
or U2604 (N_2604,N_1520,N_1976);
nor U2605 (N_2605,N_1162,N_1103);
nor U2606 (N_2606,N_1262,N_1633);
nor U2607 (N_2607,N_1567,N_1696);
and U2608 (N_2608,N_1130,N_1053);
nand U2609 (N_2609,N_1636,N_1432);
and U2610 (N_2610,N_1821,N_1642);
nor U2611 (N_2611,N_1386,N_1003);
and U2612 (N_2612,N_1834,N_1903);
or U2613 (N_2613,N_1998,N_1068);
or U2614 (N_2614,N_1377,N_1047);
nand U2615 (N_2615,N_1202,N_1953);
nor U2616 (N_2616,N_1624,N_1247);
or U2617 (N_2617,N_1707,N_1136);
or U2618 (N_2618,N_1074,N_1353);
nand U2619 (N_2619,N_1620,N_1225);
nor U2620 (N_2620,N_1261,N_1580);
nand U2621 (N_2621,N_1042,N_1632);
nand U2622 (N_2622,N_1796,N_1472);
nand U2623 (N_2623,N_1541,N_1487);
nand U2624 (N_2624,N_1227,N_1577);
or U2625 (N_2625,N_1547,N_1182);
and U2626 (N_2626,N_1609,N_1169);
or U2627 (N_2627,N_1980,N_1364);
and U2628 (N_2628,N_1984,N_1632);
and U2629 (N_2629,N_1747,N_1650);
nor U2630 (N_2630,N_1210,N_1012);
nor U2631 (N_2631,N_1109,N_1481);
nand U2632 (N_2632,N_1542,N_1832);
xnor U2633 (N_2633,N_1791,N_1326);
nor U2634 (N_2634,N_1178,N_1111);
nand U2635 (N_2635,N_1008,N_1796);
or U2636 (N_2636,N_1730,N_1020);
nand U2637 (N_2637,N_1259,N_1851);
and U2638 (N_2638,N_1538,N_1030);
and U2639 (N_2639,N_1425,N_1664);
nand U2640 (N_2640,N_1900,N_1065);
xor U2641 (N_2641,N_1745,N_1780);
nand U2642 (N_2642,N_1944,N_1784);
nor U2643 (N_2643,N_1941,N_1883);
and U2644 (N_2644,N_1361,N_1053);
xor U2645 (N_2645,N_1124,N_1485);
and U2646 (N_2646,N_1034,N_1480);
nor U2647 (N_2647,N_1170,N_1222);
nor U2648 (N_2648,N_1335,N_1886);
and U2649 (N_2649,N_1447,N_1010);
or U2650 (N_2650,N_1269,N_1678);
and U2651 (N_2651,N_1212,N_1416);
nand U2652 (N_2652,N_1280,N_1933);
nand U2653 (N_2653,N_1414,N_1502);
nand U2654 (N_2654,N_1340,N_1695);
and U2655 (N_2655,N_1018,N_1811);
and U2656 (N_2656,N_1466,N_1896);
and U2657 (N_2657,N_1480,N_1292);
and U2658 (N_2658,N_1817,N_1654);
or U2659 (N_2659,N_1380,N_1732);
or U2660 (N_2660,N_1611,N_1991);
and U2661 (N_2661,N_1758,N_1472);
nand U2662 (N_2662,N_1164,N_1330);
and U2663 (N_2663,N_1050,N_1615);
nor U2664 (N_2664,N_1388,N_1771);
or U2665 (N_2665,N_1326,N_1180);
or U2666 (N_2666,N_1267,N_1789);
and U2667 (N_2667,N_1735,N_1604);
and U2668 (N_2668,N_1108,N_1190);
nor U2669 (N_2669,N_1888,N_1492);
nand U2670 (N_2670,N_1709,N_1016);
and U2671 (N_2671,N_1136,N_1804);
nor U2672 (N_2672,N_1107,N_1881);
or U2673 (N_2673,N_1924,N_1572);
nor U2674 (N_2674,N_1095,N_1257);
nand U2675 (N_2675,N_1516,N_1523);
nand U2676 (N_2676,N_1158,N_1134);
and U2677 (N_2677,N_1296,N_1093);
nor U2678 (N_2678,N_1273,N_1887);
and U2679 (N_2679,N_1150,N_1546);
or U2680 (N_2680,N_1881,N_1206);
or U2681 (N_2681,N_1829,N_1792);
or U2682 (N_2682,N_1030,N_1772);
or U2683 (N_2683,N_1536,N_1021);
nor U2684 (N_2684,N_1787,N_1826);
or U2685 (N_2685,N_1590,N_1923);
and U2686 (N_2686,N_1816,N_1686);
nand U2687 (N_2687,N_1298,N_1601);
nand U2688 (N_2688,N_1977,N_1465);
or U2689 (N_2689,N_1893,N_1285);
or U2690 (N_2690,N_1781,N_1009);
nor U2691 (N_2691,N_1808,N_1030);
or U2692 (N_2692,N_1841,N_1043);
nor U2693 (N_2693,N_1613,N_1831);
nand U2694 (N_2694,N_1824,N_1819);
and U2695 (N_2695,N_1083,N_1538);
nand U2696 (N_2696,N_1418,N_1766);
nor U2697 (N_2697,N_1010,N_1817);
nand U2698 (N_2698,N_1826,N_1418);
and U2699 (N_2699,N_1870,N_1038);
and U2700 (N_2700,N_1103,N_1000);
or U2701 (N_2701,N_1880,N_1800);
or U2702 (N_2702,N_1385,N_1538);
nand U2703 (N_2703,N_1761,N_1850);
nand U2704 (N_2704,N_1039,N_1654);
nor U2705 (N_2705,N_1316,N_1917);
nand U2706 (N_2706,N_1288,N_1653);
and U2707 (N_2707,N_1471,N_1514);
or U2708 (N_2708,N_1802,N_1246);
nor U2709 (N_2709,N_1214,N_1818);
nand U2710 (N_2710,N_1751,N_1623);
and U2711 (N_2711,N_1722,N_1365);
or U2712 (N_2712,N_1334,N_1693);
or U2713 (N_2713,N_1676,N_1828);
xnor U2714 (N_2714,N_1604,N_1253);
nand U2715 (N_2715,N_1057,N_1065);
nand U2716 (N_2716,N_1202,N_1437);
and U2717 (N_2717,N_1059,N_1900);
or U2718 (N_2718,N_1071,N_1124);
nor U2719 (N_2719,N_1161,N_1957);
or U2720 (N_2720,N_1400,N_1116);
nor U2721 (N_2721,N_1680,N_1129);
nor U2722 (N_2722,N_1972,N_1037);
nor U2723 (N_2723,N_1809,N_1599);
nand U2724 (N_2724,N_1727,N_1776);
nor U2725 (N_2725,N_1469,N_1676);
or U2726 (N_2726,N_1392,N_1247);
nand U2727 (N_2727,N_1143,N_1670);
or U2728 (N_2728,N_1047,N_1097);
and U2729 (N_2729,N_1474,N_1602);
nor U2730 (N_2730,N_1504,N_1928);
nor U2731 (N_2731,N_1868,N_1269);
nand U2732 (N_2732,N_1689,N_1785);
or U2733 (N_2733,N_1489,N_1152);
and U2734 (N_2734,N_1460,N_1952);
or U2735 (N_2735,N_1774,N_1668);
nand U2736 (N_2736,N_1822,N_1251);
nor U2737 (N_2737,N_1948,N_1782);
or U2738 (N_2738,N_1510,N_1206);
or U2739 (N_2739,N_1797,N_1339);
nand U2740 (N_2740,N_1945,N_1442);
nand U2741 (N_2741,N_1103,N_1300);
nand U2742 (N_2742,N_1431,N_1850);
and U2743 (N_2743,N_1021,N_1422);
nor U2744 (N_2744,N_1174,N_1865);
nand U2745 (N_2745,N_1540,N_1473);
and U2746 (N_2746,N_1697,N_1051);
or U2747 (N_2747,N_1399,N_1800);
and U2748 (N_2748,N_1998,N_1278);
nor U2749 (N_2749,N_1860,N_1759);
and U2750 (N_2750,N_1746,N_1310);
nand U2751 (N_2751,N_1760,N_1323);
nand U2752 (N_2752,N_1584,N_1655);
and U2753 (N_2753,N_1568,N_1957);
nand U2754 (N_2754,N_1654,N_1072);
nand U2755 (N_2755,N_1361,N_1082);
nand U2756 (N_2756,N_1375,N_1448);
nand U2757 (N_2757,N_1111,N_1244);
nor U2758 (N_2758,N_1293,N_1243);
and U2759 (N_2759,N_1524,N_1683);
or U2760 (N_2760,N_1626,N_1614);
and U2761 (N_2761,N_1561,N_1601);
and U2762 (N_2762,N_1181,N_1355);
or U2763 (N_2763,N_1333,N_1600);
nor U2764 (N_2764,N_1060,N_1851);
and U2765 (N_2765,N_1805,N_1249);
nor U2766 (N_2766,N_1893,N_1054);
nand U2767 (N_2767,N_1861,N_1858);
or U2768 (N_2768,N_1539,N_1255);
nand U2769 (N_2769,N_1822,N_1350);
or U2770 (N_2770,N_1729,N_1601);
and U2771 (N_2771,N_1984,N_1271);
nand U2772 (N_2772,N_1386,N_1772);
or U2773 (N_2773,N_1130,N_1468);
or U2774 (N_2774,N_1610,N_1345);
and U2775 (N_2775,N_1808,N_1741);
and U2776 (N_2776,N_1077,N_1109);
or U2777 (N_2777,N_1197,N_1113);
or U2778 (N_2778,N_1647,N_1468);
or U2779 (N_2779,N_1598,N_1550);
xor U2780 (N_2780,N_1800,N_1977);
xnor U2781 (N_2781,N_1976,N_1649);
or U2782 (N_2782,N_1649,N_1539);
and U2783 (N_2783,N_1551,N_1049);
nand U2784 (N_2784,N_1596,N_1806);
and U2785 (N_2785,N_1955,N_1157);
and U2786 (N_2786,N_1342,N_1991);
or U2787 (N_2787,N_1126,N_1358);
nand U2788 (N_2788,N_1803,N_1377);
nor U2789 (N_2789,N_1394,N_1900);
xnor U2790 (N_2790,N_1855,N_1556);
or U2791 (N_2791,N_1696,N_1467);
or U2792 (N_2792,N_1529,N_1907);
nor U2793 (N_2793,N_1205,N_1656);
or U2794 (N_2794,N_1571,N_1963);
xor U2795 (N_2795,N_1402,N_1828);
nand U2796 (N_2796,N_1329,N_1546);
nor U2797 (N_2797,N_1270,N_1979);
and U2798 (N_2798,N_1169,N_1223);
nor U2799 (N_2799,N_1378,N_1366);
and U2800 (N_2800,N_1972,N_1254);
or U2801 (N_2801,N_1364,N_1456);
or U2802 (N_2802,N_1664,N_1180);
nor U2803 (N_2803,N_1105,N_1765);
and U2804 (N_2804,N_1535,N_1445);
nand U2805 (N_2805,N_1060,N_1673);
xnor U2806 (N_2806,N_1975,N_1373);
nand U2807 (N_2807,N_1810,N_1510);
nand U2808 (N_2808,N_1528,N_1341);
or U2809 (N_2809,N_1285,N_1282);
nor U2810 (N_2810,N_1174,N_1094);
xnor U2811 (N_2811,N_1085,N_1670);
nor U2812 (N_2812,N_1841,N_1729);
and U2813 (N_2813,N_1041,N_1156);
nand U2814 (N_2814,N_1985,N_1739);
or U2815 (N_2815,N_1092,N_1673);
and U2816 (N_2816,N_1407,N_1398);
or U2817 (N_2817,N_1097,N_1872);
or U2818 (N_2818,N_1381,N_1516);
nand U2819 (N_2819,N_1339,N_1660);
nand U2820 (N_2820,N_1254,N_1452);
nor U2821 (N_2821,N_1170,N_1792);
nand U2822 (N_2822,N_1376,N_1318);
nand U2823 (N_2823,N_1850,N_1931);
nand U2824 (N_2824,N_1918,N_1070);
and U2825 (N_2825,N_1861,N_1087);
nand U2826 (N_2826,N_1248,N_1894);
or U2827 (N_2827,N_1049,N_1745);
nor U2828 (N_2828,N_1713,N_1536);
nor U2829 (N_2829,N_1799,N_1024);
nand U2830 (N_2830,N_1779,N_1021);
nand U2831 (N_2831,N_1935,N_1374);
nor U2832 (N_2832,N_1973,N_1846);
nor U2833 (N_2833,N_1093,N_1411);
and U2834 (N_2834,N_1343,N_1720);
nand U2835 (N_2835,N_1313,N_1132);
nor U2836 (N_2836,N_1079,N_1802);
or U2837 (N_2837,N_1075,N_1408);
nor U2838 (N_2838,N_1158,N_1118);
and U2839 (N_2839,N_1036,N_1945);
xnor U2840 (N_2840,N_1075,N_1942);
nor U2841 (N_2841,N_1752,N_1943);
nand U2842 (N_2842,N_1382,N_1356);
or U2843 (N_2843,N_1722,N_1310);
nand U2844 (N_2844,N_1806,N_1438);
and U2845 (N_2845,N_1921,N_1820);
and U2846 (N_2846,N_1959,N_1652);
or U2847 (N_2847,N_1449,N_1575);
nor U2848 (N_2848,N_1205,N_1602);
and U2849 (N_2849,N_1334,N_1958);
nand U2850 (N_2850,N_1622,N_1562);
or U2851 (N_2851,N_1575,N_1596);
and U2852 (N_2852,N_1976,N_1055);
or U2853 (N_2853,N_1265,N_1471);
nand U2854 (N_2854,N_1647,N_1519);
and U2855 (N_2855,N_1774,N_1650);
nand U2856 (N_2856,N_1962,N_1011);
and U2857 (N_2857,N_1882,N_1915);
or U2858 (N_2858,N_1488,N_1733);
or U2859 (N_2859,N_1864,N_1313);
nand U2860 (N_2860,N_1723,N_1003);
nor U2861 (N_2861,N_1591,N_1471);
and U2862 (N_2862,N_1568,N_1836);
nand U2863 (N_2863,N_1478,N_1175);
nand U2864 (N_2864,N_1993,N_1988);
nand U2865 (N_2865,N_1730,N_1604);
or U2866 (N_2866,N_1548,N_1325);
and U2867 (N_2867,N_1410,N_1284);
nand U2868 (N_2868,N_1519,N_1920);
nand U2869 (N_2869,N_1062,N_1218);
nand U2870 (N_2870,N_1199,N_1039);
nor U2871 (N_2871,N_1137,N_1263);
nor U2872 (N_2872,N_1747,N_1890);
nor U2873 (N_2873,N_1844,N_1425);
or U2874 (N_2874,N_1605,N_1967);
nand U2875 (N_2875,N_1894,N_1633);
nand U2876 (N_2876,N_1726,N_1610);
nand U2877 (N_2877,N_1924,N_1231);
nand U2878 (N_2878,N_1916,N_1954);
and U2879 (N_2879,N_1578,N_1574);
and U2880 (N_2880,N_1952,N_1106);
nor U2881 (N_2881,N_1595,N_1669);
nor U2882 (N_2882,N_1567,N_1124);
xnor U2883 (N_2883,N_1499,N_1489);
nand U2884 (N_2884,N_1626,N_1267);
or U2885 (N_2885,N_1536,N_1587);
nand U2886 (N_2886,N_1516,N_1814);
nor U2887 (N_2887,N_1641,N_1268);
nor U2888 (N_2888,N_1544,N_1200);
nor U2889 (N_2889,N_1734,N_1337);
nor U2890 (N_2890,N_1973,N_1340);
nor U2891 (N_2891,N_1314,N_1136);
nand U2892 (N_2892,N_1350,N_1699);
nand U2893 (N_2893,N_1036,N_1598);
nand U2894 (N_2894,N_1113,N_1480);
nand U2895 (N_2895,N_1717,N_1937);
nand U2896 (N_2896,N_1492,N_1948);
and U2897 (N_2897,N_1670,N_1371);
nand U2898 (N_2898,N_1460,N_1682);
or U2899 (N_2899,N_1034,N_1612);
and U2900 (N_2900,N_1484,N_1697);
and U2901 (N_2901,N_1623,N_1697);
and U2902 (N_2902,N_1008,N_1122);
nor U2903 (N_2903,N_1148,N_1058);
nor U2904 (N_2904,N_1981,N_1774);
nand U2905 (N_2905,N_1781,N_1038);
or U2906 (N_2906,N_1632,N_1255);
or U2907 (N_2907,N_1184,N_1346);
nand U2908 (N_2908,N_1150,N_1378);
nor U2909 (N_2909,N_1062,N_1734);
nor U2910 (N_2910,N_1016,N_1334);
nand U2911 (N_2911,N_1083,N_1036);
and U2912 (N_2912,N_1050,N_1974);
nor U2913 (N_2913,N_1157,N_1483);
or U2914 (N_2914,N_1412,N_1721);
or U2915 (N_2915,N_1996,N_1151);
and U2916 (N_2916,N_1388,N_1351);
nor U2917 (N_2917,N_1296,N_1146);
and U2918 (N_2918,N_1610,N_1211);
or U2919 (N_2919,N_1636,N_1166);
nand U2920 (N_2920,N_1218,N_1473);
nor U2921 (N_2921,N_1039,N_1486);
nor U2922 (N_2922,N_1283,N_1933);
or U2923 (N_2923,N_1957,N_1368);
and U2924 (N_2924,N_1762,N_1903);
nand U2925 (N_2925,N_1206,N_1332);
and U2926 (N_2926,N_1209,N_1966);
or U2927 (N_2927,N_1787,N_1615);
nor U2928 (N_2928,N_1066,N_1390);
nand U2929 (N_2929,N_1175,N_1916);
and U2930 (N_2930,N_1901,N_1843);
xor U2931 (N_2931,N_1510,N_1784);
nor U2932 (N_2932,N_1627,N_1063);
xnor U2933 (N_2933,N_1559,N_1632);
nor U2934 (N_2934,N_1271,N_1447);
or U2935 (N_2935,N_1952,N_1084);
nand U2936 (N_2936,N_1126,N_1038);
nand U2937 (N_2937,N_1292,N_1108);
nor U2938 (N_2938,N_1830,N_1871);
nand U2939 (N_2939,N_1033,N_1215);
and U2940 (N_2940,N_1845,N_1207);
nand U2941 (N_2941,N_1683,N_1301);
nor U2942 (N_2942,N_1644,N_1783);
and U2943 (N_2943,N_1681,N_1371);
and U2944 (N_2944,N_1232,N_1782);
or U2945 (N_2945,N_1938,N_1973);
and U2946 (N_2946,N_1183,N_1562);
nand U2947 (N_2947,N_1241,N_1453);
or U2948 (N_2948,N_1700,N_1733);
nand U2949 (N_2949,N_1920,N_1278);
nand U2950 (N_2950,N_1358,N_1080);
nand U2951 (N_2951,N_1238,N_1716);
and U2952 (N_2952,N_1520,N_1477);
nand U2953 (N_2953,N_1251,N_1249);
and U2954 (N_2954,N_1666,N_1461);
nor U2955 (N_2955,N_1777,N_1506);
or U2956 (N_2956,N_1614,N_1750);
or U2957 (N_2957,N_1465,N_1456);
and U2958 (N_2958,N_1269,N_1017);
nor U2959 (N_2959,N_1440,N_1385);
and U2960 (N_2960,N_1732,N_1534);
nor U2961 (N_2961,N_1619,N_1745);
and U2962 (N_2962,N_1019,N_1654);
and U2963 (N_2963,N_1878,N_1937);
nor U2964 (N_2964,N_1836,N_1927);
and U2965 (N_2965,N_1512,N_1431);
nand U2966 (N_2966,N_1554,N_1711);
nor U2967 (N_2967,N_1347,N_1850);
nor U2968 (N_2968,N_1606,N_1320);
and U2969 (N_2969,N_1369,N_1053);
or U2970 (N_2970,N_1689,N_1258);
and U2971 (N_2971,N_1076,N_1349);
nand U2972 (N_2972,N_1471,N_1941);
nor U2973 (N_2973,N_1396,N_1288);
or U2974 (N_2974,N_1002,N_1102);
and U2975 (N_2975,N_1888,N_1931);
nor U2976 (N_2976,N_1607,N_1915);
nor U2977 (N_2977,N_1829,N_1950);
nor U2978 (N_2978,N_1100,N_1606);
nand U2979 (N_2979,N_1755,N_1921);
nor U2980 (N_2980,N_1710,N_1606);
nor U2981 (N_2981,N_1195,N_1011);
nand U2982 (N_2982,N_1530,N_1618);
nor U2983 (N_2983,N_1821,N_1210);
or U2984 (N_2984,N_1992,N_1932);
and U2985 (N_2985,N_1846,N_1612);
xnor U2986 (N_2986,N_1019,N_1917);
and U2987 (N_2987,N_1522,N_1830);
nor U2988 (N_2988,N_1775,N_1064);
or U2989 (N_2989,N_1309,N_1039);
and U2990 (N_2990,N_1819,N_1211);
or U2991 (N_2991,N_1353,N_1585);
nor U2992 (N_2992,N_1047,N_1479);
nor U2993 (N_2993,N_1144,N_1226);
and U2994 (N_2994,N_1818,N_1015);
or U2995 (N_2995,N_1778,N_1740);
and U2996 (N_2996,N_1309,N_1474);
or U2997 (N_2997,N_1179,N_1178);
nand U2998 (N_2998,N_1362,N_1842);
and U2999 (N_2999,N_1827,N_1356);
xor UO_0 (O_0,N_2290,N_2712);
and UO_1 (O_1,N_2232,N_2765);
nand UO_2 (O_2,N_2278,N_2953);
or UO_3 (O_3,N_2663,N_2872);
or UO_4 (O_4,N_2309,N_2222);
nand UO_5 (O_5,N_2142,N_2073);
and UO_6 (O_6,N_2137,N_2514);
nand UO_7 (O_7,N_2373,N_2093);
or UO_8 (O_8,N_2828,N_2587);
or UO_9 (O_9,N_2105,N_2380);
nor UO_10 (O_10,N_2383,N_2374);
or UO_11 (O_11,N_2002,N_2476);
nand UO_12 (O_12,N_2288,N_2504);
nor UO_13 (O_13,N_2990,N_2647);
nor UO_14 (O_14,N_2541,N_2867);
or UO_15 (O_15,N_2273,N_2513);
and UO_16 (O_16,N_2148,N_2890);
or UO_17 (O_17,N_2671,N_2972);
and UO_18 (O_18,N_2857,N_2451);
nand UO_19 (O_19,N_2930,N_2202);
and UO_20 (O_20,N_2092,N_2564);
nor UO_21 (O_21,N_2882,N_2796);
and UO_22 (O_22,N_2929,N_2711);
and UO_23 (O_23,N_2899,N_2943);
nand UO_24 (O_24,N_2651,N_2086);
nand UO_25 (O_25,N_2279,N_2790);
nor UO_26 (O_26,N_2859,N_2730);
or UO_27 (O_27,N_2988,N_2897);
nand UO_28 (O_28,N_2455,N_2303);
nor UO_29 (O_29,N_2694,N_2153);
nor UO_30 (O_30,N_2447,N_2179);
nand UO_31 (O_31,N_2428,N_2047);
or UO_32 (O_32,N_2237,N_2933);
nor UO_33 (O_33,N_2617,N_2660);
or UO_34 (O_34,N_2408,N_2421);
or UO_35 (O_35,N_2205,N_2847);
nor UO_36 (O_36,N_2611,N_2007);
and UO_37 (O_37,N_2597,N_2117);
or UO_38 (O_38,N_2225,N_2684);
or UO_39 (O_39,N_2794,N_2250);
or UO_40 (O_40,N_2324,N_2434);
or UO_41 (O_41,N_2572,N_2316);
nor UO_42 (O_42,N_2576,N_2082);
or UO_43 (O_43,N_2128,N_2813);
or UO_44 (O_44,N_2615,N_2718);
xnor UO_45 (O_45,N_2887,N_2444);
or UO_46 (O_46,N_2581,N_2157);
nor UO_47 (O_47,N_2553,N_2212);
nand UO_48 (O_48,N_2259,N_2844);
nand UO_49 (O_49,N_2479,N_2526);
nor UO_50 (O_50,N_2995,N_2670);
and UO_51 (O_51,N_2679,N_2401);
nor UO_52 (O_52,N_2777,N_2060);
and UO_53 (O_53,N_2644,N_2919);
nand UO_54 (O_54,N_2762,N_2193);
nor UO_55 (O_55,N_2865,N_2135);
nor UO_56 (O_56,N_2336,N_2826);
or UO_57 (O_57,N_2438,N_2822);
nand UO_58 (O_58,N_2666,N_2530);
nor UO_59 (O_59,N_2633,N_2160);
nand UO_60 (O_60,N_2700,N_2422);
and UO_61 (O_61,N_2902,N_2456);
and UO_62 (O_62,N_2731,N_2646);
nand UO_63 (O_63,N_2390,N_2920);
or UO_64 (O_64,N_2307,N_2889);
nand UO_65 (O_65,N_2207,N_2604);
and UO_66 (O_66,N_2816,N_2687);
nand UO_67 (O_67,N_2511,N_2272);
or UO_68 (O_68,N_2292,N_2323);
nor UO_69 (O_69,N_2090,N_2505);
nand UO_70 (O_70,N_2643,N_2426);
or UO_71 (O_71,N_2131,N_2625);
nand UO_72 (O_72,N_2532,N_2430);
or UO_73 (O_73,N_2419,N_2874);
nor UO_74 (O_74,N_2605,N_2125);
nand UO_75 (O_75,N_2562,N_2343);
or UO_76 (O_76,N_2558,N_2856);
xnor UO_77 (O_77,N_2833,N_2123);
nor UO_78 (O_78,N_2043,N_2664);
nand UO_79 (O_79,N_2785,N_2668);
or UO_80 (O_80,N_2612,N_2321);
and UO_81 (O_81,N_2496,N_2406);
nand UO_82 (O_82,N_2989,N_2334);
nand UO_83 (O_83,N_2294,N_2437);
nor UO_84 (O_84,N_2230,N_2876);
nor UO_85 (O_85,N_2720,N_2064);
nor UO_86 (O_86,N_2853,N_2399);
or UO_87 (O_87,N_2282,N_2517);
xnor UO_88 (O_88,N_2599,N_2168);
and UO_89 (O_89,N_2678,N_2405);
and UO_90 (O_90,N_2855,N_2170);
or UO_91 (O_91,N_2531,N_2048);
or UO_92 (O_92,N_2969,N_2404);
nor UO_93 (O_93,N_2979,N_2896);
nand UO_94 (O_94,N_2242,N_2962);
nand UO_95 (O_95,N_2078,N_2848);
nand UO_96 (O_96,N_2649,N_2821);
nor UO_97 (O_97,N_2487,N_2264);
nand UO_98 (O_98,N_2165,N_2369);
xor UO_99 (O_99,N_2509,N_2389);
or UO_100 (O_100,N_2544,N_2598);
and UO_101 (O_101,N_2573,N_2771);
nand UO_102 (O_102,N_2376,N_2787);
and UO_103 (O_103,N_2276,N_2555);
nor UO_104 (O_104,N_2934,N_2901);
and UO_105 (O_105,N_2269,N_2616);
and UO_106 (O_106,N_2782,N_2675);
nand UO_107 (O_107,N_2708,N_2769);
or UO_108 (O_108,N_2546,N_2803);
nor UO_109 (O_109,N_2861,N_2233);
and UO_110 (O_110,N_2843,N_2850);
and UO_111 (O_111,N_2554,N_2780);
and UO_112 (O_112,N_2885,N_2956);
or UO_113 (O_113,N_2158,N_2341);
and UO_114 (O_114,N_2792,N_2226);
nand UO_115 (O_115,N_2880,N_2465);
nand UO_116 (O_116,N_2959,N_2436);
nand UO_117 (O_117,N_2199,N_2370);
nor UO_118 (O_118,N_2963,N_2018);
and UO_119 (O_119,N_2851,N_2819);
nand UO_120 (O_120,N_2274,N_2674);
nor UO_121 (O_121,N_2662,N_2049);
nor UO_122 (O_122,N_2519,N_2707);
nor UO_123 (O_123,N_2468,N_2755);
nor UO_124 (O_124,N_2566,N_2775);
nor UO_125 (O_125,N_2906,N_2525);
nand UO_126 (O_126,N_2032,N_2764);
nand UO_127 (O_127,N_2940,N_2834);
nand UO_128 (O_128,N_2459,N_2055);
xnor UO_129 (O_129,N_2198,N_2799);
nand UO_130 (O_130,N_2098,N_2866);
nor UO_131 (O_131,N_2427,N_2372);
nor UO_132 (O_132,N_2485,N_2724);
nor UO_133 (O_133,N_2354,N_2021);
nor UO_134 (O_134,N_2578,N_2713);
nor UO_135 (O_135,N_2155,N_2143);
nor UO_136 (O_136,N_2881,N_2584);
and UO_137 (O_137,N_2841,N_2085);
and UO_138 (O_138,N_2768,N_2392);
nand UO_139 (O_139,N_2689,N_2395);
or UO_140 (O_140,N_2905,N_2163);
nand UO_141 (O_141,N_2188,N_2375);
nand UO_142 (O_142,N_2508,N_2669);
nand UO_143 (O_143,N_2462,N_2409);
or UO_144 (O_144,N_2502,N_2283);
and UO_145 (O_145,N_2521,N_2246);
nand UO_146 (O_146,N_2493,N_2773);
or UO_147 (O_147,N_2215,N_2045);
and UO_148 (O_148,N_2417,N_2356);
and UO_149 (O_149,N_2154,N_2591);
or UO_150 (O_150,N_2361,N_2868);
and UO_151 (O_151,N_2650,N_2838);
or UO_152 (O_152,N_2397,N_2619);
or UO_153 (O_153,N_2008,N_2330);
or UO_154 (O_154,N_2196,N_2063);
nand UO_155 (O_155,N_2824,N_2875);
or UO_156 (O_156,N_2091,N_2745);
nor UO_157 (O_157,N_2031,N_2363);
nor UO_158 (O_158,N_2482,N_2029);
or UO_159 (O_159,N_2862,N_2015);
nand UO_160 (O_160,N_2034,N_2475);
or UO_161 (O_161,N_2277,N_2115);
xor UO_162 (O_162,N_2596,N_2441);
nand UO_163 (O_163,N_2012,N_2410);
nor UO_164 (O_164,N_2335,N_2297);
and UO_165 (O_165,N_2805,N_2543);
or UO_166 (O_166,N_2568,N_2507);
nor UO_167 (O_167,N_2384,N_2839);
and UO_168 (O_168,N_2197,N_2106);
and UO_169 (O_169,N_2187,N_2345);
nand UO_170 (O_170,N_2977,N_2467);
xnor UO_171 (O_171,N_2173,N_2968);
or UO_172 (O_172,N_2339,N_2067);
nand UO_173 (O_173,N_2463,N_2355);
xnor UO_174 (O_174,N_2414,N_2539);
and UO_175 (O_175,N_2642,N_2837);
nand UO_176 (O_176,N_2315,N_2931);
and UO_177 (O_177,N_2991,N_2314);
or UO_178 (O_178,N_2985,N_2119);
or UO_179 (O_179,N_2299,N_2020);
nor UO_180 (O_180,N_2911,N_2638);
nor UO_181 (O_181,N_2676,N_2879);
nand UO_182 (O_182,N_2697,N_2585);
and UO_183 (O_183,N_2527,N_2784);
nand UO_184 (O_184,N_2066,N_2677);
nor UO_185 (O_185,N_2024,N_2001);
nor UO_186 (O_186,N_2445,N_2104);
nor UO_187 (O_187,N_2975,N_2758);
nand UO_188 (O_188,N_2331,N_2738);
nand UO_189 (O_189,N_2858,N_2068);
nor UO_190 (O_190,N_2888,N_2680);
nor UO_191 (O_191,N_2377,N_2037);
and UO_192 (O_192,N_2348,N_2310);
or UO_193 (O_193,N_2739,N_2565);
nor UO_194 (O_194,N_2652,N_2023);
or UO_195 (O_195,N_2322,N_2027);
and UO_196 (O_196,N_2191,N_2035);
and UO_197 (O_197,N_2192,N_2965);
xnor UO_198 (O_198,N_2912,N_2312);
nor UO_199 (O_199,N_2924,N_2698);
and UO_200 (O_200,N_2057,N_2172);
nand UO_201 (O_201,N_2996,N_2326);
or UO_202 (O_202,N_2522,N_2705);
nand UO_203 (O_203,N_2219,N_2797);
and UO_204 (O_204,N_2512,N_2545);
and UO_205 (O_205,N_2061,N_2084);
and UO_206 (O_206,N_2898,N_2506);
or UO_207 (O_207,N_2171,N_2823);
nor UO_208 (O_208,N_2709,N_2520);
or UO_209 (O_209,N_2448,N_2893);
and UO_210 (O_210,N_2583,N_2261);
nand UO_211 (O_211,N_2329,N_2754);
nor UO_212 (O_212,N_2247,N_2382);
nor UO_213 (O_213,N_2683,N_2159);
nand UO_214 (O_214,N_2088,N_2100);
nand UO_215 (O_215,N_2648,N_2239);
and UO_216 (O_216,N_2767,N_2113);
or UO_217 (O_217,N_2808,N_2999);
and UO_218 (O_218,N_2812,N_2721);
nand UO_219 (O_219,N_2916,N_2289);
or UO_220 (O_220,N_2726,N_2238);
nor UO_221 (O_221,N_2470,N_2588);
nand UO_222 (O_222,N_2510,N_2804);
nand UO_223 (O_223,N_2243,N_2460);
or UO_224 (O_224,N_2516,N_2590);
nand UO_225 (O_225,N_2575,N_2936);
or UO_226 (O_226,N_2005,N_2832);
xor UO_227 (O_227,N_2440,N_2120);
nor UO_228 (O_228,N_2435,N_2184);
and UO_229 (O_229,N_2469,N_2820);
nand UO_230 (O_230,N_2079,N_2500);
nor UO_231 (O_231,N_2715,N_2846);
and UO_232 (O_232,N_2495,N_2110);
nand UO_233 (O_233,N_2103,N_2559);
nand UO_234 (O_234,N_2998,N_2056);
nor UO_235 (O_235,N_2870,N_2254);
and UO_236 (O_236,N_2151,N_2194);
or UO_237 (O_237,N_2014,N_2234);
or UO_238 (O_238,N_2699,N_2150);
and UO_239 (O_239,N_2976,N_2706);
and UO_240 (O_240,N_2645,N_2814);
nand UO_241 (O_241,N_2608,N_2306);
nand UO_242 (O_242,N_2957,N_2019);
xor UO_243 (O_243,N_2641,N_2909);
nor UO_244 (O_244,N_2954,N_2682);
and UO_245 (O_245,N_2478,N_2691);
or UO_246 (O_246,N_2556,N_2665);
or UO_247 (O_247,N_2213,N_2908);
nand UO_248 (O_248,N_2203,N_2696);
and UO_249 (O_249,N_2571,N_2431);
or UO_250 (O_250,N_2621,N_2102);
nor UO_251 (O_251,N_2141,N_2256);
or UO_252 (O_252,N_2340,N_2835);
nand UO_253 (O_253,N_2964,N_2221);
and UO_254 (O_254,N_2371,N_2260);
nor UO_255 (O_255,N_2877,N_2728);
and UO_256 (O_256,N_2791,N_2702);
nand UO_257 (O_257,N_2413,N_2756);
nor UO_258 (O_258,N_2829,N_2842);
nand UO_259 (O_259,N_2942,N_2174);
or UO_260 (O_260,N_2074,N_2951);
or UO_261 (O_261,N_2800,N_2603);
xor UO_262 (O_262,N_2333,N_2627);
or UO_263 (O_263,N_2201,N_2164);
or UO_264 (O_264,N_2200,N_2244);
nand UO_265 (O_265,N_2903,N_2127);
nand UO_266 (O_266,N_2458,N_2904);
nand UO_267 (O_267,N_2752,N_2815);
or UO_268 (O_268,N_2654,N_2537);
and UO_269 (O_269,N_2280,N_2941);
or UO_270 (O_270,N_2549,N_2653);
xnor UO_271 (O_271,N_2097,N_2983);
or UO_272 (O_272,N_2618,N_2026);
nand UO_273 (O_273,N_2845,N_2783);
nand UO_274 (O_274,N_2320,N_2253);
nand UO_275 (O_275,N_2950,N_2347);
and UO_276 (O_276,N_2122,N_2825);
nand UO_277 (O_277,N_2921,N_2656);
nand UO_278 (O_278,N_2925,N_2725);
nand UO_279 (O_279,N_2304,N_2096);
nand UO_280 (O_280,N_2932,N_2116);
or UO_281 (O_281,N_2353,N_2039);
and UO_282 (O_282,N_2966,N_2582);
or UO_283 (O_283,N_2761,N_2381);
nand UO_284 (O_284,N_2614,N_2723);
nand UO_285 (O_285,N_2044,N_2542);
nand UO_286 (O_286,N_2766,N_2255);
or UO_287 (O_287,N_2220,N_2129);
and UO_288 (O_288,N_2042,N_2301);
or UO_289 (O_289,N_2251,N_2795);
nor UO_290 (O_290,N_2631,N_2971);
or UO_291 (O_291,N_2442,N_2852);
or UO_292 (O_292,N_2393,N_2138);
or UO_293 (O_293,N_2017,N_2010);
and UO_294 (O_294,N_2350,N_2368);
nand UO_295 (O_295,N_2305,N_2809);
or UO_296 (O_296,N_2658,N_2801);
nor UO_297 (O_297,N_2515,N_2149);
nor UO_298 (O_298,N_2268,N_2432);
nand UO_299 (O_299,N_2152,N_2275);
or UO_300 (O_300,N_2265,N_2107);
nor UO_301 (O_301,N_2501,N_2217);
or UO_302 (O_302,N_2869,N_2394);
nor UO_303 (O_303,N_2536,N_2692);
nor UO_304 (O_304,N_2236,N_2358);
and UO_305 (O_305,N_2494,N_2425);
nand UO_306 (O_306,N_2147,N_2411);
nand UO_307 (O_307,N_2673,N_2686);
nor UO_308 (O_308,N_2036,N_2992);
or UO_309 (O_309,N_2743,N_2332);
or UO_310 (O_310,N_2849,N_2751);
nand UO_311 (O_311,N_2811,N_2227);
nor UO_312 (O_312,N_2252,N_2607);
or UO_313 (O_313,N_2928,N_2051);
and UO_314 (O_314,N_2630,N_2302);
or UO_315 (O_315,N_2560,N_2806);
or UO_316 (O_316,N_2291,N_2922);
or UO_317 (O_317,N_2121,N_2181);
or UO_318 (O_318,N_2228,N_2831);
nor UO_319 (O_319,N_2997,N_2473);
nand UO_320 (O_320,N_2072,N_2840);
or UO_321 (O_321,N_2567,N_2781);
nand UO_322 (O_322,N_2087,N_2111);
or UO_323 (O_323,N_2481,N_2094);
nor UO_324 (O_324,N_2634,N_2130);
or UO_325 (O_325,N_2917,N_2224);
nand UO_326 (O_326,N_2955,N_2540);
or UO_327 (O_327,N_2945,N_2420);
or UO_328 (O_328,N_2727,N_2214);
or UO_329 (O_329,N_2863,N_2817);
and UO_330 (O_330,N_2241,N_2041);
nand UO_331 (O_331,N_2385,N_2362);
nand UO_332 (O_332,N_2503,N_2970);
nand UO_333 (O_333,N_2145,N_2750);
and UO_334 (O_334,N_2574,N_2364);
or UO_335 (O_335,N_2325,N_2748);
nand UO_336 (O_336,N_2589,N_2740);
nor UO_337 (O_337,N_2285,N_2454);
nor UO_338 (O_338,N_2266,N_2763);
and UO_339 (O_339,N_2894,N_2357);
and UO_340 (O_340,N_2065,N_2439);
xnor UO_341 (O_341,N_2011,N_2552);
and UO_342 (O_342,N_2742,N_2760);
and UO_343 (O_343,N_2810,N_2004);
and UO_344 (O_344,N_2918,N_2871);
xnor UO_345 (O_345,N_2786,N_2714);
nor UO_346 (O_346,N_2058,N_2788);
or UO_347 (O_347,N_2789,N_2703);
and UO_348 (O_348,N_2551,N_2003);
and UO_349 (O_349,N_2025,N_2182);
nor UO_350 (O_350,N_2183,N_2248);
or UO_351 (O_351,N_2218,N_2360);
or UO_352 (O_352,N_2774,N_2579);
or UO_353 (O_353,N_2593,N_2210);
nor UO_354 (O_354,N_2124,N_2146);
and UO_355 (O_355,N_2497,N_2308);
and UO_356 (O_356,N_2594,N_2296);
nand UO_357 (O_357,N_2480,N_2472);
or UO_358 (O_358,N_2717,N_2009);
and UO_359 (O_359,N_2349,N_2327);
and UO_360 (O_360,N_2258,N_2557);
and UO_361 (O_361,N_2229,N_2013);
or UO_362 (O_362,N_2533,N_2561);
or UO_363 (O_363,N_2352,N_2022);
and UO_364 (O_364,N_2211,N_2344);
or UO_365 (O_365,N_2006,N_2592);
nor UO_366 (O_366,N_2623,N_2586);
nand UO_367 (O_367,N_2613,N_2600);
nand UO_368 (O_368,N_2466,N_2878);
or UO_369 (O_369,N_2313,N_2655);
or UO_370 (O_370,N_2547,N_2033);
nor UO_371 (O_371,N_2529,N_2524);
and UO_372 (O_372,N_2538,N_2457);
nand UO_373 (O_373,N_2719,N_2099);
nand UO_374 (O_374,N_2563,N_2778);
nand UO_375 (O_375,N_2949,N_2109);
nor UO_376 (O_376,N_2860,N_2209);
nand UO_377 (O_377,N_2947,N_2262);
or UO_378 (O_378,N_2293,N_2534);
nor UO_379 (O_379,N_2081,N_2367);
or UO_380 (O_380,N_2701,N_2548);
and UO_381 (O_381,N_2915,N_2418);
nand UO_382 (O_382,N_2746,N_2722);
nor UO_383 (O_383,N_2059,N_2484);
nor UO_384 (O_384,N_2854,N_2595);
and UO_385 (O_385,N_2704,N_2873);
nand UO_386 (O_386,N_2747,N_2779);
or UO_387 (O_387,N_2836,N_2914);
and UO_388 (O_388,N_2175,N_2492);
or UO_389 (O_389,N_2772,N_2446);
or UO_390 (O_390,N_2359,N_2491);
nor UO_391 (O_391,N_2973,N_2980);
nand UO_392 (O_392,N_2391,N_2298);
nand UO_393 (O_393,N_2450,N_2681);
nand UO_394 (O_394,N_2400,N_2640);
nor UO_395 (O_395,N_2926,N_2449);
or UO_396 (O_396,N_2365,N_2295);
nand UO_397 (O_397,N_2672,N_2967);
or UO_398 (O_398,N_2161,N_2189);
or UO_399 (O_399,N_2733,N_2076);
or UO_400 (O_400,N_2351,N_2095);
nand UO_401 (O_401,N_2622,N_2378);
and UO_402 (O_402,N_2328,N_2249);
nor UO_403 (O_403,N_2978,N_2030);
and UO_404 (O_404,N_2342,N_2910);
and UO_405 (O_405,N_2190,N_2913);
and UO_406 (O_406,N_2223,N_2038);
nor UO_407 (O_407,N_2069,N_2053);
or UO_408 (O_408,N_2601,N_2606);
or UO_409 (O_409,N_2240,N_2398);
nand UO_410 (O_410,N_2287,N_2518);
nand UO_411 (O_411,N_2499,N_2317);
nand UO_412 (O_412,N_2667,N_2080);
nor UO_413 (O_413,N_2628,N_2284);
nand UO_414 (O_414,N_2028,N_2052);
or UO_415 (O_415,N_2178,N_2452);
nand UO_416 (O_416,N_2054,N_2162);
and UO_417 (O_417,N_2802,N_2402);
and UO_418 (O_418,N_2108,N_2000);
or UO_419 (O_419,N_2016,N_2883);
nor UO_420 (O_420,N_2101,N_2486);
nor UO_421 (O_421,N_2040,N_2661);
or UO_422 (O_422,N_2134,N_2464);
nor UO_423 (O_423,N_2632,N_2577);
and UO_424 (O_424,N_2891,N_2195);
and UO_425 (O_425,N_2884,N_2216);
or UO_426 (O_426,N_2994,N_2270);
and UO_427 (O_427,N_2952,N_2729);
nor UO_428 (O_428,N_2948,N_2089);
and UO_429 (O_429,N_2639,N_2281);
nor UO_430 (O_430,N_2071,N_2620);
and UO_431 (O_431,N_2118,N_2114);
or UO_432 (O_432,N_2489,N_2984);
and UO_433 (O_433,N_2483,N_2477);
nor UO_434 (O_434,N_2245,N_2412);
nand UO_435 (O_435,N_2626,N_2338);
nand UO_436 (O_436,N_2180,N_2659);
nor UO_437 (O_437,N_2423,N_2830);
or UO_438 (O_438,N_2528,N_2416);
nand UO_439 (O_439,N_2946,N_2471);
nor UO_440 (O_440,N_2166,N_2271);
nor UO_441 (O_441,N_2864,N_2987);
or UO_442 (O_442,N_2083,N_2488);
and UO_443 (O_443,N_2132,N_2749);
or UO_444 (O_444,N_2300,N_2523);
and UO_445 (O_445,N_2818,N_2070);
nand UO_446 (O_446,N_2535,N_2629);
or UO_447 (O_447,N_2144,N_2734);
nand UO_448 (O_448,N_2737,N_2167);
or UO_449 (O_449,N_2741,N_2938);
nand UO_450 (O_450,N_2610,N_2403);
nor UO_451 (O_451,N_2757,N_2807);
nor UO_452 (O_452,N_2474,N_2396);
nand UO_453 (O_453,N_2433,N_2235);
and UO_454 (O_454,N_2636,N_2944);
and UO_455 (O_455,N_2206,N_2133);
nand UO_456 (O_456,N_2744,N_2231);
nor UO_457 (O_457,N_2710,N_2993);
and UO_458 (O_458,N_2337,N_2657);
nand UO_459 (O_459,N_2267,N_2886);
or UO_460 (O_460,N_2693,N_2177);
nor UO_461 (O_461,N_2318,N_2974);
and UO_462 (O_462,N_2960,N_2311);
or UO_463 (O_463,N_2075,N_2387);
nor UO_464 (O_464,N_2379,N_2982);
nand UO_465 (O_465,N_2388,N_2895);
nor UO_466 (O_466,N_2569,N_2461);
nor UO_467 (O_467,N_2570,N_2046);
nor UO_468 (O_468,N_2685,N_2732);
nand UO_469 (O_469,N_2156,N_2429);
and UO_470 (O_470,N_2346,N_2490);
and UO_471 (O_471,N_2981,N_2986);
or UO_472 (O_472,N_2776,N_2498);
nand UO_473 (O_473,N_2937,N_2136);
xor UO_474 (O_474,N_2690,N_2935);
and UO_475 (O_475,N_2892,N_2927);
nand UO_476 (O_476,N_2176,N_2958);
nor UO_477 (O_477,N_2759,N_2923);
nand UO_478 (O_478,N_2637,N_2112);
nor UO_479 (O_479,N_2140,N_2263);
xor UO_480 (O_480,N_2580,N_2735);
nand UO_481 (O_481,N_2257,N_2386);
or UO_482 (O_482,N_2550,N_2695);
and UO_483 (O_483,N_2827,N_2286);
or UO_484 (O_484,N_2407,N_2716);
nand UO_485 (O_485,N_2126,N_2753);
nand UO_486 (O_486,N_2186,N_2453);
or UO_487 (O_487,N_2415,N_2319);
and UO_488 (O_488,N_2961,N_2169);
or UO_489 (O_489,N_2900,N_2688);
and UO_490 (O_490,N_2062,N_2443);
and UO_491 (O_491,N_2635,N_2624);
nor UO_492 (O_492,N_2424,N_2609);
nand UO_493 (O_493,N_2793,N_2208);
or UO_494 (O_494,N_2907,N_2185);
nor UO_495 (O_495,N_2939,N_2770);
nand UO_496 (O_496,N_2798,N_2736);
xor UO_497 (O_497,N_2050,N_2077);
nor UO_498 (O_498,N_2366,N_2204);
nor UO_499 (O_499,N_2139,N_2602);
endmodule