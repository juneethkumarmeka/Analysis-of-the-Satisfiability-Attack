module basic_500_3000_500_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_51,In_19);
and U1 (N_1,In_268,In_74);
or U2 (N_2,In_222,In_285);
and U3 (N_3,In_465,In_329);
nand U4 (N_4,In_290,In_429);
nand U5 (N_5,In_207,In_368);
or U6 (N_6,In_45,In_160);
and U7 (N_7,In_122,In_351);
nand U8 (N_8,In_406,In_40);
nor U9 (N_9,In_489,In_103);
or U10 (N_10,In_95,In_302);
nor U11 (N_11,In_66,In_476);
nand U12 (N_12,In_186,In_265);
or U13 (N_13,In_445,In_125);
and U14 (N_14,In_57,In_286);
xnor U15 (N_15,In_34,In_120);
or U16 (N_16,In_91,In_403);
nor U17 (N_17,In_4,In_480);
xnor U18 (N_18,In_372,In_36);
nand U19 (N_19,In_23,In_341);
and U20 (N_20,In_297,In_439);
nor U21 (N_21,In_484,In_176);
nand U22 (N_22,In_294,In_188);
xor U23 (N_23,In_24,In_401);
nor U24 (N_24,In_144,In_300);
or U25 (N_25,In_140,In_166);
and U26 (N_26,In_387,In_382);
or U27 (N_27,In_255,In_203);
nor U28 (N_28,In_195,In_497);
nor U29 (N_29,In_216,In_423);
or U30 (N_30,In_427,In_309);
nor U31 (N_31,In_426,In_250);
or U32 (N_32,In_114,In_93);
or U33 (N_33,In_128,In_230);
xnor U34 (N_34,In_337,In_116);
or U35 (N_35,In_320,In_12);
or U36 (N_36,In_156,In_228);
nand U37 (N_37,In_18,In_436);
or U38 (N_38,In_173,In_377);
and U39 (N_39,In_80,In_213);
nor U40 (N_40,In_152,In_204);
nand U41 (N_41,In_183,In_123);
nor U42 (N_42,In_81,In_360);
and U43 (N_43,In_181,In_459);
nand U44 (N_44,In_494,In_308);
nand U45 (N_45,In_118,In_424);
nand U46 (N_46,In_299,In_146);
or U47 (N_47,In_150,In_194);
or U48 (N_48,In_244,In_327);
xnor U49 (N_49,In_240,In_102);
nor U50 (N_50,In_344,In_31);
nor U51 (N_51,In_440,In_433);
nand U52 (N_52,In_192,In_253);
xnor U53 (N_53,In_217,In_132);
nor U54 (N_54,In_395,In_165);
nor U55 (N_55,In_187,In_223);
and U56 (N_56,In_190,In_291);
nand U57 (N_57,In_227,In_311);
nand U58 (N_58,In_493,In_295);
nand U59 (N_59,In_259,In_96);
nand U60 (N_60,In_212,In_328);
nor U61 (N_61,N_37,In_296);
xnor U62 (N_62,In_14,In_306);
or U63 (N_63,In_282,In_417);
xnor U64 (N_64,In_88,In_85);
nand U65 (N_65,In_314,In_214);
xor U66 (N_66,N_24,In_68);
nand U67 (N_67,N_26,N_19);
nor U68 (N_68,In_389,In_324);
or U69 (N_69,In_474,In_77);
or U70 (N_70,In_243,In_388);
and U71 (N_71,In_371,In_0);
and U72 (N_72,N_38,In_28);
and U73 (N_73,In_272,In_50);
nand U74 (N_74,In_248,In_422);
nor U75 (N_75,In_364,N_5);
xnor U76 (N_76,In_464,In_148);
nor U77 (N_77,In_356,N_16);
or U78 (N_78,In_399,In_30);
and U79 (N_79,In_393,In_63);
xor U80 (N_80,In_266,In_451);
nor U81 (N_81,In_269,In_167);
and U82 (N_82,In_298,In_373);
xnor U83 (N_83,In_257,In_319);
nand U84 (N_84,In_53,In_70);
and U85 (N_85,In_75,In_376);
nor U86 (N_86,In_58,In_164);
nor U87 (N_87,In_444,In_49);
nor U88 (N_88,In_234,In_8);
nor U89 (N_89,In_407,In_496);
or U90 (N_90,In_15,N_51);
or U91 (N_91,In_239,In_2);
or U92 (N_92,In_447,In_115);
nor U93 (N_93,In_492,In_21);
nand U94 (N_94,N_50,N_9);
or U95 (N_95,In_270,In_38);
xor U96 (N_96,In_25,In_416);
and U97 (N_97,In_131,In_461);
nor U98 (N_98,In_54,In_281);
xor U99 (N_99,In_274,N_41);
and U100 (N_100,In_247,In_155);
xor U101 (N_101,In_71,In_108);
xor U102 (N_102,In_437,In_149);
nand U103 (N_103,In_193,In_452);
and U104 (N_104,In_315,In_52);
xor U105 (N_105,In_6,In_462);
and U106 (N_106,In_226,In_60);
or U107 (N_107,In_7,In_105);
xnor U108 (N_108,In_487,In_26);
xor U109 (N_109,In_151,In_402);
and U110 (N_110,In_316,In_370);
xor U111 (N_111,In_415,In_301);
and U112 (N_112,In_335,N_49);
nand U113 (N_113,In_343,In_495);
and U114 (N_114,In_430,In_184);
or U115 (N_115,N_53,N_23);
xnor U116 (N_116,In_43,In_169);
xnor U117 (N_117,In_236,In_200);
and U118 (N_118,In_17,In_267);
nand U119 (N_119,In_143,In_69);
nand U120 (N_120,N_39,In_211);
nand U121 (N_121,In_264,In_5);
nor U122 (N_122,N_75,In_442);
nand U123 (N_123,In_421,In_78);
xor U124 (N_124,In_432,N_60);
and U125 (N_125,In_3,N_10);
nand U126 (N_126,In_163,In_326);
or U127 (N_127,In_279,In_202);
and U128 (N_128,N_55,In_420);
or U129 (N_129,N_3,N_14);
or U130 (N_130,In_305,In_413);
xnor U131 (N_131,N_44,N_45);
xnor U132 (N_132,In_22,In_408);
nor U133 (N_133,In_137,N_84);
nand U134 (N_134,In_446,N_92);
nand U135 (N_135,N_119,N_104);
nand U136 (N_136,In_411,N_82);
nor U137 (N_137,In_225,In_42);
nand U138 (N_138,In_454,In_92);
and U139 (N_139,In_271,N_27);
nand U140 (N_140,In_210,In_472);
or U141 (N_141,In_443,In_482);
nor U142 (N_142,In_157,In_251);
or U143 (N_143,In_27,N_34);
nand U144 (N_144,In_374,In_313);
and U145 (N_145,In_303,N_18);
nor U146 (N_146,In_470,In_384);
xor U147 (N_147,In_55,In_273);
nand U148 (N_148,In_209,In_1);
xor U149 (N_149,N_68,N_71);
nor U150 (N_150,In_357,In_410);
and U151 (N_151,In_127,In_380);
and U152 (N_152,In_242,In_307);
nand U153 (N_153,In_20,In_142);
xor U154 (N_154,N_13,In_352);
xnor U155 (N_155,In_353,N_98);
nand U156 (N_156,In_256,N_57);
and U157 (N_157,N_20,In_121);
nand U158 (N_158,In_392,In_232);
xor U159 (N_159,In_350,N_63);
nand U160 (N_160,In_62,In_134);
or U161 (N_161,In_189,In_486);
xor U162 (N_162,In_87,In_381);
and U163 (N_163,N_0,In_278);
or U164 (N_164,In_277,In_107);
xor U165 (N_165,In_378,In_359);
and U166 (N_166,In_16,N_8);
or U167 (N_167,In_218,N_12);
and U168 (N_168,In_129,In_383);
xnor U169 (N_169,In_477,In_400);
nor U170 (N_170,In_177,N_29);
xnor U171 (N_171,N_102,In_483);
or U172 (N_172,In_44,N_36);
nand U173 (N_173,In_467,N_80);
and U174 (N_174,In_418,In_260);
nor U175 (N_175,N_30,In_398);
or U176 (N_176,N_94,In_138);
xor U177 (N_177,In_224,In_221);
or U178 (N_178,N_110,In_412);
or U179 (N_179,N_35,In_67);
or U180 (N_180,In_37,In_318);
nand U181 (N_181,N_124,In_170);
and U182 (N_182,In_29,In_73);
nand U183 (N_183,In_174,In_197);
nand U184 (N_184,N_58,N_120);
xor U185 (N_185,In_48,In_246);
or U186 (N_186,In_339,N_100);
nor U187 (N_187,N_131,In_365);
or U188 (N_188,N_166,In_419);
or U189 (N_189,In_133,In_453);
and U190 (N_190,In_154,In_47);
nand U191 (N_191,In_229,N_116);
xor U192 (N_192,In_101,In_394);
or U193 (N_193,N_107,N_59);
xor U194 (N_194,N_88,N_150);
and U195 (N_195,In_434,In_141);
nor U196 (N_196,In_145,In_56);
and U197 (N_197,N_95,In_178);
or U198 (N_198,In_64,N_117);
nand U199 (N_199,N_140,In_438);
or U200 (N_200,In_61,In_206);
nor U201 (N_201,N_105,N_22);
nor U202 (N_202,N_97,In_179);
or U203 (N_203,N_96,In_205);
nand U204 (N_204,In_431,In_245);
nor U205 (N_205,In_83,N_72);
xnor U206 (N_206,In_46,N_111);
or U207 (N_207,N_173,N_142);
nand U208 (N_208,N_31,In_32);
or U209 (N_209,In_111,In_396);
or U210 (N_210,In_345,In_468);
or U211 (N_211,In_13,In_304);
nor U212 (N_212,N_101,In_89);
and U213 (N_213,In_79,N_114);
and U214 (N_214,N_91,In_435);
nand U215 (N_215,In_312,N_158);
nor U216 (N_216,In_491,In_198);
xnor U217 (N_217,N_52,In_82);
or U218 (N_218,N_127,In_106);
and U219 (N_219,N_115,In_478);
xnor U220 (N_220,In_386,In_110);
nor U221 (N_221,N_56,N_43);
or U222 (N_222,In_263,In_385);
and U223 (N_223,N_78,N_46);
xnor U224 (N_224,In_488,In_414);
and U225 (N_225,N_28,In_130);
or U226 (N_226,In_258,N_159);
nor U227 (N_227,In_369,N_149);
nand U228 (N_228,In_185,N_179);
and U229 (N_229,In_97,N_62);
or U230 (N_230,In_499,In_10);
xnor U231 (N_231,In_84,In_441);
xnor U232 (N_232,N_69,In_332);
or U233 (N_233,N_89,N_139);
nand U234 (N_234,N_129,In_168);
nor U235 (N_235,In_99,In_35);
nor U236 (N_236,In_126,In_201);
xnor U237 (N_237,In_458,In_117);
or U238 (N_238,N_138,N_66);
nor U239 (N_239,N_160,In_448);
nand U240 (N_240,In_471,N_238);
and U241 (N_241,N_134,In_367);
or U242 (N_242,In_220,N_143);
xnor U243 (N_243,N_141,N_106);
nor U244 (N_244,In_235,In_76);
nor U245 (N_245,N_234,In_119);
xor U246 (N_246,N_212,N_200);
or U247 (N_247,N_199,N_76);
nor U248 (N_248,N_153,In_280);
nor U249 (N_249,In_330,N_2);
nand U250 (N_250,N_182,N_224);
nand U251 (N_251,In_171,N_73);
nand U252 (N_252,In_98,In_254);
xnor U253 (N_253,N_170,N_174);
nand U254 (N_254,In_379,N_81);
nor U255 (N_255,N_90,N_183);
nor U256 (N_256,In_347,In_11);
nor U257 (N_257,N_54,N_135);
nor U258 (N_258,N_147,N_65);
or U259 (N_259,N_228,In_409);
and U260 (N_260,In_293,In_153);
and U261 (N_261,In_284,In_65);
or U262 (N_262,In_196,N_77);
and U263 (N_263,In_182,N_202);
nor U264 (N_264,N_225,In_233);
nand U265 (N_265,In_340,In_262);
and U266 (N_266,N_4,In_390);
xor U267 (N_267,In_490,In_9);
xor U268 (N_268,N_167,In_348);
and U269 (N_269,In_94,N_145);
nand U270 (N_270,In_90,N_189);
nand U271 (N_271,In_355,N_83);
nor U272 (N_272,In_100,In_208);
xnor U273 (N_273,In_289,N_239);
or U274 (N_274,In_238,N_186);
and U275 (N_275,N_227,In_231);
xor U276 (N_276,N_184,In_336);
xor U277 (N_277,N_137,N_118);
or U278 (N_278,N_128,N_237);
xor U279 (N_279,In_172,N_47);
nor U280 (N_280,N_132,In_322);
xor U281 (N_281,N_74,N_122);
nor U282 (N_282,In_366,N_205);
xor U283 (N_283,N_148,N_230);
xor U284 (N_284,N_171,N_220);
or U285 (N_285,N_165,N_164);
xor U286 (N_286,In_288,N_21);
xnor U287 (N_287,In_404,N_172);
or U288 (N_288,N_103,In_466);
nor U289 (N_289,N_70,N_144);
nor U290 (N_290,N_168,In_159);
and U291 (N_291,In_449,N_197);
or U292 (N_292,N_32,In_460);
nand U293 (N_293,N_236,N_176);
xor U294 (N_294,In_310,In_104);
nand U295 (N_295,N_42,In_39);
nor U296 (N_296,N_204,In_346);
xor U297 (N_297,In_252,N_191);
and U298 (N_298,N_194,N_218);
nand U299 (N_299,In_283,N_109);
nand U300 (N_300,N_217,N_206);
or U301 (N_301,In_109,N_175);
xor U302 (N_302,N_258,In_475);
xnor U303 (N_303,In_479,N_267);
or U304 (N_304,N_245,N_249);
nor U305 (N_305,N_264,N_93);
and U306 (N_306,N_209,In_215);
or U307 (N_307,N_178,N_155);
or U308 (N_308,N_290,N_192);
xor U309 (N_309,N_283,In_199);
nor U310 (N_310,N_231,N_246);
nand U311 (N_311,In_219,N_275);
nand U312 (N_312,N_196,N_40);
or U313 (N_313,In_162,N_6);
nor U314 (N_314,N_87,N_297);
and U315 (N_315,N_195,N_61);
nor U316 (N_316,N_281,N_203);
nand U317 (N_317,N_270,In_498);
xnor U318 (N_318,In_33,N_48);
and U319 (N_319,N_208,N_284);
xor U320 (N_320,N_298,In_455);
or U321 (N_321,N_279,In_361);
nand U322 (N_322,In_463,In_191);
or U323 (N_323,N_251,N_193);
nor U324 (N_324,N_274,N_222);
or U325 (N_325,N_180,N_219);
nand U326 (N_326,In_287,N_240);
nor U327 (N_327,N_252,N_287);
and U328 (N_328,N_126,In_241);
or U329 (N_329,In_139,In_331);
or U330 (N_330,N_226,N_157);
xnor U331 (N_331,N_241,In_428);
nor U332 (N_332,N_272,N_112);
nand U333 (N_333,N_294,N_280);
nor U334 (N_334,N_262,N_278);
and U335 (N_335,N_64,N_125);
nand U336 (N_336,N_291,N_266);
nor U337 (N_337,N_133,In_261);
nor U338 (N_338,N_121,In_86);
or U339 (N_339,N_11,In_59);
and U340 (N_340,N_99,N_295);
or U341 (N_341,N_221,N_25);
nor U342 (N_342,N_235,N_113);
xnor U343 (N_343,In_342,N_242);
nor U344 (N_344,N_1,In_275);
or U345 (N_345,In_450,In_334);
and U346 (N_346,N_156,N_130);
or U347 (N_347,N_247,In_349);
nor U348 (N_348,N_292,N_271);
xor U349 (N_349,N_233,N_15);
nand U350 (N_350,N_282,N_162);
and U351 (N_351,N_215,In_469);
xor U352 (N_352,N_86,N_289);
or U353 (N_353,N_268,N_273);
and U354 (N_354,In_41,N_259);
and U355 (N_355,N_296,In_457);
xor U356 (N_356,In_136,In_481);
nor U357 (N_357,In_323,N_181);
xnor U358 (N_358,N_108,N_67);
or U359 (N_359,In_338,N_210);
nand U360 (N_360,N_342,In_358);
or U361 (N_361,N_315,N_254);
nand U362 (N_362,N_351,N_255);
or U363 (N_363,N_344,N_243);
and U364 (N_364,N_185,N_256);
or U365 (N_365,N_146,In_147);
nand U366 (N_366,In_249,In_473);
xnor U367 (N_367,N_177,In_161);
xor U368 (N_368,N_321,In_112);
xor U369 (N_369,N_323,N_356);
xor U370 (N_370,N_314,N_304);
nor U371 (N_371,N_311,N_347);
and U372 (N_372,N_232,N_305);
and U373 (N_373,N_327,N_265);
or U374 (N_374,N_188,N_244);
xor U375 (N_375,In_333,In_391);
nor U376 (N_376,N_357,N_322);
and U377 (N_377,In_124,N_317);
nand U378 (N_378,N_123,N_349);
nor U379 (N_379,In_237,N_335);
xnor U380 (N_380,In_375,N_85);
or U381 (N_381,N_248,N_312);
and U382 (N_382,N_211,N_313);
and U383 (N_383,N_341,N_263);
nor U384 (N_384,N_33,In_485);
or U385 (N_385,N_352,N_355);
xnor U386 (N_386,In_135,N_300);
nand U387 (N_387,In_321,N_187);
or U388 (N_388,N_340,N_151);
xor U389 (N_389,N_331,N_310);
and U390 (N_390,N_7,N_336);
or U391 (N_391,N_261,In_362);
or U392 (N_392,N_354,N_223);
nor U393 (N_393,In_354,In_317);
xnor U394 (N_394,N_328,N_318);
nor U395 (N_395,N_253,N_330);
and U396 (N_396,In_175,In_158);
nand U397 (N_397,N_277,N_276);
and U398 (N_398,N_79,N_332);
xnor U399 (N_399,N_316,N_319);
nor U400 (N_400,In_456,N_325);
nor U401 (N_401,N_306,In_425);
or U402 (N_402,N_169,N_17);
nor U403 (N_403,N_309,In_276);
xor U404 (N_404,N_329,N_348);
and U405 (N_405,N_337,In_397);
or U406 (N_406,N_257,N_353);
or U407 (N_407,N_213,N_260);
xor U408 (N_408,N_339,In_72);
nor U409 (N_409,N_250,N_326);
nand U410 (N_410,N_163,In_325);
or U411 (N_411,N_207,N_269);
nand U412 (N_412,In_363,In_113);
xor U413 (N_413,In_292,N_154);
nor U414 (N_414,N_324,N_229);
xnor U415 (N_415,N_161,In_405);
or U416 (N_416,N_302,N_359);
and U417 (N_417,N_343,N_198);
or U418 (N_418,N_345,N_358);
nand U419 (N_419,N_288,In_180);
or U420 (N_420,N_299,N_136);
or U421 (N_421,N_397,N_417);
xor U422 (N_422,N_303,N_403);
nand U423 (N_423,N_376,N_350);
nor U424 (N_424,N_377,N_285);
and U425 (N_425,N_373,N_363);
and U426 (N_426,N_388,N_406);
and U427 (N_427,N_362,N_412);
nand U428 (N_428,N_378,N_201);
nand U429 (N_429,N_416,N_402);
nand U430 (N_430,N_413,N_386);
nand U431 (N_431,N_414,N_367);
nor U432 (N_432,N_383,N_387);
xor U433 (N_433,N_366,N_401);
or U434 (N_434,N_380,N_398);
nor U435 (N_435,N_385,N_365);
nor U436 (N_436,N_364,N_384);
and U437 (N_437,N_360,N_379);
nor U438 (N_438,N_407,N_381);
and U439 (N_439,N_214,N_361);
xor U440 (N_440,N_399,N_409);
nor U441 (N_441,N_390,N_333);
nand U442 (N_442,N_371,N_346);
and U443 (N_443,N_415,N_404);
xnor U444 (N_444,N_396,N_308);
xor U445 (N_445,N_405,N_411);
and U446 (N_446,N_393,N_410);
xnor U447 (N_447,N_375,N_400);
nor U448 (N_448,N_392,N_370);
and U449 (N_449,N_307,N_293);
and U450 (N_450,N_419,N_301);
nor U451 (N_451,N_369,N_408);
nand U452 (N_452,N_382,N_334);
nand U453 (N_453,N_286,N_389);
nor U454 (N_454,N_391,N_338);
nand U455 (N_455,N_395,N_368);
nor U456 (N_456,N_374,N_152);
nor U457 (N_457,N_418,N_320);
xor U458 (N_458,N_394,N_216);
and U459 (N_459,N_190,N_372);
or U460 (N_460,N_346,N_402);
xor U461 (N_461,N_365,N_369);
nand U462 (N_462,N_363,N_299);
and U463 (N_463,N_136,N_391);
or U464 (N_464,N_363,N_385);
and U465 (N_465,N_293,N_405);
and U466 (N_466,N_301,N_385);
xor U467 (N_467,N_408,N_393);
nand U468 (N_468,N_370,N_405);
and U469 (N_469,N_385,N_377);
nor U470 (N_470,N_379,N_381);
and U471 (N_471,N_362,N_365);
nand U472 (N_472,N_372,N_410);
or U473 (N_473,N_299,N_395);
nor U474 (N_474,N_416,N_368);
and U475 (N_475,N_412,N_384);
xor U476 (N_476,N_376,N_375);
xnor U477 (N_477,N_366,N_365);
nor U478 (N_478,N_407,N_405);
nor U479 (N_479,N_152,N_386);
or U480 (N_480,N_443,N_431);
and U481 (N_481,N_467,N_427);
and U482 (N_482,N_424,N_421);
nand U483 (N_483,N_454,N_470);
nor U484 (N_484,N_471,N_465);
nand U485 (N_485,N_448,N_449);
nand U486 (N_486,N_458,N_441);
and U487 (N_487,N_450,N_428);
nor U488 (N_488,N_457,N_456);
or U489 (N_489,N_436,N_451);
or U490 (N_490,N_460,N_446);
or U491 (N_491,N_420,N_479);
and U492 (N_492,N_445,N_478);
or U493 (N_493,N_474,N_473);
and U494 (N_494,N_461,N_444);
nand U495 (N_495,N_432,N_464);
xor U496 (N_496,N_463,N_469);
xnor U497 (N_497,N_466,N_477);
and U498 (N_498,N_434,N_455);
xnor U499 (N_499,N_439,N_476);
nor U500 (N_500,N_459,N_472);
or U501 (N_501,N_442,N_452);
and U502 (N_502,N_433,N_438);
nor U503 (N_503,N_426,N_468);
and U504 (N_504,N_423,N_462);
nor U505 (N_505,N_440,N_447);
and U506 (N_506,N_422,N_453);
nand U507 (N_507,N_430,N_429);
nand U508 (N_508,N_425,N_437);
and U509 (N_509,N_435,N_475);
nand U510 (N_510,N_423,N_468);
nor U511 (N_511,N_436,N_470);
nor U512 (N_512,N_429,N_442);
or U513 (N_513,N_474,N_437);
and U514 (N_514,N_433,N_453);
xor U515 (N_515,N_438,N_432);
or U516 (N_516,N_437,N_454);
nand U517 (N_517,N_466,N_453);
and U518 (N_518,N_459,N_474);
or U519 (N_519,N_464,N_428);
nor U520 (N_520,N_444,N_428);
and U521 (N_521,N_476,N_441);
nand U522 (N_522,N_439,N_451);
or U523 (N_523,N_472,N_468);
nand U524 (N_524,N_432,N_467);
and U525 (N_525,N_424,N_434);
or U526 (N_526,N_441,N_472);
or U527 (N_527,N_448,N_474);
nand U528 (N_528,N_466,N_461);
nand U529 (N_529,N_420,N_431);
nor U530 (N_530,N_429,N_425);
and U531 (N_531,N_445,N_433);
xor U532 (N_532,N_459,N_422);
xor U533 (N_533,N_451,N_433);
and U534 (N_534,N_425,N_462);
nand U535 (N_535,N_451,N_455);
nand U536 (N_536,N_432,N_466);
or U537 (N_537,N_437,N_424);
xor U538 (N_538,N_420,N_424);
xnor U539 (N_539,N_442,N_446);
nand U540 (N_540,N_485,N_519);
nand U541 (N_541,N_534,N_508);
xor U542 (N_542,N_505,N_522);
nand U543 (N_543,N_490,N_531);
nor U544 (N_544,N_510,N_491);
xor U545 (N_545,N_489,N_492);
xnor U546 (N_546,N_501,N_530);
nor U547 (N_547,N_538,N_523);
nor U548 (N_548,N_536,N_484);
xor U549 (N_549,N_529,N_509);
nor U550 (N_550,N_488,N_498);
nor U551 (N_551,N_537,N_526);
nand U552 (N_552,N_497,N_516);
or U553 (N_553,N_483,N_524);
nand U554 (N_554,N_512,N_493);
nor U555 (N_555,N_525,N_495);
and U556 (N_556,N_539,N_500);
or U557 (N_557,N_513,N_496);
and U558 (N_558,N_521,N_481);
xnor U559 (N_559,N_527,N_502);
xor U560 (N_560,N_518,N_487);
nand U561 (N_561,N_507,N_533);
and U562 (N_562,N_506,N_480);
and U563 (N_563,N_494,N_482);
nand U564 (N_564,N_486,N_504);
and U565 (N_565,N_517,N_532);
and U566 (N_566,N_535,N_528);
nand U567 (N_567,N_515,N_503);
nor U568 (N_568,N_511,N_514);
nor U569 (N_569,N_499,N_520);
xnor U570 (N_570,N_494,N_502);
or U571 (N_571,N_532,N_499);
xor U572 (N_572,N_517,N_505);
nand U573 (N_573,N_517,N_535);
or U574 (N_574,N_515,N_500);
nand U575 (N_575,N_499,N_513);
nor U576 (N_576,N_483,N_526);
and U577 (N_577,N_482,N_487);
xor U578 (N_578,N_529,N_510);
nor U579 (N_579,N_499,N_502);
or U580 (N_580,N_496,N_480);
xnor U581 (N_581,N_517,N_527);
nor U582 (N_582,N_498,N_535);
xnor U583 (N_583,N_497,N_486);
nor U584 (N_584,N_531,N_520);
and U585 (N_585,N_522,N_509);
or U586 (N_586,N_514,N_527);
nand U587 (N_587,N_513,N_511);
nor U588 (N_588,N_514,N_488);
nor U589 (N_589,N_525,N_493);
or U590 (N_590,N_501,N_528);
xnor U591 (N_591,N_529,N_499);
nand U592 (N_592,N_510,N_487);
nor U593 (N_593,N_531,N_491);
nor U594 (N_594,N_502,N_503);
nor U595 (N_595,N_491,N_537);
or U596 (N_596,N_518,N_530);
and U597 (N_597,N_493,N_517);
and U598 (N_598,N_527,N_488);
nand U599 (N_599,N_521,N_505);
nor U600 (N_600,N_585,N_594);
or U601 (N_601,N_593,N_598);
or U602 (N_602,N_553,N_583);
nor U603 (N_603,N_540,N_587);
and U604 (N_604,N_564,N_554);
xor U605 (N_605,N_550,N_542);
or U606 (N_606,N_546,N_590);
or U607 (N_607,N_552,N_575);
nand U608 (N_608,N_571,N_563);
and U609 (N_609,N_566,N_541);
and U610 (N_610,N_597,N_544);
and U611 (N_611,N_577,N_570);
nor U612 (N_612,N_548,N_574);
nor U613 (N_613,N_588,N_586);
and U614 (N_614,N_591,N_579);
nor U615 (N_615,N_565,N_547);
nor U616 (N_616,N_569,N_551);
nand U617 (N_617,N_560,N_562);
or U618 (N_618,N_589,N_576);
nor U619 (N_619,N_578,N_596);
xnor U620 (N_620,N_581,N_561);
or U621 (N_621,N_582,N_580);
nand U622 (N_622,N_545,N_556);
and U623 (N_623,N_558,N_572);
or U624 (N_624,N_557,N_549);
nor U625 (N_625,N_592,N_573);
or U626 (N_626,N_568,N_555);
nand U627 (N_627,N_543,N_559);
or U628 (N_628,N_584,N_595);
and U629 (N_629,N_567,N_599);
nand U630 (N_630,N_573,N_580);
xor U631 (N_631,N_544,N_583);
nor U632 (N_632,N_544,N_551);
and U633 (N_633,N_553,N_585);
nand U634 (N_634,N_588,N_581);
xnor U635 (N_635,N_572,N_595);
nand U636 (N_636,N_549,N_592);
or U637 (N_637,N_590,N_544);
nor U638 (N_638,N_558,N_555);
nand U639 (N_639,N_572,N_551);
nand U640 (N_640,N_560,N_544);
and U641 (N_641,N_550,N_549);
or U642 (N_642,N_591,N_571);
and U643 (N_643,N_572,N_588);
nand U644 (N_644,N_594,N_558);
nor U645 (N_645,N_540,N_565);
xor U646 (N_646,N_540,N_599);
and U647 (N_647,N_568,N_591);
nand U648 (N_648,N_595,N_588);
nor U649 (N_649,N_593,N_586);
xor U650 (N_650,N_598,N_588);
nor U651 (N_651,N_547,N_544);
nand U652 (N_652,N_598,N_597);
and U653 (N_653,N_596,N_585);
xnor U654 (N_654,N_557,N_592);
nor U655 (N_655,N_590,N_597);
nor U656 (N_656,N_588,N_545);
nand U657 (N_657,N_568,N_562);
nor U658 (N_658,N_587,N_580);
or U659 (N_659,N_553,N_592);
xnor U660 (N_660,N_634,N_655);
nand U661 (N_661,N_625,N_632);
xor U662 (N_662,N_603,N_600);
nand U663 (N_663,N_647,N_631);
or U664 (N_664,N_635,N_642);
and U665 (N_665,N_601,N_636);
nand U666 (N_666,N_633,N_628);
and U667 (N_667,N_630,N_654);
or U668 (N_668,N_639,N_650);
nor U669 (N_669,N_611,N_651);
nand U670 (N_670,N_604,N_622);
and U671 (N_671,N_614,N_606);
xnor U672 (N_672,N_627,N_644);
nand U673 (N_673,N_623,N_609);
and U674 (N_674,N_615,N_649);
or U675 (N_675,N_619,N_610);
xnor U676 (N_676,N_617,N_659);
and U677 (N_677,N_637,N_620);
nor U678 (N_678,N_657,N_626);
or U679 (N_679,N_645,N_638);
and U680 (N_680,N_643,N_612);
nor U681 (N_681,N_656,N_621);
nand U682 (N_682,N_616,N_629);
or U683 (N_683,N_648,N_602);
and U684 (N_684,N_653,N_640);
xnor U685 (N_685,N_618,N_641);
nor U686 (N_686,N_652,N_613);
and U687 (N_687,N_605,N_624);
nand U688 (N_688,N_646,N_607);
or U689 (N_689,N_658,N_608);
and U690 (N_690,N_603,N_636);
nor U691 (N_691,N_646,N_610);
and U692 (N_692,N_620,N_654);
or U693 (N_693,N_621,N_633);
xor U694 (N_694,N_650,N_602);
nor U695 (N_695,N_602,N_616);
nor U696 (N_696,N_601,N_606);
or U697 (N_697,N_639,N_629);
nor U698 (N_698,N_634,N_651);
xor U699 (N_699,N_614,N_629);
nand U700 (N_700,N_625,N_627);
nand U701 (N_701,N_604,N_651);
nor U702 (N_702,N_615,N_625);
nand U703 (N_703,N_657,N_651);
nand U704 (N_704,N_627,N_604);
and U705 (N_705,N_621,N_627);
or U706 (N_706,N_659,N_651);
xnor U707 (N_707,N_619,N_615);
and U708 (N_708,N_606,N_611);
nor U709 (N_709,N_628,N_651);
xnor U710 (N_710,N_608,N_638);
nor U711 (N_711,N_658,N_632);
nor U712 (N_712,N_604,N_612);
or U713 (N_713,N_632,N_609);
or U714 (N_714,N_632,N_638);
xnor U715 (N_715,N_620,N_629);
and U716 (N_716,N_605,N_639);
nand U717 (N_717,N_628,N_615);
or U718 (N_718,N_612,N_624);
or U719 (N_719,N_659,N_650);
or U720 (N_720,N_714,N_697);
or U721 (N_721,N_710,N_687);
or U722 (N_722,N_698,N_713);
xor U723 (N_723,N_684,N_695);
xor U724 (N_724,N_715,N_705);
xor U725 (N_725,N_692,N_699);
and U726 (N_726,N_675,N_669);
nand U727 (N_727,N_700,N_676);
and U728 (N_728,N_677,N_685);
nand U729 (N_729,N_711,N_666);
or U730 (N_730,N_668,N_702);
nand U731 (N_731,N_662,N_663);
or U732 (N_732,N_706,N_712);
xor U733 (N_733,N_673,N_696);
nor U734 (N_734,N_661,N_689);
nor U735 (N_735,N_694,N_701);
or U736 (N_736,N_709,N_717);
and U737 (N_737,N_718,N_704);
or U738 (N_738,N_708,N_707);
or U739 (N_739,N_719,N_679);
nand U740 (N_740,N_681,N_660);
nor U741 (N_741,N_680,N_672);
nor U742 (N_742,N_665,N_678);
nand U743 (N_743,N_690,N_667);
nor U744 (N_744,N_683,N_716);
nor U745 (N_745,N_703,N_688);
or U746 (N_746,N_670,N_691);
nand U747 (N_747,N_693,N_674);
nor U748 (N_748,N_682,N_686);
nand U749 (N_749,N_671,N_664);
or U750 (N_750,N_701,N_673);
xor U751 (N_751,N_676,N_673);
xnor U752 (N_752,N_688,N_714);
nor U753 (N_753,N_710,N_671);
nand U754 (N_754,N_662,N_707);
xor U755 (N_755,N_698,N_678);
or U756 (N_756,N_717,N_671);
xnor U757 (N_757,N_665,N_704);
or U758 (N_758,N_708,N_704);
nor U759 (N_759,N_710,N_701);
nand U760 (N_760,N_700,N_661);
or U761 (N_761,N_675,N_673);
and U762 (N_762,N_675,N_666);
or U763 (N_763,N_664,N_695);
xor U764 (N_764,N_705,N_692);
xnor U765 (N_765,N_716,N_713);
nand U766 (N_766,N_696,N_694);
xnor U767 (N_767,N_719,N_702);
or U768 (N_768,N_671,N_675);
nand U769 (N_769,N_683,N_665);
xnor U770 (N_770,N_661,N_715);
and U771 (N_771,N_694,N_709);
or U772 (N_772,N_669,N_712);
or U773 (N_773,N_684,N_660);
and U774 (N_774,N_686,N_664);
and U775 (N_775,N_672,N_716);
or U776 (N_776,N_717,N_683);
nand U777 (N_777,N_680,N_664);
or U778 (N_778,N_691,N_669);
nor U779 (N_779,N_690,N_704);
and U780 (N_780,N_752,N_732);
nor U781 (N_781,N_776,N_773);
xnor U782 (N_782,N_777,N_762);
xor U783 (N_783,N_770,N_765);
and U784 (N_784,N_729,N_735);
or U785 (N_785,N_748,N_728);
and U786 (N_786,N_760,N_774);
or U787 (N_787,N_767,N_775);
and U788 (N_788,N_727,N_757);
or U789 (N_789,N_740,N_768);
xnor U790 (N_790,N_736,N_763);
nand U791 (N_791,N_723,N_720);
xor U792 (N_792,N_741,N_749);
xnor U793 (N_793,N_738,N_764);
nand U794 (N_794,N_724,N_761);
and U795 (N_795,N_769,N_746);
and U796 (N_796,N_734,N_751);
and U797 (N_797,N_756,N_772);
nand U798 (N_798,N_753,N_745);
nor U799 (N_799,N_742,N_725);
and U800 (N_800,N_759,N_737);
or U801 (N_801,N_758,N_744);
nand U802 (N_802,N_739,N_747);
and U803 (N_803,N_733,N_754);
and U804 (N_804,N_730,N_743);
nand U805 (N_805,N_750,N_771);
xnor U806 (N_806,N_766,N_778);
nand U807 (N_807,N_721,N_755);
nand U808 (N_808,N_726,N_731);
xor U809 (N_809,N_779,N_722);
and U810 (N_810,N_764,N_723);
xor U811 (N_811,N_747,N_766);
or U812 (N_812,N_755,N_773);
or U813 (N_813,N_768,N_743);
or U814 (N_814,N_730,N_745);
and U815 (N_815,N_749,N_779);
nand U816 (N_816,N_736,N_766);
nor U817 (N_817,N_737,N_731);
or U818 (N_818,N_760,N_752);
and U819 (N_819,N_722,N_731);
xnor U820 (N_820,N_721,N_776);
nor U821 (N_821,N_763,N_766);
nand U822 (N_822,N_721,N_730);
xor U823 (N_823,N_775,N_725);
nand U824 (N_824,N_730,N_765);
or U825 (N_825,N_749,N_721);
or U826 (N_826,N_778,N_747);
nand U827 (N_827,N_778,N_740);
and U828 (N_828,N_728,N_758);
xnor U829 (N_829,N_742,N_758);
xnor U830 (N_830,N_755,N_778);
nand U831 (N_831,N_768,N_739);
or U832 (N_832,N_778,N_768);
or U833 (N_833,N_775,N_761);
nand U834 (N_834,N_752,N_736);
nand U835 (N_835,N_735,N_753);
nand U836 (N_836,N_735,N_764);
nor U837 (N_837,N_743,N_722);
nand U838 (N_838,N_741,N_757);
xor U839 (N_839,N_767,N_756);
xor U840 (N_840,N_801,N_820);
xnor U841 (N_841,N_785,N_838);
and U842 (N_842,N_825,N_806);
or U843 (N_843,N_802,N_831);
and U844 (N_844,N_791,N_827);
or U845 (N_845,N_794,N_826);
and U846 (N_846,N_834,N_811);
or U847 (N_847,N_807,N_823);
or U848 (N_848,N_783,N_809);
nor U849 (N_849,N_835,N_786);
nand U850 (N_850,N_788,N_790);
nor U851 (N_851,N_832,N_822);
or U852 (N_852,N_810,N_793);
or U853 (N_853,N_839,N_833);
nor U854 (N_854,N_816,N_828);
nand U855 (N_855,N_819,N_813);
nand U856 (N_856,N_817,N_797);
nand U857 (N_857,N_792,N_780);
nor U858 (N_858,N_815,N_836);
nor U859 (N_859,N_789,N_829);
nor U860 (N_860,N_818,N_837);
or U861 (N_861,N_812,N_795);
and U862 (N_862,N_814,N_830);
and U863 (N_863,N_821,N_781);
nand U864 (N_864,N_804,N_803);
xnor U865 (N_865,N_808,N_782);
or U866 (N_866,N_787,N_799);
xnor U867 (N_867,N_800,N_805);
or U868 (N_868,N_824,N_798);
and U869 (N_869,N_796,N_784);
and U870 (N_870,N_812,N_825);
nor U871 (N_871,N_809,N_829);
or U872 (N_872,N_827,N_786);
nand U873 (N_873,N_803,N_815);
nand U874 (N_874,N_788,N_809);
and U875 (N_875,N_782,N_793);
nor U876 (N_876,N_783,N_822);
nor U877 (N_877,N_790,N_821);
and U878 (N_878,N_802,N_835);
or U879 (N_879,N_789,N_795);
and U880 (N_880,N_828,N_810);
and U881 (N_881,N_818,N_806);
xnor U882 (N_882,N_780,N_830);
xnor U883 (N_883,N_816,N_823);
or U884 (N_884,N_828,N_792);
and U885 (N_885,N_828,N_826);
and U886 (N_886,N_822,N_801);
nor U887 (N_887,N_781,N_804);
nor U888 (N_888,N_793,N_790);
or U889 (N_889,N_823,N_797);
or U890 (N_890,N_802,N_833);
nor U891 (N_891,N_809,N_837);
xor U892 (N_892,N_830,N_803);
xor U893 (N_893,N_808,N_790);
xnor U894 (N_894,N_802,N_829);
nor U895 (N_895,N_809,N_813);
and U896 (N_896,N_799,N_783);
nand U897 (N_897,N_813,N_839);
or U898 (N_898,N_788,N_823);
nor U899 (N_899,N_794,N_786);
xnor U900 (N_900,N_874,N_854);
and U901 (N_901,N_845,N_865);
xor U902 (N_902,N_844,N_849);
xnor U903 (N_903,N_856,N_841);
nand U904 (N_904,N_869,N_846);
and U905 (N_905,N_840,N_842);
and U906 (N_906,N_866,N_864);
nand U907 (N_907,N_872,N_882);
nor U908 (N_908,N_859,N_892);
nor U909 (N_909,N_861,N_878);
or U910 (N_910,N_867,N_858);
nor U911 (N_911,N_852,N_868);
or U912 (N_912,N_877,N_895);
xor U913 (N_913,N_875,N_851);
or U914 (N_914,N_863,N_894);
and U915 (N_915,N_857,N_898);
nor U916 (N_916,N_876,N_873);
nor U917 (N_917,N_885,N_890);
or U918 (N_918,N_884,N_893);
xor U919 (N_919,N_886,N_891);
nand U920 (N_920,N_899,N_881);
xnor U921 (N_921,N_870,N_880);
or U922 (N_922,N_843,N_879);
nor U923 (N_923,N_896,N_853);
and U924 (N_924,N_847,N_871);
or U925 (N_925,N_848,N_883);
and U926 (N_926,N_889,N_855);
nor U927 (N_927,N_888,N_887);
nand U928 (N_928,N_862,N_860);
or U929 (N_929,N_850,N_897);
nor U930 (N_930,N_898,N_883);
or U931 (N_931,N_883,N_893);
xor U932 (N_932,N_864,N_848);
and U933 (N_933,N_894,N_892);
xnor U934 (N_934,N_895,N_844);
nor U935 (N_935,N_868,N_846);
and U936 (N_936,N_861,N_876);
and U937 (N_937,N_845,N_878);
and U938 (N_938,N_899,N_887);
or U939 (N_939,N_897,N_852);
and U940 (N_940,N_895,N_886);
nor U941 (N_941,N_846,N_885);
and U942 (N_942,N_860,N_863);
and U943 (N_943,N_899,N_840);
nor U944 (N_944,N_841,N_873);
or U945 (N_945,N_849,N_840);
xnor U946 (N_946,N_862,N_876);
nand U947 (N_947,N_841,N_842);
or U948 (N_948,N_844,N_851);
and U949 (N_949,N_851,N_894);
and U950 (N_950,N_840,N_883);
or U951 (N_951,N_866,N_880);
or U952 (N_952,N_873,N_850);
xor U953 (N_953,N_874,N_884);
or U954 (N_954,N_844,N_843);
xnor U955 (N_955,N_878,N_897);
and U956 (N_956,N_870,N_859);
xnor U957 (N_957,N_878,N_868);
and U958 (N_958,N_876,N_855);
xor U959 (N_959,N_841,N_861);
or U960 (N_960,N_949,N_921);
nor U961 (N_961,N_903,N_936);
and U962 (N_962,N_917,N_944);
xnor U963 (N_963,N_905,N_918);
nand U964 (N_964,N_934,N_907);
nor U965 (N_965,N_908,N_932);
or U966 (N_966,N_922,N_926);
nor U967 (N_967,N_928,N_909);
and U968 (N_968,N_939,N_940);
xor U969 (N_969,N_900,N_933);
nand U970 (N_970,N_942,N_919);
and U971 (N_971,N_916,N_947);
and U972 (N_972,N_902,N_952);
or U973 (N_973,N_911,N_937);
nand U974 (N_974,N_957,N_956);
xnor U975 (N_975,N_954,N_935);
or U976 (N_976,N_953,N_938);
or U977 (N_977,N_931,N_913);
or U978 (N_978,N_914,N_906);
xnor U979 (N_979,N_951,N_930);
or U980 (N_980,N_950,N_901);
xor U981 (N_981,N_915,N_910);
nand U982 (N_982,N_925,N_948);
or U983 (N_983,N_920,N_941);
or U984 (N_984,N_904,N_924);
or U985 (N_985,N_943,N_945);
xnor U986 (N_986,N_959,N_923);
xor U987 (N_987,N_958,N_927);
nand U988 (N_988,N_929,N_946);
nand U989 (N_989,N_912,N_955);
nor U990 (N_990,N_953,N_951);
xor U991 (N_991,N_948,N_922);
or U992 (N_992,N_958,N_955);
xor U993 (N_993,N_909,N_938);
nor U994 (N_994,N_922,N_953);
or U995 (N_995,N_920,N_915);
nor U996 (N_996,N_949,N_904);
nor U997 (N_997,N_952,N_957);
nor U998 (N_998,N_905,N_908);
or U999 (N_999,N_914,N_920);
nor U1000 (N_1000,N_953,N_909);
or U1001 (N_1001,N_908,N_927);
xnor U1002 (N_1002,N_919,N_914);
nor U1003 (N_1003,N_903,N_939);
and U1004 (N_1004,N_952,N_951);
xnor U1005 (N_1005,N_942,N_954);
nand U1006 (N_1006,N_919,N_907);
or U1007 (N_1007,N_946,N_944);
xnor U1008 (N_1008,N_912,N_909);
and U1009 (N_1009,N_944,N_932);
or U1010 (N_1010,N_925,N_934);
nor U1011 (N_1011,N_913,N_935);
xnor U1012 (N_1012,N_903,N_924);
nand U1013 (N_1013,N_956,N_934);
nand U1014 (N_1014,N_947,N_942);
or U1015 (N_1015,N_903,N_944);
nand U1016 (N_1016,N_914,N_958);
and U1017 (N_1017,N_909,N_903);
and U1018 (N_1018,N_912,N_906);
nor U1019 (N_1019,N_932,N_905);
nand U1020 (N_1020,N_1014,N_1018);
nor U1021 (N_1021,N_961,N_1019);
or U1022 (N_1022,N_995,N_985);
nor U1023 (N_1023,N_980,N_977);
nor U1024 (N_1024,N_971,N_1002);
and U1025 (N_1025,N_968,N_997);
nor U1026 (N_1026,N_982,N_1009);
or U1027 (N_1027,N_976,N_970);
nor U1028 (N_1028,N_967,N_996);
or U1029 (N_1029,N_1003,N_972);
nor U1030 (N_1030,N_962,N_1006);
xnor U1031 (N_1031,N_974,N_983);
nor U1032 (N_1032,N_991,N_1015);
or U1033 (N_1033,N_979,N_981);
nand U1034 (N_1034,N_1008,N_964);
xor U1035 (N_1035,N_1012,N_986);
nand U1036 (N_1036,N_978,N_960);
nand U1037 (N_1037,N_963,N_1000);
nand U1038 (N_1038,N_1016,N_992);
and U1039 (N_1039,N_999,N_1011);
xnor U1040 (N_1040,N_989,N_1013);
nand U1041 (N_1041,N_969,N_988);
nor U1042 (N_1042,N_975,N_998);
or U1043 (N_1043,N_973,N_965);
nand U1044 (N_1044,N_1007,N_987);
xor U1045 (N_1045,N_1005,N_994);
nor U1046 (N_1046,N_1010,N_1004);
xnor U1047 (N_1047,N_1001,N_990);
nor U1048 (N_1048,N_984,N_1017);
xnor U1049 (N_1049,N_993,N_966);
xor U1050 (N_1050,N_983,N_999);
xnor U1051 (N_1051,N_1000,N_981);
and U1052 (N_1052,N_996,N_966);
xnor U1053 (N_1053,N_971,N_981);
nand U1054 (N_1054,N_964,N_985);
or U1055 (N_1055,N_988,N_964);
nand U1056 (N_1056,N_979,N_1018);
nor U1057 (N_1057,N_1016,N_1015);
xnor U1058 (N_1058,N_976,N_981);
xnor U1059 (N_1059,N_975,N_982);
and U1060 (N_1060,N_984,N_1003);
and U1061 (N_1061,N_1003,N_1012);
and U1062 (N_1062,N_1002,N_987);
or U1063 (N_1063,N_964,N_984);
nand U1064 (N_1064,N_1009,N_975);
or U1065 (N_1065,N_1003,N_999);
nand U1066 (N_1066,N_995,N_1017);
nand U1067 (N_1067,N_1004,N_966);
or U1068 (N_1068,N_983,N_965);
xnor U1069 (N_1069,N_968,N_967);
nor U1070 (N_1070,N_962,N_978);
nor U1071 (N_1071,N_1006,N_1018);
nand U1072 (N_1072,N_1002,N_980);
xnor U1073 (N_1073,N_1013,N_990);
xor U1074 (N_1074,N_961,N_987);
nand U1075 (N_1075,N_994,N_992);
and U1076 (N_1076,N_993,N_965);
and U1077 (N_1077,N_1009,N_997);
and U1078 (N_1078,N_974,N_1001);
nand U1079 (N_1079,N_1019,N_995);
or U1080 (N_1080,N_1023,N_1079);
or U1081 (N_1081,N_1054,N_1031);
nor U1082 (N_1082,N_1052,N_1061);
or U1083 (N_1083,N_1057,N_1043);
xnor U1084 (N_1084,N_1053,N_1041);
xor U1085 (N_1085,N_1065,N_1030);
xor U1086 (N_1086,N_1074,N_1076);
and U1087 (N_1087,N_1062,N_1042);
xor U1088 (N_1088,N_1046,N_1067);
nor U1089 (N_1089,N_1032,N_1044);
xnor U1090 (N_1090,N_1049,N_1026);
xnor U1091 (N_1091,N_1070,N_1068);
and U1092 (N_1092,N_1077,N_1047);
or U1093 (N_1093,N_1075,N_1063);
xor U1094 (N_1094,N_1073,N_1037);
nand U1095 (N_1095,N_1078,N_1025);
xnor U1096 (N_1096,N_1071,N_1036);
nand U1097 (N_1097,N_1039,N_1028);
nor U1098 (N_1098,N_1034,N_1027);
and U1099 (N_1099,N_1045,N_1058);
nor U1100 (N_1100,N_1035,N_1060);
nand U1101 (N_1101,N_1059,N_1021);
nor U1102 (N_1102,N_1020,N_1022);
and U1103 (N_1103,N_1048,N_1066);
xnor U1104 (N_1104,N_1029,N_1033);
xor U1105 (N_1105,N_1069,N_1050);
or U1106 (N_1106,N_1055,N_1051);
xnor U1107 (N_1107,N_1072,N_1038);
nand U1108 (N_1108,N_1064,N_1040);
or U1109 (N_1109,N_1024,N_1056);
nand U1110 (N_1110,N_1057,N_1062);
xor U1111 (N_1111,N_1068,N_1032);
or U1112 (N_1112,N_1049,N_1025);
xor U1113 (N_1113,N_1075,N_1045);
nand U1114 (N_1114,N_1051,N_1024);
nand U1115 (N_1115,N_1021,N_1039);
or U1116 (N_1116,N_1049,N_1043);
and U1117 (N_1117,N_1046,N_1048);
nand U1118 (N_1118,N_1053,N_1023);
nand U1119 (N_1119,N_1055,N_1034);
nand U1120 (N_1120,N_1057,N_1074);
xnor U1121 (N_1121,N_1042,N_1036);
or U1122 (N_1122,N_1036,N_1074);
nand U1123 (N_1123,N_1051,N_1031);
and U1124 (N_1124,N_1058,N_1050);
and U1125 (N_1125,N_1074,N_1071);
nand U1126 (N_1126,N_1041,N_1070);
and U1127 (N_1127,N_1039,N_1075);
nor U1128 (N_1128,N_1034,N_1033);
xor U1129 (N_1129,N_1053,N_1068);
nand U1130 (N_1130,N_1040,N_1054);
xor U1131 (N_1131,N_1025,N_1068);
xnor U1132 (N_1132,N_1068,N_1030);
and U1133 (N_1133,N_1052,N_1047);
nor U1134 (N_1134,N_1045,N_1054);
nor U1135 (N_1135,N_1026,N_1078);
nand U1136 (N_1136,N_1073,N_1022);
or U1137 (N_1137,N_1078,N_1079);
nand U1138 (N_1138,N_1067,N_1058);
nand U1139 (N_1139,N_1079,N_1038);
xnor U1140 (N_1140,N_1114,N_1132);
xor U1141 (N_1141,N_1122,N_1104);
nand U1142 (N_1142,N_1097,N_1111);
or U1143 (N_1143,N_1115,N_1089);
and U1144 (N_1144,N_1110,N_1101);
nor U1145 (N_1145,N_1087,N_1092);
nand U1146 (N_1146,N_1098,N_1085);
and U1147 (N_1147,N_1088,N_1127);
nor U1148 (N_1148,N_1094,N_1082);
or U1149 (N_1149,N_1096,N_1125);
xor U1150 (N_1150,N_1138,N_1126);
or U1151 (N_1151,N_1102,N_1113);
or U1152 (N_1152,N_1095,N_1100);
nor U1153 (N_1153,N_1128,N_1124);
or U1154 (N_1154,N_1107,N_1105);
and U1155 (N_1155,N_1131,N_1103);
and U1156 (N_1156,N_1135,N_1109);
xor U1157 (N_1157,N_1137,N_1099);
nor U1158 (N_1158,N_1106,N_1119);
nor U1159 (N_1159,N_1129,N_1091);
or U1160 (N_1160,N_1139,N_1136);
nand U1161 (N_1161,N_1130,N_1123);
nand U1162 (N_1162,N_1090,N_1133);
nand U1163 (N_1163,N_1086,N_1083);
xnor U1164 (N_1164,N_1116,N_1081);
nand U1165 (N_1165,N_1117,N_1093);
or U1166 (N_1166,N_1120,N_1118);
or U1167 (N_1167,N_1108,N_1121);
or U1168 (N_1168,N_1112,N_1134);
and U1169 (N_1169,N_1084,N_1080);
and U1170 (N_1170,N_1128,N_1131);
xnor U1171 (N_1171,N_1138,N_1112);
or U1172 (N_1172,N_1090,N_1082);
or U1173 (N_1173,N_1110,N_1083);
xor U1174 (N_1174,N_1106,N_1108);
nor U1175 (N_1175,N_1091,N_1090);
and U1176 (N_1176,N_1112,N_1100);
and U1177 (N_1177,N_1098,N_1123);
and U1178 (N_1178,N_1084,N_1088);
or U1179 (N_1179,N_1085,N_1095);
or U1180 (N_1180,N_1121,N_1101);
nor U1181 (N_1181,N_1114,N_1098);
nor U1182 (N_1182,N_1089,N_1082);
nand U1183 (N_1183,N_1095,N_1110);
nand U1184 (N_1184,N_1091,N_1130);
xnor U1185 (N_1185,N_1116,N_1133);
and U1186 (N_1186,N_1096,N_1083);
nor U1187 (N_1187,N_1100,N_1117);
nor U1188 (N_1188,N_1129,N_1096);
or U1189 (N_1189,N_1111,N_1119);
nand U1190 (N_1190,N_1121,N_1109);
and U1191 (N_1191,N_1105,N_1111);
nand U1192 (N_1192,N_1114,N_1106);
nand U1193 (N_1193,N_1115,N_1082);
or U1194 (N_1194,N_1114,N_1105);
or U1195 (N_1195,N_1081,N_1133);
xnor U1196 (N_1196,N_1138,N_1106);
or U1197 (N_1197,N_1121,N_1084);
and U1198 (N_1198,N_1124,N_1135);
nor U1199 (N_1199,N_1089,N_1114);
nand U1200 (N_1200,N_1142,N_1170);
xnor U1201 (N_1201,N_1145,N_1166);
xor U1202 (N_1202,N_1187,N_1197);
or U1203 (N_1203,N_1154,N_1140);
and U1204 (N_1204,N_1198,N_1188);
and U1205 (N_1205,N_1184,N_1161);
and U1206 (N_1206,N_1165,N_1143);
and U1207 (N_1207,N_1158,N_1156);
and U1208 (N_1208,N_1148,N_1159);
or U1209 (N_1209,N_1179,N_1153);
xor U1210 (N_1210,N_1151,N_1168);
xor U1211 (N_1211,N_1174,N_1194);
nand U1212 (N_1212,N_1164,N_1175);
xor U1213 (N_1213,N_1163,N_1191);
and U1214 (N_1214,N_1171,N_1155);
nor U1215 (N_1215,N_1199,N_1150);
xor U1216 (N_1216,N_1169,N_1183);
xor U1217 (N_1217,N_1172,N_1192);
nor U1218 (N_1218,N_1178,N_1149);
or U1219 (N_1219,N_1176,N_1196);
nand U1220 (N_1220,N_1173,N_1181);
nand U1221 (N_1221,N_1144,N_1177);
or U1222 (N_1222,N_1157,N_1189);
nand U1223 (N_1223,N_1141,N_1182);
xor U1224 (N_1224,N_1167,N_1190);
and U1225 (N_1225,N_1193,N_1162);
or U1226 (N_1226,N_1147,N_1180);
and U1227 (N_1227,N_1185,N_1186);
nor U1228 (N_1228,N_1195,N_1146);
and U1229 (N_1229,N_1152,N_1160);
or U1230 (N_1230,N_1163,N_1169);
or U1231 (N_1231,N_1195,N_1168);
and U1232 (N_1232,N_1187,N_1176);
and U1233 (N_1233,N_1140,N_1182);
nand U1234 (N_1234,N_1173,N_1192);
nand U1235 (N_1235,N_1170,N_1152);
xnor U1236 (N_1236,N_1196,N_1179);
nand U1237 (N_1237,N_1143,N_1188);
and U1238 (N_1238,N_1198,N_1186);
nand U1239 (N_1239,N_1194,N_1148);
nor U1240 (N_1240,N_1144,N_1172);
xor U1241 (N_1241,N_1149,N_1174);
xor U1242 (N_1242,N_1183,N_1143);
xor U1243 (N_1243,N_1194,N_1153);
or U1244 (N_1244,N_1180,N_1150);
nor U1245 (N_1245,N_1141,N_1196);
and U1246 (N_1246,N_1161,N_1190);
nor U1247 (N_1247,N_1157,N_1186);
nor U1248 (N_1248,N_1181,N_1166);
xnor U1249 (N_1249,N_1193,N_1178);
nor U1250 (N_1250,N_1199,N_1142);
xor U1251 (N_1251,N_1178,N_1144);
or U1252 (N_1252,N_1147,N_1145);
xnor U1253 (N_1253,N_1197,N_1141);
or U1254 (N_1254,N_1189,N_1145);
and U1255 (N_1255,N_1193,N_1197);
and U1256 (N_1256,N_1175,N_1171);
and U1257 (N_1257,N_1173,N_1186);
nor U1258 (N_1258,N_1162,N_1147);
xor U1259 (N_1259,N_1153,N_1168);
nor U1260 (N_1260,N_1247,N_1216);
and U1261 (N_1261,N_1236,N_1257);
xor U1262 (N_1262,N_1258,N_1254);
nand U1263 (N_1263,N_1240,N_1205);
nand U1264 (N_1264,N_1251,N_1245);
and U1265 (N_1265,N_1208,N_1204);
nand U1266 (N_1266,N_1225,N_1228);
nor U1267 (N_1267,N_1235,N_1222);
xnor U1268 (N_1268,N_1255,N_1232);
xnor U1269 (N_1269,N_1206,N_1220);
nor U1270 (N_1270,N_1234,N_1231);
xnor U1271 (N_1271,N_1248,N_1219);
and U1272 (N_1272,N_1214,N_1223);
xor U1273 (N_1273,N_1215,N_1207);
or U1274 (N_1274,N_1211,N_1202);
xnor U1275 (N_1275,N_1209,N_1256);
nand U1276 (N_1276,N_1203,N_1242);
and U1277 (N_1277,N_1229,N_1233);
and U1278 (N_1278,N_1249,N_1210);
xnor U1279 (N_1279,N_1259,N_1243);
and U1280 (N_1280,N_1213,N_1217);
and U1281 (N_1281,N_1241,N_1226);
and U1282 (N_1282,N_1244,N_1253);
xor U1283 (N_1283,N_1200,N_1239);
nand U1284 (N_1284,N_1246,N_1227);
or U1285 (N_1285,N_1237,N_1212);
xnor U1286 (N_1286,N_1250,N_1230);
or U1287 (N_1287,N_1238,N_1224);
nand U1288 (N_1288,N_1252,N_1218);
nor U1289 (N_1289,N_1221,N_1201);
xnor U1290 (N_1290,N_1256,N_1255);
nand U1291 (N_1291,N_1244,N_1240);
xnor U1292 (N_1292,N_1207,N_1259);
nand U1293 (N_1293,N_1223,N_1202);
nor U1294 (N_1294,N_1219,N_1256);
nor U1295 (N_1295,N_1253,N_1239);
or U1296 (N_1296,N_1228,N_1229);
xor U1297 (N_1297,N_1229,N_1240);
xor U1298 (N_1298,N_1236,N_1227);
and U1299 (N_1299,N_1202,N_1200);
nor U1300 (N_1300,N_1211,N_1244);
nor U1301 (N_1301,N_1209,N_1257);
xnor U1302 (N_1302,N_1231,N_1235);
nor U1303 (N_1303,N_1216,N_1217);
and U1304 (N_1304,N_1251,N_1211);
and U1305 (N_1305,N_1225,N_1236);
xnor U1306 (N_1306,N_1222,N_1255);
nand U1307 (N_1307,N_1210,N_1201);
and U1308 (N_1308,N_1244,N_1249);
and U1309 (N_1309,N_1251,N_1216);
nand U1310 (N_1310,N_1220,N_1234);
nand U1311 (N_1311,N_1226,N_1248);
nand U1312 (N_1312,N_1232,N_1233);
nor U1313 (N_1313,N_1238,N_1209);
and U1314 (N_1314,N_1209,N_1217);
xnor U1315 (N_1315,N_1215,N_1237);
and U1316 (N_1316,N_1228,N_1250);
and U1317 (N_1317,N_1256,N_1227);
and U1318 (N_1318,N_1251,N_1222);
and U1319 (N_1319,N_1207,N_1231);
nand U1320 (N_1320,N_1304,N_1302);
or U1321 (N_1321,N_1315,N_1272);
nor U1322 (N_1322,N_1296,N_1295);
or U1323 (N_1323,N_1273,N_1288);
nand U1324 (N_1324,N_1262,N_1303);
nand U1325 (N_1325,N_1301,N_1294);
xor U1326 (N_1326,N_1308,N_1261);
nand U1327 (N_1327,N_1318,N_1316);
and U1328 (N_1328,N_1263,N_1287);
and U1329 (N_1329,N_1292,N_1281);
or U1330 (N_1330,N_1310,N_1293);
xor U1331 (N_1331,N_1317,N_1299);
xnor U1332 (N_1332,N_1290,N_1275);
and U1333 (N_1333,N_1305,N_1267);
or U1334 (N_1334,N_1306,N_1282);
or U1335 (N_1335,N_1319,N_1313);
xnor U1336 (N_1336,N_1284,N_1277);
nand U1337 (N_1337,N_1297,N_1265);
nand U1338 (N_1338,N_1283,N_1269);
xnor U1339 (N_1339,N_1286,N_1307);
xnor U1340 (N_1340,N_1266,N_1309);
nor U1341 (N_1341,N_1312,N_1260);
and U1342 (N_1342,N_1314,N_1271);
xnor U1343 (N_1343,N_1298,N_1268);
or U1344 (N_1344,N_1274,N_1279);
or U1345 (N_1345,N_1285,N_1276);
xnor U1346 (N_1346,N_1300,N_1278);
nor U1347 (N_1347,N_1289,N_1280);
nand U1348 (N_1348,N_1311,N_1291);
xor U1349 (N_1349,N_1264,N_1270);
nand U1350 (N_1350,N_1266,N_1301);
or U1351 (N_1351,N_1314,N_1315);
nor U1352 (N_1352,N_1311,N_1297);
nor U1353 (N_1353,N_1270,N_1281);
and U1354 (N_1354,N_1310,N_1267);
nor U1355 (N_1355,N_1308,N_1311);
nand U1356 (N_1356,N_1271,N_1312);
xnor U1357 (N_1357,N_1261,N_1312);
and U1358 (N_1358,N_1308,N_1263);
or U1359 (N_1359,N_1314,N_1302);
and U1360 (N_1360,N_1318,N_1277);
nor U1361 (N_1361,N_1308,N_1278);
nor U1362 (N_1362,N_1314,N_1299);
and U1363 (N_1363,N_1278,N_1261);
nand U1364 (N_1364,N_1264,N_1296);
nor U1365 (N_1365,N_1278,N_1262);
nor U1366 (N_1366,N_1311,N_1312);
xor U1367 (N_1367,N_1281,N_1273);
or U1368 (N_1368,N_1289,N_1286);
and U1369 (N_1369,N_1287,N_1291);
and U1370 (N_1370,N_1268,N_1282);
nor U1371 (N_1371,N_1313,N_1296);
nand U1372 (N_1372,N_1268,N_1304);
nand U1373 (N_1373,N_1291,N_1260);
nor U1374 (N_1374,N_1298,N_1292);
nor U1375 (N_1375,N_1314,N_1306);
and U1376 (N_1376,N_1319,N_1283);
xor U1377 (N_1377,N_1271,N_1289);
or U1378 (N_1378,N_1301,N_1287);
and U1379 (N_1379,N_1305,N_1278);
nor U1380 (N_1380,N_1338,N_1369);
xnor U1381 (N_1381,N_1343,N_1371);
and U1382 (N_1382,N_1376,N_1336);
nand U1383 (N_1383,N_1366,N_1320);
and U1384 (N_1384,N_1353,N_1337);
nand U1385 (N_1385,N_1372,N_1377);
nor U1386 (N_1386,N_1325,N_1345);
nor U1387 (N_1387,N_1351,N_1355);
nor U1388 (N_1388,N_1365,N_1342);
or U1389 (N_1389,N_1326,N_1364);
and U1390 (N_1390,N_1356,N_1378);
nor U1391 (N_1391,N_1354,N_1368);
nor U1392 (N_1392,N_1344,N_1352);
and U1393 (N_1393,N_1349,N_1357);
nor U1394 (N_1394,N_1341,N_1370);
and U1395 (N_1395,N_1340,N_1339);
and U1396 (N_1396,N_1323,N_1358);
or U1397 (N_1397,N_1327,N_1322);
nand U1398 (N_1398,N_1329,N_1331);
or U1399 (N_1399,N_1328,N_1332);
or U1400 (N_1400,N_1346,N_1359);
and U1401 (N_1401,N_1347,N_1379);
or U1402 (N_1402,N_1348,N_1367);
nor U1403 (N_1403,N_1375,N_1335);
nor U1404 (N_1404,N_1350,N_1333);
or U1405 (N_1405,N_1321,N_1362);
xnor U1406 (N_1406,N_1330,N_1373);
nand U1407 (N_1407,N_1361,N_1334);
xnor U1408 (N_1408,N_1363,N_1324);
xor U1409 (N_1409,N_1374,N_1360);
or U1410 (N_1410,N_1378,N_1341);
nor U1411 (N_1411,N_1346,N_1351);
nand U1412 (N_1412,N_1337,N_1378);
and U1413 (N_1413,N_1333,N_1370);
nand U1414 (N_1414,N_1343,N_1350);
nand U1415 (N_1415,N_1356,N_1326);
and U1416 (N_1416,N_1330,N_1332);
and U1417 (N_1417,N_1336,N_1323);
nor U1418 (N_1418,N_1352,N_1356);
nor U1419 (N_1419,N_1322,N_1356);
nand U1420 (N_1420,N_1352,N_1354);
nor U1421 (N_1421,N_1364,N_1339);
and U1422 (N_1422,N_1360,N_1367);
nor U1423 (N_1423,N_1338,N_1360);
nor U1424 (N_1424,N_1374,N_1347);
and U1425 (N_1425,N_1329,N_1324);
nor U1426 (N_1426,N_1373,N_1379);
nand U1427 (N_1427,N_1363,N_1348);
nor U1428 (N_1428,N_1331,N_1375);
nor U1429 (N_1429,N_1339,N_1378);
or U1430 (N_1430,N_1324,N_1377);
nand U1431 (N_1431,N_1378,N_1325);
nor U1432 (N_1432,N_1342,N_1373);
xnor U1433 (N_1433,N_1376,N_1333);
xnor U1434 (N_1434,N_1366,N_1329);
xor U1435 (N_1435,N_1355,N_1361);
and U1436 (N_1436,N_1378,N_1368);
nor U1437 (N_1437,N_1348,N_1353);
nor U1438 (N_1438,N_1324,N_1364);
or U1439 (N_1439,N_1369,N_1349);
and U1440 (N_1440,N_1400,N_1382);
nor U1441 (N_1441,N_1407,N_1381);
nand U1442 (N_1442,N_1392,N_1427);
xnor U1443 (N_1443,N_1396,N_1393);
and U1444 (N_1444,N_1424,N_1390);
nor U1445 (N_1445,N_1437,N_1401);
nor U1446 (N_1446,N_1415,N_1425);
or U1447 (N_1447,N_1429,N_1409);
nor U1448 (N_1448,N_1402,N_1439);
nor U1449 (N_1449,N_1391,N_1403);
or U1450 (N_1450,N_1404,N_1417);
nor U1451 (N_1451,N_1416,N_1423);
xnor U1452 (N_1452,N_1411,N_1436);
xnor U1453 (N_1453,N_1389,N_1395);
nor U1454 (N_1454,N_1398,N_1426);
nand U1455 (N_1455,N_1399,N_1397);
nand U1456 (N_1456,N_1435,N_1414);
or U1457 (N_1457,N_1428,N_1406);
xor U1458 (N_1458,N_1386,N_1420);
and U1459 (N_1459,N_1408,N_1432);
nor U1460 (N_1460,N_1405,N_1418);
nor U1461 (N_1461,N_1434,N_1387);
nor U1462 (N_1462,N_1383,N_1385);
xnor U1463 (N_1463,N_1380,N_1430);
nand U1464 (N_1464,N_1431,N_1384);
or U1465 (N_1465,N_1410,N_1421);
or U1466 (N_1466,N_1438,N_1433);
or U1467 (N_1467,N_1422,N_1413);
xor U1468 (N_1468,N_1412,N_1388);
nand U1469 (N_1469,N_1394,N_1419);
and U1470 (N_1470,N_1429,N_1425);
xnor U1471 (N_1471,N_1396,N_1409);
nor U1472 (N_1472,N_1400,N_1387);
or U1473 (N_1473,N_1403,N_1387);
xor U1474 (N_1474,N_1414,N_1424);
nand U1475 (N_1475,N_1417,N_1438);
and U1476 (N_1476,N_1389,N_1394);
or U1477 (N_1477,N_1428,N_1381);
or U1478 (N_1478,N_1401,N_1398);
or U1479 (N_1479,N_1387,N_1398);
xnor U1480 (N_1480,N_1389,N_1390);
or U1481 (N_1481,N_1432,N_1438);
nand U1482 (N_1482,N_1422,N_1426);
xor U1483 (N_1483,N_1418,N_1412);
nor U1484 (N_1484,N_1395,N_1436);
xor U1485 (N_1485,N_1381,N_1429);
or U1486 (N_1486,N_1418,N_1429);
or U1487 (N_1487,N_1434,N_1409);
nor U1488 (N_1488,N_1438,N_1414);
nand U1489 (N_1489,N_1387,N_1402);
or U1490 (N_1490,N_1432,N_1382);
and U1491 (N_1491,N_1395,N_1417);
xnor U1492 (N_1492,N_1438,N_1439);
and U1493 (N_1493,N_1410,N_1403);
nor U1494 (N_1494,N_1381,N_1406);
xnor U1495 (N_1495,N_1432,N_1395);
xor U1496 (N_1496,N_1414,N_1405);
nor U1497 (N_1497,N_1419,N_1381);
and U1498 (N_1498,N_1387,N_1408);
and U1499 (N_1499,N_1395,N_1403);
xnor U1500 (N_1500,N_1441,N_1484);
nand U1501 (N_1501,N_1462,N_1454);
and U1502 (N_1502,N_1494,N_1450);
nor U1503 (N_1503,N_1474,N_1486);
and U1504 (N_1504,N_1469,N_1472);
and U1505 (N_1505,N_1452,N_1455);
nand U1506 (N_1506,N_1467,N_1476);
nor U1507 (N_1507,N_1461,N_1447);
or U1508 (N_1508,N_1475,N_1495);
nor U1509 (N_1509,N_1471,N_1470);
nor U1510 (N_1510,N_1464,N_1451);
xor U1511 (N_1511,N_1492,N_1457);
nor U1512 (N_1512,N_1440,N_1478);
and U1513 (N_1513,N_1496,N_1444);
nand U1514 (N_1514,N_1458,N_1488);
nand U1515 (N_1515,N_1466,N_1489);
xor U1516 (N_1516,N_1459,N_1493);
or U1517 (N_1517,N_1443,N_1460);
or U1518 (N_1518,N_1473,N_1465);
nand U1519 (N_1519,N_1487,N_1499);
xnor U1520 (N_1520,N_1482,N_1480);
or U1521 (N_1521,N_1456,N_1477);
xor U1522 (N_1522,N_1468,N_1481);
xor U1523 (N_1523,N_1446,N_1449);
xnor U1524 (N_1524,N_1497,N_1498);
nand U1525 (N_1525,N_1490,N_1442);
nand U1526 (N_1526,N_1491,N_1479);
and U1527 (N_1527,N_1445,N_1453);
nor U1528 (N_1528,N_1485,N_1483);
and U1529 (N_1529,N_1448,N_1463);
and U1530 (N_1530,N_1444,N_1492);
or U1531 (N_1531,N_1469,N_1480);
and U1532 (N_1532,N_1495,N_1491);
nor U1533 (N_1533,N_1456,N_1492);
nand U1534 (N_1534,N_1465,N_1451);
and U1535 (N_1535,N_1491,N_1468);
nor U1536 (N_1536,N_1449,N_1445);
nor U1537 (N_1537,N_1496,N_1468);
nand U1538 (N_1538,N_1462,N_1460);
or U1539 (N_1539,N_1481,N_1483);
xor U1540 (N_1540,N_1463,N_1475);
nor U1541 (N_1541,N_1488,N_1487);
or U1542 (N_1542,N_1470,N_1452);
xnor U1543 (N_1543,N_1457,N_1494);
and U1544 (N_1544,N_1473,N_1461);
xnor U1545 (N_1545,N_1467,N_1453);
xnor U1546 (N_1546,N_1443,N_1446);
xor U1547 (N_1547,N_1451,N_1489);
nor U1548 (N_1548,N_1490,N_1451);
and U1549 (N_1549,N_1454,N_1456);
or U1550 (N_1550,N_1492,N_1482);
and U1551 (N_1551,N_1465,N_1498);
nand U1552 (N_1552,N_1461,N_1446);
and U1553 (N_1553,N_1484,N_1472);
or U1554 (N_1554,N_1483,N_1498);
nor U1555 (N_1555,N_1440,N_1471);
nand U1556 (N_1556,N_1444,N_1459);
or U1557 (N_1557,N_1481,N_1450);
nand U1558 (N_1558,N_1455,N_1443);
nor U1559 (N_1559,N_1479,N_1457);
and U1560 (N_1560,N_1541,N_1557);
or U1561 (N_1561,N_1501,N_1536);
or U1562 (N_1562,N_1531,N_1513);
or U1563 (N_1563,N_1545,N_1534);
nor U1564 (N_1564,N_1511,N_1510);
or U1565 (N_1565,N_1542,N_1519);
and U1566 (N_1566,N_1532,N_1556);
nand U1567 (N_1567,N_1530,N_1520);
and U1568 (N_1568,N_1506,N_1554);
and U1569 (N_1569,N_1523,N_1514);
nand U1570 (N_1570,N_1555,N_1508);
xor U1571 (N_1571,N_1559,N_1549);
or U1572 (N_1572,N_1504,N_1535);
nor U1573 (N_1573,N_1518,N_1507);
nor U1574 (N_1574,N_1552,N_1502);
or U1575 (N_1575,N_1524,N_1543);
and U1576 (N_1576,N_1528,N_1503);
xnor U1577 (N_1577,N_1550,N_1529);
nand U1578 (N_1578,N_1537,N_1512);
or U1579 (N_1579,N_1540,N_1526);
xor U1580 (N_1580,N_1525,N_1547);
xnor U1581 (N_1581,N_1515,N_1516);
xor U1582 (N_1582,N_1553,N_1521);
nor U1583 (N_1583,N_1522,N_1505);
xnor U1584 (N_1584,N_1551,N_1544);
nor U1585 (N_1585,N_1517,N_1533);
nand U1586 (N_1586,N_1509,N_1539);
xnor U1587 (N_1587,N_1527,N_1500);
nor U1588 (N_1588,N_1558,N_1548);
nor U1589 (N_1589,N_1538,N_1546);
nor U1590 (N_1590,N_1538,N_1514);
and U1591 (N_1591,N_1540,N_1501);
nand U1592 (N_1592,N_1521,N_1552);
xor U1593 (N_1593,N_1546,N_1514);
nor U1594 (N_1594,N_1532,N_1508);
and U1595 (N_1595,N_1556,N_1514);
and U1596 (N_1596,N_1505,N_1501);
and U1597 (N_1597,N_1509,N_1554);
and U1598 (N_1598,N_1553,N_1519);
or U1599 (N_1599,N_1511,N_1559);
xor U1600 (N_1600,N_1543,N_1549);
nor U1601 (N_1601,N_1500,N_1509);
xnor U1602 (N_1602,N_1531,N_1517);
and U1603 (N_1603,N_1513,N_1507);
or U1604 (N_1604,N_1553,N_1508);
xor U1605 (N_1605,N_1557,N_1546);
xnor U1606 (N_1606,N_1500,N_1526);
or U1607 (N_1607,N_1538,N_1520);
xor U1608 (N_1608,N_1535,N_1500);
xor U1609 (N_1609,N_1503,N_1536);
nor U1610 (N_1610,N_1527,N_1504);
xor U1611 (N_1611,N_1500,N_1552);
or U1612 (N_1612,N_1518,N_1555);
nand U1613 (N_1613,N_1519,N_1506);
xnor U1614 (N_1614,N_1501,N_1500);
nand U1615 (N_1615,N_1517,N_1519);
xor U1616 (N_1616,N_1557,N_1527);
nor U1617 (N_1617,N_1504,N_1516);
nor U1618 (N_1618,N_1533,N_1515);
nor U1619 (N_1619,N_1557,N_1522);
and U1620 (N_1620,N_1602,N_1615);
nor U1621 (N_1621,N_1606,N_1582);
nand U1622 (N_1622,N_1591,N_1596);
xnor U1623 (N_1623,N_1610,N_1589);
or U1624 (N_1624,N_1609,N_1561);
and U1625 (N_1625,N_1587,N_1616);
nand U1626 (N_1626,N_1601,N_1612);
xor U1627 (N_1627,N_1571,N_1619);
and U1628 (N_1628,N_1581,N_1614);
xnor U1629 (N_1629,N_1578,N_1575);
and U1630 (N_1630,N_1585,N_1618);
nand U1631 (N_1631,N_1611,N_1573);
nor U1632 (N_1632,N_1608,N_1617);
nor U1633 (N_1633,N_1605,N_1592);
xor U1634 (N_1634,N_1590,N_1588);
or U1635 (N_1635,N_1577,N_1570);
or U1636 (N_1636,N_1567,N_1580);
nor U1637 (N_1637,N_1594,N_1584);
or U1638 (N_1638,N_1597,N_1564);
nand U1639 (N_1639,N_1599,N_1579);
and U1640 (N_1640,N_1569,N_1613);
nand U1641 (N_1641,N_1560,N_1563);
nand U1642 (N_1642,N_1568,N_1583);
or U1643 (N_1643,N_1593,N_1566);
nand U1644 (N_1644,N_1607,N_1562);
nand U1645 (N_1645,N_1572,N_1565);
nand U1646 (N_1646,N_1598,N_1604);
and U1647 (N_1647,N_1595,N_1574);
or U1648 (N_1648,N_1576,N_1603);
nand U1649 (N_1649,N_1586,N_1600);
nor U1650 (N_1650,N_1562,N_1612);
nor U1651 (N_1651,N_1569,N_1602);
and U1652 (N_1652,N_1617,N_1577);
nand U1653 (N_1653,N_1619,N_1578);
nor U1654 (N_1654,N_1617,N_1585);
nand U1655 (N_1655,N_1591,N_1606);
xor U1656 (N_1656,N_1570,N_1597);
and U1657 (N_1657,N_1578,N_1618);
xor U1658 (N_1658,N_1598,N_1574);
and U1659 (N_1659,N_1577,N_1573);
xor U1660 (N_1660,N_1584,N_1589);
xnor U1661 (N_1661,N_1566,N_1586);
nor U1662 (N_1662,N_1599,N_1595);
and U1663 (N_1663,N_1616,N_1584);
nand U1664 (N_1664,N_1595,N_1565);
nor U1665 (N_1665,N_1601,N_1613);
or U1666 (N_1666,N_1582,N_1590);
or U1667 (N_1667,N_1580,N_1564);
xor U1668 (N_1668,N_1581,N_1562);
or U1669 (N_1669,N_1575,N_1570);
and U1670 (N_1670,N_1560,N_1604);
nor U1671 (N_1671,N_1613,N_1577);
or U1672 (N_1672,N_1618,N_1592);
nor U1673 (N_1673,N_1617,N_1591);
and U1674 (N_1674,N_1588,N_1572);
or U1675 (N_1675,N_1581,N_1563);
nand U1676 (N_1676,N_1589,N_1565);
and U1677 (N_1677,N_1610,N_1588);
and U1678 (N_1678,N_1563,N_1567);
nand U1679 (N_1679,N_1575,N_1560);
xnor U1680 (N_1680,N_1654,N_1640);
nand U1681 (N_1681,N_1674,N_1638);
and U1682 (N_1682,N_1630,N_1668);
xnor U1683 (N_1683,N_1634,N_1670);
nor U1684 (N_1684,N_1658,N_1672);
nor U1685 (N_1685,N_1655,N_1677);
and U1686 (N_1686,N_1659,N_1664);
and U1687 (N_1687,N_1628,N_1660);
nor U1688 (N_1688,N_1663,N_1673);
nand U1689 (N_1689,N_1647,N_1632);
nor U1690 (N_1690,N_1637,N_1633);
xor U1691 (N_1691,N_1629,N_1649);
nor U1692 (N_1692,N_1621,N_1651);
xnor U1693 (N_1693,N_1624,N_1625);
xor U1694 (N_1694,N_1645,N_1661);
and U1695 (N_1695,N_1639,N_1669);
nor U1696 (N_1696,N_1626,N_1641);
xor U1697 (N_1697,N_1662,N_1666);
nor U1698 (N_1698,N_1665,N_1657);
xnor U1699 (N_1699,N_1653,N_1642);
or U1700 (N_1700,N_1644,N_1622);
xnor U1701 (N_1701,N_1643,N_1675);
or U1702 (N_1702,N_1636,N_1667);
nor U1703 (N_1703,N_1676,N_1635);
nor U1704 (N_1704,N_1623,N_1648);
nor U1705 (N_1705,N_1627,N_1646);
nor U1706 (N_1706,N_1679,N_1650);
xor U1707 (N_1707,N_1631,N_1656);
nand U1708 (N_1708,N_1620,N_1652);
nand U1709 (N_1709,N_1671,N_1678);
and U1710 (N_1710,N_1676,N_1645);
nor U1711 (N_1711,N_1639,N_1633);
and U1712 (N_1712,N_1657,N_1644);
nor U1713 (N_1713,N_1678,N_1645);
xnor U1714 (N_1714,N_1644,N_1632);
or U1715 (N_1715,N_1632,N_1673);
nand U1716 (N_1716,N_1633,N_1667);
and U1717 (N_1717,N_1660,N_1646);
or U1718 (N_1718,N_1667,N_1675);
or U1719 (N_1719,N_1659,N_1675);
xnor U1720 (N_1720,N_1634,N_1668);
xor U1721 (N_1721,N_1653,N_1649);
nor U1722 (N_1722,N_1665,N_1674);
nand U1723 (N_1723,N_1664,N_1670);
nand U1724 (N_1724,N_1653,N_1635);
or U1725 (N_1725,N_1635,N_1632);
or U1726 (N_1726,N_1621,N_1652);
nand U1727 (N_1727,N_1679,N_1627);
or U1728 (N_1728,N_1630,N_1626);
nor U1729 (N_1729,N_1621,N_1655);
and U1730 (N_1730,N_1656,N_1671);
and U1731 (N_1731,N_1627,N_1635);
nand U1732 (N_1732,N_1654,N_1639);
and U1733 (N_1733,N_1623,N_1630);
or U1734 (N_1734,N_1631,N_1638);
and U1735 (N_1735,N_1641,N_1639);
or U1736 (N_1736,N_1631,N_1624);
nand U1737 (N_1737,N_1669,N_1657);
and U1738 (N_1738,N_1678,N_1646);
nor U1739 (N_1739,N_1675,N_1638);
nor U1740 (N_1740,N_1717,N_1715);
nor U1741 (N_1741,N_1686,N_1681);
nor U1742 (N_1742,N_1723,N_1704);
and U1743 (N_1743,N_1727,N_1697);
xnor U1744 (N_1744,N_1734,N_1688);
nand U1745 (N_1745,N_1730,N_1694);
xor U1746 (N_1746,N_1703,N_1707);
xnor U1747 (N_1747,N_1689,N_1693);
nor U1748 (N_1748,N_1708,N_1696);
and U1749 (N_1749,N_1682,N_1729);
nor U1750 (N_1750,N_1712,N_1736);
xnor U1751 (N_1751,N_1709,N_1724);
and U1752 (N_1752,N_1721,N_1699);
or U1753 (N_1753,N_1713,N_1711);
or U1754 (N_1754,N_1725,N_1722);
nor U1755 (N_1755,N_1692,N_1684);
or U1756 (N_1756,N_1698,N_1714);
nand U1757 (N_1757,N_1690,N_1718);
and U1758 (N_1758,N_1687,N_1732);
xor U1759 (N_1759,N_1726,N_1738);
nand U1760 (N_1760,N_1737,N_1710);
nor U1761 (N_1761,N_1735,N_1706);
or U1762 (N_1762,N_1719,N_1728);
or U1763 (N_1763,N_1695,N_1720);
or U1764 (N_1764,N_1702,N_1733);
nand U1765 (N_1765,N_1731,N_1685);
nor U1766 (N_1766,N_1705,N_1691);
or U1767 (N_1767,N_1739,N_1700);
and U1768 (N_1768,N_1680,N_1716);
xnor U1769 (N_1769,N_1701,N_1683);
nor U1770 (N_1770,N_1720,N_1685);
xnor U1771 (N_1771,N_1698,N_1735);
or U1772 (N_1772,N_1712,N_1717);
and U1773 (N_1773,N_1697,N_1738);
nand U1774 (N_1774,N_1680,N_1687);
xor U1775 (N_1775,N_1734,N_1730);
and U1776 (N_1776,N_1724,N_1733);
or U1777 (N_1777,N_1716,N_1700);
xor U1778 (N_1778,N_1704,N_1729);
nand U1779 (N_1779,N_1691,N_1735);
or U1780 (N_1780,N_1693,N_1736);
nor U1781 (N_1781,N_1727,N_1719);
xnor U1782 (N_1782,N_1722,N_1706);
and U1783 (N_1783,N_1719,N_1683);
xnor U1784 (N_1784,N_1686,N_1702);
or U1785 (N_1785,N_1705,N_1693);
xor U1786 (N_1786,N_1734,N_1695);
or U1787 (N_1787,N_1732,N_1725);
nand U1788 (N_1788,N_1736,N_1705);
and U1789 (N_1789,N_1716,N_1711);
and U1790 (N_1790,N_1697,N_1737);
and U1791 (N_1791,N_1727,N_1706);
nor U1792 (N_1792,N_1727,N_1684);
or U1793 (N_1793,N_1729,N_1693);
xor U1794 (N_1794,N_1685,N_1737);
xnor U1795 (N_1795,N_1726,N_1683);
nand U1796 (N_1796,N_1683,N_1685);
nand U1797 (N_1797,N_1703,N_1708);
and U1798 (N_1798,N_1739,N_1697);
nor U1799 (N_1799,N_1680,N_1695);
and U1800 (N_1800,N_1773,N_1793);
nand U1801 (N_1801,N_1760,N_1754);
nor U1802 (N_1802,N_1788,N_1787);
or U1803 (N_1803,N_1778,N_1797);
or U1804 (N_1804,N_1744,N_1782);
or U1805 (N_1805,N_1765,N_1785);
or U1806 (N_1806,N_1759,N_1769);
nand U1807 (N_1807,N_1770,N_1786);
xnor U1808 (N_1808,N_1757,N_1761);
xnor U1809 (N_1809,N_1767,N_1751);
xor U1810 (N_1810,N_1750,N_1749);
xor U1811 (N_1811,N_1776,N_1772);
xnor U1812 (N_1812,N_1752,N_1755);
or U1813 (N_1813,N_1764,N_1763);
nor U1814 (N_1814,N_1784,N_1774);
nor U1815 (N_1815,N_1758,N_1748);
or U1816 (N_1816,N_1771,N_1796);
xor U1817 (N_1817,N_1741,N_1795);
and U1818 (N_1818,N_1766,N_1742);
nand U1819 (N_1819,N_1791,N_1779);
and U1820 (N_1820,N_1756,N_1762);
and U1821 (N_1821,N_1780,N_1740);
xor U1822 (N_1822,N_1781,N_1743);
nor U1823 (N_1823,N_1753,N_1775);
and U1824 (N_1824,N_1794,N_1746);
or U1825 (N_1825,N_1745,N_1777);
nor U1826 (N_1826,N_1792,N_1789);
xor U1827 (N_1827,N_1799,N_1747);
and U1828 (N_1828,N_1798,N_1783);
and U1829 (N_1829,N_1790,N_1768);
or U1830 (N_1830,N_1754,N_1762);
nor U1831 (N_1831,N_1778,N_1742);
nand U1832 (N_1832,N_1783,N_1741);
or U1833 (N_1833,N_1741,N_1755);
nor U1834 (N_1834,N_1741,N_1765);
xor U1835 (N_1835,N_1768,N_1785);
nand U1836 (N_1836,N_1794,N_1792);
xor U1837 (N_1837,N_1747,N_1785);
and U1838 (N_1838,N_1747,N_1751);
and U1839 (N_1839,N_1758,N_1788);
xor U1840 (N_1840,N_1753,N_1781);
or U1841 (N_1841,N_1783,N_1772);
nor U1842 (N_1842,N_1772,N_1771);
or U1843 (N_1843,N_1747,N_1760);
nor U1844 (N_1844,N_1770,N_1757);
or U1845 (N_1845,N_1741,N_1780);
or U1846 (N_1846,N_1782,N_1763);
nand U1847 (N_1847,N_1781,N_1750);
xnor U1848 (N_1848,N_1749,N_1740);
xnor U1849 (N_1849,N_1763,N_1794);
xor U1850 (N_1850,N_1797,N_1773);
nand U1851 (N_1851,N_1769,N_1779);
or U1852 (N_1852,N_1784,N_1791);
or U1853 (N_1853,N_1791,N_1787);
and U1854 (N_1854,N_1743,N_1753);
nor U1855 (N_1855,N_1764,N_1771);
or U1856 (N_1856,N_1797,N_1794);
nor U1857 (N_1857,N_1789,N_1795);
nor U1858 (N_1858,N_1798,N_1760);
and U1859 (N_1859,N_1745,N_1766);
nor U1860 (N_1860,N_1855,N_1821);
or U1861 (N_1861,N_1856,N_1854);
or U1862 (N_1862,N_1808,N_1830);
or U1863 (N_1863,N_1846,N_1828);
nand U1864 (N_1864,N_1805,N_1845);
xor U1865 (N_1865,N_1801,N_1833);
nand U1866 (N_1866,N_1822,N_1852);
nand U1867 (N_1867,N_1818,N_1827);
nor U1868 (N_1868,N_1817,N_1844);
nand U1869 (N_1869,N_1848,N_1825);
nand U1870 (N_1870,N_1816,N_1813);
or U1871 (N_1871,N_1832,N_1849);
xnor U1872 (N_1872,N_1843,N_1851);
or U1873 (N_1873,N_1853,N_1847);
or U1874 (N_1874,N_1858,N_1814);
or U1875 (N_1875,N_1809,N_1857);
xor U1876 (N_1876,N_1819,N_1804);
nand U1877 (N_1877,N_1826,N_1842);
xnor U1878 (N_1878,N_1831,N_1803);
nor U1879 (N_1879,N_1823,N_1807);
nor U1880 (N_1880,N_1850,N_1810);
nor U1881 (N_1881,N_1841,N_1838);
and U1882 (N_1882,N_1839,N_1829);
nand U1883 (N_1883,N_1820,N_1812);
nor U1884 (N_1884,N_1859,N_1837);
and U1885 (N_1885,N_1840,N_1815);
xnor U1886 (N_1886,N_1811,N_1834);
nor U1887 (N_1887,N_1835,N_1802);
nor U1888 (N_1888,N_1806,N_1800);
nand U1889 (N_1889,N_1836,N_1824);
xnor U1890 (N_1890,N_1841,N_1835);
nand U1891 (N_1891,N_1840,N_1825);
or U1892 (N_1892,N_1844,N_1837);
xor U1893 (N_1893,N_1859,N_1842);
nor U1894 (N_1894,N_1839,N_1802);
or U1895 (N_1895,N_1841,N_1847);
and U1896 (N_1896,N_1829,N_1846);
xor U1897 (N_1897,N_1827,N_1855);
nor U1898 (N_1898,N_1834,N_1809);
and U1899 (N_1899,N_1808,N_1813);
xor U1900 (N_1900,N_1854,N_1812);
nand U1901 (N_1901,N_1800,N_1805);
xor U1902 (N_1902,N_1846,N_1808);
nand U1903 (N_1903,N_1846,N_1820);
or U1904 (N_1904,N_1813,N_1811);
and U1905 (N_1905,N_1842,N_1828);
nor U1906 (N_1906,N_1804,N_1832);
or U1907 (N_1907,N_1842,N_1817);
and U1908 (N_1908,N_1846,N_1815);
and U1909 (N_1909,N_1839,N_1824);
nand U1910 (N_1910,N_1814,N_1805);
xnor U1911 (N_1911,N_1830,N_1812);
nor U1912 (N_1912,N_1837,N_1857);
xor U1913 (N_1913,N_1851,N_1806);
nand U1914 (N_1914,N_1839,N_1807);
xnor U1915 (N_1915,N_1839,N_1852);
nand U1916 (N_1916,N_1843,N_1846);
or U1917 (N_1917,N_1804,N_1812);
and U1918 (N_1918,N_1853,N_1821);
nand U1919 (N_1919,N_1825,N_1854);
nand U1920 (N_1920,N_1870,N_1909);
nand U1921 (N_1921,N_1911,N_1918);
or U1922 (N_1922,N_1862,N_1880);
or U1923 (N_1923,N_1916,N_1919);
xor U1924 (N_1924,N_1913,N_1882);
and U1925 (N_1925,N_1871,N_1881);
xor U1926 (N_1926,N_1887,N_1899);
and U1927 (N_1927,N_1885,N_1905);
or U1928 (N_1928,N_1901,N_1861);
and U1929 (N_1929,N_1878,N_1886);
and U1930 (N_1930,N_1906,N_1900);
nor U1931 (N_1931,N_1891,N_1902);
nand U1932 (N_1932,N_1904,N_1892);
nor U1933 (N_1933,N_1917,N_1884);
nand U1934 (N_1934,N_1893,N_1908);
nand U1935 (N_1935,N_1866,N_1898);
xnor U1936 (N_1936,N_1894,N_1863);
and U1937 (N_1937,N_1889,N_1890);
nand U1938 (N_1938,N_1869,N_1895);
and U1939 (N_1939,N_1879,N_1875);
xnor U1940 (N_1940,N_1873,N_1896);
and U1941 (N_1941,N_1874,N_1865);
nor U1942 (N_1942,N_1910,N_1914);
nor U1943 (N_1943,N_1864,N_1888);
and U1944 (N_1944,N_1907,N_1912);
nand U1945 (N_1945,N_1877,N_1860);
and U1946 (N_1946,N_1897,N_1883);
xor U1947 (N_1947,N_1903,N_1872);
or U1948 (N_1948,N_1915,N_1867);
xnor U1949 (N_1949,N_1868,N_1876);
or U1950 (N_1950,N_1868,N_1896);
xnor U1951 (N_1951,N_1918,N_1865);
or U1952 (N_1952,N_1870,N_1866);
and U1953 (N_1953,N_1888,N_1876);
nand U1954 (N_1954,N_1903,N_1911);
and U1955 (N_1955,N_1879,N_1915);
nand U1956 (N_1956,N_1872,N_1910);
or U1957 (N_1957,N_1864,N_1860);
xor U1958 (N_1958,N_1867,N_1906);
and U1959 (N_1959,N_1871,N_1865);
xnor U1960 (N_1960,N_1891,N_1871);
or U1961 (N_1961,N_1863,N_1862);
or U1962 (N_1962,N_1876,N_1903);
nor U1963 (N_1963,N_1881,N_1890);
and U1964 (N_1964,N_1881,N_1893);
or U1965 (N_1965,N_1908,N_1913);
nand U1966 (N_1966,N_1908,N_1918);
nor U1967 (N_1967,N_1917,N_1862);
xnor U1968 (N_1968,N_1885,N_1906);
nand U1969 (N_1969,N_1861,N_1894);
nor U1970 (N_1970,N_1915,N_1896);
and U1971 (N_1971,N_1890,N_1914);
xor U1972 (N_1972,N_1873,N_1898);
nor U1973 (N_1973,N_1861,N_1886);
nand U1974 (N_1974,N_1907,N_1873);
nand U1975 (N_1975,N_1863,N_1919);
xor U1976 (N_1976,N_1870,N_1894);
nor U1977 (N_1977,N_1906,N_1886);
xnor U1978 (N_1978,N_1894,N_1868);
and U1979 (N_1979,N_1901,N_1885);
xor U1980 (N_1980,N_1965,N_1952);
nand U1981 (N_1981,N_1926,N_1975);
nor U1982 (N_1982,N_1937,N_1961);
or U1983 (N_1983,N_1971,N_1936);
or U1984 (N_1984,N_1966,N_1948);
nand U1985 (N_1985,N_1923,N_1931);
xor U1986 (N_1986,N_1968,N_1922);
and U1987 (N_1987,N_1940,N_1943);
nand U1988 (N_1988,N_1963,N_1945);
xnor U1989 (N_1989,N_1938,N_1974);
or U1990 (N_1990,N_1924,N_1978);
nor U1991 (N_1991,N_1939,N_1928);
or U1992 (N_1992,N_1935,N_1934);
and U1993 (N_1993,N_1941,N_1953);
nand U1994 (N_1994,N_1958,N_1954);
nand U1995 (N_1995,N_1960,N_1969);
xnor U1996 (N_1996,N_1951,N_1970);
xor U1997 (N_1997,N_1921,N_1955);
xnor U1998 (N_1998,N_1944,N_1956);
or U1999 (N_1999,N_1950,N_1959);
nand U2000 (N_2000,N_1972,N_1962);
and U2001 (N_2001,N_1964,N_1920);
and U2002 (N_2002,N_1929,N_1930);
xnor U2003 (N_2003,N_1946,N_1947);
nor U2004 (N_2004,N_1933,N_1942);
xnor U2005 (N_2005,N_1949,N_1957);
xnor U2006 (N_2006,N_1976,N_1973);
and U2007 (N_2007,N_1927,N_1979);
or U2008 (N_2008,N_1977,N_1967);
nand U2009 (N_2009,N_1925,N_1932);
xor U2010 (N_2010,N_1939,N_1964);
nand U2011 (N_2011,N_1972,N_1921);
xnor U2012 (N_2012,N_1953,N_1965);
nor U2013 (N_2013,N_1951,N_1956);
xnor U2014 (N_2014,N_1950,N_1951);
xor U2015 (N_2015,N_1931,N_1947);
nor U2016 (N_2016,N_1957,N_1971);
or U2017 (N_2017,N_1966,N_1945);
or U2018 (N_2018,N_1928,N_1954);
nor U2019 (N_2019,N_1958,N_1963);
xnor U2020 (N_2020,N_1933,N_1978);
nand U2021 (N_2021,N_1929,N_1945);
nand U2022 (N_2022,N_1940,N_1959);
or U2023 (N_2023,N_1963,N_1979);
or U2024 (N_2024,N_1947,N_1942);
and U2025 (N_2025,N_1942,N_1930);
xnor U2026 (N_2026,N_1972,N_1922);
nor U2027 (N_2027,N_1947,N_1925);
or U2028 (N_2028,N_1944,N_1962);
nor U2029 (N_2029,N_1973,N_1934);
xor U2030 (N_2030,N_1940,N_1956);
nand U2031 (N_2031,N_1937,N_1975);
nand U2032 (N_2032,N_1924,N_1960);
or U2033 (N_2033,N_1935,N_1951);
xnor U2034 (N_2034,N_1932,N_1923);
and U2035 (N_2035,N_1958,N_1978);
and U2036 (N_2036,N_1979,N_1977);
xor U2037 (N_2037,N_1945,N_1972);
nor U2038 (N_2038,N_1954,N_1940);
nor U2039 (N_2039,N_1927,N_1926);
xor U2040 (N_2040,N_1984,N_2018);
nand U2041 (N_2041,N_2028,N_2006);
or U2042 (N_2042,N_2031,N_1983);
xnor U2043 (N_2043,N_2009,N_2012);
and U2044 (N_2044,N_1990,N_2026);
nand U2045 (N_2045,N_2027,N_1985);
nor U2046 (N_2046,N_1982,N_2017);
or U2047 (N_2047,N_2034,N_2035);
xnor U2048 (N_2048,N_2030,N_1980);
or U2049 (N_2049,N_1991,N_1987);
nor U2050 (N_2050,N_2038,N_2024);
or U2051 (N_2051,N_2013,N_2001);
nor U2052 (N_2052,N_1981,N_1992);
nor U2053 (N_2053,N_1997,N_1996);
xor U2054 (N_2054,N_2002,N_2020);
xor U2055 (N_2055,N_2036,N_1995);
nand U2056 (N_2056,N_2008,N_2016);
or U2057 (N_2057,N_1998,N_2011);
and U2058 (N_2058,N_1993,N_1988);
and U2059 (N_2059,N_2014,N_2007);
xnor U2060 (N_2060,N_2005,N_2022);
and U2061 (N_2061,N_2000,N_2023);
and U2062 (N_2062,N_2019,N_1999);
xnor U2063 (N_2063,N_1989,N_2033);
nor U2064 (N_2064,N_2004,N_2039);
nand U2065 (N_2065,N_2025,N_2010);
nand U2066 (N_2066,N_2032,N_2029);
xnor U2067 (N_2067,N_2037,N_1994);
or U2068 (N_2068,N_2021,N_1986);
or U2069 (N_2069,N_2015,N_2003);
or U2070 (N_2070,N_2007,N_2010);
nand U2071 (N_2071,N_1996,N_1983);
nand U2072 (N_2072,N_2038,N_2000);
nor U2073 (N_2073,N_2023,N_2008);
nand U2074 (N_2074,N_1990,N_2011);
and U2075 (N_2075,N_2038,N_2020);
xor U2076 (N_2076,N_2034,N_2039);
nand U2077 (N_2077,N_1991,N_2034);
nand U2078 (N_2078,N_2001,N_2017);
xnor U2079 (N_2079,N_2029,N_1996);
xor U2080 (N_2080,N_1987,N_2037);
xnor U2081 (N_2081,N_2006,N_1997);
xor U2082 (N_2082,N_2007,N_2029);
nor U2083 (N_2083,N_2030,N_2029);
nand U2084 (N_2084,N_2036,N_2006);
and U2085 (N_2085,N_2002,N_1995);
nor U2086 (N_2086,N_1987,N_2039);
nand U2087 (N_2087,N_1989,N_2020);
xnor U2088 (N_2088,N_2038,N_2031);
nor U2089 (N_2089,N_1980,N_2018);
xor U2090 (N_2090,N_1994,N_1982);
nand U2091 (N_2091,N_2005,N_2032);
and U2092 (N_2092,N_1993,N_2034);
nor U2093 (N_2093,N_2035,N_1995);
and U2094 (N_2094,N_2031,N_1982);
nand U2095 (N_2095,N_2036,N_2023);
nand U2096 (N_2096,N_2037,N_2027);
xnor U2097 (N_2097,N_2000,N_2026);
and U2098 (N_2098,N_2037,N_1990);
and U2099 (N_2099,N_2010,N_2004);
nand U2100 (N_2100,N_2049,N_2089);
xor U2101 (N_2101,N_2093,N_2045);
nor U2102 (N_2102,N_2065,N_2085);
nand U2103 (N_2103,N_2052,N_2078);
or U2104 (N_2104,N_2043,N_2060);
and U2105 (N_2105,N_2068,N_2069);
or U2106 (N_2106,N_2067,N_2071);
and U2107 (N_2107,N_2054,N_2070);
nor U2108 (N_2108,N_2084,N_2048);
xor U2109 (N_2109,N_2050,N_2046);
nand U2110 (N_2110,N_2096,N_2083);
or U2111 (N_2111,N_2075,N_2081);
xnor U2112 (N_2112,N_2074,N_2044);
nor U2113 (N_2113,N_2056,N_2090);
nor U2114 (N_2114,N_2073,N_2082);
or U2115 (N_2115,N_2076,N_2047);
or U2116 (N_2116,N_2057,N_2055);
nand U2117 (N_2117,N_2053,N_2040);
or U2118 (N_2118,N_2092,N_2051);
or U2119 (N_2119,N_2079,N_2097);
and U2120 (N_2120,N_2066,N_2086);
xor U2121 (N_2121,N_2088,N_2062);
or U2122 (N_2122,N_2091,N_2095);
xor U2123 (N_2123,N_2041,N_2064);
nor U2124 (N_2124,N_2094,N_2077);
nand U2125 (N_2125,N_2087,N_2098);
and U2126 (N_2126,N_2080,N_2063);
xnor U2127 (N_2127,N_2058,N_2042);
xnor U2128 (N_2128,N_2061,N_2059);
and U2129 (N_2129,N_2072,N_2099);
nand U2130 (N_2130,N_2064,N_2044);
xnor U2131 (N_2131,N_2087,N_2056);
nand U2132 (N_2132,N_2044,N_2070);
nand U2133 (N_2133,N_2044,N_2046);
and U2134 (N_2134,N_2088,N_2097);
nor U2135 (N_2135,N_2068,N_2055);
and U2136 (N_2136,N_2072,N_2061);
and U2137 (N_2137,N_2053,N_2073);
nand U2138 (N_2138,N_2093,N_2075);
and U2139 (N_2139,N_2057,N_2086);
nor U2140 (N_2140,N_2064,N_2097);
or U2141 (N_2141,N_2051,N_2083);
or U2142 (N_2142,N_2060,N_2061);
or U2143 (N_2143,N_2071,N_2072);
xor U2144 (N_2144,N_2058,N_2090);
nand U2145 (N_2145,N_2097,N_2068);
or U2146 (N_2146,N_2096,N_2064);
xnor U2147 (N_2147,N_2094,N_2063);
and U2148 (N_2148,N_2062,N_2073);
xnor U2149 (N_2149,N_2063,N_2050);
nor U2150 (N_2150,N_2079,N_2089);
nand U2151 (N_2151,N_2087,N_2059);
xor U2152 (N_2152,N_2074,N_2063);
or U2153 (N_2153,N_2073,N_2040);
nand U2154 (N_2154,N_2095,N_2045);
xor U2155 (N_2155,N_2066,N_2045);
nor U2156 (N_2156,N_2050,N_2052);
and U2157 (N_2157,N_2043,N_2079);
nor U2158 (N_2158,N_2070,N_2089);
or U2159 (N_2159,N_2058,N_2085);
and U2160 (N_2160,N_2126,N_2110);
xnor U2161 (N_2161,N_2115,N_2148);
xnor U2162 (N_2162,N_2155,N_2109);
nand U2163 (N_2163,N_2113,N_2116);
nand U2164 (N_2164,N_2111,N_2128);
nand U2165 (N_2165,N_2102,N_2135);
and U2166 (N_2166,N_2125,N_2127);
or U2167 (N_2167,N_2147,N_2151);
or U2168 (N_2168,N_2156,N_2150);
xnor U2169 (N_2169,N_2149,N_2146);
nand U2170 (N_2170,N_2130,N_2139);
nand U2171 (N_2171,N_2143,N_2142);
and U2172 (N_2172,N_2138,N_2105);
or U2173 (N_2173,N_2103,N_2119);
nor U2174 (N_2174,N_2106,N_2153);
xor U2175 (N_2175,N_2140,N_2122);
nor U2176 (N_2176,N_2157,N_2118);
xnor U2177 (N_2177,N_2108,N_2141);
xnor U2178 (N_2178,N_2104,N_2154);
nand U2179 (N_2179,N_2101,N_2114);
and U2180 (N_2180,N_2132,N_2120);
nand U2181 (N_2181,N_2131,N_2145);
xor U2182 (N_2182,N_2121,N_2159);
or U2183 (N_2183,N_2134,N_2129);
or U2184 (N_2184,N_2112,N_2158);
and U2185 (N_2185,N_2107,N_2124);
or U2186 (N_2186,N_2137,N_2100);
and U2187 (N_2187,N_2136,N_2117);
nand U2188 (N_2188,N_2133,N_2123);
nor U2189 (N_2189,N_2152,N_2144);
or U2190 (N_2190,N_2125,N_2131);
xnor U2191 (N_2191,N_2149,N_2135);
nor U2192 (N_2192,N_2111,N_2150);
nand U2193 (N_2193,N_2143,N_2103);
and U2194 (N_2194,N_2133,N_2155);
xnor U2195 (N_2195,N_2145,N_2141);
and U2196 (N_2196,N_2147,N_2125);
nand U2197 (N_2197,N_2144,N_2135);
or U2198 (N_2198,N_2138,N_2141);
and U2199 (N_2199,N_2115,N_2111);
nand U2200 (N_2200,N_2142,N_2153);
nor U2201 (N_2201,N_2148,N_2105);
and U2202 (N_2202,N_2157,N_2143);
nor U2203 (N_2203,N_2152,N_2106);
xor U2204 (N_2204,N_2103,N_2106);
nor U2205 (N_2205,N_2111,N_2141);
xor U2206 (N_2206,N_2147,N_2109);
nand U2207 (N_2207,N_2154,N_2149);
or U2208 (N_2208,N_2113,N_2133);
and U2209 (N_2209,N_2123,N_2117);
xnor U2210 (N_2210,N_2141,N_2143);
nand U2211 (N_2211,N_2125,N_2156);
and U2212 (N_2212,N_2143,N_2136);
and U2213 (N_2213,N_2132,N_2145);
xnor U2214 (N_2214,N_2141,N_2121);
nor U2215 (N_2215,N_2136,N_2108);
or U2216 (N_2216,N_2116,N_2108);
xnor U2217 (N_2217,N_2105,N_2119);
nand U2218 (N_2218,N_2112,N_2159);
nand U2219 (N_2219,N_2158,N_2116);
or U2220 (N_2220,N_2185,N_2219);
xnor U2221 (N_2221,N_2175,N_2215);
or U2222 (N_2222,N_2188,N_2210);
nand U2223 (N_2223,N_2162,N_2191);
nor U2224 (N_2224,N_2186,N_2170);
nor U2225 (N_2225,N_2184,N_2201);
nand U2226 (N_2226,N_2167,N_2177);
nor U2227 (N_2227,N_2181,N_2197);
nand U2228 (N_2228,N_2174,N_2192);
nand U2229 (N_2229,N_2189,N_2183);
and U2230 (N_2230,N_2213,N_2182);
xnor U2231 (N_2231,N_2205,N_2200);
or U2232 (N_2232,N_2178,N_2216);
or U2233 (N_2233,N_2198,N_2202);
or U2234 (N_2234,N_2165,N_2169);
xor U2235 (N_2235,N_2208,N_2212);
and U2236 (N_2236,N_2204,N_2163);
and U2237 (N_2237,N_2214,N_2160);
and U2238 (N_2238,N_2164,N_2190);
nor U2239 (N_2239,N_2166,N_2218);
xor U2240 (N_2240,N_2194,N_2173);
nand U2241 (N_2241,N_2211,N_2161);
nand U2242 (N_2242,N_2199,N_2180);
xor U2243 (N_2243,N_2179,N_2217);
nor U2244 (N_2244,N_2206,N_2203);
nor U2245 (N_2245,N_2209,N_2168);
and U2246 (N_2246,N_2172,N_2196);
xnor U2247 (N_2247,N_2176,N_2195);
or U2248 (N_2248,N_2171,N_2193);
or U2249 (N_2249,N_2207,N_2187);
xnor U2250 (N_2250,N_2219,N_2163);
xor U2251 (N_2251,N_2168,N_2218);
and U2252 (N_2252,N_2196,N_2219);
and U2253 (N_2253,N_2212,N_2163);
nor U2254 (N_2254,N_2161,N_2203);
or U2255 (N_2255,N_2188,N_2187);
and U2256 (N_2256,N_2193,N_2185);
nand U2257 (N_2257,N_2190,N_2210);
xnor U2258 (N_2258,N_2206,N_2198);
xor U2259 (N_2259,N_2199,N_2189);
and U2260 (N_2260,N_2160,N_2168);
and U2261 (N_2261,N_2196,N_2199);
xor U2262 (N_2262,N_2192,N_2200);
nand U2263 (N_2263,N_2190,N_2191);
and U2264 (N_2264,N_2187,N_2182);
nand U2265 (N_2265,N_2194,N_2163);
or U2266 (N_2266,N_2204,N_2167);
nand U2267 (N_2267,N_2216,N_2188);
xor U2268 (N_2268,N_2204,N_2192);
xor U2269 (N_2269,N_2167,N_2176);
or U2270 (N_2270,N_2161,N_2171);
nand U2271 (N_2271,N_2161,N_2216);
xnor U2272 (N_2272,N_2174,N_2212);
or U2273 (N_2273,N_2199,N_2184);
nor U2274 (N_2274,N_2173,N_2175);
xnor U2275 (N_2275,N_2215,N_2207);
nor U2276 (N_2276,N_2181,N_2196);
xor U2277 (N_2277,N_2169,N_2167);
nor U2278 (N_2278,N_2201,N_2212);
nor U2279 (N_2279,N_2189,N_2204);
or U2280 (N_2280,N_2267,N_2266);
nor U2281 (N_2281,N_2252,N_2276);
or U2282 (N_2282,N_2279,N_2270);
and U2283 (N_2283,N_2222,N_2229);
xnor U2284 (N_2284,N_2237,N_2273);
nor U2285 (N_2285,N_2272,N_2246);
and U2286 (N_2286,N_2238,N_2227);
nor U2287 (N_2287,N_2242,N_2253);
nand U2288 (N_2288,N_2228,N_2230);
and U2289 (N_2289,N_2251,N_2275);
and U2290 (N_2290,N_2225,N_2234);
nor U2291 (N_2291,N_2226,N_2250);
and U2292 (N_2292,N_2271,N_2258);
nor U2293 (N_2293,N_2224,N_2220);
xnor U2294 (N_2294,N_2265,N_2247);
xor U2295 (N_2295,N_2263,N_2248);
and U2296 (N_2296,N_2278,N_2260);
xor U2297 (N_2297,N_2239,N_2255);
nor U2298 (N_2298,N_2259,N_2264);
nand U2299 (N_2299,N_2236,N_2244);
nand U2300 (N_2300,N_2233,N_2268);
nor U2301 (N_2301,N_2241,N_2240);
nand U2302 (N_2302,N_2257,N_2235);
or U2303 (N_2303,N_2277,N_2254);
or U2304 (N_2304,N_2223,N_2221);
nor U2305 (N_2305,N_2232,N_2256);
nor U2306 (N_2306,N_2261,N_2249);
nand U2307 (N_2307,N_2262,N_2231);
and U2308 (N_2308,N_2243,N_2245);
xnor U2309 (N_2309,N_2274,N_2269);
or U2310 (N_2310,N_2272,N_2242);
and U2311 (N_2311,N_2222,N_2227);
xor U2312 (N_2312,N_2266,N_2263);
or U2313 (N_2313,N_2248,N_2254);
nor U2314 (N_2314,N_2238,N_2263);
xor U2315 (N_2315,N_2223,N_2256);
nand U2316 (N_2316,N_2279,N_2225);
xnor U2317 (N_2317,N_2263,N_2240);
nor U2318 (N_2318,N_2220,N_2222);
or U2319 (N_2319,N_2233,N_2237);
and U2320 (N_2320,N_2225,N_2274);
and U2321 (N_2321,N_2278,N_2235);
nand U2322 (N_2322,N_2276,N_2254);
nand U2323 (N_2323,N_2245,N_2267);
and U2324 (N_2324,N_2268,N_2277);
or U2325 (N_2325,N_2237,N_2250);
nor U2326 (N_2326,N_2241,N_2263);
nand U2327 (N_2327,N_2222,N_2225);
or U2328 (N_2328,N_2258,N_2236);
nand U2329 (N_2329,N_2233,N_2247);
xor U2330 (N_2330,N_2256,N_2221);
nand U2331 (N_2331,N_2229,N_2263);
nor U2332 (N_2332,N_2243,N_2234);
nand U2333 (N_2333,N_2247,N_2251);
xnor U2334 (N_2334,N_2237,N_2255);
nor U2335 (N_2335,N_2246,N_2233);
xnor U2336 (N_2336,N_2267,N_2260);
or U2337 (N_2337,N_2261,N_2247);
nand U2338 (N_2338,N_2275,N_2232);
nand U2339 (N_2339,N_2246,N_2227);
xnor U2340 (N_2340,N_2297,N_2284);
and U2341 (N_2341,N_2332,N_2311);
and U2342 (N_2342,N_2290,N_2323);
nand U2343 (N_2343,N_2291,N_2302);
xnor U2344 (N_2344,N_2285,N_2327);
and U2345 (N_2345,N_2280,N_2300);
and U2346 (N_2346,N_2318,N_2314);
xnor U2347 (N_2347,N_2293,N_2321);
xor U2348 (N_2348,N_2304,N_2324);
or U2349 (N_2349,N_2301,N_2295);
nor U2350 (N_2350,N_2289,N_2331);
nor U2351 (N_2351,N_2310,N_2316);
nand U2352 (N_2352,N_2325,N_2305);
xnor U2353 (N_2353,N_2296,N_2328);
nor U2354 (N_2354,N_2281,N_2338);
nand U2355 (N_2355,N_2306,N_2322);
xor U2356 (N_2356,N_2315,N_2303);
or U2357 (N_2357,N_2326,N_2299);
and U2358 (N_2358,N_2329,N_2330);
nor U2359 (N_2359,N_2335,N_2312);
or U2360 (N_2360,N_2319,N_2320);
and U2361 (N_2361,N_2317,N_2334);
or U2362 (N_2362,N_2288,N_2287);
nand U2363 (N_2363,N_2298,N_2283);
and U2364 (N_2364,N_2294,N_2339);
xor U2365 (N_2365,N_2309,N_2307);
xor U2366 (N_2366,N_2282,N_2308);
nand U2367 (N_2367,N_2286,N_2292);
or U2368 (N_2368,N_2313,N_2336);
or U2369 (N_2369,N_2333,N_2337);
and U2370 (N_2370,N_2308,N_2319);
nand U2371 (N_2371,N_2321,N_2299);
or U2372 (N_2372,N_2337,N_2290);
or U2373 (N_2373,N_2334,N_2292);
and U2374 (N_2374,N_2288,N_2293);
or U2375 (N_2375,N_2303,N_2322);
nand U2376 (N_2376,N_2328,N_2316);
xnor U2377 (N_2377,N_2280,N_2291);
nand U2378 (N_2378,N_2332,N_2296);
nor U2379 (N_2379,N_2305,N_2304);
or U2380 (N_2380,N_2334,N_2283);
or U2381 (N_2381,N_2322,N_2285);
xnor U2382 (N_2382,N_2307,N_2310);
and U2383 (N_2383,N_2289,N_2310);
or U2384 (N_2384,N_2288,N_2286);
nor U2385 (N_2385,N_2302,N_2334);
and U2386 (N_2386,N_2305,N_2336);
and U2387 (N_2387,N_2330,N_2325);
and U2388 (N_2388,N_2280,N_2308);
nor U2389 (N_2389,N_2317,N_2304);
nand U2390 (N_2390,N_2298,N_2335);
and U2391 (N_2391,N_2303,N_2302);
and U2392 (N_2392,N_2304,N_2326);
nand U2393 (N_2393,N_2297,N_2315);
and U2394 (N_2394,N_2338,N_2326);
nor U2395 (N_2395,N_2293,N_2323);
nor U2396 (N_2396,N_2281,N_2321);
nor U2397 (N_2397,N_2284,N_2294);
nand U2398 (N_2398,N_2310,N_2296);
nor U2399 (N_2399,N_2304,N_2290);
nand U2400 (N_2400,N_2354,N_2345);
nand U2401 (N_2401,N_2364,N_2384);
or U2402 (N_2402,N_2378,N_2388);
xor U2403 (N_2403,N_2387,N_2376);
or U2404 (N_2404,N_2365,N_2352);
and U2405 (N_2405,N_2397,N_2394);
xor U2406 (N_2406,N_2368,N_2349);
nor U2407 (N_2407,N_2343,N_2357);
and U2408 (N_2408,N_2389,N_2363);
xor U2409 (N_2409,N_2340,N_2350);
xor U2410 (N_2410,N_2346,N_2370);
xnor U2411 (N_2411,N_2369,N_2379);
nand U2412 (N_2412,N_2382,N_2351);
or U2413 (N_2413,N_2347,N_2392);
nor U2414 (N_2414,N_2385,N_2391);
xor U2415 (N_2415,N_2375,N_2371);
or U2416 (N_2416,N_2367,N_2373);
nor U2417 (N_2417,N_2383,N_2372);
xor U2418 (N_2418,N_2355,N_2358);
nand U2419 (N_2419,N_2344,N_2360);
and U2420 (N_2420,N_2361,N_2396);
nand U2421 (N_2421,N_2399,N_2341);
or U2422 (N_2422,N_2386,N_2377);
nand U2423 (N_2423,N_2393,N_2380);
nor U2424 (N_2424,N_2374,N_2353);
nand U2425 (N_2425,N_2398,N_2390);
nand U2426 (N_2426,N_2356,N_2362);
xor U2427 (N_2427,N_2359,N_2342);
nor U2428 (N_2428,N_2381,N_2395);
or U2429 (N_2429,N_2366,N_2348);
or U2430 (N_2430,N_2372,N_2373);
or U2431 (N_2431,N_2385,N_2362);
or U2432 (N_2432,N_2355,N_2398);
or U2433 (N_2433,N_2367,N_2362);
nor U2434 (N_2434,N_2390,N_2343);
or U2435 (N_2435,N_2353,N_2360);
xnor U2436 (N_2436,N_2351,N_2384);
or U2437 (N_2437,N_2346,N_2398);
nand U2438 (N_2438,N_2382,N_2360);
nand U2439 (N_2439,N_2354,N_2376);
nor U2440 (N_2440,N_2374,N_2354);
and U2441 (N_2441,N_2355,N_2383);
or U2442 (N_2442,N_2390,N_2347);
and U2443 (N_2443,N_2393,N_2345);
and U2444 (N_2444,N_2376,N_2357);
and U2445 (N_2445,N_2393,N_2376);
nor U2446 (N_2446,N_2375,N_2359);
or U2447 (N_2447,N_2353,N_2377);
xnor U2448 (N_2448,N_2377,N_2345);
or U2449 (N_2449,N_2385,N_2379);
xor U2450 (N_2450,N_2377,N_2343);
nor U2451 (N_2451,N_2395,N_2380);
nor U2452 (N_2452,N_2394,N_2396);
xnor U2453 (N_2453,N_2367,N_2399);
or U2454 (N_2454,N_2391,N_2355);
or U2455 (N_2455,N_2349,N_2361);
nand U2456 (N_2456,N_2394,N_2357);
or U2457 (N_2457,N_2395,N_2358);
and U2458 (N_2458,N_2356,N_2347);
nor U2459 (N_2459,N_2373,N_2390);
nand U2460 (N_2460,N_2431,N_2443);
xor U2461 (N_2461,N_2417,N_2432);
xor U2462 (N_2462,N_2456,N_2427);
and U2463 (N_2463,N_2408,N_2428);
nor U2464 (N_2464,N_2405,N_2404);
and U2465 (N_2465,N_2413,N_2448);
and U2466 (N_2466,N_2442,N_2429);
xnor U2467 (N_2467,N_2421,N_2420);
and U2468 (N_2468,N_2446,N_2457);
nor U2469 (N_2469,N_2423,N_2458);
and U2470 (N_2470,N_2459,N_2419);
and U2471 (N_2471,N_2437,N_2411);
nor U2472 (N_2472,N_2425,N_2451);
or U2473 (N_2473,N_2410,N_2440);
or U2474 (N_2474,N_2426,N_2414);
nand U2475 (N_2475,N_2449,N_2401);
and U2476 (N_2476,N_2418,N_2452);
and U2477 (N_2477,N_2435,N_2424);
xnor U2478 (N_2478,N_2450,N_2403);
or U2479 (N_2479,N_2455,N_2453);
xor U2480 (N_2480,N_2422,N_2430);
or U2481 (N_2481,N_2400,N_2433);
nand U2482 (N_2482,N_2412,N_2447);
and U2483 (N_2483,N_2445,N_2438);
and U2484 (N_2484,N_2454,N_2416);
xor U2485 (N_2485,N_2407,N_2406);
and U2486 (N_2486,N_2409,N_2402);
xnor U2487 (N_2487,N_2415,N_2441);
nor U2488 (N_2488,N_2434,N_2444);
nand U2489 (N_2489,N_2436,N_2439);
nor U2490 (N_2490,N_2432,N_2405);
nor U2491 (N_2491,N_2403,N_2404);
or U2492 (N_2492,N_2416,N_2433);
xnor U2493 (N_2493,N_2419,N_2456);
xnor U2494 (N_2494,N_2455,N_2428);
or U2495 (N_2495,N_2433,N_2449);
and U2496 (N_2496,N_2449,N_2437);
nand U2497 (N_2497,N_2434,N_2443);
or U2498 (N_2498,N_2427,N_2451);
or U2499 (N_2499,N_2452,N_2444);
xor U2500 (N_2500,N_2426,N_2447);
xor U2501 (N_2501,N_2414,N_2452);
or U2502 (N_2502,N_2434,N_2408);
nor U2503 (N_2503,N_2410,N_2409);
nand U2504 (N_2504,N_2418,N_2421);
nand U2505 (N_2505,N_2400,N_2451);
and U2506 (N_2506,N_2427,N_2452);
or U2507 (N_2507,N_2435,N_2403);
xor U2508 (N_2508,N_2449,N_2421);
xor U2509 (N_2509,N_2433,N_2455);
or U2510 (N_2510,N_2420,N_2438);
or U2511 (N_2511,N_2453,N_2411);
or U2512 (N_2512,N_2456,N_2416);
nor U2513 (N_2513,N_2442,N_2434);
xor U2514 (N_2514,N_2405,N_2450);
and U2515 (N_2515,N_2406,N_2458);
or U2516 (N_2516,N_2438,N_2457);
and U2517 (N_2517,N_2441,N_2411);
and U2518 (N_2518,N_2440,N_2433);
nor U2519 (N_2519,N_2453,N_2434);
xnor U2520 (N_2520,N_2498,N_2508);
nand U2521 (N_2521,N_2505,N_2518);
nand U2522 (N_2522,N_2492,N_2473);
nand U2523 (N_2523,N_2460,N_2470);
nor U2524 (N_2524,N_2475,N_2472);
nand U2525 (N_2525,N_2488,N_2513);
nand U2526 (N_2526,N_2471,N_2463);
or U2527 (N_2527,N_2476,N_2497);
or U2528 (N_2528,N_2484,N_2495);
xnor U2529 (N_2529,N_2486,N_2464);
or U2530 (N_2530,N_2519,N_2465);
nor U2531 (N_2531,N_2462,N_2467);
xor U2532 (N_2532,N_2506,N_2480);
or U2533 (N_2533,N_2494,N_2485);
and U2534 (N_2534,N_2512,N_2491);
nor U2535 (N_2535,N_2503,N_2517);
or U2536 (N_2536,N_2466,N_2496);
nor U2537 (N_2537,N_2490,N_2489);
nor U2538 (N_2538,N_2502,N_2479);
or U2539 (N_2539,N_2500,N_2514);
and U2540 (N_2540,N_2516,N_2507);
or U2541 (N_2541,N_2483,N_2461);
or U2542 (N_2542,N_2511,N_2487);
or U2543 (N_2543,N_2510,N_2515);
nor U2544 (N_2544,N_2481,N_2509);
nand U2545 (N_2545,N_2504,N_2477);
or U2546 (N_2546,N_2493,N_2499);
nand U2547 (N_2547,N_2501,N_2468);
nand U2548 (N_2548,N_2469,N_2478);
xnor U2549 (N_2549,N_2482,N_2474);
xor U2550 (N_2550,N_2467,N_2480);
xor U2551 (N_2551,N_2514,N_2483);
nor U2552 (N_2552,N_2492,N_2477);
nor U2553 (N_2553,N_2471,N_2467);
nand U2554 (N_2554,N_2477,N_2481);
or U2555 (N_2555,N_2481,N_2501);
and U2556 (N_2556,N_2489,N_2461);
nand U2557 (N_2557,N_2489,N_2499);
and U2558 (N_2558,N_2480,N_2481);
or U2559 (N_2559,N_2517,N_2469);
nor U2560 (N_2560,N_2469,N_2462);
and U2561 (N_2561,N_2478,N_2461);
nand U2562 (N_2562,N_2486,N_2469);
xnor U2563 (N_2563,N_2511,N_2478);
nand U2564 (N_2564,N_2465,N_2505);
nand U2565 (N_2565,N_2497,N_2519);
and U2566 (N_2566,N_2498,N_2473);
nor U2567 (N_2567,N_2504,N_2517);
or U2568 (N_2568,N_2501,N_2503);
nand U2569 (N_2569,N_2519,N_2492);
or U2570 (N_2570,N_2472,N_2490);
xnor U2571 (N_2571,N_2464,N_2499);
nor U2572 (N_2572,N_2514,N_2506);
xnor U2573 (N_2573,N_2475,N_2492);
xnor U2574 (N_2574,N_2470,N_2481);
and U2575 (N_2575,N_2470,N_2486);
or U2576 (N_2576,N_2471,N_2503);
nand U2577 (N_2577,N_2483,N_2498);
nand U2578 (N_2578,N_2469,N_2518);
and U2579 (N_2579,N_2499,N_2502);
and U2580 (N_2580,N_2523,N_2531);
and U2581 (N_2581,N_2561,N_2522);
or U2582 (N_2582,N_2530,N_2574);
nand U2583 (N_2583,N_2545,N_2547);
or U2584 (N_2584,N_2566,N_2524);
and U2585 (N_2585,N_2563,N_2562);
and U2586 (N_2586,N_2544,N_2533);
nor U2587 (N_2587,N_2559,N_2550);
xnor U2588 (N_2588,N_2532,N_2539);
or U2589 (N_2589,N_2573,N_2554);
nor U2590 (N_2590,N_2579,N_2521);
and U2591 (N_2591,N_2540,N_2577);
nor U2592 (N_2592,N_2572,N_2549);
or U2593 (N_2593,N_2560,N_2567);
and U2594 (N_2594,N_2546,N_2536);
nand U2595 (N_2595,N_2552,N_2525);
and U2596 (N_2596,N_2548,N_2526);
and U2597 (N_2597,N_2534,N_2553);
or U2598 (N_2598,N_2576,N_2537);
nor U2599 (N_2599,N_2558,N_2538);
and U2600 (N_2600,N_2565,N_2535);
nor U2601 (N_2601,N_2520,N_2556);
nand U2602 (N_2602,N_2569,N_2543);
or U2603 (N_2603,N_2527,N_2578);
nor U2604 (N_2604,N_2542,N_2571);
and U2605 (N_2605,N_2570,N_2564);
nor U2606 (N_2606,N_2568,N_2529);
and U2607 (N_2607,N_2575,N_2557);
nor U2608 (N_2608,N_2555,N_2541);
and U2609 (N_2609,N_2528,N_2551);
or U2610 (N_2610,N_2522,N_2575);
nand U2611 (N_2611,N_2565,N_2523);
and U2612 (N_2612,N_2564,N_2521);
nand U2613 (N_2613,N_2543,N_2567);
nor U2614 (N_2614,N_2567,N_2531);
or U2615 (N_2615,N_2575,N_2563);
xnor U2616 (N_2616,N_2560,N_2550);
nand U2617 (N_2617,N_2537,N_2565);
or U2618 (N_2618,N_2568,N_2566);
xnor U2619 (N_2619,N_2576,N_2541);
nor U2620 (N_2620,N_2528,N_2522);
nor U2621 (N_2621,N_2575,N_2545);
or U2622 (N_2622,N_2541,N_2567);
nand U2623 (N_2623,N_2535,N_2577);
and U2624 (N_2624,N_2575,N_2576);
or U2625 (N_2625,N_2523,N_2576);
and U2626 (N_2626,N_2573,N_2562);
or U2627 (N_2627,N_2528,N_2524);
nor U2628 (N_2628,N_2548,N_2535);
or U2629 (N_2629,N_2534,N_2551);
nor U2630 (N_2630,N_2533,N_2575);
or U2631 (N_2631,N_2575,N_2551);
and U2632 (N_2632,N_2576,N_2561);
xor U2633 (N_2633,N_2569,N_2530);
nand U2634 (N_2634,N_2545,N_2577);
or U2635 (N_2635,N_2569,N_2563);
xnor U2636 (N_2636,N_2525,N_2530);
or U2637 (N_2637,N_2548,N_2545);
nand U2638 (N_2638,N_2532,N_2544);
or U2639 (N_2639,N_2545,N_2568);
and U2640 (N_2640,N_2614,N_2590);
and U2641 (N_2641,N_2598,N_2586);
and U2642 (N_2642,N_2628,N_2633);
xor U2643 (N_2643,N_2594,N_2589);
or U2644 (N_2644,N_2583,N_2617);
xnor U2645 (N_2645,N_2591,N_2581);
or U2646 (N_2646,N_2582,N_2580);
xor U2647 (N_2647,N_2636,N_2619);
nand U2648 (N_2648,N_2600,N_2604);
and U2649 (N_2649,N_2587,N_2601);
nor U2650 (N_2650,N_2595,N_2585);
or U2651 (N_2651,N_2597,N_2596);
nand U2652 (N_2652,N_2608,N_2635);
or U2653 (N_2653,N_2634,N_2629);
or U2654 (N_2654,N_2603,N_2627);
and U2655 (N_2655,N_2602,N_2615);
xor U2656 (N_2656,N_2593,N_2637);
and U2657 (N_2657,N_2618,N_2631);
xor U2658 (N_2658,N_2630,N_2620);
nand U2659 (N_2659,N_2623,N_2625);
nand U2660 (N_2660,N_2638,N_2621);
xnor U2661 (N_2661,N_2607,N_2613);
and U2662 (N_2662,N_2612,N_2592);
nor U2663 (N_2663,N_2639,N_2609);
nor U2664 (N_2664,N_2626,N_2611);
and U2665 (N_2665,N_2622,N_2632);
and U2666 (N_2666,N_2605,N_2599);
or U2667 (N_2667,N_2610,N_2588);
or U2668 (N_2668,N_2624,N_2616);
nand U2669 (N_2669,N_2584,N_2606);
xnor U2670 (N_2670,N_2619,N_2626);
and U2671 (N_2671,N_2613,N_2618);
or U2672 (N_2672,N_2617,N_2590);
nor U2673 (N_2673,N_2580,N_2587);
nor U2674 (N_2674,N_2625,N_2599);
xor U2675 (N_2675,N_2633,N_2593);
nor U2676 (N_2676,N_2594,N_2581);
nor U2677 (N_2677,N_2610,N_2583);
nand U2678 (N_2678,N_2619,N_2581);
nor U2679 (N_2679,N_2611,N_2599);
and U2680 (N_2680,N_2581,N_2603);
nand U2681 (N_2681,N_2596,N_2625);
xnor U2682 (N_2682,N_2598,N_2613);
nand U2683 (N_2683,N_2634,N_2606);
or U2684 (N_2684,N_2636,N_2624);
or U2685 (N_2685,N_2633,N_2589);
nor U2686 (N_2686,N_2629,N_2626);
nor U2687 (N_2687,N_2600,N_2585);
nand U2688 (N_2688,N_2601,N_2630);
and U2689 (N_2689,N_2611,N_2581);
xnor U2690 (N_2690,N_2602,N_2619);
or U2691 (N_2691,N_2604,N_2610);
or U2692 (N_2692,N_2631,N_2593);
nor U2693 (N_2693,N_2596,N_2615);
or U2694 (N_2694,N_2624,N_2587);
or U2695 (N_2695,N_2631,N_2584);
nand U2696 (N_2696,N_2608,N_2614);
nor U2697 (N_2697,N_2629,N_2587);
nor U2698 (N_2698,N_2636,N_2585);
xor U2699 (N_2699,N_2619,N_2604);
nor U2700 (N_2700,N_2668,N_2659);
nand U2701 (N_2701,N_2657,N_2677);
nand U2702 (N_2702,N_2640,N_2651);
nor U2703 (N_2703,N_2662,N_2653);
nand U2704 (N_2704,N_2666,N_2647);
xnor U2705 (N_2705,N_2655,N_2679);
and U2706 (N_2706,N_2669,N_2693);
and U2707 (N_2707,N_2671,N_2663);
or U2708 (N_2708,N_2697,N_2650);
nand U2709 (N_2709,N_2660,N_2642);
nor U2710 (N_2710,N_2695,N_2686);
nand U2711 (N_2711,N_2673,N_2661);
or U2712 (N_2712,N_2688,N_2690);
and U2713 (N_2713,N_2691,N_2645);
nand U2714 (N_2714,N_2641,N_2664);
nor U2715 (N_2715,N_2656,N_2675);
nor U2716 (N_2716,N_2694,N_2646);
nand U2717 (N_2717,N_2692,N_2665);
xor U2718 (N_2718,N_2681,N_2696);
nand U2719 (N_2719,N_2685,N_2654);
and U2720 (N_2720,N_2676,N_2698);
nor U2721 (N_2721,N_2672,N_2699);
nand U2722 (N_2722,N_2674,N_2687);
nor U2723 (N_2723,N_2680,N_2667);
or U2724 (N_2724,N_2683,N_2643);
or U2725 (N_2725,N_2689,N_2644);
nand U2726 (N_2726,N_2652,N_2682);
xor U2727 (N_2727,N_2670,N_2648);
xor U2728 (N_2728,N_2658,N_2684);
or U2729 (N_2729,N_2678,N_2649);
nor U2730 (N_2730,N_2665,N_2679);
and U2731 (N_2731,N_2641,N_2687);
and U2732 (N_2732,N_2649,N_2647);
or U2733 (N_2733,N_2660,N_2654);
and U2734 (N_2734,N_2689,N_2693);
nor U2735 (N_2735,N_2694,N_2674);
or U2736 (N_2736,N_2685,N_2682);
or U2737 (N_2737,N_2663,N_2678);
nand U2738 (N_2738,N_2656,N_2645);
nor U2739 (N_2739,N_2661,N_2691);
nand U2740 (N_2740,N_2691,N_2647);
xor U2741 (N_2741,N_2691,N_2689);
or U2742 (N_2742,N_2675,N_2679);
and U2743 (N_2743,N_2664,N_2686);
xor U2744 (N_2744,N_2695,N_2688);
xor U2745 (N_2745,N_2654,N_2677);
nand U2746 (N_2746,N_2642,N_2648);
or U2747 (N_2747,N_2651,N_2699);
and U2748 (N_2748,N_2650,N_2643);
nand U2749 (N_2749,N_2699,N_2674);
nor U2750 (N_2750,N_2671,N_2654);
or U2751 (N_2751,N_2659,N_2641);
nand U2752 (N_2752,N_2696,N_2688);
or U2753 (N_2753,N_2681,N_2651);
xnor U2754 (N_2754,N_2689,N_2651);
or U2755 (N_2755,N_2667,N_2692);
xnor U2756 (N_2756,N_2686,N_2685);
nor U2757 (N_2757,N_2650,N_2691);
nor U2758 (N_2758,N_2666,N_2665);
or U2759 (N_2759,N_2699,N_2662);
nor U2760 (N_2760,N_2712,N_2713);
xnor U2761 (N_2761,N_2753,N_2720);
and U2762 (N_2762,N_2755,N_2741);
and U2763 (N_2763,N_2757,N_2704);
xnor U2764 (N_2764,N_2710,N_2705);
or U2765 (N_2765,N_2727,N_2702);
and U2766 (N_2766,N_2723,N_2740);
and U2767 (N_2767,N_2724,N_2722);
and U2768 (N_2768,N_2735,N_2701);
nor U2769 (N_2769,N_2746,N_2758);
or U2770 (N_2770,N_2707,N_2745);
nand U2771 (N_2771,N_2728,N_2716);
and U2772 (N_2772,N_2731,N_2750);
and U2773 (N_2773,N_2749,N_2737);
nor U2774 (N_2774,N_2711,N_2706);
and U2775 (N_2775,N_2726,N_2752);
and U2776 (N_2776,N_2730,N_2747);
xnor U2777 (N_2777,N_2732,N_2715);
nand U2778 (N_2778,N_2738,N_2714);
nand U2779 (N_2779,N_2743,N_2754);
nand U2780 (N_2780,N_2708,N_2709);
nor U2781 (N_2781,N_2733,N_2718);
and U2782 (N_2782,N_2703,N_2756);
nand U2783 (N_2783,N_2700,N_2759);
nand U2784 (N_2784,N_2739,N_2742);
nand U2785 (N_2785,N_2744,N_2719);
nand U2786 (N_2786,N_2717,N_2721);
nand U2787 (N_2787,N_2736,N_2748);
and U2788 (N_2788,N_2725,N_2734);
nor U2789 (N_2789,N_2751,N_2729);
and U2790 (N_2790,N_2756,N_2717);
nand U2791 (N_2791,N_2741,N_2724);
or U2792 (N_2792,N_2710,N_2706);
or U2793 (N_2793,N_2750,N_2747);
nand U2794 (N_2794,N_2729,N_2703);
nor U2795 (N_2795,N_2758,N_2739);
or U2796 (N_2796,N_2744,N_2706);
nand U2797 (N_2797,N_2721,N_2727);
and U2798 (N_2798,N_2747,N_2724);
nor U2799 (N_2799,N_2715,N_2746);
xnor U2800 (N_2800,N_2719,N_2712);
xnor U2801 (N_2801,N_2734,N_2754);
nor U2802 (N_2802,N_2729,N_2743);
nand U2803 (N_2803,N_2717,N_2749);
xor U2804 (N_2804,N_2707,N_2744);
or U2805 (N_2805,N_2748,N_2727);
or U2806 (N_2806,N_2759,N_2758);
or U2807 (N_2807,N_2739,N_2704);
xor U2808 (N_2808,N_2758,N_2736);
nor U2809 (N_2809,N_2754,N_2711);
and U2810 (N_2810,N_2732,N_2711);
nand U2811 (N_2811,N_2724,N_2716);
nor U2812 (N_2812,N_2727,N_2706);
nor U2813 (N_2813,N_2718,N_2732);
xnor U2814 (N_2814,N_2711,N_2756);
nor U2815 (N_2815,N_2740,N_2708);
and U2816 (N_2816,N_2726,N_2742);
nand U2817 (N_2817,N_2711,N_2733);
nand U2818 (N_2818,N_2751,N_2711);
nor U2819 (N_2819,N_2713,N_2708);
xnor U2820 (N_2820,N_2804,N_2817);
nand U2821 (N_2821,N_2798,N_2775);
nor U2822 (N_2822,N_2762,N_2791);
or U2823 (N_2823,N_2806,N_2760);
nand U2824 (N_2824,N_2789,N_2765);
or U2825 (N_2825,N_2777,N_2807);
nor U2826 (N_2826,N_2763,N_2761);
xor U2827 (N_2827,N_2802,N_2782);
xor U2828 (N_2828,N_2784,N_2801);
xor U2829 (N_2829,N_2813,N_2787);
and U2830 (N_2830,N_2800,N_2788);
nor U2831 (N_2831,N_2797,N_2781);
nand U2832 (N_2832,N_2816,N_2786);
xor U2833 (N_2833,N_2805,N_2814);
and U2834 (N_2834,N_2792,N_2803);
nor U2835 (N_2835,N_2808,N_2772);
or U2836 (N_2836,N_2773,N_2812);
xnor U2837 (N_2837,N_2769,N_2815);
nand U2838 (N_2838,N_2810,N_2809);
nand U2839 (N_2839,N_2818,N_2774);
xor U2840 (N_2840,N_2764,N_2794);
xnor U2841 (N_2841,N_2776,N_2767);
xor U2842 (N_2842,N_2785,N_2771);
xor U2843 (N_2843,N_2795,N_2766);
xor U2844 (N_2844,N_2796,N_2783);
xnor U2845 (N_2845,N_2790,N_2811);
and U2846 (N_2846,N_2768,N_2778);
or U2847 (N_2847,N_2779,N_2780);
or U2848 (N_2848,N_2799,N_2819);
nor U2849 (N_2849,N_2770,N_2793);
and U2850 (N_2850,N_2773,N_2772);
or U2851 (N_2851,N_2783,N_2808);
nand U2852 (N_2852,N_2819,N_2765);
or U2853 (N_2853,N_2771,N_2805);
nor U2854 (N_2854,N_2765,N_2806);
or U2855 (N_2855,N_2764,N_2779);
nand U2856 (N_2856,N_2761,N_2796);
and U2857 (N_2857,N_2767,N_2805);
xnor U2858 (N_2858,N_2768,N_2809);
or U2859 (N_2859,N_2797,N_2789);
nand U2860 (N_2860,N_2803,N_2807);
and U2861 (N_2861,N_2796,N_2785);
or U2862 (N_2862,N_2796,N_2772);
nand U2863 (N_2863,N_2799,N_2785);
and U2864 (N_2864,N_2812,N_2802);
and U2865 (N_2865,N_2779,N_2782);
xnor U2866 (N_2866,N_2779,N_2801);
nor U2867 (N_2867,N_2787,N_2775);
nand U2868 (N_2868,N_2783,N_2790);
or U2869 (N_2869,N_2774,N_2795);
nor U2870 (N_2870,N_2760,N_2813);
and U2871 (N_2871,N_2787,N_2793);
nand U2872 (N_2872,N_2794,N_2806);
nand U2873 (N_2873,N_2814,N_2774);
and U2874 (N_2874,N_2812,N_2814);
or U2875 (N_2875,N_2791,N_2767);
and U2876 (N_2876,N_2760,N_2773);
nand U2877 (N_2877,N_2762,N_2810);
or U2878 (N_2878,N_2768,N_2786);
xnor U2879 (N_2879,N_2777,N_2818);
nor U2880 (N_2880,N_2869,N_2825);
or U2881 (N_2881,N_2826,N_2823);
or U2882 (N_2882,N_2862,N_2863);
xnor U2883 (N_2883,N_2832,N_2836);
or U2884 (N_2884,N_2870,N_2833);
and U2885 (N_2885,N_2822,N_2878);
nor U2886 (N_2886,N_2875,N_2850);
or U2887 (N_2887,N_2855,N_2866);
nand U2888 (N_2888,N_2841,N_2824);
nor U2889 (N_2889,N_2837,N_2846);
or U2890 (N_2890,N_2834,N_2872);
and U2891 (N_2891,N_2859,N_2827);
nand U2892 (N_2892,N_2844,N_2830);
nor U2893 (N_2893,N_2865,N_2845);
xnor U2894 (N_2894,N_2858,N_2847);
nor U2895 (N_2895,N_2842,N_2828);
nor U2896 (N_2896,N_2876,N_2856);
and U2897 (N_2897,N_2874,N_2871);
xor U2898 (N_2898,N_2849,N_2839);
nor U2899 (N_2899,N_2835,N_2860);
and U2900 (N_2900,N_2829,N_2852);
xor U2901 (N_2901,N_2840,N_2854);
nand U2902 (N_2902,N_2867,N_2843);
or U2903 (N_2903,N_2861,N_2820);
nand U2904 (N_2904,N_2831,N_2857);
nand U2905 (N_2905,N_2877,N_2879);
nand U2906 (N_2906,N_2864,N_2821);
nor U2907 (N_2907,N_2851,N_2848);
nor U2908 (N_2908,N_2873,N_2868);
or U2909 (N_2909,N_2853,N_2838);
or U2910 (N_2910,N_2852,N_2850);
and U2911 (N_2911,N_2868,N_2862);
or U2912 (N_2912,N_2879,N_2833);
nand U2913 (N_2913,N_2855,N_2826);
nand U2914 (N_2914,N_2866,N_2863);
or U2915 (N_2915,N_2866,N_2844);
nor U2916 (N_2916,N_2849,N_2853);
or U2917 (N_2917,N_2824,N_2853);
nor U2918 (N_2918,N_2871,N_2876);
nand U2919 (N_2919,N_2835,N_2866);
nor U2920 (N_2920,N_2844,N_2846);
and U2921 (N_2921,N_2858,N_2860);
and U2922 (N_2922,N_2822,N_2840);
xor U2923 (N_2923,N_2859,N_2834);
nand U2924 (N_2924,N_2879,N_2867);
nor U2925 (N_2925,N_2836,N_2865);
nand U2926 (N_2926,N_2870,N_2838);
xnor U2927 (N_2927,N_2855,N_2842);
xor U2928 (N_2928,N_2831,N_2876);
nor U2929 (N_2929,N_2864,N_2873);
nor U2930 (N_2930,N_2870,N_2839);
or U2931 (N_2931,N_2853,N_2846);
or U2932 (N_2932,N_2836,N_2875);
xor U2933 (N_2933,N_2864,N_2835);
and U2934 (N_2934,N_2824,N_2859);
nand U2935 (N_2935,N_2870,N_2821);
or U2936 (N_2936,N_2844,N_2851);
xor U2937 (N_2937,N_2849,N_2865);
or U2938 (N_2938,N_2852,N_2851);
nand U2939 (N_2939,N_2841,N_2834);
or U2940 (N_2940,N_2917,N_2889);
nand U2941 (N_2941,N_2935,N_2903);
nand U2942 (N_2942,N_2931,N_2904);
xnor U2943 (N_2943,N_2936,N_2890);
nor U2944 (N_2944,N_2883,N_2934);
nand U2945 (N_2945,N_2881,N_2938);
xnor U2946 (N_2946,N_2929,N_2884);
and U2947 (N_2947,N_2913,N_2907);
nor U2948 (N_2948,N_2882,N_2886);
xor U2949 (N_2949,N_2927,N_2885);
or U2950 (N_2950,N_2902,N_2900);
nor U2951 (N_2951,N_2901,N_2896);
nor U2952 (N_2952,N_2887,N_2937);
xor U2953 (N_2953,N_2891,N_2919);
or U2954 (N_2954,N_2928,N_2924);
xnor U2955 (N_2955,N_2918,N_2894);
nand U2956 (N_2956,N_2926,N_2910);
xor U2957 (N_2957,N_2939,N_2906);
xor U2958 (N_2958,N_2925,N_2915);
or U2959 (N_2959,N_2893,N_2911);
nand U2960 (N_2960,N_2914,N_2908);
and U2961 (N_2961,N_2898,N_2895);
nand U2962 (N_2962,N_2920,N_2880);
or U2963 (N_2963,N_2923,N_2916);
and U2964 (N_2964,N_2932,N_2912);
xor U2965 (N_2965,N_2922,N_2897);
nor U2966 (N_2966,N_2899,N_2933);
xor U2967 (N_2967,N_2888,N_2892);
nand U2968 (N_2968,N_2905,N_2921);
nor U2969 (N_2969,N_2930,N_2909);
or U2970 (N_2970,N_2910,N_2892);
xnor U2971 (N_2971,N_2931,N_2934);
and U2972 (N_2972,N_2928,N_2903);
or U2973 (N_2973,N_2885,N_2906);
and U2974 (N_2974,N_2935,N_2912);
xnor U2975 (N_2975,N_2909,N_2895);
and U2976 (N_2976,N_2884,N_2914);
and U2977 (N_2977,N_2938,N_2906);
nand U2978 (N_2978,N_2907,N_2900);
nor U2979 (N_2979,N_2903,N_2912);
or U2980 (N_2980,N_2939,N_2894);
or U2981 (N_2981,N_2927,N_2938);
and U2982 (N_2982,N_2917,N_2921);
nor U2983 (N_2983,N_2880,N_2911);
and U2984 (N_2984,N_2920,N_2935);
or U2985 (N_2985,N_2896,N_2894);
nor U2986 (N_2986,N_2920,N_2919);
and U2987 (N_2987,N_2880,N_2921);
xor U2988 (N_2988,N_2892,N_2928);
nor U2989 (N_2989,N_2916,N_2936);
and U2990 (N_2990,N_2906,N_2908);
or U2991 (N_2991,N_2928,N_2912);
xor U2992 (N_2992,N_2918,N_2892);
and U2993 (N_2993,N_2916,N_2897);
nor U2994 (N_2994,N_2880,N_2917);
nand U2995 (N_2995,N_2890,N_2898);
nor U2996 (N_2996,N_2889,N_2899);
or U2997 (N_2997,N_2925,N_2937);
nor U2998 (N_2998,N_2912,N_2920);
and U2999 (N_2999,N_2900,N_2893);
xnor UO_0 (O_0,N_2955,N_2946);
nor UO_1 (O_1,N_2991,N_2997);
nand UO_2 (O_2,N_2950,N_2943);
xor UO_3 (O_3,N_2948,N_2999);
and UO_4 (O_4,N_2978,N_2979);
nand UO_5 (O_5,N_2956,N_2988);
nand UO_6 (O_6,N_2945,N_2992);
nand UO_7 (O_7,N_2982,N_2989);
or UO_8 (O_8,N_2957,N_2990);
or UO_9 (O_9,N_2993,N_2976);
or UO_10 (O_10,N_2954,N_2949);
and UO_11 (O_11,N_2940,N_2983);
nor UO_12 (O_12,N_2942,N_2944);
and UO_13 (O_13,N_2994,N_2941);
nor UO_14 (O_14,N_2973,N_2987);
xnor UO_15 (O_15,N_2961,N_2971);
nor UO_16 (O_16,N_2996,N_2952);
nand UO_17 (O_17,N_2965,N_2968);
nand UO_18 (O_18,N_2977,N_2962);
nor UO_19 (O_19,N_2986,N_2972);
nor UO_20 (O_20,N_2984,N_2995);
nand UO_21 (O_21,N_2980,N_2947);
or UO_22 (O_22,N_2970,N_2998);
and UO_23 (O_23,N_2964,N_2969);
or UO_24 (O_24,N_2958,N_2966);
nand UO_25 (O_25,N_2951,N_2963);
and UO_26 (O_26,N_2953,N_2959);
nand UO_27 (O_27,N_2974,N_2967);
or UO_28 (O_28,N_2975,N_2985);
xnor UO_29 (O_29,N_2960,N_2981);
nand UO_30 (O_30,N_2973,N_2985);
xnor UO_31 (O_31,N_2987,N_2946);
xnor UO_32 (O_32,N_2972,N_2961);
nor UO_33 (O_33,N_2985,N_2960);
and UO_34 (O_34,N_2967,N_2995);
nor UO_35 (O_35,N_2951,N_2992);
or UO_36 (O_36,N_2969,N_2976);
and UO_37 (O_37,N_2942,N_2963);
or UO_38 (O_38,N_2946,N_2967);
or UO_39 (O_39,N_2965,N_2988);
and UO_40 (O_40,N_2954,N_2983);
or UO_41 (O_41,N_2997,N_2996);
or UO_42 (O_42,N_2950,N_2960);
nor UO_43 (O_43,N_2969,N_2989);
and UO_44 (O_44,N_2983,N_2993);
and UO_45 (O_45,N_2977,N_2972);
or UO_46 (O_46,N_2949,N_2965);
xor UO_47 (O_47,N_2944,N_2949);
and UO_48 (O_48,N_2970,N_2999);
xnor UO_49 (O_49,N_2943,N_2957);
nor UO_50 (O_50,N_2980,N_2975);
or UO_51 (O_51,N_2961,N_2942);
xnor UO_52 (O_52,N_2993,N_2949);
and UO_53 (O_53,N_2972,N_2953);
or UO_54 (O_54,N_2993,N_2945);
and UO_55 (O_55,N_2966,N_2948);
or UO_56 (O_56,N_2945,N_2976);
or UO_57 (O_57,N_2967,N_2964);
xnor UO_58 (O_58,N_2957,N_2959);
nand UO_59 (O_59,N_2995,N_2994);
nand UO_60 (O_60,N_2975,N_2964);
nand UO_61 (O_61,N_2968,N_2977);
nand UO_62 (O_62,N_2944,N_2982);
and UO_63 (O_63,N_2958,N_2957);
and UO_64 (O_64,N_2987,N_2956);
nand UO_65 (O_65,N_2974,N_2973);
xor UO_66 (O_66,N_2944,N_2983);
or UO_67 (O_67,N_2950,N_2983);
nand UO_68 (O_68,N_2995,N_2950);
or UO_69 (O_69,N_2951,N_2956);
xnor UO_70 (O_70,N_2982,N_2985);
and UO_71 (O_71,N_2985,N_2948);
or UO_72 (O_72,N_2953,N_2975);
and UO_73 (O_73,N_2986,N_2943);
and UO_74 (O_74,N_2979,N_2963);
xnor UO_75 (O_75,N_2998,N_2990);
or UO_76 (O_76,N_2995,N_2990);
nand UO_77 (O_77,N_2960,N_2997);
or UO_78 (O_78,N_2972,N_2984);
xnor UO_79 (O_79,N_2977,N_2958);
and UO_80 (O_80,N_2944,N_2980);
xnor UO_81 (O_81,N_2990,N_2961);
nor UO_82 (O_82,N_2997,N_2967);
and UO_83 (O_83,N_2949,N_2953);
or UO_84 (O_84,N_2992,N_2998);
xnor UO_85 (O_85,N_2949,N_2940);
nand UO_86 (O_86,N_2942,N_2995);
xnor UO_87 (O_87,N_2982,N_2957);
nor UO_88 (O_88,N_2973,N_2978);
nand UO_89 (O_89,N_2985,N_2952);
xnor UO_90 (O_90,N_2963,N_2991);
xor UO_91 (O_91,N_2991,N_2973);
or UO_92 (O_92,N_2975,N_2951);
or UO_93 (O_93,N_2949,N_2942);
and UO_94 (O_94,N_2999,N_2984);
nor UO_95 (O_95,N_2978,N_2990);
nand UO_96 (O_96,N_2990,N_2969);
nor UO_97 (O_97,N_2974,N_2961);
or UO_98 (O_98,N_2952,N_2948);
nand UO_99 (O_99,N_2946,N_2944);
nor UO_100 (O_100,N_2993,N_2967);
or UO_101 (O_101,N_2968,N_2983);
xor UO_102 (O_102,N_2954,N_2996);
xor UO_103 (O_103,N_2978,N_2974);
nor UO_104 (O_104,N_2990,N_2966);
nand UO_105 (O_105,N_2967,N_2951);
and UO_106 (O_106,N_2945,N_2952);
xnor UO_107 (O_107,N_2951,N_2990);
or UO_108 (O_108,N_2990,N_2971);
and UO_109 (O_109,N_2979,N_2954);
or UO_110 (O_110,N_2979,N_2967);
and UO_111 (O_111,N_2979,N_2984);
nor UO_112 (O_112,N_2966,N_2978);
or UO_113 (O_113,N_2946,N_2959);
nor UO_114 (O_114,N_2976,N_2984);
nor UO_115 (O_115,N_2984,N_2961);
and UO_116 (O_116,N_2980,N_2978);
xor UO_117 (O_117,N_2957,N_2964);
xnor UO_118 (O_118,N_2971,N_2999);
and UO_119 (O_119,N_2945,N_2964);
and UO_120 (O_120,N_2996,N_2955);
nand UO_121 (O_121,N_2991,N_2995);
xor UO_122 (O_122,N_2974,N_2994);
xnor UO_123 (O_123,N_2944,N_2979);
and UO_124 (O_124,N_2972,N_2993);
or UO_125 (O_125,N_2995,N_2955);
nor UO_126 (O_126,N_2992,N_2987);
nand UO_127 (O_127,N_2952,N_2961);
xnor UO_128 (O_128,N_2946,N_2963);
nor UO_129 (O_129,N_2956,N_2953);
and UO_130 (O_130,N_2952,N_2992);
or UO_131 (O_131,N_2947,N_2971);
nor UO_132 (O_132,N_2976,N_2944);
nand UO_133 (O_133,N_2986,N_2983);
nor UO_134 (O_134,N_2993,N_2988);
xnor UO_135 (O_135,N_2973,N_2968);
xor UO_136 (O_136,N_2989,N_2993);
nor UO_137 (O_137,N_2983,N_2994);
or UO_138 (O_138,N_2951,N_2961);
xor UO_139 (O_139,N_2966,N_2943);
xnor UO_140 (O_140,N_2992,N_2968);
xnor UO_141 (O_141,N_2967,N_2941);
nor UO_142 (O_142,N_2947,N_2941);
xnor UO_143 (O_143,N_2996,N_2982);
and UO_144 (O_144,N_2980,N_2981);
xnor UO_145 (O_145,N_2996,N_2998);
and UO_146 (O_146,N_2981,N_2942);
and UO_147 (O_147,N_2977,N_2992);
nand UO_148 (O_148,N_2964,N_2956);
nand UO_149 (O_149,N_2994,N_2982);
xor UO_150 (O_150,N_2947,N_2984);
nor UO_151 (O_151,N_2982,N_2980);
or UO_152 (O_152,N_2975,N_2973);
nand UO_153 (O_153,N_2966,N_2996);
nand UO_154 (O_154,N_2953,N_2989);
nor UO_155 (O_155,N_2970,N_2978);
xor UO_156 (O_156,N_2973,N_2966);
and UO_157 (O_157,N_2954,N_2980);
nand UO_158 (O_158,N_2965,N_2989);
xnor UO_159 (O_159,N_2986,N_2961);
nor UO_160 (O_160,N_2979,N_2996);
or UO_161 (O_161,N_2942,N_2979);
or UO_162 (O_162,N_2940,N_2964);
or UO_163 (O_163,N_2947,N_2952);
nand UO_164 (O_164,N_2999,N_2968);
nand UO_165 (O_165,N_2962,N_2941);
or UO_166 (O_166,N_2995,N_2956);
nor UO_167 (O_167,N_2952,N_2995);
nor UO_168 (O_168,N_2957,N_2946);
nor UO_169 (O_169,N_2940,N_2959);
xnor UO_170 (O_170,N_2956,N_2970);
and UO_171 (O_171,N_2991,N_2941);
xnor UO_172 (O_172,N_2962,N_2976);
xnor UO_173 (O_173,N_2948,N_2943);
xor UO_174 (O_174,N_2968,N_2947);
nor UO_175 (O_175,N_2967,N_2973);
nor UO_176 (O_176,N_2941,N_2940);
and UO_177 (O_177,N_2998,N_2980);
and UO_178 (O_178,N_2947,N_2979);
nor UO_179 (O_179,N_2983,N_2947);
xor UO_180 (O_180,N_2981,N_2990);
or UO_181 (O_181,N_2999,N_2985);
nand UO_182 (O_182,N_2992,N_2966);
and UO_183 (O_183,N_2979,N_2959);
xnor UO_184 (O_184,N_2957,N_2960);
nand UO_185 (O_185,N_2947,N_2955);
nand UO_186 (O_186,N_2948,N_2940);
nand UO_187 (O_187,N_2979,N_2956);
or UO_188 (O_188,N_2941,N_2975);
and UO_189 (O_189,N_2956,N_2991);
nor UO_190 (O_190,N_2984,N_2989);
and UO_191 (O_191,N_2995,N_2977);
or UO_192 (O_192,N_2991,N_2943);
and UO_193 (O_193,N_2948,N_2992);
and UO_194 (O_194,N_2998,N_2982);
nor UO_195 (O_195,N_2997,N_2956);
nand UO_196 (O_196,N_2949,N_2967);
or UO_197 (O_197,N_2978,N_2993);
or UO_198 (O_198,N_2997,N_2992);
and UO_199 (O_199,N_2963,N_2976);
and UO_200 (O_200,N_2960,N_2954);
nand UO_201 (O_201,N_2968,N_2991);
xor UO_202 (O_202,N_2977,N_2951);
and UO_203 (O_203,N_2946,N_2981);
and UO_204 (O_204,N_2997,N_2977);
nand UO_205 (O_205,N_2948,N_2961);
nor UO_206 (O_206,N_2985,N_2998);
or UO_207 (O_207,N_2940,N_2953);
and UO_208 (O_208,N_2972,N_2981);
or UO_209 (O_209,N_2949,N_2968);
nand UO_210 (O_210,N_2963,N_2987);
nor UO_211 (O_211,N_2942,N_2954);
nand UO_212 (O_212,N_2983,N_2964);
nand UO_213 (O_213,N_2970,N_2979);
or UO_214 (O_214,N_2963,N_2970);
xnor UO_215 (O_215,N_2944,N_2969);
nand UO_216 (O_216,N_2949,N_2963);
or UO_217 (O_217,N_2976,N_2965);
nor UO_218 (O_218,N_2982,N_2975);
nor UO_219 (O_219,N_2981,N_2999);
and UO_220 (O_220,N_2964,N_2951);
xnor UO_221 (O_221,N_2998,N_2995);
xor UO_222 (O_222,N_2991,N_2984);
nand UO_223 (O_223,N_2971,N_2941);
or UO_224 (O_224,N_2988,N_2970);
or UO_225 (O_225,N_2949,N_2941);
and UO_226 (O_226,N_2974,N_2940);
nand UO_227 (O_227,N_2994,N_2942);
and UO_228 (O_228,N_2945,N_2987);
nor UO_229 (O_229,N_2964,N_2988);
nand UO_230 (O_230,N_2957,N_2944);
and UO_231 (O_231,N_2990,N_2973);
xnor UO_232 (O_232,N_2995,N_2972);
nand UO_233 (O_233,N_2991,N_2980);
and UO_234 (O_234,N_2956,N_2982);
nand UO_235 (O_235,N_2969,N_2958);
nor UO_236 (O_236,N_2994,N_2980);
nand UO_237 (O_237,N_2984,N_2953);
nand UO_238 (O_238,N_2972,N_2948);
or UO_239 (O_239,N_2943,N_2962);
and UO_240 (O_240,N_2950,N_2963);
or UO_241 (O_241,N_2972,N_2970);
nand UO_242 (O_242,N_2959,N_2980);
xor UO_243 (O_243,N_2966,N_2995);
or UO_244 (O_244,N_2985,N_2942);
and UO_245 (O_245,N_2983,N_2941);
nand UO_246 (O_246,N_2960,N_2956);
nor UO_247 (O_247,N_2950,N_2968);
nand UO_248 (O_248,N_2962,N_2966);
nor UO_249 (O_249,N_2953,N_2986);
nor UO_250 (O_250,N_2947,N_2965);
or UO_251 (O_251,N_2972,N_2966);
nor UO_252 (O_252,N_2975,N_2954);
or UO_253 (O_253,N_2999,N_2993);
nand UO_254 (O_254,N_2943,N_2977);
and UO_255 (O_255,N_2992,N_2996);
nor UO_256 (O_256,N_2974,N_2942);
nand UO_257 (O_257,N_2978,N_2963);
nand UO_258 (O_258,N_2967,N_2955);
nand UO_259 (O_259,N_2943,N_2941);
or UO_260 (O_260,N_2952,N_2973);
nand UO_261 (O_261,N_2943,N_2972);
xor UO_262 (O_262,N_2970,N_2961);
or UO_263 (O_263,N_2966,N_2980);
xor UO_264 (O_264,N_2964,N_2973);
and UO_265 (O_265,N_2991,N_2982);
xnor UO_266 (O_266,N_2987,N_2976);
nor UO_267 (O_267,N_2968,N_2993);
nor UO_268 (O_268,N_2948,N_2969);
and UO_269 (O_269,N_2969,N_2997);
and UO_270 (O_270,N_2980,N_2953);
nand UO_271 (O_271,N_2942,N_2993);
nor UO_272 (O_272,N_2969,N_2986);
nand UO_273 (O_273,N_2987,N_2952);
nor UO_274 (O_274,N_2957,N_2977);
and UO_275 (O_275,N_2994,N_2968);
nand UO_276 (O_276,N_2979,N_2971);
nand UO_277 (O_277,N_2982,N_2963);
nand UO_278 (O_278,N_2992,N_2950);
xnor UO_279 (O_279,N_2981,N_2974);
nor UO_280 (O_280,N_2952,N_2960);
nand UO_281 (O_281,N_2946,N_2940);
and UO_282 (O_282,N_2949,N_2957);
or UO_283 (O_283,N_2943,N_2944);
nand UO_284 (O_284,N_2950,N_2985);
nor UO_285 (O_285,N_2962,N_2963);
and UO_286 (O_286,N_2940,N_2965);
or UO_287 (O_287,N_2956,N_2948);
nor UO_288 (O_288,N_2966,N_2961);
and UO_289 (O_289,N_2988,N_2995);
or UO_290 (O_290,N_2948,N_2996);
xor UO_291 (O_291,N_2977,N_2975);
and UO_292 (O_292,N_2966,N_2983);
nand UO_293 (O_293,N_2985,N_2958);
or UO_294 (O_294,N_2968,N_2984);
xor UO_295 (O_295,N_2971,N_2946);
and UO_296 (O_296,N_2978,N_2989);
xnor UO_297 (O_297,N_2952,N_2986);
nor UO_298 (O_298,N_2990,N_2947);
or UO_299 (O_299,N_2997,N_2947);
nand UO_300 (O_300,N_2941,N_2984);
or UO_301 (O_301,N_2985,N_2954);
nand UO_302 (O_302,N_2951,N_2984);
xor UO_303 (O_303,N_2961,N_2968);
xor UO_304 (O_304,N_2960,N_2978);
nand UO_305 (O_305,N_2960,N_2998);
nor UO_306 (O_306,N_2989,N_2960);
or UO_307 (O_307,N_2975,N_2999);
and UO_308 (O_308,N_2987,N_2948);
nand UO_309 (O_309,N_2960,N_2999);
nor UO_310 (O_310,N_2985,N_2987);
nor UO_311 (O_311,N_2992,N_2969);
or UO_312 (O_312,N_2999,N_2944);
nand UO_313 (O_313,N_2946,N_2960);
or UO_314 (O_314,N_2999,N_2963);
and UO_315 (O_315,N_2984,N_2983);
xor UO_316 (O_316,N_2942,N_2962);
nor UO_317 (O_317,N_2959,N_2949);
nor UO_318 (O_318,N_2968,N_2967);
and UO_319 (O_319,N_2977,N_2966);
or UO_320 (O_320,N_2952,N_2953);
and UO_321 (O_321,N_2944,N_2963);
nand UO_322 (O_322,N_2946,N_2961);
xnor UO_323 (O_323,N_2960,N_2964);
xnor UO_324 (O_324,N_2985,N_2947);
xnor UO_325 (O_325,N_2950,N_2945);
and UO_326 (O_326,N_2998,N_2975);
nand UO_327 (O_327,N_2959,N_2941);
and UO_328 (O_328,N_2978,N_2954);
and UO_329 (O_329,N_2978,N_2986);
xor UO_330 (O_330,N_2944,N_2948);
nand UO_331 (O_331,N_2990,N_2999);
nand UO_332 (O_332,N_2960,N_2990);
xnor UO_333 (O_333,N_2998,N_2949);
nor UO_334 (O_334,N_2941,N_2989);
nor UO_335 (O_335,N_2960,N_2974);
or UO_336 (O_336,N_2969,N_2959);
or UO_337 (O_337,N_2941,N_2968);
nand UO_338 (O_338,N_2988,N_2999);
nand UO_339 (O_339,N_2974,N_2970);
and UO_340 (O_340,N_2974,N_2987);
or UO_341 (O_341,N_2960,N_2969);
nor UO_342 (O_342,N_2989,N_2983);
nor UO_343 (O_343,N_2978,N_2981);
and UO_344 (O_344,N_2949,N_2976);
nor UO_345 (O_345,N_2955,N_2988);
xor UO_346 (O_346,N_2954,N_2973);
or UO_347 (O_347,N_2983,N_2946);
nand UO_348 (O_348,N_2941,N_2944);
nor UO_349 (O_349,N_2955,N_2966);
and UO_350 (O_350,N_2972,N_2964);
nor UO_351 (O_351,N_2943,N_2990);
and UO_352 (O_352,N_2940,N_2954);
xnor UO_353 (O_353,N_2987,N_2991);
or UO_354 (O_354,N_2950,N_2967);
and UO_355 (O_355,N_2984,N_2944);
and UO_356 (O_356,N_2951,N_2965);
nor UO_357 (O_357,N_2970,N_2997);
nand UO_358 (O_358,N_2971,N_2967);
nor UO_359 (O_359,N_2997,N_2995);
or UO_360 (O_360,N_2943,N_2971);
nor UO_361 (O_361,N_2967,N_2987);
and UO_362 (O_362,N_2992,N_2985);
nor UO_363 (O_363,N_2976,N_2983);
and UO_364 (O_364,N_2990,N_2982);
or UO_365 (O_365,N_2969,N_2965);
or UO_366 (O_366,N_2945,N_2940);
nor UO_367 (O_367,N_2994,N_2988);
or UO_368 (O_368,N_2977,N_2950);
nand UO_369 (O_369,N_2983,N_2961);
nor UO_370 (O_370,N_2947,N_2964);
or UO_371 (O_371,N_2982,N_2943);
nand UO_372 (O_372,N_2979,N_2988);
nor UO_373 (O_373,N_2966,N_2951);
and UO_374 (O_374,N_2943,N_2946);
nand UO_375 (O_375,N_2957,N_2994);
or UO_376 (O_376,N_2969,N_2988);
or UO_377 (O_377,N_2951,N_2979);
and UO_378 (O_378,N_2976,N_2973);
nand UO_379 (O_379,N_2957,N_2972);
or UO_380 (O_380,N_2944,N_2967);
and UO_381 (O_381,N_2972,N_2944);
or UO_382 (O_382,N_2950,N_2951);
and UO_383 (O_383,N_2957,N_2968);
or UO_384 (O_384,N_2955,N_2998);
nor UO_385 (O_385,N_2960,N_2951);
xnor UO_386 (O_386,N_2987,N_2990);
nor UO_387 (O_387,N_2953,N_2954);
xor UO_388 (O_388,N_2965,N_2967);
nor UO_389 (O_389,N_2954,N_2955);
nand UO_390 (O_390,N_2991,N_2985);
nand UO_391 (O_391,N_2972,N_2979);
nor UO_392 (O_392,N_2953,N_2970);
and UO_393 (O_393,N_2984,N_2952);
and UO_394 (O_394,N_2975,N_2965);
xnor UO_395 (O_395,N_2970,N_2960);
nor UO_396 (O_396,N_2963,N_2947);
and UO_397 (O_397,N_2951,N_2969);
nand UO_398 (O_398,N_2951,N_2942);
xor UO_399 (O_399,N_2967,N_2981);
xnor UO_400 (O_400,N_2950,N_2941);
nor UO_401 (O_401,N_2991,N_2993);
or UO_402 (O_402,N_2973,N_2940);
xor UO_403 (O_403,N_2987,N_2962);
or UO_404 (O_404,N_2947,N_2991);
or UO_405 (O_405,N_2986,N_2984);
nor UO_406 (O_406,N_2945,N_2959);
nor UO_407 (O_407,N_2947,N_2982);
or UO_408 (O_408,N_2970,N_2952);
and UO_409 (O_409,N_2944,N_2994);
nand UO_410 (O_410,N_2985,N_2959);
or UO_411 (O_411,N_2978,N_2995);
or UO_412 (O_412,N_2958,N_2984);
or UO_413 (O_413,N_2958,N_2971);
and UO_414 (O_414,N_2989,N_2962);
xnor UO_415 (O_415,N_2971,N_2980);
nor UO_416 (O_416,N_2975,N_2957);
nor UO_417 (O_417,N_2997,N_2961);
and UO_418 (O_418,N_2959,N_2995);
xnor UO_419 (O_419,N_2956,N_2941);
and UO_420 (O_420,N_2965,N_2953);
xor UO_421 (O_421,N_2986,N_2992);
xnor UO_422 (O_422,N_2991,N_2961);
xnor UO_423 (O_423,N_2971,N_2991);
nand UO_424 (O_424,N_2959,N_2964);
xnor UO_425 (O_425,N_2947,N_2946);
nand UO_426 (O_426,N_2973,N_2996);
xnor UO_427 (O_427,N_2941,N_2952);
nand UO_428 (O_428,N_2943,N_2994);
xnor UO_429 (O_429,N_2980,N_2992);
nor UO_430 (O_430,N_2974,N_2985);
nor UO_431 (O_431,N_2955,N_2963);
xnor UO_432 (O_432,N_2998,N_2969);
nor UO_433 (O_433,N_2987,N_2959);
nand UO_434 (O_434,N_2974,N_2999);
nand UO_435 (O_435,N_2974,N_2965);
nor UO_436 (O_436,N_2995,N_2971);
nand UO_437 (O_437,N_2992,N_2978);
xnor UO_438 (O_438,N_2982,N_2987);
nor UO_439 (O_439,N_2989,N_2972);
and UO_440 (O_440,N_2953,N_2977);
nand UO_441 (O_441,N_2998,N_2972);
or UO_442 (O_442,N_2979,N_2966);
or UO_443 (O_443,N_2974,N_2959);
nor UO_444 (O_444,N_2998,N_2978);
and UO_445 (O_445,N_2991,N_2942);
xnor UO_446 (O_446,N_2987,N_2944);
nand UO_447 (O_447,N_2995,N_2982);
nor UO_448 (O_448,N_2999,N_2976);
nor UO_449 (O_449,N_2952,N_2994);
or UO_450 (O_450,N_2974,N_2941);
nand UO_451 (O_451,N_2944,N_2960);
and UO_452 (O_452,N_2960,N_2991);
or UO_453 (O_453,N_2965,N_2972);
nand UO_454 (O_454,N_2953,N_2987);
or UO_455 (O_455,N_2950,N_2989);
nor UO_456 (O_456,N_2978,N_2951);
nor UO_457 (O_457,N_2952,N_2982);
nor UO_458 (O_458,N_2974,N_2955);
xnor UO_459 (O_459,N_2998,N_2953);
nor UO_460 (O_460,N_2988,N_2966);
xor UO_461 (O_461,N_2984,N_2959);
or UO_462 (O_462,N_2955,N_2968);
xnor UO_463 (O_463,N_2967,N_2963);
and UO_464 (O_464,N_2949,N_2960);
xnor UO_465 (O_465,N_2985,N_2962);
nor UO_466 (O_466,N_2947,N_2994);
and UO_467 (O_467,N_2964,N_2990);
xnor UO_468 (O_468,N_2979,N_2946);
nor UO_469 (O_469,N_2982,N_2969);
nor UO_470 (O_470,N_2985,N_2977);
nand UO_471 (O_471,N_2963,N_2981);
or UO_472 (O_472,N_2961,N_2995);
or UO_473 (O_473,N_2975,N_2984);
or UO_474 (O_474,N_2974,N_2995);
nand UO_475 (O_475,N_2977,N_2990);
nand UO_476 (O_476,N_2997,N_2982);
nor UO_477 (O_477,N_2996,N_2963);
nand UO_478 (O_478,N_2974,N_2951);
nor UO_479 (O_479,N_2982,N_2967);
xor UO_480 (O_480,N_2985,N_2946);
nand UO_481 (O_481,N_2969,N_2949);
xnor UO_482 (O_482,N_2944,N_2940);
xor UO_483 (O_483,N_2962,N_2983);
nand UO_484 (O_484,N_2979,N_2981);
or UO_485 (O_485,N_2973,N_2992);
nor UO_486 (O_486,N_2969,N_2954);
nand UO_487 (O_487,N_2947,N_2956);
xnor UO_488 (O_488,N_2995,N_2969);
and UO_489 (O_489,N_2989,N_2946);
and UO_490 (O_490,N_2973,N_2941);
or UO_491 (O_491,N_2957,N_2992);
or UO_492 (O_492,N_2940,N_2999);
nor UO_493 (O_493,N_2973,N_2958);
xnor UO_494 (O_494,N_2964,N_2971);
xor UO_495 (O_495,N_2953,N_2962);
or UO_496 (O_496,N_2978,N_2999);
nand UO_497 (O_497,N_2962,N_2996);
or UO_498 (O_498,N_2966,N_2954);
nand UO_499 (O_499,N_2951,N_2949);
endmodule