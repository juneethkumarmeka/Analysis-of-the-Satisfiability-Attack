module basic_1000_10000_1500_2_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5002,N_5003,N_5005,N_5006,N_5007,N_5008,N_5010,N_5011,N_5012,N_5013,N_5014,N_5016,N_5017,N_5018,N_5019,N_5021,N_5025,N_5026,N_5027,N_5029,N_5032,N_5033,N_5034,N_5037,N_5039,N_5040,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5052,N_5054,N_5056,N_5058,N_5059,N_5060,N_5062,N_5065,N_5067,N_5068,N_5073,N_5076,N_5078,N_5080,N_5084,N_5085,N_5087,N_5091,N_5096,N_5098,N_5100,N_5101,N_5102,N_5103,N_5106,N_5108,N_5109,N_5113,N_5115,N_5117,N_5118,N_5119,N_5121,N_5123,N_5124,N_5125,N_5127,N_5129,N_5130,N_5134,N_5138,N_5139,N_5143,N_5145,N_5147,N_5148,N_5149,N_5150,N_5152,N_5153,N_5154,N_5155,N_5157,N_5158,N_5159,N_5161,N_5162,N_5164,N_5165,N_5166,N_5167,N_5169,N_5170,N_5172,N_5173,N_5176,N_5177,N_5179,N_5180,N_5181,N_5183,N_5185,N_5186,N_5187,N_5189,N_5190,N_5193,N_5195,N_5196,N_5198,N_5199,N_5200,N_5202,N_5203,N_5204,N_5209,N_5211,N_5213,N_5214,N_5216,N_5217,N_5219,N_5221,N_5223,N_5224,N_5225,N_5226,N_5229,N_5231,N_5234,N_5236,N_5237,N_5238,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5250,N_5252,N_5254,N_5255,N_5256,N_5263,N_5265,N_5269,N_5270,N_5271,N_5272,N_5273,N_5277,N_5278,N_5279,N_5281,N_5282,N_5283,N_5284,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5294,N_5296,N_5297,N_5298,N_5299,N_5303,N_5304,N_5306,N_5307,N_5308,N_5309,N_5310,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5321,N_5325,N_5326,N_5327,N_5330,N_5331,N_5334,N_5335,N_5336,N_5337,N_5339,N_5340,N_5342,N_5343,N_5345,N_5346,N_5347,N_5348,N_5351,N_5352,N_5353,N_5355,N_5356,N_5357,N_5359,N_5360,N_5361,N_5362,N_5364,N_5365,N_5368,N_5369,N_5370,N_5371,N_5374,N_5375,N_5376,N_5377,N_5379,N_5382,N_5383,N_5385,N_5386,N_5387,N_5388,N_5391,N_5392,N_5396,N_5398,N_5399,N_5400,N_5402,N_5403,N_5404,N_5405,N_5407,N_5409,N_5412,N_5414,N_5415,N_5416,N_5417,N_5418,N_5421,N_5425,N_5426,N_5436,N_5437,N_5439,N_5443,N_5444,N_5446,N_5447,N_5448,N_5449,N_5451,N_5452,N_5453,N_5455,N_5456,N_5457,N_5463,N_5465,N_5466,N_5467,N_5468,N_5470,N_5471,N_5472,N_5473,N_5476,N_5483,N_5491,N_5492,N_5493,N_5495,N_5496,N_5497,N_5498,N_5500,N_5503,N_5505,N_5506,N_5508,N_5509,N_5510,N_5511,N_5513,N_5514,N_5515,N_5516,N_5518,N_5519,N_5520,N_5521,N_5525,N_5527,N_5528,N_5530,N_5532,N_5533,N_5534,N_5535,N_5536,N_5539,N_5541,N_5542,N_5543,N_5545,N_5547,N_5548,N_5549,N_5552,N_5554,N_5558,N_5560,N_5561,N_5562,N_5564,N_5565,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5576,N_5577,N_5578,N_5582,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5596,N_5599,N_5600,N_5602,N_5604,N_5605,N_5607,N_5608,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5620,N_5624,N_5625,N_5627,N_5630,N_5631,N_5632,N_5634,N_5637,N_5639,N_5640,N_5641,N_5642,N_5643,N_5645,N_5646,N_5651,N_5652,N_5653,N_5656,N_5659,N_5663,N_5664,N_5665,N_5666,N_5672,N_5675,N_5676,N_5678,N_5679,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5689,N_5692,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5702,N_5704,N_5705,N_5706,N_5709,N_5710,N_5713,N_5716,N_5717,N_5719,N_5720,N_5722,N_5723,N_5725,N_5726,N_5727,N_5728,N_5733,N_5734,N_5735,N_5737,N_5738,N_5739,N_5741,N_5742,N_5743,N_5747,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5760,N_5761,N_5762,N_5766,N_5767,N_5768,N_5769,N_5770,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5797,N_5799,N_5800,N_5802,N_5805,N_5806,N_5807,N_5810,N_5811,N_5812,N_5814,N_5815,N_5816,N_5817,N_5821,N_5822,N_5824,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5835,N_5836,N_5838,N_5839,N_5840,N_5843,N_5844,N_5846,N_5847,N_5848,N_5850,N_5852,N_5853,N_5856,N_5857,N_5860,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5872,N_5873,N_5875,N_5876,N_5877,N_5880,N_5882,N_5883,N_5885,N_5886,N_5888,N_5889,N_5890,N_5892,N_5893,N_5895,N_5896,N_5900,N_5901,N_5904,N_5905,N_5906,N_5909,N_5911,N_5912,N_5914,N_5915,N_5916,N_5919,N_5920,N_5921,N_5922,N_5923,N_5925,N_5926,N_5928,N_5929,N_5931,N_5933,N_5936,N_5938,N_5942,N_5945,N_5946,N_5947,N_5951,N_5952,N_5953,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5962,N_5963,N_5964,N_5965,N_5966,N_5969,N_5970,N_5972,N_5974,N_5976,N_5978,N_5981,N_5987,N_5988,N_5989,N_5991,N_5994,N_5997,N_5998,N_5999,N_6000,N_6005,N_6006,N_6008,N_6010,N_6014,N_6015,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6024,N_6025,N_6026,N_6028,N_6030,N_6032,N_6033,N_6037,N_6039,N_6043,N_6044,N_6045,N_6052,N_6054,N_6055,N_6056,N_6057,N_6059,N_6060,N_6061,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6071,N_6074,N_6075,N_6076,N_6078,N_6080,N_6082,N_6083,N_6084,N_6087,N_6088,N_6089,N_6090,N_6091,N_6094,N_6095,N_6096,N_6097,N_6100,N_6101,N_6102,N_6103,N_6104,N_6106,N_6107,N_6108,N_6111,N_6112,N_6113,N_6114,N_6116,N_6118,N_6119,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6132,N_6133,N_6135,N_6136,N_6140,N_6142,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6159,N_6160,N_6162,N_6164,N_6168,N_6170,N_6171,N_6174,N_6175,N_6176,N_6177,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6188,N_6189,N_6190,N_6195,N_6196,N_6197,N_6201,N_6202,N_6203,N_6204,N_6205,N_6209,N_6211,N_6213,N_6214,N_6215,N_6218,N_6220,N_6221,N_6222,N_6224,N_6225,N_6227,N_6228,N_6229,N_6230,N_6232,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6245,N_6246,N_6248,N_6249,N_6250,N_6254,N_6255,N_6256,N_6257,N_6258,N_6260,N_6263,N_6265,N_6266,N_6269,N_6271,N_6272,N_6273,N_6275,N_6277,N_6279,N_6280,N_6282,N_6285,N_6286,N_6296,N_6298,N_6303,N_6304,N_6305,N_6306,N_6308,N_6309,N_6314,N_6315,N_6316,N_6319,N_6321,N_6322,N_6324,N_6325,N_6326,N_6328,N_6329,N_6330,N_6333,N_6334,N_6336,N_6337,N_6340,N_6341,N_6342,N_6343,N_6347,N_6348,N_6351,N_6352,N_6355,N_6356,N_6358,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6381,N_6385,N_6386,N_6387,N_6388,N_6389,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6399,N_6402,N_6404,N_6405,N_6406,N_6407,N_6408,N_6412,N_6414,N_6415,N_6416,N_6419,N_6422,N_6424,N_6426,N_6428,N_6429,N_6431,N_6432,N_6433,N_6434,N_6436,N_6437,N_6440,N_6441,N_6442,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6454,N_6456,N_6457,N_6459,N_6462,N_6463,N_6464,N_6465,N_6467,N_6470,N_6471,N_6473,N_6474,N_6478,N_6479,N_6481,N_6483,N_6484,N_6485,N_6486,N_6487,N_6489,N_6490,N_6493,N_6494,N_6495,N_6496,N_6497,N_6499,N_6502,N_6503,N_6504,N_6505,N_6506,N_6508,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6518,N_6519,N_6524,N_6525,N_6527,N_6528,N_6531,N_6535,N_6536,N_6537,N_6539,N_6541,N_6543,N_6544,N_6545,N_6547,N_6549,N_6552,N_6553,N_6554,N_6556,N_6557,N_6561,N_6562,N_6563,N_6564,N_6566,N_6567,N_6569,N_6571,N_6573,N_6574,N_6578,N_6579,N_6581,N_6583,N_6584,N_6587,N_6589,N_6592,N_6596,N_6597,N_6598,N_6602,N_6604,N_6605,N_6606,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6617,N_6618,N_6621,N_6622,N_6624,N_6627,N_6631,N_6632,N_6634,N_6637,N_6638,N_6639,N_6640,N_6645,N_6647,N_6648,N_6649,N_6650,N_6651,N_6653,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6666,N_6668,N_6669,N_6670,N_6671,N_6673,N_6675,N_6676,N_6677,N_6679,N_6681,N_6685,N_6686,N_6687,N_6690,N_6691,N_6692,N_6694,N_6695,N_6696,N_6697,N_6702,N_6705,N_6706,N_6707,N_6709,N_6710,N_6714,N_6715,N_6718,N_6719,N_6724,N_6725,N_6729,N_6731,N_6732,N_6734,N_6737,N_6740,N_6741,N_6742,N_6743,N_6744,N_6746,N_6748,N_6749,N_6750,N_6752,N_6753,N_6754,N_6757,N_6759,N_6760,N_6761,N_6762,N_6765,N_6767,N_6768,N_6771,N_6772,N_6773,N_6775,N_6781,N_6782,N_6783,N_6784,N_6785,N_6788,N_6789,N_6790,N_6791,N_6792,N_6794,N_6796,N_6797,N_6801,N_6805,N_6806,N_6807,N_6812,N_6814,N_6816,N_6817,N_6819,N_6821,N_6823,N_6824,N_6826,N_6827,N_6828,N_6830,N_6833,N_6834,N_6835,N_6836,N_6837,N_6839,N_6842,N_6843,N_6846,N_6847,N_6848,N_6849,N_6853,N_6854,N_6856,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6868,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6881,N_6882,N_6883,N_6885,N_6888,N_6889,N_6890,N_6891,N_6892,N_6894,N_6896,N_6897,N_6900,N_6901,N_6902,N_6904,N_6906,N_6908,N_6909,N_6912,N_6913,N_6914,N_6916,N_6919,N_6920,N_6921,N_6924,N_6925,N_6926,N_6927,N_6930,N_6932,N_6933,N_6935,N_6936,N_6937,N_6938,N_6941,N_6942,N_6946,N_6947,N_6948,N_6950,N_6951,N_6952,N_6953,N_6955,N_6956,N_6958,N_6960,N_6961,N_6963,N_6964,N_6965,N_6966,N_6967,N_6969,N_6970,N_6972,N_6973,N_6974,N_6976,N_6977,N_6978,N_6979,N_6980,N_6984,N_6986,N_6987,N_6988,N_6989,N_6991,N_6992,N_6993,N_6995,N_6996,N_6997,N_6998,N_7000,N_7001,N_7002,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7021,N_7022,N_7023,N_7025,N_7026,N_7029,N_7031,N_7033,N_7034,N_7035,N_7043,N_7044,N_7045,N_7046,N_7048,N_7050,N_7052,N_7054,N_7055,N_7057,N_7058,N_7059,N_7060,N_7063,N_7064,N_7067,N_7068,N_7069,N_7070,N_7072,N_7073,N_7075,N_7077,N_7079,N_7080,N_7083,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7095,N_7096,N_7097,N_7098,N_7101,N_7103,N_7104,N_7105,N_7107,N_7110,N_7114,N_7119,N_7124,N_7126,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7140,N_7142,N_7144,N_7145,N_7146,N_7147,N_7148,N_7150,N_7152,N_7154,N_7155,N_7156,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7173,N_7174,N_7178,N_7179,N_7181,N_7182,N_7183,N_7184,N_7185,N_7188,N_7189,N_7190,N_7191,N_7194,N_7195,N_7196,N_7197,N_7198,N_7202,N_7203,N_7205,N_7207,N_7209,N_7210,N_7211,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7221,N_7225,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7235,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7246,N_7247,N_7249,N_7256,N_7258,N_7259,N_7263,N_7264,N_7265,N_7267,N_7268,N_7269,N_7271,N_7272,N_7274,N_7277,N_7278,N_7279,N_7280,N_7281,N_7284,N_7287,N_7289,N_7291,N_7293,N_7294,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7306,N_7307,N_7310,N_7315,N_7316,N_7321,N_7324,N_7326,N_7330,N_7333,N_7335,N_7336,N_7338,N_7339,N_7342,N_7343,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7352,N_7353,N_7356,N_7358,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7376,N_7378,N_7379,N_7380,N_7382,N_7383,N_7385,N_7386,N_7387,N_7388,N_7390,N_7391,N_7392,N_7393,N_7395,N_7397,N_7399,N_7400,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7410,N_7411,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7424,N_7426,N_7427,N_7428,N_7429,N_7431,N_7433,N_7434,N_7436,N_7438,N_7440,N_7441,N_7442,N_7443,N_7444,N_7446,N_7447,N_7448,N_7450,N_7451,N_7452,N_7453,N_7454,N_7456,N_7457,N_7458,N_7460,N_7461,N_7462,N_7464,N_7465,N_7466,N_7467,N_7469,N_7470,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7483,N_7485,N_7486,N_7488,N_7489,N_7490,N_7491,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7501,N_7505,N_7506,N_7513,N_7519,N_7521,N_7524,N_7526,N_7527,N_7529,N_7532,N_7533,N_7534,N_7537,N_7538,N_7539,N_7541,N_7542,N_7543,N_7546,N_7548,N_7549,N_7553,N_7554,N_7556,N_7560,N_7561,N_7562,N_7563,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7578,N_7579,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7597,N_7598,N_7600,N_7602,N_7605,N_7606,N_7607,N_7608,N_7609,N_7612,N_7613,N_7614,N_7615,N_7616,N_7620,N_7621,N_7622,N_7623,N_7624,N_7626,N_7629,N_7635,N_7636,N_7637,N_7640,N_7643,N_7645,N_7646,N_7649,N_7650,N_7651,N_7652,N_7653,N_7655,N_7656,N_7657,N_7659,N_7660,N_7664,N_7665,N_7667,N_7668,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7682,N_7683,N_7686,N_7691,N_7692,N_7693,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7705,N_7706,N_7707,N_7708,N_7712,N_7714,N_7715,N_7716,N_7717,N_7718,N_7724,N_7727,N_7729,N_7732,N_7733,N_7734,N_7738,N_7739,N_7740,N_7741,N_7742,N_7745,N_7746,N_7748,N_7749,N_7750,N_7753,N_7754,N_7755,N_7757,N_7758,N_7761,N_7764,N_7766,N_7769,N_7770,N_7772,N_7773,N_7774,N_7776,N_7777,N_7779,N_7780,N_7782,N_7787,N_7788,N_7789,N_7790,N_7792,N_7796,N_7798,N_7799,N_7801,N_7802,N_7803,N_7804,N_7806,N_7808,N_7809,N_7811,N_7814,N_7816,N_7817,N_7818,N_7820,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7829,N_7830,N_7832,N_7833,N_7834,N_7839,N_7841,N_7842,N_7843,N_7844,N_7847,N_7852,N_7854,N_7855,N_7857,N_7858,N_7859,N_7862,N_7863,N_7864,N_7865,N_7868,N_7873,N_7879,N_7880,N_7882,N_7883,N_7884,N_7886,N_7887,N_7888,N_7889,N_7891,N_7892,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7901,N_7903,N_7904,N_7908,N_7909,N_7911,N_7912,N_7913,N_7915,N_7916,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7928,N_7929,N_7931,N_7932,N_7933,N_7934,N_7935,N_7937,N_7939,N_7940,N_7941,N_7942,N_7943,N_7945,N_7946,N_7948,N_7951,N_7952,N_7953,N_7954,N_7955,N_7958,N_7959,N_7961,N_7965,N_7966,N_7968,N_7970,N_7971,N_7973,N_7974,N_7975,N_7976,N_7977,N_7979,N_7981,N_7982,N_7984,N_7985,N_7993,N_7994,N_7997,N_7998,N_8000,N_8001,N_8003,N_8004,N_8009,N_8011,N_8012,N_8013,N_8015,N_8016,N_8020,N_8022,N_8024,N_8027,N_8029,N_8032,N_8037,N_8038,N_8039,N_8041,N_8045,N_8046,N_8047,N_8049,N_8050,N_8054,N_8055,N_8056,N_8057,N_8059,N_8060,N_8061,N_8062,N_8064,N_8065,N_8070,N_8072,N_8074,N_8076,N_8077,N_8078,N_8080,N_8083,N_8085,N_8086,N_8089,N_8091,N_8093,N_8094,N_8095,N_8097,N_8099,N_8101,N_8104,N_8105,N_8106,N_8107,N_8108,N_8110,N_8111,N_8113,N_8116,N_8117,N_8119,N_8121,N_8127,N_8131,N_8132,N_8133,N_8136,N_8137,N_8138,N_8140,N_8143,N_8144,N_8145,N_8148,N_8149,N_8150,N_8151,N_8153,N_8158,N_8159,N_8160,N_8166,N_8167,N_8169,N_8170,N_8172,N_8173,N_8176,N_8177,N_8178,N_8179,N_8182,N_8183,N_8184,N_8186,N_8187,N_8189,N_8190,N_8192,N_8193,N_8194,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8203,N_8204,N_8207,N_8208,N_8209,N_8210,N_8212,N_8213,N_8215,N_8216,N_8219,N_8220,N_8221,N_8222,N_8224,N_8225,N_8226,N_8227,N_8229,N_8230,N_8231,N_8234,N_8236,N_8239,N_8240,N_8241,N_8247,N_8248,N_8251,N_8252,N_8254,N_8255,N_8256,N_8257,N_8261,N_8262,N_8265,N_8267,N_8269,N_8271,N_8272,N_8277,N_8278,N_8279,N_8280,N_8285,N_8286,N_8288,N_8291,N_8293,N_8296,N_8297,N_8298,N_8299,N_8301,N_8302,N_8306,N_8307,N_8308,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8323,N_8324,N_8328,N_8329,N_8330,N_8331,N_8332,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8344,N_8345,N_8347,N_8351,N_8352,N_8356,N_8358,N_8360,N_8362,N_8364,N_8365,N_8366,N_8367,N_8374,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8383,N_8385,N_8387,N_8389,N_8392,N_8395,N_8397,N_8399,N_8400,N_8401,N_8402,N_8403,N_8406,N_8407,N_8408,N_8410,N_8411,N_8412,N_8413,N_8414,N_8416,N_8418,N_8419,N_8420,N_8421,N_8422,N_8424,N_8425,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8438,N_8440,N_8442,N_8443,N_8444,N_8445,N_8446,N_8449,N_8450,N_8452,N_8453,N_8454,N_8457,N_8459,N_8460,N_8461,N_8465,N_8466,N_8469,N_8470,N_8472,N_8477,N_8478,N_8479,N_8480,N_8482,N_8483,N_8484,N_8486,N_8487,N_8488,N_8490,N_8491,N_8492,N_8495,N_8496,N_8499,N_8505,N_8507,N_8508,N_8509,N_8510,N_8511,N_8513,N_8514,N_8515,N_8516,N_8517,N_8519,N_8520,N_8521,N_8522,N_8524,N_8525,N_8527,N_8530,N_8534,N_8535,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8547,N_8548,N_8549,N_8552,N_8553,N_8554,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8569,N_8570,N_8572,N_8573,N_8574,N_8575,N_8577,N_8580,N_8582,N_8583,N_8584,N_8585,N_8588,N_8589,N_8590,N_8591,N_8594,N_8596,N_8597,N_8598,N_8599,N_8602,N_8603,N_8604,N_8605,N_8607,N_8609,N_8611,N_8612,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8640,N_8644,N_8645,N_8647,N_8648,N_8649,N_8653,N_8654,N_8657,N_8659,N_8661,N_8663,N_8664,N_8667,N_8669,N_8673,N_8674,N_8677,N_8679,N_8681,N_8683,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8697,N_8698,N_8699,N_8700,N_8701,N_8703,N_8704,N_8705,N_8706,N_8707,N_8709,N_8710,N_8712,N_8714,N_8715,N_8716,N_8717,N_8719,N_8720,N_8721,N_8722,N_8723,N_8726,N_8727,N_8729,N_8731,N_8732,N_8733,N_8734,N_8737,N_8741,N_8742,N_8743,N_8744,N_8745,N_8747,N_8748,N_8749,N_8750,N_8754,N_8756,N_8757,N_8758,N_8759,N_8761,N_8762,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8775,N_8776,N_8778,N_8779,N_8780,N_8785,N_8786,N_8787,N_8788,N_8789,N_8791,N_8792,N_8794,N_8798,N_8800,N_8801,N_8803,N_8804,N_8806,N_8807,N_8810,N_8811,N_8812,N_8814,N_8815,N_8816,N_8817,N_8820,N_8821,N_8822,N_8823,N_8824,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8838,N_8840,N_8843,N_8846,N_8847,N_8848,N_8851,N_8857,N_8859,N_8860,N_8862,N_8863,N_8865,N_8866,N_8867,N_8870,N_8872,N_8876,N_8877,N_8878,N_8880,N_8881,N_8884,N_8885,N_8886,N_8887,N_8888,N_8890,N_8891,N_8892,N_8894,N_8895,N_8896,N_8897,N_8902,N_8903,N_8904,N_8906,N_8908,N_8909,N_8910,N_8912,N_8913,N_8914,N_8916,N_8921,N_8922,N_8924,N_8926,N_8927,N_8929,N_8931,N_8933,N_8936,N_8937,N_8939,N_8940,N_8942,N_8943,N_8946,N_8949,N_8950,N_8951,N_8953,N_8954,N_8956,N_8957,N_8958,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8969,N_8971,N_8972,N_8973,N_8975,N_8978,N_8982,N_8984,N_8985,N_8987,N_8989,N_8990,N_8993,N_8994,N_8995,N_8996,N_8997,N_8999,N_9004,N_9005,N_9006,N_9007,N_9008,N_9011,N_9013,N_9014,N_9015,N_9017,N_9018,N_9019,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9029,N_9030,N_9031,N_9036,N_9037,N_9041,N_9042,N_9045,N_9048,N_9049,N_9050,N_9052,N_9053,N_9057,N_9059,N_9060,N_9062,N_9064,N_9065,N_9067,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9079,N_9080,N_9081,N_9084,N_9085,N_9086,N_9087,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9100,N_9101,N_9102,N_9103,N_9105,N_9108,N_9109,N_9111,N_9112,N_9113,N_9116,N_9118,N_9119,N_9120,N_9122,N_9123,N_9127,N_9130,N_9131,N_9132,N_9134,N_9135,N_9137,N_9139,N_9140,N_9142,N_9143,N_9145,N_9146,N_9147,N_9148,N_9150,N_9153,N_9156,N_9157,N_9158,N_9160,N_9162,N_9164,N_9165,N_9168,N_9169,N_9173,N_9174,N_9175,N_9177,N_9179,N_9180,N_9181,N_9184,N_9185,N_9188,N_9192,N_9196,N_9198,N_9199,N_9200,N_9201,N_9202,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9213,N_9216,N_9217,N_9219,N_9220,N_9222,N_9223,N_9224,N_9225,N_9226,N_9228,N_9231,N_9234,N_9238,N_9240,N_9242,N_9243,N_9246,N_9247,N_9253,N_9256,N_9257,N_9258,N_9259,N_9261,N_9262,N_9264,N_9266,N_9267,N_9268,N_9269,N_9273,N_9274,N_9275,N_9278,N_9280,N_9284,N_9285,N_9286,N_9287,N_9288,N_9290,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9301,N_9302,N_9303,N_9304,N_9305,N_9307,N_9309,N_9310,N_9311,N_9312,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9326,N_9328,N_9329,N_9330,N_9331,N_9333,N_9334,N_9335,N_9336,N_9339,N_9340,N_9342,N_9343,N_9346,N_9348,N_9349,N_9351,N_9352,N_9353,N_9354,N_9355,N_9357,N_9358,N_9363,N_9364,N_9365,N_9366,N_9367,N_9369,N_9371,N_9373,N_9375,N_9377,N_9378,N_9379,N_9381,N_9383,N_9384,N_9385,N_9386,N_9388,N_9389,N_9391,N_9392,N_9394,N_9396,N_9397,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9408,N_9409,N_9414,N_9415,N_9416,N_9417,N_9418,N_9420,N_9422,N_9423,N_9426,N_9429,N_9430,N_9433,N_9434,N_9435,N_9437,N_9438,N_9440,N_9441,N_9442,N_9445,N_9447,N_9448,N_9450,N_9452,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9462,N_9464,N_9467,N_9471,N_9474,N_9475,N_9476,N_9478,N_9479,N_9480,N_9482,N_9485,N_9488,N_9489,N_9490,N_9493,N_9494,N_9495,N_9498,N_9500,N_9504,N_9506,N_9507,N_9508,N_9511,N_9513,N_9514,N_9515,N_9516,N_9519,N_9520,N_9521,N_9522,N_9523,N_9525,N_9526,N_9528,N_9529,N_9530,N_9532,N_9533,N_9536,N_9537,N_9538,N_9539,N_9541,N_9543,N_9545,N_9547,N_9549,N_9550,N_9552,N_9555,N_9556,N_9561,N_9562,N_9566,N_9567,N_9568,N_9569,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9578,N_9579,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9599,N_9604,N_9605,N_9606,N_9607,N_9608,N_9610,N_9612,N_9613,N_9615,N_9617,N_9619,N_9620,N_9622,N_9624,N_9625,N_9626,N_9628,N_9629,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9648,N_9649,N_9651,N_9652,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9661,N_9662,N_9663,N_9665,N_9666,N_9668,N_9670,N_9674,N_9677,N_9681,N_9682,N_9684,N_9685,N_9688,N_9689,N_9690,N_9691,N_9693,N_9698,N_9701,N_9702,N_9703,N_9704,N_9705,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9717,N_9718,N_9719,N_9722,N_9723,N_9729,N_9731,N_9732,N_9733,N_9734,N_9735,N_9739,N_9740,N_9741,N_9742,N_9744,N_9747,N_9748,N_9749,N_9751,N_9753,N_9755,N_9756,N_9758,N_9759,N_9760,N_9763,N_9764,N_9767,N_9768,N_9769,N_9770,N_9772,N_9773,N_9774,N_9775,N_9777,N_9779,N_9781,N_9783,N_9785,N_9789,N_9790,N_9792,N_9793,N_9795,N_9797,N_9798,N_9799,N_9800,N_9804,N_9805,N_9806,N_9810,N_9812,N_9814,N_9815,N_9818,N_9819,N_9820,N_9822,N_9823,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9834,N_9835,N_9836,N_9837,N_9839,N_9840,N_9843,N_9845,N_9846,N_9849,N_9850,N_9851,N_9852,N_9854,N_9857,N_9859,N_9860,N_9862,N_9863,N_9864,N_9865,N_9866,N_9868,N_9873,N_9874,N_9875,N_9877,N_9879,N_9880,N_9881,N_9883,N_9884,N_9885,N_9886,N_9888,N_9889,N_9890,N_9894,N_9895,N_9896,N_9897,N_9899,N_9901,N_9904,N_9906,N_9908,N_9909,N_9910,N_9912,N_9913,N_9914,N_9917,N_9918,N_9919,N_9920,N_9922,N_9923,N_9924,N_9925,N_9926,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9936,N_9937,N_9938,N_9940,N_9942,N_9944,N_9945,N_9947,N_9949,N_9952,N_9954,N_9955,N_9956,N_9958,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9971,N_9972,N_9974,N_9975,N_9977,N_9978,N_9979,N_9981,N_9982,N_9984,N_9988,N_9989,N_9990,N_9992,N_9993,N_9994,N_9995,N_9998;
and U0 (N_0,In_286,In_275);
nor U1 (N_1,In_955,In_942);
nor U2 (N_2,In_480,In_361);
and U3 (N_3,In_358,In_193);
or U4 (N_4,In_490,In_717);
nand U5 (N_5,In_157,In_887);
nor U6 (N_6,In_300,In_336);
nand U7 (N_7,In_702,In_243);
or U8 (N_8,In_20,In_73);
or U9 (N_9,In_0,In_134);
xor U10 (N_10,In_640,In_291);
xnor U11 (N_11,In_927,In_666);
nor U12 (N_12,In_914,In_109);
and U13 (N_13,In_888,In_372);
or U14 (N_14,In_11,In_45);
xor U15 (N_15,In_630,In_209);
xor U16 (N_16,In_428,In_186);
nand U17 (N_17,In_341,In_941);
nor U18 (N_18,In_738,In_346);
nand U19 (N_19,In_660,In_279);
xnor U20 (N_20,In_687,In_535);
xnor U21 (N_21,In_858,In_135);
and U22 (N_22,In_443,In_735);
nor U23 (N_23,In_661,In_68);
or U24 (N_24,In_655,In_552);
nor U25 (N_25,In_442,In_620);
and U26 (N_26,In_69,In_445);
xnor U27 (N_27,In_67,In_161);
or U28 (N_28,In_387,In_618);
nand U29 (N_29,In_409,In_250);
or U30 (N_30,In_893,In_196);
nor U31 (N_31,In_197,In_78);
or U32 (N_32,In_897,In_921);
nand U33 (N_33,In_939,In_844);
nor U34 (N_34,In_945,In_802);
nor U35 (N_35,In_534,In_904);
nand U36 (N_36,In_987,In_83);
nand U37 (N_37,In_288,In_784);
nand U38 (N_38,In_555,In_16);
or U39 (N_39,In_65,In_453);
and U40 (N_40,In_369,In_347);
and U41 (N_41,In_155,In_416);
nor U42 (N_42,In_616,In_648);
xnor U43 (N_43,In_800,In_406);
nor U44 (N_44,In_184,In_837);
and U45 (N_45,In_169,In_145);
nor U46 (N_46,In_342,In_228);
and U47 (N_47,In_632,In_707);
nand U48 (N_48,In_567,In_441);
nand U49 (N_49,In_494,In_107);
nor U50 (N_50,In_973,In_895);
nor U51 (N_51,In_561,In_192);
or U52 (N_52,In_482,In_518);
xnor U53 (N_53,In_423,In_515);
nor U54 (N_54,In_556,In_175);
or U55 (N_55,In_14,In_875);
nand U56 (N_56,In_407,In_321);
or U57 (N_57,In_664,In_812);
nor U58 (N_58,In_230,In_103);
xnor U59 (N_59,In_586,In_225);
nand U60 (N_60,In_662,In_131);
nor U61 (N_61,In_191,In_512);
xnor U62 (N_62,In_79,In_199);
or U63 (N_63,In_591,In_201);
or U64 (N_64,In_801,In_594);
nand U65 (N_65,In_479,In_990);
xor U66 (N_66,In_373,In_469);
nand U67 (N_67,In_88,In_302);
xor U68 (N_68,In_468,In_345);
and U69 (N_69,In_823,In_422);
xor U70 (N_70,In_628,In_141);
nand U71 (N_71,In_6,In_439);
and U72 (N_72,In_557,In_349);
or U73 (N_73,In_639,In_375);
nor U74 (N_74,In_313,In_585);
xnor U75 (N_75,In_524,In_128);
xnor U76 (N_76,In_502,In_23);
xnor U77 (N_77,In_37,In_357);
nor U78 (N_78,In_674,In_19);
nor U79 (N_79,In_467,In_545);
nand U80 (N_80,In_762,In_785);
nor U81 (N_81,In_968,In_722);
nor U82 (N_82,In_562,In_280);
and U83 (N_83,In_36,In_158);
nand U84 (N_84,In_98,In_590);
nor U85 (N_85,In_381,In_755);
and U86 (N_86,In_473,In_581);
or U87 (N_87,In_143,In_380);
nand U88 (N_88,In_260,In_690);
and U89 (N_89,In_262,In_343);
xor U90 (N_90,In_621,In_991);
nand U91 (N_91,In_181,In_398);
nand U92 (N_92,In_7,In_388);
nand U93 (N_93,In_334,In_274);
nand U94 (N_94,In_124,In_351);
xor U95 (N_95,In_610,In_237);
xnor U96 (N_96,In_241,In_127);
or U97 (N_97,In_878,In_960);
nand U98 (N_98,In_865,In_2);
or U99 (N_99,In_712,In_852);
nor U100 (N_100,In_356,In_438);
xor U101 (N_101,In_133,In_91);
nor U102 (N_102,In_763,In_958);
nand U103 (N_103,In_56,In_99);
nor U104 (N_104,In_781,In_456);
xor U105 (N_105,In_101,In_170);
nand U106 (N_106,In_983,In_10);
and U107 (N_107,In_910,In_956);
and U108 (N_108,In_394,In_319);
nand U109 (N_109,In_836,In_706);
nor U110 (N_110,In_203,In_753);
xor U111 (N_111,In_283,In_601);
nand U112 (N_112,In_675,In_129);
or U113 (N_113,In_337,In_360);
xor U114 (N_114,In_385,In_495);
and U115 (N_115,In_726,In_139);
nor U116 (N_116,In_376,In_70);
nand U117 (N_117,In_460,In_885);
xor U118 (N_118,In_164,In_348);
or U119 (N_119,In_177,In_588);
or U120 (N_120,In_154,In_234);
nand U121 (N_121,In_259,In_327);
xor U122 (N_122,In_732,In_806);
and U123 (N_123,In_115,In_148);
nor U124 (N_124,In_111,In_344);
nand U125 (N_125,In_948,In_805);
nor U126 (N_126,In_391,In_47);
or U127 (N_127,In_435,In_108);
nor U128 (N_128,In_908,In_807);
nand U129 (N_129,In_365,In_304);
and U130 (N_130,In_913,In_57);
or U131 (N_131,In_672,In_13);
or U132 (N_132,In_957,In_924);
nand U133 (N_133,In_481,In_838);
and U134 (N_134,In_764,In_476);
nor U135 (N_135,In_720,In_613);
nand U136 (N_136,In_450,In_740);
nor U137 (N_137,In_508,In_163);
and U138 (N_138,In_174,In_403);
nand U139 (N_139,In_268,In_694);
xnor U140 (N_140,In_151,In_754);
nand U141 (N_141,In_724,In_41);
and U142 (N_142,In_827,In_959);
and U143 (N_143,In_411,In_117);
and U144 (N_144,In_452,In_35);
or U145 (N_145,In_570,In_950);
and U146 (N_146,In_606,In_658);
nand U147 (N_147,In_751,In_371);
or U148 (N_148,In_206,In_217);
and U149 (N_149,In_821,In_95);
and U150 (N_150,In_529,In_454);
nand U151 (N_151,In_251,In_214);
or U152 (N_152,In_743,In_605);
nor U153 (N_153,In_253,In_22);
and U154 (N_154,In_305,In_267);
xor U155 (N_155,In_771,In_532);
xor U156 (N_156,In_565,In_121);
and U157 (N_157,In_572,In_287);
nor U158 (N_158,In_440,In_355);
and U159 (N_159,In_890,In_142);
nor U160 (N_160,In_190,In_848);
and U161 (N_161,In_860,In_77);
xnor U162 (N_162,In_389,In_316);
nor U163 (N_163,In_229,In_593);
xor U164 (N_164,In_841,In_528);
and U165 (N_165,In_52,In_278);
nand U166 (N_166,In_309,In_798);
xor U167 (N_167,In_988,In_410);
nand U168 (N_168,In_644,In_239);
and U169 (N_169,In_87,In_367);
xor U170 (N_170,In_659,In_102);
nor U171 (N_171,In_831,In_232);
nand U172 (N_172,In_140,In_937);
and U173 (N_173,In_49,In_150);
nor U174 (N_174,In_680,In_338);
or U175 (N_175,In_402,In_946);
nor U176 (N_176,In_270,In_944);
nor U177 (N_177,In_513,In_856);
nand U178 (N_178,In_136,In_213);
and U179 (N_179,In_76,In_627);
nand U180 (N_180,In_44,In_879);
nor U181 (N_181,In_202,In_951);
nor U182 (N_182,In_651,In_714);
or U183 (N_183,In_297,In_850);
nand U184 (N_184,In_589,In_30);
xnor U185 (N_185,In_679,In_668);
and U186 (N_186,In_8,In_779);
nor U187 (N_187,In_693,In_749);
and U188 (N_188,In_298,In_641);
nand U189 (N_189,In_900,In_855);
nand U190 (N_190,In_769,In_929);
xor U191 (N_191,In_501,In_113);
nand U192 (N_192,In_160,In_700);
and U193 (N_193,In_62,In_459);
or U194 (N_194,In_932,In_797);
xnor U195 (N_195,In_500,In_61);
nor U196 (N_196,In_293,In_211);
and U197 (N_197,In_851,In_713);
xor U198 (N_198,In_474,In_363);
or U199 (N_199,In_611,In_943);
or U200 (N_200,In_55,In_461);
nand U201 (N_201,In_974,In_81);
nand U202 (N_202,In_979,In_730);
xor U203 (N_203,In_840,In_725);
or U204 (N_204,In_218,In_105);
or U205 (N_205,In_835,In_153);
xor U206 (N_206,In_624,In_80);
and U207 (N_207,In_156,In_984);
xor U208 (N_208,In_208,In_971);
nor U209 (N_209,In_303,In_263);
nand U210 (N_210,In_727,In_825);
nor U211 (N_211,In_66,In_272);
xor U212 (N_212,In_82,In_434);
or U213 (N_213,In_692,In_284);
or U214 (N_214,In_965,In_324);
and U215 (N_215,In_162,In_379);
and U216 (N_216,In_326,In_466);
nor U217 (N_217,In_311,In_832);
and U218 (N_218,In_673,In_182);
xor U219 (N_219,In_881,In_993);
and U220 (N_220,In_992,In_701);
nand U221 (N_221,In_366,In_859);
and U222 (N_222,In_637,In_188);
nor U223 (N_223,In_339,In_359);
or U224 (N_224,In_905,In_166);
or U225 (N_225,In_332,In_401);
nand U226 (N_226,In_207,In_608);
xor U227 (N_227,In_533,In_446);
nor U228 (N_228,In_246,In_683);
and U229 (N_229,In_558,In_750);
xor U230 (N_230,In_216,In_235);
or U231 (N_231,In_273,In_396);
and U232 (N_232,In_809,In_455);
nor U233 (N_233,In_90,In_575);
nor U234 (N_234,In_966,In_677);
and U235 (N_235,In_27,In_537);
xor U236 (N_236,In_42,In_778);
nor U237 (N_237,In_180,In_982);
nor U238 (N_238,In_954,In_176);
nand U239 (N_239,In_195,In_547);
xnor U240 (N_240,In_104,In_144);
and U241 (N_241,In_231,In_866);
xor U242 (N_242,In_912,In_252);
nor U243 (N_243,In_475,In_978);
nand U244 (N_244,In_564,In_917);
nand U245 (N_245,In_498,In_292);
nor U246 (N_246,In_870,In_884);
and U247 (N_247,In_39,In_970);
and U248 (N_248,In_657,In_464);
nor U249 (N_249,In_514,In_808);
or U250 (N_250,In_421,In_447);
or U251 (N_251,In_1,In_472);
or U252 (N_252,In_775,In_554);
or U253 (N_253,In_744,In_503);
and U254 (N_254,In_695,In_519);
nand U255 (N_255,In_704,In_776);
nand U256 (N_256,In_418,In_486);
nand U257 (N_257,In_645,In_663);
nand U258 (N_258,In_696,In_931);
and U259 (N_259,In_597,In_863);
nand U260 (N_260,In_566,In_492);
xor U261 (N_261,In_697,In_861);
and U262 (N_262,In_483,In_625);
nand U263 (N_263,In_669,In_803);
nand U264 (N_264,In_891,In_489);
nor U265 (N_265,In_783,In_523);
nand U266 (N_266,In_854,In_215);
xor U267 (N_267,In_986,In_622);
nand U268 (N_268,In_643,In_236);
nor U269 (N_269,In_509,In_510);
nand U270 (N_270,In_811,In_431);
and U271 (N_271,In_839,In_609);
or U272 (N_272,In_934,In_340);
xor U273 (N_273,In_901,In_737);
or U274 (N_274,In_171,In_427);
xor U275 (N_275,In_352,In_204);
xor U276 (N_276,In_48,In_165);
or U277 (N_277,In_33,In_377);
nand U278 (N_278,In_617,In_777);
or U279 (N_279,In_289,In_71);
nand U280 (N_280,In_308,In_698);
or U281 (N_281,In_719,In_395);
and U282 (N_282,In_676,In_255);
nor U283 (N_283,In_742,In_652);
nand U284 (N_284,In_172,In_623);
nor U285 (N_285,In_918,In_462);
or U286 (N_286,In_59,In_43);
xnor U287 (N_287,In_147,In_770);
nand U288 (N_288,In_210,In_374);
nor U289 (N_289,In_224,In_963);
xnor U290 (N_290,In_782,In_846);
nor U291 (N_291,In_74,In_896);
and U292 (N_292,In_179,In_198);
xor U293 (N_293,In_412,In_767);
and U294 (N_294,In_364,In_146);
and U295 (N_295,In_185,In_889);
nor U296 (N_296,In_392,In_540);
nand U297 (N_297,In_768,In_953);
or U298 (N_298,In_223,In_996);
nand U299 (N_299,In_994,In_384);
or U300 (N_300,In_682,In_458);
nand U301 (N_301,In_686,In_488);
xor U302 (N_302,In_429,In_323);
xor U303 (N_303,In_245,In_84);
nor U304 (N_304,In_189,In_819);
and U305 (N_305,In_592,In_728);
nand U306 (N_306,In_386,In_168);
xor U307 (N_307,In_26,In_173);
nand U308 (N_308,In_969,In_869);
and U309 (N_309,In_595,In_650);
and U310 (N_310,In_862,In_600);
nand U311 (N_311,In_603,In_985);
nand U312 (N_312,In_187,In_578);
nand U313 (N_313,In_813,In_233);
or U314 (N_314,In_315,In_551);
and U315 (N_315,In_899,In_938);
nand U316 (N_316,In_322,In_546);
and U317 (N_317,In_525,In_817);
xnor U318 (N_318,In_933,In_200);
and U319 (N_319,In_583,In_829);
nand U320 (N_320,In_28,In_766);
nor U321 (N_321,In_419,In_997);
or U322 (N_322,In_867,In_282);
xnor U323 (N_323,In_906,In_85);
or U324 (N_324,In_898,In_178);
xor U325 (N_325,In_542,In_792);
nand U326 (N_326,In_925,In_4);
or U327 (N_327,In_656,In_574);
xor U328 (N_328,In_810,In_119);
xor U329 (N_329,In_607,In_559);
or U330 (N_330,In_935,In_312);
xor U331 (N_331,In_868,In_923);
or U332 (N_332,In_307,In_820);
and U333 (N_333,In_873,In_799);
nor U334 (N_334,In_612,In_484);
nor U335 (N_335,In_238,In_249);
nand U336 (N_336,In_746,In_15);
nor U337 (N_337,In_998,In_437);
and U338 (N_338,In_631,In_538);
or U339 (N_339,In_522,In_772);
nand U340 (N_340,In_794,In_444);
and U341 (N_341,In_125,In_417);
or U342 (N_342,In_100,In_505);
and U343 (N_343,In_667,In_212);
xnor U344 (N_344,In_399,In_705);
nand U345 (N_345,In_633,In_818);
nor U346 (N_346,In_977,In_451);
nand U347 (N_347,In_629,In_874);
or U348 (N_348,In_449,In_688);
nor U349 (N_349,In_353,In_110);
xor U350 (N_350,In_789,In_220);
or U351 (N_351,In_132,In_106);
nand U352 (N_352,In_40,In_50);
or U353 (N_353,In_487,In_734);
xnor U354 (N_354,In_828,In_247);
or U355 (N_355,In_759,In_795);
and U356 (N_356,In_75,In_244);
and U357 (N_357,In_788,In_814);
nand U358 (N_358,In_573,In_549);
or U359 (N_359,In_167,In_383);
xor U360 (N_360,In_415,In_425);
nor U361 (N_361,In_847,In_465);
nor U362 (N_362,In_122,In_86);
nand U363 (N_363,In_967,In_318);
and U364 (N_364,In_433,In_12);
or U365 (N_365,In_331,In_277);
nand U366 (N_366,In_853,In_635);
and U367 (N_367,In_834,In_568);
nor U368 (N_368,In_92,In_63);
nand U369 (N_369,In_715,In_457);
xor U370 (N_370,In_424,In_709);
and U371 (N_371,In_38,In_587);
xor U372 (N_372,In_504,In_93);
xor U373 (N_373,In_882,In_527);
and U374 (N_374,In_786,In_892);
nand U375 (N_375,In_400,In_584);
or U376 (N_376,In_646,In_582);
nand U377 (N_377,In_310,In_741);
nand U378 (N_378,In_29,In_947);
nor U379 (N_379,In_649,In_857);
and U380 (N_380,In_830,In_599);
and U381 (N_381,In_301,In_520);
and U382 (N_382,In_748,In_880);
and U383 (N_383,In_24,In_902);
nand U384 (N_384,In_149,In_773);
or U385 (N_385,In_408,In_485);
nor U386 (N_386,In_31,In_756);
and U387 (N_387,In_137,In_975);
and U388 (N_388,In_97,In_876);
nand U389 (N_389,In_816,In_670);
and U390 (N_390,In_493,In_94);
and U391 (N_391,In_261,In_264);
xor U392 (N_392,In_222,In_915);
or U393 (N_393,In_414,In_18);
nor U394 (N_394,In_295,In_114);
nor U395 (N_395,In_926,In_463);
and U396 (N_396,In_491,In_678);
nor U397 (N_397,In_580,In_496);
xnor U398 (N_398,In_711,In_320);
and U399 (N_399,In_362,In_708);
nand U400 (N_400,In_903,In_940);
or U401 (N_401,In_922,In_471);
nand U402 (N_402,In_265,In_511);
or U403 (N_403,In_886,In_329);
nand U404 (N_404,In_314,In_736);
or U405 (N_405,In_790,In_685);
xnor U406 (N_406,In_636,In_995);
nor U407 (N_407,In_699,In_120);
and U408 (N_408,In_89,In_21);
nand U409 (N_409,In_328,In_96);
xor U410 (N_410,In_413,In_571);
nand U411 (N_411,In_536,In_138);
nor U412 (N_412,In_521,In_647);
or U413 (N_413,In_723,In_248);
nor U414 (N_414,In_989,In_843);
nand U415 (N_415,In_325,In_526);
nor U416 (N_416,In_703,In_72);
nor U417 (N_417,In_949,In_370);
xor U418 (N_418,In_761,In_604);
nand U419 (N_419,In_689,In_553);
nor U420 (N_420,In_257,In_368);
nand U421 (N_421,In_930,In_826);
nor U422 (N_422,In_420,In_665);
and U423 (N_423,In_563,In_152);
and U424 (N_424,In_430,In_638);
xnor U425 (N_425,In_497,In_739);
and U426 (N_426,In_920,In_507);
or U427 (N_427,In_596,In_378);
xor U428 (N_428,In_506,In_517);
nand U429 (N_429,In_227,In_123);
or U430 (N_430,In_757,In_615);
nand U431 (N_431,In_226,In_393);
or U432 (N_432,In_354,In_269);
xor U433 (N_433,In_691,In_271);
nand U434 (N_434,In_5,In_436);
nand U435 (N_435,In_53,In_710);
xnor U436 (N_436,In_530,In_448);
and U437 (N_437,In_787,In_330);
nand U438 (N_438,In_34,In_221);
and U439 (N_439,In_877,In_382);
or U440 (N_440,In_550,In_980);
nor U441 (N_441,In_183,In_849);
or U442 (N_442,In_602,In_962);
nor U443 (N_443,In_654,In_240);
xnor U444 (N_444,In_833,In_579);
xor U445 (N_445,In_159,In_478);
nand U446 (N_446,In_290,In_194);
nor U447 (N_447,In_432,In_928);
and U448 (N_448,In_118,In_681);
nor U449 (N_449,In_907,In_205);
xnor U450 (N_450,In_634,In_916);
xnor U451 (N_451,In_745,In_793);
and U452 (N_452,In_299,In_780);
or U453 (N_453,In_804,In_306);
or U454 (N_454,In_3,In_976);
nand U455 (N_455,In_684,In_58);
and U456 (N_456,In_721,In_350);
nor U457 (N_457,In_543,In_285);
or U458 (N_458,In_335,In_9);
and U459 (N_459,In_822,In_569);
nand U460 (N_460,In_242,In_516);
nor U461 (N_461,In_999,In_883);
nand U462 (N_462,In_824,In_32);
and U463 (N_463,In_845,In_281);
nand U464 (N_464,In_470,In_598);
or U465 (N_465,In_294,In_116);
or U466 (N_466,In_716,In_266);
nor U467 (N_467,In_404,In_54);
and U468 (N_468,In_25,In_17);
or U469 (N_469,In_765,In_219);
xor U470 (N_470,In_671,In_541);
nor U471 (N_471,In_256,In_731);
and U472 (N_472,In_796,In_51);
xor U473 (N_473,In_752,In_791);
or U474 (N_474,In_126,In_842);
xor U475 (N_475,In_619,In_296);
or U476 (N_476,In_747,In_872);
nor U477 (N_477,In_539,In_548);
xor U478 (N_478,In_130,In_919);
or U479 (N_479,In_815,In_718);
xor U480 (N_480,In_871,In_317);
xor U481 (N_481,In_499,In_544);
nor U482 (N_482,In_577,In_909);
or U483 (N_483,In_911,In_477);
nor U484 (N_484,In_333,In_560);
or U485 (N_485,In_936,In_614);
and U486 (N_486,In_390,In_653);
nor U487 (N_487,In_254,In_46);
xnor U488 (N_488,In_258,In_642);
or U489 (N_489,In_276,In_60);
xnor U490 (N_490,In_626,In_729);
xnor U491 (N_491,In_972,In_981);
nand U492 (N_492,In_952,In_426);
nand U493 (N_493,In_774,In_733);
and U494 (N_494,In_760,In_961);
xnor U495 (N_495,In_64,In_397);
nand U496 (N_496,In_576,In_405);
nor U497 (N_497,In_758,In_894);
nand U498 (N_498,In_531,In_112);
or U499 (N_499,In_964,In_864);
xnor U500 (N_500,In_141,In_413);
xnor U501 (N_501,In_915,In_737);
nand U502 (N_502,In_517,In_248);
or U503 (N_503,In_556,In_773);
nor U504 (N_504,In_909,In_85);
or U505 (N_505,In_683,In_362);
or U506 (N_506,In_719,In_40);
nor U507 (N_507,In_552,In_641);
xnor U508 (N_508,In_9,In_183);
nor U509 (N_509,In_326,In_433);
nor U510 (N_510,In_950,In_471);
or U511 (N_511,In_554,In_791);
nor U512 (N_512,In_751,In_704);
xor U513 (N_513,In_404,In_931);
nor U514 (N_514,In_747,In_609);
xor U515 (N_515,In_211,In_685);
xnor U516 (N_516,In_613,In_151);
nor U517 (N_517,In_996,In_335);
or U518 (N_518,In_530,In_257);
and U519 (N_519,In_696,In_243);
and U520 (N_520,In_579,In_852);
or U521 (N_521,In_308,In_20);
nor U522 (N_522,In_499,In_126);
and U523 (N_523,In_352,In_460);
xor U524 (N_524,In_806,In_181);
xor U525 (N_525,In_145,In_324);
nor U526 (N_526,In_58,In_666);
nand U527 (N_527,In_37,In_550);
xnor U528 (N_528,In_247,In_23);
nand U529 (N_529,In_645,In_864);
xor U530 (N_530,In_162,In_873);
or U531 (N_531,In_186,In_201);
or U532 (N_532,In_401,In_69);
nand U533 (N_533,In_304,In_275);
and U534 (N_534,In_26,In_999);
nand U535 (N_535,In_943,In_22);
nor U536 (N_536,In_92,In_544);
or U537 (N_537,In_749,In_774);
xor U538 (N_538,In_298,In_792);
and U539 (N_539,In_640,In_960);
nand U540 (N_540,In_604,In_250);
nand U541 (N_541,In_266,In_636);
and U542 (N_542,In_16,In_755);
xor U543 (N_543,In_944,In_48);
xor U544 (N_544,In_422,In_698);
xnor U545 (N_545,In_66,In_699);
nand U546 (N_546,In_852,In_619);
and U547 (N_547,In_188,In_401);
nand U548 (N_548,In_605,In_329);
nor U549 (N_549,In_502,In_652);
or U550 (N_550,In_90,In_892);
xnor U551 (N_551,In_508,In_991);
and U552 (N_552,In_533,In_958);
and U553 (N_553,In_831,In_877);
nor U554 (N_554,In_327,In_170);
or U555 (N_555,In_871,In_893);
nand U556 (N_556,In_88,In_970);
or U557 (N_557,In_111,In_572);
and U558 (N_558,In_562,In_676);
or U559 (N_559,In_163,In_68);
or U560 (N_560,In_98,In_740);
nand U561 (N_561,In_344,In_313);
xor U562 (N_562,In_254,In_901);
xnor U563 (N_563,In_350,In_434);
or U564 (N_564,In_363,In_249);
or U565 (N_565,In_483,In_449);
xnor U566 (N_566,In_979,In_244);
nand U567 (N_567,In_879,In_338);
xnor U568 (N_568,In_829,In_785);
nor U569 (N_569,In_995,In_538);
and U570 (N_570,In_775,In_786);
and U571 (N_571,In_406,In_352);
and U572 (N_572,In_287,In_94);
nor U573 (N_573,In_640,In_892);
nor U574 (N_574,In_231,In_507);
or U575 (N_575,In_710,In_510);
xor U576 (N_576,In_26,In_379);
or U577 (N_577,In_741,In_918);
or U578 (N_578,In_177,In_815);
and U579 (N_579,In_281,In_763);
and U580 (N_580,In_224,In_70);
xor U581 (N_581,In_821,In_446);
nand U582 (N_582,In_742,In_45);
or U583 (N_583,In_807,In_931);
xor U584 (N_584,In_955,In_986);
xnor U585 (N_585,In_114,In_617);
and U586 (N_586,In_241,In_711);
nand U587 (N_587,In_804,In_762);
and U588 (N_588,In_181,In_844);
xnor U589 (N_589,In_499,In_516);
nand U590 (N_590,In_191,In_429);
or U591 (N_591,In_692,In_748);
or U592 (N_592,In_722,In_477);
and U593 (N_593,In_338,In_293);
xnor U594 (N_594,In_659,In_116);
and U595 (N_595,In_1,In_537);
nand U596 (N_596,In_317,In_267);
nand U597 (N_597,In_380,In_195);
nor U598 (N_598,In_799,In_370);
and U599 (N_599,In_972,In_171);
nand U600 (N_600,In_881,In_392);
xnor U601 (N_601,In_756,In_335);
or U602 (N_602,In_77,In_250);
nor U603 (N_603,In_515,In_890);
and U604 (N_604,In_660,In_87);
and U605 (N_605,In_820,In_119);
nand U606 (N_606,In_987,In_571);
or U607 (N_607,In_821,In_355);
nor U608 (N_608,In_818,In_778);
xnor U609 (N_609,In_867,In_947);
nand U610 (N_610,In_487,In_396);
or U611 (N_611,In_378,In_68);
nor U612 (N_612,In_211,In_28);
and U613 (N_613,In_118,In_870);
and U614 (N_614,In_532,In_643);
nand U615 (N_615,In_687,In_495);
xnor U616 (N_616,In_616,In_970);
nand U617 (N_617,In_164,In_762);
nand U618 (N_618,In_760,In_179);
xor U619 (N_619,In_866,In_569);
nand U620 (N_620,In_977,In_242);
and U621 (N_621,In_714,In_243);
nor U622 (N_622,In_690,In_939);
and U623 (N_623,In_248,In_358);
and U624 (N_624,In_577,In_318);
nand U625 (N_625,In_481,In_686);
and U626 (N_626,In_182,In_895);
nor U627 (N_627,In_341,In_259);
nand U628 (N_628,In_390,In_690);
or U629 (N_629,In_53,In_677);
and U630 (N_630,In_535,In_111);
or U631 (N_631,In_185,In_531);
or U632 (N_632,In_317,In_182);
or U633 (N_633,In_588,In_370);
and U634 (N_634,In_942,In_472);
nor U635 (N_635,In_3,In_655);
nand U636 (N_636,In_396,In_369);
nand U637 (N_637,In_148,In_947);
xnor U638 (N_638,In_452,In_974);
nor U639 (N_639,In_391,In_75);
and U640 (N_640,In_545,In_105);
nor U641 (N_641,In_628,In_856);
nor U642 (N_642,In_791,In_751);
and U643 (N_643,In_341,In_526);
and U644 (N_644,In_243,In_212);
nand U645 (N_645,In_102,In_561);
and U646 (N_646,In_45,In_99);
nand U647 (N_647,In_295,In_661);
nand U648 (N_648,In_36,In_308);
nand U649 (N_649,In_458,In_8);
and U650 (N_650,In_149,In_910);
nor U651 (N_651,In_168,In_194);
nor U652 (N_652,In_908,In_231);
nand U653 (N_653,In_585,In_672);
nand U654 (N_654,In_116,In_495);
or U655 (N_655,In_233,In_642);
xnor U656 (N_656,In_567,In_542);
and U657 (N_657,In_133,In_692);
or U658 (N_658,In_604,In_590);
and U659 (N_659,In_401,In_806);
xnor U660 (N_660,In_839,In_264);
xor U661 (N_661,In_260,In_18);
nor U662 (N_662,In_178,In_400);
or U663 (N_663,In_233,In_839);
and U664 (N_664,In_647,In_784);
or U665 (N_665,In_676,In_341);
and U666 (N_666,In_848,In_669);
xor U667 (N_667,In_732,In_843);
or U668 (N_668,In_849,In_868);
xor U669 (N_669,In_572,In_812);
or U670 (N_670,In_434,In_577);
nand U671 (N_671,In_217,In_349);
nand U672 (N_672,In_922,In_407);
nor U673 (N_673,In_352,In_82);
xnor U674 (N_674,In_367,In_858);
and U675 (N_675,In_147,In_660);
xnor U676 (N_676,In_947,In_864);
nor U677 (N_677,In_563,In_642);
and U678 (N_678,In_243,In_239);
nand U679 (N_679,In_257,In_994);
nor U680 (N_680,In_500,In_387);
and U681 (N_681,In_602,In_477);
and U682 (N_682,In_338,In_224);
nor U683 (N_683,In_447,In_579);
nor U684 (N_684,In_91,In_767);
and U685 (N_685,In_226,In_30);
or U686 (N_686,In_893,In_666);
and U687 (N_687,In_765,In_284);
nand U688 (N_688,In_770,In_153);
or U689 (N_689,In_530,In_269);
or U690 (N_690,In_53,In_363);
or U691 (N_691,In_493,In_647);
nand U692 (N_692,In_992,In_308);
or U693 (N_693,In_591,In_722);
nor U694 (N_694,In_65,In_375);
nand U695 (N_695,In_1,In_941);
xnor U696 (N_696,In_406,In_188);
nor U697 (N_697,In_285,In_459);
nor U698 (N_698,In_598,In_673);
or U699 (N_699,In_474,In_727);
or U700 (N_700,In_677,In_923);
xor U701 (N_701,In_93,In_680);
xor U702 (N_702,In_788,In_22);
and U703 (N_703,In_575,In_564);
nand U704 (N_704,In_410,In_57);
xor U705 (N_705,In_296,In_518);
xnor U706 (N_706,In_936,In_461);
or U707 (N_707,In_657,In_123);
and U708 (N_708,In_949,In_128);
and U709 (N_709,In_782,In_567);
xor U710 (N_710,In_474,In_207);
and U711 (N_711,In_764,In_433);
nand U712 (N_712,In_246,In_601);
or U713 (N_713,In_471,In_390);
xor U714 (N_714,In_140,In_250);
nor U715 (N_715,In_738,In_104);
nand U716 (N_716,In_983,In_168);
xnor U717 (N_717,In_139,In_749);
xor U718 (N_718,In_516,In_316);
nand U719 (N_719,In_828,In_237);
nor U720 (N_720,In_589,In_701);
nand U721 (N_721,In_513,In_780);
nand U722 (N_722,In_62,In_262);
xor U723 (N_723,In_300,In_650);
or U724 (N_724,In_911,In_541);
nand U725 (N_725,In_860,In_684);
nor U726 (N_726,In_312,In_680);
or U727 (N_727,In_684,In_160);
nand U728 (N_728,In_263,In_793);
and U729 (N_729,In_175,In_920);
and U730 (N_730,In_892,In_499);
nand U731 (N_731,In_573,In_651);
or U732 (N_732,In_149,In_591);
xor U733 (N_733,In_896,In_744);
xor U734 (N_734,In_121,In_302);
xnor U735 (N_735,In_121,In_66);
nor U736 (N_736,In_681,In_119);
and U737 (N_737,In_946,In_240);
nor U738 (N_738,In_717,In_74);
and U739 (N_739,In_509,In_355);
or U740 (N_740,In_536,In_197);
nor U741 (N_741,In_197,In_244);
and U742 (N_742,In_650,In_311);
nand U743 (N_743,In_42,In_680);
nand U744 (N_744,In_410,In_109);
nand U745 (N_745,In_206,In_363);
or U746 (N_746,In_823,In_771);
and U747 (N_747,In_269,In_847);
and U748 (N_748,In_552,In_279);
xor U749 (N_749,In_660,In_576);
and U750 (N_750,In_312,In_440);
xnor U751 (N_751,In_667,In_351);
nor U752 (N_752,In_85,In_449);
or U753 (N_753,In_784,In_515);
nand U754 (N_754,In_668,In_316);
xnor U755 (N_755,In_640,In_562);
xor U756 (N_756,In_189,In_679);
nand U757 (N_757,In_355,In_143);
nand U758 (N_758,In_383,In_218);
and U759 (N_759,In_265,In_915);
nand U760 (N_760,In_788,In_732);
nor U761 (N_761,In_899,In_320);
xnor U762 (N_762,In_17,In_285);
nor U763 (N_763,In_519,In_545);
and U764 (N_764,In_781,In_954);
nand U765 (N_765,In_404,In_892);
or U766 (N_766,In_654,In_10);
nand U767 (N_767,In_405,In_460);
xnor U768 (N_768,In_545,In_83);
or U769 (N_769,In_198,In_326);
and U770 (N_770,In_172,In_243);
nor U771 (N_771,In_667,In_265);
xnor U772 (N_772,In_35,In_843);
nor U773 (N_773,In_782,In_561);
and U774 (N_774,In_416,In_539);
xnor U775 (N_775,In_14,In_817);
nor U776 (N_776,In_710,In_90);
nand U777 (N_777,In_982,In_932);
nand U778 (N_778,In_763,In_883);
nor U779 (N_779,In_575,In_16);
nor U780 (N_780,In_204,In_43);
or U781 (N_781,In_845,In_450);
nand U782 (N_782,In_528,In_521);
and U783 (N_783,In_436,In_877);
and U784 (N_784,In_910,In_294);
nand U785 (N_785,In_419,In_746);
nor U786 (N_786,In_498,In_458);
or U787 (N_787,In_819,In_102);
xor U788 (N_788,In_998,In_146);
and U789 (N_789,In_65,In_871);
xor U790 (N_790,In_306,In_106);
nand U791 (N_791,In_30,In_984);
xor U792 (N_792,In_595,In_131);
and U793 (N_793,In_438,In_337);
and U794 (N_794,In_27,In_808);
and U795 (N_795,In_196,In_33);
or U796 (N_796,In_679,In_566);
nand U797 (N_797,In_292,In_930);
nor U798 (N_798,In_833,In_682);
nand U799 (N_799,In_461,In_370);
xnor U800 (N_800,In_812,In_116);
nand U801 (N_801,In_40,In_475);
or U802 (N_802,In_288,In_510);
xnor U803 (N_803,In_193,In_278);
xnor U804 (N_804,In_951,In_77);
nor U805 (N_805,In_643,In_371);
or U806 (N_806,In_417,In_942);
nand U807 (N_807,In_9,In_52);
nor U808 (N_808,In_249,In_171);
xnor U809 (N_809,In_758,In_611);
or U810 (N_810,In_567,In_372);
or U811 (N_811,In_217,In_584);
nand U812 (N_812,In_27,In_191);
nor U813 (N_813,In_326,In_643);
or U814 (N_814,In_226,In_802);
xor U815 (N_815,In_284,In_90);
nand U816 (N_816,In_937,In_837);
xnor U817 (N_817,In_292,In_411);
nor U818 (N_818,In_88,In_496);
nor U819 (N_819,In_691,In_585);
nand U820 (N_820,In_179,In_539);
nor U821 (N_821,In_839,In_752);
or U822 (N_822,In_335,In_125);
nand U823 (N_823,In_149,In_880);
nand U824 (N_824,In_36,In_399);
nand U825 (N_825,In_396,In_898);
and U826 (N_826,In_864,In_407);
or U827 (N_827,In_246,In_88);
xor U828 (N_828,In_101,In_924);
or U829 (N_829,In_755,In_163);
nand U830 (N_830,In_976,In_227);
nand U831 (N_831,In_433,In_670);
xnor U832 (N_832,In_272,In_274);
nor U833 (N_833,In_811,In_408);
xnor U834 (N_834,In_486,In_937);
nand U835 (N_835,In_860,In_347);
nand U836 (N_836,In_51,In_823);
nor U837 (N_837,In_42,In_710);
nand U838 (N_838,In_354,In_812);
and U839 (N_839,In_727,In_892);
xnor U840 (N_840,In_464,In_333);
or U841 (N_841,In_487,In_447);
and U842 (N_842,In_721,In_959);
xor U843 (N_843,In_357,In_604);
and U844 (N_844,In_330,In_205);
xor U845 (N_845,In_398,In_546);
nor U846 (N_846,In_382,In_453);
nand U847 (N_847,In_654,In_273);
nor U848 (N_848,In_757,In_567);
nand U849 (N_849,In_700,In_92);
and U850 (N_850,In_202,In_38);
nand U851 (N_851,In_238,In_290);
and U852 (N_852,In_279,In_911);
xor U853 (N_853,In_410,In_347);
and U854 (N_854,In_905,In_694);
nand U855 (N_855,In_282,In_563);
and U856 (N_856,In_768,In_606);
or U857 (N_857,In_324,In_679);
nand U858 (N_858,In_610,In_65);
xor U859 (N_859,In_61,In_751);
and U860 (N_860,In_909,In_67);
xor U861 (N_861,In_792,In_361);
xor U862 (N_862,In_795,In_767);
xor U863 (N_863,In_168,In_889);
and U864 (N_864,In_641,In_944);
xor U865 (N_865,In_404,In_460);
xnor U866 (N_866,In_711,In_466);
nand U867 (N_867,In_406,In_63);
xor U868 (N_868,In_406,In_855);
or U869 (N_869,In_284,In_313);
xor U870 (N_870,In_956,In_988);
nand U871 (N_871,In_606,In_333);
xor U872 (N_872,In_698,In_902);
nor U873 (N_873,In_548,In_920);
nand U874 (N_874,In_28,In_351);
xnor U875 (N_875,In_982,In_16);
xnor U876 (N_876,In_568,In_750);
and U877 (N_877,In_871,In_940);
and U878 (N_878,In_575,In_865);
nand U879 (N_879,In_721,In_480);
or U880 (N_880,In_195,In_198);
nand U881 (N_881,In_875,In_384);
xnor U882 (N_882,In_230,In_740);
nor U883 (N_883,In_477,In_759);
or U884 (N_884,In_537,In_793);
or U885 (N_885,In_661,In_828);
nor U886 (N_886,In_71,In_903);
nand U887 (N_887,In_268,In_513);
or U888 (N_888,In_243,In_623);
nor U889 (N_889,In_670,In_115);
xnor U890 (N_890,In_565,In_430);
xnor U891 (N_891,In_433,In_671);
and U892 (N_892,In_523,In_679);
nor U893 (N_893,In_806,In_50);
xnor U894 (N_894,In_12,In_114);
xnor U895 (N_895,In_198,In_32);
xor U896 (N_896,In_21,In_681);
nand U897 (N_897,In_346,In_685);
or U898 (N_898,In_366,In_455);
nor U899 (N_899,In_267,In_469);
nand U900 (N_900,In_321,In_397);
xnor U901 (N_901,In_766,In_5);
nor U902 (N_902,In_681,In_267);
nand U903 (N_903,In_445,In_162);
xnor U904 (N_904,In_590,In_295);
or U905 (N_905,In_424,In_428);
and U906 (N_906,In_381,In_687);
or U907 (N_907,In_714,In_619);
or U908 (N_908,In_692,In_877);
nand U909 (N_909,In_760,In_662);
or U910 (N_910,In_108,In_935);
and U911 (N_911,In_65,In_9);
or U912 (N_912,In_528,In_48);
and U913 (N_913,In_998,In_699);
and U914 (N_914,In_95,In_669);
or U915 (N_915,In_640,In_985);
or U916 (N_916,In_29,In_42);
nor U917 (N_917,In_556,In_650);
or U918 (N_918,In_362,In_909);
or U919 (N_919,In_232,In_265);
xor U920 (N_920,In_707,In_425);
or U921 (N_921,In_994,In_764);
and U922 (N_922,In_586,In_815);
xor U923 (N_923,In_779,In_206);
or U924 (N_924,In_960,In_353);
nor U925 (N_925,In_988,In_913);
or U926 (N_926,In_668,In_746);
or U927 (N_927,In_155,In_881);
and U928 (N_928,In_209,In_389);
or U929 (N_929,In_678,In_347);
xor U930 (N_930,In_203,In_836);
nand U931 (N_931,In_343,In_946);
or U932 (N_932,In_871,In_464);
nand U933 (N_933,In_848,In_567);
xnor U934 (N_934,In_592,In_113);
nand U935 (N_935,In_295,In_966);
nand U936 (N_936,In_625,In_79);
nand U937 (N_937,In_983,In_569);
and U938 (N_938,In_511,In_281);
nand U939 (N_939,In_29,In_505);
nand U940 (N_940,In_542,In_276);
and U941 (N_941,In_952,In_448);
xnor U942 (N_942,In_964,In_884);
or U943 (N_943,In_227,In_725);
nor U944 (N_944,In_722,In_61);
or U945 (N_945,In_331,In_878);
or U946 (N_946,In_131,In_775);
nand U947 (N_947,In_465,In_187);
nor U948 (N_948,In_971,In_462);
xor U949 (N_949,In_980,In_315);
and U950 (N_950,In_57,In_467);
or U951 (N_951,In_48,In_365);
nor U952 (N_952,In_556,In_493);
xnor U953 (N_953,In_266,In_758);
or U954 (N_954,In_839,In_988);
xnor U955 (N_955,In_78,In_851);
xnor U956 (N_956,In_137,In_257);
nand U957 (N_957,In_908,In_25);
xnor U958 (N_958,In_334,In_379);
nand U959 (N_959,In_751,In_364);
and U960 (N_960,In_136,In_419);
or U961 (N_961,In_38,In_76);
nor U962 (N_962,In_433,In_172);
or U963 (N_963,In_974,In_671);
or U964 (N_964,In_144,In_546);
or U965 (N_965,In_362,In_811);
and U966 (N_966,In_24,In_699);
or U967 (N_967,In_759,In_771);
or U968 (N_968,In_421,In_42);
nor U969 (N_969,In_452,In_790);
and U970 (N_970,In_978,In_865);
nor U971 (N_971,In_698,In_982);
or U972 (N_972,In_509,In_629);
nor U973 (N_973,In_772,In_505);
and U974 (N_974,In_672,In_389);
nand U975 (N_975,In_856,In_595);
nand U976 (N_976,In_602,In_791);
nand U977 (N_977,In_180,In_489);
nand U978 (N_978,In_94,In_657);
and U979 (N_979,In_786,In_988);
and U980 (N_980,In_173,In_386);
xnor U981 (N_981,In_394,In_704);
xnor U982 (N_982,In_43,In_124);
and U983 (N_983,In_155,In_395);
and U984 (N_984,In_840,In_768);
nand U985 (N_985,In_96,In_438);
and U986 (N_986,In_198,In_814);
nand U987 (N_987,In_718,In_697);
and U988 (N_988,In_540,In_349);
and U989 (N_989,In_911,In_79);
or U990 (N_990,In_307,In_806);
and U991 (N_991,In_235,In_356);
or U992 (N_992,In_888,In_124);
or U993 (N_993,In_868,In_910);
nand U994 (N_994,In_646,In_623);
or U995 (N_995,In_134,In_500);
nand U996 (N_996,In_13,In_797);
xnor U997 (N_997,In_888,In_758);
nand U998 (N_998,In_884,In_253);
nor U999 (N_999,In_247,In_465);
and U1000 (N_1000,In_42,In_839);
and U1001 (N_1001,In_784,In_991);
nand U1002 (N_1002,In_664,In_166);
or U1003 (N_1003,In_566,In_173);
xnor U1004 (N_1004,In_181,In_892);
nor U1005 (N_1005,In_502,In_980);
xnor U1006 (N_1006,In_266,In_625);
nand U1007 (N_1007,In_915,In_240);
or U1008 (N_1008,In_873,In_32);
xnor U1009 (N_1009,In_141,In_323);
or U1010 (N_1010,In_337,In_18);
nand U1011 (N_1011,In_262,In_431);
nor U1012 (N_1012,In_153,In_664);
nor U1013 (N_1013,In_614,In_571);
xnor U1014 (N_1014,In_438,In_576);
nand U1015 (N_1015,In_73,In_799);
nor U1016 (N_1016,In_868,In_973);
or U1017 (N_1017,In_794,In_841);
xnor U1018 (N_1018,In_602,In_481);
nor U1019 (N_1019,In_79,In_366);
nand U1020 (N_1020,In_394,In_167);
and U1021 (N_1021,In_324,In_630);
nand U1022 (N_1022,In_303,In_282);
nand U1023 (N_1023,In_618,In_949);
xor U1024 (N_1024,In_675,In_303);
and U1025 (N_1025,In_108,In_618);
xnor U1026 (N_1026,In_743,In_553);
and U1027 (N_1027,In_854,In_824);
and U1028 (N_1028,In_430,In_51);
or U1029 (N_1029,In_868,In_764);
xnor U1030 (N_1030,In_179,In_748);
nor U1031 (N_1031,In_712,In_67);
xnor U1032 (N_1032,In_42,In_596);
xor U1033 (N_1033,In_819,In_860);
or U1034 (N_1034,In_276,In_123);
nand U1035 (N_1035,In_822,In_214);
xnor U1036 (N_1036,In_898,In_237);
or U1037 (N_1037,In_938,In_250);
and U1038 (N_1038,In_877,In_211);
nor U1039 (N_1039,In_781,In_466);
and U1040 (N_1040,In_720,In_48);
nor U1041 (N_1041,In_321,In_618);
or U1042 (N_1042,In_935,In_225);
nand U1043 (N_1043,In_31,In_221);
nor U1044 (N_1044,In_683,In_202);
nor U1045 (N_1045,In_794,In_214);
and U1046 (N_1046,In_290,In_270);
nor U1047 (N_1047,In_792,In_192);
and U1048 (N_1048,In_849,In_78);
and U1049 (N_1049,In_148,In_843);
or U1050 (N_1050,In_727,In_686);
or U1051 (N_1051,In_691,In_980);
and U1052 (N_1052,In_783,In_109);
or U1053 (N_1053,In_609,In_777);
xnor U1054 (N_1054,In_852,In_281);
or U1055 (N_1055,In_952,In_617);
xnor U1056 (N_1056,In_1,In_352);
nand U1057 (N_1057,In_235,In_678);
nor U1058 (N_1058,In_711,In_796);
xor U1059 (N_1059,In_723,In_191);
or U1060 (N_1060,In_646,In_784);
xnor U1061 (N_1061,In_165,In_981);
and U1062 (N_1062,In_126,In_992);
xor U1063 (N_1063,In_111,In_406);
xnor U1064 (N_1064,In_72,In_356);
nor U1065 (N_1065,In_408,In_440);
nand U1066 (N_1066,In_371,In_674);
xor U1067 (N_1067,In_831,In_859);
or U1068 (N_1068,In_202,In_305);
nand U1069 (N_1069,In_352,In_335);
xor U1070 (N_1070,In_17,In_734);
and U1071 (N_1071,In_750,In_529);
and U1072 (N_1072,In_708,In_946);
nor U1073 (N_1073,In_52,In_60);
and U1074 (N_1074,In_540,In_820);
nand U1075 (N_1075,In_208,In_654);
nand U1076 (N_1076,In_514,In_109);
xor U1077 (N_1077,In_202,In_88);
xor U1078 (N_1078,In_304,In_28);
xor U1079 (N_1079,In_209,In_440);
nand U1080 (N_1080,In_907,In_557);
nand U1081 (N_1081,In_899,In_630);
nand U1082 (N_1082,In_977,In_988);
nor U1083 (N_1083,In_406,In_867);
nor U1084 (N_1084,In_517,In_551);
nor U1085 (N_1085,In_501,In_416);
xnor U1086 (N_1086,In_36,In_711);
nand U1087 (N_1087,In_951,In_326);
and U1088 (N_1088,In_403,In_806);
nor U1089 (N_1089,In_323,In_368);
nor U1090 (N_1090,In_139,In_970);
nand U1091 (N_1091,In_750,In_97);
xnor U1092 (N_1092,In_410,In_969);
or U1093 (N_1093,In_312,In_614);
nand U1094 (N_1094,In_165,In_302);
or U1095 (N_1095,In_559,In_945);
nor U1096 (N_1096,In_633,In_606);
xnor U1097 (N_1097,In_560,In_149);
and U1098 (N_1098,In_685,In_691);
nand U1099 (N_1099,In_422,In_979);
and U1100 (N_1100,In_766,In_895);
nand U1101 (N_1101,In_796,In_899);
or U1102 (N_1102,In_836,In_310);
and U1103 (N_1103,In_214,In_645);
xnor U1104 (N_1104,In_501,In_511);
nor U1105 (N_1105,In_158,In_9);
and U1106 (N_1106,In_190,In_596);
xnor U1107 (N_1107,In_526,In_933);
nor U1108 (N_1108,In_651,In_23);
xnor U1109 (N_1109,In_891,In_287);
or U1110 (N_1110,In_923,In_27);
and U1111 (N_1111,In_31,In_943);
and U1112 (N_1112,In_128,In_65);
xnor U1113 (N_1113,In_899,In_820);
nand U1114 (N_1114,In_890,In_788);
nand U1115 (N_1115,In_41,In_96);
nand U1116 (N_1116,In_937,In_216);
xor U1117 (N_1117,In_724,In_830);
nand U1118 (N_1118,In_165,In_805);
nand U1119 (N_1119,In_314,In_561);
nand U1120 (N_1120,In_719,In_838);
nand U1121 (N_1121,In_553,In_281);
or U1122 (N_1122,In_93,In_949);
and U1123 (N_1123,In_764,In_3);
or U1124 (N_1124,In_784,In_664);
xor U1125 (N_1125,In_272,In_960);
or U1126 (N_1126,In_896,In_988);
nand U1127 (N_1127,In_703,In_253);
nand U1128 (N_1128,In_383,In_998);
nor U1129 (N_1129,In_579,In_92);
and U1130 (N_1130,In_765,In_160);
xnor U1131 (N_1131,In_643,In_82);
or U1132 (N_1132,In_563,In_649);
and U1133 (N_1133,In_600,In_675);
xnor U1134 (N_1134,In_156,In_823);
nand U1135 (N_1135,In_431,In_107);
nor U1136 (N_1136,In_115,In_363);
nand U1137 (N_1137,In_206,In_780);
or U1138 (N_1138,In_878,In_891);
nand U1139 (N_1139,In_254,In_633);
and U1140 (N_1140,In_245,In_944);
or U1141 (N_1141,In_778,In_554);
nand U1142 (N_1142,In_874,In_995);
or U1143 (N_1143,In_751,In_674);
or U1144 (N_1144,In_195,In_654);
nand U1145 (N_1145,In_929,In_562);
and U1146 (N_1146,In_227,In_534);
nor U1147 (N_1147,In_311,In_173);
nand U1148 (N_1148,In_848,In_644);
and U1149 (N_1149,In_765,In_383);
nand U1150 (N_1150,In_374,In_408);
or U1151 (N_1151,In_634,In_63);
or U1152 (N_1152,In_709,In_693);
or U1153 (N_1153,In_639,In_609);
xor U1154 (N_1154,In_440,In_918);
xnor U1155 (N_1155,In_762,In_672);
or U1156 (N_1156,In_427,In_477);
nor U1157 (N_1157,In_396,In_117);
or U1158 (N_1158,In_723,In_967);
or U1159 (N_1159,In_436,In_586);
nand U1160 (N_1160,In_324,In_789);
and U1161 (N_1161,In_420,In_43);
or U1162 (N_1162,In_47,In_919);
nor U1163 (N_1163,In_508,In_347);
nand U1164 (N_1164,In_788,In_42);
nor U1165 (N_1165,In_253,In_500);
nor U1166 (N_1166,In_706,In_805);
or U1167 (N_1167,In_485,In_386);
and U1168 (N_1168,In_715,In_655);
nor U1169 (N_1169,In_479,In_31);
xor U1170 (N_1170,In_913,In_633);
xnor U1171 (N_1171,In_88,In_504);
nor U1172 (N_1172,In_968,In_817);
and U1173 (N_1173,In_101,In_129);
nand U1174 (N_1174,In_31,In_456);
nor U1175 (N_1175,In_708,In_395);
nand U1176 (N_1176,In_671,In_567);
xor U1177 (N_1177,In_542,In_526);
and U1178 (N_1178,In_668,In_625);
nor U1179 (N_1179,In_394,In_310);
or U1180 (N_1180,In_714,In_890);
nand U1181 (N_1181,In_616,In_709);
xnor U1182 (N_1182,In_690,In_801);
and U1183 (N_1183,In_129,In_970);
nand U1184 (N_1184,In_345,In_384);
or U1185 (N_1185,In_745,In_266);
and U1186 (N_1186,In_449,In_636);
and U1187 (N_1187,In_775,In_430);
or U1188 (N_1188,In_473,In_626);
and U1189 (N_1189,In_308,In_366);
xor U1190 (N_1190,In_36,In_20);
and U1191 (N_1191,In_776,In_935);
or U1192 (N_1192,In_894,In_485);
nor U1193 (N_1193,In_200,In_946);
nand U1194 (N_1194,In_130,In_954);
xnor U1195 (N_1195,In_15,In_326);
xor U1196 (N_1196,In_581,In_667);
nand U1197 (N_1197,In_367,In_449);
xor U1198 (N_1198,In_391,In_290);
xor U1199 (N_1199,In_889,In_649);
nor U1200 (N_1200,In_595,In_407);
or U1201 (N_1201,In_7,In_127);
and U1202 (N_1202,In_212,In_537);
and U1203 (N_1203,In_41,In_575);
nand U1204 (N_1204,In_788,In_551);
nand U1205 (N_1205,In_576,In_603);
nand U1206 (N_1206,In_757,In_349);
nor U1207 (N_1207,In_492,In_156);
and U1208 (N_1208,In_469,In_961);
nor U1209 (N_1209,In_427,In_245);
xor U1210 (N_1210,In_673,In_490);
xnor U1211 (N_1211,In_480,In_338);
xor U1212 (N_1212,In_326,In_665);
nand U1213 (N_1213,In_248,In_477);
and U1214 (N_1214,In_635,In_830);
or U1215 (N_1215,In_618,In_975);
and U1216 (N_1216,In_795,In_324);
nor U1217 (N_1217,In_723,In_701);
and U1218 (N_1218,In_51,In_520);
and U1219 (N_1219,In_591,In_338);
nand U1220 (N_1220,In_571,In_937);
or U1221 (N_1221,In_911,In_898);
and U1222 (N_1222,In_642,In_954);
nand U1223 (N_1223,In_145,In_711);
nand U1224 (N_1224,In_129,In_271);
nand U1225 (N_1225,In_923,In_749);
xor U1226 (N_1226,In_347,In_208);
and U1227 (N_1227,In_302,In_215);
xor U1228 (N_1228,In_845,In_846);
or U1229 (N_1229,In_193,In_725);
nor U1230 (N_1230,In_168,In_801);
nor U1231 (N_1231,In_349,In_914);
xor U1232 (N_1232,In_665,In_205);
and U1233 (N_1233,In_979,In_255);
nor U1234 (N_1234,In_883,In_200);
nand U1235 (N_1235,In_482,In_113);
or U1236 (N_1236,In_493,In_541);
and U1237 (N_1237,In_906,In_138);
xor U1238 (N_1238,In_211,In_460);
or U1239 (N_1239,In_584,In_936);
and U1240 (N_1240,In_877,In_545);
nand U1241 (N_1241,In_543,In_783);
nand U1242 (N_1242,In_29,In_46);
nand U1243 (N_1243,In_539,In_21);
or U1244 (N_1244,In_100,In_833);
and U1245 (N_1245,In_146,In_974);
and U1246 (N_1246,In_284,In_737);
and U1247 (N_1247,In_962,In_157);
and U1248 (N_1248,In_917,In_493);
nor U1249 (N_1249,In_435,In_177);
and U1250 (N_1250,In_819,In_878);
nand U1251 (N_1251,In_381,In_768);
or U1252 (N_1252,In_939,In_507);
nand U1253 (N_1253,In_66,In_580);
xor U1254 (N_1254,In_885,In_48);
and U1255 (N_1255,In_8,In_584);
or U1256 (N_1256,In_893,In_418);
or U1257 (N_1257,In_714,In_843);
and U1258 (N_1258,In_881,In_934);
or U1259 (N_1259,In_82,In_767);
nor U1260 (N_1260,In_175,In_428);
and U1261 (N_1261,In_829,In_390);
and U1262 (N_1262,In_313,In_632);
nor U1263 (N_1263,In_467,In_320);
nand U1264 (N_1264,In_185,In_389);
or U1265 (N_1265,In_989,In_129);
or U1266 (N_1266,In_980,In_123);
nand U1267 (N_1267,In_806,In_944);
xnor U1268 (N_1268,In_630,In_154);
nand U1269 (N_1269,In_702,In_400);
xnor U1270 (N_1270,In_536,In_947);
nand U1271 (N_1271,In_306,In_6);
and U1272 (N_1272,In_843,In_465);
nor U1273 (N_1273,In_5,In_426);
or U1274 (N_1274,In_517,In_26);
and U1275 (N_1275,In_356,In_512);
nand U1276 (N_1276,In_724,In_181);
or U1277 (N_1277,In_436,In_445);
nor U1278 (N_1278,In_387,In_282);
xnor U1279 (N_1279,In_308,In_897);
or U1280 (N_1280,In_27,In_888);
nand U1281 (N_1281,In_283,In_804);
nor U1282 (N_1282,In_664,In_957);
nand U1283 (N_1283,In_565,In_109);
or U1284 (N_1284,In_613,In_832);
and U1285 (N_1285,In_478,In_379);
and U1286 (N_1286,In_106,In_209);
nor U1287 (N_1287,In_851,In_712);
or U1288 (N_1288,In_238,In_483);
or U1289 (N_1289,In_308,In_354);
or U1290 (N_1290,In_208,In_19);
or U1291 (N_1291,In_200,In_447);
or U1292 (N_1292,In_115,In_689);
nor U1293 (N_1293,In_877,In_419);
xor U1294 (N_1294,In_575,In_309);
xor U1295 (N_1295,In_410,In_138);
nand U1296 (N_1296,In_180,In_710);
nor U1297 (N_1297,In_432,In_77);
xor U1298 (N_1298,In_160,In_101);
or U1299 (N_1299,In_167,In_91);
nand U1300 (N_1300,In_745,In_852);
nand U1301 (N_1301,In_831,In_324);
xnor U1302 (N_1302,In_133,In_216);
nor U1303 (N_1303,In_24,In_379);
nor U1304 (N_1304,In_896,In_476);
xor U1305 (N_1305,In_323,In_563);
and U1306 (N_1306,In_959,In_737);
xnor U1307 (N_1307,In_324,In_925);
and U1308 (N_1308,In_359,In_700);
xnor U1309 (N_1309,In_522,In_992);
xnor U1310 (N_1310,In_602,In_66);
xor U1311 (N_1311,In_445,In_648);
nor U1312 (N_1312,In_673,In_358);
nor U1313 (N_1313,In_744,In_653);
nor U1314 (N_1314,In_268,In_97);
nor U1315 (N_1315,In_26,In_757);
nand U1316 (N_1316,In_697,In_456);
or U1317 (N_1317,In_721,In_695);
xnor U1318 (N_1318,In_313,In_11);
xnor U1319 (N_1319,In_27,In_836);
nand U1320 (N_1320,In_945,In_771);
nand U1321 (N_1321,In_602,In_789);
xor U1322 (N_1322,In_515,In_75);
and U1323 (N_1323,In_784,In_621);
nor U1324 (N_1324,In_638,In_634);
nor U1325 (N_1325,In_935,In_190);
and U1326 (N_1326,In_772,In_609);
xnor U1327 (N_1327,In_260,In_251);
nor U1328 (N_1328,In_989,In_159);
and U1329 (N_1329,In_716,In_648);
nand U1330 (N_1330,In_210,In_865);
and U1331 (N_1331,In_64,In_601);
or U1332 (N_1332,In_639,In_921);
nor U1333 (N_1333,In_731,In_423);
and U1334 (N_1334,In_611,In_643);
xnor U1335 (N_1335,In_374,In_937);
nand U1336 (N_1336,In_762,In_691);
and U1337 (N_1337,In_432,In_840);
xor U1338 (N_1338,In_211,In_786);
or U1339 (N_1339,In_478,In_351);
nor U1340 (N_1340,In_892,In_270);
nor U1341 (N_1341,In_37,In_65);
nand U1342 (N_1342,In_807,In_976);
nor U1343 (N_1343,In_572,In_701);
xnor U1344 (N_1344,In_573,In_302);
xnor U1345 (N_1345,In_79,In_42);
nor U1346 (N_1346,In_991,In_147);
or U1347 (N_1347,In_938,In_370);
nand U1348 (N_1348,In_377,In_257);
or U1349 (N_1349,In_986,In_409);
nor U1350 (N_1350,In_517,In_836);
or U1351 (N_1351,In_672,In_945);
nand U1352 (N_1352,In_307,In_881);
nand U1353 (N_1353,In_753,In_847);
nor U1354 (N_1354,In_383,In_569);
xor U1355 (N_1355,In_390,In_306);
xnor U1356 (N_1356,In_856,In_203);
or U1357 (N_1357,In_936,In_444);
nor U1358 (N_1358,In_997,In_403);
nand U1359 (N_1359,In_787,In_512);
xor U1360 (N_1360,In_322,In_656);
xnor U1361 (N_1361,In_874,In_668);
or U1362 (N_1362,In_93,In_33);
nand U1363 (N_1363,In_621,In_563);
nor U1364 (N_1364,In_697,In_883);
nor U1365 (N_1365,In_87,In_610);
nor U1366 (N_1366,In_860,In_859);
or U1367 (N_1367,In_969,In_403);
xnor U1368 (N_1368,In_161,In_798);
xnor U1369 (N_1369,In_478,In_999);
or U1370 (N_1370,In_799,In_471);
or U1371 (N_1371,In_611,In_938);
and U1372 (N_1372,In_937,In_197);
xor U1373 (N_1373,In_660,In_516);
xor U1374 (N_1374,In_850,In_705);
nor U1375 (N_1375,In_401,In_26);
nor U1376 (N_1376,In_561,In_241);
nand U1377 (N_1377,In_484,In_74);
xnor U1378 (N_1378,In_481,In_824);
or U1379 (N_1379,In_76,In_184);
or U1380 (N_1380,In_818,In_966);
nor U1381 (N_1381,In_543,In_222);
nand U1382 (N_1382,In_862,In_582);
nand U1383 (N_1383,In_552,In_330);
nor U1384 (N_1384,In_524,In_879);
nor U1385 (N_1385,In_95,In_579);
and U1386 (N_1386,In_136,In_200);
nor U1387 (N_1387,In_327,In_192);
or U1388 (N_1388,In_991,In_879);
and U1389 (N_1389,In_445,In_807);
or U1390 (N_1390,In_3,In_14);
and U1391 (N_1391,In_906,In_561);
and U1392 (N_1392,In_512,In_16);
xnor U1393 (N_1393,In_546,In_529);
nand U1394 (N_1394,In_202,In_168);
and U1395 (N_1395,In_214,In_975);
xnor U1396 (N_1396,In_108,In_775);
or U1397 (N_1397,In_870,In_52);
nor U1398 (N_1398,In_832,In_234);
xor U1399 (N_1399,In_338,In_996);
or U1400 (N_1400,In_409,In_105);
xor U1401 (N_1401,In_162,In_175);
and U1402 (N_1402,In_86,In_694);
nand U1403 (N_1403,In_842,In_648);
and U1404 (N_1404,In_476,In_997);
xor U1405 (N_1405,In_13,In_404);
xor U1406 (N_1406,In_370,In_766);
or U1407 (N_1407,In_839,In_303);
xor U1408 (N_1408,In_619,In_563);
or U1409 (N_1409,In_260,In_878);
nand U1410 (N_1410,In_230,In_649);
and U1411 (N_1411,In_849,In_333);
and U1412 (N_1412,In_138,In_330);
nand U1413 (N_1413,In_218,In_687);
and U1414 (N_1414,In_339,In_630);
or U1415 (N_1415,In_842,In_689);
nor U1416 (N_1416,In_63,In_843);
xnor U1417 (N_1417,In_635,In_828);
nor U1418 (N_1418,In_882,In_502);
nor U1419 (N_1419,In_31,In_896);
or U1420 (N_1420,In_205,In_883);
nor U1421 (N_1421,In_345,In_125);
xor U1422 (N_1422,In_220,In_329);
nor U1423 (N_1423,In_611,In_464);
nor U1424 (N_1424,In_290,In_938);
nand U1425 (N_1425,In_95,In_101);
and U1426 (N_1426,In_334,In_541);
and U1427 (N_1427,In_843,In_245);
and U1428 (N_1428,In_766,In_538);
nor U1429 (N_1429,In_710,In_761);
nand U1430 (N_1430,In_738,In_753);
nor U1431 (N_1431,In_390,In_750);
xor U1432 (N_1432,In_374,In_768);
nor U1433 (N_1433,In_737,In_5);
nand U1434 (N_1434,In_670,In_891);
nand U1435 (N_1435,In_566,In_576);
and U1436 (N_1436,In_182,In_62);
or U1437 (N_1437,In_661,In_741);
nor U1438 (N_1438,In_962,In_612);
nand U1439 (N_1439,In_376,In_169);
nor U1440 (N_1440,In_114,In_543);
or U1441 (N_1441,In_954,In_914);
and U1442 (N_1442,In_963,In_484);
and U1443 (N_1443,In_593,In_677);
and U1444 (N_1444,In_262,In_213);
nor U1445 (N_1445,In_768,In_73);
or U1446 (N_1446,In_991,In_478);
nand U1447 (N_1447,In_472,In_591);
and U1448 (N_1448,In_496,In_573);
nand U1449 (N_1449,In_576,In_551);
and U1450 (N_1450,In_504,In_582);
xnor U1451 (N_1451,In_981,In_35);
or U1452 (N_1452,In_392,In_970);
nand U1453 (N_1453,In_238,In_693);
and U1454 (N_1454,In_658,In_230);
nand U1455 (N_1455,In_523,In_652);
or U1456 (N_1456,In_17,In_496);
nor U1457 (N_1457,In_651,In_462);
nand U1458 (N_1458,In_444,In_903);
nor U1459 (N_1459,In_902,In_615);
nor U1460 (N_1460,In_62,In_21);
xor U1461 (N_1461,In_603,In_984);
nand U1462 (N_1462,In_927,In_758);
nor U1463 (N_1463,In_597,In_897);
and U1464 (N_1464,In_72,In_802);
nor U1465 (N_1465,In_479,In_468);
and U1466 (N_1466,In_308,In_191);
or U1467 (N_1467,In_83,In_640);
or U1468 (N_1468,In_494,In_267);
and U1469 (N_1469,In_956,In_304);
or U1470 (N_1470,In_281,In_325);
or U1471 (N_1471,In_725,In_996);
nand U1472 (N_1472,In_652,In_229);
nor U1473 (N_1473,In_666,In_635);
xor U1474 (N_1474,In_541,In_994);
xnor U1475 (N_1475,In_341,In_774);
and U1476 (N_1476,In_785,In_184);
or U1477 (N_1477,In_692,In_994);
nor U1478 (N_1478,In_484,In_288);
nand U1479 (N_1479,In_181,In_609);
nor U1480 (N_1480,In_669,In_856);
xnor U1481 (N_1481,In_409,In_307);
or U1482 (N_1482,In_739,In_476);
nand U1483 (N_1483,In_840,In_514);
xnor U1484 (N_1484,In_656,In_70);
nor U1485 (N_1485,In_1,In_34);
or U1486 (N_1486,In_519,In_462);
and U1487 (N_1487,In_601,In_426);
xor U1488 (N_1488,In_910,In_654);
nand U1489 (N_1489,In_683,In_825);
nand U1490 (N_1490,In_126,In_87);
and U1491 (N_1491,In_905,In_211);
xnor U1492 (N_1492,In_388,In_562);
xor U1493 (N_1493,In_135,In_747);
and U1494 (N_1494,In_291,In_122);
nand U1495 (N_1495,In_616,In_581);
and U1496 (N_1496,In_848,In_929);
and U1497 (N_1497,In_178,In_693);
nand U1498 (N_1498,In_452,In_920);
or U1499 (N_1499,In_870,In_926);
or U1500 (N_1500,In_467,In_251);
nor U1501 (N_1501,In_685,In_147);
or U1502 (N_1502,In_989,In_149);
or U1503 (N_1503,In_970,In_650);
xnor U1504 (N_1504,In_459,In_193);
nand U1505 (N_1505,In_822,In_598);
or U1506 (N_1506,In_312,In_299);
nand U1507 (N_1507,In_500,In_266);
xnor U1508 (N_1508,In_453,In_510);
or U1509 (N_1509,In_551,In_930);
and U1510 (N_1510,In_915,In_353);
xnor U1511 (N_1511,In_237,In_114);
nand U1512 (N_1512,In_705,In_824);
and U1513 (N_1513,In_527,In_714);
nor U1514 (N_1514,In_916,In_483);
and U1515 (N_1515,In_371,In_486);
nor U1516 (N_1516,In_232,In_452);
nor U1517 (N_1517,In_360,In_975);
or U1518 (N_1518,In_260,In_882);
and U1519 (N_1519,In_822,In_363);
nand U1520 (N_1520,In_623,In_909);
nand U1521 (N_1521,In_798,In_630);
xnor U1522 (N_1522,In_772,In_596);
nand U1523 (N_1523,In_897,In_14);
or U1524 (N_1524,In_691,In_437);
and U1525 (N_1525,In_436,In_369);
nand U1526 (N_1526,In_473,In_726);
and U1527 (N_1527,In_573,In_451);
nor U1528 (N_1528,In_952,In_551);
nand U1529 (N_1529,In_975,In_603);
nand U1530 (N_1530,In_265,In_319);
xnor U1531 (N_1531,In_434,In_564);
or U1532 (N_1532,In_600,In_22);
nor U1533 (N_1533,In_485,In_496);
nand U1534 (N_1534,In_627,In_534);
xnor U1535 (N_1535,In_12,In_725);
nor U1536 (N_1536,In_224,In_422);
xnor U1537 (N_1537,In_427,In_249);
and U1538 (N_1538,In_856,In_523);
and U1539 (N_1539,In_550,In_939);
xnor U1540 (N_1540,In_924,In_711);
xnor U1541 (N_1541,In_22,In_784);
or U1542 (N_1542,In_558,In_723);
and U1543 (N_1543,In_259,In_858);
nand U1544 (N_1544,In_534,In_628);
nor U1545 (N_1545,In_406,In_929);
or U1546 (N_1546,In_233,In_337);
nor U1547 (N_1547,In_229,In_122);
nor U1548 (N_1548,In_100,In_281);
xor U1549 (N_1549,In_229,In_129);
xnor U1550 (N_1550,In_941,In_392);
nor U1551 (N_1551,In_960,In_626);
or U1552 (N_1552,In_304,In_258);
nand U1553 (N_1553,In_826,In_125);
and U1554 (N_1554,In_734,In_175);
xor U1555 (N_1555,In_677,In_494);
nor U1556 (N_1556,In_79,In_635);
xor U1557 (N_1557,In_817,In_893);
and U1558 (N_1558,In_821,In_827);
nand U1559 (N_1559,In_397,In_42);
or U1560 (N_1560,In_901,In_432);
xor U1561 (N_1561,In_958,In_70);
nand U1562 (N_1562,In_5,In_758);
nand U1563 (N_1563,In_15,In_28);
and U1564 (N_1564,In_153,In_113);
xor U1565 (N_1565,In_621,In_905);
nand U1566 (N_1566,In_760,In_569);
nand U1567 (N_1567,In_881,In_607);
nand U1568 (N_1568,In_169,In_965);
xnor U1569 (N_1569,In_13,In_10);
and U1570 (N_1570,In_30,In_175);
nand U1571 (N_1571,In_21,In_353);
nand U1572 (N_1572,In_180,In_233);
xor U1573 (N_1573,In_305,In_920);
and U1574 (N_1574,In_580,In_377);
nor U1575 (N_1575,In_6,In_692);
xnor U1576 (N_1576,In_692,In_793);
or U1577 (N_1577,In_784,In_609);
or U1578 (N_1578,In_528,In_450);
and U1579 (N_1579,In_909,In_940);
xor U1580 (N_1580,In_872,In_973);
xor U1581 (N_1581,In_580,In_607);
nor U1582 (N_1582,In_207,In_663);
or U1583 (N_1583,In_393,In_721);
or U1584 (N_1584,In_532,In_187);
nand U1585 (N_1585,In_354,In_193);
or U1586 (N_1586,In_248,In_671);
nor U1587 (N_1587,In_9,In_509);
and U1588 (N_1588,In_603,In_376);
xor U1589 (N_1589,In_917,In_728);
xnor U1590 (N_1590,In_233,In_127);
nor U1591 (N_1591,In_236,In_739);
nand U1592 (N_1592,In_454,In_231);
nor U1593 (N_1593,In_549,In_308);
xor U1594 (N_1594,In_502,In_144);
or U1595 (N_1595,In_578,In_332);
or U1596 (N_1596,In_491,In_289);
or U1597 (N_1597,In_909,In_950);
nand U1598 (N_1598,In_575,In_732);
or U1599 (N_1599,In_492,In_786);
nand U1600 (N_1600,In_654,In_183);
and U1601 (N_1601,In_158,In_892);
or U1602 (N_1602,In_798,In_489);
or U1603 (N_1603,In_898,In_624);
nand U1604 (N_1604,In_381,In_523);
or U1605 (N_1605,In_886,In_394);
nor U1606 (N_1606,In_468,In_30);
or U1607 (N_1607,In_391,In_365);
xnor U1608 (N_1608,In_792,In_764);
or U1609 (N_1609,In_652,In_592);
xor U1610 (N_1610,In_953,In_856);
nor U1611 (N_1611,In_335,In_897);
nor U1612 (N_1612,In_935,In_176);
nand U1613 (N_1613,In_221,In_944);
or U1614 (N_1614,In_49,In_242);
nor U1615 (N_1615,In_64,In_880);
and U1616 (N_1616,In_711,In_981);
nand U1617 (N_1617,In_538,In_306);
and U1618 (N_1618,In_280,In_905);
and U1619 (N_1619,In_11,In_554);
and U1620 (N_1620,In_26,In_40);
nor U1621 (N_1621,In_545,In_314);
nor U1622 (N_1622,In_827,In_594);
and U1623 (N_1623,In_735,In_744);
and U1624 (N_1624,In_681,In_462);
nand U1625 (N_1625,In_16,In_275);
or U1626 (N_1626,In_905,In_151);
nor U1627 (N_1627,In_404,In_58);
xor U1628 (N_1628,In_617,In_88);
xor U1629 (N_1629,In_151,In_570);
nor U1630 (N_1630,In_277,In_64);
nand U1631 (N_1631,In_490,In_31);
xnor U1632 (N_1632,In_412,In_576);
and U1633 (N_1633,In_497,In_690);
and U1634 (N_1634,In_700,In_127);
xor U1635 (N_1635,In_339,In_1);
and U1636 (N_1636,In_935,In_542);
or U1637 (N_1637,In_550,In_689);
nor U1638 (N_1638,In_97,In_28);
and U1639 (N_1639,In_749,In_336);
or U1640 (N_1640,In_486,In_396);
nor U1641 (N_1641,In_525,In_798);
xor U1642 (N_1642,In_430,In_434);
nand U1643 (N_1643,In_428,In_139);
nand U1644 (N_1644,In_254,In_902);
nand U1645 (N_1645,In_377,In_80);
and U1646 (N_1646,In_202,In_467);
nand U1647 (N_1647,In_724,In_730);
nand U1648 (N_1648,In_170,In_761);
nand U1649 (N_1649,In_492,In_653);
nand U1650 (N_1650,In_800,In_532);
nand U1651 (N_1651,In_859,In_343);
and U1652 (N_1652,In_215,In_367);
and U1653 (N_1653,In_547,In_205);
xor U1654 (N_1654,In_796,In_218);
nand U1655 (N_1655,In_153,In_969);
nor U1656 (N_1656,In_906,In_466);
nand U1657 (N_1657,In_292,In_501);
or U1658 (N_1658,In_189,In_976);
xor U1659 (N_1659,In_845,In_215);
xor U1660 (N_1660,In_34,In_26);
nand U1661 (N_1661,In_505,In_119);
or U1662 (N_1662,In_992,In_30);
or U1663 (N_1663,In_334,In_311);
xnor U1664 (N_1664,In_3,In_95);
xnor U1665 (N_1665,In_396,In_588);
nor U1666 (N_1666,In_668,In_291);
nand U1667 (N_1667,In_740,In_77);
and U1668 (N_1668,In_729,In_589);
nand U1669 (N_1669,In_298,In_213);
or U1670 (N_1670,In_614,In_238);
and U1671 (N_1671,In_195,In_821);
or U1672 (N_1672,In_783,In_58);
and U1673 (N_1673,In_20,In_61);
nor U1674 (N_1674,In_961,In_152);
and U1675 (N_1675,In_363,In_618);
nor U1676 (N_1676,In_269,In_972);
and U1677 (N_1677,In_53,In_28);
and U1678 (N_1678,In_64,In_667);
and U1679 (N_1679,In_473,In_261);
nor U1680 (N_1680,In_849,In_580);
nor U1681 (N_1681,In_427,In_548);
nand U1682 (N_1682,In_622,In_198);
nand U1683 (N_1683,In_752,In_108);
nand U1684 (N_1684,In_538,In_74);
nand U1685 (N_1685,In_685,In_528);
xnor U1686 (N_1686,In_751,In_174);
nand U1687 (N_1687,In_866,In_321);
xnor U1688 (N_1688,In_833,In_451);
nor U1689 (N_1689,In_3,In_954);
and U1690 (N_1690,In_675,In_549);
xnor U1691 (N_1691,In_527,In_253);
xnor U1692 (N_1692,In_0,In_629);
or U1693 (N_1693,In_230,In_8);
nor U1694 (N_1694,In_80,In_899);
and U1695 (N_1695,In_676,In_8);
nand U1696 (N_1696,In_683,In_850);
nand U1697 (N_1697,In_290,In_210);
and U1698 (N_1698,In_506,In_726);
nand U1699 (N_1699,In_823,In_865);
or U1700 (N_1700,In_286,In_994);
or U1701 (N_1701,In_291,In_437);
nand U1702 (N_1702,In_546,In_221);
xor U1703 (N_1703,In_934,In_671);
xor U1704 (N_1704,In_146,In_837);
and U1705 (N_1705,In_132,In_454);
nor U1706 (N_1706,In_173,In_62);
or U1707 (N_1707,In_496,In_178);
or U1708 (N_1708,In_510,In_49);
nand U1709 (N_1709,In_429,In_411);
and U1710 (N_1710,In_925,In_119);
nand U1711 (N_1711,In_729,In_706);
or U1712 (N_1712,In_324,In_272);
or U1713 (N_1713,In_641,In_775);
and U1714 (N_1714,In_967,In_847);
and U1715 (N_1715,In_720,In_353);
or U1716 (N_1716,In_935,In_680);
xor U1717 (N_1717,In_340,In_853);
and U1718 (N_1718,In_7,In_500);
nand U1719 (N_1719,In_484,In_858);
nand U1720 (N_1720,In_419,In_58);
and U1721 (N_1721,In_376,In_970);
xnor U1722 (N_1722,In_217,In_650);
xor U1723 (N_1723,In_421,In_462);
nand U1724 (N_1724,In_705,In_93);
and U1725 (N_1725,In_623,In_778);
xor U1726 (N_1726,In_232,In_579);
nand U1727 (N_1727,In_344,In_703);
or U1728 (N_1728,In_28,In_668);
nor U1729 (N_1729,In_629,In_521);
or U1730 (N_1730,In_416,In_500);
nor U1731 (N_1731,In_817,In_701);
nor U1732 (N_1732,In_864,In_208);
nand U1733 (N_1733,In_394,In_278);
or U1734 (N_1734,In_571,In_58);
nor U1735 (N_1735,In_478,In_226);
xnor U1736 (N_1736,In_978,In_306);
xnor U1737 (N_1737,In_446,In_127);
nand U1738 (N_1738,In_325,In_192);
nor U1739 (N_1739,In_486,In_322);
xnor U1740 (N_1740,In_402,In_588);
and U1741 (N_1741,In_765,In_917);
nor U1742 (N_1742,In_914,In_408);
nor U1743 (N_1743,In_635,In_748);
and U1744 (N_1744,In_224,In_87);
nor U1745 (N_1745,In_730,In_541);
or U1746 (N_1746,In_754,In_261);
or U1747 (N_1747,In_12,In_388);
nand U1748 (N_1748,In_497,In_543);
nand U1749 (N_1749,In_555,In_670);
or U1750 (N_1750,In_644,In_593);
xor U1751 (N_1751,In_530,In_917);
xor U1752 (N_1752,In_640,In_926);
or U1753 (N_1753,In_647,In_416);
nand U1754 (N_1754,In_834,In_470);
and U1755 (N_1755,In_754,In_492);
xnor U1756 (N_1756,In_455,In_964);
and U1757 (N_1757,In_517,In_256);
nand U1758 (N_1758,In_853,In_833);
xor U1759 (N_1759,In_298,In_871);
xor U1760 (N_1760,In_927,In_585);
or U1761 (N_1761,In_472,In_133);
or U1762 (N_1762,In_97,In_247);
nor U1763 (N_1763,In_319,In_371);
nor U1764 (N_1764,In_404,In_137);
and U1765 (N_1765,In_853,In_257);
nor U1766 (N_1766,In_988,In_904);
nor U1767 (N_1767,In_833,In_771);
or U1768 (N_1768,In_553,In_955);
nand U1769 (N_1769,In_181,In_270);
and U1770 (N_1770,In_956,In_67);
nand U1771 (N_1771,In_233,In_544);
nor U1772 (N_1772,In_24,In_364);
xnor U1773 (N_1773,In_365,In_510);
or U1774 (N_1774,In_802,In_584);
or U1775 (N_1775,In_999,In_188);
xnor U1776 (N_1776,In_322,In_194);
nor U1777 (N_1777,In_927,In_204);
or U1778 (N_1778,In_718,In_985);
or U1779 (N_1779,In_164,In_260);
or U1780 (N_1780,In_482,In_65);
and U1781 (N_1781,In_351,In_647);
nand U1782 (N_1782,In_370,In_896);
or U1783 (N_1783,In_532,In_198);
and U1784 (N_1784,In_984,In_610);
xor U1785 (N_1785,In_872,In_665);
and U1786 (N_1786,In_540,In_744);
nor U1787 (N_1787,In_655,In_860);
nand U1788 (N_1788,In_318,In_925);
or U1789 (N_1789,In_995,In_786);
nand U1790 (N_1790,In_585,In_952);
xnor U1791 (N_1791,In_419,In_975);
or U1792 (N_1792,In_844,In_721);
and U1793 (N_1793,In_358,In_262);
or U1794 (N_1794,In_364,In_706);
nor U1795 (N_1795,In_540,In_802);
xnor U1796 (N_1796,In_130,In_156);
xor U1797 (N_1797,In_396,In_238);
xnor U1798 (N_1798,In_339,In_254);
xnor U1799 (N_1799,In_25,In_621);
or U1800 (N_1800,In_693,In_752);
nand U1801 (N_1801,In_256,In_412);
nor U1802 (N_1802,In_447,In_852);
xor U1803 (N_1803,In_876,In_570);
nand U1804 (N_1804,In_19,In_408);
xor U1805 (N_1805,In_532,In_931);
or U1806 (N_1806,In_757,In_890);
or U1807 (N_1807,In_624,In_587);
and U1808 (N_1808,In_213,In_783);
or U1809 (N_1809,In_198,In_893);
and U1810 (N_1810,In_925,In_888);
and U1811 (N_1811,In_934,In_174);
and U1812 (N_1812,In_221,In_86);
xor U1813 (N_1813,In_287,In_838);
nand U1814 (N_1814,In_132,In_862);
and U1815 (N_1815,In_963,In_770);
nand U1816 (N_1816,In_501,In_400);
or U1817 (N_1817,In_381,In_765);
xnor U1818 (N_1818,In_810,In_882);
or U1819 (N_1819,In_245,In_338);
xor U1820 (N_1820,In_199,In_862);
nand U1821 (N_1821,In_808,In_478);
nor U1822 (N_1822,In_299,In_669);
xor U1823 (N_1823,In_19,In_926);
nand U1824 (N_1824,In_152,In_301);
or U1825 (N_1825,In_68,In_876);
nor U1826 (N_1826,In_815,In_584);
xor U1827 (N_1827,In_95,In_375);
nand U1828 (N_1828,In_261,In_514);
xor U1829 (N_1829,In_973,In_706);
or U1830 (N_1830,In_837,In_45);
nor U1831 (N_1831,In_299,In_381);
and U1832 (N_1832,In_513,In_752);
xnor U1833 (N_1833,In_209,In_813);
xor U1834 (N_1834,In_18,In_466);
and U1835 (N_1835,In_357,In_576);
and U1836 (N_1836,In_330,In_179);
nor U1837 (N_1837,In_793,In_262);
nor U1838 (N_1838,In_171,In_826);
nor U1839 (N_1839,In_20,In_502);
and U1840 (N_1840,In_530,In_966);
or U1841 (N_1841,In_771,In_394);
nor U1842 (N_1842,In_211,In_776);
xor U1843 (N_1843,In_308,In_527);
and U1844 (N_1844,In_663,In_812);
nand U1845 (N_1845,In_553,In_573);
nor U1846 (N_1846,In_68,In_981);
nand U1847 (N_1847,In_729,In_470);
xor U1848 (N_1848,In_84,In_574);
and U1849 (N_1849,In_66,In_986);
xor U1850 (N_1850,In_411,In_705);
xnor U1851 (N_1851,In_920,In_887);
xnor U1852 (N_1852,In_424,In_208);
xnor U1853 (N_1853,In_69,In_145);
or U1854 (N_1854,In_981,In_594);
nand U1855 (N_1855,In_620,In_997);
xor U1856 (N_1856,In_472,In_338);
xnor U1857 (N_1857,In_166,In_438);
nand U1858 (N_1858,In_870,In_777);
nor U1859 (N_1859,In_678,In_710);
and U1860 (N_1860,In_379,In_719);
and U1861 (N_1861,In_433,In_64);
nor U1862 (N_1862,In_330,In_219);
nor U1863 (N_1863,In_7,In_514);
nor U1864 (N_1864,In_719,In_638);
nor U1865 (N_1865,In_815,In_841);
and U1866 (N_1866,In_254,In_640);
nor U1867 (N_1867,In_112,In_778);
and U1868 (N_1868,In_16,In_22);
and U1869 (N_1869,In_580,In_712);
or U1870 (N_1870,In_945,In_15);
nor U1871 (N_1871,In_263,In_494);
or U1872 (N_1872,In_622,In_191);
xor U1873 (N_1873,In_209,In_260);
or U1874 (N_1874,In_613,In_893);
or U1875 (N_1875,In_257,In_884);
and U1876 (N_1876,In_968,In_646);
xor U1877 (N_1877,In_658,In_672);
nor U1878 (N_1878,In_371,In_530);
nand U1879 (N_1879,In_517,In_526);
nand U1880 (N_1880,In_699,In_570);
nor U1881 (N_1881,In_693,In_385);
or U1882 (N_1882,In_412,In_173);
and U1883 (N_1883,In_843,In_825);
and U1884 (N_1884,In_822,In_218);
or U1885 (N_1885,In_104,In_237);
and U1886 (N_1886,In_182,In_772);
and U1887 (N_1887,In_206,In_258);
nor U1888 (N_1888,In_14,In_422);
xnor U1889 (N_1889,In_891,In_586);
and U1890 (N_1890,In_752,In_639);
nand U1891 (N_1891,In_117,In_28);
nor U1892 (N_1892,In_492,In_69);
nand U1893 (N_1893,In_665,In_512);
nor U1894 (N_1894,In_455,In_200);
xnor U1895 (N_1895,In_247,In_807);
or U1896 (N_1896,In_347,In_372);
and U1897 (N_1897,In_532,In_607);
or U1898 (N_1898,In_872,In_783);
and U1899 (N_1899,In_704,In_468);
nand U1900 (N_1900,In_629,In_666);
or U1901 (N_1901,In_242,In_77);
nand U1902 (N_1902,In_383,In_176);
and U1903 (N_1903,In_106,In_389);
and U1904 (N_1904,In_323,In_57);
xnor U1905 (N_1905,In_661,In_576);
xnor U1906 (N_1906,In_783,In_607);
or U1907 (N_1907,In_16,In_95);
nor U1908 (N_1908,In_675,In_650);
nand U1909 (N_1909,In_369,In_670);
and U1910 (N_1910,In_866,In_660);
nand U1911 (N_1911,In_697,In_281);
nand U1912 (N_1912,In_381,In_598);
and U1913 (N_1913,In_643,In_884);
xnor U1914 (N_1914,In_688,In_757);
or U1915 (N_1915,In_413,In_181);
and U1916 (N_1916,In_654,In_172);
xnor U1917 (N_1917,In_983,In_55);
or U1918 (N_1918,In_303,In_685);
nand U1919 (N_1919,In_863,In_352);
nand U1920 (N_1920,In_640,In_462);
xor U1921 (N_1921,In_377,In_259);
nor U1922 (N_1922,In_254,In_391);
nor U1923 (N_1923,In_720,In_636);
nor U1924 (N_1924,In_491,In_429);
or U1925 (N_1925,In_602,In_40);
or U1926 (N_1926,In_87,In_38);
or U1927 (N_1927,In_589,In_135);
and U1928 (N_1928,In_284,In_488);
nor U1929 (N_1929,In_822,In_761);
nor U1930 (N_1930,In_524,In_373);
and U1931 (N_1931,In_799,In_451);
and U1932 (N_1932,In_301,In_759);
nor U1933 (N_1933,In_551,In_477);
or U1934 (N_1934,In_23,In_106);
xor U1935 (N_1935,In_708,In_71);
and U1936 (N_1936,In_621,In_590);
and U1937 (N_1937,In_926,In_571);
and U1938 (N_1938,In_615,In_135);
and U1939 (N_1939,In_471,In_307);
and U1940 (N_1940,In_299,In_779);
or U1941 (N_1941,In_243,In_85);
nor U1942 (N_1942,In_832,In_906);
and U1943 (N_1943,In_830,In_275);
and U1944 (N_1944,In_883,In_821);
nand U1945 (N_1945,In_795,In_793);
and U1946 (N_1946,In_41,In_244);
and U1947 (N_1947,In_565,In_708);
nand U1948 (N_1948,In_950,In_497);
nand U1949 (N_1949,In_340,In_913);
and U1950 (N_1950,In_591,In_6);
and U1951 (N_1951,In_772,In_144);
and U1952 (N_1952,In_313,In_461);
xnor U1953 (N_1953,In_973,In_644);
or U1954 (N_1954,In_529,In_56);
nor U1955 (N_1955,In_3,In_461);
and U1956 (N_1956,In_34,In_818);
xnor U1957 (N_1957,In_78,In_838);
nor U1958 (N_1958,In_288,In_111);
or U1959 (N_1959,In_908,In_26);
and U1960 (N_1960,In_706,In_213);
xnor U1961 (N_1961,In_342,In_408);
nand U1962 (N_1962,In_506,In_688);
nand U1963 (N_1963,In_820,In_325);
xnor U1964 (N_1964,In_418,In_802);
nor U1965 (N_1965,In_920,In_30);
or U1966 (N_1966,In_454,In_871);
or U1967 (N_1967,In_551,In_69);
nor U1968 (N_1968,In_798,In_23);
nor U1969 (N_1969,In_151,In_125);
nand U1970 (N_1970,In_960,In_109);
or U1971 (N_1971,In_304,In_67);
xor U1972 (N_1972,In_799,In_606);
nand U1973 (N_1973,In_288,In_536);
nor U1974 (N_1974,In_827,In_296);
xor U1975 (N_1975,In_680,In_894);
xor U1976 (N_1976,In_656,In_120);
and U1977 (N_1977,In_491,In_94);
or U1978 (N_1978,In_880,In_635);
nand U1979 (N_1979,In_253,In_100);
xnor U1980 (N_1980,In_680,In_974);
nor U1981 (N_1981,In_602,In_95);
nor U1982 (N_1982,In_497,In_285);
or U1983 (N_1983,In_528,In_476);
nand U1984 (N_1984,In_296,In_33);
or U1985 (N_1985,In_44,In_31);
xnor U1986 (N_1986,In_996,In_929);
nand U1987 (N_1987,In_706,In_38);
nand U1988 (N_1988,In_447,In_400);
nor U1989 (N_1989,In_803,In_187);
nand U1990 (N_1990,In_993,In_88);
or U1991 (N_1991,In_25,In_154);
nor U1992 (N_1992,In_138,In_421);
and U1993 (N_1993,In_740,In_350);
and U1994 (N_1994,In_11,In_603);
xnor U1995 (N_1995,In_380,In_376);
and U1996 (N_1996,In_472,In_139);
and U1997 (N_1997,In_945,In_795);
xnor U1998 (N_1998,In_538,In_398);
nand U1999 (N_1999,In_252,In_254);
or U2000 (N_2000,In_672,In_256);
and U2001 (N_2001,In_942,In_849);
nand U2002 (N_2002,In_254,In_192);
xnor U2003 (N_2003,In_412,In_751);
nand U2004 (N_2004,In_453,In_576);
nand U2005 (N_2005,In_657,In_154);
nand U2006 (N_2006,In_976,In_406);
xor U2007 (N_2007,In_242,In_869);
xnor U2008 (N_2008,In_505,In_708);
nor U2009 (N_2009,In_527,In_633);
or U2010 (N_2010,In_791,In_195);
and U2011 (N_2011,In_852,In_144);
xnor U2012 (N_2012,In_213,In_864);
and U2013 (N_2013,In_336,In_754);
or U2014 (N_2014,In_817,In_179);
or U2015 (N_2015,In_542,In_566);
xnor U2016 (N_2016,In_180,In_101);
nor U2017 (N_2017,In_985,In_655);
or U2018 (N_2018,In_378,In_476);
and U2019 (N_2019,In_173,In_375);
xor U2020 (N_2020,In_674,In_814);
nor U2021 (N_2021,In_756,In_215);
nand U2022 (N_2022,In_735,In_368);
or U2023 (N_2023,In_237,In_513);
and U2024 (N_2024,In_246,In_114);
nor U2025 (N_2025,In_60,In_734);
nand U2026 (N_2026,In_785,In_814);
or U2027 (N_2027,In_735,In_575);
xnor U2028 (N_2028,In_673,In_447);
xor U2029 (N_2029,In_914,In_658);
nand U2030 (N_2030,In_677,In_556);
xor U2031 (N_2031,In_340,In_362);
and U2032 (N_2032,In_745,In_785);
xnor U2033 (N_2033,In_340,In_686);
nand U2034 (N_2034,In_917,In_388);
or U2035 (N_2035,In_646,In_647);
nor U2036 (N_2036,In_367,In_984);
and U2037 (N_2037,In_986,In_513);
nor U2038 (N_2038,In_593,In_214);
nand U2039 (N_2039,In_492,In_417);
nand U2040 (N_2040,In_90,In_597);
nor U2041 (N_2041,In_833,In_169);
and U2042 (N_2042,In_194,In_763);
nand U2043 (N_2043,In_940,In_262);
xor U2044 (N_2044,In_912,In_641);
xor U2045 (N_2045,In_50,In_484);
or U2046 (N_2046,In_501,In_766);
nor U2047 (N_2047,In_710,In_733);
xnor U2048 (N_2048,In_617,In_161);
or U2049 (N_2049,In_643,In_415);
and U2050 (N_2050,In_54,In_533);
nor U2051 (N_2051,In_578,In_444);
or U2052 (N_2052,In_386,In_372);
nor U2053 (N_2053,In_1,In_840);
and U2054 (N_2054,In_265,In_286);
nor U2055 (N_2055,In_480,In_681);
or U2056 (N_2056,In_446,In_390);
or U2057 (N_2057,In_84,In_567);
or U2058 (N_2058,In_267,In_174);
or U2059 (N_2059,In_55,In_424);
or U2060 (N_2060,In_698,In_86);
or U2061 (N_2061,In_79,In_282);
nor U2062 (N_2062,In_388,In_891);
xor U2063 (N_2063,In_605,In_851);
or U2064 (N_2064,In_943,In_917);
or U2065 (N_2065,In_623,In_264);
and U2066 (N_2066,In_936,In_64);
xnor U2067 (N_2067,In_827,In_179);
nand U2068 (N_2068,In_322,In_879);
xnor U2069 (N_2069,In_858,In_762);
and U2070 (N_2070,In_856,In_250);
nand U2071 (N_2071,In_873,In_615);
or U2072 (N_2072,In_386,In_608);
or U2073 (N_2073,In_7,In_161);
or U2074 (N_2074,In_406,In_79);
nand U2075 (N_2075,In_122,In_908);
nand U2076 (N_2076,In_37,In_163);
nand U2077 (N_2077,In_654,In_870);
or U2078 (N_2078,In_381,In_155);
and U2079 (N_2079,In_612,In_311);
xnor U2080 (N_2080,In_743,In_487);
nand U2081 (N_2081,In_402,In_809);
and U2082 (N_2082,In_350,In_573);
and U2083 (N_2083,In_256,In_382);
and U2084 (N_2084,In_94,In_546);
xnor U2085 (N_2085,In_513,In_157);
or U2086 (N_2086,In_868,In_172);
nand U2087 (N_2087,In_134,In_855);
xor U2088 (N_2088,In_253,In_451);
or U2089 (N_2089,In_350,In_528);
nand U2090 (N_2090,In_681,In_810);
or U2091 (N_2091,In_150,In_168);
nor U2092 (N_2092,In_195,In_388);
nand U2093 (N_2093,In_159,In_909);
and U2094 (N_2094,In_275,In_350);
nor U2095 (N_2095,In_647,In_482);
nor U2096 (N_2096,In_816,In_709);
or U2097 (N_2097,In_533,In_151);
xor U2098 (N_2098,In_107,In_652);
and U2099 (N_2099,In_669,In_80);
and U2100 (N_2100,In_792,In_141);
xnor U2101 (N_2101,In_155,In_555);
xor U2102 (N_2102,In_277,In_545);
nor U2103 (N_2103,In_858,In_466);
and U2104 (N_2104,In_584,In_403);
and U2105 (N_2105,In_464,In_366);
nor U2106 (N_2106,In_282,In_200);
nand U2107 (N_2107,In_598,In_946);
nand U2108 (N_2108,In_23,In_50);
nor U2109 (N_2109,In_882,In_480);
or U2110 (N_2110,In_102,In_296);
and U2111 (N_2111,In_691,In_788);
xor U2112 (N_2112,In_606,In_831);
or U2113 (N_2113,In_13,In_142);
or U2114 (N_2114,In_690,In_92);
xor U2115 (N_2115,In_132,In_895);
nand U2116 (N_2116,In_469,In_870);
nor U2117 (N_2117,In_830,In_593);
xnor U2118 (N_2118,In_131,In_62);
or U2119 (N_2119,In_79,In_741);
nand U2120 (N_2120,In_765,In_414);
xor U2121 (N_2121,In_458,In_305);
or U2122 (N_2122,In_440,In_538);
nand U2123 (N_2123,In_3,In_139);
xor U2124 (N_2124,In_248,In_293);
nand U2125 (N_2125,In_892,In_487);
nor U2126 (N_2126,In_966,In_802);
nor U2127 (N_2127,In_345,In_139);
and U2128 (N_2128,In_58,In_435);
nand U2129 (N_2129,In_922,In_473);
and U2130 (N_2130,In_683,In_337);
nand U2131 (N_2131,In_101,In_912);
nand U2132 (N_2132,In_394,In_119);
or U2133 (N_2133,In_461,In_167);
or U2134 (N_2134,In_463,In_136);
or U2135 (N_2135,In_106,In_242);
nand U2136 (N_2136,In_598,In_12);
and U2137 (N_2137,In_718,In_467);
xnor U2138 (N_2138,In_276,In_752);
nand U2139 (N_2139,In_803,In_756);
nor U2140 (N_2140,In_551,In_839);
xnor U2141 (N_2141,In_157,In_945);
nor U2142 (N_2142,In_10,In_751);
or U2143 (N_2143,In_95,In_682);
nand U2144 (N_2144,In_625,In_165);
or U2145 (N_2145,In_170,In_808);
nand U2146 (N_2146,In_213,In_80);
nand U2147 (N_2147,In_712,In_238);
nor U2148 (N_2148,In_301,In_736);
and U2149 (N_2149,In_155,In_976);
or U2150 (N_2150,In_178,In_703);
nor U2151 (N_2151,In_372,In_487);
nor U2152 (N_2152,In_999,In_869);
or U2153 (N_2153,In_133,In_874);
and U2154 (N_2154,In_223,In_282);
nor U2155 (N_2155,In_270,In_998);
xor U2156 (N_2156,In_781,In_155);
nor U2157 (N_2157,In_770,In_225);
nor U2158 (N_2158,In_758,In_896);
xor U2159 (N_2159,In_377,In_756);
nor U2160 (N_2160,In_173,In_134);
and U2161 (N_2161,In_897,In_452);
and U2162 (N_2162,In_778,In_34);
nor U2163 (N_2163,In_222,In_795);
and U2164 (N_2164,In_714,In_222);
nand U2165 (N_2165,In_679,In_824);
nand U2166 (N_2166,In_233,In_573);
xnor U2167 (N_2167,In_164,In_741);
and U2168 (N_2168,In_978,In_162);
or U2169 (N_2169,In_470,In_256);
nor U2170 (N_2170,In_856,In_845);
or U2171 (N_2171,In_206,In_415);
and U2172 (N_2172,In_545,In_798);
nand U2173 (N_2173,In_1,In_726);
nand U2174 (N_2174,In_10,In_908);
xnor U2175 (N_2175,In_222,In_615);
or U2176 (N_2176,In_820,In_551);
nor U2177 (N_2177,In_661,In_701);
or U2178 (N_2178,In_74,In_522);
and U2179 (N_2179,In_212,In_618);
and U2180 (N_2180,In_361,In_467);
nor U2181 (N_2181,In_933,In_958);
or U2182 (N_2182,In_311,In_42);
nor U2183 (N_2183,In_654,In_989);
or U2184 (N_2184,In_165,In_879);
nand U2185 (N_2185,In_169,In_559);
nor U2186 (N_2186,In_393,In_976);
nand U2187 (N_2187,In_6,In_984);
and U2188 (N_2188,In_213,In_888);
nand U2189 (N_2189,In_674,In_274);
or U2190 (N_2190,In_862,In_875);
nand U2191 (N_2191,In_334,In_862);
and U2192 (N_2192,In_4,In_835);
or U2193 (N_2193,In_402,In_265);
and U2194 (N_2194,In_101,In_4);
or U2195 (N_2195,In_524,In_779);
nand U2196 (N_2196,In_987,In_296);
nand U2197 (N_2197,In_648,In_896);
and U2198 (N_2198,In_694,In_135);
and U2199 (N_2199,In_21,In_434);
xnor U2200 (N_2200,In_92,In_233);
xnor U2201 (N_2201,In_510,In_259);
nand U2202 (N_2202,In_431,In_866);
xnor U2203 (N_2203,In_98,In_9);
nand U2204 (N_2204,In_866,In_109);
or U2205 (N_2205,In_427,In_844);
or U2206 (N_2206,In_583,In_773);
nand U2207 (N_2207,In_566,In_120);
nor U2208 (N_2208,In_880,In_911);
or U2209 (N_2209,In_643,In_632);
nand U2210 (N_2210,In_931,In_149);
nand U2211 (N_2211,In_949,In_828);
or U2212 (N_2212,In_894,In_431);
or U2213 (N_2213,In_823,In_136);
or U2214 (N_2214,In_374,In_477);
or U2215 (N_2215,In_959,In_126);
nand U2216 (N_2216,In_797,In_529);
nor U2217 (N_2217,In_363,In_383);
nor U2218 (N_2218,In_864,In_483);
nor U2219 (N_2219,In_54,In_634);
or U2220 (N_2220,In_811,In_623);
and U2221 (N_2221,In_66,In_305);
nor U2222 (N_2222,In_941,In_606);
xor U2223 (N_2223,In_921,In_168);
nor U2224 (N_2224,In_142,In_935);
xor U2225 (N_2225,In_689,In_2);
and U2226 (N_2226,In_224,In_179);
nand U2227 (N_2227,In_688,In_59);
xor U2228 (N_2228,In_506,In_586);
nand U2229 (N_2229,In_142,In_587);
and U2230 (N_2230,In_222,In_46);
nor U2231 (N_2231,In_775,In_29);
xor U2232 (N_2232,In_396,In_505);
xor U2233 (N_2233,In_534,In_886);
and U2234 (N_2234,In_644,In_276);
and U2235 (N_2235,In_999,In_147);
nand U2236 (N_2236,In_661,In_745);
nand U2237 (N_2237,In_793,In_487);
nor U2238 (N_2238,In_346,In_572);
or U2239 (N_2239,In_543,In_346);
and U2240 (N_2240,In_332,In_779);
and U2241 (N_2241,In_243,In_526);
nand U2242 (N_2242,In_933,In_30);
nand U2243 (N_2243,In_122,In_883);
and U2244 (N_2244,In_374,In_754);
and U2245 (N_2245,In_458,In_888);
nor U2246 (N_2246,In_140,In_404);
nor U2247 (N_2247,In_374,In_668);
nor U2248 (N_2248,In_320,In_929);
xor U2249 (N_2249,In_251,In_389);
and U2250 (N_2250,In_657,In_854);
and U2251 (N_2251,In_945,In_814);
nand U2252 (N_2252,In_963,In_303);
nand U2253 (N_2253,In_4,In_347);
nor U2254 (N_2254,In_965,In_189);
nor U2255 (N_2255,In_828,In_780);
or U2256 (N_2256,In_848,In_137);
or U2257 (N_2257,In_245,In_538);
or U2258 (N_2258,In_46,In_825);
xor U2259 (N_2259,In_841,In_757);
nor U2260 (N_2260,In_501,In_494);
nor U2261 (N_2261,In_89,In_368);
and U2262 (N_2262,In_478,In_736);
nor U2263 (N_2263,In_166,In_881);
and U2264 (N_2264,In_864,In_251);
xnor U2265 (N_2265,In_150,In_328);
and U2266 (N_2266,In_739,In_988);
nor U2267 (N_2267,In_741,In_569);
and U2268 (N_2268,In_883,In_920);
or U2269 (N_2269,In_983,In_629);
and U2270 (N_2270,In_832,In_754);
nor U2271 (N_2271,In_662,In_934);
and U2272 (N_2272,In_873,In_947);
nand U2273 (N_2273,In_676,In_462);
nor U2274 (N_2274,In_128,In_431);
and U2275 (N_2275,In_564,In_9);
or U2276 (N_2276,In_279,In_523);
xor U2277 (N_2277,In_115,In_962);
or U2278 (N_2278,In_747,In_647);
or U2279 (N_2279,In_912,In_612);
and U2280 (N_2280,In_149,In_209);
and U2281 (N_2281,In_552,In_286);
xor U2282 (N_2282,In_326,In_429);
nand U2283 (N_2283,In_883,In_440);
nand U2284 (N_2284,In_379,In_936);
nand U2285 (N_2285,In_623,In_397);
nand U2286 (N_2286,In_244,In_845);
xnor U2287 (N_2287,In_603,In_844);
nand U2288 (N_2288,In_620,In_74);
nand U2289 (N_2289,In_1,In_718);
or U2290 (N_2290,In_656,In_825);
nor U2291 (N_2291,In_129,In_890);
nand U2292 (N_2292,In_775,In_117);
or U2293 (N_2293,In_287,In_806);
or U2294 (N_2294,In_852,In_691);
nand U2295 (N_2295,In_495,In_455);
and U2296 (N_2296,In_430,In_658);
nand U2297 (N_2297,In_24,In_924);
or U2298 (N_2298,In_692,In_969);
xnor U2299 (N_2299,In_459,In_90);
nand U2300 (N_2300,In_715,In_969);
nor U2301 (N_2301,In_657,In_846);
or U2302 (N_2302,In_718,In_704);
nand U2303 (N_2303,In_244,In_644);
xnor U2304 (N_2304,In_993,In_6);
nor U2305 (N_2305,In_58,In_852);
and U2306 (N_2306,In_974,In_270);
nand U2307 (N_2307,In_458,In_423);
xnor U2308 (N_2308,In_785,In_743);
nand U2309 (N_2309,In_625,In_127);
nand U2310 (N_2310,In_452,In_15);
and U2311 (N_2311,In_832,In_420);
xor U2312 (N_2312,In_48,In_772);
nor U2313 (N_2313,In_989,In_751);
nand U2314 (N_2314,In_24,In_484);
and U2315 (N_2315,In_131,In_92);
or U2316 (N_2316,In_468,In_577);
or U2317 (N_2317,In_644,In_910);
nand U2318 (N_2318,In_73,In_28);
xnor U2319 (N_2319,In_675,In_559);
nor U2320 (N_2320,In_331,In_533);
and U2321 (N_2321,In_252,In_803);
nor U2322 (N_2322,In_490,In_720);
nor U2323 (N_2323,In_642,In_354);
nor U2324 (N_2324,In_220,In_751);
xnor U2325 (N_2325,In_650,In_162);
or U2326 (N_2326,In_271,In_418);
or U2327 (N_2327,In_617,In_802);
xnor U2328 (N_2328,In_697,In_335);
and U2329 (N_2329,In_278,In_982);
or U2330 (N_2330,In_716,In_27);
and U2331 (N_2331,In_982,In_385);
nor U2332 (N_2332,In_33,In_706);
xor U2333 (N_2333,In_502,In_706);
and U2334 (N_2334,In_540,In_508);
nand U2335 (N_2335,In_893,In_103);
and U2336 (N_2336,In_246,In_355);
nand U2337 (N_2337,In_884,In_717);
nand U2338 (N_2338,In_621,In_727);
nand U2339 (N_2339,In_57,In_880);
and U2340 (N_2340,In_588,In_441);
or U2341 (N_2341,In_638,In_366);
nor U2342 (N_2342,In_959,In_109);
nor U2343 (N_2343,In_527,In_26);
and U2344 (N_2344,In_461,In_102);
nor U2345 (N_2345,In_574,In_568);
or U2346 (N_2346,In_104,In_204);
and U2347 (N_2347,In_825,In_980);
xor U2348 (N_2348,In_954,In_989);
or U2349 (N_2349,In_946,In_789);
and U2350 (N_2350,In_187,In_522);
nand U2351 (N_2351,In_807,In_928);
nor U2352 (N_2352,In_751,In_369);
nand U2353 (N_2353,In_849,In_230);
xor U2354 (N_2354,In_717,In_692);
xor U2355 (N_2355,In_846,In_461);
xor U2356 (N_2356,In_509,In_838);
nor U2357 (N_2357,In_912,In_449);
xnor U2358 (N_2358,In_507,In_296);
and U2359 (N_2359,In_800,In_703);
nor U2360 (N_2360,In_244,In_739);
nand U2361 (N_2361,In_829,In_652);
xor U2362 (N_2362,In_475,In_650);
or U2363 (N_2363,In_122,In_769);
nor U2364 (N_2364,In_47,In_48);
nand U2365 (N_2365,In_759,In_715);
nand U2366 (N_2366,In_318,In_310);
and U2367 (N_2367,In_149,In_725);
nand U2368 (N_2368,In_559,In_270);
and U2369 (N_2369,In_130,In_439);
nor U2370 (N_2370,In_406,In_606);
nor U2371 (N_2371,In_44,In_735);
nor U2372 (N_2372,In_38,In_187);
and U2373 (N_2373,In_964,In_19);
or U2374 (N_2374,In_994,In_867);
and U2375 (N_2375,In_145,In_304);
and U2376 (N_2376,In_582,In_376);
and U2377 (N_2377,In_620,In_661);
nand U2378 (N_2378,In_376,In_950);
and U2379 (N_2379,In_61,In_268);
xor U2380 (N_2380,In_654,In_317);
nor U2381 (N_2381,In_112,In_188);
nor U2382 (N_2382,In_768,In_302);
and U2383 (N_2383,In_741,In_52);
or U2384 (N_2384,In_437,In_519);
and U2385 (N_2385,In_429,In_291);
and U2386 (N_2386,In_531,In_592);
nor U2387 (N_2387,In_742,In_705);
xor U2388 (N_2388,In_811,In_299);
or U2389 (N_2389,In_460,In_694);
nor U2390 (N_2390,In_785,In_45);
xor U2391 (N_2391,In_46,In_804);
or U2392 (N_2392,In_754,In_134);
nor U2393 (N_2393,In_233,In_158);
or U2394 (N_2394,In_745,In_186);
nor U2395 (N_2395,In_270,In_831);
xor U2396 (N_2396,In_545,In_158);
xor U2397 (N_2397,In_97,In_417);
nand U2398 (N_2398,In_961,In_364);
nor U2399 (N_2399,In_404,In_457);
nand U2400 (N_2400,In_7,In_145);
nor U2401 (N_2401,In_966,In_157);
and U2402 (N_2402,In_999,In_959);
nand U2403 (N_2403,In_753,In_698);
nand U2404 (N_2404,In_184,In_580);
or U2405 (N_2405,In_98,In_289);
or U2406 (N_2406,In_463,In_77);
or U2407 (N_2407,In_364,In_354);
or U2408 (N_2408,In_659,In_593);
or U2409 (N_2409,In_695,In_963);
and U2410 (N_2410,In_300,In_278);
and U2411 (N_2411,In_617,In_922);
and U2412 (N_2412,In_802,In_157);
nand U2413 (N_2413,In_317,In_918);
nor U2414 (N_2414,In_755,In_390);
xnor U2415 (N_2415,In_182,In_250);
and U2416 (N_2416,In_422,In_97);
and U2417 (N_2417,In_849,In_63);
nor U2418 (N_2418,In_333,In_804);
and U2419 (N_2419,In_426,In_270);
or U2420 (N_2420,In_925,In_583);
nand U2421 (N_2421,In_768,In_675);
xnor U2422 (N_2422,In_629,In_282);
nor U2423 (N_2423,In_587,In_948);
nand U2424 (N_2424,In_273,In_804);
or U2425 (N_2425,In_192,In_624);
or U2426 (N_2426,In_259,In_260);
xnor U2427 (N_2427,In_186,In_172);
nor U2428 (N_2428,In_721,In_136);
and U2429 (N_2429,In_742,In_692);
nor U2430 (N_2430,In_637,In_103);
nand U2431 (N_2431,In_198,In_516);
xnor U2432 (N_2432,In_587,In_469);
or U2433 (N_2433,In_288,In_971);
nor U2434 (N_2434,In_332,In_334);
or U2435 (N_2435,In_656,In_805);
nand U2436 (N_2436,In_967,In_99);
xnor U2437 (N_2437,In_522,In_342);
and U2438 (N_2438,In_793,In_925);
or U2439 (N_2439,In_327,In_180);
nand U2440 (N_2440,In_226,In_681);
and U2441 (N_2441,In_514,In_672);
nand U2442 (N_2442,In_939,In_168);
or U2443 (N_2443,In_325,In_749);
and U2444 (N_2444,In_189,In_242);
nor U2445 (N_2445,In_237,In_16);
and U2446 (N_2446,In_498,In_225);
nor U2447 (N_2447,In_281,In_501);
nand U2448 (N_2448,In_515,In_663);
nor U2449 (N_2449,In_120,In_509);
or U2450 (N_2450,In_303,In_585);
nor U2451 (N_2451,In_588,In_332);
nand U2452 (N_2452,In_503,In_161);
or U2453 (N_2453,In_746,In_37);
xnor U2454 (N_2454,In_365,In_321);
or U2455 (N_2455,In_96,In_947);
and U2456 (N_2456,In_69,In_880);
nor U2457 (N_2457,In_61,In_857);
nor U2458 (N_2458,In_161,In_983);
nor U2459 (N_2459,In_222,In_442);
xor U2460 (N_2460,In_889,In_494);
nor U2461 (N_2461,In_987,In_825);
nand U2462 (N_2462,In_126,In_941);
nand U2463 (N_2463,In_444,In_295);
and U2464 (N_2464,In_208,In_713);
nor U2465 (N_2465,In_605,In_34);
nor U2466 (N_2466,In_983,In_301);
nand U2467 (N_2467,In_979,In_783);
and U2468 (N_2468,In_382,In_501);
or U2469 (N_2469,In_382,In_282);
nor U2470 (N_2470,In_625,In_261);
and U2471 (N_2471,In_186,In_738);
or U2472 (N_2472,In_771,In_499);
nor U2473 (N_2473,In_14,In_104);
nand U2474 (N_2474,In_458,In_11);
xor U2475 (N_2475,In_631,In_885);
or U2476 (N_2476,In_190,In_861);
nand U2477 (N_2477,In_672,In_425);
or U2478 (N_2478,In_262,In_347);
nor U2479 (N_2479,In_471,In_778);
xnor U2480 (N_2480,In_67,In_409);
and U2481 (N_2481,In_944,In_602);
nand U2482 (N_2482,In_252,In_895);
nor U2483 (N_2483,In_111,In_930);
xnor U2484 (N_2484,In_552,In_752);
nand U2485 (N_2485,In_553,In_292);
nand U2486 (N_2486,In_237,In_23);
nor U2487 (N_2487,In_585,In_525);
nand U2488 (N_2488,In_568,In_358);
xor U2489 (N_2489,In_738,In_319);
nor U2490 (N_2490,In_610,In_523);
and U2491 (N_2491,In_864,In_664);
xor U2492 (N_2492,In_968,In_856);
nor U2493 (N_2493,In_123,In_626);
xnor U2494 (N_2494,In_878,In_152);
or U2495 (N_2495,In_827,In_640);
and U2496 (N_2496,In_813,In_101);
nand U2497 (N_2497,In_651,In_387);
and U2498 (N_2498,In_661,In_868);
or U2499 (N_2499,In_182,In_734);
and U2500 (N_2500,In_812,In_40);
or U2501 (N_2501,In_616,In_593);
xnor U2502 (N_2502,In_889,In_692);
and U2503 (N_2503,In_310,In_876);
nand U2504 (N_2504,In_933,In_1);
xor U2505 (N_2505,In_985,In_739);
nor U2506 (N_2506,In_508,In_263);
nor U2507 (N_2507,In_70,In_558);
nor U2508 (N_2508,In_474,In_349);
xnor U2509 (N_2509,In_188,In_385);
xor U2510 (N_2510,In_671,In_52);
and U2511 (N_2511,In_232,In_934);
xor U2512 (N_2512,In_668,In_179);
nand U2513 (N_2513,In_461,In_257);
xor U2514 (N_2514,In_944,In_354);
or U2515 (N_2515,In_909,In_65);
and U2516 (N_2516,In_779,In_236);
nand U2517 (N_2517,In_740,In_733);
or U2518 (N_2518,In_68,In_39);
nor U2519 (N_2519,In_348,In_946);
or U2520 (N_2520,In_235,In_182);
xnor U2521 (N_2521,In_36,In_826);
xor U2522 (N_2522,In_806,In_107);
nand U2523 (N_2523,In_780,In_892);
or U2524 (N_2524,In_288,In_151);
nand U2525 (N_2525,In_214,In_914);
nor U2526 (N_2526,In_613,In_225);
xor U2527 (N_2527,In_345,In_941);
and U2528 (N_2528,In_578,In_240);
nand U2529 (N_2529,In_118,In_372);
nor U2530 (N_2530,In_770,In_337);
nand U2531 (N_2531,In_582,In_549);
and U2532 (N_2532,In_323,In_363);
xor U2533 (N_2533,In_590,In_138);
xnor U2534 (N_2534,In_706,In_612);
and U2535 (N_2535,In_664,In_167);
or U2536 (N_2536,In_297,In_527);
or U2537 (N_2537,In_350,In_945);
xnor U2538 (N_2538,In_4,In_629);
nand U2539 (N_2539,In_631,In_66);
and U2540 (N_2540,In_936,In_909);
xor U2541 (N_2541,In_453,In_20);
nand U2542 (N_2542,In_443,In_288);
xnor U2543 (N_2543,In_686,In_285);
or U2544 (N_2544,In_726,In_535);
and U2545 (N_2545,In_138,In_210);
and U2546 (N_2546,In_330,In_315);
or U2547 (N_2547,In_454,In_891);
xor U2548 (N_2548,In_389,In_429);
nand U2549 (N_2549,In_985,In_28);
or U2550 (N_2550,In_647,In_575);
or U2551 (N_2551,In_713,In_985);
nand U2552 (N_2552,In_607,In_634);
nand U2553 (N_2553,In_766,In_441);
nor U2554 (N_2554,In_881,In_164);
or U2555 (N_2555,In_584,In_214);
and U2556 (N_2556,In_221,In_410);
nand U2557 (N_2557,In_28,In_884);
xnor U2558 (N_2558,In_762,In_29);
nand U2559 (N_2559,In_993,In_821);
nor U2560 (N_2560,In_951,In_38);
nand U2561 (N_2561,In_719,In_619);
or U2562 (N_2562,In_619,In_815);
nor U2563 (N_2563,In_15,In_704);
or U2564 (N_2564,In_481,In_426);
and U2565 (N_2565,In_254,In_696);
nor U2566 (N_2566,In_384,In_771);
and U2567 (N_2567,In_438,In_411);
and U2568 (N_2568,In_532,In_411);
nand U2569 (N_2569,In_293,In_698);
or U2570 (N_2570,In_330,In_190);
nor U2571 (N_2571,In_345,In_55);
or U2572 (N_2572,In_743,In_588);
xnor U2573 (N_2573,In_619,In_79);
nand U2574 (N_2574,In_945,In_68);
xnor U2575 (N_2575,In_871,In_528);
nand U2576 (N_2576,In_486,In_809);
or U2577 (N_2577,In_890,In_431);
xor U2578 (N_2578,In_640,In_535);
or U2579 (N_2579,In_55,In_344);
nor U2580 (N_2580,In_206,In_529);
xnor U2581 (N_2581,In_975,In_737);
nor U2582 (N_2582,In_215,In_386);
nand U2583 (N_2583,In_259,In_813);
or U2584 (N_2584,In_646,In_105);
and U2585 (N_2585,In_30,In_171);
and U2586 (N_2586,In_986,In_113);
or U2587 (N_2587,In_220,In_787);
and U2588 (N_2588,In_745,In_644);
xnor U2589 (N_2589,In_343,In_41);
and U2590 (N_2590,In_461,In_154);
nand U2591 (N_2591,In_261,In_423);
nor U2592 (N_2592,In_755,In_67);
nand U2593 (N_2593,In_272,In_222);
and U2594 (N_2594,In_654,In_135);
or U2595 (N_2595,In_967,In_574);
nor U2596 (N_2596,In_357,In_891);
nor U2597 (N_2597,In_331,In_435);
nand U2598 (N_2598,In_836,In_752);
nand U2599 (N_2599,In_614,In_37);
or U2600 (N_2600,In_311,In_764);
nor U2601 (N_2601,In_811,In_593);
nand U2602 (N_2602,In_926,In_570);
nor U2603 (N_2603,In_447,In_44);
nand U2604 (N_2604,In_764,In_849);
xor U2605 (N_2605,In_929,In_39);
or U2606 (N_2606,In_549,In_569);
nor U2607 (N_2607,In_163,In_206);
xor U2608 (N_2608,In_108,In_251);
xnor U2609 (N_2609,In_872,In_489);
nor U2610 (N_2610,In_939,In_238);
nand U2611 (N_2611,In_712,In_524);
nor U2612 (N_2612,In_299,In_385);
or U2613 (N_2613,In_385,In_737);
nor U2614 (N_2614,In_46,In_83);
nor U2615 (N_2615,In_117,In_794);
nor U2616 (N_2616,In_404,In_980);
or U2617 (N_2617,In_856,In_165);
and U2618 (N_2618,In_85,In_762);
nor U2619 (N_2619,In_163,In_957);
nor U2620 (N_2620,In_523,In_763);
nand U2621 (N_2621,In_801,In_215);
or U2622 (N_2622,In_115,In_596);
nand U2623 (N_2623,In_328,In_42);
and U2624 (N_2624,In_289,In_666);
or U2625 (N_2625,In_802,In_11);
nand U2626 (N_2626,In_688,In_209);
nor U2627 (N_2627,In_395,In_913);
and U2628 (N_2628,In_58,In_366);
xnor U2629 (N_2629,In_148,In_262);
and U2630 (N_2630,In_575,In_244);
and U2631 (N_2631,In_405,In_553);
and U2632 (N_2632,In_311,In_196);
nor U2633 (N_2633,In_130,In_75);
xor U2634 (N_2634,In_852,In_278);
and U2635 (N_2635,In_541,In_764);
nor U2636 (N_2636,In_684,In_441);
and U2637 (N_2637,In_373,In_157);
nand U2638 (N_2638,In_786,In_654);
nand U2639 (N_2639,In_844,In_60);
nand U2640 (N_2640,In_676,In_931);
xor U2641 (N_2641,In_807,In_744);
or U2642 (N_2642,In_945,In_699);
nand U2643 (N_2643,In_54,In_108);
nor U2644 (N_2644,In_442,In_267);
nor U2645 (N_2645,In_880,In_336);
or U2646 (N_2646,In_169,In_623);
xor U2647 (N_2647,In_205,In_334);
nand U2648 (N_2648,In_311,In_854);
or U2649 (N_2649,In_705,In_282);
and U2650 (N_2650,In_284,In_568);
nand U2651 (N_2651,In_274,In_452);
xor U2652 (N_2652,In_964,In_70);
nand U2653 (N_2653,In_932,In_477);
nor U2654 (N_2654,In_892,In_885);
nor U2655 (N_2655,In_130,In_785);
or U2656 (N_2656,In_331,In_266);
nor U2657 (N_2657,In_178,In_99);
nand U2658 (N_2658,In_692,In_733);
nor U2659 (N_2659,In_370,In_379);
nor U2660 (N_2660,In_996,In_840);
nand U2661 (N_2661,In_452,In_875);
and U2662 (N_2662,In_584,In_216);
or U2663 (N_2663,In_585,In_566);
or U2664 (N_2664,In_574,In_279);
nand U2665 (N_2665,In_785,In_113);
and U2666 (N_2666,In_756,In_7);
xor U2667 (N_2667,In_219,In_402);
nand U2668 (N_2668,In_928,In_640);
and U2669 (N_2669,In_968,In_524);
and U2670 (N_2670,In_130,In_244);
nand U2671 (N_2671,In_134,In_652);
or U2672 (N_2672,In_295,In_290);
and U2673 (N_2673,In_633,In_54);
nand U2674 (N_2674,In_552,In_661);
and U2675 (N_2675,In_996,In_418);
xor U2676 (N_2676,In_507,In_382);
and U2677 (N_2677,In_652,In_360);
or U2678 (N_2678,In_43,In_165);
nor U2679 (N_2679,In_514,In_148);
nor U2680 (N_2680,In_97,In_477);
nor U2681 (N_2681,In_81,In_827);
and U2682 (N_2682,In_46,In_175);
nor U2683 (N_2683,In_439,In_462);
or U2684 (N_2684,In_887,In_851);
xnor U2685 (N_2685,In_891,In_30);
nor U2686 (N_2686,In_448,In_284);
and U2687 (N_2687,In_748,In_250);
and U2688 (N_2688,In_438,In_38);
xor U2689 (N_2689,In_102,In_210);
nor U2690 (N_2690,In_255,In_335);
and U2691 (N_2691,In_524,In_64);
and U2692 (N_2692,In_828,In_203);
or U2693 (N_2693,In_81,In_40);
and U2694 (N_2694,In_928,In_89);
and U2695 (N_2695,In_781,In_551);
or U2696 (N_2696,In_17,In_211);
and U2697 (N_2697,In_916,In_310);
or U2698 (N_2698,In_694,In_144);
nand U2699 (N_2699,In_41,In_142);
nand U2700 (N_2700,In_587,In_570);
xor U2701 (N_2701,In_141,In_775);
nand U2702 (N_2702,In_495,In_397);
xor U2703 (N_2703,In_992,In_794);
and U2704 (N_2704,In_387,In_614);
or U2705 (N_2705,In_74,In_443);
or U2706 (N_2706,In_612,In_732);
nand U2707 (N_2707,In_674,In_703);
or U2708 (N_2708,In_389,In_669);
or U2709 (N_2709,In_550,In_85);
or U2710 (N_2710,In_35,In_689);
nor U2711 (N_2711,In_859,In_201);
nand U2712 (N_2712,In_599,In_756);
and U2713 (N_2713,In_239,In_581);
nor U2714 (N_2714,In_784,In_236);
nor U2715 (N_2715,In_988,In_74);
and U2716 (N_2716,In_991,In_282);
nor U2717 (N_2717,In_600,In_712);
and U2718 (N_2718,In_780,In_185);
or U2719 (N_2719,In_561,In_547);
xor U2720 (N_2720,In_220,In_76);
and U2721 (N_2721,In_316,In_689);
nor U2722 (N_2722,In_627,In_847);
nand U2723 (N_2723,In_644,In_982);
nor U2724 (N_2724,In_478,In_479);
or U2725 (N_2725,In_259,In_448);
or U2726 (N_2726,In_66,In_263);
xor U2727 (N_2727,In_20,In_576);
xnor U2728 (N_2728,In_869,In_936);
xnor U2729 (N_2729,In_992,In_316);
and U2730 (N_2730,In_322,In_235);
and U2731 (N_2731,In_917,In_250);
xnor U2732 (N_2732,In_271,In_640);
xnor U2733 (N_2733,In_192,In_618);
xor U2734 (N_2734,In_79,In_588);
nor U2735 (N_2735,In_750,In_375);
and U2736 (N_2736,In_909,In_923);
or U2737 (N_2737,In_605,In_476);
xor U2738 (N_2738,In_692,In_343);
xor U2739 (N_2739,In_631,In_554);
and U2740 (N_2740,In_158,In_796);
nand U2741 (N_2741,In_262,In_835);
or U2742 (N_2742,In_67,In_249);
nand U2743 (N_2743,In_274,In_966);
and U2744 (N_2744,In_699,In_302);
or U2745 (N_2745,In_418,In_186);
or U2746 (N_2746,In_836,In_287);
or U2747 (N_2747,In_334,In_250);
xnor U2748 (N_2748,In_754,In_856);
nand U2749 (N_2749,In_983,In_685);
or U2750 (N_2750,In_83,In_459);
nor U2751 (N_2751,In_477,In_888);
or U2752 (N_2752,In_941,In_22);
nand U2753 (N_2753,In_349,In_623);
nand U2754 (N_2754,In_147,In_846);
xor U2755 (N_2755,In_887,In_55);
nor U2756 (N_2756,In_916,In_893);
and U2757 (N_2757,In_669,In_840);
xor U2758 (N_2758,In_663,In_337);
nor U2759 (N_2759,In_580,In_181);
and U2760 (N_2760,In_910,In_593);
or U2761 (N_2761,In_595,In_904);
nor U2762 (N_2762,In_556,In_723);
or U2763 (N_2763,In_500,In_189);
xor U2764 (N_2764,In_857,In_267);
nor U2765 (N_2765,In_852,In_140);
or U2766 (N_2766,In_898,In_648);
and U2767 (N_2767,In_627,In_523);
xnor U2768 (N_2768,In_98,In_273);
xor U2769 (N_2769,In_496,In_2);
nor U2770 (N_2770,In_182,In_288);
or U2771 (N_2771,In_535,In_218);
or U2772 (N_2772,In_896,In_114);
xor U2773 (N_2773,In_810,In_629);
or U2774 (N_2774,In_432,In_679);
and U2775 (N_2775,In_472,In_694);
nand U2776 (N_2776,In_484,In_397);
and U2777 (N_2777,In_287,In_876);
or U2778 (N_2778,In_205,In_336);
or U2779 (N_2779,In_164,In_486);
nand U2780 (N_2780,In_779,In_739);
xor U2781 (N_2781,In_52,In_861);
or U2782 (N_2782,In_816,In_349);
nand U2783 (N_2783,In_772,In_669);
nand U2784 (N_2784,In_304,In_164);
xnor U2785 (N_2785,In_271,In_334);
nor U2786 (N_2786,In_930,In_153);
nand U2787 (N_2787,In_636,In_224);
nor U2788 (N_2788,In_139,In_103);
nor U2789 (N_2789,In_758,In_229);
and U2790 (N_2790,In_565,In_690);
nor U2791 (N_2791,In_850,In_773);
nor U2792 (N_2792,In_937,In_178);
nor U2793 (N_2793,In_842,In_62);
and U2794 (N_2794,In_229,In_628);
or U2795 (N_2795,In_883,In_952);
or U2796 (N_2796,In_492,In_475);
and U2797 (N_2797,In_582,In_681);
nor U2798 (N_2798,In_606,In_378);
xor U2799 (N_2799,In_126,In_570);
xnor U2800 (N_2800,In_338,In_894);
nand U2801 (N_2801,In_753,In_359);
and U2802 (N_2802,In_391,In_640);
nand U2803 (N_2803,In_927,In_424);
nand U2804 (N_2804,In_974,In_593);
or U2805 (N_2805,In_98,In_608);
and U2806 (N_2806,In_555,In_227);
nor U2807 (N_2807,In_146,In_417);
xnor U2808 (N_2808,In_262,In_657);
or U2809 (N_2809,In_604,In_525);
xnor U2810 (N_2810,In_209,In_315);
nand U2811 (N_2811,In_163,In_6);
xnor U2812 (N_2812,In_321,In_843);
xnor U2813 (N_2813,In_697,In_77);
or U2814 (N_2814,In_398,In_561);
nor U2815 (N_2815,In_638,In_307);
and U2816 (N_2816,In_469,In_776);
or U2817 (N_2817,In_477,In_813);
nor U2818 (N_2818,In_799,In_332);
or U2819 (N_2819,In_481,In_433);
nor U2820 (N_2820,In_448,In_921);
nor U2821 (N_2821,In_223,In_327);
nand U2822 (N_2822,In_751,In_593);
nor U2823 (N_2823,In_113,In_86);
or U2824 (N_2824,In_193,In_941);
and U2825 (N_2825,In_503,In_743);
and U2826 (N_2826,In_446,In_486);
xor U2827 (N_2827,In_888,In_340);
nor U2828 (N_2828,In_422,In_894);
or U2829 (N_2829,In_705,In_924);
nor U2830 (N_2830,In_357,In_905);
or U2831 (N_2831,In_323,In_755);
nor U2832 (N_2832,In_305,In_657);
nor U2833 (N_2833,In_239,In_906);
or U2834 (N_2834,In_804,In_354);
xor U2835 (N_2835,In_309,In_248);
and U2836 (N_2836,In_664,In_417);
xor U2837 (N_2837,In_698,In_427);
nor U2838 (N_2838,In_133,In_894);
or U2839 (N_2839,In_22,In_27);
or U2840 (N_2840,In_678,In_694);
or U2841 (N_2841,In_395,In_249);
or U2842 (N_2842,In_752,In_797);
and U2843 (N_2843,In_347,In_353);
or U2844 (N_2844,In_499,In_9);
and U2845 (N_2845,In_15,In_563);
nor U2846 (N_2846,In_577,In_290);
and U2847 (N_2847,In_691,In_408);
nand U2848 (N_2848,In_767,In_992);
xor U2849 (N_2849,In_385,In_266);
nor U2850 (N_2850,In_797,In_845);
or U2851 (N_2851,In_419,In_737);
nand U2852 (N_2852,In_971,In_49);
xor U2853 (N_2853,In_494,In_205);
or U2854 (N_2854,In_304,In_351);
and U2855 (N_2855,In_417,In_475);
xnor U2856 (N_2856,In_49,In_822);
or U2857 (N_2857,In_727,In_320);
and U2858 (N_2858,In_25,In_899);
xor U2859 (N_2859,In_942,In_8);
nand U2860 (N_2860,In_500,In_451);
xor U2861 (N_2861,In_409,In_345);
or U2862 (N_2862,In_661,In_516);
and U2863 (N_2863,In_772,In_252);
nand U2864 (N_2864,In_684,In_451);
nand U2865 (N_2865,In_542,In_508);
xor U2866 (N_2866,In_277,In_980);
or U2867 (N_2867,In_553,In_659);
nand U2868 (N_2868,In_525,In_30);
and U2869 (N_2869,In_81,In_755);
or U2870 (N_2870,In_626,In_790);
nand U2871 (N_2871,In_830,In_914);
xnor U2872 (N_2872,In_509,In_12);
nor U2873 (N_2873,In_239,In_242);
xnor U2874 (N_2874,In_714,In_784);
or U2875 (N_2875,In_284,In_400);
xor U2876 (N_2876,In_728,In_932);
or U2877 (N_2877,In_898,In_421);
nor U2878 (N_2878,In_482,In_600);
nor U2879 (N_2879,In_599,In_940);
nor U2880 (N_2880,In_934,In_554);
xor U2881 (N_2881,In_320,In_906);
and U2882 (N_2882,In_769,In_25);
or U2883 (N_2883,In_809,In_821);
nand U2884 (N_2884,In_940,In_623);
and U2885 (N_2885,In_507,In_634);
or U2886 (N_2886,In_333,In_218);
xnor U2887 (N_2887,In_577,In_72);
nand U2888 (N_2888,In_82,In_903);
nor U2889 (N_2889,In_421,In_717);
and U2890 (N_2890,In_22,In_24);
and U2891 (N_2891,In_769,In_680);
xnor U2892 (N_2892,In_914,In_351);
xor U2893 (N_2893,In_644,In_947);
xor U2894 (N_2894,In_211,In_671);
nor U2895 (N_2895,In_723,In_411);
nand U2896 (N_2896,In_166,In_503);
nand U2897 (N_2897,In_960,In_70);
xnor U2898 (N_2898,In_189,In_376);
or U2899 (N_2899,In_390,In_994);
nor U2900 (N_2900,In_24,In_692);
nand U2901 (N_2901,In_502,In_271);
or U2902 (N_2902,In_48,In_495);
xor U2903 (N_2903,In_96,In_330);
xor U2904 (N_2904,In_124,In_313);
xnor U2905 (N_2905,In_450,In_909);
nor U2906 (N_2906,In_731,In_5);
xor U2907 (N_2907,In_206,In_291);
nand U2908 (N_2908,In_787,In_718);
xor U2909 (N_2909,In_508,In_675);
or U2910 (N_2910,In_155,In_288);
xnor U2911 (N_2911,In_703,In_809);
nor U2912 (N_2912,In_354,In_452);
xnor U2913 (N_2913,In_318,In_433);
nor U2914 (N_2914,In_950,In_673);
nor U2915 (N_2915,In_428,In_378);
xor U2916 (N_2916,In_232,In_310);
and U2917 (N_2917,In_349,In_288);
nand U2918 (N_2918,In_852,In_741);
xnor U2919 (N_2919,In_57,In_938);
nand U2920 (N_2920,In_381,In_632);
and U2921 (N_2921,In_685,In_816);
nand U2922 (N_2922,In_278,In_530);
and U2923 (N_2923,In_640,In_326);
nor U2924 (N_2924,In_127,In_552);
nand U2925 (N_2925,In_142,In_263);
nor U2926 (N_2926,In_231,In_46);
nand U2927 (N_2927,In_533,In_975);
or U2928 (N_2928,In_221,In_8);
or U2929 (N_2929,In_720,In_685);
nand U2930 (N_2930,In_296,In_964);
or U2931 (N_2931,In_737,In_266);
xor U2932 (N_2932,In_28,In_301);
nor U2933 (N_2933,In_18,In_586);
xnor U2934 (N_2934,In_551,In_206);
nor U2935 (N_2935,In_302,In_388);
nand U2936 (N_2936,In_572,In_443);
and U2937 (N_2937,In_767,In_42);
xnor U2938 (N_2938,In_283,In_1);
nor U2939 (N_2939,In_627,In_893);
nand U2940 (N_2940,In_972,In_222);
nand U2941 (N_2941,In_365,In_945);
and U2942 (N_2942,In_521,In_20);
or U2943 (N_2943,In_432,In_508);
xor U2944 (N_2944,In_252,In_188);
and U2945 (N_2945,In_84,In_156);
or U2946 (N_2946,In_316,In_314);
nand U2947 (N_2947,In_395,In_733);
or U2948 (N_2948,In_401,In_136);
nand U2949 (N_2949,In_648,In_533);
xor U2950 (N_2950,In_60,In_665);
nor U2951 (N_2951,In_588,In_251);
nor U2952 (N_2952,In_797,In_683);
nor U2953 (N_2953,In_521,In_958);
nand U2954 (N_2954,In_628,In_151);
xnor U2955 (N_2955,In_897,In_514);
or U2956 (N_2956,In_281,In_267);
or U2957 (N_2957,In_951,In_362);
and U2958 (N_2958,In_145,In_222);
xnor U2959 (N_2959,In_406,In_630);
and U2960 (N_2960,In_312,In_487);
nand U2961 (N_2961,In_107,In_868);
nand U2962 (N_2962,In_481,In_1);
and U2963 (N_2963,In_444,In_546);
and U2964 (N_2964,In_955,In_35);
nand U2965 (N_2965,In_993,In_78);
nand U2966 (N_2966,In_10,In_157);
or U2967 (N_2967,In_761,In_393);
nor U2968 (N_2968,In_63,In_585);
xor U2969 (N_2969,In_635,In_215);
and U2970 (N_2970,In_819,In_755);
or U2971 (N_2971,In_312,In_51);
nand U2972 (N_2972,In_368,In_372);
nand U2973 (N_2973,In_312,In_455);
nand U2974 (N_2974,In_667,In_675);
xnor U2975 (N_2975,In_578,In_337);
xnor U2976 (N_2976,In_534,In_921);
or U2977 (N_2977,In_608,In_45);
and U2978 (N_2978,In_897,In_497);
or U2979 (N_2979,In_273,In_755);
xor U2980 (N_2980,In_759,In_924);
and U2981 (N_2981,In_830,In_610);
xor U2982 (N_2982,In_421,In_854);
or U2983 (N_2983,In_756,In_323);
nor U2984 (N_2984,In_821,In_672);
or U2985 (N_2985,In_625,In_674);
xnor U2986 (N_2986,In_355,In_60);
and U2987 (N_2987,In_614,In_786);
nor U2988 (N_2988,In_10,In_863);
and U2989 (N_2989,In_535,In_533);
or U2990 (N_2990,In_808,In_611);
and U2991 (N_2991,In_710,In_662);
nor U2992 (N_2992,In_990,In_627);
nor U2993 (N_2993,In_490,In_316);
nand U2994 (N_2994,In_790,In_787);
nor U2995 (N_2995,In_884,In_681);
or U2996 (N_2996,In_867,In_686);
and U2997 (N_2997,In_624,In_691);
or U2998 (N_2998,In_842,In_319);
nor U2999 (N_2999,In_128,In_948);
and U3000 (N_3000,In_53,In_641);
and U3001 (N_3001,In_480,In_322);
xnor U3002 (N_3002,In_873,In_972);
or U3003 (N_3003,In_6,In_166);
or U3004 (N_3004,In_27,In_712);
nor U3005 (N_3005,In_220,In_937);
xor U3006 (N_3006,In_991,In_569);
and U3007 (N_3007,In_384,In_66);
xor U3008 (N_3008,In_134,In_906);
xor U3009 (N_3009,In_776,In_738);
nand U3010 (N_3010,In_298,In_150);
nor U3011 (N_3011,In_899,In_340);
or U3012 (N_3012,In_71,In_420);
nor U3013 (N_3013,In_473,In_152);
and U3014 (N_3014,In_282,In_445);
xor U3015 (N_3015,In_816,In_80);
and U3016 (N_3016,In_756,In_636);
and U3017 (N_3017,In_191,In_391);
nor U3018 (N_3018,In_903,In_386);
or U3019 (N_3019,In_412,In_73);
or U3020 (N_3020,In_561,In_842);
or U3021 (N_3021,In_713,In_64);
xnor U3022 (N_3022,In_707,In_236);
nor U3023 (N_3023,In_919,In_60);
or U3024 (N_3024,In_270,In_163);
nor U3025 (N_3025,In_611,In_144);
or U3026 (N_3026,In_841,In_689);
and U3027 (N_3027,In_247,In_429);
and U3028 (N_3028,In_48,In_829);
or U3029 (N_3029,In_136,In_919);
nor U3030 (N_3030,In_739,In_274);
nor U3031 (N_3031,In_796,In_869);
or U3032 (N_3032,In_890,In_810);
and U3033 (N_3033,In_783,In_385);
and U3034 (N_3034,In_492,In_307);
xnor U3035 (N_3035,In_982,In_530);
xnor U3036 (N_3036,In_984,In_644);
nor U3037 (N_3037,In_203,In_880);
xnor U3038 (N_3038,In_857,In_289);
and U3039 (N_3039,In_515,In_805);
xor U3040 (N_3040,In_287,In_129);
or U3041 (N_3041,In_437,In_563);
xnor U3042 (N_3042,In_555,In_349);
and U3043 (N_3043,In_452,In_303);
and U3044 (N_3044,In_588,In_51);
nor U3045 (N_3045,In_884,In_91);
and U3046 (N_3046,In_902,In_649);
and U3047 (N_3047,In_256,In_25);
xor U3048 (N_3048,In_255,In_454);
xnor U3049 (N_3049,In_164,In_932);
or U3050 (N_3050,In_624,In_302);
and U3051 (N_3051,In_425,In_960);
nand U3052 (N_3052,In_984,In_358);
nand U3053 (N_3053,In_613,In_2);
and U3054 (N_3054,In_957,In_279);
xor U3055 (N_3055,In_938,In_517);
and U3056 (N_3056,In_623,In_848);
xor U3057 (N_3057,In_543,In_236);
or U3058 (N_3058,In_468,In_184);
xor U3059 (N_3059,In_649,In_361);
nor U3060 (N_3060,In_953,In_372);
and U3061 (N_3061,In_363,In_349);
or U3062 (N_3062,In_282,In_551);
nand U3063 (N_3063,In_233,In_842);
nor U3064 (N_3064,In_206,In_593);
nor U3065 (N_3065,In_430,In_903);
or U3066 (N_3066,In_773,In_769);
or U3067 (N_3067,In_55,In_321);
nor U3068 (N_3068,In_900,In_518);
or U3069 (N_3069,In_543,In_747);
nor U3070 (N_3070,In_657,In_821);
or U3071 (N_3071,In_17,In_664);
xor U3072 (N_3072,In_192,In_262);
and U3073 (N_3073,In_622,In_74);
or U3074 (N_3074,In_484,In_117);
and U3075 (N_3075,In_973,In_713);
or U3076 (N_3076,In_290,In_129);
nand U3077 (N_3077,In_758,In_780);
nor U3078 (N_3078,In_909,In_783);
and U3079 (N_3079,In_0,In_968);
nor U3080 (N_3080,In_593,In_545);
and U3081 (N_3081,In_994,In_613);
nand U3082 (N_3082,In_72,In_400);
or U3083 (N_3083,In_104,In_267);
nor U3084 (N_3084,In_587,In_299);
and U3085 (N_3085,In_754,In_961);
xor U3086 (N_3086,In_803,In_696);
xnor U3087 (N_3087,In_978,In_681);
nand U3088 (N_3088,In_87,In_744);
and U3089 (N_3089,In_674,In_378);
xnor U3090 (N_3090,In_38,In_973);
nand U3091 (N_3091,In_784,In_700);
and U3092 (N_3092,In_555,In_133);
nand U3093 (N_3093,In_242,In_60);
nor U3094 (N_3094,In_555,In_366);
xnor U3095 (N_3095,In_422,In_567);
and U3096 (N_3096,In_783,In_696);
nor U3097 (N_3097,In_555,In_999);
and U3098 (N_3098,In_513,In_903);
xnor U3099 (N_3099,In_703,In_380);
xor U3100 (N_3100,In_211,In_175);
and U3101 (N_3101,In_51,In_171);
nor U3102 (N_3102,In_778,In_375);
or U3103 (N_3103,In_544,In_706);
nand U3104 (N_3104,In_214,In_783);
nand U3105 (N_3105,In_376,In_257);
xor U3106 (N_3106,In_778,In_409);
xor U3107 (N_3107,In_97,In_259);
and U3108 (N_3108,In_814,In_614);
and U3109 (N_3109,In_41,In_197);
xor U3110 (N_3110,In_189,In_300);
and U3111 (N_3111,In_571,In_216);
xor U3112 (N_3112,In_559,In_638);
xnor U3113 (N_3113,In_378,In_598);
nand U3114 (N_3114,In_871,In_861);
nand U3115 (N_3115,In_789,In_37);
xnor U3116 (N_3116,In_731,In_185);
and U3117 (N_3117,In_897,In_849);
nand U3118 (N_3118,In_419,In_673);
xnor U3119 (N_3119,In_211,In_802);
nor U3120 (N_3120,In_372,In_34);
nor U3121 (N_3121,In_749,In_593);
and U3122 (N_3122,In_158,In_705);
and U3123 (N_3123,In_191,In_315);
nor U3124 (N_3124,In_35,In_367);
xnor U3125 (N_3125,In_392,In_303);
nor U3126 (N_3126,In_447,In_886);
or U3127 (N_3127,In_460,In_762);
nand U3128 (N_3128,In_14,In_469);
nor U3129 (N_3129,In_696,In_553);
nor U3130 (N_3130,In_23,In_84);
and U3131 (N_3131,In_788,In_538);
xnor U3132 (N_3132,In_115,In_642);
or U3133 (N_3133,In_102,In_333);
nand U3134 (N_3134,In_374,In_110);
nand U3135 (N_3135,In_415,In_97);
or U3136 (N_3136,In_486,In_144);
or U3137 (N_3137,In_213,In_344);
and U3138 (N_3138,In_801,In_752);
and U3139 (N_3139,In_433,In_755);
xnor U3140 (N_3140,In_915,In_41);
nor U3141 (N_3141,In_710,In_213);
and U3142 (N_3142,In_514,In_721);
xnor U3143 (N_3143,In_7,In_679);
and U3144 (N_3144,In_603,In_615);
xor U3145 (N_3145,In_640,In_228);
or U3146 (N_3146,In_107,In_166);
xor U3147 (N_3147,In_677,In_158);
xnor U3148 (N_3148,In_438,In_639);
xor U3149 (N_3149,In_183,In_168);
xnor U3150 (N_3150,In_815,In_791);
nand U3151 (N_3151,In_790,In_585);
and U3152 (N_3152,In_958,In_33);
nor U3153 (N_3153,In_379,In_997);
nor U3154 (N_3154,In_403,In_476);
xnor U3155 (N_3155,In_191,In_637);
nand U3156 (N_3156,In_881,In_361);
xnor U3157 (N_3157,In_71,In_121);
xnor U3158 (N_3158,In_521,In_833);
or U3159 (N_3159,In_336,In_981);
nor U3160 (N_3160,In_385,In_2);
xor U3161 (N_3161,In_415,In_126);
nand U3162 (N_3162,In_114,In_841);
and U3163 (N_3163,In_837,In_252);
and U3164 (N_3164,In_330,In_120);
or U3165 (N_3165,In_8,In_872);
nor U3166 (N_3166,In_987,In_516);
or U3167 (N_3167,In_11,In_146);
xnor U3168 (N_3168,In_222,In_624);
nand U3169 (N_3169,In_660,In_967);
or U3170 (N_3170,In_373,In_861);
and U3171 (N_3171,In_94,In_646);
xor U3172 (N_3172,In_190,In_898);
xnor U3173 (N_3173,In_118,In_980);
xor U3174 (N_3174,In_17,In_36);
or U3175 (N_3175,In_894,In_913);
or U3176 (N_3176,In_116,In_434);
or U3177 (N_3177,In_707,In_853);
and U3178 (N_3178,In_144,In_279);
and U3179 (N_3179,In_792,In_603);
and U3180 (N_3180,In_299,In_132);
nor U3181 (N_3181,In_752,In_16);
and U3182 (N_3182,In_977,In_765);
nand U3183 (N_3183,In_129,In_499);
nand U3184 (N_3184,In_35,In_345);
xor U3185 (N_3185,In_308,In_507);
and U3186 (N_3186,In_568,In_171);
nor U3187 (N_3187,In_877,In_169);
and U3188 (N_3188,In_665,In_950);
or U3189 (N_3189,In_535,In_617);
and U3190 (N_3190,In_504,In_403);
nand U3191 (N_3191,In_14,In_973);
and U3192 (N_3192,In_322,In_931);
nor U3193 (N_3193,In_592,In_536);
and U3194 (N_3194,In_630,In_468);
nor U3195 (N_3195,In_165,In_901);
nand U3196 (N_3196,In_900,In_534);
nor U3197 (N_3197,In_210,In_116);
nor U3198 (N_3198,In_615,In_88);
nor U3199 (N_3199,In_38,In_61);
nor U3200 (N_3200,In_870,In_715);
nand U3201 (N_3201,In_362,In_949);
and U3202 (N_3202,In_585,In_275);
or U3203 (N_3203,In_976,In_12);
nor U3204 (N_3204,In_969,In_218);
nor U3205 (N_3205,In_401,In_474);
nor U3206 (N_3206,In_107,In_795);
xnor U3207 (N_3207,In_800,In_831);
xor U3208 (N_3208,In_665,In_711);
xor U3209 (N_3209,In_871,In_570);
and U3210 (N_3210,In_224,In_39);
nand U3211 (N_3211,In_255,In_205);
and U3212 (N_3212,In_101,In_137);
or U3213 (N_3213,In_448,In_203);
xor U3214 (N_3214,In_876,In_165);
nor U3215 (N_3215,In_168,In_90);
nand U3216 (N_3216,In_560,In_82);
or U3217 (N_3217,In_635,In_429);
and U3218 (N_3218,In_377,In_134);
or U3219 (N_3219,In_453,In_196);
nand U3220 (N_3220,In_99,In_472);
nand U3221 (N_3221,In_313,In_286);
xnor U3222 (N_3222,In_834,In_799);
or U3223 (N_3223,In_124,In_782);
nand U3224 (N_3224,In_708,In_543);
nand U3225 (N_3225,In_483,In_950);
and U3226 (N_3226,In_31,In_518);
xnor U3227 (N_3227,In_855,In_381);
xnor U3228 (N_3228,In_906,In_666);
xnor U3229 (N_3229,In_593,In_22);
nor U3230 (N_3230,In_838,In_100);
or U3231 (N_3231,In_250,In_691);
and U3232 (N_3232,In_938,In_65);
nand U3233 (N_3233,In_831,In_858);
nor U3234 (N_3234,In_411,In_739);
or U3235 (N_3235,In_427,In_264);
nand U3236 (N_3236,In_889,In_352);
or U3237 (N_3237,In_598,In_129);
and U3238 (N_3238,In_934,In_116);
and U3239 (N_3239,In_13,In_102);
nand U3240 (N_3240,In_952,In_344);
xnor U3241 (N_3241,In_974,In_445);
or U3242 (N_3242,In_569,In_450);
nor U3243 (N_3243,In_685,In_409);
nand U3244 (N_3244,In_470,In_810);
xor U3245 (N_3245,In_729,In_84);
xnor U3246 (N_3246,In_140,In_757);
xnor U3247 (N_3247,In_32,In_863);
and U3248 (N_3248,In_213,In_60);
and U3249 (N_3249,In_548,In_404);
and U3250 (N_3250,In_380,In_810);
nand U3251 (N_3251,In_329,In_540);
and U3252 (N_3252,In_776,In_306);
nand U3253 (N_3253,In_669,In_160);
or U3254 (N_3254,In_115,In_444);
nor U3255 (N_3255,In_872,In_41);
or U3256 (N_3256,In_6,In_605);
or U3257 (N_3257,In_169,In_431);
nand U3258 (N_3258,In_532,In_105);
or U3259 (N_3259,In_898,In_884);
nor U3260 (N_3260,In_721,In_808);
nand U3261 (N_3261,In_846,In_556);
nor U3262 (N_3262,In_552,In_984);
and U3263 (N_3263,In_744,In_693);
nand U3264 (N_3264,In_58,In_470);
nand U3265 (N_3265,In_791,In_771);
nand U3266 (N_3266,In_852,In_615);
xor U3267 (N_3267,In_279,In_314);
nor U3268 (N_3268,In_759,In_85);
or U3269 (N_3269,In_420,In_688);
xnor U3270 (N_3270,In_697,In_206);
or U3271 (N_3271,In_347,In_76);
or U3272 (N_3272,In_533,In_760);
or U3273 (N_3273,In_860,In_315);
nand U3274 (N_3274,In_866,In_78);
nand U3275 (N_3275,In_410,In_793);
nand U3276 (N_3276,In_351,In_782);
nand U3277 (N_3277,In_534,In_204);
or U3278 (N_3278,In_658,In_352);
xnor U3279 (N_3279,In_607,In_710);
nor U3280 (N_3280,In_431,In_72);
nand U3281 (N_3281,In_463,In_337);
nand U3282 (N_3282,In_448,In_113);
nor U3283 (N_3283,In_966,In_849);
xor U3284 (N_3284,In_433,In_228);
nand U3285 (N_3285,In_944,In_286);
or U3286 (N_3286,In_439,In_589);
xor U3287 (N_3287,In_38,In_135);
nand U3288 (N_3288,In_91,In_194);
nor U3289 (N_3289,In_380,In_460);
nor U3290 (N_3290,In_754,In_107);
nor U3291 (N_3291,In_242,In_693);
and U3292 (N_3292,In_809,In_302);
and U3293 (N_3293,In_491,In_277);
nor U3294 (N_3294,In_705,In_684);
or U3295 (N_3295,In_917,In_837);
nor U3296 (N_3296,In_563,In_833);
nand U3297 (N_3297,In_970,In_53);
and U3298 (N_3298,In_738,In_371);
xor U3299 (N_3299,In_926,In_29);
xor U3300 (N_3300,In_432,In_991);
or U3301 (N_3301,In_912,In_435);
and U3302 (N_3302,In_946,In_73);
and U3303 (N_3303,In_972,In_687);
or U3304 (N_3304,In_118,In_640);
or U3305 (N_3305,In_276,In_592);
and U3306 (N_3306,In_965,In_575);
and U3307 (N_3307,In_940,In_174);
and U3308 (N_3308,In_421,In_73);
or U3309 (N_3309,In_189,In_845);
and U3310 (N_3310,In_313,In_326);
nor U3311 (N_3311,In_852,In_625);
or U3312 (N_3312,In_391,In_403);
or U3313 (N_3313,In_957,In_450);
and U3314 (N_3314,In_238,In_45);
nand U3315 (N_3315,In_397,In_57);
or U3316 (N_3316,In_574,In_834);
xnor U3317 (N_3317,In_714,In_566);
and U3318 (N_3318,In_545,In_665);
and U3319 (N_3319,In_808,In_960);
xnor U3320 (N_3320,In_339,In_940);
or U3321 (N_3321,In_910,In_750);
xor U3322 (N_3322,In_294,In_663);
nand U3323 (N_3323,In_505,In_845);
xor U3324 (N_3324,In_192,In_964);
nand U3325 (N_3325,In_408,In_253);
nand U3326 (N_3326,In_54,In_758);
xnor U3327 (N_3327,In_104,In_509);
and U3328 (N_3328,In_716,In_767);
or U3329 (N_3329,In_120,In_708);
and U3330 (N_3330,In_465,In_821);
and U3331 (N_3331,In_89,In_268);
and U3332 (N_3332,In_954,In_131);
and U3333 (N_3333,In_364,In_368);
nand U3334 (N_3334,In_574,In_228);
xor U3335 (N_3335,In_198,In_563);
nand U3336 (N_3336,In_592,In_100);
or U3337 (N_3337,In_338,In_304);
xnor U3338 (N_3338,In_784,In_465);
nor U3339 (N_3339,In_395,In_355);
and U3340 (N_3340,In_301,In_979);
xnor U3341 (N_3341,In_912,In_465);
xor U3342 (N_3342,In_240,In_428);
or U3343 (N_3343,In_265,In_221);
and U3344 (N_3344,In_73,In_126);
and U3345 (N_3345,In_561,In_789);
or U3346 (N_3346,In_596,In_90);
nor U3347 (N_3347,In_497,In_616);
and U3348 (N_3348,In_172,In_626);
nor U3349 (N_3349,In_801,In_197);
nand U3350 (N_3350,In_618,In_536);
and U3351 (N_3351,In_51,In_260);
nor U3352 (N_3352,In_181,In_260);
nor U3353 (N_3353,In_845,In_182);
nor U3354 (N_3354,In_774,In_754);
and U3355 (N_3355,In_265,In_301);
or U3356 (N_3356,In_848,In_911);
or U3357 (N_3357,In_452,In_306);
and U3358 (N_3358,In_615,In_988);
and U3359 (N_3359,In_795,In_348);
nand U3360 (N_3360,In_46,In_724);
or U3361 (N_3361,In_311,In_807);
nor U3362 (N_3362,In_429,In_18);
and U3363 (N_3363,In_870,In_605);
nor U3364 (N_3364,In_295,In_683);
xnor U3365 (N_3365,In_948,In_366);
nor U3366 (N_3366,In_644,In_940);
or U3367 (N_3367,In_339,In_207);
nand U3368 (N_3368,In_783,In_88);
nor U3369 (N_3369,In_897,In_901);
or U3370 (N_3370,In_972,In_481);
xor U3371 (N_3371,In_173,In_250);
nand U3372 (N_3372,In_839,In_132);
and U3373 (N_3373,In_891,In_10);
or U3374 (N_3374,In_875,In_988);
or U3375 (N_3375,In_61,In_107);
or U3376 (N_3376,In_949,In_909);
or U3377 (N_3377,In_586,In_190);
xor U3378 (N_3378,In_462,In_933);
nor U3379 (N_3379,In_308,In_754);
and U3380 (N_3380,In_988,In_730);
xnor U3381 (N_3381,In_853,In_932);
nand U3382 (N_3382,In_346,In_436);
and U3383 (N_3383,In_632,In_61);
nor U3384 (N_3384,In_141,In_466);
nor U3385 (N_3385,In_250,In_657);
nand U3386 (N_3386,In_158,In_706);
and U3387 (N_3387,In_209,In_607);
and U3388 (N_3388,In_352,In_473);
nand U3389 (N_3389,In_394,In_881);
and U3390 (N_3390,In_361,In_9);
or U3391 (N_3391,In_965,In_223);
nor U3392 (N_3392,In_634,In_433);
and U3393 (N_3393,In_601,In_833);
xnor U3394 (N_3394,In_412,In_840);
or U3395 (N_3395,In_663,In_27);
or U3396 (N_3396,In_888,In_348);
nor U3397 (N_3397,In_436,In_220);
xnor U3398 (N_3398,In_827,In_417);
or U3399 (N_3399,In_793,In_960);
nor U3400 (N_3400,In_885,In_259);
or U3401 (N_3401,In_388,In_379);
and U3402 (N_3402,In_670,In_609);
xnor U3403 (N_3403,In_970,In_633);
nor U3404 (N_3404,In_506,In_432);
nor U3405 (N_3405,In_195,In_116);
and U3406 (N_3406,In_505,In_604);
xor U3407 (N_3407,In_371,In_655);
and U3408 (N_3408,In_412,In_750);
and U3409 (N_3409,In_204,In_655);
nand U3410 (N_3410,In_359,In_680);
and U3411 (N_3411,In_434,In_30);
or U3412 (N_3412,In_951,In_227);
nand U3413 (N_3413,In_47,In_747);
and U3414 (N_3414,In_95,In_856);
nor U3415 (N_3415,In_297,In_554);
and U3416 (N_3416,In_282,In_161);
and U3417 (N_3417,In_627,In_220);
nor U3418 (N_3418,In_255,In_402);
and U3419 (N_3419,In_972,In_211);
xnor U3420 (N_3420,In_990,In_303);
and U3421 (N_3421,In_823,In_397);
or U3422 (N_3422,In_242,In_840);
xnor U3423 (N_3423,In_362,In_940);
nor U3424 (N_3424,In_473,In_423);
xnor U3425 (N_3425,In_399,In_224);
nand U3426 (N_3426,In_325,In_159);
nand U3427 (N_3427,In_168,In_574);
nand U3428 (N_3428,In_895,In_714);
xor U3429 (N_3429,In_886,In_627);
nor U3430 (N_3430,In_303,In_568);
nor U3431 (N_3431,In_90,In_984);
nand U3432 (N_3432,In_828,In_856);
or U3433 (N_3433,In_768,In_243);
nor U3434 (N_3434,In_68,In_169);
and U3435 (N_3435,In_119,In_24);
and U3436 (N_3436,In_338,In_781);
and U3437 (N_3437,In_45,In_449);
nor U3438 (N_3438,In_519,In_956);
nor U3439 (N_3439,In_729,In_50);
nand U3440 (N_3440,In_884,In_789);
and U3441 (N_3441,In_773,In_355);
or U3442 (N_3442,In_139,In_361);
nor U3443 (N_3443,In_225,In_584);
xnor U3444 (N_3444,In_212,In_300);
nor U3445 (N_3445,In_603,In_358);
nand U3446 (N_3446,In_402,In_840);
or U3447 (N_3447,In_484,In_624);
nor U3448 (N_3448,In_774,In_166);
or U3449 (N_3449,In_184,In_898);
and U3450 (N_3450,In_599,In_42);
nand U3451 (N_3451,In_799,In_649);
xor U3452 (N_3452,In_828,In_970);
nor U3453 (N_3453,In_745,In_288);
xor U3454 (N_3454,In_44,In_579);
and U3455 (N_3455,In_587,In_256);
nand U3456 (N_3456,In_915,In_282);
nand U3457 (N_3457,In_984,In_894);
or U3458 (N_3458,In_370,In_28);
or U3459 (N_3459,In_133,In_867);
xor U3460 (N_3460,In_790,In_960);
and U3461 (N_3461,In_494,In_585);
xnor U3462 (N_3462,In_825,In_495);
nand U3463 (N_3463,In_917,In_940);
nor U3464 (N_3464,In_685,In_630);
xnor U3465 (N_3465,In_620,In_532);
nor U3466 (N_3466,In_498,In_457);
xor U3467 (N_3467,In_173,In_278);
or U3468 (N_3468,In_922,In_822);
nand U3469 (N_3469,In_344,In_797);
and U3470 (N_3470,In_151,In_300);
xor U3471 (N_3471,In_780,In_597);
xor U3472 (N_3472,In_416,In_871);
and U3473 (N_3473,In_221,In_791);
xor U3474 (N_3474,In_312,In_828);
or U3475 (N_3475,In_227,In_168);
nand U3476 (N_3476,In_661,In_199);
or U3477 (N_3477,In_976,In_399);
and U3478 (N_3478,In_710,In_207);
and U3479 (N_3479,In_596,In_860);
xor U3480 (N_3480,In_109,In_376);
xnor U3481 (N_3481,In_493,In_969);
xor U3482 (N_3482,In_230,In_104);
nor U3483 (N_3483,In_598,In_13);
nor U3484 (N_3484,In_523,In_849);
xor U3485 (N_3485,In_438,In_487);
or U3486 (N_3486,In_136,In_229);
nand U3487 (N_3487,In_247,In_698);
or U3488 (N_3488,In_262,In_574);
and U3489 (N_3489,In_637,In_599);
xor U3490 (N_3490,In_22,In_927);
xnor U3491 (N_3491,In_700,In_456);
xor U3492 (N_3492,In_639,In_2);
nor U3493 (N_3493,In_441,In_25);
xnor U3494 (N_3494,In_368,In_313);
xnor U3495 (N_3495,In_32,In_89);
nand U3496 (N_3496,In_797,In_774);
or U3497 (N_3497,In_137,In_103);
and U3498 (N_3498,In_970,In_785);
and U3499 (N_3499,In_320,In_795);
nor U3500 (N_3500,In_388,In_34);
and U3501 (N_3501,In_725,In_765);
or U3502 (N_3502,In_236,In_923);
or U3503 (N_3503,In_943,In_686);
xnor U3504 (N_3504,In_926,In_606);
and U3505 (N_3505,In_348,In_643);
nand U3506 (N_3506,In_892,In_311);
nand U3507 (N_3507,In_758,In_183);
xor U3508 (N_3508,In_705,In_26);
nand U3509 (N_3509,In_560,In_793);
or U3510 (N_3510,In_116,In_159);
nand U3511 (N_3511,In_849,In_328);
or U3512 (N_3512,In_238,In_308);
and U3513 (N_3513,In_695,In_790);
nor U3514 (N_3514,In_690,In_930);
nand U3515 (N_3515,In_791,In_558);
or U3516 (N_3516,In_138,In_685);
xor U3517 (N_3517,In_643,In_983);
and U3518 (N_3518,In_658,In_791);
xnor U3519 (N_3519,In_422,In_626);
and U3520 (N_3520,In_880,In_830);
nor U3521 (N_3521,In_558,In_665);
xnor U3522 (N_3522,In_441,In_909);
and U3523 (N_3523,In_72,In_987);
xor U3524 (N_3524,In_518,In_285);
nor U3525 (N_3525,In_48,In_196);
nand U3526 (N_3526,In_344,In_340);
nor U3527 (N_3527,In_699,In_775);
nand U3528 (N_3528,In_490,In_13);
nand U3529 (N_3529,In_466,In_833);
xnor U3530 (N_3530,In_755,In_930);
xnor U3531 (N_3531,In_668,In_868);
and U3532 (N_3532,In_778,In_452);
nand U3533 (N_3533,In_872,In_931);
nor U3534 (N_3534,In_952,In_208);
nand U3535 (N_3535,In_642,In_667);
nor U3536 (N_3536,In_569,In_275);
or U3537 (N_3537,In_642,In_962);
nor U3538 (N_3538,In_523,In_692);
or U3539 (N_3539,In_348,In_44);
or U3540 (N_3540,In_848,In_0);
nor U3541 (N_3541,In_153,In_422);
and U3542 (N_3542,In_177,In_296);
nand U3543 (N_3543,In_484,In_777);
and U3544 (N_3544,In_997,In_932);
nor U3545 (N_3545,In_199,In_918);
and U3546 (N_3546,In_290,In_469);
or U3547 (N_3547,In_860,In_816);
and U3548 (N_3548,In_660,In_127);
xnor U3549 (N_3549,In_594,In_26);
and U3550 (N_3550,In_162,In_758);
or U3551 (N_3551,In_414,In_933);
or U3552 (N_3552,In_847,In_971);
nand U3553 (N_3553,In_852,In_282);
and U3554 (N_3554,In_897,In_952);
xor U3555 (N_3555,In_627,In_515);
nand U3556 (N_3556,In_401,In_85);
and U3557 (N_3557,In_803,In_219);
and U3558 (N_3558,In_415,In_306);
or U3559 (N_3559,In_831,In_718);
nor U3560 (N_3560,In_995,In_782);
xnor U3561 (N_3561,In_693,In_945);
and U3562 (N_3562,In_123,In_963);
nor U3563 (N_3563,In_676,In_73);
and U3564 (N_3564,In_985,In_698);
and U3565 (N_3565,In_218,In_314);
or U3566 (N_3566,In_650,In_952);
or U3567 (N_3567,In_677,In_656);
nand U3568 (N_3568,In_356,In_858);
or U3569 (N_3569,In_810,In_411);
nor U3570 (N_3570,In_34,In_50);
nor U3571 (N_3571,In_415,In_175);
or U3572 (N_3572,In_528,In_178);
nor U3573 (N_3573,In_296,In_273);
nor U3574 (N_3574,In_39,In_190);
nor U3575 (N_3575,In_0,In_985);
and U3576 (N_3576,In_875,In_406);
xnor U3577 (N_3577,In_567,In_160);
nand U3578 (N_3578,In_330,In_414);
xnor U3579 (N_3579,In_891,In_531);
and U3580 (N_3580,In_317,In_569);
and U3581 (N_3581,In_134,In_945);
or U3582 (N_3582,In_672,In_96);
or U3583 (N_3583,In_875,In_989);
and U3584 (N_3584,In_526,In_705);
and U3585 (N_3585,In_829,In_937);
and U3586 (N_3586,In_243,In_196);
and U3587 (N_3587,In_113,In_965);
nand U3588 (N_3588,In_901,In_232);
nor U3589 (N_3589,In_35,In_392);
nor U3590 (N_3590,In_10,In_659);
or U3591 (N_3591,In_707,In_582);
xnor U3592 (N_3592,In_312,In_909);
nor U3593 (N_3593,In_168,In_190);
xor U3594 (N_3594,In_484,In_894);
nand U3595 (N_3595,In_30,In_237);
nand U3596 (N_3596,In_977,In_996);
or U3597 (N_3597,In_739,In_313);
xor U3598 (N_3598,In_856,In_623);
xor U3599 (N_3599,In_175,In_677);
nor U3600 (N_3600,In_659,In_411);
or U3601 (N_3601,In_420,In_391);
nor U3602 (N_3602,In_774,In_692);
or U3603 (N_3603,In_875,In_785);
nand U3604 (N_3604,In_240,In_919);
nand U3605 (N_3605,In_537,In_784);
or U3606 (N_3606,In_193,In_661);
xor U3607 (N_3607,In_887,In_408);
or U3608 (N_3608,In_34,In_209);
nor U3609 (N_3609,In_588,In_850);
nand U3610 (N_3610,In_6,In_904);
xor U3611 (N_3611,In_676,In_861);
and U3612 (N_3612,In_821,In_43);
and U3613 (N_3613,In_528,In_856);
nor U3614 (N_3614,In_499,In_691);
xor U3615 (N_3615,In_388,In_732);
xor U3616 (N_3616,In_400,In_679);
xnor U3617 (N_3617,In_939,In_558);
nor U3618 (N_3618,In_816,In_644);
nor U3619 (N_3619,In_9,In_419);
nand U3620 (N_3620,In_197,In_58);
nor U3621 (N_3621,In_938,In_2);
or U3622 (N_3622,In_786,In_548);
or U3623 (N_3623,In_522,In_594);
and U3624 (N_3624,In_415,In_472);
nand U3625 (N_3625,In_144,In_621);
nor U3626 (N_3626,In_234,In_344);
and U3627 (N_3627,In_804,In_631);
or U3628 (N_3628,In_633,In_480);
nor U3629 (N_3629,In_475,In_674);
nand U3630 (N_3630,In_991,In_973);
nand U3631 (N_3631,In_401,In_372);
nor U3632 (N_3632,In_441,In_656);
or U3633 (N_3633,In_246,In_523);
and U3634 (N_3634,In_591,In_918);
xnor U3635 (N_3635,In_910,In_939);
and U3636 (N_3636,In_422,In_841);
nand U3637 (N_3637,In_319,In_480);
or U3638 (N_3638,In_831,In_763);
and U3639 (N_3639,In_486,In_220);
nor U3640 (N_3640,In_486,In_707);
nand U3641 (N_3641,In_894,In_270);
and U3642 (N_3642,In_767,In_32);
or U3643 (N_3643,In_200,In_133);
nor U3644 (N_3644,In_365,In_598);
nand U3645 (N_3645,In_328,In_731);
and U3646 (N_3646,In_350,In_188);
nor U3647 (N_3647,In_488,In_23);
xnor U3648 (N_3648,In_571,In_450);
and U3649 (N_3649,In_967,In_710);
or U3650 (N_3650,In_545,In_358);
and U3651 (N_3651,In_329,In_188);
nand U3652 (N_3652,In_725,In_960);
xor U3653 (N_3653,In_462,In_265);
and U3654 (N_3654,In_78,In_426);
and U3655 (N_3655,In_923,In_565);
and U3656 (N_3656,In_829,In_59);
and U3657 (N_3657,In_3,In_567);
or U3658 (N_3658,In_411,In_287);
nand U3659 (N_3659,In_254,In_626);
nor U3660 (N_3660,In_448,In_458);
xor U3661 (N_3661,In_435,In_465);
nor U3662 (N_3662,In_980,In_435);
and U3663 (N_3663,In_398,In_949);
xor U3664 (N_3664,In_916,In_858);
nor U3665 (N_3665,In_581,In_44);
nor U3666 (N_3666,In_706,In_880);
and U3667 (N_3667,In_120,In_559);
or U3668 (N_3668,In_299,In_572);
or U3669 (N_3669,In_445,In_584);
xor U3670 (N_3670,In_426,In_869);
and U3671 (N_3671,In_987,In_254);
nand U3672 (N_3672,In_920,In_14);
or U3673 (N_3673,In_356,In_396);
nand U3674 (N_3674,In_843,In_174);
xnor U3675 (N_3675,In_687,In_70);
nand U3676 (N_3676,In_947,In_799);
nand U3677 (N_3677,In_197,In_378);
or U3678 (N_3678,In_977,In_952);
or U3679 (N_3679,In_837,In_803);
or U3680 (N_3680,In_50,In_405);
nor U3681 (N_3681,In_463,In_863);
xor U3682 (N_3682,In_739,In_806);
xor U3683 (N_3683,In_401,In_638);
nor U3684 (N_3684,In_465,In_896);
xor U3685 (N_3685,In_612,In_559);
nor U3686 (N_3686,In_399,In_747);
or U3687 (N_3687,In_780,In_242);
nand U3688 (N_3688,In_957,In_481);
and U3689 (N_3689,In_697,In_823);
xnor U3690 (N_3690,In_635,In_449);
nor U3691 (N_3691,In_209,In_479);
or U3692 (N_3692,In_832,In_983);
nand U3693 (N_3693,In_28,In_788);
and U3694 (N_3694,In_504,In_286);
or U3695 (N_3695,In_812,In_150);
nand U3696 (N_3696,In_992,In_35);
xor U3697 (N_3697,In_551,In_452);
nand U3698 (N_3698,In_698,In_424);
xor U3699 (N_3699,In_588,In_130);
and U3700 (N_3700,In_240,In_309);
or U3701 (N_3701,In_832,In_41);
nand U3702 (N_3702,In_874,In_748);
nand U3703 (N_3703,In_441,In_26);
nor U3704 (N_3704,In_947,In_950);
and U3705 (N_3705,In_605,In_710);
nor U3706 (N_3706,In_778,In_726);
nor U3707 (N_3707,In_828,In_494);
xnor U3708 (N_3708,In_156,In_901);
nor U3709 (N_3709,In_688,In_576);
nor U3710 (N_3710,In_625,In_190);
xor U3711 (N_3711,In_640,In_675);
or U3712 (N_3712,In_352,In_464);
nor U3713 (N_3713,In_538,In_946);
or U3714 (N_3714,In_714,In_635);
and U3715 (N_3715,In_654,In_488);
and U3716 (N_3716,In_917,In_470);
and U3717 (N_3717,In_641,In_697);
xor U3718 (N_3718,In_541,In_35);
or U3719 (N_3719,In_888,In_205);
xor U3720 (N_3720,In_870,In_432);
nor U3721 (N_3721,In_284,In_131);
nor U3722 (N_3722,In_203,In_513);
or U3723 (N_3723,In_752,In_359);
or U3724 (N_3724,In_430,In_442);
xnor U3725 (N_3725,In_327,In_852);
and U3726 (N_3726,In_451,In_980);
nand U3727 (N_3727,In_855,In_308);
and U3728 (N_3728,In_858,In_906);
and U3729 (N_3729,In_988,In_925);
nand U3730 (N_3730,In_553,In_394);
and U3731 (N_3731,In_125,In_270);
or U3732 (N_3732,In_209,In_347);
and U3733 (N_3733,In_976,In_890);
or U3734 (N_3734,In_270,In_715);
nor U3735 (N_3735,In_761,In_579);
or U3736 (N_3736,In_56,In_594);
and U3737 (N_3737,In_747,In_878);
xor U3738 (N_3738,In_395,In_975);
and U3739 (N_3739,In_60,In_426);
and U3740 (N_3740,In_346,In_413);
and U3741 (N_3741,In_699,In_421);
xnor U3742 (N_3742,In_584,In_931);
or U3743 (N_3743,In_584,In_789);
xnor U3744 (N_3744,In_829,In_517);
and U3745 (N_3745,In_890,In_931);
xnor U3746 (N_3746,In_940,In_481);
or U3747 (N_3747,In_852,In_514);
and U3748 (N_3748,In_530,In_955);
or U3749 (N_3749,In_203,In_566);
and U3750 (N_3750,In_912,In_328);
and U3751 (N_3751,In_557,In_492);
xor U3752 (N_3752,In_489,In_915);
and U3753 (N_3753,In_933,In_509);
or U3754 (N_3754,In_737,In_569);
nand U3755 (N_3755,In_174,In_37);
nor U3756 (N_3756,In_218,In_954);
xnor U3757 (N_3757,In_550,In_220);
nor U3758 (N_3758,In_614,In_855);
nand U3759 (N_3759,In_446,In_14);
and U3760 (N_3760,In_416,In_106);
nor U3761 (N_3761,In_92,In_698);
nor U3762 (N_3762,In_1,In_741);
nand U3763 (N_3763,In_733,In_506);
or U3764 (N_3764,In_443,In_19);
and U3765 (N_3765,In_174,In_108);
or U3766 (N_3766,In_120,In_631);
nor U3767 (N_3767,In_445,In_274);
xnor U3768 (N_3768,In_403,In_452);
nand U3769 (N_3769,In_785,In_625);
xnor U3770 (N_3770,In_233,In_429);
nor U3771 (N_3771,In_342,In_285);
or U3772 (N_3772,In_595,In_902);
xor U3773 (N_3773,In_698,In_925);
nand U3774 (N_3774,In_493,In_736);
xor U3775 (N_3775,In_480,In_411);
xnor U3776 (N_3776,In_332,In_364);
or U3777 (N_3777,In_606,In_23);
nor U3778 (N_3778,In_160,In_710);
nor U3779 (N_3779,In_389,In_71);
xor U3780 (N_3780,In_688,In_804);
xor U3781 (N_3781,In_695,In_177);
or U3782 (N_3782,In_728,In_436);
and U3783 (N_3783,In_247,In_473);
or U3784 (N_3784,In_663,In_928);
nor U3785 (N_3785,In_520,In_363);
nor U3786 (N_3786,In_649,In_971);
nor U3787 (N_3787,In_61,In_338);
nand U3788 (N_3788,In_397,In_649);
xnor U3789 (N_3789,In_841,In_325);
nor U3790 (N_3790,In_630,In_467);
nor U3791 (N_3791,In_625,In_992);
xnor U3792 (N_3792,In_153,In_241);
or U3793 (N_3793,In_292,In_24);
nor U3794 (N_3794,In_23,In_331);
nor U3795 (N_3795,In_451,In_889);
xnor U3796 (N_3796,In_286,In_892);
nor U3797 (N_3797,In_87,In_831);
and U3798 (N_3798,In_39,In_885);
or U3799 (N_3799,In_830,In_568);
or U3800 (N_3800,In_127,In_879);
nor U3801 (N_3801,In_700,In_934);
xor U3802 (N_3802,In_103,In_600);
nor U3803 (N_3803,In_613,In_336);
nor U3804 (N_3804,In_626,In_574);
or U3805 (N_3805,In_638,In_325);
nor U3806 (N_3806,In_244,In_217);
and U3807 (N_3807,In_931,In_553);
xnor U3808 (N_3808,In_710,In_474);
or U3809 (N_3809,In_917,In_954);
and U3810 (N_3810,In_867,In_831);
or U3811 (N_3811,In_330,In_112);
and U3812 (N_3812,In_485,In_168);
or U3813 (N_3813,In_632,In_821);
and U3814 (N_3814,In_436,In_935);
nand U3815 (N_3815,In_148,In_573);
xnor U3816 (N_3816,In_590,In_766);
or U3817 (N_3817,In_545,In_727);
xnor U3818 (N_3818,In_503,In_939);
nand U3819 (N_3819,In_741,In_854);
nor U3820 (N_3820,In_615,In_439);
or U3821 (N_3821,In_82,In_0);
nand U3822 (N_3822,In_278,In_821);
and U3823 (N_3823,In_581,In_840);
and U3824 (N_3824,In_980,In_334);
xnor U3825 (N_3825,In_534,In_845);
nor U3826 (N_3826,In_343,In_221);
or U3827 (N_3827,In_635,In_434);
and U3828 (N_3828,In_252,In_795);
nand U3829 (N_3829,In_153,In_600);
xor U3830 (N_3830,In_970,In_414);
or U3831 (N_3831,In_975,In_767);
xnor U3832 (N_3832,In_428,In_989);
nand U3833 (N_3833,In_849,In_853);
and U3834 (N_3834,In_517,In_714);
nand U3835 (N_3835,In_31,In_61);
xor U3836 (N_3836,In_10,In_497);
and U3837 (N_3837,In_274,In_26);
nand U3838 (N_3838,In_792,In_328);
xor U3839 (N_3839,In_360,In_420);
or U3840 (N_3840,In_737,In_704);
nor U3841 (N_3841,In_16,In_35);
nand U3842 (N_3842,In_179,In_602);
nor U3843 (N_3843,In_298,In_758);
nand U3844 (N_3844,In_84,In_236);
nand U3845 (N_3845,In_290,In_234);
or U3846 (N_3846,In_405,In_203);
nand U3847 (N_3847,In_944,In_824);
nand U3848 (N_3848,In_775,In_237);
nor U3849 (N_3849,In_239,In_21);
nor U3850 (N_3850,In_54,In_917);
xnor U3851 (N_3851,In_817,In_619);
nor U3852 (N_3852,In_683,In_553);
nor U3853 (N_3853,In_680,In_592);
nand U3854 (N_3854,In_645,In_454);
and U3855 (N_3855,In_939,In_408);
nor U3856 (N_3856,In_231,In_416);
and U3857 (N_3857,In_655,In_981);
or U3858 (N_3858,In_914,In_108);
nand U3859 (N_3859,In_260,In_504);
nor U3860 (N_3860,In_734,In_278);
xor U3861 (N_3861,In_751,In_199);
nand U3862 (N_3862,In_673,In_560);
nand U3863 (N_3863,In_939,In_267);
or U3864 (N_3864,In_291,In_463);
nor U3865 (N_3865,In_464,In_533);
or U3866 (N_3866,In_424,In_99);
nand U3867 (N_3867,In_419,In_429);
or U3868 (N_3868,In_881,In_490);
xor U3869 (N_3869,In_53,In_692);
xnor U3870 (N_3870,In_819,In_470);
and U3871 (N_3871,In_980,In_131);
or U3872 (N_3872,In_38,In_684);
xnor U3873 (N_3873,In_268,In_721);
xnor U3874 (N_3874,In_518,In_289);
nor U3875 (N_3875,In_700,In_250);
xor U3876 (N_3876,In_766,In_421);
nand U3877 (N_3877,In_342,In_354);
xnor U3878 (N_3878,In_775,In_245);
xnor U3879 (N_3879,In_926,In_404);
nor U3880 (N_3880,In_93,In_352);
nand U3881 (N_3881,In_261,In_166);
or U3882 (N_3882,In_644,In_348);
or U3883 (N_3883,In_866,In_168);
and U3884 (N_3884,In_933,In_503);
xor U3885 (N_3885,In_992,In_773);
nand U3886 (N_3886,In_797,In_159);
nand U3887 (N_3887,In_345,In_528);
or U3888 (N_3888,In_895,In_362);
xor U3889 (N_3889,In_138,In_667);
nor U3890 (N_3890,In_369,In_704);
xor U3891 (N_3891,In_743,In_863);
nand U3892 (N_3892,In_939,In_68);
and U3893 (N_3893,In_729,In_935);
nor U3894 (N_3894,In_975,In_653);
xnor U3895 (N_3895,In_104,In_15);
or U3896 (N_3896,In_422,In_952);
nor U3897 (N_3897,In_193,In_268);
and U3898 (N_3898,In_340,In_740);
xnor U3899 (N_3899,In_779,In_288);
or U3900 (N_3900,In_271,In_333);
nand U3901 (N_3901,In_815,In_319);
nor U3902 (N_3902,In_902,In_802);
nor U3903 (N_3903,In_471,In_423);
or U3904 (N_3904,In_19,In_845);
nor U3905 (N_3905,In_712,In_676);
and U3906 (N_3906,In_336,In_832);
and U3907 (N_3907,In_476,In_522);
xnor U3908 (N_3908,In_647,In_279);
nand U3909 (N_3909,In_789,In_552);
nand U3910 (N_3910,In_775,In_114);
nand U3911 (N_3911,In_708,In_503);
xnor U3912 (N_3912,In_712,In_653);
xor U3913 (N_3913,In_99,In_718);
nor U3914 (N_3914,In_293,In_925);
or U3915 (N_3915,In_202,In_96);
or U3916 (N_3916,In_950,In_631);
xnor U3917 (N_3917,In_841,In_598);
xor U3918 (N_3918,In_830,In_328);
xor U3919 (N_3919,In_553,In_623);
nand U3920 (N_3920,In_577,In_754);
xnor U3921 (N_3921,In_417,In_874);
and U3922 (N_3922,In_507,In_206);
nor U3923 (N_3923,In_389,In_328);
or U3924 (N_3924,In_943,In_938);
or U3925 (N_3925,In_376,In_238);
xor U3926 (N_3926,In_335,In_132);
xnor U3927 (N_3927,In_467,In_414);
xor U3928 (N_3928,In_610,In_70);
and U3929 (N_3929,In_727,In_680);
nor U3930 (N_3930,In_363,In_106);
nand U3931 (N_3931,In_525,In_620);
and U3932 (N_3932,In_868,In_381);
nand U3933 (N_3933,In_947,In_225);
nand U3934 (N_3934,In_999,In_294);
nor U3935 (N_3935,In_938,In_322);
nor U3936 (N_3936,In_337,In_289);
xor U3937 (N_3937,In_255,In_959);
nand U3938 (N_3938,In_563,In_272);
xnor U3939 (N_3939,In_406,In_98);
nor U3940 (N_3940,In_807,In_653);
nor U3941 (N_3941,In_946,In_427);
and U3942 (N_3942,In_79,In_191);
or U3943 (N_3943,In_634,In_896);
or U3944 (N_3944,In_272,In_338);
nand U3945 (N_3945,In_552,In_555);
nor U3946 (N_3946,In_888,In_262);
and U3947 (N_3947,In_322,In_292);
nor U3948 (N_3948,In_628,In_917);
and U3949 (N_3949,In_2,In_50);
or U3950 (N_3950,In_158,In_678);
nand U3951 (N_3951,In_364,In_716);
or U3952 (N_3952,In_239,In_34);
xnor U3953 (N_3953,In_847,In_35);
nor U3954 (N_3954,In_226,In_82);
nand U3955 (N_3955,In_122,In_188);
and U3956 (N_3956,In_679,In_639);
xnor U3957 (N_3957,In_27,In_745);
xnor U3958 (N_3958,In_62,In_994);
nor U3959 (N_3959,In_854,In_675);
nand U3960 (N_3960,In_217,In_26);
and U3961 (N_3961,In_778,In_968);
and U3962 (N_3962,In_770,In_17);
xnor U3963 (N_3963,In_873,In_781);
xor U3964 (N_3964,In_310,In_497);
and U3965 (N_3965,In_199,In_216);
nor U3966 (N_3966,In_471,In_903);
nor U3967 (N_3967,In_800,In_446);
or U3968 (N_3968,In_748,In_62);
nor U3969 (N_3969,In_228,In_976);
or U3970 (N_3970,In_228,In_454);
nand U3971 (N_3971,In_480,In_979);
xnor U3972 (N_3972,In_482,In_858);
and U3973 (N_3973,In_898,In_213);
nor U3974 (N_3974,In_51,In_438);
xor U3975 (N_3975,In_596,In_517);
xnor U3976 (N_3976,In_290,In_632);
nand U3977 (N_3977,In_862,In_140);
xor U3978 (N_3978,In_325,In_173);
nor U3979 (N_3979,In_107,In_997);
and U3980 (N_3980,In_199,In_352);
nand U3981 (N_3981,In_966,In_27);
nand U3982 (N_3982,In_698,In_136);
and U3983 (N_3983,In_160,In_303);
or U3984 (N_3984,In_978,In_138);
and U3985 (N_3985,In_650,In_448);
or U3986 (N_3986,In_821,In_33);
nand U3987 (N_3987,In_667,In_237);
nand U3988 (N_3988,In_6,In_866);
nor U3989 (N_3989,In_960,In_247);
xor U3990 (N_3990,In_671,In_261);
and U3991 (N_3991,In_14,In_543);
and U3992 (N_3992,In_791,In_774);
or U3993 (N_3993,In_261,In_561);
or U3994 (N_3994,In_361,In_466);
nand U3995 (N_3995,In_620,In_236);
xor U3996 (N_3996,In_805,In_585);
xnor U3997 (N_3997,In_706,In_813);
nand U3998 (N_3998,In_557,In_886);
nand U3999 (N_3999,In_808,In_322);
nor U4000 (N_4000,In_54,In_852);
xnor U4001 (N_4001,In_443,In_620);
and U4002 (N_4002,In_664,In_839);
nor U4003 (N_4003,In_969,In_369);
nand U4004 (N_4004,In_761,In_182);
nand U4005 (N_4005,In_728,In_216);
xor U4006 (N_4006,In_996,In_948);
nand U4007 (N_4007,In_518,In_555);
xor U4008 (N_4008,In_441,In_739);
nor U4009 (N_4009,In_452,In_291);
nand U4010 (N_4010,In_835,In_910);
nor U4011 (N_4011,In_828,In_509);
nand U4012 (N_4012,In_443,In_784);
nor U4013 (N_4013,In_360,In_262);
and U4014 (N_4014,In_679,In_411);
xnor U4015 (N_4015,In_27,In_614);
nand U4016 (N_4016,In_515,In_791);
and U4017 (N_4017,In_250,In_574);
nor U4018 (N_4018,In_468,In_862);
xnor U4019 (N_4019,In_876,In_862);
nor U4020 (N_4020,In_657,In_502);
nand U4021 (N_4021,In_665,In_320);
nor U4022 (N_4022,In_129,In_498);
or U4023 (N_4023,In_739,In_391);
xor U4024 (N_4024,In_773,In_814);
and U4025 (N_4025,In_162,In_198);
nand U4026 (N_4026,In_557,In_72);
nor U4027 (N_4027,In_321,In_425);
xor U4028 (N_4028,In_704,In_412);
or U4029 (N_4029,In_668,In_477);
xnor U4030 (N_4030,In_173,In_378);
xor U4031 (N_4031,In_333,In_629);
xnor U4032 (N_4032,In_966,In_79);
nor U4033 (N_4033,In_629,In_424);
nor U4034 (N_4034,In_166,In_790);
and U4035 (N_4035,In_221,In_564);
xor U4036 (N_4036,In_399,In_121);
and U4037 (N_4037,In_731,In_96);
and U4038 (N_4038,In_197,In_439);
and U4039 (N_4039,In_630,In_933);
nand U4040 (N_4040,In_263,In_60);
nand U4041 (N_4041,In_579,In_764);
xnor U4042 (N_4042,In_404,In_800);
xor U4043 (N_4043,In_332,In_718);
xor U4044 (N_4044,In_12,In_348);
and U4045 (N_4045,In_200,In_824);
and U4046 (N_4046,In_395,In_350);
xor U4047 (N_4047,In_975,In_271);
nor U4048 (N_4048,In_224,In_887);
and U4049 (N_4049,In_794,In_928);
or U4050 (N_4050,In_555,In_768);
and U4051 (N_4051,In_524,In_95);
xnor U4052 (N_4052,In_791,In_670);
nor U4053 (N_4053,In_50,In_403);
xor U4054 (N_4054,In_328,In_119);
nor U4055 (N_4055,In_301,In_118);
xor U4056 (N_4056,In_575,In_475);
or U4057 (N_4057,In_439,In_669);
nand U4058 (N_4058,In_451,In_976);
xor U4059 (N_4059,In_648,In_419);
or U4060 (N_4060,In_986,In_521);
and U4061 (N_4061,In_788,In_56);
xnor U4062 (N_4062,In_258,In_12);
and U4063 (N_4063,In_256,In_711);
or U4064 (N_4064,In_781,In_34);
and U4065 (N_4065,In_673,In_267);
nor U4066 (N_4066,In_456,In_695);
xnor U4067 (N_4067,In_711,In_357);
and U4068 (N_4068,In_905,In_949);
nand U4069 (N_4069,In_256,In_404);
and U4070 (N_4070,In_214,In_330);
or U4071 (N_4071,In_444,In_37);
xor U4072 (N_4072,In_458,In_394);
nor U4073 (N_4073,In_917,In_81);
and U4074 (N_4074,In_189,In_910);
xnor U4075 (N_4075,In_501,In_723);
xnor U4076 (N_4076,In_580,In_298);
xor U4077 (N_4077,In_412,In_871);
xnor U4078 (N_4078,In_265,In_321);
nor U4079 (N_4079,In_284,In_797);
xor U4080 (N_4080,In_18,In_742);
nand U4081 (N_4081,In_205,In_160);
and U4082 (N_4082,In_141,In_830);
and U4083 (N_4083,In_429,In_106);
or U4084 (N_4084,In_578,In_302);
nand U4085 (N_4085,In_347,In_725);
nand U4086 (N_4086,In_977,In_687);
nand U4087 (N_4087,In_507,In_335);
nor U4088 (N_4088,In_170,In_639);
or U4089 (N_4089,In_458,In_117);
and U4090 (N_4090,In_301,In_884);
nor U4091 (N_4091,In_949,In_256);
nand U4092 (N_4092,In_718,In_699);
xor U4093 (N_4093,In_680,In_447);
and U4094 (N_4094,In_309,In_15);
nor U4095 (N_4095,In_366,In_791);
nor U4096 (N_4096,In_815,In_115);
xor U4097 (N_4097,In_118,In_138);
or U4098 (N_4098,In_994,In_320);
nor U4099 (N_4099,In_646,In_220);
xnor U4100 (N_4100,In_893,In_235);
nor U4101 (N_4101,In_479,In_156);
and U4102 (N_4102,In_366,In_959);
nand U4103 (N_4103,In_994,In_617);
nor U4104 (N_4104,In_114,In_346);
nand U4105 (N_4105,In_16,In_203);
nand U4106 (N_4106,In_311,In_20);
and U4107 (N_4107,In_687,In_365);
nor U4108 (N_4108,In_329,In_989);
nand U4109 (N_4109,In_753,In_238);
xor U4110 (N_4110,In_829,In_601);
nor U4111 (N_4111,In_400,In_252);
xnor U4112 (N_4112,In_363,In_639);
xnor U4113 (N_4113,In_664,In_163);
and U4114 (N_4114,In_930,In_917);
nand U4115 (N_4115,In_177,In_577);
or U4116 (N_4116,In_61,In_763);
xor U4117 (N_4117,In_168,In_836);
and U4118 (N_4118,In_410,In_870);
xnor U4119 (N_4119,In_744,In_534);
or U4120 (N_4120,In_784,In_503);
and U4121 (N_4121,In_895,In_104);
nor U4122 (N_4122,In_567,In_272);
and U4123 (N_4123,In_664,In_695);
xor U4124 (N_4124,In_359,In_228);
and U4125 (N_4125,In_116,In_162);
and U4126 (N_4126,In_539,In_350);
nor U4127 (N_4127,In_256,In_561);
and U4128 (N_4128,In_971,In_881);
nand U4129 (N_4129,In_507,In_217);
xor U4130 (N_4130,In_699,In_601);
nand U4131 (N_4131,In_402,In_380);
and U4132 (N_4132,In_390,In_67);
xnor U4133 (N_4133,In_770,In_637);
or U4134 (N_4134,In_878,In_567);
or U4135 (N_4135,In_928,In_207);
xnor U4136 (N_4136,In_800,In_797);
and U4137 (N_4137,In_770,In_669);
nand U4138 (N_4138,In_927,In_670);
nand U4139 (N_4139,In_414,In_341);
xor U4140 (N_4140,In_974,In_311);
or U4141 (N_4141,In_336,In_934);
or U4142 (N_4142,In_497,In_422);
or U4143 (N_4143,In_757,In_213);
nor U4144 (N_4144,In_853,In_503);
xor U4145 (N_4145,In_195,In_822);
xor U4146 (N_4146,In_79,In_684);
nor U4147 (N_4147,In_937,In_955);
and U4148 (N_4148,In_606,In_685);
or U4149 (N_4149,In_412,In_671);
nor U4150 (N_4150,In_996,In_245);
xnor U4151 (N_4151,In_428,In_819);
and U4152 (N_4152,In_920,In_205);
nor U4153 (N_4153,In_808,In_670);
nand U4154 (N_4154,In_270,In_716);
and U4155 (N_4155,In_872,In_459);
nor U4156 (N_4156,In_600,In_822);
or U4157 (N_4157,In_751,In_232);
and U4158 (N_4158,In_769,In_50);
or U4159 (N_4159,In_884,In_940);
and U4160 (N_4160,In_324,In_407);
nand U4161 (N_4161,In_218,In_462);
nor U4162 (N_4162,In_395,In_497);
nand U4163 (N_4163,In_66,In_886);
or U4164 (N_4164,In_458,In_82);
and U4165 (N_4165,In_734,In_517);
or U4166 (N_4166,In_583,In_400);
nand U4167 (N_4167,In_172,In_330);
nand U4168 (N_4168,In_929,In_441);
nor U4169 (N_4169,In_51,In_583);
or U4170 (N_4170,In_711,In_627);
nand U4171 (N_4171,In_850,In_199);
xnor U4172 (N_4172,In_665,In_879);
xor U4173 (N_4173,In_391,In_920);
and U4174 (N_4174,In_865,In_571);
and U4175 (N_4175,In_14,In_198);
and U4176 (N_4176,In_607,In_38);
or U4177 (N_4177,In_264,In_491);
nand U4178 (N_4178,In_238,In_498);
and U4179 (N_4179,In_169,In_455);
nand U4180 (N_4180,In_658,In_322);
or U4181 (N_4181,In_932,In_806);
xnor U4182 (N_4182,In_855,In_380);
or U4183 (N_4183,In_718,In_982);
and U4184 (N_4184,In_734,In_47);
xor U4185 (N_4185,In_655,In_240);
nand U4186 (N_4186,In_871,In_421);
nor U4187 (N_4187,In_173,In_695);
xnor U4188 (N_4188,In_612,In_119);
and U4189 (N_4189,In_339,In_473);
or U4190 (N_4190,In_642,In_935);
or U4191 (N_4191,In_516,In_811);
or U4192 (N_4192,In_457,In_869);
or U4193 (N_4193,In_938,In_856);
or U4194 (N_4194,In_596,In_61);
nand U4195 (N_4195,In_11,In_590);
or U4196 (N_4196,In_228,In_490);
nor U4197 (N_4197,In_474,In_536);
nor U4198 (N_4198,In_533,In_992);
xnor U4199 (N_4199,In_966,In_216);
nand U4200 (N_4200,In_728,In_678);
nand U4201 (N_4201,In_768,In_169);
and U4202 (N_4202,In_947,In_131);
and U4203 (N_4203,In_723,In_751);
or U4204 (N_4204,In_644,In_151);
and U4205 (N_4205,In_125,In_254);
nand U4206 (N_4206,In_854,In_554);
or U4207 (N_4207,In_477,In_417);
xnor U4208 (N_4208,In_266,In_483);
nand U4209 (N_4209,In_484,In_259);
nor U4210 (N_4210,In_631,In_301);
and U4211 (N_4211,In_339,In_512);
xnor U4212 (N_4212,In_563,In_546);
nand U4213 (N_4213,In_612,In_585);
xor U4214 (N_4214,In_884,In_504);
nand U4215 (N_4215,In_22,In_459);
nand U4216 (N_4216,In_974,In_812);
nor U4217 (N_4217,In_680,In_205);
nand U4218 (N_4218,In_585,In_977);
or U4219 (N_4219,In_701,In_720);
or U4220 (N_4220,In_869,In_671);
nor U4221 (N_4221,In_111,In_773);
and U4222 (N_4222,In_172,In_953);
and U4223 (N_4223,In_563,In_821);
or U4224 (N_4224,In_783,In_301);
xnor U4225 (N_4225,In_388,In_873);
and U4226 (N_4226,In_332,In_659);
or U4227 (N_4227,In_891,In_695);
nor U4228 (N_4228,In_97,In_301);
and U4229 (N_4229,In_703,In_900);
xor U4230 (N_4230,In_642,In_364);
and U4231 (N_4231,In_658,In_347);
nor U4232 (N_4232,In_828,In_977);
or U4233 (N_4233,In_936,In_763);
nor U4234 (N_4234,In_89,In_409);
or U4235 (N_4235,In_123,In_849);
nand U4236 (N_4236,In_874,In_640);
nand U4237 (N_4237,In_655,In_659);
and U4238 (N_4238,In_81,In_791);
and U4239 (N_4239,In_485,In_966);
xor U4240 (N_4240,In_838,In_811);
xnor U4241 (N_4241,In_561,In_217);
nand U4242 (N_4242,In_626,In_890);
xnor U4243 (N_4243,In_352,In_811);
nand U4244 (N_4244,In_504,In_58);
or U4245 (N_4245,In_754,In_66);
or U4246 (N_4246,In_840,In_824);
and U4247 (N_4247,In_42,In_271);
nand U4248 (N_4248,In_220,In_636);
or U4249 (N_4249,In_267,In_709);
and U4250 (N_4250,In_862,In_33);
or U4251 (N_4251,In_434,In_854);
nand U4252 (N_4252,In_7,In_851);
nor U4253 (N_4253,In_77,In_923);
and U4254 (N_4254,In_578,In_528);
and U4255 (N_4255,In_978,In_117);
nor U4256 (N_4256,In_785,In_645);
or U4257 (N_4257,In_98,In_103);
xnor U4258 (N_4258,In_600,In_156);
and U4259 (N_4259,In_380,In_894);
nor U4260 (N_4260,In_459,In_598);
and U4261 (N_4261,In_408,In_415);
and U4262 (N_4262,In_637,In_108);
xor U4263 (N_4263,In_72,In_697);
nand U4264 (N_4264,In_81,In_302);
and U4265 (N_4265,In_467,In_174);
nor U4266 (N_4266,In_935,In_469);
xor U4267 (N_4267,In_157,In_448);
xor U4268 (N_4268,In_710,In_396);
and U4269 (N_4269,In_896,In_100);
nor U4270 (N_4270,In_664,In_426);
xor U4271 (N_4271,In_520,In_92);
xnor U4272 (N_4272,In_517,In_310);
xnor U4273 (N_4273,In_7,In_116);
or U4274 (N_4274,In_431,In_538);
and U4275 (N_4275,In_68,In_772);
or U4276 (N_4276,In_974,In_876);
or U4277 (N_4277,In_201,In_682);
or U4278 (N_4278,In_792,In_389);
and U4279 (N_4279,In_765,In_516);
and U4280 (N_4280,In_702,In_253);
xor U4281 (N_4281,In_896,In_863);
xnor U4282 (N_4282,In_766,In_531);
or U4283 (N_4283,In_815,In_333);
nand U4284 (N_4284,In_145,In_973);
or U4285 (N_4285,In_768,In_120);
nand U4286 (N_4286,In_516,In_202);
or U4287 (N_4287,In_218,In_609);
nor U4288 (N_4288,In_186,In_841);
and U4289 (N_4289,In_810,In_747);
and U4290 (N_4290,In_189,In_640);
xor U4291 (N_4291,In_779,In_826);
nand U4292 (N_4292,In_110,In_482);
and U4293 (N_4293,In_582,In_669);
nor U4294 (N_4294,In_523,In_262);
nor U4295 (N_4295,In_312,In_362);
or U4296 (N_4296,In_394,In_59);
and U4297 (N_4297,In_795,In_170);
and U4298 (N_4298,In_678,In_572);
xnor U4299 (N_4299,In_59,In_430);
nor U4300 (N_4300,In_77,In_967);
or U4301 (N_4301,In_236,In_229);
or U4302 (N_4302,In_851,In_48);
xnor U4303 (N_4303,In_919,In_971);
nand U4304 (N_4304,In_894,In_689);
nor U4305 (N_4305,In_809,In_785);
xor U4306 (N_4306,In_820,In_541);
nand U4307 (N_4307,In_129,In_871);
nand U4308 (N_4308,In_978,In_845);
or U4309 (N_4309,In_259,In_395);
or U4310 (N_4310,In_670,In_768);
or U4311 (N_4311,In_415,In_229);
nand U4312 (N_4312,In_837,In_620);
xnor U4313 (N_4313,In_268,In_463);
and U4314 (N_4314,In_988,In_715);
and U4315 (N_4315,In_15,In_832);
and U4316 (N_4316,In_867,In_566);
nor U4317 (N_4317,In_801,In_953);
nor U4318 (N_4318,In_345,In_233);
nand U4319 (N_4319,In_234,In_813);
nor U4320 (N_4320,In_416,In_606);
nand U4321 (N_4321,In_176,In_397);
or U4322 (N_4322,In_910,In_967);
or U4323 (N_4323,In_706,In_775);
or U4324 (N_4324,In_845,In_831);
or U4325 (N_4325,In_292,In_165);
nor U4326 (N_4326,In_147,In_94);
nor U4327 (N_4327,In_746,In_167);
nand U4328 (N_4328,In_867,In_878);
xor U4329 (N_4329,In_410,In_164);
nand U4330 (N_4330,In_189,In_514);
nand U4331 (N_4331,In_660,In_663);
nor U4332 (N_4332,In_17,In_396);
nor U4333 (N_4333,In_767,In_810);
or U4334 (N_4334,In_766,In_247);
nor U4335 (N_4335,In_810,In_449);
nand U4336 (N_4336,In_671,In_702);
nor U4337 (N_4337,In_720,In_547);
xnor U4338 (N_4338,In_402,In_384);
nand U4339 (N_4339,In_60,In_211);
nand U4340 (N_4340,In_62,In_896);
and U4341 (N_4341,In_590,In_64);
nor U4342 (N_4342,In_186,In_743);
xor U4343 (N_4343,In_314,In_383);
or U4344 (N_4344,In_11,In_150);
and U4345 (N_4345,In_75,In_99);
nand U4346 (N_4346,In_188,In_107);
xnor U4347 (N_4347,In_385,In_601);
or U4348 (N_4348,In_363,In_762);
nand U4349 (N_4349,In_325,In_528);
and U4350 (N_4350,In_794,In_812);
xor U4351 (N_4351,In_152,In_667);
or U4352 (N_4352,In_680,In_342);
nand U4353 (N_4353,In_571,In_86);
and U4354 (N_4354,In_354,In_838);
and U4355 (N_4355,In_542,In_352);
xor U4356 (N_4356,In_631,In_582);
xor U4357 (N_4357,In_801,In_742);
nor U4358 (N_4358,In_14,In_325);
xnor U4359 (N_4359,In_426,In_698);
nor U4360 (N_4360,In_113,In_882);
nand U4361 (N_4361,In_606,In_591);
xor U4362 (N_4362,In_539,In_813);
nor U4363 (N_4363,In_318,In_16);
nor U4364 (N_4364,In_547,In_808);
and U4365 (N_4365,In_460,In_742);
nand U4366 (N_4366,In_895,In_155);
and U4367 (N_4367,In_744,In_510);
nor U4368 (N_4368,In_124,In_122);
nand U4369 (N_4369,In_657,In_422);
and U4370 (N_4370,In_254,In_762);
xor U4371 (N_4371,In_653,In_722);
or U4372 (N_4372,In_714,In_999);
and U4373 (N_4373,In_372,In_724);
xor U4374 (N_4374,In_687,In_658);
xnor U4375 (N_4375,In_842,In_903);
or U4376 (N_4376,In_588,In_438);
nor U4377 (N_4377,In_8,In_191);
and U4378 (N_4378,In_426,In_2);
and U4379 (N_4379,In_505,In_294);
nand U4380 (N_4380,In_649,In_685);
xor U4381 (N_4381,In_240,In_832);
or U4382 (N_4382,In_257,In_50);
nand U4383 (N_4383,In_524,In_35);
nand U4384 (N_4384,In_21,In_850);
nor U4385 (N_4385,In_671,In_982);
and U4386 (N_4386,In_575,In_48);
xnor U4387 (N_4387,In_586,In_35);
xor U4388 (N_4388,In_418,In_559);
xor U4389 (N_4389,In_387,In_881);
and U4390 (N_4390,In_904,In_772);
and U4391 (N_4391,In_679,In_856);
and U4392 (N_4392,In_944,In_621);
nand U4393 (N_4393,In_673,In_502);
nand U4394 (N_4394,In_816,In_551);
nand U4395 (N_4395,In_371,In_553);
nor U4396 (N_4396,In_838,In_476);
or U4397 (N_4397,In_276,In_923);
nand U4398 (N_4398,In_305,In_290);
nand U4399 (N_4399,In_842,In_387);
nand U4400 (N_4400,In_344,In_669);
xor U4401 (N_4401,In_928,In_517);
xnor U4402 (N_4402,In_919,In_344);
nand U4403 (N_4403,In_777,In_934);
xor U4404 (N_4404,In_820,In_916);
or U4405 (N_4405,In_434,In_636);
nand U4406 (N_4406,In_738,In_866);
and U4407 (N_4407,In_973,In_450);
and U4408 (N_4408,In_509,In_218);
or U4409 (N_4409,In_5,In_438);
or U4410 (N_4410,In_732,In_980);
nor U4411 (N_4411,In_132,In_183);
or U4412 (N_4412,In_373,In_739);
and U4413 (N_4413,In_988,In_724);
nand U4414 (N_4414,In_440,In_735);
nor U4415 (N_4415,In_959,In_106);
nor U4416 (N_4416,In_271,In_81);
xor U4417 (N_4417,In_269,In_416);
xor U4418 (N_4418,In_136,In_839);
or U4419 (N_4419,In_24,In_679);
nor U4420 (N_4420,In_477,In_245);
nand U4421 (N_4421,In_717,In_943);
or U4422 (N_4422,In_370,In_57);
xor U4423 (N_4423,In_385,In_558);
xnor U4424 (N_4424,In_43,In_560);
and U4425 (N_4425,In_505,In_766);
and U4426 (N_4426,In_505,In_862);
nor U4427 (N_4427,In_923,In_412);
nand U4428 (N_4428,In_681,In_940);
and U4429 (N_4429,In_610,In_505);
xor U4430 (N_4430,In_378,In_324);
xor U4431 (N_4431,In_323,In_657);
and U4432 (N_4432,In_135,In_794);
xnor U4433 (N_4433,In_607,In_130);
nand U4434 (N_4434,In_873,In_410);
or U4435 (N_4435,In_877,In_931);
nand U4436 (N_4436,In_979,In_315);
nor U4437 (N_4437,In_322,In_487);
xnor U4438 (N_4438,In_199,In_101);
xor U4439 (N_4439,In_135,In_479);
or U4440 (N_4440,In_6,In_93);
nand U4441 (N_4441,In_137,In_480);
nand U4442 (N_4442,In_994,In_968);
and U4443 (N_4443,In_991,In_172);
or U4444 (N_4444,In_750,In_807);
and U4445 (N_4445,In_829,In_531);
xor U4446 (N_4446,In_320,In_237);
and U4447 (N_4447,In_605,In_403);
nor U4448 (N_4448,In_65,In_86);
or U4449 (N_4449,In_269,In_965);
xnor U4450 (N_4450,In_112,In_359);
and U4451 (N_4451,In_554,In_640);
or U4452 (N_4452,In_315,In_845);
nand U4453 (N_4453,In_286,In_434);
or U4454 (N_4454,In_225,In_569);
nand U4455 (N_4455,In_617,In_769);
nand U4456 (N_4456,In_358,In_866);
and U4457 (N_4457,In_447,In_610);
and U4458 (N_4458,In_928,In_249);
and U4459 (N_4459,In_676,In_956);
nor U4460 (N_4460,In_762,In_605);
or U4461 (N_4461,In_911,In_959);
nand U4462 (N_4462,In_888,In_602);
or U4463 (N_4463,In_708,In_223);
xor U4464 (N_4464,In_328,In_117);
and U4465 (N_4465,In_888,In_41);
nor U4466 (N_4466,In_208,In_488);
and U4467 (N_4467,In_626,In_812);
and U4468 (N_4468,In_460,In_942);
nor U4469 (N_4469,In_233,In_224);
nor U4470 (N_4470,In_536,In_166);
nand U4471 (N_4471,In_461,In_640);
and U4472 (N_4472,In_115,In_874);
nand U4473 (N_4473,In_847,In_919);
or U4474 (N_4474,In_467,In_380);
nor U4475 (N_4475,In_386,In_800);
or U4476 (N_4476,In_422,In_443);
nand U4477 (N_4477,In_13,In_922);
nor U4478 (N_4478,In_273,In_277);
or U4479 (N_4479,In_561,In_879);
nor U4480 (N_4480,In_967,In_52);
and U4481 (N_4481,In_790,In_729);
xnor U4482 (N_4482,In_986,In_341);
and U4483 (N_4483,In_149,In_955);
nor U4484 (N_4484,In_635,In_756);
nor U4485 (N_4485,In_539,In_300);
xor U4486 (N_4486,In_155,In_900);
nor U4487 (N_4487,In_309,In_147);
nor U4488 (N_4488,In_909,In_985);
or U4489 (N_4489,In_972,In_120);
and U4490 (N_4490,In_366,In_316);
and U4491 (N_4491,In_813,In_893);
xnor U4492 (N_4492,In_574,In_720);
and U4493 (N_4493,In_270,In_772);
xor U4494 (N_4494,In_957,In_810);
or U4495 (N_4495,In_818,In_259);
and U4496 (N_4496,In_479,In_530);
nor U4497 (N_4497,In_258,In_197);
xnor U4498 (N_4498,In_777,In_613);
or U4499 (N_4499,In_205,In_309);
or U4500 (N_4500,In_272,In_239);
nand U4501 (N_4501,In_280,In_298);
and U4502 (N_4502,In_589,In_433);
or U4503 (N_4503,In_475,In_190);
and U4504 (N_4504,In_428,In_195);
or U4505 (N_4505,In_764,In_349);
nand U4506 (N_4506,In_553,In_19);
and U4507 (N_4507,In_510,In_269);
and U4508 (N_4508,In_11,In_536);
nor U4509 (N_4509,In_468,In_295);
nand U4510 (N_4510,In_319,In_222);
nor U4511 (N_4511,In_684,In_225);
and U4512 (N_4512,In_259,In_788);
xor U4513 (N_4513,In_748,In_290);
or U4514 (N_4514,In_941,In_63);
nand U4515 (N_4515,In_423,In_62);
or U4516 (N_4516,In_167,In_530);
xnor U4517 (N_4517,In_231,In_330);
and U4518 (N_4518,In_912,In_646);
and U4519 (N_4519,In_533,In_420);
and U4520 (N_4520,In_590,In_356);
or U4521 (N_4521,In_130,In_345);
xor U4522 (N_4522,In_696,In_594);
and U4523 (N_4523,In_550,In_973);
and U4524 (N_4524,In_565,In_788);
or U4525 (N_4525,In_893,In_298);
and U4526 (N_4526,In_539,In_686);
nor U4527 (N_4527,In_790,In_737);
and U4528 (N_4528,In_90,In_771);
or U4529 (N_4529,In_220,In_121);
nor U4530 (N_4530,In_704,In_919);
nand U4531 (N_4531,In_18,In_635);
nor U4532 (N_4532,In_292,In_20);
or U4533 (N_4533,In_721,In_389);
xnor U4534 (N_4534,In_337,In_669);
or U4535 (N_4535,In_844,In_433);
or U4536 (N_4536,In_79,In_349);
xor U4537 (N_4537,In_894,In_899);
and U4538 (N_4538,In_604,In_430);
and U4539 (N_4539,In_984,In_287);
or U4540 (N_4540,In_276,In_869);
nor U4541 (N_4541,In_52,In_445);
nand U4542 (N_4542,In_941,In_703);
or U4543 (N_4543,In_303,In_273);
and U4544 (N_4544,In_990,In_152);
nor U4545 (N_4545,In_40,In_317);
nor U4546 (N_4546,In_704,In_839);
nand U4547 (N_4547,In_532,In_433);
nor U4548 (N_4548,In_152,In_774);
nand U4549 (N_4549,In_124,In_774);
or U4550 (N_4550,In_4,In_366);
nand U4551 (N_4551,In_972,In_659);
and U4552 (N_4552,In_628,In_906);
nand U4553 (N_4553,In_451,In_759);
and U4554 (N_4554,In_778,In_113);
nor U4555 (N_4555,In_751,In_644);
or U4556 (N_4556,In_135,In_596);
nor U4557 (N_4557,In_96,In_971);
nand U4558 (N_4558,In_671,In_506);
or U4559 (N_4559,In_740,In_656);
or U4560 (N_4560,In_297,In_33);
and U4561 (N_4561,In_618,In_453);
xor U4562 (N_4562,In_288,In_690);
nand U4563 (N_4563,In_42,In_306);
and U4564 (N_4564,In_983,In_572);
nand U4565 (N_4565,In_747,In_885);
and U4566 (N_4566,In_246,In_129);
and U4567 (N_4567,In_971,In_842);
or U4568 (N_4568,In_846,In_32);
or U4569 (N_4569,In_959,In_511);
xor U4570 (N_4570,In_762,In_399);
nor U4571 (N_4571,In_947,In_592);
nand U4572 (N_4572,In_89,In_60);
nor U4573 (N_4573,In_258,In_200);
and U4574 (N_4574,In_996,In_997);
or U4575 (N_4575,In_17,In_412);
nand U4576 (N_4576,In_585,In_263);
or U4577 (N_4577,In_620,In_77);
or U4578 (N_4578,In_613,In_261);
xnor U4579 (N_4579,In_6,In_429);
nand U4580 (N_4580,In_257,In_383);
nand U4581 (N_4581,In_243,In_756);
nand U4582 (N_4582,In_841,In_675);
xnor U4583 (N_4583,In_205,In_603);
nand U4584 (N_4584,In_189,In_136);
xnor U4585 (N_4585,In_616,In_349);
nor U4586 (N_4586,In_453,In_89);
nor U4587 (N_4587,In_824,In_142);
and U4588 (N_4588,In_221,In_191);
and U4589 (N_4589,In_735,In_394);
xnor U4590 (N_4590,In_192,In_336);
and U4591 (N_4591,In_851,In_939);
or U4592 (N_4592,In_848,In_867);
and U4593 (N_4593,In_717,In_80);
nand U4594 (N_4594,In_955,In_491);
and U4595 (N_4595,In_837,In_576);
nand U4596 (N_4596,In_611,In_294);
xor U4597 (N_4597,In_717,In_559);
and U4598 (N_4598,In_973,In_523);
or U4599 (N_4599,In_111,In_518);
nor U4600 (N_4600,In_29,In_853);
nand U4601 (N_4601,In_942,In_53);
or U4602 (N_4602,In_868,In_401);
and U4603 (N_4603,In_711,In_892);
xnor U4604 (N_4604,In_265,In_226);
nand U4605 (N_4605,In_431,In_423);
and U4606 (N_4606,In_70,In_94);
and U4607 (N_4607,In_578,In_886);
or U4608 (N_4608,In_654,In_460);
nor U4609 (N_4609,In_776,In_140);
nand U4610 (N_4610,In_66,In_75);
and U4611 (N_4611,In_949,In_733);
xnor U4612 (N_4612,In_160,In_300);
xnor U4613 (N_4613,In_737,In_33);
or U4614 (N_4614,In_75,In_50);
nand U4615 (N_4615,In_668,In_521);
nor U4616 (N_4616,In_968,In_414);
nand U4617 (N_4617,In_384,In_152);
nor U4618 (N_4618,In_438,In_820);
nor U4619 (N_4619,In_590,In_176);
or U4620 (N_4620,In_422,In_984);
nor U4621 (N_4621,In_890,In_848);
nor U4622 (N_4622,In_964,In_947);
xnor U4623 (N_4623,In_384,In_92);
nand U4624 (N_4624,In_727,In_353);
or U4625 (N_4625,In_692,In_996);
nand U4626 (N_4626,In_488,In_593);
nor U4627 (N_4627,In_334,In_55);
xnor U4628 (N_4628,In_473,In_102);
xor U4629 (N_4629,In_824,In_989);
and U4630 (N_4630,In_176,In_117);
or U4631 (N_4631,In_559,In_650);
or U4632 (N_4632,In_851,In_300);
xnor U4633 (N_4633,In_925,In_609);
and U4634 (N_4634,In_375,In_983);
and U4635 (N_4635,In_148,In_668);
nor U4636 (N_4636,In_340,In_49);
nor U4637 (N_4637,In_867,In_138);
or U4638 (N_4638,In_309,In_973);
xor U4639 (N_4639,In_336,In_92);
or U4640 (N_4640,In_116,In_945);
xnor U4641 (N_4641,In_638,In_500);
xor U4642 (N_4642,In_882,In_834);
xor U4643 (N_4643,In_474,In_697);
nor U4644 (N_4644,In_806,In_765);
or U4645 (N_4645,In_51,In_530);
nand U4646 (N_4646,In_133,In_938);
and U4647 (N_4647,In_382,In_985);
and U4648 (N_4648,In_939,In_420);
nand U4649 (N_4649,In_420,In_814);
nand U4650 (N_4650,In_433,In_570);
and U4651 (N_4651,In_12,In_550);
or U4652 (N_4652,In_536,In_268);
nand U4653 (N_4653,In_940,In_468);
and U4654 (N_4654,In_605,In_46);
and U4655 (N_4655,In_34,In_735);
and U4656 (N_4656,In_141,In_79);
xor U4657 (N_4657,In_232,In_323);
nor U4658 (N_4658,In_636,In_320);
xnor U4659 (N_4659,In_919,In_822);
nand U4660 (N_4660,In_13,In_127);
nor U4661 (N_4661,In_352,In_142);
nand U4662 (N_4662,In_915,In_52);
xor U4663 (N_4663,In_824,In_801);
and U4664 (N_4664,In_819,In_133);
and U4665 (N_4665,In_402,In_257);
and U4666 (N_4666,In_830,In_608);
xor U4667 (N_4667,In_213,In_32);
or U4668 (N_4668,In_342,In_715);
or U4669 (N_4669,In_918,In_425);
or U4670 (N_4670,In_763,In_564);
or U4671 (N_4671,In_180,In_557);
xnor U4672 (N_4672,In_380,In_475);
nand U4673 (N_4673,In_50,In_61);
nand U4674 (N_4674,In_752,In_140);
and U4675 (N_4675,In_544,In_355);
xnor U4676 (N_4676,In_402,In_8);
nor U4677 (N_4677,In_966,In_83);
nand U4678 (N_4678,In_78,In_806);
and U4679 (N_4679,In_973,In_656);
nand U4680 (N_4680,In_479,In_834);
xnor U4681 (N_4681,In_365,In_468);
nand U4682 (N_4682,In_328,In_704);
or U4683 (N_4683,In_909,In_153);
or U4684 (N_4684,In_83,In_944);
nor U4685 (N_4685,In_224,In_79);
nand U4686 (N_4686,In_209,In_943);
nor U4687 (N_4687,In_683,In_282);
and U4688 (N_4688,In_864,In_789);
and U4689 (N_4689,In_98,In_890);
nor U4690 (N_4690,In_514,In_565);
nor U4691 (N_4691,In_321,In_306);
and U4692 (N_4692,In_129,In_185);
nor U4693 (N_4693,In_745,In_908);
and U4694 (N_4694,In_104,In_184);
or U4695 (N_4695,In_556,In_168);
and U4696 (N_4696,In_450,In_495);
nor U4697 (N_4697,In_949,In_956);
nor U4698 (N_4698,In_535,In_271);
nand U4699 (N_4699,In_83,In_531);
nor U4700 (N_4700,In_232,In_924);
nor U4701 (N_4701,In_3,In_81);
nor U4702 (N_4702,In_663,In_671);
nand U4703 (N_4703,In_316,In_884);
xor U4704 (N_4704,In_423,In_792);
nand U4705 (N_4705,In_86,In_371);
xnor U4706 (N_4706,In_648,In_357);
nor U4707 (N_4707,In_454,In_419);
nand U4708 (N_4708,In_133,In_663);
or U4709 (N_4709,In_54,In_446);
nor U4710 (N_4710,In_118,In_747);
or U4711 (N_4711,In_372,In_868);
nand U4712 (N_4712,In_5,In_113);
xor U4713 (N_4713,In_732,In_527);
nor U4714 (N_4714,In_264,In_606);
and U4715 (N_4715,In_343,In_835);
and U4716 (N_4716,In_668,In_226);
nor U4717 (N_4717,In_326,In_518);
or U4718 (N_4718,In_638,In_380);
or U4719 (N_4719,In_903,In_635);
or U4720 (N_4720,In_987,In_906);
or U4721 (N_4721,In_88,In_156);
nor U4722 (N_4722,In_533,In_23);
nor U4723 (N_4723,In_916,In_983);
xor U4724 (N_4724,In_832,In_322);
xnor U4725 (N_4725,In_654,In_280);
or U4726 (N_4726,In_90,In_241);
and U4727 (N_4727,In_704,In_892);
xnor U4728 (N_4728,In_24,In_400);
nand U4729 (N_4729,In_195,In_878);
or U4730 (N_4730,In_183,In_139);
and U4731 (N_4731,In_722,In_779);
and U4732 (N_4732,In_944,In_982);
xnor U4733 (N_4733,In_314,In_367);
and U4734 (N_4734,In_532,In_599);
nor U4735 (N_4735,In_380,In_284);
and U4736 (N_4736,In_443,In_374);
nor U4737 (N_4737,In_942,In_730);
xor U4738 (N_4738,In_245,In_152);
nor U4739 (N_4739,In_621,In_926);
or U4740 (N_4740,In_890,In_229);
nor U4741 (N_4741,In_82,In_582);
and U4742 (N_4742,In_598,In_193);
nand U4743 (N_4743,In_856,In_841);
and U4744 (N_4744,In_80,In_617);
nor U4745 (N_4745,In_750,In_700);
xnor U4746 (N_4746,In_200,In_669);
xnor U4747 (N_4747,In_401,In_348);
or U4748 (N_4748,In_322,In_671);
or U4749 (N_4749,In_327,In_487);
nand U4750 (N_4750,In_569,In_515);
nand U4751 (N_4751,In_150,In_964);
xnor U4752 (N_4752,In_426,In_542);
nand U4753 (N_4753,In_405,In_546);
xnor U4754 (N_4754,In_510,In_308);
and U4755 (N_4755,In_116,In_977);
or U4756 (N_4756,In_204,In_986);
and U4757 (N_4757,In_608,In_95);
xor U4758 (N_4758,In_22,In_806);
xor U4759 (N_4759,In_368,In_640);
nand U4760 (N_4760,In_635,In_608);
and U4761 (N_4761,In_406,In_518);
nand U4762 (N_4762,In_659,In_690);
or U4763 (N_4763,In_114,In_755);
or U4764 (N_4764,In_996,In_786);
xnor U4765 (N_4765,In_930,In_274);
xnor U4766 (N_4766,In_302,In_361);
nor U4767 (N_4767,In_316,In_573);
and U4768 (N_4768,In_711,In_760);
xnor U4769 (N_4769,In_268,In_992);
or U4770 (N_4770,In_417,In_49);
nand U4771 (N_4771,In_139,In_617);
and U4772 (N_4772,In_131,In_443);
nand U4773 (N_4773,In_951,In_95);
and U4774 (N_4774,In_688,In_330);
nor U4775 (N_4775,In_623,In_685);
nor U4776 (N_4776,In_444,In_790);
and U4777 (N_4777,In_954,In_353);
xor U4778 (N_4778,In_569,In_815);
xnor U4779 (N_4779,In_499,In_733);
or U4780 (N_4780,In_538,In_134);
and U4781 (N_4781,In_435,In_767);
nor U4782 (N_4782,In_790,In_657);
and U4783 (N_4783,In_715,In_956);
or U4784 (N_4784,In_679,In_985);
xnor U4785 (N_4785,In_763,In_413);
nand U4786 (N_4786,In_616,In_229);
nand U4787 (N_4787,In_548,In_349);
or U4788 (N_4788,In_644,In_909);
xnor U4789 (N_4789,In_9,In_747);
or U4790 (N_4790,In_188,In_568);
nor U4791 (N_4791,In_415,In_54);
nand U4792 (N_4792,In_252,In_222);
xor U4793 (N_4793,In_631,In_427);
and U4794 (N_4794,In_253,In_904);
nor U4795 (N_4795,In_796,In_830);
or U4796 (N_4796,In_235,In_222);
nand U4797 (N_4797,In_708,In_9);
nand U4798 (N_4798,In_828,In_738);
and U4799 (N_4799,In_787,In_176);
nand U4800 (N_4800,In_558,In_529);
or U4801 (N_4801,In_835,In_854);
or U4802 (N_4802,In_352,In_651);
or U4803 (N_4803,In_360,In_658);
and U4804 (N_4804,In_702,In_320);
nor U4805 (N_4805,In_481,In_200);
xor U4806 (N_4806,In_269,In_60);
or U4807 (N_4807,In_888,In_537);
or U4808 (N_4808,In_666,In_138);
nand U4809 (N_4809,In_901,In_906);
xor U4810 (N_4810,In_443,In_913);
and U4811 (N_4811,In_426,In_833);
or U4812 (N_4812,In_548,In_632);
or U4813 (N_4813,In_772,In_500);
nand U4814 (N_4814,In_284,In_449);
and U4815 (N_4815,In_983,In_818);
and U4816 (N_4816,In_476,In_637);
nor U4817 (N_4817,In_541,In_503);
and U4818 (N_4818,In_752,In_287);
nand U4819 (N_4819,In_767,In_296);
or U4820 (N_4820,In_217,In_13);
nor U4821 (N_4821,In_785,In_212);
nand U4822 (N_4822,In_340,In_805);
or U4823 (N_4823,In_637,In_399);
xnor U4824 (N_4824,In_475,In_343);
or U4825 (N_4825,In_58,In_533);
nand U4826 (N_4826,In_888,In_997);
nor U4827 (N_4827,In_677,In_575);
and U4828 (N_4828,In_544,In_318);
xnor U4829 (N_4829,In_169,In_481);
or U4830 (N_4830,In_819,In_253);
nand U4831 (N_4831,In_504,In_945);
nor U4832 (N_4832,In_870,In_31);
or U4833 (N_4833,In_6,In_810);
nor U4834 (N_4834,In_60,In_671);
or U4835 (N_4835,In_972,In_813);
or U4836 (N_4836,In_298,In_192);
nand U4837 (N_4837,In_757,In_607);
and U4838 (N_4838,In_680,In_544);
or U4839 (N_4839,In_638,In_955);
or U4840 (N_4840,In_406,In_970);
nor U4841 (N_4841,In_987,In_131);
or U4842 (N_4842,In_590,In_942);
xnor U4843 (N_4843,In_594,In_336);
or U4844 (N_4844,In_574,In_920);
or U4845 (N_4845,In_349,In_541);
or U4846 (N_4846,In_509,In_306);
xor U4847 (N_4847,In_773,In_453);
nor U4848 (N_4848,In_319,In_229);
xor U4849 (N_4849,In_205,In_737);
or U4850 (N_4850,In_273,In_109);
xnor U4851 (N_4851,In_903,In_257);
and U4852 (N_4852,In_812,In_356);
or U4853 (N_4853,In_287,In_834);
nor U4854 (N_4854,In_969,In_871);
nand U4855 (N_4855,In_709,In_786);
or U4856 (N_4856,In_803,In_270);
xnor U4857 (N_4857,In_880,In_109);
and U4858 (N_4858,In_638,In_186);
xor U4859 (N_4859,In_322,In_82);
or U4860 (N_4860,In_842,In_0);
or U4861 (N_4861,In_649,In_816);
or U4862 (N_4862,In_918,In_920);
xor U4863 (N_4863,In_888,In_36);
xor U4864 (N_4864,In_564,In_72);
or U4865 (N_4865,In_557,In_448);
or U4866 (N_4866,In_52,In_202);
nor U4867 (N_4867,In_23,In_315);
nand U4868 (N_4868,In_40,In_451);
xor U4869 (N_4869,In_640,In_656);
or U4870 (N_4870,In_423,In_670);
and U4871 (N_4871,In_303,In_521);
and U4872 (N_4872,In_439,In_431);
nor U4873 (N_4873,In_524,In_621);
or U4874 (N_4874,In_570,In_956);
nor U4875 (N_4875,In_562,In_890);
and U4876 (N_4876,In_895,In_299);
xnor U4877 (N_4877,In_719,In_150);
nand U4878 (N_4878,In_178,In_928);
xnor U4879 (N_4879,In_387,In_63);
xor U4880 (N_4880,In_435,In_618);
xnor U4881 (N_4881,In_315,In_539);
or U4882 (N_4882,In_711,In_307);
xnor U4883 (N_4883,In_379,In_54);
xor U4884 (N_4884,In_860,In_938);
xor U4885 (N_4885,In_608,In_5);
xnor U4886 (N_4886,In_582,In_487);
xor U4887 (N_4887,In_683,In_949);
xnor U4888 (N_4888,In_4,In_413);
nand U4889 (N_4889,In_320,In_445);
nor U4890 (N_4890,In_339,In_282);
and U4891 (N_4891,In_41,In_230);
or U4892 (N_4892,In_2,In_179);
xnor U4893 (N_4893,In_968,In_650);
nor U4894 (N_4894,In_783,In_216);
or U4895 (N_4895,In_864,In_509);
nand U4896 (N_4896,In_102,In_134);
xnor U4897 (N_4897,In_353,In_547);
nand U4898 (N_4898,In_992,In_114);
nor U4899 (N_4899,In_181,In_34);
xnor U4900 (N_4900,In_608,In_285);
or U4901 (N_4901,In_502,In_884);
nor U4902 (N_4902,In_142,In_416);
xnor U4903 (N_4903,In_565,In_423);
nand U4904 (N_4904,In_959,In_538);
xnor U4905 (N_4905,In_973,In_710);
nor U4906 (N_4906,In_19,In_12);
nand U4907 (N_4907,In_709,In_239);
nor U4908 (N_4908,In_9,In_452);
nand U4909 (N_4909,In_939,In_744);
nor U4910 (N_4910,In_27,In_197);
xnor U4911 (N_4911,In_538,In_396);
nand U4912 (N_4912,In_796,In_802);
or U4913 (N_4913,In_98,In_648);
nor U4914 (N_4914,In_491,In_96);
nor U4915 (N_4915,In_839,In_769);
and U4916 (N_4916,In_659,In_175);
and U4917 (N_4917,In_739,In_412);
nor U4918 (N_4918,In_583,In_700);
and U4919 (N_4919,In_287,In_381);
and U4920 (N_4920,In_872,In_738);
nand U4921 (N_4921,In_676,In_922);
or U4922 (N_4922,In_846,In_403);
or U4923 (N_4923,In_869,In_940);
or U4924 (N_4924,In_856,In_346);
or U4925 (N_4925,In_896,In_495);
and U4926 (N_4926,In_404,In_605);
nor U4927 (N_4927,In_283,In_620);
nor U4928 (N_4928,In_663,In_586);
nand U4929 (N_4929,In_997,In_914);
or U4930 (N_4930,In_157,In_929);
nand U4931 (N_4931,In_410,In_168);
or U4932 (N_4932,In_438,In_479);
and U4933 (N_4933,In_274,In_819);
nand U4934 (N_4934,In_551,In_167);
or U4935 (N_4935,In_372,In_239);
nand U4936 (N_4936,In_223,In_288);
or U4937 (N_4937,In_469,In_283);
nor U4938 (N_4938,In_819,In_994);
and U4939 (N_4939,In_877,In_530);
or U4940 (N_4940,In_441,In_317);
and U4941 (N_4941,In_373,In_960);
nor U4942 (N_4942,In_306,In_412);
or U4943 (N_4943,In_650,In_614);
and U4944 (N_4944,In_872,In_44);
xor U4945 (N_4945,In_637,In_302);
or U4946 (N_4946,In_918,In_88);
and U4947 (N_4947,In_436,In_773);
nor U4948 (N_4948,In_140,In_343);
nor U4949 (N_4949,In_149,In_948);
or U4950 (N_4950,In_646,In_702);
and U4951 (N_4951,In_758,In_849);
nor U4952 (N_4952,In_519,In_107);
xor U4953 (N_4953,In_495,In_257);
xor U4954 (N_4954,In_869,In_807);
and U4955 (N_4955,In_447,In_981);
or U4956 (N_4956,In_176,In_258);
nand U4957 (N_4957,In_248,In_567);
or U4958 (N_4958,In_7,In_403);
nor U4959 (N_4959,In_492,In_144);
and U4960 (N_4960,In_292,In_412);
and U4961 (N_4961,In_130,In_423);
or U4962 (N_4962,In_703,In_217);
nor U4963 (N_4963,In_455,In_536);
and U4964 (N_4964,In_264,In_236);
and U4965 (N_4965,In_364,In_994);
or U4966 (N_4966,In_241,In_920);
nor U4967 (N_4967,In_280,In_105);
xor U4968 (N_4968,In_263,In_757);
nor U4969 (N_4969,In_7,In_996);
xnor U4970 (N_4970,In_118,In_946);
and U4971 (N_4971,In_70,In_957);
xor U4972 (N_4972,In_772,In_767);
or U4973 (N_4973,In_468,In_209);
nor U4974 (N_4974,In_158,In_485);
nand U4975 (N_4975,In_867,In_85);
and U4976 (N_4976,In_616,In_524);
or U4977 (N_4977,In_157,In_212);
or U4978 (N_4978,In_238,In_795);
and U4979 (N_4979,In_286,In_52);
nand U4980 (N_4980,In_301,In_829);
nand U4981 (N_4981,In_978,In_987);
xnor U4982 (N_4982,In_696,In_42);
nor U4983 (N_4983,In_13,In_401);
nor U4984 (N_4984,In_897,In_765);
xor U4985 (N_4985,In_927,In_970);
nand U4986 (N_4986,In_528,In_232);
nand U4987 (N_4987,In_539,In_753);
xnor U4988 (N_4988,In_880,In_565);
nor U4989 (N_4989,In_133,In_55);
or U4990 (N_4990,In_875,In_794);
xor U4991 (N_4991,In_137,In_401);
and U4992 (N_4992,In_95,In_630);
xnor U4993 (N_4993,In_447,In_801);
and U4994 (N_4994,In_439,In_36);
or U4995 (N_4995,In_685,In_478);
or U4996 (N_4996,In_627,In_480);
xnor U4997 (N_4997,In_194,In_803);
and U4998 (N_4998,In_752,In_55);
nor U4999 (N_4999,In_583,In_705);
and U5000 (N_5000,N_755,N_2905);
and U5001 (N_5001,N_100,N_368);
xor U5002 (N_5002,N_4205,N_2033);
or U5003 (N_5003,N_4141,N_328);
xnor U5004 (N_5004,N_474,N_810);
and U5005 (N_5005,N_4779,N_2133);
nor U5006 (N_5006,N_1230,N_511);
or U5007 (N_5007,N_3151,N_4295);
nand U5008 (N_5008,N_994,N_4886);
nor U5009 (N_5009,N_1808,N_2249);
and U5010 (N_5010,N_3641,N_1803);
or U5011 (N_5011,N_2195,N_2982);
and U5012 (N_5012,N_2794,N_1760);
and U5013 (N_5013,N_2956,N_2731);
and U5014 (N_5014,N_4327,N_4876);
nand U5015 (N_5015,N_3174,N_4284);
and U5016 (N_5016,N_4861,N_3224);
xor U5017 (N_5017,N_145,N_3901);
nor U5018 (N_5018,N_4572,N_3361);
or U5019 (N_5019,N_415,N_298);
nor U5020 (N_5020,N_898,N_1470);
xnor U5021 (N_5021,N_3044,N_3021);
xor U5022 (N_5022,N_1981,N_1231);
nand U5023 (N_5023,N_3980,N_549);
or U5024 (N_5024,N_334,N_466);
nor U5025 (N_5025,N_3928,N_4985);
nand U5026 (N_5026,N_969,N_4880);
and U5027 (N_5027,N_1621,N_2899);
nor U5028 (N_5028,N_4470,N_3691);
or U5029 (N_5029,N_750,N_1194);
or U5030 (N_5030,N_2366,N_1991);
nor U5031 (N_5031,N_3406,N_3240);
or U5032 (N_5032,N_1419,N_3636);
nor U5033 (N_5033,N_3043,N_3790);
and U5034 (N_5034,N_1137,N_3781);
and U5035 (N_5035,N_4850,N_805);
nand U5036 (N_5036,N_2386,N_1340);
nor U5037 (N_5037,N_4366,N_276);
and U5038 (N_5038,N_3315,N_4591);
xor U5039 (N_5039,N_1712,N_4391);
nor U5040 (N_5040,N_4988,N_3339);
nand U5041 (N_5041,N_2745,N_4469);
nor U5042 (N_5042,N_2970,N_200);
nor U5043 (N_5043,N_385,N_4481);
and U5044 (N_5044,N_1906,N_3030);
or U5045 (N_5045,N_691,N_1829);
or U5046 (N_5046,N_586,N_1001);
or U5047 (N_5047,N_1792,N_3565);
nor U5048 (N_5048,N_2364,N_782);
xor U5049 (N_5049,N_624,N_1176);
or U5050 (N_5050,N_4101,N_4598);
xnor U5051 (N_5051,N_2517,N_1774);
nand U5052 (N_5052,N_768,N_1051);
nor U5053 (N_5053,N_4786,N_2499);
nor U5054 (N_5054,N_4055,N_1607);
nor U5055 (N_5055,N_275,N_272);
and U5056 (N_5056,N_3326,N_233);
nand U5057 (N_5057,N_4232,N_1322);
nor U5058 (N_5058,N_889,N_4049);
and U5059 (N_5059,N_1400,N_3727);
and U5060 (N_5060,N_4342,N_1102);
nor U5061 (N_5061,N_2670,N_3945);
and U5062 (N_5062,N_1057,N_3515);
nor U5063 (N_5063,N_1560,N_2363);
or U5064 (N_5064,N_2415,N_217);
and U5065 (N_5065,N_3772,N_4667);
nor U5066 (N_5066,N_273,N_2354);
and U5067 (N_5067,N_4912,N_2062);
nand U5068 (N_5068,N_3733,N_2466);
or U5069 (N_5069,N_3723,N_1933);
nand U5070 (N_5070,N_4977,N_2128);
nand U5071 (N_5071,N_2305,N_4854);
xor U5072 (N_5072,N_1853,N_2320);
or U5073 (N_5073,N_1645,N_1476);
and U5074 (N_5074,N_4245,N_581);
xor U5075 (N_5075,N_2586,N_235);
or U5076 (N_5076,N_899,N_201);
nor U5077 (N_5077,N_2471,N_1148);
or U5078 (N_5078,N_3197,N_1518);
nand U5079 (N_5079,N_2625,N_4766);
nand U5080 (N_5080,N_540,N_3485);
nor U5081 (N_5081,N_1611,N_353);
nand U5082 (N_5082,N_464,N_1542);
or U5083 (N_5083,N_3989,N_3101);
xor U5084 (N_5084,N_3711,N_1074);
and U5085 (N_5085,N_3512,N_1003);
or U5086 (N_5086,N_1869,N_319);
and U5087 (N_5087,N_1827,N_1602);
nor U5088 (N_5088,N_2056,N_73);
and U5089 (N_5089,N_2820,N_461);
nand U5090 (N_5090,N_1559,N_4337);
and U5091 (N_5091,N_2132,N_4976);
and U5092 (N_5092,N_4445,N_3715);
and U5093 (N_5093,N_672,N_527);
nor U5094 (N_5094,N_4581,N_1885);
nand U5095 (N_5095,N_1583,N_3075);
or U5096 (N_5096,N_408,N_3333);
nand U5097 (N_5097,N_4701,N_4484);
nor U5098 (N_5098,N_611,N_584);
and U5099 (N_5099,N_4459,N_4440);
or U5100 (N_5100,N_1737,N_4962);
nor U5101 (N_5101,N_4460,N_1601);
nand U5102 (N_5102,N_1442,N_971);
nand U5103 (N_5103,N_3698,N_836);
nor U5104 (N_5104,N_943,N_4240);
nor U5105 (N_5105,N_620,N_2325);
or U5106 (N_5106,N_490,N_1545);
xor U5107 (N_5107,N_4318,N_1263);
nand U5108 (N_5108,N_2252,N_1311);
or U5109 (N_5109,N_1278,N_3903);
xnor U5110 (N_5110,N_325,N_3201);
and U5111 (N_5111,N_1140,N_91);
and U5112 (N_5112,N_829,N_1091);
xor U5113 (N_5113,N_3494,N_4326);
nand U5114 (N_5114,N_4673,N_659);
and U5115 (N_5115,N_2263,N_4899);
nand U5116 (N_5116,N_1673,N_2702);
xor U5117 (N_5117,N_913,N_1095);
or U5118 (N_5118,N_118,N_4213);
and U5119 (N_5119,N_1153,N_996);
nand U5120 (N_5120,N_3425,N_2894);
and U5121 (N_5121,N_4688,N_4528);
and U5122 (N_5122,N_4200,N_4718);
xnor U5123 (N_5123,N_3161,N_3492);
and U5124 (N_5124,N_3705,N_4379);
xor U5125 (N_5125,N_2661,N_3517);
nor U5126 (N_5126,N_1546,N_2689);
or U5127 (N_5127,N_1550,N_1082);
or U5128 (N_5128,N_4785,N_974);
and U5129 (N_5129,N_1493,N_4751);
and U5130 (N_5130,N_2273,N_3622);
and U5131 (N_5131,N_2506,N_4154);
nor U5132 (N_5132,N_2999,N_4601);
xnor U5133 (N_5133,N_2412,N_3583);
or U5134 (N_5134,N_3371,N_3440);
nand U5135 (N_5135,N_4378,N_4171);
nand U5136 (N_5136,N_3412,N_2888);
nand U5137 (N_5137,N_1844,N_401);
or U5138 (N_5138,N_3884,N_1783);
xor U5139 (N_5139,N_955,N_3629);
nand U5140 (N_5140,N_378,N_2308);
or U5141 (N_5141,N_525,N_1762);
or U5142 (N_5142,N_4864,N_695);
xnor U5143 (N_5143,N_841,N_3567);
and U5144 (N_5144,N_1732,N_4216);
and U5145 (N_5145,N_3159,N_3531);
nand U5146 (N_5146,N_1608,N_2573);
nand U5147 (N_5147,N_4927,N_569);
xnor U5148 (N_5148,N_1328,N_4402);
xor U5149 (N_5149,N_242,N_1454);
nand U5150 (N_5150,N_638,N_3788);
or U5151 (N_5151,N_3031,N_3195);
or U5152 (N_5152,N_3179,N_1466);
or U5153 (N_5153,N_4239,N_3287);
xor U5154 (N_5154,N_45,N_2685);
nor U5155 (N_5155,N_1767,N_4717);
nand U5156 (N_5156,N_4056,N_4332);
nor U5157 (N_5157,N_4994,N_3115);
or U5158 (N_5158,N_4400,N_3346);
nor U5159 (N_5159,N_891,N_3049);
or U5160 (N_5160,N_119,N_3285);
and U5161 (N_5161,N_326,N_293);
nor U5162 (N_5162,N_3038,N_789);
or U5163 (N_5163,N_2954,N_3245);
nand U5164 (N_5164,N_3569,N_2251);
nand U5165 (N_5165,N_3740,N_2553);
xor U5166 (N_5166,N_1930,N_2748);
xnor U5167 (N_5167,N_4291,N_2516);
xor U5168 (N_5168,N_95,N_510);
nor U5169 (N_5169,N_1994,N_3035);
nand U5170 (N_5170,N_1689,N_2280);
nor U5171 (N_5171,N_397,N_3267);
and U5172 (N_5172,N_3480,N_3123);
nor U5173 (N_5173,N_909,N_1505);
nor U5174 (N_5174,N_3695,N_2452);
nand U5175 (N_5175,N_2546,N_4077);
nor U5176 (N_5176,N_3748,N_4600);
xor U5177 (N_5177,N_3602,N_2779);
nor U5178 (N_5178,N_2226,N_802);
xnor U5179 (N_5179,N_109,N_770);
nand U5180 (N_5180,N_3717,N_1150);
nand U5181 (N_5181,N_808,N_4594);
or U5182 (N_5182,N_4421,N_130);
or U5183 (N_5183,N_998,N_877);
nor U5184 (N_5184,N_1374,N_2981);
or U5185 (N_5185,N_1554,N_4110);
nor U5186 (N_5186,N_467,N_3437);
nand U5187 (N_5187,N_1226,N_2081);
and U5188 (N_5188,N_1432,N_2436);
nand U5189 (N_5189,N_3911,N_3783);
nor U5190 (N_5190,N_820,N_1144);
and U5191 (N_5191,N_3904,N_2846);
nand U5192 (N_5192,N_373,N_4944);
and U5193 (N_5193,N_4658,N_1857);
and U5194 (N_5194,N_4403,N_2526);
xnor U5195 (N_5195,N_872,N_3754);
nor U5196 (N_5196,N_3228,N_3550);
and U5197 (N_5197,N_1478,N_1572);
nor U5198 (N_5198,N_2148,N_4040);
nor U5199 (N_5199,N_2938,N_930);
nor U5200 (N_5200,N_486,N_1066);
nand U5201 (N_5201,N_1490,N_1507);
nand U5202 (N_5202,N_3447,N_925);
and U5203 (N_5203,N_556,N_1142);
nor U5204 (N_5204,N_1175,N_3807);
and U5205 (N_5205,N_4159,N_3538);
xnor U5206 (N_5206,N_3999,N_1145);
and U5207 (N_5207,N_2446,N_3786);
or U5208 (N_5208,N_796,N_2800);
or U5209 (N_5209,N_975,N_1119);
nand U5210 (N_5210,N_4569,N_4943);
xor U5211 (N_5211,N_3072,N_2222);
xnor U5212 (N_5212,N_2806,N_3493);
or U5213 (N_5213,N_2311,N_4259);
nand U5214 (N_5214,N_2127,N_662);
or U5215 (N_5215,N_1480,N_658);
nand U5216 (N_5216,N_3796,N_357);
nand U5217 (N_5217,N_205,N_688);
xnor U5218 (N_5218,N_3861,N_2609);
nand U5219 (N_5219,N_1812,N_4522);
nor U5220 (N_5220,N_1786,N_2299);
or U5221 (N_5221,N_4914,N_2350);
nor U5222 (N_5222,N_1818,N_628);
and U5223 (N_5223,N_124,N_2074);
nand U5224 (N_5224,N_3433,N_4755);
and U5225 (N_5225,N_626,N_4565);
xnor U5226 (N_5226,N_1959,N_3968);
or U5227 (N_5227,N_4230,N_20);
or U5228 (N_5228,N_4848,N_1884);
xnor U5229 (N_5229,N_386,N_2260);
nor U5230 (N_5230,N_4094,N_451);
xor U5231 (N_5231,N_702,N_3458);
nor U5232 (N_5232,N_355,N_1438);
or U5233 (N_5233,N_166,N_2259);
xor U5234 (N_5234,N_533,N_1726);
xnor U5235 (N_5235,N_1811,N_4472);
xnor U5236 (N_5236,N_4080,N_2037);
or U5237 (N_5237,N_1355,N_4517);
xnor U5238 (N_5238,N_4903,N_1071);
and U5239 (N_5239,N_2986,N_4852);
xnor U5240 (N_5240,N_2706,N_2833);
nor U5241 (N_5241,N_2399,N_4115);
nor U5242 (N_5242,N_3002,N_1060);
xor U5243 (N_5243,N_1464,N_2844);
nand U5244 (N_5244,N_3478,N_1138);
xnor U5245 (N_5245,N_3652,N_2442);
nand U5246 (N_5246,N_3080,N_4248);
nor U5247 (N_5247,N_4193,N_2435);
xnor U5248 (N_5248,N_4748,N_3252);
xnor U5249 (N_5249,N_19,N_1562);
nor U5250 (N_5250,N_4277,N_4794);
nor U5251 (N_5251,N_4693,N_230);
xor U5252 (N_5252,N_1850,N_547);
nand U5253 (N_5253,N_2911,N_2796);
nand U5254 (N_5254,N_3832,N_2505);
or U5255 (N_5255,N_4137,N_4253);
and U5256 (N_5256,N_4729,N_4426);
and U5257 (N_5257,N_2021,N_2687);
and U5258 (N_5258,N_1566,N_3686);
xnor U5259 (N_5259,N_3153,N_4335);
nor U5260 (N_5260,N_3133,N_1791);
and U5261 (N_5261,N_2790,N_4406);
or U5262 (N_5262,N_3771,N_1483);
nor U5263 (N_5263,N_274,N_827);
xnor U5264 (N_5264,N_2218,N_2443);
nand U5265 (N_5265,N_1233,N_3286);
nand U5266 (N_5266,N_512,N_3657);
nor U5267 (N_5267,N_3768,N_2409);
xnor U5268 (N_5268,N_3836,N_4288);
nor U5269 (N_5269,N_202,N_4561);
nor U5270 (N_5270,N_632,N_3124);
and U5271 (N_5271,N_3455,N_2361);
nand U5272 (N_5272,N_2686,N_2980);
or U5273 (N_5273,N_1370,N_4995);
or U5274 (N_5274,N_3548,N_886);
xor U5275 (N_5275,N_2893,N_3918);
and U5276 (N_5276,N_689,N_3353);
nor U5277 (N_5277,N_423,N_459);
xor U5278 (N_5278,N_4499,N_4936);
or U5279 (N_5279,N_460,N_3831);
and U5280 (N_5280,N_1512,N_3546);
xor U5281 (N_5281,N_2859,N_3857);
and U5282 (N_5282,N_1882,N_1899);
or U5283 (N_5283,N_830,N_3022);
or U5284 (N_5284,N_3572,N_3415);
or U5285 (N_5285,N_383,N_1042);
or U5286 (N_5286,N_4461,N_522);
or U5287 (N_5287,N_1484,N_2777);
and U5288 (N_5288,N_1963,N_4182);
xor U5289 (N_5289,N_3894,N_1260);
or U5290 (N_5290,N_1841,N_4832);
or U5291 (N_5291,N_3155,N_2935);
nor U5292 (N_5292,N_1964,N_2303);
xnor U5293 (N_5293,N_4915,N_1492);
or U5294 (N_5294,N_4802,N_193);
nor U5295 (N_5295,N_4412,N_4136);
or U5296 (N_5296,N_4628,N_582);
nand U5297 (N_5297,N_2632,N_4466);
and U5298 (N_5298,N_3676,N_2229);
and U5299 (N_5299,N_1851,N_2297);
nand U5300 (N_5300,N_3725,N_4651);
or U5301 (N_5301,N_2194,N_1946);
xor U5302 (N_5302,N_1942,N_2246);
xnor U5303 (N_5303,N_311,N_2000);
xnor U5304 (N_5304,N_669,N_1659);
nand U5305 (N_5305,N_4933,N_2590);
nand U5306 (N_5306,N_678,N_1460);
nand U5307 (N_5307,N_3793,N_1469);
and U5308 (N_5308,N_2003,N_3509);
nand U5309 (N_5309,N_3812,N_4971);
xor U5310 (N_5310,N_1907,N_3242);
or U5311 (N_5311,N_1598,N_2667);
nand U5312 (N_5312,N_2549,N_1614);
nand U5313 (N_5313,N_912,N_4145);
nand U5314 (N_5314,N_1660,N_2727);
or U5315 (N_5315,N_2795,N_879);
or U5316 (N_5316,N_36,N_3764);
and U5317 (N_5317,N_639,N_1761);
nor U5318 (N_5318,N_3281,N_4817);
nand U5319 (N_5319,N_3874,N_18);
or U5320 (N_5320,N_32,N_3063);
and U5321 (N_5321,N_552,N_416);
xor U5322 (N_5322,N_788,N_4105);
nor U5323 (N_5323,N_4874,N_1005);
nand U5324 (N_5324,N_1014,N_3845);
xor U5325 (N_5325,N_3370,N_3470);
xnor U5326 (N_5326,N_2428,N_356);
and U5327 (N_5327,N_3656,N_4507);
xor U5328 (N_5328,N_3940,N_381);
nor U5329 (N_5329,N_2184,N_3580);
or U5330 (N_5330,N_4293,N_3510);
xor U5331 (N_5331,N_2508,N_4855);
nand U5332 (N_5332,N_4262,N_1427);
and U5333 (N_5333,N_3443,N_455);
xor U5334 (N_5334,N_2697,N_697);
and U5335 (N_5335,N_4131,N_4908);
or U5336 (N_5336,N_2847,N_1364);
nor U5337 (N_5337,N_2459,N_1232);
or U5338 (N_5338,N_745,N_647);
nor U5339 (N_5339,N_939,N_758);
or U5340 (N_5340,N_4317,N_675);
xor U5341 (N_5341,N_3731,N_3843);
or U5342 (N_5342,N_67,N_3489);
or U5343 (N_5343,N_3034,N_2574);
and U5344 (N_5344,N_4282,N_4109);
and U5345 (N_5345,N_2425,N_1842);
nor U5346 (N_5346,N_4893,N_1475);
xnor U5347 (N_5347,N_2611,N_4334);
nand U5348 (N_5348,N_2943,N_404);
and U5349 (N_5349,N_3936,N_1411);
xnor U5350 (N_5350,N_2090,N_3895);
or U5351 (N_5351,N_1993,N_410);
nor U5352 (N_5352,N_4663,N_2877);
nand U5353 (N_5353,N_778,N_3524);
and U5354 (N_5354,N_2395,N_4249);
nor U5355 (N_5355,N_3840,N_852);
nand U5356 (N_5356,N_2371,N_2649);
nor U5357 (N_5357,N_1152,N_3611);
xor U5358 (N_5358,N_809,N_1831);
nor U5359 (N_5359,N_414,N_82);
xnor U5360 (N_5360,N_2873,N_3551);
and U5361 (N_5361,N_893,N_4341);
xor U5362 (N_5362,N_4800,N_2657);
nor U5363 (N_5363,N_4415,N_2676);
and U5364 (N_5364,N_4924,N_1391);
or U5365 (N_5365,N_3718,N_3738);
and U5366 (N_5366,N_3759,N_2340);
xnor U5367 (N_5367,N_2151,N_643);
nor U5368 (N_5368,N_3187,N_736);
nand U5369 (N_5369,N_4895,N_3853);
nand U5370 (N_5370,N_158,N_567);
nand U5371 (N_5371,N_2124,N_2129);
nor U5372 (N_5372,N_1903,N_2942);
nand U5373 (N_5373,N_294,N_849);
nor U5374 (N_5374,N_4273,N_2560);
or U5375 (N_5375,N_1229,N_2176);
or U5376 (N_5376,N_2801,N_1861);
nor U5377 (N_5377,N_4227,N_1863);
nor U5378 (N_5378,N_3780,N_2708);
or U5379 (N_5379,N_3017,N_3053);
nor U5380 (N_5380,N_3357,N_3402);
xnor U5381 (N_5381,N_2357,N_4827);
nor U5382 (N_5382,N_1250,N_1336);
xnor U5383 (N_5383,N_1543,N_1805);
nor U5384 (N_5384,N_989,N_2304);
xnor U5385 (N_5385,N_926,N_4928);
nor U5386 (N_5386,N_421,N_114);
xnor U5387 (N_5387,N_3445,N_3844);
or U5388 (N_5388,N_3774,N_4602);
nor U5389 (N_5389,N_536,N_4791);
and U5390 (N_5390,N_2921,N_1021);
xnor U5391 (N_5391,N_767,N_1718);
nand U5392 (N_5392,N_3975,N_3972);
and U5393 (N_5393,N_3007,N_4694);
or U5394 (N_5394,N_3331,N_2211);
and U5395 (N_5395,N_4149,N_2726);
and U5396 (N_5396,N_4552,N_2694);
xor U5397 (N_5397,N_1113,N_2022);
nand U5398 (N_5398,N_693,N_1700);
nand U5399 (N_5399,N_2589,N_187);
and U5400 (N_5400,N_1276,N_2855);
nor U5401 (N_5401,N_722,N_3024);
and U5402 (N_5402,N_3981,N_2396);
nor U5403 (N_5403,N_3970,N_1187);
or U5404 (N_5404,N_3677,N_1481);
and U5405 (N_5405,N_4423,N_1154);
nor U5406 (N_5406,N_1925,N_3720);
and U5407 (N_5407,N_4735,N_4554);
xnor U5408 (N_5408,N_881,N_3878);
xor U5409 (N_5409,N_1671,N_760);
or U5410 (N_5410,N_3506,N_3332);
nand U5411 (N_5411,N_2843,N_3355);
xnor U5412 (N_5412,N_4405,N_443);
nand U5413 (N_5413,N_3454,N_358);
nor U5414 (N_5414,N_3871,N_1526);
nor U5415 (N_5415,N_1000,N_2046);
and U5416 (N_5416,N_2643,N_4532);
or U5417 (N_5417,N_4442,N_701);
nor U5418 (N_5418,N_2821,N_3107);
xnor U5419 (N_5419,N_794,N_2239);
or U5420 (N_5420,N_2461,N_308);
xor U5421 (N_5421,N_1445,N_2881);
xor U5422 (N_5422,N_2701,N_4413);
xnor U5423 (N_5423,N_3309,N_409);
and U5424 (N_5424,N_4087,N_1637);
nand U5425 (N_5425,N_4384,N_417);
nor U5426 (N_5426,N_4313,N_4330);
nand U5427 (N_5427,N_1688,N_515);
nand U5428 (N_5428,N_4257,N_3303);
xor U5429 (N_5429,N_761,N_2617);
and U5430 (N_5430,N_2417,N_2974);
xnor U5431 (N_5431,N_1300,N_4290);
and U5432 (N_5432,N_1032,N_168);
nand U5433 (N_5433,N_2952,N_4617);
nor U5434 (N_5434,N_4652,N_4531);
and U5435 (N_5435,N_2167,N_182);
nor U5436 (N_5436,N_1305,N_1349);
nand U5437 (N_5437,N_305,N_1749);
xnor U5438 (N_5438,N_3291,N_216);
nand U5439 (N_5439,N_3690,N_3993);
nor U5440 (N_5440,N_729,N_3672);
nor U5441 (N_5441,N_2052,N_2217);
nand U5442 (N_5442,N_2141,N_2460);
nor U5443 (N_5443,N_4134,N_4215);
or U5444 (N_5444,N_1415,N_6);
nand U5445 (N_5445,N_985,N_4887);
and U5446 (N_5446,N_1630,N_3585);
and U5447 (N_5447,N_3459,N_2163);
or U5448 (N_5448,N_98,N_4163);
nand U5449 (N_5449,N_4206,N_3753);
or U5450 (N_5450,N_3841,N_713);
nor U5451 (N_5451,N_3553,N_3888);
xor U5452 (N_5452,N_4382,N_1618);
or U5453 (N_5453,N_2121,N_376);
or U5454 (N_5454,N_553,N_3964);
xor U5455 (N_5455,N_610,N_2889);
nor U5456 (N_5456,N_159,N_1301);
nor U5457 (N_5457,N_1223,N_1500);
nand U5458 (N_5458,N_751,N_359);
or U5459 (N_5459,N_765,N_4002);
xor U5460 (N_5460,N_4185,N_4130);
and U5461 (N_5461,N_3941,N_1662);
nand U5462 (N_5462,N_3104,N_1318);
nor U5463 (N_5463,N_2413,N_1306);
nand U5464 (N_5464,N_1107,N_2822);
or U5465 (N_5465,N_3092,N_577);
nor U5466 (N_5466,N_3609,N_997);
or U5467 (N_5467,N_742,N_3801);
nor U5468 (N_5468,N_1800,N_1339);
nand U5469 (N_5469,N_3687,N_3891);
or U5470 (N_5470,N_1025,N_1372);
or U5471 (N_5471,N_3463,N_4024);
and U5472 (N_5472,N_3164,N_1677);
and U5473 (N_5473,N_1321,N_3037);
nand U5474 (N_5474,N_2112,N_1976);
and U5475 (N_5475,N_4029,N_2870);
nand U5476 (N_5476,N_249,N_1781);
or U5477 (N_5477,N_1213,N_4011);
nand U5478 (N_5478,N_3108,N_94);
xnor U5479 (N_5479,N_208,N_3141);
xnor U5480 (N_5480,N_1736,N_3144);
or U5481 (N_5481,N_222,N_2307);
nand U5482 (N_5482,N_4860,N_4099);
nor U5483 (N_5483,N_3887,N_3077);
nand U5484 (N_5484,N_3876,N_650);
xnor U5485 (N_5485,N_1271,N_4901);
nand U5486 (N_5486,N_151,N_2012);
or U5487 (N_5487,N_2674,N_35);
nor U5488 (N_5488,N_2856,N_1817);
nor U5489 (N_5489,N_2780,N_3089);
and U5490 (N_5490,N_3689,N_4979);
and U5491 (N_5491,N_4097,N_2178);
xor U5492 (N_5492,N_3213,N_4709);
xnor U5493 (N_5493,N_4167,N_921);
xor U5494 (N_5494,N_2627,N_1126);
or U5495 (N_5495,N_3003,N_2886);
and U5496 (N_5496,N_2498,N_4926);
xor U5497 (N_5497,N_2671,N_4890);
xor U5498 (N_5498,N_4749,N_4180);
xor U5499 (N_5499,N_3631,N_2600);
and U5500 (N_5500,N_1384,N_1825);
xor U5501 (N_5501,N_2282,N_4542);
or U5502 (N_5502,N_4082,N_1290);
and U5503 (N_5503,N_1734,N_4734);
xor U5504 (N_5504,N_725,N_2375);
or U5505 (N_5505,N_377,N_1446);
and U5506 (N_5506,N_3314,N_3797);
xor U5507 (N_5507,N_739,N_2512);
nor U5508 (N_5508,N_1072,N_142);
or U5509 (N_5509,N_607,N_3671);
nand U5510 (N_5510,N_433,N_3653);
and U5511 (N_5511,N_198,N_919);
and U5512 (N_5512,N_573,N_1722);
nand U5513 (N_5513,N_3387,N_2169);
xnor U5514 (N_5514,N_4446,N_2143);
nand U5515 (N_5515,N_445,N_2931);
or U5516 (N_5516,N_630,N_3637);
and U5517 (N_5517,N_2370,N_4435);
xnor U5518 (N_5518,N_1685,N_2620);
xnor U5519 (N_5519,N_860,N_4774);
nor U5520 (N_5520,N_772,N_825);
nand U5521 (N_5521,N_3015,N_2593);
or U5522 (N_5522,N_2243,N_1004);
and U5523 (N_5523,N_4408,N_3360);
nand U5524 (N_5524,N_1646,N_2079);
nand U5525 (N_5525,N_1888,N_2971);
nor U5526 (N_5526,N_2991,N_4836);
nand U5527 (N_5527,N_3419,N_3352);
xor U5528 (N_5528,N_1958,N_4972);
nand U5529 (N_5529,N_4820,N_1010);
nor U5530 (N_5530,N_4967,N_3369);
nor U5531 (N_5531,N_3721,N_4111);
nand U5532 (N_5532,N_4819,N_26);
or U5533 (N_5533,N_4642,N_199);
nor U5534 (N_5534,N_640,N_4235);
nand U5535 (N_5535,N_2637,N_2563);
xor U5536 (N_5536,N_3040,N_2737);
nor U5537 (N_5537,N_3914,N_3958);
or U5538 (N_5538,N_933,N_4883);
xor U5539 (N_5539,N_1296,N_1116);
nand U5540 (N_5540,N_795,N_2783);
and U5541 (N_5541,N_4923,N_266);
nand U5542 (N_5542,N_1801,N_4328);
xnor U5543 (N_5543,N_1746,N_1105);
xor U5544 (N_5544,N_4496,N_2122);
nand U5545 (N_5545,N_4917,N_161);
or U5546 (N_5546,N_37,N_1508);
and U5547 (N_5547,N_288,N_4942);
xnor U5548 (N_5548,N_4455,N_1338);
xnor U5549 (N_5549,N_3603,N_4147);
nand U5550 (N_5550,N_2897,N_674);
xnor U5551 (N_5551,N_4653,N_3800);
or U5552 (N_5552,N_1380,N_1016);
xor U5553 (N_5553,N_1742,N_901);
or U5554 (N_5554,N_2717,N_2746);
xor U5555 (N_5555,N_2232,N_503);
and U5556 (N_5556,N_4038,N_4989);
or U5557 (N_5557,N_313,N_1960);
nor U5558 (N_5558,N_2103,N_904);
and U5559 (N_5559,N_2300,N_2724);
nor U5560 (N_5560,N_1333,N_4054);
or U5561 (N_5561,N_3465,N_3500);
and U5562 (N_5562,N_4960,N_4173);
or U5563 (N_5563,N_2319,N_1987);
nand U5564 (N_5564,N_3694,N_3496);
nand U5565 (N_5565,N_147,N_2057);
or U5566 (N_5566,N_1120,N_4813);
nand U5567 (N_5567,N_4298,N_4872);
nand U5568 (N_5568,N_1855,N_4025);
nand U5569 (N_5569,N_2402,N_2048);
or U5570 (N_5570,N_47,N_2392);
and U5571 (N_5571,N_3280,N_1193);
and U5572 (N_5572,N_3349,N_3409);
nand U5573 (N_5573,N_4372,N_3587);
or U5574 (N_5574,N_595,N_660);
and U5575 (N_5575,N_4896,N_1373);
and U5576 (N_5576,N_603,N_1310);
and U5577 (N_5577,N_1622,N_4708);
nor U5578 (N_5578,N_1839,N_394);
nand U5579 (N_5579,N_1541,N_458);
nor U5580 (N_5580,N_472,N_462);
and U5581 (N_5581,N_3703,N_4608);
or U5582 (N_5582,N_4364,N_4938);
xnor U5583 (N_5583,N_1949,N_2945);
and U5584 (N_5584,N_2064,N_3648);
and U5585 (N_5585,N_2950,N_137);
xor U5586 (N_5586,N_2695,N_2482);
or U5587 (N_5587,N_4904,N_4612);
or U5588 (N_5588,N_961,N_1241);
nand U5589 (N_5589,N_4916,N_86);
nor U5590 (N_5590,N_2664,N_1195);
xor U5591 (N_5591,N_1948,N_1575);
and U5592 (N_5592,N_1747,N_4053);
nand U5593 (N_5593,N_441,N_4140);
xor U5594 (N_5594,N_419,N_1519);
or U5595 (N_5595,N_2220,N_4108);
xor U5596 (N_5596,N_3010,N_2346);
xor U5597 (N_5597,N_4234,N_1254);
and U5598 (N_5598,N_1569,N_4012);
or U5599 (N_5599,N_344,N_4789);
nand U5600 (N_5600,N_4801,N_30);
nor U5601 (N_5601,N_4778,N_4279);
nand U5602 (N_5602,N_2776,N_944);
nor U5603 (N_5603,N_3816,N_4568);
nor U5604 (N_5604,N_2278,N_2457);
nor U5605 (N_5605,N_3110,N_2377);
xnor U5606 (N_5606,N_1798,N_2015);
and U5607 (N_5607,N_2922,N_4319);
nor U5608 (N_5608,N_2315,N_3448);
nor U5609 (N_5609,N_4706,N_56);
nand U5610 (N_5610,N_3655,N_1935);
or U5611 (N_5611,N_3305,N_776);
nand U5612 (N_5612,N_654,N_1127);
xor U5613 (N_5613,N_3190,N_1365);
xnor U5614 (N_5614,N_2383,N_2367);
nand U5615 (N_5615,N_4952,N_1972);
xnor U5616 (N_5616,N_4634,N_1967);
nor U5617 (N_5617,N_43,N_3097);
xnor U5618 (N_5618,N_4746,N_1489);
nor U5619 (N_5619,N_3033,N_3250);
nor U5620 (N_5620,N_3917,N_4905);
and U5621 (N_5621,N_1369,N_2047);
and U5622 (N_5622,N_3621,N_2787);
nor U5623 (N_5623,N_811,N_4278);
xor U5624 (N_5624,N_3544,N_312);
nand U5625 (N_5625,N_4476,N_3564);
xnor U5626 (N_5626,N_4236,N_2421);
and U5627 (N_5627,N_3837,N_4090);
or U5628 (N_5628,N_1239,N_4558);
xnor U5629 (N_5629,N_2290,N_3916);
and U5630 (N_5630,N_4566,N_237);
nand U5631 (N_5631,N_4524,N_65);
and U5632 (N_5632,N_133,N_2998);
xnor U5633 (N_5633,N_2359,N_1146);
nand U5634 (N_5634,N_1281,N_2996);
and U5635 (N_5635,N_3613,N_3724);
or U5636 (N_5636,N_371,N_2110);
nor U5637 (N_5637,N_3167,N_953);
xor U5638 (N_5638,N_3570,N_733);
xor U5639 (N_5639,N_3390,N_1216);
nand U5640 (N_5640,N_320,N_4003);
nor U5641 (N_5641,N_4750,N_4399);
nand U5642 (N_5642,N_3020,N_456);
nand U5643 (N_5643,N_2204,N_4189);
nand U5644 (N_5644,N_668,N_3680);
xor U5645 (N_5645,N_2418,N_942);
and U5646 (N_5646,N_3826,N_2106);
nand U5647 (N_5647,N_744,N_3126);
nand U5648 (N_5648,N_485,N_207);
and U5649 (N_5649,N_2650,N_3769);
nand U5650 (N_5650,N_4562,N_1651);
or U5651 (N_5651,N_3176,N_4879);
nand U5652 (N_5652,N_1367,N_4513);
or U5653 (N_5653,N_2720,N_2522);
and U5654 (N_5654,N_2994,N_1157);
nor U5655 (N_5655,N_4393,N_629);
nor U5656 (N_5656,N_59,N_2937);
xnor U5657 (N_5657,N_2131,N_1494);
xnor U5658 (N_5658,N_3867,N_1324);
or U5659 (N_5659,N_2732,N_594);
xor U5660 (N_5660,N_2788,N_2181);
xor U5661 (N_5661,N_1280,N_1864);
nand U5662 (N_5662,N_3520,N_625);
nand U5663 (N_5663,N_2043,N_2102);
nor U5664 (N_5664,N_709,N_766);
or U5665 (N_5665,N_1787,N_4676);
nand U5666 (N_5666,N_2656,N_4668);
nor U5667 (N_5667,N_613,N_2108);
nand U5668 (N_5668,N_387,N_4756);
xnor U5669 (N_5669,N_941,N_1390);
nor U5670 (N_5670,N_2713,N_4218);
or U5671 (N_5671,N_3199,N_2266);
or U5672 (N_5672,N_2224,N_2154);
or U5673 (N_5673,N_380,N_4268);
xor U5674 (N_5674,N_1092,N_8);
nand U5675 (N_5675,N_3340,N_4760);
nand U5676 (N_5676,N_3362,N_4741);
nand U5677 (N_5677,N_4981,N_4478);
nor U5678 (N_5678,N_934,N_1330);
or U5679 (N_5679,N_2468,N_2890);
nand U5680 (N_5680,N_1439,N_4361);
nand U5681 (N_5681,N_916,N_4884);
nor U5682 (N_5682,N_3117,N_2279);
or U5683 (N_5683,N_2042,N_2973);
xor U5684 (N_5684,N_4252,N_430);
and U5685 (N_5685,N_2918,N_1309);
nor U5686 (N_5686,N_2934,N_488);
or U5687 (N_5687,N_3348,N_1838);
xnor U5688 (N_5688,N_3441,N_2534);
xnor U5689 (N_5689,N_3890,N_2509);
or U5690 (N_5690,N_3259,N_1617);
nand U5691 (N_5691,N_2985,N_2744);
or U5692 (N_5692,N_4743,N_3701);
and U5693 (N_5693,N_3646,N_4247);
nor U5694 (N_5694,N_2652,N_3873);
nor U5695 (N_5695,N_3739,N_4103);
xor U5696 (N_5696,N_773,N_4847);
nor U5697 (N_5697,N_1770,N_165);
xnor U5698 (N_5698,N_4351,N_602);
nand U5699 (N_5699,N_3967,N_491);
xor U5700 (N_5700,N_976,N_84);
or U5701 (N_5701,N_11,N_2698);
or U5702 (N_5702,N_1764,N_3498);
and U5703 (N_5703,N_2317,N_3414);
xor U5704 (N_5704,N_3354,N_336);
nand U5705 (N_5705,N_2453,N_4659);
and U5706 (N_5706,N_1944,N_2219);
and U5707 (N_5707,N_3529,N_3351);
and U5708 (N_5708,N_1418,N_2255);
or U5709 (N_5709,N_2665,N_927);
nand U5710 (N_5710,N_1430,N_3102);
xor U5711 (N_5711,N_3233,N_1392);
xor U5712 (N_5712,N_2854,N_4856);
or U5713 (N_5713,N_3854,N_1307);
nor U5714 (N_5714,N_92,N_3659);
or U5715 (N_5715,N_2580,N_2292);
nor U5716 (N_5716,N_609,N_1548);
nor U5717 (N_5717,N_792,N_4219);
and U5718 (N_5718,N_329,N_4450);
or U5719 (N_5719,N_884,N_2120);
nand U5720 (N_5720,N_2663,N_4563);
nor U5721 (N_5721,N_4968,N_4493);
xnor U5722 (N_5722,N_1556,N_3986);
nand U5723 (N_5723,N_2721,N_1420);
or U5724 (N_5724,N_546,N_861);
nand U5725 (N_5725,N_2944,N_3858);
nand U5726 (N_5726,N_3424,N_493);
xor U5727 (N_5727,N_4867,N_484);
nand U5728 (N_5728,N_988,N_914);
xor U5729 (N_5729,N_1974,N_1093);
xor U5730 (N_5730,N_4669,N_10);
or U5731 (N_5731,N_1743,N_4151);
or U5732 (N_5732,N_1775,N_260);
and U5733 (N_5733,N_3523,N_1412);
nand U5734 (N_5734,N_2976,N_554);
and U5735 (N_5735,N_3112,N_2830);
xnor U5736 (N_5736,N_243,N_1125);
and U5737 (N_5737,N_4680,N_3707);
nand U5738 (N_5738,N_4119,N_4689);
nand U5739 (N_5739,N_4818,N_2929);
nand U5740 (N_5740,N_150,N_120);
xor U5741 (N_5741,N_4223,N_1690);
nor U5742 (N_5742,N_4485,N_2345);
and U5743 (N_5743,N_3863,N_2610);
and U5744 (N_5744,N_1047,N_866);
xnor U5745 (N_5745,N_4649,N_3761);
and U5746 (N_5746,N_3575,N_4675);
xor U5747 (N_5747,N_388,N_1344);
nor U5748 (N_5748,N_3552,N_504);
xor U5749 (N_5749,N_2815,N_2535);
xor U5750 (N_5750,N_2262,N_2451);
nor U5751 (N_5751,N_2761,N_1756);
and U5752 (N_5752,N_1204,N_1581);
xor U5753 (N_5753,N_1180,N_4434);
xnor U5754 (N_5754,N_327,N_3347);
nor U5755 (N_5755,N_3094,N_3025);
nor U5756 (N_5756,N_3956,N_1613);
nor U5757 (N_5757,N_2193,N_478);
and U5758 (N_5758,N_4354,N_4772);
nand U5759 (N_5759,N_44,N_3760);
nor U5760 (N_5760,N_3795,N_4350);
xor U5761 (N_5761,N_17,N_3896);
nand U5762 (N_5762,N_4842,N_4974);
nor U5763 (N_5763,N_2158,N_366);
nand U5764 (N_5764,N_3047,N_2565);
and U5765 (N_5765,N_1679,N_1080);
xnor U5766 (N_5766,N_3221,N_561);
or U5767 (N_5767,N_132,N_936);
xnor U5768 (N_5768,N_3943,N_3254);
and U5769 (N_5769,N_1269,N_3157);
or U5770 (N_5770,N_4587,N_3392);
and U5771 (N_5771,N_4921,N_3734);
nand U5772 (N_5772,N_1849,N_228);
nand U5773 (N_5773,N_4212,N_341);
nand U5774 (N_5774,N_826,N_1788);
xor U5775 (N_5775,N_2480,N_1347);
or U5776 (N_5776,N_2486,N_2884);
or U5777 (N_5777,N_492,N_447);
nor U5778 (N_5778,N_3143,N_3706);
and U5779 (N_5779,N_4834,N_1606);
or U5780 (N_5780,N_3775,N_72);
nor U5781 (N_5781,N_497,N_3055);
nand U5782 (N_5782,N_4196,N_3987);
nor U5783 (N_5783,N_2411,N_2175);
nor U5784 (N_5784,N_1823,N_1018);
and U5785 (N_5785,N_4004,N_1450);
nand U5786 (N_5786,N_3951,N_1158);
xor U5787 (N_5787,N_2039,N_4102);
nor U5788 (N_5788,N_3545,N_3184);
nand U5789 (N_5789,N_3650,N_1129);
or U5790 (N_5790,N_4000,N_3557);
xor U5791 (N_5791,N_476,N_3984);
nor U5792 (N_5792,N_1376,N_2149);
xor U5793 (N_5793,N_3258,N_878);
nor U5794 (N_5794,N_2891,N_3532);
or U5795 (N_5795,N_2955,N_1794);
xor U5796 (N_5796,N_3411,N_3487);
or U5797 (N_5797,N_3211,N_1937);
nand U5798 (N_5798,N_197,N_3815);
nor U5799 (N_5799,N_2764,N_757);
or U5800 (N_5800,N_4021,N_4868);
nor U5801 (N_5801,N_4037,N_2203);
nand U5802 (N_5802,N_2007,N_3595);
or U5803 (N_5803,N_3839,N_3978);
nor U5804 (N_5804,N_2857,N_4333);
xor U5805 (N_5805,N_1491,N_428);
or U5806 (N_5806,N_931,N_4707);
nand U5807 (N_5807,N_390,N_4892);
xor U5808 (N_5808,N_3490,N_4999);
and U5809 (N_5809,N_2144,N_1225);
and U5810 (N_5810,N_1769,N_212);
and U5811 (N_5811,N_3922,N_3670);
nand U5812 (N_5812,N_2547,N_3612);
nor U5813 (N_5813,N_1530,N_3386);
and U5814 (N_5814,N_4505,N_4128);
xnor U5815 (N_5815,N_869,N_170);
or U5816 (N_5816,N_3913,N_615);
nor U5817 (N_5817,N_281,N_3654);
xnor U5818 (N_5818,N_3434,N_2438);
nand U5819 (N_5819,N_3732,N_4686);
nor U5820 (N_5820,N_2373,N_2006);
nor U5821 (N_5821,N_3954,N_2867);
nor U5822 (N_5822,N_3965,N_4919);
and U5823 (N_5823,N_1727,N_173);
or U5824 (N_5824,N_816,N_2646);
nor U5825 (N_5825,N_125,N_2055);
and U5826 (N_5826,N_4670,N_1094);
and U5827 (N_5827,N_3651,N_1683);
nor U5828 (N_5828,N_4704,N_190);
and U5829 (N_5829,N_4592,N_720);
nor U5830 (N_5830,N_420,N_3090);
or U5831 (N_5831,N_834,N_4201);
or U5832 (N_5832,N_2675,N_4465);
or U5833 (N_5833,N_402,N_1046);
and U5834 (N_5834,N_4611,N_3316);
nand U5835 (N_5835,N_1407,N_4866);
xnor U5836 (N_5836,N_4371,N_1763);
or U5837 (N_5837,N_929,N_102);
nor U5838 (N_5838,N_2,N_821);
xnor U5839 (N_5839,N_3068,N_3308);
nand U5840 (N_5840,N_3824,N_4006);
or U5841 (N_5841,N_1579,N_4837);
nand U5842 (N_5842,N_2678,N_450);
xnor U5843 (N_5843,N_302,N_3926);
nor U5844 (N_5844,N_4824,N_4641);
xnor U5845 (N_5845,N_309,N_571);
and U5846 (N_5846,N_951,N_1745);
nand U5847 (N_5847,N_2502,N_1468);
or U5848 (N_5848,N_568,N_239);
or U5849 (N_5849,N_2958,N_1623);
and U5850 (N_5850,N_685,N_3920);
nor U5851 (N_5851,N_1558,N_2378);
nand U5852 (N_5852,N_4324,N_3236);
xnor U5853 (N_5853,N_3942,N_4503);
or U5854 (N_5854,N_1635,N_3061);
nor U5855 (N_5855,N_3708,N_2592);
and U5856 (N_5856,N_4017,N_4389);
nor U5857 (N_5857,N_1279,N_3713);
nand U5858 (N_5858,N_1947,N_2053);
nor U5859 (N_5859,N_4031,N_835);
nand U5860 (N_5860,N_2807,N_1198);
xor U5861 (N_5861,N_3632,N_347);
or U5862 (N_5862,N_1182,N_2734);
nor U5863 (N_5863,N_4156,N_2640);
nor U5864 (N_5864,N_1143,N_1398);
nor U5865 (N_5865,N_1843,N_2268);
nor U5866 (N_5866,N_2543,N_4488);
or U5867 (N_5867,N_2188,N_1270);
or U5868 (N_5868,N_3450,N_2115);
nand U5869 (N_5869,N_333,N_3266);
nor U5870 (N_5870,N_2594,N_1642);
or U5871 (N_5871,N_3821,N_4918);
nor U5872 (N_5872,N_3421,N_2237);
nor U5873 (N_5873,N_726,N_3931);
nand U5874 (N_5874,N_498,N_247);
xor U5875 (N_5875,N_4081,N_4187);
and U5876 (N_5876,N_1227,N_2076);
xnor U5877 (N_5877,N_452,N_4947);
and U5878 (N_5878,N_1929,N_2878);
and U5879 (N_5879,N_2083,N_297);
or U5880 (N_5880,N_4489,N_740);
nor U5881 (N_5881,N_4932,N_480);
nor U5882 (N_5882,N_4416,N_3855);
xor U5883 (N_5883,N_932,N_61);
or U5884 (N_5884,N_1431,N_4072);
nor U5885 (N_5885,N_1252,N_3057);
nor U5886 (N_5886,N_4865,N_1840);
or U5887 (N_5887,N_3248,N_2322);
nand U5888 (N_5888,N_1222,N_2798);
nand U5889 (N_5889,N_1852,N_3842);
or U5890 (N_5890,N_3513,N_255);
nor U5891 (N_5891,N_1165,N_4085);
or U5892 (N_5892,N_4875,N_3806);
nand U5893 (N_5893,N_2683,N_3905);
or U5894 (N_5894,N_1996,N_894);
and U5895 (N_5895,N_2318,N_694);
nand U5896 (N_5896,N_2636,N_2716);
nand U5897 (N_5897,N_3969,N_57);
xnor U5898 (N_5898,N_1536,N_2874);
xor U5899 (N_5899,N_2005,N_3304);
and U5900 (N_5900,N_3799,N_4498);
xnor U5901 (N_5901,N_2205,N_1990);
or U5902 (N_5902,N_2368,N_3137);
nand U5903 (N_5903,N_4477,N_2601);
nand U5904 (N_5904,N_2736,N_3745);
nand U5905 (N_5905,N_3483,N_33);
xnor U5906 (N_5906,N_1654,N_2351);
xnor U5907 (N_5907,N_3495,N_2080);
or U5908 (N_5908,N_4646,N_666);
or U5909 (N_5909,N_1997,N_90);
and U5910 (N_5910,N_4703,N_1352);
xnor U5911 (N_5911,N_4208,N_115);
nor U5912 (N_5912,N_4061,N_3401);
nand U5913 (N_5913,N_4700,N_1219);
nor U5914 (N_5914,N_2523,N_1804);
nand U5915 (N_5915,N_1462,N_2034);
or U5916 (N_5916,N_3404,N_2422);
xor U5917 (N_5917,N_2880,N_4630);
nand U5918 (N_5918,N_4050,N_2387);
xnor U5919 (N_5919,N_2858,N_4474);
and U5920 (N_5920,N_3435,N_2758);
or U5921 (N_5921,N_1022,N_231);
xnor U5922 (N_5922,N_605,N_1302);
nor U5923 (N_5923,N_2781,N_4160);
nor U5924 (N_5924,N_1246,N_4297);
xnor U5925 (N_5925,N_4195,N_4312);
nor U5926 (N_5926,N_1482,N_2085);
xnor U5927 (N_5927,N_2146,N_4010);
and U5928 (N_5928,N_87,N_453);
and U5929 (N_5929,N_2916,N_88);
xnor U5930 (N_5930,N_2380,N_1294);
xnor U5931 (N_5931,N_64,N_1323);
or U5932 (N_5932,N_2247,N_3451);
or U5933 (N_5933,N_2602,N_238);
or U5934 (N_5934,N_591,N_3222);
or U5935 (N_5935,N_4664,N_1658);
or U5936 (N_5936,N_3519,N_4992);
nor U5937 (N_5937,N_1585,N_3073);
nand U5938 (N_5938,N_3358,N_1002);
nand U5939 (N_5939,N_4894,N_621);
nand U5940 (N_5940,N_4048,N_1992);
nor U5941 (N_5941,N_593,N_4539);
and U5942 (N_5942,N_4124,N_2651);
or U5943 (N_5943,N_1159,N_2036);
and U5944 (N_5944,N_824,N_4345);
or U5945 (N_5945,N_1291,N_973);
and U5946 (N_5946,N_4051,N_4486);
or U5947 (N_5947,N_4272,N_4747);
nor U5948 (N_5948,N_3013,N_1707);
or U5949 (N_5949,N_1121,N_2839);
and U5950 (N_5950,N_2932,N_2928);
nor U5951 (N_5951,N_4728,N_902);
xnor U5952 (N_5952,N_4662,N_798);
xnor U5953 (N_5953,N_4754,N_978);
or U5954 (N_5954,N_1504,N_1331);
nand U5955 (N_5955,N_3730,N_4433);
nand U5956 (N_5956,N_3449,N_4381);
and U5957 (N_5957,N_3518,N_4849);
nand U5958 (N_5958,N_4233,N_3507);
nor U5959 (N_5959,N_1604,N_1923);
nand U5960 (N_5960,N_2677,N_3095);
and U5961 (N_5961,N_2088,N_2882);
xor U5962 (N_5962,N_4092,N_4740);
and U5963 (N_5963,N_1035,N_448);
nor U5964 (N_5964,N_749,N_4888);
xor U5965 (N_5965,N_3321,N_3296);
nor U5966 (N_5966,N_2647,N_831);
nand U5967 (N_5967,N_1173,N_4194);
nand U5968 (N_5968,N_908,N_4016);
or U5969 (N_5969,N_995,N_680);
xnor U5970 (N_5970,N_1053,N_3383);
nand U5971 (N_5971,N_4621,N_4192);
nand U5972 (N_5972,N_711,N_2027);
nor U5973 (N_5973,N_1437,N_4183);
nand U5974 (N_5974,N_2514,N_2841);
xnor U5975 (N_5975,N_1178,N_786);
nand U5976 (N_5976,N_2044,N_576);
or U5977 (N_5977,N_2500,N_1771);
nand U5978 (N_5978,N_4270,N_2804);
or U5979 (N_5979,N_2904,N_851);
nor U5980 (N_5980,N_4762,N_2770);
nor U5981 (N_5981,N_4098,N_897);
and U5982 (N_5982,N_1013,N_4390);
and U5983 (N_5983,N_4521,N_1034);
and U5984 (N_5984,N_2430,N_1495);
nand U5985 (N_5985,N_2965,N_494);
nand U5986 (N_5986,N_317,N_1027);
or U5987 (N_5987,N_3814,N_1297);
nand U5988 (N_5988,N_3220,N_3086);
xnor U5989 (N_5989,N_2775,N_4636);
nor U5990 (N_5990,N_2388,N_3504);
and U5991 (N_5991,N_3709,N_2741);
xnor U5992 (N_5992,N_3462,N_735);
nand U5993 (N_5993,N_4419,N_2432);
xor U5994 (N_5994,N_1813,N_4677);
xor U5995 (N_5995,N_4609,N_3399);
or U5996 (N_5996,N_4104,N_4576);
nand U5997 (N_5997,N_1968,N_41);
nand U5998 (N_5998,N_4070,N_2372);
or U5999 (N_5999,N_1358,N_4432);
nor U6000 (N_6000,N_3737,N_4530);
nand U6001 (N_6001,N_2691,N_3864);
or U6002 (N_6002,N_3319,N_1312);
xnor U6003 (N_6003,N_815,N_3960);
xnor U6004 (N_6004,N_1100,N_3635);
nor U6005 (N_6005,N_2426,N_1386);
xnor U6006 (N_6006,N_3577,N_2189);
xor U6007 (N_6007,N_2615,N_2391);
and U6008 (N_6008,N_888,N_708);
xor U6009 (N_6009,N_1551,N_2635);
or U6010 (N_6010,N_4626,N_2216);
nor U6011 (N_6011,N_1527,N_4527);
xnor U6012 (N_6012,N_4808,N_4244);
nand U6013 (N_6013,N_3307,N_1218);
or U6014 (N_6014,N_4121,N_3566);
or U6015 (N_6015,N_1759,N_4133);
or U6016 (N_6016,N_3907,N_1354);
nand U6017 (N_6017,N_2915,N_848);
xnor U6018 (N_6018,N_3643,N_3219);
or U6019 (N_6019,N_3147,N_4052);
nor U6020 (N_6020,N_1534,N_4068);
nor U6021 (N_6021,N_3559,N_1315);
or U6022 (N_6022,N_1345,N_444);
xor U6023 (N_6023,N_1628,N_3881);
nor U6024 (N_6024,N_1510,N_747);
or U6025 (N_6025,N_2871,N_2476);
nand U6026 (N_6026,N_3755,N_3277);
and U6027 (N_6027,N_1485,N_4221);
or U6028 (N_6028,N_2242,N_3952);
and U6029 (N_6029,N_529,N_4036);
nand U6030 (N_6030,N_648,N_1387);
and U6031 (N_6031,N_2828,N_2993);
and U6032 (N_6032,N_580,N_345);
nor U6033 (N_6033,N_4306,N_2571);
xor U6034 (N_6034,N_4490,N_3974);
nor U6035 (N_6035,N_3540,N_2228);
and U6036 (N_6036,N_1784,N_156);
nand U6037 (N_6037,N_2089,N_4595);
and U6038 (N_6038,N_3173,N_3088);
xor U6039 (N_6039,N_27,N_566);
or U6040 (N_6040,N_3403,N_1098);
and U6041 (N_6041,N_2389,N_4603);
and U6042 (N_6042,N_1668,N_3869);
xnor U6043 (N_6043,N_3852,N_2963);
nand U6044 (N_6044,N_2530,N_784);
or U6045 (N_6045,N_2754,N_4840);
nor U6046 (N_6046,N_2824,N_2562);
xnor U6047 (N_6047,N_1220,N_2778);
nor U6048 (N_6048,N_2362,N_3085);
nand U6049 (N_6049,N_2612,N_4069);
nor U6050 (N_6050,N_2078,N_587);
xor U6051 (N_6051,N_4925,N_1191);
or U6052 (N_6052,N_2087,N_828);
and U6053 (N_6053,N_3180,N_686);
xnor U6054 (N_6054,N_4533,N_1982);
nor U6055 (N_6055,N_4744,N_714);
or U6056 (N_6056,N_4736,N_4095);
and U6057 (N_6057,N_3479,N_2316);
and U6058 (N_6058,N_4770,N_4074);
or U6059 (N_6059,N_39,N_4311);
or U6060 (N_6060,N_2957,N_517);
or U6061 (N_6061,N_1078,N_1461);
xor U6062 (N_6062,N_3663,N_523);
or U6063 (N_6063,N_3381,N_3644);
and U6064 (N_6064,N_945,N_1750);
nor U6065 (N_6065,N_3289,N_2271);
or U6066 (N_6066,N_2557,N_3662);
nand U6067 (N_6067,N_562,N_3264);
nor U6068 (N_6068,N_3743,N_4501);
and U6069 (N_6069,N_4773,N_1049);
xor U6070 (N_6070,N_4714,N_542);
or U6071 (N_6071,N_4640,N_339);
xor U6072 (N_6072,N_1876,N_783);
and U6073 (N_6073,N_4480,N_1978);
xor U6074 (N_6074,N_1299,N_3924);
nor U6075 (N_6075,N_2287,N_2139);
xnor U6076 (N_6076,N_2208,N_435);
or U6077 (N_6077,N_3626,N_465);
or U6078 (N_6078,N_1273,N_3834);
and U6079 (N_6079,N_746,N_1128);
xor U6080 (N_6080,N_3464,N_867);
and U6081 (N_6081,N_3599,N_1169);
and U6082 (N_6082,N_405,N_301);
nand U6083 (N_6083,N_2433,N_863);
nor U6084 (N_6084,N_1103,N_1414);
and U6085 (N_6085,N_538,N_3165);
xor U6086 (N_6086,N_2862,N_4788);
nand U6087 (N_6087,N_4650,N_2513);
xor U6088 (N_6088,N_3961,N_2616);
or U6089 (N_6089,N_1350,N_900);
xnor U6090 (N_6090,N_543,N_323);
and U6091 (N_6091,N_871,N_1676);
or U6092 (N_6092,N_3060,N_2049);
and U6093 (N_6093,N_66,N_219);
nand U6094 (N_6094,N_1117,N_2423);
and U6095 (N_6095,N_1871,N_1719);
or U6096 (N_6096,N_4654,N_752);
nor U6097 (N_6097,N_1610,N_4671);
nand U6098 (N_6098,N_3198,N_2623);
nor U6099 (N_6099,N_2084,N_2805);
nand U6100 (N_6100,N_411,N_3491);
or U6101 (N_6101,N_2397,N_3027);
or U6102 (N_6102,N_2023,N_4737);
nor U6103 (N_6103,N_1809,N_3325);
nor U6104 (N_6104,N_1036,N_1408);
nand U6105 (N_6105,N_2861,N_1911);
or U6106 (N_6106,N_352,N_1711);
xor U6107 (N_6107,N_1023,N_2567);
xor U6108 (N_6108,N_3050,N_4519);
and U6109 (N_6109,N_75,N_4067);
and U6110 (N_6110,N_2641,N_4158);
xor U6111 (N_6111,N_1957,N_2933);
and U6112 (N_6112,N_1147,N_938);
xor U6113 (N_6113,N_2173,N_3808);
nor U6114 (N_6114,N_3722,N_4957);
nand U6115 (N_6115,N_4246,N_2926);
nor U6116 (N_6116,N_3408,N_4739);
nand U6117 (N_6117,N_551,N_4543);
and U6118 (N_6118,N_3139,N_206);
nor U6119 (N_6119,N_1912,N_2093);
nor U6120 (N_6120,N_463,N_731);
xnor U6121 (N_6121,N_684,N_2289);
xor U6122 (N_6122,N_1185,N_3113);
nor U6123 (N_6123,N_4348,N_531);
and U6124 (N_6124,N_1520,N_1332);
nand U6125 (N_6125,N_1740,N_53);
nor U6126 (N_6126,N_4560,N_3130);
nand U6127 (N_6127,N_598,N_1962);
nor U6128 (N_6128,N_1983,N_3607);
and U6129 (N_6129,N_362,N_4889);
xnor U6130 (N_6130,N_3202,N_1939);
and U6131 (N_6131,N_1674,N_254);
and U6132 (N_6132,N_42,N_4084);
or U6133 (N_6133,N_1909,N_2728);
or U6134 (N_6134,N_1636,N_2284);
nand U6135 (N_6135,N_4615,N_2537);
or U6136 (N_6136,N_2544,N_3923);
nor U6137 (N_6137,N_1985,N_1619);
xnor U6138 (N_6138,N_4178,N_3601);
or U6139 (N_6139,N_3062,N_4363);
or U6140 (N_6140,N_4264,N_1631);
or U6141 (N_6141,N_4666,N_3959);
nor U6142 (N_6142,N_3818,N_1063);
xor U6143 (N_6143,N_1830,N_2020);
xor U6144 (N_6144,N_9,N_2054);
nor U6145 (N_6145,N_1591,N_2114);
nor U6146 (N_6146,N_920,N_349);
xnor U6147 (N_6147,N_4858,N_4229);
and U6148 (N_6148,N_4321,N_3310);
nor U6149 (N_6149,N_3938,N_530);
and U6150 (N_6150,N_3791,N_2356);
and U6151 (N_6151,N_2197,N_2863);
xnor U6152 (N_6152,N_4966,N_3368);
and U6153 (N_6153,N_4209,N_4713);
nand U6154 (N_6154,N_2872,N_85);
xor U6155 (N_6155,N_3789,N_1692);
xnor U6156 (N_6156,N_2086,N_3776);
nand U6157 (N_6157,N_4964,N_2756);
nand U6158 (N_6158,N_762,N_4112);
or U6159 (N_6159,N_1247,N_2925);
xor U6160 (N_6160,N_3541,N_983);
nor U6161 (N_6161,N_1207,N_129);
nor U6162 (N_6162,N_570,N_2723);
nor U6163 (N_6163,N_1731,N_2939);
or U6164 (N_6164,N_4088,N_2735);
or U6165 (N_6165,N_4804,N_3948);
nor U6166 (N_6166,N_1041,N_2556);
or U6167 (N_6167,N_38,N_719);
nand U6168 (N_6168,N_1089,N_4276);
nand U6169 (N_6169,N_2337,N_3582);
xor U6170 (N_6170,N_3885,N_3785);
and U6171 (N_6171,N_732,N_1123);
nand U6172 (N_6172,N_4930,N_49);
nor U6173 (N_6173,N_3395,N_918);
and U6174 (N_6174,N_3,N_2265);
and U6175 (N_6175,N_3669,N_710);
xnor U6176 (N_6176,N_4705,N_4285);
nor U6177 (N_6177,N_2107,N_3527);
nor U6178 (N_6178,N_4020,N_3282);
nor U6179 (N_6179,N_2866,N_2393);
or U6180 (N_6180,N_1678,N_3023);
or U6181 (N_6181,N_1471,N_2869);
nand U6182 (N_6182,N_982,N_2603);
or U6183 (N_6183,N_1015,N_4660);
nand U6184 (N_6184,N_2967,N_4575);
or U6185 (N_6185,N_363,N_3243);
or U6186 (N_6186,N_122,N_1563);
or U6187 (N_6187,N_1069,N_1895);
nor U6188 (N_6188,N_1951,N_1245);
xnor U6189 (N_6189,N_4873,N_372);
and U6190 (N_6190,N_957,N_3428);
and U6191 (N_6191,N_3042,N_1580);
or U6192 (N_6192,N_105,N_906);
and U6193 (N_6193,N_3973,N_2598);
xnor U6194 (N_6194,N_4534,N_4959);
and U6195 (N_6195,N_3944,N_2997);
nand U6196 (N_6196,N_3946,N_2398);
nor U6197 (N_6197,N_664,N_4441);
nor U6198 (N_6198,N_544,N_1875);
xnor U6199 (N_6199,N_3262,N_1824);
and U6200 (N_6200,N_3350,N_2038);
xor U6201 (N_6201,N_1977,N_924);
nor U6202 (N_6202,N_1684,N_4692);
nand U6203 (N_6203,N_4627,N_1209);
nand U6204 (N_6204,N_3615,N_2155);
nand U6205 (N_6205,N_3474,N_513);
nand U6206 (N_6206,N_1807,N_3140);
nand U6207 (N_6207,N_1135,N_244);
nor U6208 (N_6208,N_2358,N_4910);
nand U6209 (N_6209,N_1612,N_4922);
nand U6210 (N_6210,N_1155,N_1261);
or U6211 (N_6211,N_178,N_392);
nand U6212 (N_6212,N_4120,N_1277);
xor U6213 (N_6213,N_946,N_2831);
nor U6214 (N_6214,N_2644,N_227);
xor U6215 (N_6215,N_3071,N_2050);
nor U6216 (N_6216,N_1934,N_911);
xnor U6217 (N_6217,N_4153,N_4580);
and U6218 (N_6218,N_3716,N_2150);
nor U6219 (N_6219,N_2504,N_1649);
and U6220 (N_6220,N_1778,N_2743);
or U6221 (N_6221,N_4217,N_2583);
nand U6222 (N_6222,N_4948,N_1341);
or U6223 (N_6223,N_154,N_2286);
and U6224 (N_6224,N_3719,N_2355);
or U6225 (N_6225,N_4355,N_681);
or U6226 (N_6226,N_887,N_3131);
and U6227 (N_6227,N_4656,N_2302);
nand U6228 (N_6228,N_717,N_3271);
and U6229 (N_6229,N_1552,N_3283);
and U6230 (N_6230,N_4199,N_4541);
or U6231 (N_6231,N_291,N_4352);
and U6232 (N_6232,N_3456,N_4076);
or U6233 (N_6233,N_1533,N_2608);
nand U6234 (N_6234,N_2628,N_4502);
xnor U6235 (N_6235,N_4869,N_1625);
nand U6236 (N_6236,N_3778,N_1256);
nor U6237 (N_6237,N_2014,N_1898);
xor U6238 (N_6238,N_1950,N_1528);
nor U6239 (N_6239,N_1285,N_1284);
or U6240 (N_6240,N_3256,N_4383);
nor U6241 (N_6241,N_3628,N_4665);
nand U6242 (N_6242,N_2236,N_1019);
nor U6243 (N_6243,N_1265,N_3215);
and U6244 (N_6244,N_3991,N_3391);
xnor U6245 (N_6245,N_968,N_2126);
and U6246 (N_6246,N_4186,N_1088);
xnor U6247 (N_6247,N_1038,N_4309);
xnor U6248 (N_6248,N_1564,N_2257);
and U6249 (N_6249,N_3823,N_2165);
nand U6250 (N_6250,N_4418,N_3605);
nor U6251 (N_6251,N_1130,N_4165);
or U6252 (N_6252,N_135,N_1557);
nor U6253 (N_6253,N_1567,N_4710);
xor U6254 (N_6254,N_69,N_3129);
and U6255 (N_6255,N_4973,N_4643);
nor U6256 (N_6256,N_3335,N_361);
xnor U6257 (N_6257,N_2177,N_2104);
xor U6258 (N_6258,N_797,N_3849);
nand U6259 (N_6259,N_3329,N_1725);
nand U6260 (N_6260,N_1796,N_952);
xor U6261 (N_6261,N_2376,N_1498);
nor U6262 (N_6262,N_1050,N_1810);
nand U6263 (N_6263,N_3301,N_1189);
xor U6264 (N_6264,N_4047,N_4681);
xor U6265 (N_6265,N_3076,N_3702);
and U6266 (N_6266,N_2123,N_3809);
nand U6267 (N_6267,N_241,N_1693);
xor U6268 (N_6268,N_1487,N_791);
xor U6269 (N_6269,N_4197,N_3488);
xnor U6270 (N_6270,N_1643,N_1877);
nand U6271 (N_6271,N_558,N_3638);
and U6272 (N_6272,N_4325,N_4965);
or U6273 (N_6273,N_3135,N_3935);
and U6274 (N_6274,N_2747,N_3070);
and U6275 (N_6275,N_169,N_3306);
nand U6276 (N_6276,N_495,N_1698);
and U6277 (N_6277,N_3216,N_4181);
xnor U6278 (N_6278,N_4997,N_3556);
nand U6279 (N_6279,N_1845,N_1938);
nand U6280 (N_6280,N_1434,N_2182);
or U6281 (N_6281,N_3046,N_4495);
nand U6282 (N_6282,N_3156,N_3249);
nor U6283 (N_6283,N_391,N_2613);
and U6284 (N_6284,N_4699,N_1111);
nand U6285 (N_6285,N_3384,N_2171);
xnor U6286 (N_6286,N_3125,N_700);
nor U6287 (N_6287,N_2814,N_3910);
and U6288 (N_6288,N_2551,N_3265);
nand U6289 (N_6289,N_812,N_25);
or U6290 (N_6290,N_424,N_4451);
nand U6291 (N_6291,N_3590,N_1956);
xnor U6292 (N_6292,N_508,N_657);
xnor U6293 (N_6293,N_1382,N_2419);
and U6294 (N_6294,N_4225,N_3146);
nand U6295 (N_6295,N_4555,N_1989);
xor U6296 (N_6296,N_1161,N_2936);
xor U6297 (N_6297,N_3688,N_1926);
nor U6298 (N_6298,N_2642,N_2692);
xor U6299 (N_6299,N_2660,N_4369);
nor U6300 (N_6300,N_4280,N_1870);
or U6301 (N_6301,N_1998,N_3835);
xnor U6302 (N_6302,N_4023,N_4823);
and U6303 (N_6303,N_3438,N_4454);
nor U6304 (N_6304,N_240,N_271);
nand U6305 (N_6305,N_15,N_3048);
nor U6306 (N_6306,N_1891,N_2138);
or U6307 (N_6307,N_2406,N_2739);
or U6308 (N_6308,N_4424,N_1887);
and U6309 (N_6309,N_2342,N_4427);
or U6310 (N_6310,N_4956,N_429);
nor U6311 (N_6311,N_4777,N_3000);
nand U6312 (N_6312,N_3225,N_24);
and U6313 (N_6313,N_3893,N_3803);
and U6314 (N_6314,N_1837,N_2130);
nand U6315 (N_6315,N_50,N_1435);
nor U6316 (N_6316,N_671,N_4881);
xor U6317 (N_6317,N_3290,N_1104);
nand U6318 (N_6318,N_2525,N_4030);
nor U6319 (N_6319,N_471,N_322);
nor U6320 (N_6320,N_3481,N_1174);
or U6321 (N_6321,N_1385,N_3342);
nor U6322 (N_6322,N_2763,N_1517);
or U6323 (N_6323,N_838,N_3484);
nand U6324 (N_6324,N_2883,N_2835);
or U6325 (N_6325,N_2481,N_4556);
nand U6326 (N_6326,N_4584,N_4909);
and U6327 (N_6327,N_707,N_400);
nand U6328 (N_6328,N_4046,N_3588);
or U6329 (N_6329,N_2075,N_4593);
xor U6330 (N_6330,N_365,N_803);
or U6331 (N_6331,N_367,N_703);
nor U6332 (N_6332,N_4396,N_1008);
or U6333 (N_6333,N_3208,N_3128);
nand U6334 (N_6334,N_407,N_2907);
and U6335 (N_6335,N_3882,N_2634);
xnor U6336 (N_6336,N_2230,N_1488);
and U6337 (N_6337,N_3526,N_2185);
or U6338 (N_6338,N_2860,N_1594);
xor U6339 (N_6339,N_1721,N_706);
nand U6340 (N_6340,N_2524,N_3618);
and U6341 (N_6341,N_1084,N_4839);
nor U6342 (N_6342,N_4633,N_3983);
and U6343 (N_6343,N_2714,N_2467);
xnor U6344 (N_6344,N_3217,N_653);
and U6345 (N_6345,N_1406,N_2407);
nand U6346 (N_6346,N_257,N_4731);
nand U6347 (N_6347,N_3728,N_2914);
and U6348 (N_6348,N_2347,N_287);
nand U6349 (N_6349,N_4753,N_2267);
and U6350 (N_6350,N_1059,N_4296);
or U6351 (N_6351,N_3442,N_3547);
and U6352 (N_6352,N_1403,N_600);
and U6353 (N_6353,N_4588,N_3270);
xnor U6354 (N_6354,N_192,N_3554);
and U6355 (N_6355,N_3511,N_3276);
and U6356 (N_6356,N_2951,N_256);
nor U6357 (N_6357,N_4803,N_4228);
or U6358 (N_6358,N_775,N_1188);
nor U6359 (N_6359,N_1709,N_3279);
xnor U6360 (N_6360,N_2576,N_2585);
and U6361 (N_6361,N_4648,N_3833);
nor U6362 (N_6362,N_3338,N_1716);
or U6363 (N_6363,N_3921,N_2294);
xnor U6364 (N_6364,N_473,N_2920);
and U6365 (N_6365,N_3617,N_2722);
or U6366 (N_6366,N_1587,N_2441);
or U6367 (N_6367,N_858,N_28);
nor U6368 (N_6368,N_1848,N_261);
or U6369 (N_6369,N_1576,N_3990);
nor U6370 (N_6370,N_822,N_4761);
nand U6371 (N_6371,N_4220,N_501);
and U6372 (N_6372,N_2638,N_3109);
nor U6373 (N_6373,N_1055,N_4805);
and U6374 (N_6374,N_2809,N_1624);
nor U6375 (N_6375,N_470,N_4845);
xor U6376 (N_6376,N_2343,N_292);
nand U6377 (N_6377,N_2812,N_2990);
and U6378 (N_6378,N_4548,N_3992);
and U6379 (N_6379,N_3345,N_3014);
xnor U6380 (N_6380,N_3295,N_1068);
nand U6381 (N_6381,N_3149,N_696);
and U6382 (N_6382,N_1832,N_3872);
nor U6383 (N_6383,N_890,N_162);
xor U6384 (N_6384,N_4411,N_4585);
nor U6385 (N_6385,N_2099,N_364);
or U6386 (N_6386,N_1704,N_4902);
nand U6387 (N_6387,N_4812,N_3822);
xnor U6388 (N_6388,N_2465,N_2187);
xor U6389 (N_6389,N_1702,N_3827);
nor U6390 (N_6390,N_4570,N_550);
nand U6391 (N_6391,N_23,N_1134);
nor U6392 (N_6392,N_4863,N_3366);
xnor U6393 (N_6393,N_1192,N_3466);
xor U6394 (N_6394,N_1366,N_3697);
nand U6395 (N_6395,N_1067,N_1416);
nor U6396 (N_6396,N_2595,N_2109);
and U6397 (N_6397,N_4398,N_4720);
nor U6398 (N_6398,N_4164,N_2826);
nor U6399 (N_6399,N_489,N_4540);
and U6400 (N_6400,N_3029,N_3170);
nor U6401 (N_6401,N_631,N_299);
nand U6402 (N_6402,N_1521,N_959);
nand U6403 (N_6403,N_1754,N_690);
nor U6404 (N_6404,N_559,N_4931);
and U6405 (N_6405,N_3649,N_3247);
and U6406 (N_6406,N_1920,N_4796);
and U6407 (N_6407,N_2533,N_2607);
or U6408 (N_6408,N_2696,N_3997);
or U6409 (N_6409,N_140,N_3185);
nor U6410 (N_6410,N_3953,N_4086);
and U6411 (N_6411,N_1395,N_1799);
nand U6412 (N_6412,N_2605,N_2331);
nor U6413 (N_6413,N_3596,N_4742);
nand U6414 (N_6414,N_2786,N_1463);
nor U6415 (N_6415,N_4444,N_876);
or U6416 (N_6416,N_1449,N_2100);
nand U6417 (N_6417,N_1011,N_2172);
nand U6418 (N_6418,N_236,N_3423);
and U6419 (N_6419,N_4438,N_1592);
nand U6420 (N_6420,N_2491,N_2227);
and U6421 (N_6421,N_4987,N_903);
and U6422 (N_6422,N_1806,N_1234);
nor U6423 (N_6423,N_4726,N_4308);
nand U6424 (N_6424,N_2496,N_1897);
nand U6425 (N_6425,N_1514,N_4300);
and U6426 (N_6426,N_1706,N_4267);
or U6427 (N_6427,N_31,N_1348);
nand U6428 (N_6428,N_139,N_2532);
nor U6429 (N_6429,N_1099,N_915);
xnor U6430 (N_6430,N_839,N_4042);
xnor U6431 (N_6431,N_4370,N_922);
nor U6432 (N_6432,N_4241,N_4961);
or U6433 (N_6433,N_3120,N_3166);
and U6434 (N_6434,N_2978,N_4806);
nor U6435 (N_6435,N_1931,N_4203);
and U6436 (N_6436,N_4607,N_2330);
nand U6437 (N_6437,N_4996,N_4064);
nor U6438 (N_6438,N_1109,N_1744);
xor U6439 (N_6439,N_2536,N_4841);
xnor U6440 (N_6440,N_967,N_4452);
and U6441 (N_6441,N_1083,N_4365);
or U6442 (N_6442,N_2906,N_2309);
nor U6443 (N_6443,N_4846,N_2385);
xor U6444 (N_6444,N_1196,N_3640);
or U6445 (N_6445,N_2408,N_3430);
nor U6446 (N_6446,N_2836,N_1286);
xnor U6447 (N_6447,N_2902,N_4397);
xor U6448 (N_6448,N_1237,N_526);
xor U6449 (N_6449,N_2454,N_3229);
or U6450 (N_6450,N_3273,N_426);
nor U6451 (N_6451,N_2654,N_3633);
xnor U6452 (N_6452,N_3624,N_3658);
xnor U6453 (N_6453,N_2245,N_1549);
or U6454 (N_6454,N_332,N_4138);
or U6455 (N_6455,N_2969,N_4005);
nand U6456 (N_6456,N_524,N_3218);
nand U6457 (N_6457,N_1076,N_21);
xnor U6458 (N_6458,N_1388,N_2898);
nor U6459 (N_6459,N_2579,N_1325);
or U6460 (N_6460,N_3083,N_3820);
or U6461 (N_6461,N_855,N_1212);
or U6462 (N_6462,N_753,N_2134);
nand U6463 (N_6463,N_1186,N_4978);
nor U6464 (N_6464,N_4473,N_2234);
nand U6465 (N_6465,N_395,N_97);
nor U6466 (N_6466,N_2680,N_548);
nor U6467 (N_6467,N_469,N_2324);
xnor U6468 (N_6468,N_3542,N_3995);
xnor U6469 (N_6469,N_3665,N_4515);
nand U6470 (N_6470,N_2733,N_2668);
nand U6471 (N_6471,N_3067,N_4123);
nor U6472 (N_6472,N_3589,N_2212);
xnor U6473 (N_6473,N_4287,N_4790);
or U6474 (N_6474,N_2669,N_3045);
nand U6475 (N_6475,N_623,N_646);
or U6476 (N_6476,N_3172,N_3018);
and U6477 (N_6477,N_4644,N_4065);
nand U6478 (N_6478,N_3418,N_2382);
xnor U6479 (N_6479,N_3235,N_4358);
or U6480 (N_6480,N_853,N_218);
and U6481 (N_6481,N_1044,N_4625);
and U6482 (N_6482,N_2328,N_4690);
or U6483 (N_6483,N_3417,N_2291);
nand U6484 (N_6484,N_2853,N_188);
or U6485 (N_6485,N_2202,N_2439);
and U6486 (N_6486,N_3762,N_1343);
and U6487 (N_6487,N_2604,N_2729);
nor U6488 (N_6488,N_128,N_4586);
and U6489 (N_6489,N_3251,N_4142);
or U6490 (N_6490,N_3324,N_1681);
and U6491 (N_6491,N_3087,N_4780);
nor U6492 (N_6492,N_1629,N_3819);
and U6493 (N_6493,N_2352,N_2750);
nand U6494 (N_6494,N_883,N_813);
nand U6495 (N_6495,N_2464,N_4177);
nand U6496 (N_6496,N_3955,N_4026);
nor U6497 (N_6497,N_2213,N_4783);
xnor U6498 (N_6498,N_439,N_535);
nor U6499 (N_6499,N_1217,N_4645);
xnor U6500 (N_6500,N_4449,N_2972);
or U6501 (N_6501,N_4941,N_4483);
and U6502 (N_6502,N_3751,N_2427);
nor U6503 (N_6503,N_2283,N_2768);
and U6504 (N_6504,N_246,N_1970);
and U6505 (N_6505,N_3525,N_850);
and U6506 (N_6506,N_393,N_3093);
nor U6507 (N_6507,N_2276,N_2135);
xor U6508 (N_6508,N_1932,N_2164);
or U6509 (N_6509,N_2403,N_4035);
nand U6510 (N_6510,N_2068,N_1272);
xnor U6511 (N_6511,N_1682,N_4014);
nand U6512 (N_6512,N_801,N_3431);
nor U6513 (N_6513,N_2335,N_111);
and U6514 (N_6514,N_248,N_3341);
xor U6515 (N_6515,N_2301,N_2390);
or U6516 (N_6516,N_3536,N_3639);
nand U6517 (N_6517,N_3446,N_2774);
nor U6518 (N_6518,N_3528,N_4439);
and U6519 (N_6519,N_4721,N_2767);
and U6520 (N_6520,N_588,N_3726);
or U6521 (N_6521,N_3004,N_194);
nor U6522 (N_6522,N_4807,N_555);
xnor U6523 (N_6523,N_1755,N_2966);
or U6524 (N_6524,N_790,N_1881);
xnor U6525 (N_6525,N_3963,N_833);
or U6526 (N_6526,N_3378,N_4500);
or U6527 (N_6527,N_2116,N_2582);
or U6528 (N_6528,N_4951,N_641);
nand U6529 (N_6529,N_3238,N_2360);
and U6530 (N_6530,N_804,N_563);
and U6531 (N_6531,N_2707,N_177);
and U6532 (N_6532,N_557,N_1156);
nor U6533 (N_6533,N_4724,N_1132);
or U6534 (N_6534,N_300,N_2298);
nand U6535 (N_6535,N_1405,N_3084);
and U6536 (N_6536,N_819,N_3111);
or U6537 (N_6537,N_1081,N_3311);
or U6538 (N_6538,N_4269,N_3427);
and U6539 (N_6539,N_3081,N_2485);
or U6540 (N_6540,N_3592,N_2827);
or U6541 (N_6541,N_2896,N_4787);
or U6542 (N_6542,N_928,N_2125);
nand U6543 (N_6543,N_4632,N_3336);
and U6544 (N_6544,N_1667,N_1499);
and U6545 (N_6545,N_652,N_1789);
or U6546 (N_6546,N_412,N_1941);
nor U6547 (N_6547,N_3191,N_1056);
nor U6548 (N_6548,N_3227,N_4258);
xor U6549 (N_6549,N_3798,N_721);
nor U6550 (N_6550,N_4289,N_2410);
or U6551 (N_6551,N_4935,N_2031);
xor U6552 (N_6552,N_1308,N_3327);
xor U6553 (N_6553,N_2771,N_895);
nor U6554 (N_6554,N_3664,N_265);
nor U6555 (N_6555,N_375,N_1873);
or U6556 (N_6556,N_787,N_2277);
or U6557 (N_6557,N_3505,N_2434);
nor U6558 (N_6558,N_1221,N_4409);
xnor U6559 (N_6559,N_3376,N_1267);
or U6560 (N_6560,N_3998,N_1440);
nand U6561 (N_6561,N_146,N_1040);
and U6562 (N_6562,N_2338,N_3979);
nor U6563 (N_6563,N_2192,N_619);
xnor U6564 (N_6564,N_1215,N_507);
xor U6565 (N_6565,N_3750,N_1210);
or U6566 (N_6566,N_3373,N_4833);
and U6567 (N_6567,N_3535,N_1588);
nor U6568 (N_6568,N_2473,N_3996);
nor U6569 (N_6569,N_225,N_1131);
xnor U6570 (N_6570,N_374,N_2850);
nor U6571 (N_6571,N_62,N_2024);
and U6572 (N_6572,N_1164,N_1168);
and U6573 (N_6573,N_4211,N_224);
and U6574 (N_6574,N_1399,N_1922);
or U6575 (N_6575,N_1695,N_160);
or U6576 (N_6576,N_4631,N_4360);
and U6577 (N_6577,N_2145,N_3848);
and U6578 (N_6578,N_541,N_2773);
and U6579 (N_6579,N_1547,N_4606);
nand U6580 (N_6580,N_2992,N_1163);
and U6581 (N_6581,N_1114,N_670);
and U6582 (N_6582,N_2159,N_4404);
nor U6583 (N_6583,N_1597,N_1052);
xor U6584 (N_6584,N_157,N_2987);
nor U6585 (N_6585,N_1136,N_4210);
xnor U6586 (N_6586,N_3313,N_3223);
nor U6587 (N_6587,N_1031,N_1283);
nor U6588 (N_6588,N_2333,N_3467);
and U6589 (N_6589,N_482,N_4019);
and U6590 (N_6590,N_1326,N_2693);
and U6591 (N_6591,N_3422,N_2353);
nand U6592 (N_6592,N_4537,N_954);
nand U6593 (N_6593,N_2682,N_1289);
nor U6594 (N_6594,N_2264,N_2013);
nand U6595 (N_6595,N_882,N_4307);
xor U6596 (N_6596,N_2416,N_3597);
nor U6597 (N_6597,N_2545,N_4202);
and U6598 (N_6598,N_817,N_3206);
nor U6599 (N_6599,N_2240,N_457);
and U6600 (N_6600,N_3232,N_3192);
or U6601 (N_6601,N_496,N_1444);
nand U6602 (N_6602,N_4368,N_2117);
and U6603 (N_6603,N_1574,N_1413);
or U6604 (N_6604,N_1584,N_910);
and U6605 (N_6605,N_220,N_2002);
nor U6606 (N_6606,N_1009,N_4698);
or U6607 (N_6607,N_3226,N_4243);
and U6608 (N_6608,N_1661,N_3947);
nand U6609 (N_6609,N_4526,N_1773);
and U6610 (N_6610,N_2575,N_4377);
nand U6611 (N_6611,N_1954,N_2584);
xor U6612 (N_6612,N_3899,N_1632);
nor U6613 (N_6613,N_3794,N_4635);
nor U6614 (N_6614,N_1525,N_3239);
or U6615 (N_6615,N_2995,N_718);
and U6616 (N_6616,N_1728,N_1275);
nand U6617 (N_6617,N_123,N_687);
nor U6618 (N_6618,N_617,N_3372);
and U6619 (N_6619,N_1568,N_253);
nand U6620 (N_6620,N_972,N_4175);
nand U6621 (N_6621,N_4367,N_2254);
and U6622 (N_6622,N_4388,N_4768);
nand U6623 (N_6623,N_2162,N_1524);
nor U6624 (N_6624,N_1058,N_4955);
or U6625 (N_6625,N_1699,N_4590);
xor U6626 (N_6626,N_1139,N_2495);
nor U6627 (N_6627,N_1757,N_4984);
nor U6628 (N_6628,N_545,N_2912);
nand U6629 (N_6629,N_1017,N_2561);
nand U6630 (N_6630,N_2487,N_3886);
or U6631 (N_6631,N_4286,N_715);
and U6632 (N_6632,N_2621,N_3098);
nor U6633 (N_6633,N_3091,N_3405);
xnor U6634 (N_6634,N_89,N_2401);
or U6635 (N_6635,N_267,N_4089);
or U6636 (N_6636,N_519,N_4538);
nor U6637 (N_6637,N_2253,N_3193);
and U6638 (N_6638,N_1640,N_213);
nand U6639 (N_6639,N_1577,N_4610);
or U6640 (N_6640,N_2270,N_3746);
xor U6641 (N_6641,N_4828,N_1075);
nor U6642 (N_6642,N_516,N_4683);
and U6643 (N_6643,N_1738,N_4765);
or U6644 (N_6644,N_4263,N_4083);
nand U6645 (N_6645,N_1819,N_40);
nand U6646 (N_6646,N_3766,N_4155);
xnor U6647 (N_6647,N_2244,N_487);
and U6648 (N_6648,N_606,N_4039);
nand U6649 (N_6649,N_2941,N_2069);
nor U6650 (N_6650,N_2310,N_268);
nor U6651 (N_6651,N_3367,N_1701);
or U6652 (N_6652,N_3257,N_3614);
nor U6653 (N_6653,N_1793,N_4702);
nor U6654 (N_6654,N_4946,N_1710);
or U6655 (N_6655,N_3008,N_3912);
and U6656 (N_6656,N_2864,N_4429);
or U6657 (N_6657,N_682,N_3502);
nor U6658 (N_6658,N_432,N_1133);
and U6659 (N_6659,N_1443,N_369);
nor U6660 (N_6660,N_4716,N_2440);
nand U6661 (N_6661,N_1359,N_2587);
xor U6662 (N_6662,N_875,N_3452);
nor U6663 (N_6663,N_1540,N_2964);
nand U6664 (N_6664,N_1242,N_665);
nand U6665 (N_6665,N_2095,N_475);
or U6666 (N_6666,N_537,N_279);
nand U6667 (N_6667,N_2541,N_4825);
nor U6668 (N_6668,N_2474,N_4771);
and U6669 (N_6669,N_2336,N_4299);
nor U6670 (N_6670,N_3763,N_3246);
nor U6671 (N_6671,N_185,N_3234);
and U6672 (N_6672,N_2045,N_330);
nand U6673 (N_6673,N_3468,N_4394);
xor U6674 (N_6674,N_3059,N_427);
nor U6675 (N_6675,N_2622,N_4497);
and U6676 (N_6676,N_4793,N_3530);
nor U6677 (N_6677,N_4057,N_734);
nand U6678 (N_6678,N_1030,N_4775);
nor U6679 (N_6679,N_4338,N_539);
or U6680 (N_6680,N_870,N_4041);
xnor U6681 (N_6681,N_993,N_2501);
nor U6682 (N_6682,N_167,N_1979);
nor U6683 (N_6683,N_4266,N_2740);
nor U6684 (N_6684,N_645,N_1503);
and U6685 (N_6685,N_907,N_1320);
nand U6686 (N_6686,N_4013,N_250);
or U6687 (N_6687,N_2913,N_1509);
nor U6688 (N_6688,N_3846,N_4844);
or U6689 (N_6689,N_2223,N_3274);
nor U6690 (N_6690,N_4647,N_3684);
xnor U6691 (N_6691,N_661,N_2759);
nand U6692 (N_6692,N_1214,N_2097);
xor U6693 (N_6693,N_1079,N_4376);
nand U6694 (N_6694,N_1313,N_104);
and U6695 (N_6695,N_2975,N_1866);
nor U6696 (N_6696,N_1975,N_3379);
or U6697 (N_6697,N_245,N_2092);
and U6698 (N_6698,N_1883,N_354);
xnor U6699 (N_6699,N_1902,N_3773);
and U6700 (N_6700,N_4582,N_4843);
xor U6701 (N_6701,N_63,N_4767);
nor U6702 (N_6702,N_112,N_4122);
and U6703 (N_6703,N_2908,N_3209);
or U6704 (N_6704,N_4514,N_1351);
nor U6705 (N_6705,N_315,N_3561);
xor U6706 (N_6706,N_3284,N_321);
xnor U6707 (N_6707,N_4549,N_4436);
xnor U6708 (N_6708,N_2507,N_716);
and U6709 (N_6709,N_4991,N_4604);
nand U6710 (N_6710,N_3735,N_4529);
and U6711 (N_6711,N_1936,N_807);
xor U6712 (N_6712,N_4174,N_1401);
nand U6713 (N_6713,N_3105,N_446);
nor U6714 (N_6714,N_76,N_1644);
or U6715 (N_6715,N_1532,N_4437);
and U6716 (N_6716,N_575,N_4314);
and U6717 (N_6717,N_1199,N_2201);
xor U6718 (N_6718,N_1523,N_3420);
xnor U6719 (N_6719,N_3508,N_4148);
or U6720 (N_6720,N_590,N_1110);
nand U6721 (N_6721,N_896,N_1316);
nand U6722 (N_6722,N_4583,N_1772);
nand U6723 (N_6723,N_4043,N_2470);
and U6724 (N_6724,N_1486,N_2577);
nand U6725 (N_6725,N_1537,N_1452);
or U6726 (N_6726,N_3883,N_1634);
and U6727 (N_6727,N_1244,N_16);
and U6728 (N_6728,N_4385,N_3162);
nand U6729 (N_6729,N_3962,N_730);
and U6730 (N_6730,N_2186,N_1202);
nand U6731 (N_6731,N_4431,N_1235);
xnor U6732 (N_6732,N_3171,N_4898);
or U6733 (N_6733,N_3939,N_844);
xnor U6734 (N_6734,N_1007,N_2570);
nor U6735 (N_6735,N_4482,N_499);
nand U6736 (N_6736,N_2374,N_2983);
nand U6737 (N_6737,N_449,N_1713);
and U6738 (N_6738,N_2058,N_2478);
nand U6739 (N_6739,N_3593,N_2140);
nand U6740 (N_6740,N_3784,N_4018);
xnor U6741 (N_6741,N_3400,N_3200);
nor U6742 (N_6742,N_3514,N_1638);
xor U6743 (N_6743,N_4599,N_4292);
and U6744 (N_6744,N_437,N_1758);
and U6745 (N_6745,N_3182,N_1337);
and U6746 (N_6746,N_1073,N_2755);
xor U6747 (N_6747,N_2684,N_1821);
and U6748 (N_6748,N_2306,N_396);
or U6749 (N_6749,N_759,N_4425);
nor U6750 (N_6750,N_3744,N_209);
xnor U6751 (N_6751,N_4797,N_3850);
xnor U6752 (N_6752,N_1596,N_3660);
nor U6753 (N_6753,N_2596,N_506);
nor U6754 (N_6754,N_4954,N_1593);
nor U6755 (N_6755,N_2659,N_4687);
and U6756 (N_6756,N_126,N_2312);
or U6757 (N_6757,N_1586,N_4564);
or U6758 (N_6758,N_1293,N_2810);
nand U6759 (N_6759,N_1203,N_0);
xor U6760 (N_6760,N_2709,N_3079);
or U6761 (N_6761,N_4346,N_4723);
or U6762 (N_6762,N_1397,N_4091);
and U6763 (N_6763,N_2161,N_2349);
or U6764 (N_6764,N_2832,N_4242);
and U6765 (N_6765,N_2953,N_4885);
or U6766 (N_6766,N_2210,N_2160);
and U6767 (N_6767,N_2344,N_1243);
nand U6768 (N_6768,N_777,N_1835);
nor U6769 (N_6769,N_4882,N_74);
nand U6770 (N_6770,N_2339,N_175);
and U6771 (N_6771,N_3269,N_2238);
nand U6772 (N_6772,N_868,N_4062);
and U6773 (N_6773,N_4150,N_2314);
and U6774 (N_6774,N_2793,N_1404);
and U6775 (N_6775,N_4557,N_2548);
xor U6776 (N_6776,N_4605,N_534);
or U6777 (N_6777,N_2293,N_2961);
xor U6778 (N_6778,N_1687,N_2511);
and U6779 (N_6779,N_1952,N_2578);
nor U6780 (N_6780,N_578,N_4316);
and U6781 (N_6781,N_4782,N_3851);
xor U6782 (N_6782,N_3163,N_4551);
nand U6783 (N_6783,N_5,N_3036);
and U6784 (N_6784,N_3937,N_3297);
xor U6785 (N_6785,N_1820,N_4757);
xnor U6786 (N_6786,N_4763,N_3661);
xor U6787 (N_6787,N_1329,N_4479);
and U6788 (N_6788,N_2105,N_1201);
nor U6789 (N_6789,N_2424,N_3692);
nor U6790 (N_6790,N_204,N_2288);
nor U6791 (N_6791,N_1924,N_520);
or U6792 (N_6792,N_4034,N_1615);
nand U6793 (N_6793,N_1892,N_3994);
nand U6794 (N_6794,N_4032,N_1037);
nor U6795 (N_6795,N_338,N_3813);
nand U6796 (N_6796,N_2988,N_3830);
and U6797 (N_6797,N_1751,N_1600);
nor U6798 (N_6798,N_1181,N_3825);
nand U6799 (N_6799,N_3875,N_2258);
or U6800 (N_6800,N_3158,N_3127);
nor U6801 (N_6801,N_2449,N_2327);
and U6802 (N_6802,N_3275,N_3011);
or U6803 (N_6803,N_1171,N_1375);
xnor U6804 (N_6804,N_399,N_1479);
nand U6805 (N_6805,N_2198,N_704);
nor U6806 (N_6806,N_2749,N_3668);
and U6807 (N_6807,N_981,N_585);
xnor U6808 (N_6808,N_4906,N_1802);
xor U6809 (N_6809,N_2630,N_1633);
nand U6810 (N_6810,N_4679,N_1953);
or U6811 (N_6811,N_4414,N_316);
or U6812 (N_6812,N_3178,N_4523);
and U6813 (N_6813,N_3856,N_342);
or U6814 (N_6814,N_2248,N_234);
or U6815 (N_6815,N_1797,N_2811);
or U6816 (N_6816,N_1228,N_4392);
xnor U6817 (N_6817,N_2119,N_4274);
or U6818 (N_6818,N_1826,N_4637);
nor U6819 (N_6819,N_806,N_229);
or U6820 (N_6820,N_1197,N_1535);
and U6821 (N_6821,N_2679,N_2472);
and U6822 (N_6822,N_2757,N_2179);
nand U6823 (N_6823,N_2923,N_4347);
and U6824 (N_6824,N_3729,N_1363);
nor U6825 (N_6825,N_3181,N_48);
and U6826 (N_6826,N_4897,N_454);
nand U6827 (N_6827,N_171,N_1394);
nand U6828 (N_6828,N_1650,N_2477);
nand U6829 (N_6829,N_1,N_1457);
and U6830 (N_6830,N_3026,N_2029);
nand U6831 (N_6831,N_2170,N_964);
or U6832 (N_6832,N_1253,N_1020);
xor U6833 (N_6833,N_155,N_1317);
xor U6834 (N_6834,N_1539,N_2738);
and U6835 (N_6835,N_4188,N_1106);
xor U6836 (N_6836,N_189,N_3385);
or U6837 (N_6837,N_3710,N_847);
xor U6838 (N_6838,N_780,N_83);
nor U6839 (N_6839,N_3294,N_2450);
nand U6840 (N_6840,N_2281,N_4166);
nand U6841 (N_6841,N_4857,N_3134);
nor U6842 (N_6842,N_3674,N_3473);
xnor U6843 (N_6843,N_1785,N_370);
nand U6844 (N_6844,N_70,N_4831);
nand U6845 (N_6845,N_4125,N_4457);
nor U6846 (N_6846,N_1342,N_1648);
nor U6847 (N_6847,N_874,N_285);
nor U6848 (N_6848,N_4214,N_4715);
or U6849 (N_6849,N_1298,N_4168);
xor U6850 (N_6850,N_1453,N_3145);
and U6851 (N_6851,N_3207,N_1973);
and U6852 (N_6852,N_2948,N_1915);
nor U6853 (N_6853,N_2760,N_2261);
xnor U6854 (N_6854,N_3749,N_2924);
or U6855 (N_6855,N_479,N_58);
nand U6856 (N_6856,N_1206,N_3880);
and U6857 (N_6857,N_3300,N_3476);
and U6858 (N_6858,N_117,N_4);
or U6859 (N_6859,N_2190,N_2949);
and U6860 (N_6860,N_642,N_3571);
nor U6861 (N_6861,N_728,N_763);
xor U6862 (N_6862,N_1472,N_1112);
nand U6863 (N_6863,N_4028,N_532);
xor U6864 (N_6864,N_1288,N_4871);
and U6865 (N_6865,N_502,N_2329);
and U6866 (N_6866,N_3317,N_4907);
and U6867 (N_6867,N_269,N_172);
and U6868 (N_6868,N_3562,N_3394);
and U6869 (N_6869,N_3877,N_3679);
or U6870 (N_6870,N_93,N_862);
and U6871 (N_6871,N_2569,N_2065);
nor U6872 (N_6872,N_3902,N_592);
or U6873 (N_6873,N_4343,N_251);
nor U6874 (N_6874,N_1496,N_1236);
nor U6875 (N_6875,N_2004,N_46);
nand U6876 (N_6876,N_2538,N_4386);
xnor U6877 (N_6877,N_3028,N_1927);
nand U6878 (N_6878,N_2784,N_4132);
or U6879 (N_6879,N_4950,N_2947);
nand U6880 (N_6880,N_2703,N_2231);
nor U6881 (N_6881,N_1458,N_4544);
nand U6882 (N_6882,N_4380,N_4007);
and U6883 (N_6883,N_1999,N_3471);
nor U6884 (N_6884,N_723,N_4172);
nor U6885 (N_6885,N_2153,N_4913);
nor U6886 (N_6886,N_4116,N_1200);
xnor U6887 (N_6887,N_2256,N_136);
xnor U6888 (N_6888,N_4344,N_4678);
nand U6889 (N_6889,N_966,N_289);
and U6890 (N_6890,N_644,N_846);
and U6891 (N_6891,N_3136,N_4176);
xnor U6892 (N_6892,N_2404,N_1969);
or U6893 (N_6893,N_649,N_379);
or U6894 (N_6894,N_4491,N_3627);
or U6895 (N_6895,N_350,N_4310);
and U6896 (N_6896,N_2559,N_3685);
nor U6897 (N_6897,N_1656,N_3477);
and U6898 (N_6898,N_2539,N_2040);
nand U6899 (N_6899,N_2456,N_3859);
nor U6900 (N_6900,N_3767,N_4231);
or U6901 (N_6901,N_4934,N_1368);
and U6902 (N_6902,N_1921,N_917);
xnor U6903 (N_6903,N_756,N_4597);
xnor U6904 (N_6904,N_1672,N_1513);
xnor U6905 (N_6905,N_1995,N_3261);
xor U6906 (N_6906,N_52,N_2803);
nor U6907 (N_6907,N_1167,N_3396);
nor U6908 (N_6908,N_837,N_1896);
nand U6909 (N_6909,N_4506,N_3263);
nand U6910 (N_6910,N_4579,N_3915);
nor U6911 (N_6911,N_2489,N_2572);
or U6912 (N_6912,N_2895,N_2848);
nor U6913 (N_6913,N_1515,N_738);
and U6914 (N_6914,N_1816,N_1665);
and U6915 (N_6915,N_3318,N_854);
and U6916 (N_6916,N_769,N_4261);
nand U6917 (N_6917,N_655,N_4940);
nand U6918 (N_6918,N_2063,N_1900);
nor U6919 (N_6919,N_4520,N_337);
and U6920 (N_6920,N_956,N_741);
or U6921 (N_6921,N_3860,N_4126);
xnor U6922 (N_6922,N_4998,N_3522);
or U6923 (N_6923,N_2405,N_636);
xor U6924 (N_6924,N_2645,N_2200);
and U6925 (N_6925,N_1729,N_3573);
nand U6926 (N_6926,N_3204,N_4545);
or U6927 (N_6927,N_880,N_277);
nand U6928 (N_6928,N_4336,N_3039);
and U6929 (N_6929,N_840,N_1448);
and U6930 (N_6930,N_1389,N_724);
or U6931 (N_6931,N_4695,N_2365);
and U6932 (N_6932,N_210,N_282);
nand U6933 (N_6933,N_1064,N_2431);
nand U6934 (N_6934,N_2542,N_4712);
nand U6935 (N_6935,N_1160,N_2772);
or U6936 (N_6936,N_295,N_2011);
nand U6937 (N_6937,N_980,N_2762);
nand U6938 (N_6938,N_940,N_977);
xnor U6939 (N_6939,N_2540,N_3497);
nor U6940 (N_6940,N_4567,N_4685);
and U6941 (N_6941,N_4733,N_2369);
and U6942 (N_6942,N_2147,N_1565);
xnor U6943 (N_6943,N_99,N_3712);
nor U6944 (N_6944,N_4508,N_2469);
or U6945 (N_6945,N_3186,N_986);
nand U6946 (N_6946,N_3188,N_51);
nor U6947 (N_6947,N_4589,N_2852);
nor U6948 (N_6948,N_1266,N_176);
or U6949 (N_6949,N_2529,N_3868);
xor U6950 (N_6950,N_1696,N_1822);
and U6951 (N_6951,N_892,N_1459);
xor U6952 (N_6952,N_4323,N_4464);
and U6953 (N_6953,N_434,N_699);
nand U6954 (N_6954,N_1511,N_1024);
or U6955 (N_6955,N_4256,N_3925);
and U6956 (N_6956,N_3253,N_2751);
or U6957 (N_6957,N_3817,N_258);
xnor U6958 (N_6958,N_3549,N_4983);
or U6959 (N_6959,N_1874,N_2025);
nand U6960 (N_6960,N_4661,N_4878);
nor U6961 (N_6961,N_14,N_2658);
nor U6962 (N_6962,N_2845,N_3103);
nand U6963 (N_6963,N_2070,N_3683);
xnor U6964 (N_6964,N_164,N_180);
or U6965 (N_6965,N_2528,N_2554);
xor U6966 (N_6966,N_3230,N_226);
nand U6967 (N_6967,N_2681,N_859);
xnor U6968 (N_6968,N_622,N_1908);
xnor U6969 (N_6969,N_3482,N_2321);
or U6970 (N_6970,N_1641,N_4990);
nand U6971 (N_6971,N_4949,N_1422);
nor U6972 (N_6972,N_2834,N_970);
or U6973 (N_6973,N_4516,N_3069);
nand U6974 (N_6974,N_29,N_1262);
xor U6975 (N_6975,N_34,N_589);
nor U6976 (N_6976,N_127,N_3397);
xor U6977 (N_6977,N_1357,N_1627);
nand U6978 (N_6978,N_2719,N_4059);
or U6979 (N_6979,N_1451,N_4060);
and U6980 (N_6980,N_3374,N_2348);
or U6981 (N_6981,N_1795,N_2455);
or U6982 (N_6982,N_1529,N_1697);
xor U6983 (N_6983,N_2960,N_4657);
or U6984 (N_6984,N_3757,N_505);
xor U6985 (N_6985,N_1790,N_134);
and U6986 (N_6986,N_1304,N_3579);
xor U6987 (N_6987,N_2823,N_1620);
or U6988 (N_6988,N_864,N_4809);
nor U6989 (N_6989,N_425,N_4430);
and U6990 (N_6990,N_764,N_2061);
and U6991 (N_6991,N_304,N_612);
nand U6992 (N_6992,N_2030,N_4204);
nor U6993 (N_6993,N_4106,N_3741);
and U6994 (N_6994,N_990,N_4638);
nand U6995 (N_6995,N_60,N_3988);
nand U6996 (N_6996,N_4117,N_4303);
xnor U6997 (N_6997,N_4463,N_4471);
or U6998 (N_6998,N_2394,N_574);
or U6999 (N_6999,N_4071,N_1077);
nand U7000 (N_7000,N_1240,N_1087);
nor U7001 (N_7001,N_1177,N_3429);
or U7002 (N_7002,N_2032,N_4401);
nand U7003 (N_7003,N_2648,N_3328);
or U7004 (N_7004,N_4302,N_2332);
nor U7005 (N_7005,N_4810,N_4373);
and U7006 (N_7006,N_3558,N_183);
or U7007 (N_7007,N_3058,N_3927);
nor U7008 (N_7008,N_1854,N_382);
nand U7009 (N_7009,N_4745,N_604);
nand U7010 (N_7010,N_436,N_2494);
or U7011 (N_7011,N_2662,N_937);
nor U7012 (N_7012,N_1039,N_4722);
nand U7013 (N_7013,N_179,N_2785);
or U7014 (N_7014,N_793,N_1184);
xnor U7015 (N_7015,N_1735,N_4237);
nand U7016 (N_7016,N_4986,N_3194);
nor U7017 (N_7017,N_1065,N_3982);
xor U7018 (N_7018,N_3293,N_4620);
or U7019 (N_7019,N_2688,N_3138);
or U7020 (N_7020,N_1303,N_3320);
and U7021 (N_7021,N_4682,N_1205);
nand U7022 (N_7022,N_948,N_2071);
or U7023 (N_7023,N_4799,N_3898);
or U7024 (N_7024,N_3169,N_4157);
and U7025 (N_7025,N_2655,N_1971);
or U7026 (N_7026,N_3278,N_2968);
nand U7027 (N_7027,N_2851,N_3066);
or U7028 (N_7028,N_4143,N_1599);
xor U7029 (N_7029,N_1327,N_4420);
and U7030 (N_7030,N_1473,N_1377);
or U7031 (N_7031,N_2797,N_13);
nor U7032 (N_7032,N_2199,N_3516);
nand U7033 (N_7033,N_116,N_1090);
nand U7034 (N_7034,N_885,N_4063);
or U7035 (N_7035,N_2766,N_3811);
nand U7036 (N_7036,N_306,N_4139);
nand U7037 (N_7037,N_1605,N_4691);
or U7038 (N_7038,N_3472,N_4100);
xor U7039 (N_7039,N_1425,N_1733);
or U7040 (N_7040,N_4349,N_2817);
nand U7041 (N_7041,N_2591,N_2077);
and U7042 (N_7042,N_1561,N_110);
and U7043 (N_7043,N_4008,N_3056);
nand U7044 (N_7044,N_4518,N_2196);
xnor U7045 (N_7045,N_3032,N_616);
xnor U7046 (N_7046,N_413,N_1383);
xnor U7047 (N_7047,N_3177,N_3804);
nor U7048 (N_7048,N_1901,N_3758);
and U7049 (N_7049,N_1705,N_2384);
xor U7050 (N_7050,N_232,N_683);
and U7051 (N_7051,N_4462,N_2887);
nand U7052 (N_7052,N_2429,N_2381);
xnor U7053 (N_7053,N_1259,N_676);
or U7054 (N_7054,N_2492,N_1768);
xnor U7055 (N_7055,N_4162,N_131);
nor U7056 (N_7056,N_3693,N_4629);
nand U7057 (N_7057,N_2445,N_4730);
or U7058 (N_7058,N_4118,N_1669);
or U7059 (N_7059,N_3122,N_1717);
and U7060 (N_7060,N_962,N_2479);
or U7061 (N_7061,N_651,N_4494);
xor U7062 (N_7062,N_290,N_77);
nor U7063 (N_7063,N_4550,N_4732);
xnor U7064 (N_7064,N_431,N_1739);
or U7065 (N_7065,N_2447,N_3682);
nor U7066 (N_7066,N_1720,N_3364);
nand U7067 (N_7067,N_3779,N_3016);
nand U7068 (N_7068,N_3678,N_4387);
or U7069 (N_7069,N_4331,N_3214);
nor U7070 (N_7070,N_2879,N_771);
nand U7071 (N_7071,N_3078,N_1531);
xnor U7072 (N_7072,N_203,N_4769);
nor U7073 (N_7073,N_2518,N_2782);
nand U7074 (N_7074,N_3892,N_514);
xnor U7075 (N_7075,N_1179,N_4357);
xor U7076 (N_7076,N_4619,N_4260);
nand U7077 (N_7077,N_2700,N_4830);
or U7078 (N_7078,N_3132,N_1752);
xor U7079 (N_7079,N_303,N_1287);
or U7080 (N_7080,N_3977,N_2940);
xor U7081 (N_7081,N_3616,N_1856);
xnor U7082 (N_7082,N_4301,N_1879);
and U7083 (N_7083,N_3934,N_184);
nand U7084 (N_7084,N_343,N_3439);
nor U7085 (N_7085,N_3393,N_4816);
nor U7086 (N_7086,N_1860,N_991);
nor U7087 (N_7087,N_4853,N_264);
nor U7088 (N_7088,N_1006,N_779);
nand U7089 (N_7089,N_389,N_1945);
xnor U7090 (N_7090,N_3802,N_2313);
or U7091 (N_7091,N_2564,N_4758);
nor U7092 (N_7092,N_4226,N_2962);
or U7093 (N_7093,N_3426,N_1680);
nand U7094 (N_7094,N_3432,N_1396);
xor U7095 (N_7095,N_800,N_2295);
nor U7096 (N_7096,N_4322,N_1421);
or U7097 (N_7097,N_2619,N_3681);
and U7098 (N_7098,N_1867,N_1815);
and U7099 (N_7099,N_3619,N_1777);
nor U7100 (N_7100,N_1714,N_2323);
nand U7101 (N_7101,N_667,N_1988);
or U7102 (N_7102,N_4407,N_1595);
and U7103 (N_7103,N_4838,N_1516);
nor U7104 (N_7104,N_3696,N_4870);
xnor U7105 (N_7105,N_3288,N_1258);
or U7106 (N_7106,N_3591,N_2712);
or U7107 (N_7107,N_2849,N_3976);
and U7108 (N_7108,N_1208,N_1703);
nor U7109 (N_7109,N_3019,N_3704);
and U7110 (N_7110,N_3667,N_3865);
and U7111 (N_7111,N_2484,N_4509);
and U7112 (N_7112,N_1115,N_3377);
xnor U7113 (N_7113,N_2588,N_2752);
nand U7114 (N_7114,N_3642,N_2174);
and U7115 (N_7115,N_2837,N_3344);
and U7116 (N_7116,N_3560,N_663);
or U7117 (N_7117,N_2018,N_340);
or U7118 (N_7118,N_1961,N_2041);
or U7119 (N_7119,N_2137,N_1170);
xor U7120 (N_7120,N_2901,N_984);
nand U7121 (N_7121,N_781,N_1553);
and U7122 (N_7122,N_318,N_1965);
xor U7123 (N_7123,N_4281,N_1862);
and U7124 (N_7124,N_4340,N_1033);
xor U7125 (N_7125,N_1502,N_4329);
nor U7126 (N_7126,N_3521,N_1477);
nor U7127 (N_7127,N_1940,N_181);
nor U7128 (N_7128,N_163,N_4015);
xnor U7129 (N_7129,N_1779,N_2597);
or U7130 (N_7130,N_1166,N_1410);
and U7131 (N_7131,N_215,N_1118);
nand U7132 (N_7132,N_2233,N_3630);
and U7133 (N_7133,N_418,N_3606);
or U7134 (N_7134,N_4859,N_346);
nor U7135 (N_7135,N_1918,N_3114);
xor U7136 (N_7136,N_483,N_3012);
or U7137 (N_7137,N_2483,N_4374);
nor U7138 (N_7138,N_3461,N_55);
nand U7139 (N_7139,N_705,N_3168);
nand U7140 (N_7140,N_4027,N_3909);
nand U7141 (N_7141,N_856,N_78);
nor U7142 (N_7142,N_1086,N_4829);
nand U7143 (N_7143,N_1724,N_1096);
nor U7144 (N_7144,N_1626,N_3460);
nor U7145 (N_7145,N_2876,N_221);
xnor U7146 (N_7146,N_4467,N_7);
and U7147 (N_7147,N_4546,N_1314);
xor U7148 (N_7148,N_477,N_1029);
nor U7149 (N_7149,N_2825,N_799);
xor U7150 (N_7150,N_1426,N_3805);
nor U7151 (N_7151,N_2725,N_3119);
nand U7152 (N_7152,N_1190,N_1858);
nand U7153 (N_7153,N_3889,N_2444);
nor U7154 (N_7154,N_4613,N_4623);
nand U7155 (N_7155,N_2214,N_3054);
or U7156 (N_7156,N_4179,N_992);
and U7157 (N_7157,N_3096,N_403);
xor U7158 (N_7158,N_2215,N_4304);
xor U7159 (N_7159,N_3534,N_2209);
nor U7160 (N_7160,N_3009,N_1346);
or U7161 (N_7161,N_3568,N_4198);
xor U7162 (N_7162,N_3365,N_2019);
xor U7163 (N_7163,N_4161,N_4759);
xnor U7164 (N_7164,N_3337,N_1151);
nand U7165 (N_7165,N_2629,N_2180);
or U7166 (N_7166,N_1814,N_4696);
or U7167 (N_7167,N_4190,N_2008);
xnor U7168 (N_7168,N_4356,N_1573);
and U7169 (N_7169,N_3985,N_108);
nand U7170 (N_7170,N_4752,N_331);
xnor U7171 (N_7171,N_3410,N_1335);
nor U7172 (N_7172,N_4738,N_2073);
xnor U7173 (N_7173,N_3765,N_2979);
or U7174 (N_7174,N_935,N_1149);
xnor U7175 (N_7175,N_1708,N_3299);
or U7176 (N_7176,N_2581,N_1828);
and U7177 (N_7177,N_3064,N_2183);
or U7178 (N_7178,N_4146,N_3475);
nor U7179 (N_7179,N_1894,N_1846);
xnor U7180 (N_7180,N_438,N_1647);
or U7181 (N_7181,N_2606,N_3099);
and U7182 (N_7182,N_3782,N_2488);
nor U7183 (N_7183,N_564,N_4265);
nor U7184 (N_7184,N_2816,N_1522);
xor U7185 (N_7185,N_2742,N_3930);
or U7186 (N_7186,N_679,N_3966);
and U7187 (N_7187,N_1652,N_4958);
or U7188 (N_7188,N_1108,N_4135);
and U7189 (N_7189,N_1356,N_4458);
xor U7190 (N_7190,N_2672,N_1603);
and U7191 (N_7191,N_1436,N_3001);
and U7192 (N_7192,N_4492,N_1657);
or U7193 (N_7193,N_1054,N_2091);
nor U7194 (N_7194,N_692,N_4900);
and U7195 (N_7195,N_2152,N_4835);
nor U7196 (N_7196,N_2274,N_4251);
or U7197 (N_7197,N_3210,N_4044);
nand U7198 (N_7198,N_2753,N_81);
nand U7199 (N_7199,N_2066,N_2010);
and U7200 (N_7200,N_351,N_2059);
nand U7201 (N_7201,N_4571,N_2618);
and U7202 (N_7202,N_4821,N_2379);
and U7203 (N_7203,N_2868,N_2009);
and U7204 (N_7204,N_4320,N_4784);
and U7205 (N_7205,N_3620,N_68);
and U7206 (N_7206,N_2631,N_440);
nor U7207 (N_7207,N_2017,N_4395);
nor U7208 (N_7208,N_3645,N_4009);
xnor U7209 (N_7209,N_262,N_923);
or U7210 (N_7210,N_865,N_2503);
xor U7211 (N_7211,N_4811,N_1715);
nand U7212 (N_7212,N_2026,N_2919);
or U7213 (N_7213,N_1880,N_3604);
nand U7214 (N_7214,N_4283,N_3268);
nand U7215 (N_7215,N_500,N_1748);
nor U7216 (N_7216,N_3407,N_1555);
nand U7217 (N_7217,N_4184,N_1655);
or U7218 (N_7218,N_4697,N_4096);
nor U7219 (N_7219,N_2035,N_579);
nand U7220 (N_7220,N_843,N_4862);
nor U7221 (N_7221,N_4443,N_4078);
or U7222 (N_7222,N_3416,N_4275);
and U7223 (N_7223,N_270,N_947);
and U7224 (N_7224,N_2458,N_1238);
nand U7225 (N_7225,N_4764,N_4776);
and U7226 (N_7226,N_3154,N_4022);
and U7227 (N_7227,N_4573,N_3594);
nor U7228 (N_7228,N_1694,N_1101);
or U7229 (N_7229,N_1670,N_4144);
or U7230 (N_7230,N_3608,N_1043);
nand U7231 (N_7231,N_1292,N_1249);
and U7232 (N_7232,N_1691,N_3121);
or U7233 (N_7233,N_113,N_1371);
and U7234 (N_7234,N_2082,N_152);
xor U7235 (N_7235,N_2250,N_3272);
nand U7236 (N_7236,N_4294,N_2326);
xnor U7237 (N_7237,N_71,N_3533);
or U7238 (N_7238,N_3343,N_2900);
xor U7239 (N_7239,N_601,N_3241);
or U7240 (N_7240,N_3756,N_2927);
xor U7241 (N_7241,N_3388,N_2531);
xnor U7242 (N_7242,N_2791,N_4254);
nand U7243 (N_7243,N_4725,N_3829);
nor U7244 (N_7244,N_138,N_999);
and U7245 (N_7245,N_54,N_960);
nand U7246 (N_7246,N_191,N_3150);
nand U7247 (N_7247,N_4512,N_2094);
or U7248 (N_7248,N_2614,N_360);
nand U7249 (N_7249,N_2527,N_3870);
nor U7250 (N_7250,N_1943,N_1582);
and U7251 (N_7251,N_3578,N_1122);
nand U7252 (N_7252,N_1905,N_3787);
nand U7253 (N_7253,N_2903,N_4093);
xor U7254 (N_7254,N_1966,N_2910);
nor U7255 (N_7255,N_4058,N_2493);
nor U7256 (N_7256,N_2699,N_4353);
and U7257 (N_7257,N_4929,N_2111);
nand U7258 (N_7258,N_4578,N_2673);
xnor U7259 (N_7259,N_1417,N_307);
and U7260 (N_7260,N_3499,N_4255);
xor U7261 (N_7261,N_4851,N_2510);
and U7262 (N_7262,N_3574,N_1045);
and U7263 (N_7263,N_3255,N_2098);
and U7264 (N_7264,N_4814,N_4169);
or U7265 (N_7265,N_1872,N_2168);
nor U7266 (N_7266,N_4448,N_4547);
or U7267 (N_7267,N_2666,N_560);
nor U7268 (N_7268,N_3334,N_1571);
xor U7269 (N_7269,N_1379,N_4191);
nand U7270 (N_7270,N_1889,N_1765);
and U7271 (N_7271,N_2818,N_949);
xnor U7272 (N_7272,N_103,N_1506);
nand U7273 (N_7273,N_1378,N_2475);
nor U7274 (N_7274,N_2420,N_3906);
xnor U7275 (N_7275,N_3469,N_2334);
and U7276 (N_7276,N_1353,N_4475);
xnor U7277 (N_7277,N_1409,N_3298);
nand U7278 (N_7278,N_2060,N_4684);
nor U7279 (N_7279,N_1834,N_3292);
xnor U7280 (N_7280,N_4487,N_1274);
and U7281 (N_7281,N_1467,N_965);
xor U7282 (N_7282,N_4410,N_3929);
or U7283 (N_7283,N_2705,N_3742);
xor U7284 (N_7284,N_481,N_2272);
nand U7285 (N_7285,N_1474,N_1538);
xor U7286 (N_7286,N_3770,N_2704);
or U7287 (N_7287,N_3634,N_4207);
xor U7288 (N_7288,N_3106,N_4674);
nor U7289 (N_7289,N_4511,N_3152);
nor U7290 (N_7290,N_174,N_1984);
xor U7291 (N_7291,N_1268,N_1455);
nand U7292 (N_7292,N_2414,N_4911);
xnor U7293 (N_7293,N_3356,N_599);
and U7294 (N_7294,N_1061,N_1251);
nand U7295 (N_7295,N_2157,N_141);
and U7296 (N_7296,N_963,N_2892);
xnor U7297 (N_7297,N_4428,N_121);
and U7298 (N_7298,N_3792,N_814);
nor U7299 (N_7299,N_4222,N_3971);
xnor U7300 (N_7300,N_1776,N_4456);
nor U7301 (N_7301,N_1986,N_3537);
nor U7302 (N_7302,N_1589,N_2653);
or U7303 (N_7303,N_1124,N_3260);
and U7304 (N_7304,N_1162,N_2840);
nor U7305 (N_7305,N_4073,N_3389);
nand U7306 (N_7306,N_3503,N_1070);
nor U7307 (N_7307,N_1904,N_2285);
or U7308 (N_7308,N_4618,N_2808);
xor U7309 (N_7309,N_1295,N_2802);
or U7310 (N_7310,N_2552,N_1980);
nor U7311 (N_7311,N_1381,N_3699);
nor U7312 (N_7312,N_677,N_3949);
nand U7313 (N_7313,N_3598,N_1264);
xnor U7314 (N_7314,N_1847,N_3501);
nand U7315 (N_7315,N_1183,N_2566);
or U7316 (N_7316,N_3586,N_3777);
nand U7317 (N_7317,N_3900,N_3555);
or U7318 (N_7318,N_1428,N_1026);
nand U7319 (N_7319,N_223,N_2136);
or U7320 (N_7320,N_2769,N_737);
nor U7321 (N_7321,N_1141,N_4920);
nor U7322 (N_7322,N_4553,N_905);
and U7323 (N_7323,N_259,N_3457);
nor U7324 (N_7324,N_1465,N_1878);
and U7325 (N_7325,N_3116,N_3322);
and U7326 (N_7326,N_4001,N_2096);
or U7327 (N_7327,N_80,N_528);
or U7328 (N_7328,N_3957,N_4114);
xnor U7329 (N_7329,N_2341,N_3382);
and U7330 (N_7330,N_263,N_2225);
xnor U7331 (N_7331,N_4453,N_727);
nor U7332 (N_7332,N_1663,N_3052);
and U7333 (N_7333,N_148,N_4980);
nor U7334 (N_7334,N_2989,N_4075);
and U7335 (N_7335,N_4170,N_1666);
and U7336 (N_7336,N_442,N_4107);
nor U7337 (N_7337,N_3205,N_1675);
and U7338 (N_7338,N_4792,N_2016);
xnor U7339 (N_7339,N_468,N_1402);
and U7340 (N_7340,N_2639,N_3212);
nor U7341 (N_7341,N_3919,N_1865);
or U7342 (N_7342,N_252,N_4781);
nand U7343 (N_7343,N_3897,N_3543);
and U7344 (N_7344,N_1955,N_1686);
nor U7345 (N_7345,N_4953,N_4815);
or U7346 (N_7346,N_3082,N_4045);
nor U7347 (N_7347,N_743,N_4596);
nor U7348 (N_7348,N_3074,N_1429);
or U7349 (N_7349,N_2113,N_2490);
and U7350 (N_7350,N_832,N_4559);
nor U7351 (N_7351,N_2550,N_195);
xor U7352 (N_7352,N_2296,N_2984);
or U7353 (N_7353,N_2977,N_4826);
and U7354 (N_7354,N_2715,N_3908);
nand U7355 (N_7355,N_4877,N_2051);
and U7356 (N_7356,N_3142,N_1544);
or U7357 (N_7357,N_4468,N_1062);
nand U7358 (N_7358,N_673,N_1928);
xnor U7359 (N_7359,N_4362,N_818);
and U7360 (N_7360,N_2437,N_3237);
nor U7361 (N_7361,N_637,N_3359);
nand U7362 (N_7362,N_3700,N_2555);
xor U7363 (N_7363,N_406,N_583);
xor U7364 (N_7364,N_2067,N_4535);
nand U7365 (N_7365,N_1753,N_3752);
or U7366 (N_7366,N_2626,N_2842);
or U7367 (N_7367,N_518,N_2875);
and U7368 (N_7368,N_2520,N_2792);
xnor U7369 (N_7369,N_2930,N_1653);
or U7370 (N_7370,N_608,N_4152);
xor U7371 (N_7371,N_3933,N_3623);
nand U7372 (N_7372,N_4969,N_596);
nand U7373 (N_7373,N_2829,N_79);
nor U7374 (N_7374,N_3323,N_2001);
nor U7375 (N_7375,N_3006,N_3714);
or U7376 (N_7376,N_12,N_1616);
nor U7377 (N_7377,N_572,N_3486);
nor U7378 (N_7378,N_1424,N_3453);
or U7379 (N_7379,N_2789,N_4305);
and U7380 (N_7380,N_3866,N_3666);
xnor U7381 (N_7381,N_3862,N_4975);
and U7382 (N_7382,N_101,N_1447);
nand U7383 (N_7383,N_284,N_1590);
xor U7384 (N_7384,N_1211,N_3398);
or U7385 (N_7385,N_2885,N_2235);
xor U7386 (N_7386,N_4359,N_1723);
nand U7387 (N_7387,N_857,N_1916);
xnor U7388 (N_7388,N_3330,N_1257);
nor U7389 (N_7389,N_2118,N_2521);
xor U7390 (N_7390,N_4422,N_3675);
and U7391 (N_7391,N_4127,N_4639);
xor U7392 (N_7392,N_748,N_2909);
nor U7393 (N_7393,N_211,N_4315);
xnor U7394 (N_7394,N_1833,N_335);
or U7395 (N_7395,N_4066,N_1097);
or U7396 (N_7396,N_3203,N_2799);
nor U7397 (N_7397,N_3413,N_1362);
or U7398 (N_7398,N_1319,N_2558);
and U7399 (N_7399,N_1910,N_296);
nor U7400 (N_7400,N_2101,N_2448);
and U7401 (N_7401,N_2599,N_4079);
nand U7402 (N_7402,N_4891,N_2633);
or U7403 (N_7403,N_2275,N_2028);
nand U7404 (N_7404,N_1639,N_873);
and U7405 (N_7405,N_2568,N_4525);
or U7406 (N_7406,N_785,N_2917);
nand U7407 (N_7407,N_3539,N_1282);
nor U7408 (N_7408,N_2959,N_4113);
nor U7409 (N_7409,N_3647,N_1012);
nand U7410 (N_7410,N_4963,N_1334);
or U7411 (N_7411,N_286,N_2462);
or U7412 (N_7412,N_2142,N_4033);
nor U7413 (N_7413,N_3005,N_2730);
xnor U7414 (N_7414,N_3610,N_2690);
or U7415 (N_7415,N_2463,N_4224);
and U7416 (N_7416,N_2765,N_4672);
nor U7417 (N_7417,N_2221,N_4375);
xor U7418 (N_7418,N_2519,N_4795);
and U7419 (N_7419,N_950,N_4447);
xor U7420 (N_7420,N_1859,N_3175);
nor U7421 (N_7421,N_3747,N_1085);
nand U7422 (N_7422,N_3065,N_509);
or U7423 (N_7423,N_774,N_2819);
nand U7424 (N_7424,N_310,N_196);
xor U7425 (N_7425,N_278,N_96);
xnor U7426 (N_7426,N_2191,N_1890);
xnor U7427 (N_7427,N_144,N_2269);
nand U7428 (N_7428,N_4937,N_987);
and U7429 (N_7429,N_4945,N_634);
and U7430 (N_7430,N_22,N_384);
nand U7431 (N_7431,N_1441,N_1919);
or U7432 (N_7432,N_565,N_3436);
or U7433 (N_7433,N_1172,N_2156);
or U7434 (N_7434,N_4614,N_3041);
nand U7435 (N_7435,N_3051,N_3189);
nor U7436 (N_7436,N_4970,N_3312);
nand U7437 (N_7437,N_3160,N_1664);
or U7438 (N_7438,N_4822,N_2206);
nor U7439 (N_7439,N_1224,N_4622);
and U7440 (N_7440,N_842,N_3444);
nand U7441 (N_7441,N_1393,N_1917);
nand U7442 (N_7442,N_3363,N_106);
or U7443 (N_7443,N_2207,N_1501);
nand U7444 (N_7444,N_3847,N_2400);
xnor U7445 (N_7445,N_3576,N_4939);
and U7446 (N_7446,N_4711,N_2241);
or U7447 (N_7447,N_2865,N_1893);
nand U7448 (N_7448,N_1766,N_1782);
nor U7449 (N_7449,N_3736,N_635);
or U7450 (N_7450,N_1248,N_214);
and U7451 (N_7451,N_1868,N_4417);
nor U7452 (N_7452,N_521,N_618);
xor U7453 (N_7453,N_3932,N_4577);
nor U7454 (N_7454,N_143,N_4624);
nor U7455 (N_7455,N_4339,N_2166);
nand U7456 (N_7456,N_398,N_3879);
and U7457 (N_7457,N_3950,N_1456);
nand U7458 (N_7458,N_4655,N_633);
xor U7459 (N_7459,N_698,N_3302);
and U7460 (N_7460,N_1578,N_1497);
and U7461 (N_7461,N_280,N_1741);
xnor U7462 (N_7462,N_2838,N_422);
nor U7463 (N_7463,N_3196,N_149);
and U7464 (N_7464,N_3183,N_1780);
nand U7465 (N_7465,N_3584,N_348);
or U7466 (N_7466,N_845,N_3625);
or U7467 (N_7467,N_3118,N_3828);
nand U7468 (N_7468,N_712,N_1609);
or U7469 (N_7469,N_1433,N_754);
nor U7470 (N_7470,N_3838,N_1886);
xnor U7471 (N_7471,N_4250,N_107);
and U7472 (N_7472,N_4982,N_1913);
nor U7473 (N_7473,N_4536,N_627);
or U7474 (N_7474,N_1048,N_2813);
and U7475 (N_7475,N_656,N_4504);
nand U7476 (N_7476,N_823,N_1423);
nor U7477 (N_7477,N_1360,N_2946);
or U7478 (N_7478,N_153,N_314);
nand U7479 (N_7479,N_3673,N_3810);
and U7480 (N_7480,N_1570,N_3375);
or U7481 (N_7481,N_3148,N_2072);
nor U7482 (N_7482,N_1836,N_4510);
and U7483 (N_7483,N_4238,N_2515);
or U7484 (N_7484,N_2718,N_1255);
xnor U7485 (N_7485,N_1028,N_186);
nor U7486 (N_7486,N_958,N_597);
xor U7487 (N_7487,N_4993,N_1914);
or U7488 (N_7488,N_3563,N_283);
or U7489 (N_7489,N_4129,N_3581);
nor U7490 (N_7490,N_2710,N_1730);
nor U7491 (N_7491,N_2711,N_3244);
nand U7492 (N_7492,N_3600,N_324);
or U7493 (N_7493,N_3380,N_979);
or U7494 (N_7494,N_4271,N_4616);
xnor U7495 (N_7495,N_2624,N_614);
or U7496 (N_7496,N_3231,N_1361);
or U7497 (N_7497,N_4574,N_2497);
nand U7498 (N_7498,N_3100,N_4719);
or U7499 (N_7499,N_4798,N_4727);
nand U7500 (N_7500,N_3603,N_374);
or U7501 (N_7501,N_2355,N_3218);
nor U7502 (N_7502,N_2156,N_2069);
nand U7503 (N_7503,N_4279,N_3478);
nand U7504 (N_7504,N_573,N_478);
and U7505 (N_7505,N_1871,N_1707);
nor U7506 (N_7506,N_1363,N_2048);
and U7507 (N_7507,N_2331,N_2611);
nor U7508 (N_7508,N_3882,N_852);
or U7509 (N_7509,N_1682,N_3915);
xnor U7510 (N_7510,N_4491,N_190);
nor U7511 (N_7511,N_3424,N_2301);
xnor U7512 (N_7512,N_1078,N_1101);
and U7513 (N_7513,N_3060,N_871);
or U7514 (N_7514,N_2177,N_4567);
or U7515 (N_7515,N_4062,N_4919);
and U7516 (N_7516,N_1245,N_3239);
nor U7517 (N_7517,N_3768,N_1518);
or U7518 (N_7518,N_3641,N_1895);
nand U7519 (N_7519,N_1561,N_397);
nand U7520 (N_7520,N_817,N_2747);
and U7521 (N_7521,N_3289,N_3337);
and U7522 (N_7522,N_4306,N_4816);
xnor U7523 (N_7523,N_1776,N_424);
or U7524 (N_7524,N_4428,N_4935);
nor U7525 (N_7525,N_2890,N_2809);
nand U7526 (N_7526,N_2116,N_3004);
xor U7527 (N_7527,N_1854,N_748);
nand U7528 (N_7528,N_2165,N_4209);
or U7529 (N_7529,N_3597,N_421);
nor U7530 (N_7530,N_4785,N_1856);
and U7531 (N_7531,N_3310,N_1146);
nand U7532 (N_7532,N_1664,N_4647);
and U7533 (N_7533,N_315,N_538);
and U7534 (N_7534,N_3298,N_3928);
or U7535 (N_7535,N_2574,N_4347);
and U7536 (N_7536,N_489,N_4051);
nand U7537 (N_7537,N_1280,N_4483);
nand U7538 (N_7538,N_799,N_683);
and U7539 (N_7539,N_4442,N_690);
and U7540 (N_7540,N_681,N_1459);
xor U7541 (N_7541,N_3111,N_2346);
xor U7542 (N_7542,N_603,N_3264);
nand U7543 (N_7543,N_2130,N_4164);
xor U7544 (N_7544,N_1908,N_2252);
or U7545 (N_7545,N_717,N_50);
nand U7546 (N_7546,N_4621,N_4892);
nand U7547 (N_7547,N_3191,N_4424);
nor U7548 (N_7548,N_1135,N_4903);
and U7549 (N_7549,N_2937,N_2692);
nand U7550 (N_7550,N_3880,N_4461);
and U7551 (N_7551,N_1599,N_1811);
or U7552 (N_7552,N_513,N_4787);
xnor U7553 (N_7553,N_3881,N_1123);
or U7554 (N_7554,N_2917,N_4658);
or U7555 (N_7555,N_4679,N_621);
or U7556 (N_7556,N_148,N_4605);
nand U7557 (N_7557,N_1748,N_2027);
and U7558 (N_7558,N_4132,N_493);
nor U7559 (N_7559,N_760,N_3263);
xnor U7560 (N_7560,N_397,N_435);
xnor U7561 (N_7561,N_4621,N_3632);
nor U7562 (N_7562,N_4644,N_673);
nand U7563 (N_7563,N_2451,N_2811);
and U7564 (N_7564,N_321,N_4513);
or U7565 (N_7565,N_617,N_2405);
xnor U7566 (N_7566,N_31,N_650);
or U7567 (N_7567,N_3186,N_3852);
xor U7568 (N_7568,N_3558,N_2364);
or U7569 (N_7569,N_1270,N_3290);
or U7570 (N_7570,N_2107,N_165);
xnor U7571 (N_7571,N_3087,N_1607);
or U7572 (N_7572,N_1603,N_1541);
xor U7573 (N_7573,N_843,N_4682);
nor U7574 (N_7574,N_707,N_1375);
or U7575 (N_7575,N_3544,N_660);
nor U7576 (N_7576,N_4423,N_3233);
or U7577 (N_7577,N_2839,N_2735);
nor U7578 (N_7578,N_3127,N_1028);
or U7579 (N_7579,N_1603,N_719);
nor U7580 (N_7580,N_3558,N_2028);
and U7581 (N_7581,N_1570,N_2638);
or U7582 (N_7582,N_618,N_3318);
nor U7583 (N_7583,N_2212,N_1226);
or U7584 (N_7584,N_4791,N_3609);
nor U7585 (N_7585,N_873,N_811);
nor U7586 (N_7586,N_3465,N_3648);
or U7587 (N_7587,N_2003,N_4319);
or U7588 (N_7588,N_4591,N_3858);
nand U7589 (N_7589,N_4908,N_3382);
and U7590 (N_7590,N_2684,N_2262);
nand U7591 (N_7591,N_2178,N_1994);
nand U7592 (N_7592,N_1651,N_1882);
or U7593 (N_7593,N_4806,N_1320);
and U7594 (N_7594,N_2444,N_3734);
or U7595 (N_7595,N_3564,N_393);
and U7596 (N_7596,N_4621,N_4268);
or U7597 (N_7597,N_786,N_2845);
or U7598 (N_7598,N_2474,N_2841);
xnor U7599 (N_7599,N_4255,N_4391);
nor U7600 (N_7600,N_3182,N_4030);
nor U7601 (N_7601,N_3124,N_4325);
nor U7602 (N_7602,N_4101,N_152);
or U7603 (N_7603,N_4880,N_3665);
and U7604 (N_7604,N_374,N_137);
and U7605 (N_7605,N_3689,N_4969);
or U7606 (N_7606,N_3241,N_732);
nor U7607 (N_7607,N_3616,N_3218);
nor U7608 (N_7608,N_4294,N_1438);
xor U7609 (N_7609,N_1211,N_2636);
nor U7610 (N_7610,N_2143,N_166);
nor U7611 (N_7611,N_3783,N_344);
nor U7612 (N_7612,N_1373,N_2432);
or U7613 (N_7613,N_1746,N_1573);
nand U7614 (N_7614,N_3503,N_2100);
nand U7615 (N_7615,N_4098,N_4748);
and U7616 (N_7616,N_771,N_2001);
nor U7617 (N_7617,N_3257,N_808);
nor U7618 (N_7618,N_529,N_640);
nand U7619 (N_7619,N_2375,N_3862);
and U7620 (N_7620,N_3921,N_2147);
or U7621 (N_7621,N_2493,N_2150);
nand U7622 (N_7622,N_4184,N_24);
xor U7623 (N_7623,N_395,N_3579);
and U7624 (N_7624,N_4763,N_4679);
nor U7625 (N_7625,N_3342,N_2935);
xor U7626 (N_7626,N_4298,N_2428);
and U7627 (N_7627,N_3407,N_491);
and U7628 (N_7628,N_4954,N_1430);
and U7629 (N_7629,N_1884,N_3974);
or U7630 (N_7630,N_2617,N_1184);
or U7631 (N_7631,N_98,N_502);
and U7632 (N_7632,N_1827,N_1364);
xor U7633 (N_7633,N_4639,N_2831);
or U7634 (N_7634,N_4539,N_8);
and U7635 (N_7635,N_930,N_3384);
nand U7636 (N_7636,N_76,N_3843);
nor U7637 (N_7637,N_319,N_749);
or U7638 (N_7638,N_4820,N_1871);
nor U7639 (N_7639,N_2408,N_2615);
and U7640 (N_7640,N_2167,N_1279);
or U7641 (N_7641,N_511,N_1026);
and U7642 (N_7642,N_4712,N_1822);
xor U7643 (N_7643,N_3735,N_3481);
or U7644 (N_7644,N_290,N_3456);
or U7645 (N_7645,N_2495,N_3019);
and U7646 (N_7646,N_45,N_3675);
nand U7647 (N_7647,N_4478,N_211);
nor U7648 (N_7648,N_700,N_3625);
or U7649 (N_7649,N_1729,N_834);
xor U7650 (N_7650,N_3781,N_3751);
nand U7651 (N_7651,N_814,N_4005);
xor U7652 (N_7652,N_4851,N_3223);
or U7653 (N_7653,N_1491,N_1886);
or U7654 (N_7654,N_2922,N_1152);
or U7655 (N_7655,N_4574,N_884);
and U7656 (N_7656,N_59,N_969);
nand U7657 (N_7657,N_4047,N_642);
nand U7658 (N_7658,N_1912,N_4037);
nor U7659 (N_7659,N_2868,N_571);
xor U7660 (N_7660,N_2227,N_1866);
and U7661 (N_7661,N_2460,N_3832);
and U7662 (N_7662,N_4068,N_1212);
or U7663 (N_7663,N_545,N_2909);
xor U7664 (N_7664,N_3380,N_4412);
or U7665 (N_7665,N_4216,N_1886);
xor U7666 (N_7666,N_638,N_4611);
or U7667 (N_7667,N_99,N_3695);
nor U7668 (N_7668,N_3521,N_2809);
and U7669 (N_7669,N_3817,N_3291);
and U7670 (N_7670,N_3052,N_4332);
or U7671 (N_7671,N_1337,N_1016);
xor U7672 (N_7672,N_4753,N_2105);
and U7673 (N_7673,N_4660,N_2910);
xnor U7674 (N_7674,N_1731,N_3966);
or U7675 (N_7675,N_4406,N_4591);
nor U7676 (N_7676,N_2126,N_1471);
or U7677 (N_7677,N_4322,N_1849);
and U7678 (N_7678,N_3247,N_4952);
or U7679 (N_7679,N_1717,N_4105);
xor U7680 (N_7680,N_4005,N_4855);
nor U7681 (N_7681,N_1221,N_2786);
nor U7682 (N_7682,N_3490,N_1189);
xor U7683 (N_7683,N_3765,N_4552);
or U7684 (N_7684,N_363,N_2997);
nor U7685 (N_7685,N_958,N_4878);
nor U7686 (N_7686,N_2296,N_3335);
xor U7687 (N_7687,N_2567,N_2508);
or U7688 (N_7688,N_1450,N_4391);
and U7689 (N_7689,N_1641,N_1097);
nor U7690 (N_7690,N_3073,N_3025);
xnor U7691 (N_7691,N_1073,N_2046);
or U7692 (N_7692,N_4990,N_2962);
xnor U7693 (N_7693,N_1154,N_1994);
xor U7694 (N_7694,N_4394,N_832);
and U7695 (N_7695,N_1094,N_2065);
nor U7696 (N_7696,N_3311,N_3684);
and U7697 (N_7697,N_3100,N_2879);
nor U7698 (N_7698,N_108,N_3721);
nand U7699 (N_7699,N_4584,N_49);
and U7700 (N_7700,N_2209,N_1743);
or U7701 (N_7701,N_4474,N_4651);
and U7702 (N_7702,N_571,N_630);
and U7703 (N_7703,N_1866,N_4116);
and U7704 (N_7704,N_3101,N_3220);
nand U7705 (N_7705,N_2020,N_4753);
nand U7706 (N_7706,N_465,N_1959);
xnor U7707 (N_7707,N_3243,N_1516);
or U7708 (N_7708,N_2662,N_576);
nor U7709 (N_7709,N_3970,N_4165);
and U7710 (N_7710,N_4964,N_4159);
or U7711 (N_7711,N_3687,N_2769);
nand U7712 (N_7712,N_2012,N_114);
and U7713 (N_7713,N_926,N_1437);
nor U7714 (N_7714,N_1172,N_4095);
and U7715 (N_7715,N_581,N_1604);
nand U7716 (N_7716,N_1639,N_121);
or U7717 (N_7717,N_1421,N_442);
nand U7718 (N_7718,N_4522,N_4856);
or U7719 (N_7719,N_1503,N_2305);
and U7720 (N_7720,N_583,N_2431);
or U7721 (N_7721,N_1957,N_1072);
nor U7722 (N_7722,N_1000,N_3887);
nor U7723 (N_7723,N_2987,N_4229);
xor U7724 (N_7724,N_464,N_4914);
xnor U7725 (N_7725,N_133,N_552);
or U7726 (N_7726,N_518,N_1071);
or U7727 (N_7727,N_3464,N_3665);
nand U7728 (N_7728,N_3476,N_1699);
nand U7729 (N_7729,N_1109,N_1875);
and U7730 (N_7730,N_2343,N_4895);
and U7731 (N_7731,N_1459,N_159);
or U7732 (N_7732,N_3243,N_4395);
and U7733 (N_7733,N_2077,N_374);
and U7734 (N_7734,N_3794,N_2779);
or U7735 (N_7735,N_3407,N_2766);
or U7736 (N_7736,N_4048,N_2957);
nand U7737 (N_7737,N_4387,N_1706);
xnor U7738 (N_7738,N_319,N_875);
nor U7739 (N_7739,N_2474,N_2623);
and U7740 (N_7740,N_279,N_3565);
and U7741 (N_7741,N_1067,N_2613);
xor U7742 (N_7742,N_735,N_2588);
nor U7743 (N_7743,N_3018,N_3725);
and U7744 (N_7744,N_3275,N_1608);
and U7745 (N_7745,N_4164,N_3776);
xor U7746 (N_7746,N_4004,N_3416);
xor U7747 (N_7747,N_2145,N_2692);
xor U7748 (N_7748,N_3609,N_918);
nor U7749 (N_7749,N_285,N_2678);
or U7750 (N_7750,N_2313,N_3846);
or U7751 (N_7751,N_4696,N_2815);
nor U7752 (N_7752,N_1055,N_2752);
or U7753 (N_7753,N_949,N_330);
and U7754 (N_7754,N_2432,N_1345);
nor U7755 (N_7755,N_2590,N_2910);
xnor U7756 (N_7756,N_4185,N_1771);
nor U7757 (N_7757,N_235,N_3233);
xnor U7758 (N_7758,N_4072,N_4377);
or U7759 (N_7759,N_322,N_2639);
xor U7760 (N_7760,N_4061,N_3195);
nand U7761 (N_7761,N_60,N_3225);
xor U7762 (N_7762,N_2466,N_2037);
xor U7763 (N_7763,N_1591,N_1317);
and U7764 (N_7764,N_3144,N_2942);
and U7765 (N_7765,N_2318,N_196);
xnor U7766 (N_7766,N_924,N_2909);
xor U7767 (N_7767,N_2084,N_3288);
and U7768 (N_7768,N_1796,N_1704);
and U7769 (N_7769,N_4095,N_1789);
and U7770 (N_7770,N_442,N_3491);
and U7771 (N_7771,N_4017,N_2128);
xnor U7772 (N_7772,N_134,N_456);
and U7773 (N_7773,N_2008,N_649);
nand U7774 (N_7774,N_1354,N_1172);
or U7775 (N_7775,N_3848,N_1900);
nor U7776 (N_7776,N_3122,N_1885);
nand U7777 (N_7777,N_3100,N_442);
xnor U7778 (N_7778,N_4041,N_4511);
nor U7779 (N_7779,N_2016,N_408);
xnor U7780 (N_7780,N_109,N_3068);
or U7781 (N_7781,N_3910,N_1036);
nand U7782 (N_7782,N_1657,N_1525);
xor U7783 (N_7783,N_4956,N_927);
or U7784 (N_7784,N_1904,N_1626);
nand U7785 (N_7785,N_1825,N_1832);
nor U7786 (N_7786,N_511,N_418);
and U7787 (N_7787,N_3860,N_1481);
nand U7788 (N_7788,N_3994,N_2813);
nand U7789 (N_7789,N_4355,N_848);
and U7790 (N_7790,N_4572,N_3264);
nor U7791 (N_7791,N_2676,N_4197);
or U7792 (N_7792,N_3568,N_1176);
xnor U7793 (N_7793,N_4387,N_1295);
xor U7794 (N_7794,N_1718,N_2633);
nand U7795 (N_7795,N_3904,N_204);
xor U7796 (N_7796,N_3936,N_2059);
nor U7797 (N_7797,N_3722,N_1914);
nand U7798 (N_7798,N_976,N_3544);
nor U7799 (N_7799,N_300,N_1743);
nor U7800 (N_7800,N_2431,N_2109);
and U7801 (N_7801,N_4300,N_4215);
xor U7802 (N_7802,N_490,N_811);
nor U7803 (N_7803,N_1249,N_102);
and U7804 (N_7804,N_84,N_1143);
nand U7805 (N_7805,N_368,N_25);
nor U7806 (N_7806,N_2711,N_2314);
nand U7807 (N_7807,N_3404,N_4486);
or U7808 (N_7808,N_2545,N_1035);
and U7809 (N_7809,N_4528,N_4133);
nand U7810 (N_7810,N_1000,N_3338);
or U7811 (N_7811,N_1432,N_1865);
and U7812 (N_7812,N_2681,N_1049);
nand U7813 (N_7813,N_4588,N_4780);
xor U7814 (N_7814,N_926,N_572);
or U7815 (N_7815,N_587,N_3631);
and U7816 (N_7816,N_2682,N_559);
nand U7817 (N_7817,N_1772,N_4575);
xor U7818 (N_7818,N_2046,N_135);
nand U7819 (N_7819,N_4365,N_1172);
xor U7820 (N_7820,N_4481,N_1308);
or U7821 (N_7821,N_4558,N_2335);
nor U7822 (N_7822,N_2678,N_325);
nor U7823 (N_7823,N_4693,N_170);
and U7824 (N_7824,N_4168,N_2135);
or U7825 (N_7825,N_422,N_4360);
or U7826 (N_7826,N_2872,N_1574);
and U7827 (N_7827,N_4820,N_4960);
nor U7828 (N_7828,N_2848,N_2429);
and U7829 (N_7829,N_4301,N_3804);
nor U7830 (N_7830,N_3427,N_4956);
and U7831 (N_7831,N_2109,N_1295);
nor U7832 (N_7832,N_4457,N_3858);
and U7833 (N_7833,N_1051,N_1400);
nand U7834 (N_7834,N_3391,N_2252);
nand U7835 (N_7835,N_3703,N_2183);
xor U7836 (N_7836,N_3342,N_886);
and U7837 (N_7837,N_4292,N_4607);
nand U7838 (N_7838,N_4012,N_3667);
and U7839 (N_7839,N_3840,N_0);
nand U7840 (N_7840,N_3144,N_3319);
or U7841 (N_7841,N_626,N_3719);
nor U7842 (N_7842,N_3884,N_1577);
nor U7843 (N_7843,N_4730,N_1392);
nor U7844 (N_7844,N_4008,N_4490);
nor U7845 (N_7845,N_4925,N_720);
xor U7846 (N_7846,N_2069,N_770);
nor U7847 (N_7847,N_4436,N_2281);
nor U7848 (N_7848,N_1556,N_553);
xor U7849 (N_7849,N_4377,N_4200);
nor U7850 (N_7850,N_1418,N_4051);
and U7851 (N_7851,N_1434,N_101);
xor U7852 (N_7852,N_3530,N_142);
or U7853 (N_7853,N_1083,N_169);
xnor U7854 (N_7854,N_4020,N_4164);
xnor U7855 (N_7855,N_4238,N_2798);
and U7856 (N_7856,N_232,N_3622);
or U7857 (N_7857,N_4327,N_2472);
or U7858 (N_7858,N_4798,N_4737);
or U7859 (N_7859,N_2590,N_3287);
nand U7860 (N_7860,N_2186,N_1727);
nor U7861 (N_7861,N_1023,N_2658);
xor U7862 (N_7862,N_2780,N_10);
nand U7863 (N_7863,N_3281,N_4749);
nor U7864 (N_7864,N_2987,N_4404);
xnor U7865 (N_7865,N_3335,N_4709);
or U7866 (N_7866,N_911,N_2713);
or U7867 (N_7867,N_4570,N_963);
or U7868 (N_7868,N_754,N_912);
and U7869 (N_7869,N_107,N_1058);
xnor U7870 (N_7870,N_3518,N_1058);
nor U7871 (N_7871,N_2226,N_3499);
nor U7872 (N_7872,N_3583,N_2958);
or U7873 (N_7873,N_3517,N_4494);
or U7874 (N_7874,N_3881,N_422);
and U7875 (N_7875,N_3333,N_1034);
or U7876 (N_7876,N_2579,N_3239);
and U7877 (N_7877,N_4798,N_2352);
or U7878 (N_7878,N_3898,N_278);
xnor U7879 (N_7879,N_3056,N_2508);
nand U7880 (N_7880,N_3567,N_3467);
nor U7881 (N_7881,N_3332,N_4588);
and U7882 (N_7882,N_3897,N_1836);
xnor U7883 (N_7883,N_441,N_3223);
nor U7884 (N_7884,N_2459,N_3885);
and U7885 (N_7885,N_3476,N_4017);
or U7886 (N_7886,N_3056,N_4662);
nor U7887 (N_7887,N_2607,N_2869);
or U7888 (N_7888,N_945,N_1552);
nor U7889 (N_7889,N_1848,N_1913);
nor U7890 (N_7890,N_2780,N_2958);
nand U7891 (N_7891,N_2833,N_3415);
nand U7892 (N_7892,N_2952,N_4828);
xnor U7893 (N_7893,N_258,N_3947);
nor U7894 (N_7894,N_3888,N_4556);
nand U7895 (N_7895,N_1399,N_3563);
and U7896 (N_7896,N_1507,N_2825);
or U7897 (N_7897,N_477,N_1409);
nand U7898 (N_7898,N_848,N_4990);
and U7899 (N_7899,N_3352,N_419);
xor U7900 (N_7900,N_4150,N_4036);
xor U7901 (N_7901,N_4763,N_2583);
or U7902 (N_7902,N_3294,N_4267);
xnor U7903 (N_7903,N_62,N_2491);
xnor U7904 (N_7904,N_394,N_1665);
and U7905 (N_7905,N_4916,N_1885);
nand U7906 (N_7906,N_4825,N_1617);
or U7907 (N_7907,N_3022,N_1922);
and U7908 (N_7908,N_906,N_1804);
xor U7909 (N_7909,N_2662,N_3134);
or U7910 (N_7910,N_1325,N_4557);
nor U7911 (N_7911,N_4029,N_2830);
xnor U7912 (N_7912,N_3595,N_4473);
or U7913 (N_7913,N_910,N_3408);
nor U7914 (N_7914,N_4381,N_9);
xor U7915 (N_7915,N_4614,N_129);
xor U7916 (N_7916,N_1678,N_1538);
nand U7917 (N_7917,N_2100,N_3861);
nor U7918 (N_7918,N_4629,N_2400);
or U7919 (N_7919,N_2222,N_3777);
nor U7920 (N_7920,N_2408,N_1347);
nand U7921 (N_7921,N_4525,N_4120);
nor U7922 (N_7922,N_361,N_3448);
xor U7923 (N_7923,N_1761,N_4311);
nand U7924 (N_7924,N_4133,N_4756);
nand U7925 (N_7925,N_179,N_1084);
nand U7926 (N_7926,N_769,N_4406);
xor U7927 (N_7927,N_4546,N_2269);
nor U7928 (N_7928,N_769,N_3618);
and U7929 (N_7929,N_4654,N_1614);
xnor U7930 (N_7930,N_1105,N_104);
nand U7931 (N_7931,N_4014,N_4789);
or U7932 (N_7932,N_2525,N_1721);
or U7933 (N_7933,N_1905,N_2648);
nor U7934 (N_7934,N_3478,N_767);
xor U7935 (N_7935,N_689,N_2497);
xor U7936 (N_7936,N_1683,N_377);
nand U7937 (N_7937,N_991,N_4461);
nand U7938 (N_7938,N_4833,N_3657);
nand U7939 (N_7939,N_4266,N_4723);
nand U7940 (N_7940,N_43,N_226);
nor U7941 (N_7941,N_4776,N_891);
or U7942 (N_7942,N_1586,N_2973);
nor U7943 (N_7943,N_4294,N_2197);
and U7944 (N_7944,N_2986,N_1179);
nand U7945 (N_7945,N_3025,N_1131);
nand U7946 (N_7946,N_1743,N_2857);
nand U7947 (N_7947,N_1185,N_3903);
nor U7948 (N_7948,N_749,N_3577);
xor U7949 (N_7949,N_4490,N_1535);
nand U7950 (N_7950,N_2367,N_3107);
or U7951 (N_7951,N_2555,N_4052);
or U7952 (N_7952,N_2013,N_3506);
nor U7953 (N_7953,N_4088,N_2079);
xnor U7954 (N_7954,N_4411,N_3334);
and U7955 (N_7955,N_7,N_1524);
nor U7956 (N_7956,N_1668,N_4967);
nand U7957 (N_7957,N_2983,N_3366);
xor U7958 (N_7958,N_1938,N_2973);
and U7959 (N_7959,N_2957,N_4945);
xnor U7960 (N_7960,N_1848,N_2254);
nand U7961 (N_7961,N_576,N_3710);
xor U7962 (N_7962,N_2091,N_2569);
or U7963 (N_7963,N_383,N_2973);
nand U7964 (N_7964,N_340,N_1542);
or U7965 (N_7965,N_3636,N_3873);
xnor U7966 (N_7966,N_576,N_4146);
xor U7967 (N_7967,N_3149,N_1420);
xor U7968 (N_7968,N_2866,N_4548);
or U7969 (N_7969,N_3276,N_3196);
nand U7970 (N_7970,N_2970,N_3855);
or U7971 (N_7971,N_3676,N_4781);
and U7972 (N_7972,N_3210,N_3172);
nand U7973 (N_7973,N_119,N_848);
and U7974 (N_7974,N_3086,N_4476);
nor U7975 (N_7975,N_2997,N_4046);
and U7976 (N_7976,N_1113,N_3330);
nor U7977 (N_7977,N_4996,N_2533);
nor U7978 (N_7978,N_3311,N_3094);
and U7979 (N_7979,N_2196,N_666);
and U7980 (N_7980,N_3027,N_4211);
nand U7981 (N_7981,N_963,N_3035);
and U7982 (N_7982,N_1997,N_3960);
xor U7983 (N_7983,N_438,N_3458);
nand U7984 (N_7984,N_1168,N_3190);
xor U7985 (N_7985,N_2155,N_2020);
nor U7986 (N_7986,N_3342,N_389);
nand U7987 (N_7987,N_3708,N_3364);
nand U7988 (N_7988,N_1980,N_196);
or U7989 (N_7989,N_3509,N_4042);
or U7990 (N_7990,N_98,N_3462);
or U7991 (N_7991,N_1574,N_3243);
and U7992 (N_7992,N_1393,N_344);
xor U7993 (N_7993,N_564,N_2178);
nand U7994 (N_7994,N_2397,N_287);
and U7995 (N_7995,N_425,N_3349);
xnor U7996 (N_7996,N_2774,N_3787);
nor U7997 (N_7997,N_2243,N_3169);
and U7998 (N_7998,N_1987,N_3543);
and U7999 (N_7999,N_4164,N_1647);
and U8000 (N_8000,N_2031,N_2723);
nand U8001 (N_8001,N_3239,N_3993);
xor U8002 (N_8002,N_2864,N_596);
xnor U8003 (N_8003,N_3093,N_3550);
xnor U8004 (N_8004,N_1157,N_4015);
xnor U8005 (N_8005,N_41,N_371);
xor U8006 (N_8006,N_4687,N_3956);
or U8007 (N_8007,N_3925,N_4950);
nor U8008 (N_8008,N_2952,N_1579);
nand U8009 (N_8009,N_529,N_3694);
xnor U8010 (N_8010,N_493,N_1893);
and U8011 (N_8011,N_729,N_4478);
nand U8012 (N_8012,N_522,N_529);
and U8013 (N_8013,N_2985,N_2684);
and U8014 (N_8014,N_3567,N_1748);
or U8015 (N_8015,N_1030,N_4551);
nor U8016 (N_8016,N_2621,N_4719);
nand U8017 (N_8017,N_4035,N_1531);
nor U8018 (N_8018,N_2253,N_3970);
or U8019 (N_8019,N_3312,N_3918);
xnor U8020 (N_8020,N_3820,N_3365);
xnor U8021 (N_8021,N_4774,N_1079);
nor U8022 (N_8022,N_4691,N_2609);
nor U8023 (N_8023,N_1190,N_2786);
nand U8024 (N_8024,N_4710,N_1289);
and U8025 (N_8025,N_2337,N_3081);
or U8026 (N_8026,N_447,N_3060);
or U8027 (N_8027,N_4406,N_705);
and U8028 (N_8028,N_2823,N_228);
nor U8029 (N_8029,N_100,N_1361);
xor U8030 (N_8030,N_231,N_3415);
xor U8031 (N_8031,N_3638,N_3677);
or U8032 (N_8032,N_2128,N_692);
or U8033 (N_8033,N_4768,N_719);
nand U8034 (N_8034,N_1315,N_2606);
nor U8035 (N_8035,N_2977,N_3070);
nor U8036 (N_8036,N_962,N_1847);
nand U8037 (N_8037,N_1179,N_131);
nand U8038 (N_8038,N_1031,N_645);
nor U8039 (N_8039,N_1571,N_1172);
or U8040 (N_8040,N_201,N_4648);
nand U8041 (N_8041,N_3469,N_2342);
nor U8042 (N_8042,N_459,N_1452);
nor U8043 (N_8043,N_686,N_2597);
xor U8044 (N_8044,N_3476,N_3637);
or U8045 (N_8045,N_4477,N_2037);
xor U8046 (N_8046,N_4676,N_3376);
nand U8047 (N_8047,N_4002,N_3829);
or U8048 (N_8048,N_1596,N_4872);
xnor U8049 (N_8049,N_1018,N_495);
and U8050 (N_8050,N_2875,N_4984);
nor U8051 (N_8051,N_2009,N_4861);
or U8052 (N_8052,N_2421,N_2070);
and U8053 (N_8053,N_2830,N_3942);
nand U8054 (N_8054,N_992,N_4293);
and U8055 (N_8055,N_2492,N_4384);
and U8056 (N_8056,N_5,N_2061);
nor U8057 (N_8057,N_1692,N_3997);
xor U8058 (N_8058,N_4402,N_2947);
nor U8059 (N_8059,N_3597,N_4067);
and U8060 (N_8060,N_2376,N_4802);
nand U8061 (N_8061,N_1162,N_352);
or U8062 (N_8062,N_1045,N_1851);
nand U8063 (N_8063,N_4896,N_2681);
nor U8064 (N_8064,N_1665,N_1752);
nor U8065 (N_8065,N_1837,N_630);
nand U8066 (N_8066,N_1523,N_2478);
xnor U8067 (N_8067,N_1542,N_1683);
or U8068 (N_8068,N_4965,N_3482);
nand U8069 (N_8069,N_4898,N_333);
xor U8070 (N_8070,N_3111,N_3360);
xnor U8071 (N_8071,N_895,N_987);
xnor U8072 (N_8072,N_4440,N_3271);
nand U8073 (N_8073,N_570,N_3089);
or U8074 (N_8074,N_3691,N_631);
nor U8075 (N_8075,N_2953,N_3118);
nor U8076 (N_8076,N_2776,N_2691);
or U8077 (N_8077,N_2445,N_4606);
or U8078 (N_8078,N_3376,N_4731);
or U8079 (N_8079,N_2578,N_956);
and U8080 (N_8080,N_4970,N_4075);
nand U8081 (N_8081,N_1241,N_4741);
xor U8082 (N_8082,N_533,N_243);
nor U8083 (N_8083,N_1741,N_984);
nor U8084 (N_8084,N_1104,N_616);
nand U8085 (N_8085,N_3152,N_4116);
and U8086 (N_8086,N_2769,N_4002);
nand U8087 (N_8087,N_1462,N_3751);
nand U8088 (N_8088,N_2919,N_587);
and U8089 (N_8089,N_3081,N_3);
nand U8090 (N_8090,N_2499,N_4888);
or U8091 (N_8091,N_3969,N_3711);
nor U8092 (N_8092,N_2075,N_3596);
and U8093 (N_8093,N_186,N_2896);
and U8094 (N_8094,N_4695,N_119);
or U8095 (N_8095,N_849,N_4666);
and U8096 (N_8096,N_2590,N_3518);
xnor U8097 (N_8097,N_3640,N_1151);
nand U8098 (N_8098,N_191,N_1249);
or U8099 (N_8099,N_4713,N_850);
nor U8100 (N_8100,N_487,N_4310);
and U8101 (N_8101,N_2618,N_207);
nand U8102 (N_8102,N_126,N_920);
xnor U8103 (N_8103,N_1473,N_4600);
and U8104 (N_8104,N_2269,N_2432);
and U8105 (N_8105,N_4925,N_1976);
and U8106 (N_8106,N_3402,N_1428);
and U8107 (N_8107,N_4629,N_1523);
and U8108 (N_8108,N_4934,N_1509);
nor U8109 (N_8109,N_2922,N_2244);
and U8110 (N_8110,N_1285,N_3748);
and U8111 (N_8111,N_4300,N_2776);
or U8112 (N_8112,N_703,N_3224);
nand U8113 (N_8113,N_1918,N_151);
nor U8114 (N_8114,N_4306,N_2896);
or U8115 (N_8115,N_3477,N_4739);
or U8116 (N_8116,N_4482,N_4227);
xnor U8117 (N_8117,N_1869,N_229);
nor U8118 (N_8118,N_1787,N_529);
xor U8119 (N_8119,N_2000,N_489);
and U8120 (N_8120,N_3305,N_4423);
nand U8121 (N_8121,N_4522,N_3311);
or U8122 (N_8122,N_3507,N_4908);
nand U8123 (N_8123,N_4201,N_2599);
nand U8124 (N_8124,N_1096,N_1961);
xnor U8125 (N_8125,N_959,N_2409);
nor U8126 (N_8126,N_2699,N_3070);
nand U8127 (N_8127,N_636,N_1556);
or U8128 (N_8128,N_2051,N_3818);
xor U8129 (N_8129,N_609,N_4892);
xnor U8130 (N_8130,N_181,N_2395);
or U8131 (N_8131,N_3213,N_4035);
or U8132 (N_8132,N_4188,N_2599);
xor U8133 (N_8133,N_2101,N_2072);
nor U8134 (N_8134,N_4413,N_1553);
xor U8135 (N_8135,N_2032,N_623);
xnor U8136 (N_8136,N_4500,N_3999);
xnor U8137 (N_8137,N_1676,N_2300);
nor U8138 (N_8138,N_2615,N_3637);
or U8139 (N_8139,N_1927,N_657);
nor U8140 (N_8140,N_306,N_3815);
xnor U8141 (N_8141,N_1526,N_4126);
nor U8142 (N_8142,N_567,N_3822);
nand U8143 (N_8143,N_3847,N_1007);
nand U8144 (N_8144,N_3925,N_1343);
and U8145 (N_8145,N_1086,N_2960);
nand U8146 (N_8146,N_1640,N_1762);
and U8147 (N_8147,N_766,N_696);
and U8148 (N_8148,N_4792,N_3182);
nor U8149 (N_8149,N_581,N_4005);
nor U8150 (N_8150,N_4196,N_1793);
and U8151 (N_8151,N_663,N_3709);
and U8152 (N_8152,N_2497,N_853);
and U8153 (N_8153,N_2547,N_2557);
or U8154 (N_8154,N_4116,N_4350);
or U8155 (N_8155,N_3364,N_3250);
xor U8156 (N_8156,N_3751,N_4334);
or U8157 (N_8157,N_827,N_4726);
xnor U8158 (N_8158,N_1069,N_3835);
and U8159 (N_8159,N_3729,N_4482);
and U8160 (N_8160,N_1458,N_1520);
and U8161 (N_8161,N_2553,N_4762);
xnor U8162 (N_8162,N_17,N_2396);
nand U8163 (N_8163,N_532,N_839);
and U8164 (N_8164,N_538,N_1538);
nor U8165 (N_8165,N_4932,N_2813);
and U8166 (N_8166,N_1939,N_4755);
or U8167 (N_8167,N_1897,N_772);
and U8168 (N_8168,N_2926,N_1117);
nand U8169 (N_8169,N_2839,N_4164);
nand U8170 (N_8170,N_808,N_4456);
xnor U8171 (N_8171,N_2258,N_2041);
and U8172 (N_8172,N_2731,N_1860);
or U8173 (N_8173,N_1544,N_3454);
and U8174 (N_8174,N_4892,N_3445);
and U8175 (N_8175,N_3409,N_3821);
and U8176 (N_8176,N_616,N_623);
or U8177 (N_8177,N_1956,N_2257);
nand U8178 (N_8178,N_907,N_1916);
nand U8179 (N_8179,N_1140,N_3788);
and U8180 (N_8180,N_1497,N_1956);
nor U8181 (N_8181,N_3713,N_2891);
and U8182 (N_8182,N_1143,N_2167);
xor U8183 (N_8183,N_2355,N_374);
or U8184 (N_8184,N_1779,N_3836);
nor U8185 (N_8185,N_4857,N_4272);
nor U8186 (N_8186,N_2315,N_2933);
xnor U8187 (N_8187,N_1860,N_2119);
nand U8188 (N_8188,N_3882,N_4567);
or U8189 (N_8189,N_2500,N_549);
and U8190 (N_8190,N_2049,N_3794);
or U8191 (N_8191,N_4211,N_2139);
nor U8192 (N_8192,N_1561,N_3101);
or U8193 (N_8193,N_3339,N_3310);
and U8194 (N_8194,N_2513,N_2805);
xor U8195 (N_8195,N_2314,N_4931);
or U8196 (N_8196,N_1192,N_2192);
or U8197 (N_8197,N_4817,N_4247);
or U8198 (N_8198,N_3627,N_3693);
and U8199 (N_8199,N_350,N_3886);
nand U8200 (N_8200,N_1198,N_2636);
and U8201 (N_8201,N_32,N_4076);
nor U8202 (N_8202,N_4935,N_2762);
xnor U8203 (N_8203,N_3683,N_288);
nand U8204 (N_8204,N_1290,N_4457);
nand U8205 (N_8205,N_116,N_3134);
xor U8206 (N_8206,N_250,N_3134);
xor U8207 (N_8207,N_2498,N_2275);
nor U8208 (N_8208,N_268,N_4628);
and U8209 (N_8209,N_1080,N_3228);
xor U8210 (N_8210,N_4873,N_1854);
nor U8211 (N_8211,N_2861,N_4821);
and U8212 (N_8212,N_1207,N_3198);
nor U8213 (N_8213,N_1508,N_3253);
xnor U8214 (N_8214,N_1445,N_484);
nor U8215 (N_8215,N_4262,N_1066);
xnor U8216 (N_8216,N_2541,N_3294);
nand U8217 (N_8217,N_4780,N_4965);
nor U8218 (N_8218,N_3822,N_677);
nand U8219 (N_8219,N_4790,N_4982);
xnor U8220 (N_8220,N_4706,N_188);
nand U8221 (N_8221,N_4527,N_2503);
xnor U8222 (N_8222,N_223,N_726);
xor U8223 (N_8223,N_876,N_2059);
nand U8224 (N_8224,N_752,N_2514);
nor U8225 (N_8225,N_2519,N_1154);
nand U8226 (N_8226,N_2969,N_4529);
xor U8227 (N_8227,N_3670,N_2737);
nor U8228 (N_8228,N_4057,N_1708);
nor U8229 (N_8229,N_3834,N_220);
or U8230 (N_8230,N_3352,N_348);
or U8231 (N_8231,N_1574,N_1651);
or U8232 (N_8232,N_18,N_1120);
and U8233 (N_8233,N_4269,N_514);
or U8234 (N_8234,N_2094,N_3395);
or U8235 (N_8235,N_1982,N_665);
nand U8236 (N_8236,N_3728,N_4797);
and U8237 (N_8237,N_4087,N_3634);
xnor U8238 (N_8238,N_2078,N_199);
xnor U8239 (N_8239,N_4866,N_666);
or U8240 (N_8240,N_3118,N_3503);
xor U8241 (N_8241,N_4490,N_767);
and U8242 (N_8242,N_772,N_4306);
xnor U8243 (N_8243,N_1479,N_1850);
and U8244 (N_8244,N_3643,N_4718);
and U8245 (N_8245,N_622,N_3412);
and U8246 (N_8246,N_3162,N_2054);
and U8247 (N_8247,N_1513,N_3972);
xnor U8248 (N_8248,N_4523,N_2908);
or U8249 (N_8249,N_3895,N_2124);
nor U8250 (N_8250,N_2453,N_1950);
xor U8251 (N_8251,N_4704,N_362);
or U8252 (N_8252,N_675,N_460);
nor U8253 (N_8253,N_540,N_2269);
xnor U8254 (N_8254,N_4430,N_1334);
xor U8255 (N_8255,N_353,N_2515);
nor U8256 (N_8256,N_2922,N_763);
and U8257 (N_8257,N_2209,N_1572);
nand U8258 (N_8258,N_2997,N_3434);
nor U8259 (N_8259,N_935,N_4821);
xnor U8260 (N_8260,N_1939,N_387);
and U8261 (N_8261,N_4131,N_2685);
nor U8262 (N_8262,N_4373,N_3281);
or U8263 (N_8263,N_315,N_260);
nor U8264 (N_8264,N_4528,N_191);
and U8265 (N_8265,N_1900,N_3528);
xor U8266 (N_8266,N_1107,N_4574);
and U8267 (N_8267,N_4471,N_3386);
and U8268 (N_8268,N_4787,N_1765);
and U8269 (N_8269,N_2046,N_1941);
and U8270 (N_8270,N_2299,N_996);
nand U8271 (N_8271,N_2254,N_1780);
nand U8272 (N_8272,N_3536,N_2070);
or U8273 (N_8273,N_1024,N_1701);
and U8274 (N_8274,N_3477,N_4178);
nor U8275 (N_8275,N_4328,N_352);
or U8276 (N_8276,N_2249,N_1823);
or U8277 (N_8277,N_1808,N_1497);
nor U8278 (N_8278,N_1440,N_1796);
nand U8279 (N_8279,N_1619,N_1761);
nor U8280 (N_8280,N_2370,N_3522);
nand U8281 (N_8281,N_2614,N_4691);
nor U8282 (N_8282,N_548,N_1046);
nand U8283 (N_8283,N_4544,N_3125);
xnor U8284 (N_8284,N_2173,N_306);
xor U8285 (N_8285,N_1065,N_3358);
or U8286 (N_8286,N_3884,N_179);
nor U8287 (N_8287,N_2199,N_2619);
xnor U8288 (N_8288,N_1295,N_394);
nor U8289 (N_8289,N_588,N_2185);
nor U8290 (N_8290,N_2946,N_1581);
and U8291 (N_8291,N_4747,N_907);
and U8292 (N_8292,N_786,N_4332);
and U8293 (N_8293,N_2390,N_2720);
xnor U8294 (N_8294,N_674,N_758);
xor U8295 (N_8295,N_63,N_27);
xnor U8296 (N_8296,N_4495,N_1216);
and U8297 (N_8297,N_4682,N_3208);
and U8298 (N_8298,N_4572,N_2596);
xnor U8299 (N_8299,N_3501,N_166);
nand U8300 (N_8300,N_4659,N_548);
xnor U8301 (N_8301,N_695,N_1478);
nor U8302 (N_8302,N_4350,N_4509);
nand U8303 (N_8303,N_3068,N_4649);
xor U8304 (N_8304,N_1920,N_4989);
nor U8305 (N_8305,N_1203,N_2804);
nor U8306 (N_8306,N_3631,N_4061);
and U8307 (N_8307,N_4656,N_2689);
xor U8308 (N_8308,N_1781,N_4557);
and U8309 (N_8309,N_2879,N_3200);
and U8310 (N_8310,N_264,N_3174);
and U8311 (N_8311,N_4659,N_4229);
nor U8312 (N_8312,N_2640,N_4799);
or U8313 (N_8313,N_3029,N_777);
xnor U8314 (N_8314,N_239,N_3610);
nor U8315 (N_8315,N_4819,N_2107);
xor U8316 (N_8316,N_3841,N_1299);
nor U8317 (N_8317,N_430,N_4637);
nand U8318 (N_8318,N_1789,N_2688);
nand U8319 (N_8319,N_2249,N_536);
nor U8320 (N_8320,N_4080,N_2498);
xnor U8321 (N_8321,N_4844,N_4496);
nor U8322 (N_8322,N_801,N_2728);
or U8323 (N_8323,N_4769,N_3362);
or U8324 (N_8324,N_3443,N_3452);
nand U8325 (N_8325,N_1836,N_2361);
or U8326 (N_8326,N_4657,N_3501);
or U8327 (N_8327,N_1544,N_359);
xnor U8328 (N_8328,N_1227,N_4671);
nor U8329 (N_8329,N_1138,N_2615);
nand U8330 (N_8330,N_3522,N_4750);
xnor U8331 (N_8331,N_243,N_4193);
nand U8332 (N_8332,N_984,N_2242);
or U8333 (N_8333,N_1228,N_1491);
and U8334 (N_8334,N_293,N_3504);
or U8335 (N_8335,N_808,N_3154);
and U8336 (N_8336,N_1398,N_1605);
or U8337 (N_8337,N_2723,N_757);
or U8338 (N_8338,N_1271,N_50);
nor U8339 (N_8339,N_3484,N_2513);
or U8340 (N_8340,N_4422,N_2821);
or U8341 (N_8341,N_1719,N_2850);
and U8342 (N_8342,N_3213,N_1405);
nor U8343 (N_8343,N_4783,N_4039);
nand U8344 (N_8344,N_3056,N_2932);
nor U8345 (N_8345,N_2757,N_1263);
nand U8346 (N_8346,N_3599,N_640);
nand U8347 (N_8347,N_2290,N_2206);
xor U8348 (N_8348,N_4470,N_2957);
nor U8349 (N_8349,N_4091,N_3349);
xnor U8350 (N_8350,N_2725,N_2200);
nand U8351 (N_8351,N_535,N_2292);
nand U8352 (N_8352,N_729,N_1466);
xnor U8353 (N_8353,N_3474,N_4076);
xnor U8354 (N_8354,N_4221,N_2171);
or U8355 (N_8355,N_4244,N_30);
or U8356 (N_8356,N_3204,N_1156);
xor U8357 (N_8357,N_4598,N_5);
nor U8358 (N_8358,N_1223,N_263);
nand U8359 (N_8359,N_2549,N_427);
xor U8360 (N_8360,N_2115,N_2301);
and U8361 (N_8361,N_3233,N_3647);
or U8362 (N_8362,N_2079,N_441);
or U8363 (N_8363,N_3271,N_2545);
and U8364 (N_8364,N_3892,N_3246);
and U8365 (N_8365,N_4739,N_3584);
or U8366 (N_8366,N_739,N_4212);
nand U8367 (N_8367,N_1488,N_4902);
or U8368 (N_8368,N_3668,N_3645);
xnor U8369 (N_8369,N_2931,N_1235);
xnor U8370 (N_8370,N_3519,N_1157);
nand U8371 (N_8371,N_3799,N_2657);
nand U8372 (N_8372,N_530,N_2949);
or U8373 (N_8373,N_4370,N_4099);
or U8374 (N_8374,N_2528,N_1903);
xor U8375 (N_8375,N_3785,N_3236);
nand U8376 (N_8376,N_421,N_2966);
nor U8377 (N_8377,N_874,N_2644);
nand U8378 (N_8378,N_1481,N_2366);
or U8379 (N_8379,N_127,N_8);
or U8380 (N_8380,N_1315,N_774);
nor U8381 (N_8381,N_4092,N_3305);
nand U8382 (N_8382,N_2869,N_2634);
nor U8383 (N_8383,N_370,N_718);
nor U8384 (N_8384,N_4702,N_938);
nor U8385 (N_8385,N_594,N_1267);
and U8386 (N_8386,N_582,N_1914);
nand U8387 (N_8387,N_1275,N_2255);
nand U8388 (N_8388,N_479,N_856);
and U8389 (N_8389,N_148,N_1223);
nand U8390 (N_8390,N_4835,N_4867);
nand U8391 (N_8391,N_4121,N_3840);
xnor U8392 (N_8392,N_2818,N_4445);
nand U8393 (N_8393,N_4229,N_334);
nor U8394 (N_8394,N_2663,N_481);
xor U8395 (N_8395,N_1653,N_4156);
and U8396 (N_8396,N_1268,N_1301);
and U8397 (N_8397,N_4593,N_458);
and U8398 (N_8398,N_2677,N_3242);
xor U8399 (N_8399,N_340,N_3820);
nor U8400 (N_8400,N_1454,N_963);
nor U8401 (N_8401,N_1288,N_1712);
and U8402 (N_8402,N_1393,N_2627);
and U8403 (N_8403,N_3862,N_4754);
nor U8404 (N_8404,N_4446,N_3324);
nor U8405 (N_8405,N_1604,N_3600);
xnor U8406 (N_8406,N_764,N_1026);
or U8407 (N_8407,N_3075,N_2199);
nor U8408 (N_8408,N_3259,N_1276);
nand U8409 (N_8409,N_1707,N_845);
xnor U8410 (N_8410,N_3537,N_856);
or U8411 (N_8411,N_3057,N_3684);
or U8412 (N_8412,N_4715,N_51);
xnor U8413 (N_8413,N_3662,N_2484);
xor U8414 (N_8414,N_3259,N_3871);
and U8415 (N_8415,N_1612,N_2680);
nand U8416 (N_8416,N_4410,N_4995);
or U8417 (N_8417,N_1415,N_2153);
and U8418 (N_8418,N_4238,N_2238);
xor U8419 (N_8419,N_878,N_219);
nand U8420 (N_8420,N_3894,N_496);
nand U8421 (N_8421,N_3773,N_722);
nand U8422 (N_8422,N_2348,N_4451);
and U8423 (N_8423,N_3430,N_4128);
xor U8424 (N_8424,N_971,N_4699);
nand U8425 (N_8425,N_1512,N_1716);
nand U8426 (N_8426,N_1760,N_1900);
and U8427 (N_8427,N_2848,N_4722);
nand U8428 (N_8428,N_4421,N_2712);
nor U8429 (N_8429,N_2235,N_3962);
or U8430 (N_8430,N_4195,N_3418);
nand U8431 (N_8431,N_4292,N_607);
xnor U8432 (N_8432,N_297,N_1335);
and U8433 (N_8433,N_2493,N_844);
xor U8434 (N_8434,N_2522,N_843);
nand U8435 (N_8435,N_4182,N_4930);
nor U8436 (N_8436,N_1398,N_4007);
or U8437 (N_8437,N_827,N_2510);
xnor U8438 (N_8438,N_1520,N_1323);
xor U8439 (N_8439,N_2003,N_596);
or U8440 (N_8440,N_3710,N_47);
xor U8441 (N_8441,N_2006,N_2040);
nand U8442 (N_8442,N_833,N_1675);
nor U8443 (N_8443,N_2922,N_537);
nor U8444 (N_8444,N_1959,N_256);
xor U8445 (N_8445,N_2527,N_731);
nand U8446 (N_8446,N_3146,N_998);
and U8447 (N_8447,N_1104,N_3295);
xor U8448 (N_8448,N_3839,N_3120);
xnor U8449 (N_8449,N_4375,N_3008);
or U8450 (N_8450,N_4175,N_3408);
and U8451 (N_8451,N_2328,N_1851);
and U8452 (N_8452,N_4961,N_2822);
xor U8453 (N_8453,N_1660,N_669);
nor U8454 (N_8454,N_1480,N_2180);
and U8455 (N_8455,N_3129,N_1122);
nor U8456 (N_8456,N_852,N_3701);
nor U8457 (N_8457,N_4143,N_4308);
and U8458 (N_8458,N_355,N_1869);
nor U8459 (N_8459,N_3374,N_957);
nor U8460 (N_8460,N_2790,N_914);
xor U8461 (N_8461,N_4164,N_1904);
xor U8462 (N_8462,N_4524,N_2362);
nor U8463 (N_8463,N_4060,N_809);
xnor U8464 (N_8464,N_24,N_3914);
xnor U8465 (N_8465,N_2720,N_1413);
xnor U8466 (N_8466,N_101,N_2180);
nand U8467 (N_8467,N_2329,N_624);
or U8468 (N_8468,N_1167,N_875);
nor U8469 (N_8469,N_2852,N_3841);
xnor U8470 (N_8470,N_572,N_2561);
xnor U8471 (N_8471,N_4266,N_558);
xor U8472 (N_8472,N_4374,N_2563);
nor U8473 (N_8473,N_186,N_3055);
xor U8474 (N_8474,N_3482,N_1981);
xor U8475 (N_8475,N_1859,N_2963);
nand U8476 (N_8476,N_4361,N_26);
nor U8477 (N_8477,N_668,N_3175);
and U8478 (N_8478,N_485,N_362);
and U8479 (N_8479,N_3146,N_2619);
nor U8480 (N_8480,N_756,N_2955);
and U8481 (N_8481,N_2580,N_2164);
nor U8482 (N_8482,N_556,N_2288);
or U8483 (N_8483,N_2329,N_460);
or U8484 (N_8484,N_4196,N_2007);
xor U8485 (N_8485,N_2175,N_3265);
and U8486 (N_8486,N_3728,N_133);
or U8487 (N_8487,N_3073,N_1026);
or U8488 (N_8488,N_4968,N_3969);
or U8489 (N_8489,N_1868,N_4985);
nand U8490 (N_8490,N_3113,N_1089);
xor U8491 (N_8491,N_1983,N_98);
nand U8492 (N_8492,N_1158,N_4255);
and U8493 (N_8493,N_2774,N_2845);
xnor U8494 (N_8494,N_3241,N_1836);
nand U8495 (N_8495,N_1706,N_311);
xnor U8496 (N_8496,N_4389,N_172);
and U8497 (N_8497,N_4648,N_3559);
nand U8498 (N_8498,N_4318,N_3682);
or U8499 (N_8499,N_4998,N_1334);
and U8500 (N_8500,N_2652,N_349);
nand U8501 (N_8501,N_1469,N_4349);
and U8502 (N_8502,N_110,N_2306);
nor U8503 (N_8503,N_1971,N_4307);
xnor U8504 (N_8504,N_2283,N_4038);
xnor U8505 (N_8505,N_4606,N_553);
and U8506 (N_8506,N_276,N_4814);
and U8507 (N_8507,N_1805,N_4192);
nor U8508 (N_8508,N_4854,N_4401);
or U8509 (N_8509,N_599,N_2159);
xnor U8510 (N_8510,N_2970,N_3469);
nand U8511 (N_8511,N_3286,N_942);
and U8512 (N_8512,N_4920,N_4614);
nand U8513 (N_8513,N_3577,N_1104);
xnor U8514 (N_8514,N_723,N_1213);
xor U8515 (N_8515,N_3073,N_2574);
nand U8516 (N_8516,N_1214,N_1699);
or U8517 (N_8517,N_1523,N_3850);
xnor U8518 (N_8518,N_4742,N_173);
and U8519 (N_8519,N_4973,N_4710);
or U8520 (N_8520,N_4733,N_3286);
nor U8521 (N_8521,N_2146,N_3763);
nor U8522 (N_8522,N_3335,N_2245);
xnor U8523 (N_8523,N_2612,N_1273);
and U8524 (N_8524,N_840,N_683);
nor U8525 (N_8525,N_698,N_4803);
or U8526 (N_8526,N_3503,N_3578);
nand U8527 (N_8527,N_3816,N_107);
and U8528 (N_8528,N_2436,N_83);
xor U8529 (N_8529,N_2541,N_1405);
nor U8530 (N_8530,N_2081,N_488);
and U8531 (N_8531,N_2012,N_1659);
xor U8532 (N_8532,N_720,N_2821);
and U8533 (N_8533,N_711,N_395);
xnor U8534 (N_8534,N_172,N_1618);
xor U8535 (N_8535,N_4702,N_3171);
nand U8536 (N_8536,N_2640,N_3377);
or U8537 (N_8537,N_1811,N_4360);
nand U8538 (N_8538,N_2903,N_3981);
xnor U8539 (N_8539,N_2874,N_1140);
xnor U8540 (N_8540,N_289,N_4580);
xnor U8541 (N_8541,N_3460,N_4188);
nand U8542 (N_8542,N_4175,N_4461);
or U8543 (N_8543,N_4290,N_873);
nand U8544 (N_8544,N_228,N_3);
nor U8545 (N_8545,N_1667,N_3280);
and U8546 (N_8546,N_221,N_1267);
or U8547 (N_8547,N_1920,N_2895);
or U8548 (N_8548,N_56,N_1211);
nand U8549 (N_8549,N_4600,N_393);
and U8550 (N_8550,N_3664,N_1223);
nor U8551 (N_8551,N_133,N_3791);
xor U8552 (N_8552,N_2930,N_1583);
or U8553 (N_8553,N_543,N_1359);
or U8554 (N_8554,N_2232,N_3091);
or U8555 (N_8555,N_4485,N_3425);
or U8556 (N_8556,N_3771,N_2148);
xnor U8557 (N_8557,N_4419,N_3801);
xor U8558 (N_8558,N_4795,N_2363);
nand U8559 (N_8559,N_2816,N_2482);
nor U8560 (N_8560,N_929,N_4187);
or U8561 (N_8561,N_1302,N_4230);
or U8562 (N_8562,N_1050,N_3593);
and U8563 (N_8563,N_2869,N_610);
and U8564 (N_8564,N_2921,N_859);
xor U8565 (N_8565,N_214,N_4228);
nor U8566 (N_8566,N_4453,N_1374);
xor U8567 (N_8567,N_3697,N_3153);
xor U8568 (N_8568,N_1771,N_1225);
or U8569 (N_8569,N_1186,N_2688);
nor U8570 (N_8570,N_1616,N_2366);
or U8571 (N_8571,N_3163,N_1743);
nand U8572 (N_8572,N_1747,N_3490);
nor U8573 (N_8573,N_4960,N_1152);
or U8574 (N_8574,N_3505,N_1991);
nor U8575 (N_8575,N_975,N_850);
or U8576 (N_8576,N_3070,N_4818);
nand U8577 (N_8577,N_2015,N_2408);
and U8578 (N_8578,N_474,N_2101);
nor U8579 (N_8579,N_4291,N_469);
nand U8580 (N_8580,N_3546,N_286);
and U8581 (N_8581,N_353,N_2153);
nand U8582 (N_8582,N_4352,N_2309);
nor U8583 (N_8583,N_2246,N_4464);
nor U8584 (N_8584,N_2316,N_3772);
or U8585 (N_8585,N_480,N_2845);
or U8586 (N_8586,N_4072,N_3018);
nand U8587 (N_8587,N_4327,N_1450);
or U8588 (N_8588,N_4154,N_1851);
or U8589 (N_8589,N_4669,N_4112);
xor U8590 (N_8590,N_3640,N_207);
nand U8591 (N_8591,N_2826,N_1261);
or U8592 (N_8592,N_570,N_2806);
nand U8593 (N_8593,N_565,N_2991);
nand U8594 (N_8594,N_3251,N_4207);
or U8595 (N_8595,N_1692,N_4784);
xor U8596 (N_8596,N_4515,N_2905);
xnor U8597 (N_8597,N_4289,N_4408);
or U8598 (N_8598,N_4433,N_965);
xnor U8599 (N_8599,N_777,N_3265);
nand U8600 (N_8600,N_3259,N_2704);
and U8601 (N_8601,N_2411,N_1855);
or U8602 (N_8602,N_4338,N_4863);
xor U8603 (N_8603,N_4100,N_3937);
and U8604 (N_8604,N_1003,N_3446);
nand U8605 (N_8605,N_757,N_3903);
nor U8606 (N_8606,N_2947,N_4618);
xor U8607 (N_8607,N_2964,N_12);
and U8608 (N_8608,N_4741,N_92);
nand U8609 (N_8609,N_3733,N_94);
nand U8610 (N_8610,N_3437,N_4866);
nand U8611 (N_8611,N_3458,N_1765);
nand U8612 (N_8612,N_328,N_3024);
nand U8613 (N_8613,N_2385,N_3268);
nor U8614 (N_8614,N_2882,N_2128);
or U8615 (N_8615,N_3070,N_656);
nor U8616 (N_8616,N_4424,N_1042);
nand U8617 (N_8617,N_3972,N_4016);
or U8618 (N_8618,N_2572,N_4251);
and U8619 (N_8619,N_2253,N_748);
and U8620 (N_8620,N_886,N_446);
nor U8621 (N_8621,N_4907,N_4070);
xnor U8622 (N_8622,N_1183,N_510);
xnor U8623 (N_8623,N_3122,N_3719);
nand U8624 (N_8624,N_1548,N_4309);
and U8625 (N_8625,N_1909,N_3501);
and U8626 (N_8626,N_1138,N_2737);
and U8627 (N_8627,N_3797,N_4443);
xnor U8628 (N_8628,N_2757,N_4571);
or U8629 (N_8629,N_1537,N_2666);
and U8630 (N_8630,N_4862,N_418);
nor U8631 (N_8631,N_2496,N_4144);
and U8632 (N_8632,N_3259,N_2345);
and U8633 (N_8633,N_2054,N_462);
xor U8634 (N_8634,N_4575,N_1156);
xor U8635 (N_8635,N_2649,N_2762);
or U8636 (N_8636,N_296,N_4597);
nor U8637 (N_8637,N_3920,N_3775);
nand U8638 (N_8638,N_2997,N_1919);
xnor U8639 (N_8639,N_768,N_2206);
nor U8640 (N_8640,N_3882,N_2090);
and U8641 (N_8641,N_4910,N_3716);
xnor U8642 (N_8642,N_4125,N_3507);
or U8643 (N_8643,N_1715,N_4693);
xor U8644 (N_8644,N_4579,N_3638);
or U8645 (N_8645,N_4425,N_3883);
nand U8646 (N_8646,N_4652,N_4280);
or U8647 (N_8647,N_3781,N_1604);
or U8648 (N_8648,N_1190,N_754);
or U8649 (N_8649,N_308,N_3100);
nand U8650 (N_8650,N_109,N_1180);
nand U8651 (N_8651,N_2493,N_4110);
and U8652 (N_8652,N_2430,N_315);
and U8653 (N_8653,N_1000,N_2533);
and U8654 (N_8654,N_2686,N_862);
xnor U8655 (N_8655,N_4513,N_3540);
xnor U8656 (N_8656,N_1007,N_1342);
and U8657 (N_8657,N_4638,N_4875);
nor U8658 (N_8658,N_4443,N_2016);
and U8659 (N_8659,N_4896,N_3857);
nor U8660 (N_8660,N_3462,N_4074);
and U8661 (N_8661,N_168,N_1988);
nor U8662 (N_8662,N_3329,N_4804);
and U8663 (N_8663,N_3101,N_1268);
or U8664 (N_8664,N_1569,N_4997);
and U8665 (N_8665,N_4736,N_69);
or U8666 (N_8666,N_781,N_2143);
nor U8667 (N_8667,N_3210,N_84);
nor U8668 (N_8668,N_1771,N_3962);
nand U8669 (N_8669,N_2443,N_2440);
or U8670 (N_8670,N_287,N_3543);
and U8671 (N_8671,N_3990,N_3386);
and U8672 (N_8672,N_1707,N_4734);
and U8673 (N_8673,N_3303,N_528);
or U8674 (N_8674,N_4285,N_587);
nand U8675 (N_8675,N_4529,N_119);
and U8676 (N_8676,N_1314,N_2668);
and U8677 (N_8677,N_767,N_2489);
and U8678 (N_8678,N_1758,N_2532);
xnor U8679 (N_8679,N_3485,N_726);
and U8680 (N_8680,N_575,N_1542);
and U8681 (N_8681,N_1287,N_2473);
xnor U8682 (N_8682,N_2594,N_4516);
and U8683 (N_8683,N_4804,N_214);
nor U8684 (N_8684,N_2840,N_1487);
or U8685 (N_8685,N_1536,N_622);
or U8686 (N_8686,N_2053,N_2285);
or U8687 (N_8687,N_2389,N_4261);
xnor U8688 (N_8688,N_2641,N_1824);
nand U8689 (N_8689,N_3207,N_199);
nor U8690 (N_8690,N_1566,N_1902);
or U8691 (N_8691,N_1415,N_2212);
and U8692 (N_8692,N_1408,N_3242);
xor U8693 (N_8693,N_1648,N_4838);
or U8694 (N_8694,N_4111,N_4459);
xnor U8695 (N_8695,N_1711,N_1843);
nor U8696 (N_8696,N_1599,N_4121);
nand U8697 (N_8697,N_4297,N_113);
xor U8698 (N_8698,N_3227,N_4028);
xor U8699 (N_8699,N_335,N_2087);
and U8700 (N_8700,N_1997,N_3334);
nand U8701 (N_8701,N_2854,N_3290);
or U8702 (N_8702,N_2275,N_2677);
nand U8703 (N_8703,N_4396,N_1044);
nand U8704 (N_8704,N_3237,N_1354);
nand U8705 (N_8705,N_858,N_2922);
or U8706 (N_8706,N_1777,N_1070);
xor U8707 (N_8707,N_928,N_2659);
or U8708 (N_8708,N_679,N_869);
or U8709 (N_8709,N_3876,N_3671);
nand U8710 (N_8710,N_2246,N_4492);
or U8711 (N_8711,N_2313,N_2274);
or U8712 (N_8712,N_389,N_895);
nor U8713 (N_8713,N_163,N_4139);
xor U8714 (N_8714,N_3765,N_4429);
and U8715 (N_8715,N_3644,N_2282);
and U8716 (N_8716,N_4915,N_3052);
and U8717 (N_8717,N_4918,N_2766);
xor U8718 (N_8718,N_2379,N_4670);
nor U8719 (N_8719,N_2702,N_3863);
and U8720 (N_8720,N_2922,N_3895);
and U8721 (N_8721,N_4612,N_2802);
and U8722 (N_8722,N_2188,N_89);
and U8723 (N_8723,N_2549,N_4954);
xor U8724 (N_8724,N_2302,N_886);
and U8725 (N_8725,N_2580,N_4640);
nor U8726 (N_8726,N_466,N_3042);
or U8727 (N_8727,N_1794,N_3841);
nand U8728 (N_8728,N_784,N_377);
nand U8729 (N_8729,N_3858,N_3133);
nand U8730 (N_8730,N_4461,N_340);
and U8731 (N_8731,N_3281,N_4682);
nand U8732 (N_8732,N_160,N_2217);
and U8733 (N_8733,N_982,N_769);
or U8734 (N_8734,N_3147,N_3750);
or U8735 (N_8735,N_767,N_2391);
nand U8736 (N_8736,N_1130,N_974);
nand U8737 (N_8737,N_563,N_1598);
xnor U8738 (N_8738,N_1728,N_3885);
nand U8739 (N_8739,N_1962,N_2372);
xor U8740 (N_8740,N_2543,N_960);
and U8741 (N_8741,N_4081,N_344);
nand U8742 (N_8742,N_3185,N_3877);
nand U8743 (N_8743,N_4223,N_3489);
xnor U8744 (N_8744,N_224,N_1300);
nand U8745 (N_8745,N_1706,N_2438);
or U8746 (N_8746,N_857,N_372);
xor U8747 (N_8747,N_971,N_25);
nand U8748 (N_8748,N_2207,N_4066);
nor U8749 (N_8749,N_4448,N_385);
nor U8750 (N_8750,N_4257,N_2308);
nand U8751 (N_8751,N_3489,N_4443);
or U8752 (N_8752,N_2,N_4153);
nand U8753 (N_8753,N_4793,N_770);
or U8754 (N_8754,N_2557,N_1059);
and U8755 (N_8755,N_2485,N_2856);
or U8756 (N_8756,N_3425,N_893);
or U8757 (N_8757,N_1309,N_2955);
or U8758 (N_8758,N_1737,N_4010);
nand U8759 (N_8759,N_1275,N_716);
and U8760 (N_8760,N_920,N_3336);
or U8761 (N_8761,N_2222,N_2101);
nor U8762 (N_8762,N_4756,N_2579);
xnor U8763 (N_8763,N_1374,N_2727);
xor U8764 (N_8764,N_4260,N_3726);
or U8765 (N_8765,N_3867,N_633);
and U8766 (N_8766,N_3426,N_2711);
nor U8767 (N_8767,N_1781,N_1744);
xor U8768 (N_8768,N_1164,N_1003);
and U8769 (N_8769,N_3892,N_1429);
nor U8770 (N_8770,N_3694,N_1701);
nor U8771 (N_8771,N_4832,N_3629);
or U8772 (N_8772,N_292,N_4872);
or U8773 (N_8773,N_2111,N_915);
xor U8774 (N_8774,N_2696,N_934);
and U8775 (N_8775,N_3148,N_4464);
and U8776 (N_8776,N_4794,N_3146);
and U8777 (N_8777,N_4232,N_2533);
and U8778 (N_8778,N_3042,N_4913);
nor U8779 (N_8779,N_1607,N_4361);
and U8780 (N_8780,N_1866,N_714);
nor U8781 (N_8781,N_2702,N_4765);
xor U8782 (N_8782,N_4258,N_1241);
nor U8783 (N_8783,N_3988,N_4616);
nand U8784 (N_8784,N_1926,N_1081);
nor U8785 (N_8785,N_4043,N_3520);
nor U8786 (N_8786,N_4204,N_82);
xor U8787 (N_8787,N_3761,N_1444);
xnor U8788 (N_8788,N_389,N_3362);
nand U8789 (N_8789,N_2638,N_3981);
or U8790 (N_8790,N_1069,N_3143);
nor U8791 (N_8791,N_4075,N_2307);
or U8792 (N_8792,N_3602,N_2921);
nor U8793 (N_8793,N_1303,N_459);
xor U8794 (N_8794,N_4541,N_2565);
nand U8795 (N_8795,N_4493,N_1506);
or U8796 (N_8796,N_4762,N_1602);
and U8797 (N_8797,N_3977,N_639);
xnor U8798 (N_8798,N_1238,N_3738);
nor U8799 (N_8799,N_3106,N_145);
nor U8800 (N_8800,N_2745,N_1987);
and U8801 (N_8801,N_4109,N_436);
and U8802 (N_8802,N_223,N_4577);
nand U8803 (N_8803,N_1235,N_413);
nor U8804 (N_8804,N_442,N_3523);
and U8805 (N_8805,N_4085,N_4442);
xor U8806 (N_8806,N_2145,N_2341);
xor U8807 (N_8807,N_1682,N_3048);
nand U8808 (N_8808,N_1286,N_319);
nand U8809 (N_8809,N_1965,N_1648);
and U8810 (N_8810,N_2509,N_3577);
nor U8811 (N_8811,N_562,N_1012);
nor U8812 (N_8812,N_1810,N_3267);
or U8813 (N_8813,N_2377,N_1628);
or U8814 (N_8814,N_4605,N_53);
nor U8815 (N_8815,N_2916,N_4587);
and U8816 (N_8816,N_4901,N_3363);
xnor U8817 (N_8817,N_438,N_3828);
or U8818 (N_8818,N_3437,N_261);
nand U8819 (N_8819,N_2825,N_1015);
and U8820 (N_8820,N_4612,N_478);
and U8821 (N_8821,N_2019,N_3868);
nor U8822 (N_8822,N_2000,N_4936);
nand U8823 (N_8823,N_2148,N_2407);
or U8824 (N_8824,N_3411,N_4574);
or U8825 (N_8825,N_2203,N_3598);
and U8826 (N_8826,N_4467,N_4336);
and U8827 (N_8827,N_4997,N_3852);
and U8828 (N_8828,N_330,N_919);
nor U8829 (N_8829,N_1233,N_4196);
and U8830 (N_8830,N_4801,N_2720);
xor U8831 (N_8831,N_1461,N_1478);
nand U8832 (N_8832,N_2240,N_2961);
xnor U8833 (N_8833,N_2136,N_997);
xnor U8834 (N_8834,N_695,N_2666);
nor U8835 (N_8835,N_1978,N_1225);
nand U8836 (N_8836,N_1638,N_2801);
nor U8837 (N_8837,N_1867,N_4874);
nand U8838 (N_8838,N_4271,N_1587);
and U8839 (N_8839,N_4271,N_4277);
nand U8840 (N_8840,N_3643,N_688);
and U8841 (N_8841,N_3257,N_2465);
xnor U8842 (N_8842,N_1474,N_347);
xor U8843 (N_8843,N_1895,N_3136);
and U8844 (N_8844,N_2827,N_1774);
and U8845 (N_8845,N_2752,N_637);
and U8846 (N_8846,N_777,N_3875);
nand U8847 (N_8847,N_3315,N_3542);
nand U8848 (N_8848,N_1954,N_478);
xor U8849 (N_8849,N_729,N_997);
nor U8850 (N_8850,N_628,N_3009);
xnor U8851 (N_8851,N_561,N_4112);
xnor U8852 (N_8852,N_690,N_3092);
xor U8853 (N_8853,N_1660,N_72);
nand U8854 (N_8854,N_2462,N_3648);
nor U8855 (N_8855,N_3751,N_2328);
or U8856 (N_8856,N_2740,N_3640);
nand U8857 (N_8857,N_4282,N_124);
xor U8858 (N_8858,N_95,N_2587);
nor U8859 (N_8859,N_4936,N_268);
and U8860 (N_8860,N_2127,N_1045);
and U8861 (N_8861,N_3781,N_2071);
nand U8862 (N_8862,N_1668,N_2682);
xor U8863 (N_8863,N_4768,N_2482);
and U8864 (N_8864,N_4205,N_125);
or U8865 (N_8865,N_2011,N_4718);
nor U8866 (N_8866,N_4362,N_1216);
or U8867 (N_8867,N_4969,N_413);
or U8868 (N_8868,N_355,N_917);
xnor U8869 (N_8869,N_2712,N_2271);
and U8870 (N_8870,N_2818,N_1829);
nor U8871 (N_8871,N_3186,N_2585);
nor U8872 (N_8872,N_2089,N_1772);
and U8873 (N_8873,N_3486,N_462);
and U8874 (N_8874,N_3970,N_2544);
nor U8875 (N_8875,N_4788,N_2132);
nand U8876 (N_8876,N_2274,N_160);
or U8877 (N_8877,N_3176,N_1324);
nor U8878 (N_8878,N_3270,N_1917);
nor U8879 (N_8879,N_990,N_1017);
nor U8880 (N_8880,N_737,N_1408);
nor U8881 (N_8881,N_761,N_4879);
nor U8882 (N_8882,N_3835,N_845);
and U8883 (N_8883,N_3539,N_4694);
xor U8884 (N_8884,N_4444,N_1804);
xnor U8885 (N_8885,N_1548,N_3566);
xnor U8886 (N_8886,N_1620,N_4122);
and U8887 (N_8887,N_3668,N_2374);
nor U8888 (N_8888,N_4048,N_745);
or U8889 (N_8889,N_4816,N_2915);
or U8890 (N_8890,N_4259,N_2536);
or U8891 (N_8891,N_3649,N_4608);
and U8892 (N_8892,N_4362,N_4685);
xor U8893 (N_8893,N_1977,N_4924);
or U8894 (N_8894,N_2979,N_4797);
and U8895 (N_8895,N_3287,N_4202);
nor U8896 (N_8896,N_1084,N_2952);
nand U8897 (N_8897,N_4795,N_4800);
xor U8898 (N_8898,N_3364,N_2991);
and U8899 (N_8899,N_1018,N_4253);
or U8900 (N_8900,N_1070,N_3607);
nand U8901 (N_8901,N_3094,N_215);
or U8902 (N_8902,N_1185,N_1426);
nor U8903 (N_8903,N_42,N_2481);
and U8904 (N_8904,N_2082,N_2595);
nor U8905 (N_8905,N_568,N_1805);
xor U8906 (N_8906,N_2373,N_4375);
and U8907 (N_8907,N_2498,N_4056);
nor U8908 (N_8908,N_46,N_4573);
or U8909 (N_8909,N_765,N_1280);
nand U8910 (N_8910,N_3793,N_1134);
nand U8911 (N_8911,N_1285,N_4533);
or U8912 (N_8912,N_840,N_715);
nand U8913 (N_8913,N_1027,N_96);
and U8914 (N_8914,N_116,N_2898);
nand U8915 (N_8915,N_2055,N_3217);
nand U8916 (N_8916,N_3709,N_4304);
and U8917 (N_8917,N_1205,N_589);
or U8918 (N_8918,N_1856,N_2472);
xnor U8919 (N_8919,N_4135,N_4537);
nor U8920 (N_8920,N_3663,N_1882);
xnor U8921 (N_8921,N_754,N_1825);
xnor U8922 (N_8922,N_3704,N_4459);
or U8923 (N_8923,N_3695,N_2931);
nor U8924 (N_8924,N_1871,N_3070);
nand U8925 (N_8925,N_553,N_2527);
nand U8926 (N_8926,N_1374,N_3223);
or U8927 (N_8927,N_617,N_1914);
and U8928 (N_8928,N_1382,N_4515);
xor U8929 (N_8929,N_322,N_4935);
and U8930 (N_8930,N_3090,N_1262);
and U8931 (N_8931,N_373,N_773);
and U8932 (N_8932,N_77,N_58);
xor U8933 (N_8933,N_3440,N_3479);
nand U8934 (N_8934,N_3038,N_3624);
nor U8935 (N_8935,N_1844,N_2849);
nor U8936 (N_8936,N_3848,N_1249);
nand U8937 (N_8937,N_1181,N_3540);
nand U8938 (N_8938,N_2557,N_1763);
and U8939 (N_8939,N_437,N_4457);
nand U8940 (N_8940,N_356,N_3950);
nand U8941 (N_8941,N_3864,N_1865);
nor U8942 (N_8942,N_2677,N_4690);
and U8943 (N_8943,N_646,N_3222);
or U8944 (N_8944,N_3768,N_2633);
or U8945 (N_8945,N_1901,N_4028);
or U8946 (N_8946,N_2002,N_2160);
xnor U8947 (N_8947,N_4910,N_70);
and U8948 (N_8948,N_4935,N_3030);
or U8949 (N_8949,N_2338,N_2105);
xnor U8950 (N_8950,N_1140,N_4896);
nor U8951 (N_8951,N_2781,N_3269);
and U8952 (N_8952,N_2410,N_4851);
nand U8953 (N_8953,N_4560,N_3542);
nor U8954 (N_8954,N_684,N_246);
nor U8955 (N_8955,N_2655,N_1869);
or U8956 (N_8956,N_3135,N_1077);
and U8957 (N_8957,N_855,N_3098);
xor U8958 (N_8958,N_2032,N_569);
nand U8959 (N_8959,N_1259,N_1228);
and U8960 (N_8960,N_3614,N_2919);
or U8961 (N_8961,N_2252,N_1701);
or U8962 (N_8962,N_3952,N_1590);
and U8963 (N_8963,N_3785,N_2764);
nand U8964 (N_8964,N_1183,N_4661);
and U8965 (N_8965,N_3429,N_3289);
or U8966 (N_8966,N_4525,N_4785);
or U8967 (N_8967,N_2406,N_1283);
nor U8968 (N_8968,N_2872,N_4387);
and U8969 (N_8969,N_1095,N_4513);
and U8970 (N_8970,N_657,N_2748);
and U8971 (N_8971,N_4078,N_967);
and U8972 (N_8972,N_3197,N_65);
or U8973 (N_8973,N_916,N_4627);
xnor U8974 (N_8974,N_4169,N_3175);
or U8975 (N_8975,N_4404,N_1537);
nor U8976 (N_8976,N_1771,N_1555);
or U8977 (N_8977,N_1811,N_3647);
nor U8978 (N_8978,N_4628,N_2939);
or U8979 (N_8979,N_2056,N_4581);
xnor U8980 (N_8980,N_48,N_3758);
xnor U8981 (N_8981,N_1515,N_212);
nor U8982 (N_8982,N_1913,N_527);
and U8983 (N_8983,N_47,N_4635);
nand U8984 (N_8984,N_2932,N_1937);
or U8985 (N_8985,N_3913,N_1626);
nand U8986 (N_8986,N_3417,N_516);
xnor U8987 (N_8987,N_243,N_4907);
xnor U8988 (N_8988,N_1464,N_2636);
nor U8989 (N_8989,N_2081,N_438);
nand U8990 (N_8990,N_3107,N_849);
or U8991 (N_8991,N_1593,N_2488);
xor U8992 (N_8992,N_1414,N_2282);
nand U8993 (N_8993,N_396,N_4668);
or U8994 (N_8994,N_949,N_219);
nor U8995 (N_8995,N_4635,N_2113);
xor U8996 (N_8996,N_1065,N_2529);
xnor U8997 (N_8997,N_3338,N_65);
and U8998 (N_8998,N_1060,N_4487);
nand U8999 (N_8999,N_1876,N_2594);
nor U9000 (N_9000,N_3893,N_1143);
nand U9001 (N_9001,N_2527,N_1848);
nor U9002 (N_9002,N_4277,N_4229);
or U9003 (N_9003,N_3597,N_1130);
xor U9004 (N_9004,N_4865,N_1017);
xnor U9005 (N_9005,N_3435,N_3851);
and U9006 (N_9006,N_395,N_4629);
or U9007 (N_9007,N_615,N_3875);
nor U9008 (N_9008,N_2464,N_2789);
xor U9009 (N_9009,N_4286,N_208);
and U9010 (N_9010,N_3300,N_1864);
nor U9011 (N_9011,N_4762,N_2129);
nand U9012 (N_9012,N_2947,N_664);
or U9013 (N_9013,N_2900,N_4254);
and U9014 (N_9014,N_1328,N_1700);
and U9015 (N_9015,N_3436,N_576);
xor U9016 (N_9016,N_3202,N_2626);
nand U9017 (N_9017,N_3400,N_2759);
or U9018 (N_9018,N_3704,N_3805);
and U9019 (N_9019,N_4863,N_1685);
or U9020 (N_9020,N_3801,N_4413);
or U9021 (N_9021,N_1779,N_497);
xor U9022 (N_9022,N_1212,N_488);
or U9023 (N_9023,N_235,N_588);
nor U9024 (N_9024,N_1935,N_4176);
nor U9025 (N_9025,N_3981,N_3596);
and U9026 (N_9026,N_229,N_3555);
or U9027 (N_9027,N_300,N_4708);
xnor U9028 (N_9028,N_430,N_4527);
nand U9029 (N_9029,N_3999,N_2524);
nand U9030 (N_9030,N_1347,N_619);
nand U9031 (N_9031,N_4509,N_43);
and U9032 (N_9032,N_3472,N_617);
nand U9033 (N_9033,N_4002,N_1748);
and U9034 (N_9034,N_937,N_3262);
nand U9035 (N_9035,N_3018,N_1065);
nand U9036 (N_9036,N_3126,N_672);
nand U9037 (N_9037,N_4970,N_1363);
xnor U9038 (N_9038,N_487,N_1006);
nand U9039 (N_9039,N_922,N_516);
and U9040 (N_9040,N_1192,N_4966);
nand U9041 (N_9041,N_4583,N_2989);
or U9042 (N_9042,N_175,N_1807);
and U9043 (N_9043,N_2083,N_856);
nand U9044 (N_9044,N_2800,N_624);
xnor U9045 (N_9045,N_3039,N_4902);
and U9046 (N_9046,N_1945,N_4799);
xnor U9047 (N_9047,N_2415,N_2318);
nor U9048 (N_9048,N_1206,N_1644);
nand U9049 (N_9049,N_637,N_4670);
xnor U9050 (N_9050,N_3882,N_33);
and U9051 (N_9051,N_2338,N_2595);
and U9052 (N_9052,N_3156,N_2529);
nand U9053 (N_9053,N_3347,N_3602);
nor U9054 (N_9054,N_3576,N_4828);
xnor U9055 (N_9055,N_3847,N_3444);
or U9056 (N_9056,N_642,N_4580);
nand U9057 (N_9057,N_852,N_383);
and U9058 (N_9058,N_3193,N_4234);
xor U9059 (N_9059,N_4652,N_4748);
xnor U9060 (N_9060,N_3146,N_2115);
nand U9061 (N_9061,N_2611,N_4510);
or U9062 (N_9062,N_2942,N_1747);
or U9063 (N_9063,N_4922,N_3123);
xnor U9064 (N_9064,N_1039,N_206);
and U9065 (N_9065,N_1101,N_1561);
and U9066 (N_9066,N_1942,N_4314);
or U9067 (N_9067,N_136,N_995);
and U9068 (N_9068,N_4449,N_3211);
nand U9069 (N_9069,N_4126,N_3730);
and U9070 (N_9070,N_1022,N_3897);
and U9071 (N_9071,N_1562,N_3674);
or U9072 (N_9072,N_204,N_2653);
and U9073 (N_9073,N_1050,N_564);
and U9074 (N_9074,N_545,N_4242);
or U9075 (N_9075,N_3,N_842);
nand U9076 (N_9076,N_789,N_1674);
xnor U9077 (N_9077,N_1776,N_1664);
nand U9078 (N_9078,N_4408,N_1058);
xor U9079 (N_9079,N_2193,N_4596);
and U9080 (N_9080,N_209,N_4697);
and U9081 (N_9081,N_3030,N_2849);
nor U9082 (N_9082,N_1207,N_1492);
nor U9083 (N_9083,N_2689,N_4389);
nand U9084 (N_9084,N_2463,N_3746);
and U9085 (N_9085,N_1710,N_3237);
or U9086 (N_9086,N_3754,N_4430);
xnor U9087 (N_9087,N_2728,N_2800);
nor U9088 (N_9088,N_4623,N_3430);
nand U9089 (N_9089,N_2753,N_1751);
or U9090 (N_9090,N_2608,N_4739);
and U9091 (N_9091,N_1380,N_1683);
or U9092 (N_9092,N_4779,N_92);
xnor U9093 (N_9093,N_4631,N_1945);
xor U9094 (N_9094,N_2738,N_1112);
xor U9095 (N_9095,N_2260,N_1885);
xor U9096 (N_9096,N_3551,N_1150);
nand U9097 (N_9097,N_4302,N_3972);
nand U9098 (N_9098,N_2990,N_2924);
nand U9099 (N_9099,N_1420,N_2040);
nand U9100 (N_9100,N_927,N_2517);
and U9101 (N_9101,N_4830,N_3148);
nand U9102 (N_9102,N_3484,N_3659);
xnor U9103 (N_9103,N_575,N_3746);
and U9104 (N_9104,N_2645,N_437);
nor U9105 (N_9105,N_2648,N_2035);
nor U9106 (N_9106,N_1273,N_1894);
nand U9107 (N_9107,N_968,N_2529);
or U9108 (N_9108,N_2301,N_3051);
and U9109 (N_9109,N_901,N_681);
xnor U9110 (N_9110,N_2852,N_2550);
and U9111 (N_9111,N_995,N_2435);
xor U9112 (N_9112,N_3466,N_4016);
and U9113 (N_9113,N_3264,N_908);
or U9114 (N_9114,N_273,N_1782);
and U9115 (N_9115,N_611,N_3086);
or U9116 (N_9116,N_108,N_3257);
and U9117 (N_9117,N_271,N_535);
xor U9118 (N_9118,N_3210,N_1041);
nor U9119 (N_9119,N_3428,N_521);
xnor U9120 (N_9120,N_2343,N_3292);
or U9121 (N_9121,N_2184,N_3862);
and U9122 (N_9122,N_4417,N_3339);
and U9123 (N_9123,N_1675,N_1218);
nor U9124 (N_9124,N_3805,N_3752);
or U9125 (N_9125,N_1460,N_208);
and U9126 (N_9126,N_4124,N_2176);
nand U9127 (N_9127,N_884,N_939);
and U9128 (N_9128,N_1628,N_4445);
xnor U9129 (N_9129,N_442,N_3875);
nor U9130 (N_9130,N_1344,N_723);
nor U9131 (N_9131,N_1746,N_454);
xor U9132 (N_9132,N_2321,N_146);
and U9133 (N_9133,N_839,N_2101);
xnor U9134 (N_9134,N_2326,N_4682);
or U9135 (N_9135,N_4762,N_2724);
xnor U9136 (N_9136,N_1946,N_2728);
nor U9137 (N_9137,N_2487,N_1113);
nor U9138 (N_9138,N_3662,N_1721);
xnor U9139 (N_9139,N_4442,N_4973);
and U9140 (N_9140,N_3150,N_4374);
xor U9141 (N_9141,N_3799,N_848);
and U9142 (N_9142,N_4574,N_3805);
nand U9143 (N_9143,N_4315,N_4250);
or U9144 (N_9144,N_3582,N_3694);
nor U9145 (N_9145,N_1173,N_4304);
nand U9146 (N_9146,N_222,N_3790);
and U9147 (N_9147,N_1862,N_493);
xnor U9148 (N_9148,N_130,N_588);
and U9149 (N_9149,N_1935,N_1579);
nor U9150 (N_9150,N_989,N_4326);
nand U9151 (N_9151,N_1296,N_1782);
nand U9152 (N_9152,N_2,N_3066);
or U9153 (N_9153,N_3289,N_3497);
and U9154 (N_9154,N_2439,N_2596);
or U9155 (N_9155,N_285,N_4725);
or U9156 (N_9156,N_3132,N_84);
or U9157 (N_9157,N_3131,N_4742);
nor U9158 (N_9158,N_4487,N_1883);
nor U9159 (N_9159,N_1022,N_567);
nand U9160 (N_9160,N_4735,N_2568);
nand U9161 (N_9161,N_3839,N_4608);
and U9162 (N_9162,N_3192,N_1180);
and U9163 (N_9163,N_3161,N_3681);
or U9164 (N_9164,N_572,N_3008);
and U9165 (N_9165,N_822,N_2619);
xnor U9166 (N_9166,N_1601,N_4411);
and U9167 (N_9167,N_1527,N_2009);
and U9168 (N_9168,N_446,N_3625);
nor U9169 (N_9169,N_621,N_4085);
and U9170 (N_9170,N_1098,N_1089);
nor U9171 (N_9171,N_363,N_3222);
nor U9172 (N_9172,N_1870,N_241);
and U9173 (N_9173,N_3274,N_1548);
nor U9174 (N_9174,N_2142,N_2497);
or U9175 (N_9175,N_4053,N_2123);
or U9176 (N_9176,N_2044,N_2221);
nor U9177 (N_9177,N_3903,N_2882);
and U9178 (N_9178,N_363,N_855);
or U9179 (N_9179,N_2764,N_1473);
xor U9180 (N_9180,N_2455,N_2176);
nand U9181 (N_9181,N_657,N_4370);
nor U9182 (N_9182,N_2896,N_4883);
nand U9183 (N_9183,N_2837,N_849);
xnor U9184 (N_9184,N_2791,N_4168);
xor U9185 (N_9185,N_2664,N_580);
nand U9186 (N_9186,N_4122,N_2647);
nor U9187 (N_9187,N_2128,N_4717);
xnor U9188 (N_9188,N_4916,N_3375);
and U9189 (N_9189,N_4299,N_4943);
or U9190 (N_9190,N_3992,N_2459);
or U9191 (N_9191,N_3252,N_1212);
xnor U9192 (N_9192,N_4989,N_3427);
and U9193 (N_9193,N_4360,N_2143);
xor U9194 (N_9194,N_4912,N_2795);
or U9195 (N_9195,N_3771,N_3548);
xor U9196 (N_9196,N_443,N_3843);
xor U9197 (N_9197,N_3509,N_1836);
xor U9198 (N_9198,N_338,N_1301);
or U9199 (N_9199,N_929,N_2255);
or U9200 (N_9200,N_3501,N_397);
nor U9201 (N_9201,N_3457,N_2498);
and U9202 (N_9202,N_4513,N_1940);
or U9203 (N_9203,N_3756,N_3644);
xor U9204 (N_9204,N_4824,N_3222);
or U9205 (N_9205,N_4715,N_3613);
and U9206 (N_9206,N_2135,N_3777);
or U9207 (N_9207,N_888,N_1957);
or U9208 (N_9208,N_2315,N_4024);
or U9209 (N_9209,N_4603,N_2840);
nor U9210 (N_9210,N_4332,N_4223);
xor U9211 (N_9211,N_3594,N_3448);
and U9212 (N_9212,N_604,N_4194);
or U9213 (N_9213,N_15,N_3023);
nand U9214 (N_9214,N_22,N_2110);
xor U9215 (N_9215,N_2576,N_4782);
xor U9216 (N_9216,N_4893,N_742);
xnor U9217 (N_9217,N_3989,N_1551);
xor U9218 (N_9218,N_3049,N_4872);
and U9219 (N_9219,N_4822,N_3505);
xnor U9220 (N_9220,N_2064,N_1773);
xor U9221 (N_9221,N_155,N_2392);
nor U9222 (N_9222,N_4781,N_38);
xor U9223 (N_9223,N_2001,N_3716);
and U9224 (N_9224,N_2987,N_1100);
or U9225 (N_9225,N_1433,N_124);
nand U9226 (N_9226,N_4475,N_3883);
xnor U9227 (N_9227,N_776,N_4448);
xor U9228 (N_9228,N_3204,N_3271);
and U9229 (N_9229,N_404,N_4139);
nor U9230 (N_9230,N_3159,N_99);
nand U9231 (N_9231,N_2952,N_3434);
xor U9232 (N_9232,N_4279,N_722);
and U9233 (N_9233,N_273,N_4886);
nand U9234 (N_9234,N_2397,N_1645);
nor U9235 (N_9235,N_1854,N_2675);
or U9236 (N_9236,N_1779,N_3468);
or U9237 (N_9237,N_2018,N_2488);
nor U9238 (N_9238,N_3472,N_3847);
nor U9239 (N_9239,N_4681,N_91);
nand U9240 (N_9240,N_1580,N_15);
nor U9241 (N_9241,N_800,N_2100);
nor U9242 (N_9242,N_3129,N_2102);
xnor U9243 (N_9243,N_3169,N_1313);
nand U9244 (N_9244,N_3178,N_744);
xor U9245 (N_9245,N_3369,N_4812);
xor U9246 (N_9246,N_3735,N_376);
nand U9247 (N_9247,N_983,N_216);
or U9248 (N_9248,N_2832,N_2559);
and U9249 (N_9249,N_2399,N_4480);
nor U9250 (N_9250,N_143,N_3643);
xor U9251 (N_9251,N_4064,N_2801);
nor U9252 (N_9252,N_1881,N_2715);
nor U9253 (N_9253,N_3756,N_4203);
nor U9254 (N_9254,N_2840,N_1481);
and U9255 (N_9255,N_2213,N_648);
nand U9256 (N_9256,N_532,N_1679);
xor U9257 (N_9257,N_352,N_830);
nand U9258 (N_9258,N_4096,N_931);
and U9259 (N_9259,N_3083,N_835);
nor U9260 (N_9260,N_3876,N_3754);
or U9261 (N_9261,N_3973,N_803);
nand U9262 (N_9262,N_4854,N_2417);
nand U9263 (N_9263,N_2100,N_310);
nand U9264 (N_9264,N_3823,N_43);
xnor U9265 (N_9265,N_1063,N_697);
xnor U9266 (N_9266,N_4385,N_1317);
and U9267 (N_9267,N_1496,N_2706);
xor U9268 (N_9268,N_1275,N_405);
or U9269 (N_9269,N_2526,N_2774);
or U9270 (N_9270,N_1380,N_2514);
and U9271 (N_9271,N_1094,N_1347);
nand U9272 (N_9272,N_4269,N_3692);
or U9273 (N_9273,N_3857,N_2986);
or U9274 (N_9274,N_202,N_1859);
nand U9275 (N_9275,N_131,N_2963);
nand U9276 (N_9276,N_2920,N_606);
nor U9277 (N_9277,N_4244,N_4501);
nand U9278 (N_9278,N_2371,N_2204);
nand U9279 (N_9279,N_51,N_3900);
or U9280 (N_9280,N_1660,N_445);
or U9281 (N_9281,N_2293,N_1472);
and U9282 (N_9282,N_3219,N_2329);
or U9283 (N_9283,N_4421,N_4580);
xnor U9284 (N_9284,N_2848,N_559);
nand U9285 (N_9285,N_1088,N_3328);
or U9286 (N_9286,N_1616,N_333);
nor U9287 (N_9287,N_2463,N_4033);
xor U9288 (N_9288,N_1085,N_2666);
nor U9289 (N_9289,N_4281,N_2711);
nand U9290 (N_9290,N_474,N_2749);
xnor U9291 (N_9291,N_3852,N_4052);
and U9292 (N_9292,N_228,N_3621);
or U9293 (N_9293,N_3386,N_2091);
or U9294 (N_9294,N_4780,N_2698);
nor U9295 (N_9295,N_2350,N_4037);
or U9296 (N_9296,N_1859,N_4894);
or U9297 (N_9297,N_1669,N_3108);
nor U9298 (N_9298,N_104,N_2739);
or U9299 (N_9299,N_3262,N_2648);
nand U9300 (N_9300,N_2341,N_4724);
xnor U9301 (N_9301,N_4437,N_4733);
and U9302 (N_9302,N_186,N_560);
xnor U9303 (N_9303,N_1852,N_377);
and U9304 (N_9304,N_763,N_3914);
xor U9305 (N_9305,N_10,N_4244);
nor U9306 (N_9306,N_2805,N_2898);
and U9307 (N_9307,N_4104,N_4645);
and U9308 (N_9308,N_3931,N_1931);
or U9309 (N_9309,N_4353,N_2563);
nor U9310 (N_9310,N_1081,N_930);
and U9311 (N_9311,N_1949,N_4123);
xor U9312 (N_9312,N_3903,N_4936);
nand U9313 (N_9313,N_4741,N_2004);
or U9314 (N_9314,N_1807,N_412);
or U9315 (N_9315,N_253,N_1388);
and U9316 (N_9316,N_4023,N_1689);
and U9317 (N_9317,N_3356,N_3206);
nor U9318 (N_9318,N_1108,N_2614);
xor U9319 (N_9319,N_2799,N_648);
nor U9320 (N_9320,N_928,N_650);
and U9321 (N_9321,N_4305,N_287);
or U9322 (N_9322,N_599,N_732);
or U9323 (N_9323,N_1829,N_4508);
nand U9324 (N_9324,N_4252,N_88);
nor U9325 (N_9325,N_1218,N_4581);
nand U9326 (N_9326,N_1196,N_441);
nor U9327 (N_9327,N_995,N_2950);
or U9328 (N_9328,N_242,N_3959);
xnor U9329 (N_9329,N_731,N_1117);
or U9330 (N_9330,N_3526,N_3778);
nor U9331 (N_9331,N_2926,N_4540);
xnor U9332 (N_9332,N_2333,N_4360);
xor U9333 (N_9333,N_2287,N_586);
and U9334 (N_9334,N_1773,N_3757);
nor U9335 (N_9335,N_3069,N_4254);
nand U9336 (N_9336,N_214,N_2067);
nor U9337 (N_9337,N_2816,N_647);
nor U9338 (N_9338,N_4269,N_3411);
and U9339 (N_9339,N_118,N_4139);
xnor U9340 (N_9340,N_3663,N_2673);
nand U9341 (N_9341,N_4889,N_994);
nor U9342 (N_9342,N_4165,N_56);
or U9343 (N_9343,N_1662,N_3656);
nand U9344 (N_9344,N_3783,N_714);
xor U9345 (N_9345,N_4151,N_4250);
nor U9346 (N_9346,N_3359,N_1309);
nand U9347 (N_9347,N_2264,N_3762);
and U9348 (N_9348,N_3075,N_1348);
nor U9349 (N_9349,N_1068,N_3358);
xor U9350 (N_9350,N_4006,N_960);
or U9351 (N_9351,N_883,N_4);
or U9352 (N_9352,N_718,N_2719);
nand U9353 (N_9353,N_1058,N_2468);
and U9354 (N_9354,N_2444,N_4097);
nand U9355 (N_9355,N_4562,N_2518);
nand U9356 (N_9356,N_3080,N_264);
nand U9357 (N_9357,N_1954,N_3619);
or U9358 (N_9358,N_2367,N_3472);
xnor U9359 (N_9359,N_1546,N_2353);
nor U9360 (N_9360,N_3948,N_3453);
and U9361 (N_9361,N_1307,N_4142);
nand U9362 (N_9362,N_502,N_1684);
and U9363 (N_9363,N_4063,N_2886);
or U9364 (N_9364,N_2174,N_802);
nor U9365 (N_9365,N_475,N_1950);
nand U9366 (N_9366,N_624,N_834);
nor U9367 (N_9367,N_3154,N_155);
nor U9368 (N_9368,N_1365,N_555);
or U9369 (N_9369,N_1560,N_4310);
or U9370 (N_9370,N_3208,N_4599);
and U9371 (N_9371,N_2141,N_2008);
nor U9372 (N_9372,N_4331,N_1030);
nor U9373 (N_9373,N_4688,N_2133);
or U9374 (N_9374,N_4493,N_4888);
xor U9375 (N_9375,N_2204,N_3829);
nor U9376 (N_9376,N_152,N_3651);
nor U9377 (N_9377,N_4859,N_4753);
nand U9378 (N_9378,N_3178,N_2637);
nor U9379 (N_9379,N_1289,N_485);
nor U9380 (N_9380,N_3023,N_1717);
or U9381 (N_9381,N_2343,N_1203);
xor U9382 (N_9382,N_1873,N_4612);
nor U9383 (N_9383,N_4178,N_4775);
and U9384 (N_9384,N_1271,N_4086);
or U9385 (N_9385,N_2132,N_255);
nor U9386 (N_9386,N_3465,N_629);
xnor U9387 (N_9387,N_3009,N_2660);
nor U9388 (N_9388,N_3021,N_235);
nor U9389 (N_9389,N_2243,N_2121);
xor U9390 (N_9390,N_2038,N_2230);
or U9391 (N_9391,N_1422,N_2599);
nand U9392 (N_9392,N_1996,N_2171);
xnor U9393 (N_9393,N_155,N_1230);
xnor U9394 (N_9394,N_1464,N_3480);
nand U9395 (N_9395,N_4521,N_2288);
nor U9396 (N_9396,N_4561,N_3452);
and U9397 (N_9397,N_4841,N_528);
or U9398 (N_9398,N_4816,N_1325);
nor U9399 (N_9399,N_4924,N_3280);
and U9400 (N_9400,N_1609,N_3732);
nand U9401 (N_9401,N_4383,N_159);
xor U9402 (N_9402,N_780,N_2284);
nor U9403 (N_9403,N_1854,N_2796);
and U9404 (N_9404,N_22,N_875);
or U9405 (N_9405,N_4068,N_196);
xor U9406 (N_9406,N_3722,N_160);
nor U9407 (N_9407,N_1671,N_4112);
or U9408 (N_9408,N_2676,N_2921);
or U9409 (N_9409,N_1449,N_4751);
or U9410 (N_9410,N_2670,N_1777);
nor U9411 (N_9411,N_1950,N_2684);
xor U9412 (N_9412,N_1427,N_4504);
nor U9413 (N_9413,N_425,N_2536);
xnor U9414 (N_9414,N_217,N_3916);
and U9415 (N_9415,N_1916,N_522);
and U9416 (N_9416,N_2602,N_1098);
xnor U9417 (N_9417,N_4169,N_2315);
or U9418 (N_9418,N_4178,N_1126);
nor U9419 (N_9419,N_4182,N_1652);
nor U9420 (N_9420,N_4517,N_2016);
xnor U9421 (N_9421,N_2709,N_4892);
nor U9422 (N_9422,N_3163,N_742);
or U9423 (N_9423,N_4977,N_836);
and U9424 (N_9424,N_4163,N_4057);
nor U9425 (N_9425,N_4054,N_4474);
xnor U9426 (N_9426,N_4761,N_232);
or U9427 (N_9427,N_4099,N_4663);
and U9428 (N_9428,N_4025,N_4775);
nand U9429 (N_9429,N_1478,N_4949);
and U9430 (N_9430,N_3357,N_2316);
and U9431 (N_9431,N_2107,N_444);
nor U9432 (N_9432,N_695,N_4398);
nor U9433 (N_9433,N_2431,N_1799);
nand U9434 (N_9434,N_3107,N_3327);
xnor U9435 (N_9435,N_4999,N_2220);
nor U9436 (N_9436,N_1893,N_1302);
nand U9437 (N_9437,N_4374,N_1630);
nand U9438 (N_9438,N_4083,N_910);
xnor U9439 (N_9439,N_4592,N_181);
xnor U9440 (N_9440,N_4714,N_4871);
xor U9441 (N_9441,N_80,N_1313);
xnor U9442 (N_9442,N_3290,N_959);
nor U9443 (N_9443,N_2165,N_2114);
nor U9444 (N_9444,N_722,N_3826);
or U9445 (N_9445,N_4476,N_4581);
nor U9446 (N_9446,N_724,N_3984);
nand U9447 (N_9447,N_3657,N_391);
nor U9448 (N_9448,N_2764,N_1697);
and U9449 (N_9449,N_2260,N_566);
or U9450 (N_9450,N_4210,N_3660);
xnor U9451 (N_9451,N_2104,N_1793);
or U9452 (N_9452,N_2475,N_868);
nand U9453 (N_9453,N_1641,N_111);
nand U9454 (N_9454,N_4035,N_2415);
and U9455 (N_9455,N_4205,N_2669);
nor U9456 (N_9456,N_1881,N_939);
nor U9457 (N_9457,N_4264,N_3268);
and U9458 (N_9458,N_4166,N_888);
or U9459 (N_9459,N_2812,N_2024);
xnor U9460 (N_9460,N_3862,N_2114);
nand U9461 (N_9461,N_4582,N_4194);
and U9462 (N_9462,N_73,N_3138);
or U9463 (N_9463,N_660,N_3242);
and U9464 (N_9464,N_4381,N_4215);
or U9465 (N_9465,N_56,N_182);
nor U9466 (N_9466,N_3073,N_3567);
or U9467 (N_9467,N_286,N_3541);
nor U9468 (N_9468,N_3938,N_2320);
xor U9469 (N_9469,N_4632,N_1531);
nand U9470 (N_9470,N_4558,N_2018);
nand U9471 (N_9471,N_4761,N_1803);
nand U9472 (N_9472,N_4797,N_569);
and U9473 (N_9473,N_3533,N_1348);
nand U9474 (N_9474,N_1701,N_3732);
nor U9475 (N_9475,N_4354,N_3177);
or U9476 (N_9476,N_4520,N_3504);
and U9477 (N_9477,N_826,N_4478);
nor U9478 (N_9478,N_2353,N_706);
nand U9479 (N_9479,N_4377,N_3920);
nor U9480 (N_9480,N_2772,N_190);
nor U9481 (N_9481,N_4792,N_2426);
nand U9482 (N_9482,N_3758,N_1915);
or U9483 (N_9483,N_3502,N_2562);
or U9484 (N_9484,N_77,N_2435);
nor U9485 (N_9485,N_1737,N_1247);
xor U9486 (N_9486,N_3754,N_3673);
nand U9487 (N_9487,N_1581,N_2461);
xnor U9488 (N_9488,N_1039,N_290);
xor U9489 (N_9489,N_3676,N_3034);
nand U9490 (N_9490,N_4097,N_4931);
or U9491 (N_9491,N_2146,N_1298);
and U9492 (N_9492,N_381,N_1444);
nor U9493 (N_9493,N_3180,N_1467);
nand U9494 (N_9494,N_79,N_3818);
nand U9495 (N_9495,N_3370,N_3483);
nor U9496 (N_9496,N_2966,N_174);
or U9497 (N_9497,N_921,N_4155);
or U9498 (N_9498,N_4240,N_14);
or U9499 (N_9499,N_2848,N_876);
or U9500 (N_9500,N_1280,N_2031);
nand U9501 (N_9501,N_4835,N_4027);
or U9502 (N_9502,N_138,N_784);
and U9503 (N_9503,N_589,N_1533);
nand U9504 (N_9504,N_2299,N_4803);
nand U9505 (N_9505,N_2540,N_1972);
xnor U9506 (N_9506,N_1151,N_4696);
or U9507 (N_9507,N_3013,N_1536);
or U9508 (N_9508,N_3193,N_1736);
nand U9509 (N_9509,N_3454,N_2184);
xnor U9510 (N_9510,N_1505,N_159);
xnor U9511 (N_9511,N_2744,N_4970);
nand U9512 (N_9512,N_4968,N_2280);
and U9513 (N_9513,N_969,N_2198);
or U9514 (N_9514,N_1783,N_1101);
or U9515 (N_9515,N_3627,N_1720);
nand U9516 (N_9516,N_1527,N_1591);
xor U9517 (N_9517,N_2547,N_1463);
or U9518 (N_9518,N_4221,N_2502);
or U9519 (N_9519,N_3669,N_2633);
or U9520 (N_9520,N_3044,N_513);
and U9521 (N_9521,N_4278,N_3245);
nor U9522 (N_9522,N_3027,N_3230);
or U9523 (N_9523,N_4090,N_2514);
nor U9524 (N_9524,N_1365,N_1489);
xor U9525 (N_9525,N_3384,N_848);
and U9526 (N_9526,N_2468,N_3123);
xnor U9527 (N_9527,N_1253,N_780);
nor U9528 (N_9528,N_1111,N_1607);
xor U9529 (N_9529,N_3661,N_1424);
and U9530 (N_9530,N_4797,N_2954);
and U9531 (N_9531,N_2084,N_2976);
and U9532 (N_9532,N_804,N_1197);
and U9533 (N_9533,N_1307,N_4989);
or U9534 (N_9534,N_4952,N_3957);
and U9535 (N_9535,N_2323,N_2414);
nor U9536 (N_9536,N_1908,N_3414);
nand U9537 (N_9537,N_4792,N_4067);
xor U9538 (N_9538,N_434,N_697);
xnor U9539 (N_9539,N_337,N_2051);
or U9540 (N_9540,N_2549,N_4392);
nor U9541 (N_9541,N_1680,N_2855);
and U9542 (N_9542,N_254,N_4359);
nand U9543 (N_9543,N_3259,N_4370);
nand U9544 (N_9544,N_2334,N_3538);
nor U9545 (N_9545,N_2297,N_2726);
and U9546 (N_9546,N_3327,N_3712);
or U9547 (N_9547,N_933,N_4625);
or U9548 (N_9548,N_4631,N_1093);
and U9549 (N_9549,N_1583,N_2249);
nor U9550 (N_9550,N_906,N_4338);
or U9551 (N_9551,N_1529,N_1851);
xor U9552 (N_9552,N_2025,N_1174);
and U9553 (N_9553,N_3254,N_4604);
or U9554 (N_9554,N_4441,N_701);
and U9555 (N_9555,N_2112,N_1829);
nand U9556 (N_9556,N_4136,N_4115);
or U9557 (N_9557,N_1953,N_2427);
xor U9558 (N_9558,N_1412,N_4694);
nor U9559 (N_9559,N_3082,N_4727);
nand U9560 (N_9560,N_928,N_4153);
or U9561 (N_9561,N_4738,N_2183);
or U9562 (N_9562,N_2347,N_3621);
and U9563 (N_9563,N_1674,N_83);
and U9564 (N_9564,N_3282,N_189);
or U9565 (N_9565,N_1045,N_1565);
nand U9566 (N_9566,N_225,N_876);
xor U9567 (N_9567,N_1926,N_13);
nor U9568 (N_9568,N_2132,N_77);
and U9569 (N_9569,N_416,N_4720);
nand U9570 (N_9570,N_878,N_236);
nand U9571 (N_9571,N_2352,N_3463);
or U9572 (N_9572,N_3481,N_3826);
nor U9573 (N_9573,N_4930,N_4009);
nor U9574 (N_9574,N_4049,N_475);
nor U9575 (N_9575,N_2017,N_272);
and U9576 (N_9576,N_3,N_4134);
xnor U9577 (N_9577,N_724,N_2544);
nor U9578 (N_9578,N_4863,N_3278);
and U9579 (N_9579,N_869,N_4293);
nor U9580 (N_9580,N_2355,N_3665);
nor U9581 (N_9581,N_2203,N_3876);
or U9582 (N_9582,N_2659,N_1984);
xor U9583 (N_9583,N_3541,N_733);
xor U9584 (N_9584,N_4727,N_3145);
nand U9585 (N_9585,N_1126,N_2267);
or U9586 (N_9586,N_2833,N_3613);
nand U9587 (N_9587,N_4306,N_4552);
and U9588 (N_9588,N_1702,N_4089);
and U9589 (N_9589,N_561,N_2416);
or U9590 (N_9590,N_496,N_3849);
and U9591 (N_9591,N_1621,N_1063);
or U9592 (N_9592,N_4950,N_2159);
nand U9593 (N_9593,N_4766,N_781);
xnor U9594 (N_9594,N_4453,N_2323);
nor U9595 (N_9595,N_2155,N_2754);
nand U9596 (N_9596,N_4333,N_33);
nand U9597 (N_9597,N_1995,N_4353);
or U9598 (N_9598,N_3057,N_3844);
nor U9599 (N_9599,N_2457,N_3326);
nand U9600 (N_9600,N_2799,N_3534);
and U9601 (N_9601,N_4544,N_2189);
or U9602 (N_9602,N_2711,N_3556);
and U9603 (N_9603,N_484,N_1309);
nand U9604 (N_9604,N_2328,N_3155);
and U9605 (N_9605,N_264,N_2712);
nor U9606 (N_9606,N_1247,N_3398);
or U9607 (N_9607,N_138,N_438);
nand U9608 (N_9608,N_2286,N_3159);
xnor U9609 (N_9609,N_1393,N_4492);
nand U9610 (N_9610,N_86,N_4782);
nand U9611 (N_9611,N_4549,N_1829);
nand U9612 (N_9612,N_4882,N_3297);
nand U9613 (N_9613,N_3027,N_340);
nand U9614 (N_9614,N_2774,N_3633);
or U9615 (N_9615,N_2965,N_2590);
xnor U9616 (N_9616,N_4238,N_2743);
nand U9617 (N_9617,N_4211,N_589);
and U9618 (N_9618,N_4516,N_4713);
nor U9619 (N_9619,N_2689,N_4144);
xor U9620 (N_9620,N_1597,N_1792);
xor U9621 (N_9621,N_1262,N_4872);
xnor U9622 (N_9622,N_359,N_1006);
xor U9623 (N_9623,N_4700,N_1485);
xor U9624 (N_9624,N_3592,N_2573);
and U9625 (N_9625,N_2196,N_3425);
xor U9626 (N_9626,N_4251,N_524);
xor U9627 (N_9627,N_2586,N_1819);
nor U9628 (N_9628,N_1416,N_438);
nor U9629 (N_9629,N_1487,N_2144);
xnor U9630 (N_9630,N_1623,N_4940);
and U9631 (N_9631,N_2839,N_2157);
or U9632 (N_9632,N_3840,N_1337);
nand U9633 (N_9633,N_393,N_3857);
or U9634 (N_9634,N_4502,N_3969);
and U9635 (N_9635,N_1812,N_1068);
and U9636 (N_9636,N_42,N_3175);
and U9637 (N_9637,N_504,N_4573);
xnor U9638 (N_9638,N_4785,N_267);
nor U9639 (N_9639,N_1134,N_2080);
nand U9640 (N_9640,N_1257,N_3973);
or U9641 (N_9641,N_802,N_4250);
nand U9642 (N_9642,N_141,N_3613);
and U9643 (N_9643,N_4290,N_3011);
nand U9644 (N_9644,N_1217,N_52);
nor U9645 (N_9645,N_2408,N_1587);
xnor U9646 (N_9646,N_1460,N_4005);
xor U9647 (N_9647,N_761,N_2371);
nand U9648 (N_9648,N_3273,N_2289);
xor U9649 (N_9649,N_167,N_1904);
and U9650 (N_9650,N_3122,N_3615);
or U9651 (N_9651,N_3938,N_4921);
and U9652 (N_9652,N_1860,N_803);
nand U9653 (N_9653,N_2625,N_2906);
nand U9654 (N_9654,N_2695,N_2560);
or U9655 (N_9655,N_4433,N_3367);
xnor U9656 (N_9656,N_4188,N_3302);
and U9657 (N_9657,N_2104,N_2210);
xor U9658 (N_9658,N_904,N_408);
or U9659 (N_9659,N_1184,N_1674);
or U9660 (N_9660,N_4225,N_3001);
or U9661 (N_9661,N_4302,N_4678);
xor U9662 (N_9662,N_686,N_4293);
xor U9663 (N_9663,N_3149,N_4604);
xnor U9664 (N_9664,N_1086,N_4442);
or U9665 (N_9665,N_384,N_4555);
nor U9666 (N_9666,N_1502,N_4067);
or U9667 (N_9667,N_2787,N_2822);
and U9668 (N_9668,N_2715,N_2336);
or U9669 (N_9669,N_4591,N_1344);
nor U9670 (N_9670,N_3058,N_1149);
and U9671 (N_9671,N_2176,N_5);
xor U9672 (N_9672,N_1599,N_444);
and U9673 (N_9673,N_2569,N_3825);
or U9674 (N_9674,N_3540,N_3841);
or U9675 (N_9675,N_3343,N_3142);
nor U9676 (N_9676,N_2234,N_2582);
nand U9677 (N_9677,N_4520,N_2980);
and U9678 (N_9678,N_4895,N_3246);
and U9679 (N_9679,N_1665,N_2494);
xor U9680 (N_9680,N_1787,N_1050);
nand U9681 (N_9681,N_1782,N_1166);
nor U9682 (N_9682,N_2799,N_2535);
nor U9683 (N_9683,N_3549,N_4276);
nand U9684 (N_9684,N_4305,N_4413);
nand U9685 (N_9685,N_4521,N_2029);
or U9686 (N_9686,N_1434,N_1570);
or U9687 (N_9687,N_2053,N_4104);
or U9688 (N_9688,N_1797,N_4038);
nand U9689 (N_9689,N_842,N_2872);
xor U9690 (N_9690,N_2204,N_4266);
or U9691 (N_9691,N_3007,N_825);
xnor U9692 (N_9692,N_2949,N_2683);
nand U9693 (N_9693,N_4515,N_3442);
or U9694 (N_9694,N_4126,N_1058);
xnor U9695 (N_9695,N_1097,N_731);
or U9696 (N_9696,N_2352,N_4512);
or U9697 (N_9697,N_2260,N_4818);
and U9698 (N_9698,N_3486,N_1454);
and U9699 (N_9699,N_3996,N_3131);
xnor U9700 (N_9700,N_4173,N_2589);
nor U9701 (N_9701,N_980,N_2754);
and U9702 (N_9702,N_3491,N_3600);
and U9703 (N_9703,N_3806,N_4155);
xnor U9704 (N_9704,N_2692,N_2947);
nand U9705 (N_9705,N_4655,N_4289);
nand U9706 (N_9706,N_2005,N_319);
or U9707 (N_9707,N_3774,N_1450);
nor U9708 (N_9708,N_3915,N_3254);
xnor U9709 (N_9709,N_784,N_2450);
xnor U9710 (N_9710,N_4198,N_4844);
and U9711 (N_9711,N_3161,N_4172);
xor U9712 (N_9712,N_4783,N_1563);
xor U9713 (N_9713,N_715,N_894);
and U9714 (N_9714,N_3904,N_3694);
nand U9715 (N_9715,N_2068,N_1540);
nand U9716 (N_9716,N_3654,N_3482);
nor U9717 (N_9717,N_2871,N_4545);
nor U9718 (N_9718,N_947,N_2090);
nor U9719 (N_9719,N_2822,N_2278);
nand U9720 (N_9720,N_3299,N_2412);
and U9721 (N_9721,N_3477,N_4196);
or U9722 (N_9722,N_1352,N_1795);
and U9723 (N_9723,N_560,N_1696);
nand U9724 (N_9724,N_2644,N_1861);
or U9725 (N_9725,N_2149,N_406);
xor U9726 (N_9726,N_434,N_2314);
nand U9727 (N_9727,N_4709,N_2914);
nor U9728 (N_9728,N_4441,N_891);
and U9729 (N_9729,N_1113,N_3798);
xnor U9730 (N_9730,N_1698,N_1940);
xnor U9731 (N_9731,N_4772,N_3290);
nand U9732 (N_9732,N_891,N_3359);
nand U9733 (N_9733,N_4119,N_751);
or U9734 (N_9734,N_2052,N_940);
nor U9735 (N_9735,N_2090,N_4190);
nor U9736 (N_9736,N_541,N_3929);
or U9737 (N_9737,N_4318,N_4740);
nand U9738 (N_9738,N_2852,N_271);
nand U9739 (N_9739,N_654,N_3974);
and U9740 (N_9740,N_1160,N_2162);
or U9741 (N_9741,N_4461,N_2549);
or U9742 (N_9742,N_2091,N_3383);
or U9743 (N_9743,N_1037,N_3649);
or U9744 (N_9744,N_2978,N_373);
or U9745 (N_9745,N_4542,N_3624);
nor U9746 (N_9746,N_861,N_2445);
nor U9747 (N_9747,N_198,N_3267);
nor U9748 (N_9748,N_2939,N_1288);
or U9749 (N_9749,N_3454,N_1229);
xor U9750 (N_9750,N_2110,N_598);
and U9751 (N_9751,N_3596,N_4237);
and U9752 (N_9752,N_3265,N_3477);
nor U9753 (N_9753,N_2335,N_207);
or U9754 (N_9754,N_4147,N_3136);
or U9755 (N_9755,N_1226,N_4606);
xnor U9756 (N_9756,N_2057,N_1430);
or U9757 (N_9757,N_4093,N_4595);
nand U9758 (N_9758,N_1017,N_248);
xnor U9759 (N_9759,N_1360,N_1560);
xor U9760 (N_9760,N_3420,N_748);
xor U9761 (N_9761,N_4981,N_1753);
nor U9762 (N_9762,N_1272,N_3665);
and U9763 (N_9763,N_2894,N_3803);
and U9764 (N_9764,N_1155,N_2395);
or U9765 (N_9765,N_4561,N_4853);
or U9766 (N_9766,N_4032,N_599);
nor U9767 (N_9767,N_4073,N_123);
nand U9768 (N_9768,N_3164,N_3753);
or U9769 (N_9769,N_1585,N_3217);
and U9770 (N_9770,N_1385,N_4769);
and U9771 (N_9771,N_4972,N_4673);
and U9772 (N_9772,N_3721,N_3243);
and U9773 (N_9773,N_2753,N_3983);
nor U9774 (N_9774,N_946,N_4857);
nor U9775 (N_9775,N_3605,N_2457);
or U9776 (N_9776,N_4794,N_2627);
nor U9777 (N_9777,N_2298,N_1185);
or U9778 (N_9778,N_2848,N_2802);
and U9779 (N_9779,N_1747,N_4471);
xor U9780 (N_9780,N_910,N_2342);
or U9781 (N_9781,N_2413,N_609);
nor U9782 (N_9782,N_835,N_2810);
or U9783 (N_9783,N_3701,N_168);
nor U9784 (N_9784,N_2903,N_433);
nand U9785 (N_9785,N_1265,N_3207);
nor U9786 (N_9786,N_548,N_2969);
nand U9787 (N_9787,N_4909,N_4828);
nand U9788 (N_9788,N_2837,N_2128);
or U9789 (N_9789,N_3619,N_1474);
nand U9790 (N_9790,N_691,N_1613);
nor U9791 (N_9791,N_268,N_92);
xnor U9792 (N_9792,N_3738,N_3999);
nand U9793 (N_9793,N_4713,N_1147);
or U9794 (N_9794,N_276,N_200);
or U9795 (N_9795,N_306,N_3976);
nand U9796 (N_9796,N_841,N_370);
xor U9797 (N_9797,N_1203,N_2580);
or U9798 (N_9798,N_1712,N_698);
and U9799 (N_9799,N_3316,N_1812);
nand U9800 (N_9800,N_2731,N_4366);
nand U9801 (N_9801,N_4094,N_3381);
xnor U9802 (N_9802,N_2162,N_3555);
nor U9803 (N_9803,N_444,N_3149);
nor U9804 (N_9804,N_496,N_2107);
and U9805 (N_9805,N_4550,N_4610);
and U9806 (N_9806,N_4815,N_3021);
nand U9807 (N_9807,N_3764,N_2133);
or U9808 (N_9808,N_1307,N_3028);
nor U9809 (N_9809,N_1150,N_935);
or U9810 (N_9810,N_4364,N_316);
xor U9811 (N_9811,N_184,N_3687);
nand U9812 (N_9812,N_1766,N_3877);
xnor U9813 (N_9813,N_4828,N_872);
and U9814 (N_9814,N_2603,N_968);
xor U9815 (N_9815,N_2681,N_2081);
nor U9816 (N_9816,N_1944,N_103);
nand U9817 (N_9817,N_4888,N_4771);
nor U9818 (N_9818,N_3266,N_442);
nand U9819 (N_9819,N_2768,N_4249);
nor U9820 (N_9820,N_401,N_2875);
xor U9821 (N_9821,N_1973,N_2682);
nor U9822 (N_9822,N_3951,N_4127);
and U9823 (N_9823,N_881,N_953);
or U9824 (N_9824,N_3104,N_1324);
xor U9825 (N_9825,N_1992,N_3963);
xor U9826 (N_9826,N_4336,N_2796);
xnor U9827 (N_9827,N_1917,N_1100);
or U9828 (N_9828,N_4925,N_58);
nor U9829 (N_9829,N_2909,N_4192);
xnor U9830 (N_9830,N_3045,N_4530);
xnor U9831 (N_9831,N_4455,N_4160);
xnor U9832 (N_9832,N_2798,N_471);
or U9833 (N_9833,N_2122,N_907);
xor U9834 (N_9834,N_4109,N_4395);
or U9835 (N_9835,N_1325,N_3390);
or U9836 (N_9836,N_4877,N_2725);
or U9837 (N_9837,N_3988,N_960);
nor U9838 (N_9838,N_1808,N_251);
and U9839 (N_9839,N_1242,N_4796);
and U9840 (N_9840,N_1880,N_4779);
nor U9841 (N_9841,N_809,N_3987);
nand U9842 (N_9842,N_3309,N_1435);
xnor U9843 (N_9843,N_2158,N_2162);
or U9844 (N_9844,N_2665,N_1448);
nand U9845 (N_9845,N_1354,N_3317);
nand U9846 (N_9846,N_3349,N_2647);
or U9847 (N_9847,N_2480,N_4980);
or U9848 (N_9848,N_4048,N_2724);
nand U9849 (N_9849,N_4480,N_1314);
xor U9850 (N_9850,N_3268,N_897);
nor U9851 (N_9851,N_2066,N_1091);
nor U9852 (N_9852,N_2010,N_2236);
and U9853 (N_9853,N_1887,N_882);
xnor U9854 (N_9854,N_740,N_3945);
or U9855 (N_9855,N_4182,N_2543);
nor U9856 (N_9856,N_1552,N_619);
xor U9857 (N_9857,N_2942,N_754);
nand U9858 (N_9858,N_1474,N_4905);
and U9859 (N_9859,N_4626,N_603);
or U9860 (N_9860,N_780,N_2948);
or U9861 (N_9861,N_1506,N_3984);
xor U9862 (N_9862,N_2332,N_547);
and U9863 (N_9863,N_471,N_4073);
nand U9864 (N_9864,N_3130,N_1481);
and U9865 (N_9865,N_2119,N_2160);
nand U9866 (N_9866,N_2839,N_4984);
or U9867 (N_9867,N_4404,N_1683);
and U9868 (N_9868,N_4051,N_1670);
xor U9869 (N_9869,N_840,N_1339);
and U9870 (N_9870,N_233,N_3825);
nand U9871 (N_9871,N_4893,N_706);
nor U9872 (N_9872,N_2110,N_4159);
and U9873 (N_9873,N_115,N_1288);
nor U9874 (N_9874,N_4381,N_166);
and U9875 (N_9875,N_1409,N_1054);
or U9876 (N_9876,N_720,N_3750);
and U9877 (N_9877,N_505,N_2066);
nor U9878 (N_9878,N_4424,N_3246);
xnor U9879 (N_9879,N_2105,N_3602);
or U9880 (N_9880,N_270,N_4775);
or U9881 (N_9881,N_989,N_4159);
or U9882 (N_9882,N_1880,N_3553);
and U9883 (N_9883,N_349,N_4608);
and U9884 (N_9884,N_3583,N_4559);
or U9885 (N_9885,N_1380,N_3611);
and U9886 (N_9886,N_336,N_2401);
or U9887 (N_9887,N_4773,N_4176);
or U9888 (N_9888,N_1918,N_3101);
nand U9889 (N_9889,N_1005,N_4599);
or U9890 (N_9890,N_4811,N_1395);
xor U9891 (N_9891,N_2532,N_3122);
nand U9892 (N_9892,N_709,N_286);
nor U9893 (N_9893,N_2219,N_1294);
or U9894 (N_9894,N_1873,N_1566);
or U9895 (N_9895,N_560,N_3956);
or U9896 (N_9896,N_2782,N_2332);
or U9897 (N_9897,N_3750,N_2603);
nand U9898 (N_9898,N_1370,N_120);
and U9899 (N_9899,N_3924,N_965);
or U9900 (N_9900,N_4691,N_4317);
nor U9901 (N_9901,N_129,N_3753);
nand U9902 (N_9902,N_3872,N_439);
or U9903 (N_9903,N_3329,N_2287);
xnor U9904 (N_9904,N_1976,N_914);
nand U9905 (N_9905,N_1069,N_2445);
or U9906 (N_9906,N_3447,N_4867);
or U9907 (N_9907,N_1506,N_1002);
nor U9908 (N_9908,N_2731,N_2988);
and U9909 (N_9909,N_2576,N_4409);
nand U9910 (N_9910,N_3435,N_1503);
xnor U9911 (N_9911,N_1823,N_3786);
nand U9912 (N_9912,N_1568,N_1166);
xnor U9913 (N_9913,N_2878,N_332);
nor U9914 (N_9914,N_1979,N_3714);
or U9915 (N_9915,N_3537,N_4295);
nor U9916 (N_9916,N_653,N_3649);
nand U9917 (N_9917,N_1732,N_1852);
nand U9918 (N_9918,N_502,N_3719);
xnor U9919 (N_9919,N_1770,N_4945);
and U9920 (N_9920,N_146,N_1986);
or U9921 (N_9921,N_501,N_4756);
and U9922 (N_9922,N_3075,N_2757);
or U9923 (N_9923,N_203,N_4103);
xor U9924 (N_9924,N_1185,N_3160);
xnor U9925 (N_9925,N_2921,N_3338);
xnor U9926 (N_9926,N_3263,N_1221);
nor U9927 (N_9927,N_1599,N_3267);
nor U9928 (N_9928,N_2892,N_4920);
nand U9929 (N_9929,N_4123,N_2309);
or U9930 (N_9930,N_4806,N_247);
or U9931 (N_9931,N_404,N_1245);
xnor U9932 (N_9932,N_1554,N_4600);
nor U9933 (N_9933,N_3681,N_4525);
or U9934 (N_9934,N_2426,N_2291);
nand U9935 (N_9935,N_3053,N_1951);
or U9936 (N_9936,N_2869,N_1966);
nor U9937 (N_9937,N_2437,N_444);
nor U9938 (N_9938,N_539,N_1228);
nor U9939 (N_9939,N_4795,N_1433);
nand U9940 (N_9940,N_3286,N_1234);
xnor U9941 (N_9941,N_2609,N_1751);
or U9942 (N_9942,N_309,N_2422);
or U9943 (N_9943,N_4416,N_2086);
nand U9944 (N_9944,N_2439,N_3773);
and U9945 (N_9945,N_4020,N_1341);
and U9946 (N_9946,N_3950,N_479);
or U9947 (N_9947,N_2457,N_602);
xor U9948 (N_9948,N_234,N_3507);
nor U9949 (N_9949,N_2981,N_3369);
nor U9950 (N_9950,N_88,N_2873);
and U9951 (N_9951,N_1739,N_4361);
nor U9952 (N_9952,N_1263,N_3211);
nand U9953 (N_9953,N_244,N_2377);
nand U9954 (N_9954,N_1689,N_4988);
xor U9955 (N_9955,N_1066,N_2074);
or U9956 (N_9956,N_3405,N_3090);
nor U9957 (N_9957,N_837,N_605);
and U9958 (N_9958,N_239,N_1880);
and U9959 (N_9959,N_2111,N_1605);
or U9960 (N_9960,N_1551,N_4133);
nand U9961 (N_9961,N_4187,N_2766);
or U9962 (N_9962,N_3387,N_2359);
or U9963 (N_9963,N_1649,N_2523);
nand U9964 (N_9964,N_4074,N_506);
nand U9965 (N_9965,N_3344,N_807);
nand U9966 (N_9966,N_4991,N_4877);
and U9967 (N_9967,N_2760,N_4945);
nor U9968 (N_9968,N_332,N_4122);
xnor U9969 (N_9969,N_3899,N_1683);
and U9970 (N_9970,N_621,N_3596);
and U9971 (N_9971,N_4823,N_4305);
or U9972 (N_9972,N_1201,N_3994);
xor U9973 (N_9973,N_732,N_3419);
nor U9974 (N_9974,N_361,N_2153);
or U9975 (N_9975,N_1209,N_4354);
nor U9976 (N_9976,N_2927,N_2398);
and U9977 (N_9977,N_4369,N_2825);
nor U9978 (N_9978,N_742,N_2831);
xnor U9979 (N_9979,N_3986,N_2813);
nand U9980 (N_9980,N_1194,N_116);
nand U9981 (N_9981,N_2659,N_2671);
nand U9982 (N_9982,N_4091,N_4182);
nor U9983 (N_9983,N_2898,N_338);
or U9984 (N_9984,N_4408,N_1677);
and U9985 (N_9985,N_2212,N_586);
or U9986 (N_9986,N_4503,N_4406);
and U9987 (N_9987,N_4524,N_3476);
xor U9988 (N_9988,N_1789,N_2291);
or U9989 (N_9989,N_254,N_2106);
nand U9990 (N_9990,N_4191,N_517);
nor U9991 (N_9991,N_4212,N_4502);
nor U9992 (N_9992,N_238,N_3756);
nor U9993 (N_9993,N_792,N_538);
and U9994 (N_9994,N_3574,N_3685);
and U9995 (N_9995,N_1337,N_4547);
and U9996 (N_9996,N_604,N_4461);
xnor U9997 (N_9997,N_2211,N_1000);
xnor U9998 (N_9998,N_3074,N_3458);
or U9999 (N_9999,N_3938,N_3246);
or UO_0 (O_0,N_8352,N_9805);
and UO_1 (O_1,N_7170,N_6275);
and UO_2 (O_2,N_5040,N_5500);
and UO_3 (O_3,N_8520,N_6028);
nand UO_4 (O_4,N_5906,N_8297);
nor UO_5 (O_5,N_7984,N_8149);
or UO_6 (O_6,N_9317,N_9026);
nor UO_7 (O_7,N_7761,N_9719);
or UO_8 (O_8,N_5059,N_6791);
nand UO_9 (O_9,N_7405,N_7790);
nand UO_10 (O_10,N_8560,N_7271);
and UO_11 (O_11,N_6861,N_5402);
and UO_12 (O_12,N_8620,N_7769);
nor UO_13 (O_13,N_9773,N_5569);
xnor UO_14 (O_14,N_7758,N_8534);
or UO_15 (O_15,N_7477,N_6950);
nand UO_16 (O_16,N_8389,N_8776);
and UO_17 (O_17,N_8715,N_6941);
nand UO_18 (O_18,N_8484,N_5955);
and UO_19 (O_19,N_5921,N_7787);
or UO_20 (O_20,N_9668,N_6592);
nand UO_21 (O_21,N_7284,N_6528);
and UO_22 (O_22,N_5101,N_6197);
nand UO_23 (O_23,N_7993,N_8807);
xnor UO_24 (O_24,N_7060,N_9769);
or UO_25 (O_25,N_8953,N_8618);
or UO_26 (O_26,N_6897,N_7868);
and UO_27 (O_27,N_6702,N_8878);
nand UO_28 (O_28,N_9945,N_7998);
and UO_29 (O_29,N_7607,N_9464);
nor UO_30 (O_30,N_6271,N_8429);
or UO_31 (O_31,N_9758,N_5738);
nor UO_32 (O_32,N_9639,N_7456);
and UO_33 (O_33,N_6734,N_7280);
and UO_34 (O_34,N_5084,N_9264);
nand UO_35 (O_35,N_5240,N_8080);
and UO_36 (O_36,N_9901,N_6938);
nand UO_37 (O_37,N_7818,N_8480);
nor UO_38 (O_38,N_5705,N_8663);
or UO_39 (O_39,N_7473,N_9042);
and UO_40 (O_40,N_6221,N_8517);
nand UO_41 (O_41,N_8460,N_7000);
nand UO_42 (O_42,N_8222,N_9586);
nand UO_43 (O_43,N_7378,N_9897);
nand UO_44 (O_44,N_9247,N_5011);
nor UO_45 (O_45,N_7235,N_6649);
xor UO_46 (O_46,N_9416,N_6581);
or UO_47 (O_47,N_6916,N_9242);
and UO_48 (O_48,N_9049,N_9456);
and UO_49 (O_49,N_5282,N_5048);
xor UO_50 (O_50,N_7823,N_9116);
xnor UO_51 (O_51,N_9617,N_7691);
xor UO_52 (O_52,N_9628,N_5155);
nand UO_53 (O_53,N_9585,N_9334);
and UO_54 (O_54,N_9894,N_5853);
nand UO_55 (O_55,N_8224,N_8511);
nand UO_56 (O_56,N_9877,N_6127);
nand UO_57 (O_57,N_8627,N_9854);
nand UO_58 (O_58,N_9052,N_5281);
nand UO_59 (O_59,N_8059,N_7562);
or UO_60 (O_60,N_9269,N_5226);
and UO_61 (O_61,N_5415,N_8179);
or UO_62 (O_62,N_5800,N_8158);
or UO_63 (O_63,N_7080,N_8516);
nor UO_64 (O_64,N_6119,N_6519);
or UO_65 (O_65,N_5945,N_9944);
xnor UO_66 (O_66,N_9006,N_5857);
and UO_67 (O_67,N_5518,N_8995);
or UO_68 (O_68,N_7865,N_5844);
nor UO_69 (O_69,N_5532,N_5615);
xnor UO_70 (O_70,N_7229,N_8634);
nand UO_71 (O_71,N_7142,N_9397);
nand UO_72 (O_72,N_6866,N_9868);
xor UO_73 (O_73,N_9305,N_9352);
or UO_74 (O_74,N_9365,N_9906);
nand UO_75 (O_75,N_5045,N_6740);
xnor UO_76 (O_76,N_6996,N_6888);
xor UO_77 (O_77,N_7652,N_5138);
nor UO_78 (O_78,N_7774,N_5637);
nand UO_79 (O_79,N_6325,N_6005);
or UO_80 (O_80,N_9498,N_7891);
nand UO_81 (O_81,N_7920,N_8499);
nor UO_82 (O_82,N_6909,N_5624);
nor UO_83 (O_83,N_8886,N_5535);
nand UO_84 (O_84,N_7665,N_6282);
xnor UO_85 (O_85,N_9749,N_7007);
nand UO_86 (O_86,N_9132,N_6405);
nand UO_87 (O_87,N_6783,N_8016);
or UO_88 (O_88,N_5204,N_5956);
or UO_89 (O_89,N_5678,N_7533);
xor UO_90 (O_90,N_9367,N_6367);
nor UO_91 (O_91,N_7075,N_6685);
and UO_92 (O_92,N_5515,N_7388);
nand UO_93 (O_93,N_5758,N_8225);
xnor UO_94 (O_94,N_6394,N_8428);
or UO_95 (O_95,N_8207,N_8607);
and UO_96 (O_96,N_7732,N_7307);
or UO_97 (O_97,N_8265,N_6008);
nand UO_98 (O_98,N_8215,N_6710);
xor UO_99 (O_99,N_5483,N_8183);
and UO_100 (O_100,N_5237,N_5176);
nand UO_101 (O_101,N_8083,N_5530);
or UO_102 (O_102,N_5905,N_5296);
nand UO_103 (O_103,N_5193,N_9165);
nor UO_104 (O_104,N_8862,N_7929);
xnor UO_105 (O_105,N_6817,N_8261);
nand UO_106 (O_106,N_7598,N_6446);
or UO_107 (O_107,N_7945,N_6992);
nor UO_108 (O_108,N_7150,N_8603);
or UO_109 (O_109,N_7146,N_8186);
nand UO_110 (O_110,N_8625,N_7961);
nand UO_111 (O_111,N_9442,N_5696);
xnor UO_112 (O_112,N_8580,N_9429);
and UO_113 (O_113,N_8213,N_8685);
or UO_114 (O_114,N_9568,N_7420);
or UO_115 (O_115,N_9815,N_9070);
xor UO_116 (O_116,N_5953,N_9085);
and UO_117 (O_117,N_9060,N_7649);
and UO_118 (O_118,N_9777,N_6037);
and UO_119 (O_119,N_5198,N_6536);
xor UO_120 (O_120,N_8888,N_8329);
nor UO_121 (O_121,N_9139,N_6788);
and UO_122 (O_122,N_9827,N_7659);
xor UO_123 (O_123,N_7343,N_6889);
and UO_124 (O_124,N_8024,N_7933);
nand UO_125 (O_125,N_9772,N_5936);
and UO_126 (O_126,N_6562,N_5592);
nor UO_127 (O_127,N_8843,N_6054);
nor UO_128 (O_128,N_9348,N_9936);
xor UO_129 (O_129,N_8420,N_5900);
nand UO_130 (O_130,N_9105,N_8815);
or UO_131 (O_131,N_5109,N_5050);
xnor UO_132 (O_132,N_5815,N_9304);
xor UO_133 (O_133,N_6160,N_5767);
and UO_134 (O_134,N_5926,N_9086);
xnor UO_135 (O_135,N_7954,N_5812);
nand UO_136 (O_136,N_6263,N_5725);
nand UO_137 (O_137,N_6653,N_5374);
and UO_138 (O_138,N_6088,N_6566);
nand UO_139 (O_139,N_5931,N_8101);
and UO_140 (O_140,N_9420,N_9008);
xor UO_141 (O_141,N_8626,N_5520);
xnor UO_142 (O_142,N_5852,N_7496);
nand UO_143 (O_143,N_9205,N_6970);
or UO_144 (O_144,N_6356,N_8962);
and UO_145 (O_145,N_8773,N_7034);
xnor UO_146 (O_146,N_5586,N_8863);
or UO_147 (O_147,N_5103,N_6552);
or UO_148 (O_148,N_7553,N_8029);
xnor UO_149 (O_149,N_7497,N_8279);
and UO_150 (O_150,N_6333,N_9275);
nor UO_151 (O_151,N_6695,N_5310);
and UO_152 (O_152,N_5173,N_6871);
nor UO_153 (O_153,N_6245,N_6485);
or UO_154 (O_154,N_5080,N_8076);
nor UO_155 (O_155,N_9422,N_6214);
nor UO_156 (O_156,N_9297,N_7101);
xor UO_157 (O_157,N_9798,N_7148);
and UO_158 (O_158,N_9226,N_5121);
nor UO_159 (O_159,N_5078,N_8590);
nand UO_160 (O_160,N_9185,N_5925);
nor UO_161 (O_161,N_5143,N_5470);
nor UO_162 (O_162,N_9545,N_7371);
and UO_163 (O_163,N_6757,N_8513);
or UO_164 (O_164,N_6322,N_7895);
or UO_165 (O_165,N_6065,N_6687);
and UO_166 (O_166,N_6308,N_7119);
and UO_167 (O_167,N_7091,N_8543);
nor UO_168 (O_168,N_6414,N_5312);
nand UO_169 (O_169,N_5213,N_8880);
xor UO_170 (O_170,N_6135,N_7297);
and UO_171 (O_171,N_6951,N_7898);
nand UO_172 (O_172,N_5039,N_6587);
or UO_173 (O_173,N_7046,N_6772);
or UO_174 (O_174,N_5370,N_6668);
nand UO_175 (O_175,N_5062,N_5511);
nor UO_176 (O_176,N_6365,N_7834);
nor UO_177 (O_177,N_7588,N_6440);
nand UO_178 (O_178,N_8541,N_9030);
nand UO_179 (O_179,N_9931,N_6490);
or UO_180 (O_180,N_5102,N_7301);
or UO_181 (O_181,N_6638,N_6211);
nor UO_182 (O_182,N_6639,N_9579);
nor UO_183 (O_183,N_8791,N_6976);
nor UO_184 (O_184,N_6052,N_6505);
nor UO_185 (O_185,N_7773,N_5318);
and UO_186 (O_186,N_7727,N_7937);
and UO_187 (O_187,N_9742,N_6634);
or UO_188 (O_188,N_9665,N_9021);
and UO_189 (O_189,N_6074,N_5054);
nand UO_190 (O_190,N_7058,N_6995);
nor UO_191 (O_191,N_5351,N_9296);
nand UO_192 (O_192,N_9908,N_5779);
nand UO_193 (O_193,N_8596,N_9222);
and UO_194 (O_194,N_9005,N_6882);
nor UO_195 (O_195,N_9731,N_5091);
and UO_196 (O_196,N_9299,N_8599);
and UO_197 (O_197,N_5403,N_6336);
xnor UO_198 (O_198,N_7521,N_7454);
xor UO_199 (O_199,N_8072,N_5810);
nand UO_200 (O_200,N_6790,N_8097);
nor UO_201 (O_201,N_7824,N_9607);
and UO_202 (O_202,N_6429,N_8964);
nor UO_203 (O_203,N_5396,N_6610);
or UO_204 (O_204,N_8890,N_7706);
nor UO_205 (O_205,N_6132,N_5283);
and UO_206 (O_206,N_8570,N_8347);
nand UO_207 (O_207,N_6180,N_7755);
nor UO_208 (O_208,N_9075,N_6988);
or UO_209 (O_209,N_8573,N_8496);
nor UO_210 (O_210,N_9612,N_9698);
nand UO_211 (O_211,N_7213,N_7780);
and UO_212 (O_212,N_6669,N_5807);
nand UO_213 (O_213,N_5846,N_6942);
nand UO_214 (O_214,N_5073,N_8483);
and UO_215 (O_215,N_5836,N_9146);
and UO_216 (O_216,N_7527,N_9715);
and UO_217 (O_217,N_9909,N_8788);
xnor UO_218 (O_218,N_7279,N_6241);
nand UO_219 (O_219,N_7416,N_6205);
or UO_220 (O_220,N_5578,N_5695);
nor UO_221 (O_221,N_9832,N_7616);
and UO_222 (O_222,N_9634,N_8419);
nand UO_223 (O_223,N_9423,N_7548);
nor UO_224 (O_224,N_8488,N_5811);
nand UO_225 (O_225,N_5570,N_8145);
xnor UO_226 (O_226,N_5244,N_6583);
nor UO_227 (O_227,N_8027,N_5177);
xor UO_228 (O_228,N_7479,N_5265);
and UO_229 (O_229,N_6714,N_6676);
nor UO_230 (O_230,N_5016,N_7764);
or UO_231 (O_231,N_5663,N_6374);
xor UO_232 (O_232,N_5252,N_7134);
xnor UO_233 (O_233,N_9448,N_8833);
and UO_234 (O_234,N_5543,N_7415);
nand UO_235 (O_235,N_5355,N_5735);
or UO_236 (O_236,N_8937,N_6696);
nor UO_237 (O_237,N_9307,N_6101);
xnor UO_238 (O_238,N_7888,N_8709);
xor UO_239 (O_239,N_9022,N_8254);
nand UO_240 (O_240,N_5610,N_6125);
nand UO_241 (O_241,N_6225,N_6201);
and UO_242 (O_242,N_8910,N_9937);
and UO_243 (O_243,N_5467,N_8891);
and UO_244 (O_244,N_5167,N_8830);
nor UO_245 (O_245,N_8846,N_5582);
and UO_246 (O_246,N_9143,N_5519);
xnor UO_247 (O_247,N_8712,N_6767);
or UO_248 (O_248,N_8169,N_6256);
and UO_249 (O_249,N_6055,N_6064);
nand UO_250 (O_250,N_7191,N_7546);
or UO_251 (O_251,N_9595,N_8301);
xnor UO_252 (O_252,N_8814,N_6724);
or UO_253 (O_253,N_5608,N_7757);
and UO_254 (O_254,N_8714,N_8280);
nand UO_255 (O_255,N_8045,N_8291);
xor UO_256 (O_256,N_5716,N_6602);
xnor UO_257 (O_257,N_5651,N_7966);
nor UO_258 (O_258,N_6979,N_7746);
or UO_259 (O_259,N_9437,N_7614);
or UO_260 (O_260,N_6108,N_5946);
nor UO_261 (O_261,N_9770,N_8402);
or UO_262 (O_262,N_8345,N_6966);
nor UO_263 (O_263,N_8089,N_5309);
or UO_264 (O_264,N_8963,N_7291);
nor UO_265 (O_265,N_6075,N_8978);
or UO_266 (O_266,N_9329,N_6066);
xor UO_267 (O_267,N_6948,N_8707);
xnor UO_268 (O_268,N_9543,N_7178);
nand UO_269 (O_269,N_5928,N_8817);
xnor UO_270 (O_270,N_6184,N_9208);
or UO_271 (O_271,N_6235,N_7806);
or UO_272 (O_272,N_7916,N_5824);
or UO_273 (O_273,N_5203,N_8099);
nor UO_274 (O_274,N_5152,N_6896);
nand UO_275 (O_275,N_8591,N_7407);
nand UO_276 (O_276,N_5827,N_7539);
or UO_277 (O_277,N_8505,N_6080);
and UO_278 (O_278,N_5989,N_7272);
nand UO_279 (O_279,N_5439,N_9926);
nor UO_280 (O_280,N_9619,N_5802);
nor UO_281 (O_281,N_9709,N_9834);
and UO_282 (O_282,N_5630,N_8729);
xor UO_283 (O_283,N_9113,N_9295);
xnor UO_284 (O_284,N_7258,N_6213);
xor UO_285 (O_285,N_7104,N_7974);
nor UO_286 (O_286,N_6239,N_9583);
and UO_287 (O_287,N_6315,N_7973);
nor UO_288 (O_288,N_5106,N_8166);
and UO_289 (O_289,N_7862,N_8050);
and UO_290 (O_290,N_8061,N_5231);
or UO_291 (O_291,N_8887,N_6707);
xnor UO_292 (O_292,N_8681,N_7724);
nand UO_293 (O_293,N_7360,N_6673);
or UO_294 (O_294,N_7277,N_6547);
nand UO_295 (O_295,N_8972,N_6372);
or UO_296 (O_296,N_6280,N_7458);
nand UO_297 (O_297,N_7069,N_6974);
or UO_298 (O_298,N_9122,N_5013);
nor UO_299 (O_299,N_6965,N_7897);
nor UO_300 (O_300,N_8465,N_5147);
and UO_301 (O_301,N_8198,N_8137);
xnor UO_302 (O_302,N_5294,N_5722);
or UO_303 (O_303,N_6883,N_5014);
nor UO_304 (O_304,N_9369,N_7179);
nand UO_305 (O_305,N_5942,N_5292);
and UO_306 (O_306,N_5574,N_8838);
or UO_307 (O_307,N_9593,N_8701);
and UO_308 (O_308,N_7397,N_8745);
nor UO_309 (O_309,N_8916,N_5870);
or UO_310 (O_310,N_9574,N_8210);
xnor UO_311 (O_311,N_8572,N_7573);
or UO_312 (O_312,N_7243,N_9375);
and UO_313 (O_313,N_6615,N_8367);
and UO_314 (O_314,N_5172,N_6107);
nor UO_315 (O_315,N_5790,N_9266);
nor UO_316 (O_316,N_6637,N_6686);
and UO_317 (O_317,N_5875,N_9223);
nand UO_318 (O_318,N_6872,N_6876);
or UO_319 (O_319,N_5364,N_8612);
nand UO_320 (O_320,N_6807,N_6597);
xor UO_321 (O_321,N_9836,N_7419);
and UO_322 (O_322,N_7830,N_6865);
nor UO_323 (O_323,N_7931,N_6044);
and UO_324 (O_324,N_7054,N_6103);
xor UO_325 (O_325,N_9342,N_7440);
xnor UO_326 (O_326,N_8231,N_8540);
and UO_327 (O_327,N_7682,N_9199);
and UO_328 (O_328,N_5957,N_8750);
nor UO_329 (O_329,N_7057,N_7833);
or UO_330 (O_330,N_6892,N_7623);
xor UO_331 (O_331,N_6731,N_9658);
nor UO_332 (O_332,N_6980,N_7494);
or UO_333 (O_333,N_7426,N_8466);
xnor UO_334 (O_334,N_8801,N_6175);
or UO_335 (O_335,N_9418,N_9826);
nor UO_336 (O_336,N_8823,N_9753);
or UO_337 (O_337,N_8296,N_6613);
xor UO_338 (O_338,N_8199,N_5256);
nor UO_339 (O_339,N_6229,N_8062);
xor UO_340 (O_340,N_7429,N_8418);
and UO_341 (O_341,N_9520,N_8859);
xnor UO_342 (O_342,N_9642,N_6677);
nor UO_343 (O_343,N_5672,N_5567);
xor UO_344 (O_344,N_8723,N_7919);
and UO_345 (O_345,N_5139,N_6508);
nor UO_346 (O_346,N_6579,N_5371);
nand UO_347 (O_347,N_5346,N_6424);
nor UO_348 (O_348,N_6835,N_6675);
nor UO_349 (O_349,N_6661,N_9298);
or UO_350 (O_350,N_7387,N_8624);
or UO_351 (O_351,N_6483,N_5457);
xor UO_352 (O_352,N_5199,N_7362);
or UO_353 (O_353,N_8999,N_9955);
and UO_354 (O_354,N_7219,N_6847);
nand UO_355 (O_355,N_5134,N_5119);
nand UO_356 (O_356,N_6454,N_5340);
xor UO_357 (O_357,N_7670,N_9302);
xnor UO_358 (O_358,N_5627,N_7227);
and UO_359 (O_359,N_6464,N_5117);
and UO_360 (O_360,N_5966,N_9701);
nand UO_361 (O_361,N_7742,N_9589);
nand UO_362 (O_362,N_5545,N_8761);
and UO_363 (O_363,N_6659,N_8432);
xnor UO_364 (O_364,N_8341,N_8942);
and UO_365 (O_365,N_7958,N_9357);
and UO_366 (O_366,N_6431,N_6340);
and UO_367 (O_367,N_9123,N_5689);
xnor UO_368 (O_368,N_7606,N_5375);
nand UO_369 (O_369,N_7707,N_9930);
nor UO_370 (O_370,N_9804,N_7952);
and UO_371 (O_371,N_6741,N_6094);
nor UO_372 (O_372,N_6442,N_8196);
xnor UO_373 (O_373,N_8113,N_9045);
nor UO_374 (O_374,N_5019,N_6631);
xnor UO_375 (O_375,N_9636,N_7537);
and UO_376 (O_376,N_8743,N_8055);
nand UO_377 (O_377,N_6033,N_9400);
and UO_378 (O_378,N_6181,N_9474);
xor UO_379 (O_379,N_9823,N_9354);
nand UO_380 (O_380,N_5728,N_5495);
nand UO_381 (O_381,N_5991,N_8140);
nor UO_382 (O_382,N_7017,N_8379);
or UO_383 (O_383,N_7566,N_8293);
and UO_384 (O_384,N_6930,N_6955);
nand UO_385 (O_385,N_9582,N_9386);
xor UO_386 (O_386,N_6045,N_6574);
and UO_387 (O_387,N_6749,N_9792);
or UO_388 (O_388,N_9702,N_8203);
nor UO_389 (O_389,N_7385,N_8602);
and UO_390 (O_390,N_7289,N_5554);
and UO_391 (O_391,N_9053,N_6863);
or UO_392 (O_392,N_9355,N_9528);
nor UO_393 (O_393,N_7072,N_8703);
nor UO_394 (O_394,N_9606,N_9097);
xor UO_395 (O_395,N_7574,N_7965);
nor UO_396 (O_396,N_6906,N_8812);
or UO_397 (O_397,N_7391,N_7534);
nand UO_398 (O_398,N_6386,N_6060);
xnor UO_399 (O_399,N_7889,N_5972);
nand UO_400 (O_400,N_5416,N_5476);
nand UO_401 (O_401,N_9880,N_5200);
and UO_402 (O_402,N_7513,N_6503);
and UO_403 (O_403,N_7264,N_9328);
nor UO_404 (O_404,N_6539,N_7571);
nor UO_405 (O_405,N_6351,N_6891);
or UO_406 (O_406,N_8119,N_8575);
and UO_407 (O_407,N_7228,N_9013);
or UO_408 (O_408,N_9080,N_5963);
and UO_409 (O_409,N_7152,N_5998);
xnor UO_410 (O_410,N_8362,N_5263);
nor UO_411 (O_411,N_9401,N_6032);
and UO_412 (O_412,N_7096,N_6083);
and UO_413 (O_413,N_6444,N_9763);
xor UO_414 (O_414,N_6496,N_8271);
and UO_415 (O_415,N_7232,N_9977);
nor UO_416 (O_416,N_9268,N_9783);
xor UO_417 (O_417,N_8604,N_9312);
and UO_418 (O_418,N_7132,N_7183);
nand UO_419 (O_419,N_8759,N_6824);
and UO_420 (O_420,N_6718,N_6228);
xnor UO_421 (O_421,N_9919,N_7137);
xor UO_422 (O_422,N_8272,N_8577);
or UO_423 (O_423,N_8758,N_7083);
nor UO_424 (O_424,N_6706,N_6436);
xor UO_425 (O_425,N_5286,N_9940);
nor UO_426 (O_426,N_5868,N_9840);
xor UO_427 (O_427,N_6958,N_9797);
xor UO_428 (O_428,N_7029,N_5539);
or UO_429 (O_429,N_5632,N_7570);
or UO_430 (O_430,N_7156,N_6497);
nor UO_431 (O_431,N_8479,N_7410);
or UO_432 (O_432,N_9508,N_8138);
nor UO_433 (O_433,N_5065,N_8876);
and UO_434 (O_434,N_5596,N_5356);
nand UO_435 (O_435,N_6535,N_5565);
and UO_436 (O_436,N_6164,N_9539);
xor UO_437 (O_437,N_6961,N_5877);
nor UO_438 (O_438,N_5361,N_7602);
and UO_439 (O_439,N_9231,N_9995);
and UO_440 (O_440,N_5377,N_6316);
and UO_441 (O_441,N_9513,N_7306);
or UO_442 (O_442,N_8926,N_7136);
xor UO_443 (O_443,N_9849,N_8387);
or UO_444 (O_444,N_7981,N_8143);
and UO_445 (O_445,N_6964,N_8775);
xor UO_446 (O_446,N_5383,N_5284);
or UO_447 (O_447,N_5999,N_9947);
xor UO_448 (O_448,N_6956,N_6022);
nor UO_449 (O_449,N_7390,N_8605);
nor UO_450 (O_450,N_5640,N_9654);
or UO_451 (O_451,N_6894,N_6760);
and UO_452 (O_452,N_5838,N_6952);
xnor UO_453 (O_453,N_9015,N_9402);
and UO_454 (O_454,N_6363,N_6527);
nor UO_455 (O_455,N_8722,N_7244);
xnor UO_456 (O_456,N_9404,N_5769);
and UO_457 (O_457,N_6486,N_5656);
xnor UO_458 (O_458,N_8990,N_5914);
or UO_459 (O_459,N_5618,N_7667);
and UO_460 (O_460,N_7624,N_8056);
xor UO_461 (O_461,N_5221,N_9093);
and UO_462 (O_462,N_9156,N_8422);
or UO_463 (O_463,N_7316,N_6203);
or UO_464 (O_464,N_7147,N_8726);
and UO_465 (O_465,N_8095,N_9626);
nor UO_466 (O_466,N_8252,N_6246);
xor UO_467 (O_467,N_9489,N_8564);
nand UO_468 (O_468,N_7015,N_7560);
nand UO_469 (O_469,N_7857,N_9843);
xnor UO_470 (O_470,N_6839,N_6329);
or UO_471 (O_471,N_7994,N_9599);
and UO_472 (O_472,N_9693,N_7174);
nor UO_473 (O_473,N_8413,N_9322);
nand UO_474 (O_474,N_9504,N_9863);
xor UO_475 (O_475,N_6285,N_8219);
and UO_476 (O_476,N_8337,N_7339);
and UO_477 (O_477,N_7087,N_7050);
and UO_478 (O_478,N_6864,N_5643);
nand UO_479 (O_479,N_5386,N_8956);
nand UO_480 (O_480,N_5864,N_5452);
and UO_481 (O_481,N_9169,N_7467);
or UO_482 (O_482,N_9666,N_5697);
and UO_483 (O_483,N_5291,N_7462);
xor UO_484 (O_484,N_9747,N_9482);
nor UO_485 (O_485,N_7045,N_9506);
and UO_486 (O_486,N_9572,N_5997);
xnor UO_487 (O_487,N_9733,N_8015);
or UO_488 (O_488,N_6789,N_9812);
nor UO_489 (O_489,N_8192,N_8226);
nand UO_490 (O_490,N_9396,N_8971);
xnor UO_491 (O_491,N_8569,N_8929);
nand UO_492 (O_492,N_6705,N_6900);
or UO_493 (O_493,N_7013,N_6543);
and UO_494 (O_494,N_7185,N_7138);
xor UO_495 (O_495,N_7214,N_9713);
or UO_496 (O_496,N_7549,N_5542);
xnor UO_497 (O_497,N_8365,N_7977);
or UO_498 (O_498,N_6095,N_5149);
nand UO_499 (O_499,N_8687,N_8450);
and UO_500 (O_500,N_9875,N_8486);
nor UO_501 (O_501,N_5360,N_7107);
xor UO_502 (O_502,N_8400,N_5448);
or UO_503 (O_503,N_6371,N_9087);
nand UO_504 (O_504,N_5681,N_8121);
or UO_505 (O_505,N_7748,N_8835);
or UO_506 (O_506,N_5068,N_6375);
or UO_507 (O_507,N_9990,N_9938);
nand UO_508 (O_508,N_8877,N_9378);
or UO_509 (O_509,N_9739,N_5885);
nand UO_510 (O_510,N_9259,N_6220);
nor UO_511 (O_511,N_8716,N_5883);
and UO_512 (O_512,N_7450,N_5211);
nor UO_513 (O_513,N_7935,N_5625);
xnor UO_514 (O_514,N_9576,N_7237);
xor UO_515 (O_515,N_8867,N_8316);
xnor UO_516 (O_516,N_7161,N_8395);
or UO_517 (O_517,N_8216,N_5505);
nand UO_518 (O_518,N_8647,N_7909);
nor UO_519 (O_519,N_7259,N_7043);
and UO_520 (O_520,N_5723,N_5399);
nor UO_521 (O_521,N_6569,N_6977);
xor UO_522 (O_522,N_5005,N_6666);
or UO_523 (O_523,N_9799,N_8770);
nor UO_524 (O_524,N_8047,N_5426);
nor UO_525 (O_525,N_8117,N_6406);
nor UO_526 (O_526,N_6640,N_7814);
xnor UO_527 (O_527,N_9988,N_6279);
and UO_528 (O_528,N_5561,N_8840);
xnor UO_529 (O_529,N_7324,N_8653);
nand UO_530 (O_530,N_6541,N_5196);
xnor UO_531 (O_531,N_6104,N_7347);
and UO_532 (O_532,N_8108,N_5446);
and UO_533 (O_533,N_9120,N_5473);
and UO_534 (O_534,N_7959,N_9835);
and UO_535 (O_535,N_9071,N_5756);
and UO_536 (O_536,N_7715,N_6927);
nand UO_537 (O_537,N_9536,N_7590);
nor UO_538 (O_538,N_9525,N_8288);
or UO_539 (O_539,N_6014,N_8262);
nand UO_540 (O_540,N_7650,N_5317);
xnor UO_541 (O_541,N_7349,N_6612);
nor UO_542 (O_542,N_7955,N_7182);
nor UO_543 (O_543,N_8954,N_5330);
nor UO_544 (O_544,N_6334,N_6404);
and UO_545 (O_545,N_5743,N_7668);
or UO_546 (O_546,N_8320,N_8104);
and UO_547 (O_547,N_8431,N_9641);
nand UO_548 (O_548,N_7103,N_5161);
and UO_549 (O_549,N_9441,N_6571);
nand UO_550 (O_550,N_9140,N_7915);
nand UO_551 (O_551,N_6504,N_8530);
xnor UO_552 (O_552,N_8403,N_9200);
nand UO_553 (O_553,N_6470,N_7209);
xnor UO_554 (O_554,N_7578,N_9984);
and UO_555 (O_555,N_7019,N_8377);
and UO_556 (O_556,N_8609,N_8335);
xnor UO_557 (O_557,N_8286,N_5387);
or UO_558 (O_558,N_8212,N_6471);
and UO_559 (O_559,N_5269,N_6185);
xnor UO_560 (O_560,N_7672,N_7438);
or UO_561 (O_561,N_9478,N_9646);
nor UO_562 (O_562,N_9781,N_9301);
xnor UO_563 (O_563,N_7683,N_5455);
and UO_564 (O_564,N_9810,N_9381);
nor UO_565 (O_565,N_8780,N_8659);
and UO_566 (O_566,N_9989,N_5981);
or UO_567 (O_567,N_7162,N_5335);
nand UO_568 (O_568,N_8424,N_8778);
or UO_569 (O_569,N_5289,N_5589);
or UO_570 (O_570,N_8847,N_9493);
xnor UO_571 (O_571,N_6314,N_7167);
and UO_572 (O_572,N_7717,N_6330);
or UO_573 (O_573,N_8407,N_8385);
and UO_574 (O_574,N_5762,N_8943);
and UO_575 (O_575,N_6502,N_7646);
nor UO_576 (O_576,N_7809,N_6746);
nand UO_577 (O_577,N_7855,N_9150);
nand UO_578 (O_578,N_9137,N_7928);
and UO_579 (O_579,N_9932,N_9433);
and UO_580 (O_580,N_7541,N_9587);
nor UO_581 (O_581,N_8969,N_8490);
nand UO_582 (O_582,N_9879,N_8330);
nand UO_583 (O_583,N_5391,N_6258);
or UO_584 (O_584,N_9532,N_7488);
xor UO_585 (O_585,N_5404,N_9258);
and UO_586 (O_586,N_9392,N_9978);
and UO_587 (O_587,N_8535,N_8803);
nand UO_588 (O_588,N_7447,N_7825);
nor UO_589 (O_589,N_8897,N_5922);
nand UO_590 (O_590,N_6823,N_9261);
nor UO_591 (O_591,N_5548,N_7635);
nor UO_592 (O_592,N_6248,N_6182);
nor UO_593 (O_593,N_7655,N_7526);
nand UO_594 (O_594,N_7660,N_7451);
or UO_595 (O_595,N_6596,N_9825);
nor UO_596 (O_596,N_8949,N_9735);
xnor UO_597 (O_597,N_9340,N_5049);
nor UO_598 (O_598,N_9522,N_7380);
xnor UO_599 (O_599,N_5492,N_7501);
or UO_600 (O_600,N_8454,N_9343);
nor UO_601 (O_601,N_5008,N_8768);
nor UO_602 (O_602,N_5216,N_7886);
xnor UO_603 (O_603,N_8902,N_5568);
and UO_604 (O_604,N_7055,N_9649);
nor UO_605 (O_605,N_9081,N_7692);
nor UO_606 (O_606,N_8779,N_6925);
nand UO_607 (O_607,N_7605,N_9098);
nand UO_608 (O_608,N_7674,N_8896);
xnor UO_609 (O_609,N_5911,N_7976);
nand UO_610 (O_610,N_7202,N_7934);
and UO_611 (O_611,N_8037,N_7766);
and UO_612 (O_612,N_7925,N_8939);
or UO_613 (O_613,N_7656,N_6902);
and UO_614 (O_614,N_9635,N_8064);
and UO_615 (O_615,N_7811,N_6152);
nor UO_616 (O_616,N_8197,N_9228);
or UO_617 (O_617,N_7090,N_6154);
nor UO_618 (O_618,N_7188,N_9711);
nand UO_619 (O_619,N_9625,N_5463);
xor UO_620 (O_620,N_8747,N_6146);
nand UO_621 (O_621,N_6660,N_7005);
and UO_622 (O_622,N_6445,N_8940);
nor UO_623 (O_623,N_8515,N_6269);
and UO_624 (O_624,N_6097,N_9059);
nor UO_625 (O_625,N_5876,N_8376);
nor UO_626 (O_626,N_7203,N_9017);
xor UO_627 (O_627,N_8430,N_8514);
nor UO_628 (O_628,N_8547,N_5316);
nand UO_629 (O_629,N_7428,N_7923);
or UO_630 (O_630,N_6651,N_5768);
xor UO_631 (O_631,N_5229,N_5034);
nor UO_632 (O_632,N_6608,N_6236);
or UO_633 (O_633,N_6140,N_6272);
and UO_634 (O_634,N_5821,N_7073);
and UO_635 (O_635,N_6124,N_9438);
nor UO_636 (O_636,N_6030,N_5003);
nor UO_637 (O_637,N_7946,N_6556);
or UO_638 (O_638,N_5525,N_9134);
and UO_639 (O_639,N_5682,N_8078);
or UO_640 (O_640,N_5780,N_5799);
xor UO_641 (O_641,N_5886,N_6209);
nor UO_642 (O_642,N_7133,N_9041);
nor UO_643 (O_643,N_5829,N_9992);
nand UO_644 (O_644,N_5219,N_6796);
nor UO_645 (O_645,N_7506,N_6459);
and UO_646 (O_646,N_9638,N_7940);
nor UO_647 (O_647,N_7941,N_7772);
or UO_648 (O_648,N_7968,N_8190);
nand UO_649 (O_649,N_9285,N_8957);
or UO_650 (O_650,N_5326,N_9175);
or UO_651 (O_651,N_8786,N_7671);
nor UO_652 (O_652,N_5830,N_6168);
and UO_653 (O_653,N_5108,N_7801);
xor UO_654 (O_654,N_5962,N_8444);
nor UO_655 (O_655,N_6518,N_9707);
nor UO_656 (O_656,N_8619,N_5970);
and UO_657 (O_657,N_9830,N_6242);
xor UO_658 (O_658,N_6553,N_9074);
and UO_659 (O_659,N_8906,N_7708);
xnor UO_660 (O_660,N_9689,N_9889);
and UO_661 (O_661,N_9759,N_5153);
and UO_662 (O_662,N_9294,N_5421);
nand UO_663 (O_663,N_6499,N_7912);
nor UO_664 (O_664,N_9158,N_6355);
or UO_665 (O_665,N_8401,N_6364);
nor UO_666 (O_666,N_6328,N_9023);
nor UO_667 (O_667,N_5398,N_9972);
xor UO_668 (O_668,N_6456,N_8193);
and UO_669 (O_669,N_8640,N_5792);
and UO_670 (O_670,N_9575,N_5056);
nor UO_671 (O_671,N_7465,N_7442);
or UO_672 (O_672,N_6914,N_7476);
nand UO_673 (O_673,N_7352,N_7436);
xor UO_674 (O_674,N_9691,N_6149);
nor UO_675 (O_675,N_7979,N_9173);
nand UO_676 (O_676,N_9979,N_5867);
nor UO_677 (O_677,N_5951,N_9655);
nor UO_678 (O_678,N_9578,N_5919);
nand UO_679 (O_679,N_8220,N_7894);
xnor UO_680 (O_680,N_9394,N_9471);
xor UO_681 (O_681,N_9581,N_9280);
xor UO_682 (O_682,N_9705,N_8931);
and UO_683 (O_683,N_6561,N_5493);
nand UO_684 (O_684,N_9690,N_8144);
or UO_685 (O_685,N_9253,N_9495);
or UO_686 (O_686,N_7392,N_7400);
nor UO_687 (O_687,N_5892,N_9688);
or UO_688 (O_688,N_6890,N_8038);
nor UO_689 (O_689,N_7716,N_8332);
nor UO_690 (O_690,N_7883,N_9615);
nand UO_691 (O_691,N_9981,N_6537);
nor UO_692 (O_692,N_5046,N_6609);
xnor UO_693 (O_693,N_6156,N_8692);
or UO_694 (O_694,N_9207,N_5067);
or UO_695 (O_695,N_6753,N_6342);
or UO_696 (O_696,N_7712,N_6972);
nor UO_697 (O_697,N_5700,N_9224);
nor UO_698 (O_698,N_5190,N_9965);
nor UO_699 (O_699,N_5379,N_5571);
nand UO_700 (O_700,N_7441,N_6946);
and UO_701 (O_701,N_5727,N_8324);
and UO_702 (O_702,N_6781,N_8323);
nor UO_703 (O_703,N_7238,N_6525);
nand UO_704 (O_704,N_5414,N_9102);
nand UO_705 (O_705,N_9458,N_7696);
nand UO_706 (O_706,N_7014,N_7753);
nor UO_707 (O_707,N_5060,N_7466);
xnor UO_708 (O_708,N_8737,N_5376);
xnor UO_709 (O_709,N_5959,N_5665);
nor UO_710 (O_710,N_6067,N_5585);
and UO_711 (O_711,N_5085,N_8558);
or UO_712 (O_712,N_7097,N_6725);
nor UO_713 (O_713,N_8719,N_5938);
nand UO_714 (O_714,N_8848,N_9974);
or UO_715 (O_715,N_6621,N_7615);
xor UO_716 (O_716,N_7904,N_9717);
nand UO_717 (O_717,N_7859,N_8487);
or UO_718 (O_718,N_7089,N_9704);
xnor UO_719 (O_719,N_8894,N_6478);
xor UO_720 (O_720,N_6388,N_7035);
or UO_721 (O_721,N_7612,N_7939);
nor UO_722 (O_722,N_5741,N_6381);
nand UO_723 (O_723,N_7498,N_7374);
xor UO_724 (O_724,N_7701,N_8446);
nand UO_725 (O_725,N_8209,N_9923);
and UO_726 (O_726,N_6729,N_6266);
or UO_727 (O_727,N_6412,N_6819);
and UO_728 (O_728,N_9547,N_5503);
xnor UO_729 (O_729,N_5465,N_6989);
or UO_730 (O_730,N_5157,N_9262);
nor UO_731 (O_731,N_9111,N_6645);
nand UO_732 (O_732,N_5314,N_6510);
xor UO_733 (O_733,N_5752,N_7240);
and UO_734 (O_734,N_5533,N_9109);
xor UO_735 (O_735,N_8699,N_9562);
and UO_736 (O_736,N_6130,N_8756);
or UO_737 (O_737,N_6862,N_7542);
or UO_738 (O_738,N_5288,N_6719);
or UO_739 (O_739,N_7803,N_5368);
nor UO_740 (O_740,N_8182,N_9353);
xor UO_741 (O_741,N_8356,N_9904);
and UO_742 (O_742,N_6511,N_9326);
nor UO_743 (O_743,N_5278,N_5076);
or UO_744 (O_744,N_7565,N_8635);
nor UO_745 (O_745,N_6399,N_8914);
nand UO_746 (O_746,N_6484,N_6554);
xor UO_747 (O_747,N_9331,N_7697);
or UO_748 (O_748,N_6142,N_5653);
nand UO_749 (O_749,N_5255,N_6102);
xor UO_750 (O_750,N_8806,N_9108);
nor UO_751 (O_751,N_8811,N_7433);
nand UO_752 (O_752,N_5115,N_6218);
and UO_753 (O_753,N_5888,N_9384);
xor UO_754 (O_754,N_8364,N_8884);
xor UO_755 (O_755,N_9569,N_5686);
or UO_756 (O_756,N_5562,N_6255);
nor UO_757 (O_757,N_6937,N_9321);
or UO_758 (O_758,N_7239,N_8201);
and UO_759 (O_759,N_7070,N_9101);
xnor UO_760 (O_760,N_9278,N_7241);
and UO_761 (O_761,N_9209,N_9608);
nor UO_762 (O_762,N_6908,N_9096);
nor UO_763 (O_763,N_9952,N_7393);
or UO_764 (O_764,N_7653,N_6415);
xnor UO_765 (O_765,N_7556,N_6387);
nand UO_766 (O_766,N_5590,N_8241);
and UO_767 (O_767,N_8810,N_5298);
xnor UO_768 (O_768,N_8674,N_8628);
and UO_769 (O_769,N_5246,N_5129);
and UO_770 (O_770,N_9303,N_7505);
nor UO_771 (O_771,N_7799,N_7461);
nand UO_772 (O_772,N_7434,N_6856);
nand UO_773 (O_773,N_6816,N_7621);
and UO_774 (O_774,N_5761,N_5528);
xor UO_775 (O_775,N_7386,N_9790);
and UO_776 (O_776,N_9708,N_6814);
and UO_777 (O_777,N_5007,N_8654);
nand UO_778 (O_778,N_9201,N_8820);
or UO_779 (O_779,N_9885,N_5098);
xor UO_780 (O_780,N_6926,N_9873);
and UO_781 (O_781,N_8629,N_8744);
nand UO_782 (O_782,N_9982,N_8669);
and UO_783 (O_783,N_5915,N_7166);
and UO_784 (O_784,N_9405,N_5642);
or UO_785 (O_785,N_7321,N_9243);
nand UO_786 (O_786,N_9685,N_8561);
nand UO_787 (O_787,N_7626,N_6133);
nand UO_788 (O_788,N_5243,N_9723);
nand UO_789 (O_789,N_9748,N_6144);
or UO_790 (O_790,N_5833,N_9656);
nor UO_791 (O_791,N_7181,N_9415);
and UO_792 (O_792,N_7453,N_5472);
xor UO_793 (O_793,N_6846,N_6924);
xnor UO_794 (O_794,N_5785,N_7460);
nor UO_795 (O_795,N_5392,N_6732);
and UO_796 (O_796,N_9822,N_9188);
nor UO_797 (O_797,N_7326,N_7532);
nor UO_798 (O_798,N_6664,N_6224);
xnor UO_799 (O_799,N_7970,N_9103);
xor UO_800 (O_800,N_6304,N_6557);
and UO_801 (O_801,N_7839,N_8022);
nor UO_802 (O_802,N_6771,N_7364);
xnor UO_803 (O_803,N_6578,N_6069);
or UO_804 (O_804,N_8438,N_8583);
xor UO_805 (O_805,N_7330,N_7942);
nor UO_806 (O_806,N_7197,N_7480);
or UO_807 (O_807,N_7446,N_8538);
or UO_808 (O_808,N_8127,N_7293);
xor UO_809 (O_809,N_5145,N_7184);
nand UO_810 (O_810,N_9445,N_8459);
nand UO_811 (O_811,N_5987,N_8966);
or UO_812 (O_812,N_6449,N_8537);
and UO_813 (O_813,N_6222,N_5026);
nand UO_814 (O_814,N_7022,N_6006);
nand UO_815 (O_815,N_8060,N_7911);
or UO_816 (O_816,N_5509,N_7464);
xor UO_817 (O_817,N_8091,N_7278);
or UO_818 (O_818,N_6487,N_8895);
nand UO_819 (O_819,N_8399,N_8461);
or UO_820 (O_820,N_7281,N_5645);
or UO_821 (O_821,N_6273,N_9584);
nor UO_822 (O_822,N_5185,N_9958);
or UO_823 (O_823,N_5737,N_8829);
nand UO_824 (O_824,N_5418,N_8200);
and UO_825 (O_825,N_5181,N_8748);
or UO_826 (O_826,N_5150,N_9014);
nor UO_827 (O_827,N_5223,N_7077);
xnor UO_828 (O_828,N_5817,N_9467);
nand UO_829 (O_829,N_7543,N_7348);
nor UO_830 (O_830,N_9538,N_6309);
or UO_831 (O_831,N_7444,N_5058);
and UO_832 (O_832,N_5037,N_7211);
and UO_833 (O_833,N_7267,N_6679);
nor UO_834 (O_834,N_9549,N_9488);
nand UO_835 (O_835,N_8622,N_9349);
or UO_836 (O_836,N_9403,N_7829);
nor UO_837 (O_837,N_9852,N_7345);
and UO_838 (O_838,N_5339,N_6061);
nor UO_839 (O_839,N_8412,N_9677);
and UO_840 (O_840,N_9645,N_8741);
xor UO_841 (O_841,N_7499,N_5786);
or UO_842 (O_842,N_8933,N_6833);
and UO_843 (O_843,N_9480,N_9490);
and UO_844 (O_844,N_5272,N_5726);
xnor UO_845 (O_845,N_6396,N_9969);
xnor UO_846 (O_846,N_5127,N_7189);
nor UO_847 (O_847,N_7903,N_9975);
nor UO_848 (O_848,N_6775,N_5287);
or UO_849 (O_849,N_5130,N_8664);
nand UO_850 (O_850,N_7064,N_9025);
nor UO_851 (O_851,N_5123,N_6647);
and UO_852 (O_852,N_5325,N_5952);
or UO_853 (O_853,N_5828,N_8792);
xor UO_854 (O_854,N_6373,N_6919);
and UO_855 (O_855,N_9839,N_5587);
and UO_856 (O_856,N_5775,N_5273);
xor UO_857 (O_857,N_9206,N_7493);
nand UO_858 (O_858,N_5359,N_6868);
and UO_859 (O_859,N_7609,N_7443);
xnor UO_860 (O_860,N_6873,N_8824);
nand UO_861 (O_861,N_7529,N_6690);
nor UO_862 (O_862,N_8383,N_7010);
xor UO_863 (O_863,N_8542,N_9507);
nor UO_864 (O_864,N_5620,N_9459);
nor UO_865 (O_865,N_6849,N_8721);
nor UO_866 (O_866,N_8697,N_5560);
and UO_867 (O_867,N_9335,N_9388);
or UO_868 (O_868,N_6936,N_8700);
nor UO_869 (O_869,N_7629,N_7572);
and UO_870 (O_870,N_7820,N_9057);
or UO_871 (O_871,N_8851,N_5534);
and UO_872 (O_872,N_6848,N_9592);
and UO_873 (O_873,N_8425,N_8105);
or UO_874 (O_874,N_9319,N_6821);
xnor UO_875 (O_875,N_5052,N_9363);
nand UO_876 (O_876,N_5471,N_5947);
xor UO_877 (O_877,N_5704,N_9426);
and UO_878 (O_878,N_7524,N_9860);
nand UO_879 (O_879,N_6963,N_5345);
nand UO_880 (O_880,N_5348,N_8705);
and UO_881 (O_881,N_9084,N_5856);
nor UO_882 (O_882,N_5616,N_5591);
or UO_883 (O_883,N_8548,N_7300);
nor UO_884 (O_884,N_9933,N_8452);
or UO_885 (O_885,N_7613,N_6128);
and UO_886 (O_886,N_9460,N_7673);
nor UO_887 (O_887,N_8598,N_6933);
or UO_888 (O_888,N_6448,N_8821);
or UO_889 (O_889,N_9942,N_7698);
and UO_890 (O_890,N_5960,N_9457);
xor UO_891 (O_891,N_6195,N_8011);
xor UO_892 (O_892,N_7586,N_8677);
nor UO_893 (O_893,N_7636,N_9274);
nand UO_894 (O_894,N_5805,N_9571);
and UO_895 (O_895,N_9127,N_9682);
or UO_896 (O_896,N_7491,N_7068);
nand UO_897 (O_897,N_9881,N_9661);
and UO_898 (O_898,N_7372,N_9414);
nor UO_899 (O_899,N_8177,N_8172);
and UO_900 (O_900,N_7841,N_7827);
nor UO_901 (O_901,N_8093,N_6451);
and UO_902 (O_902,N_6506,N_8597);
xor UO_903 (O_903,N_7733,N_8184);
nand UO_904 (O_904,N_9073,N_6395);
nor UO_905 (O_905,N_5604,N_7754);
and UO_906 (O_906,N_7368,N_8706);
nor UO_907 (O_907,N_5599,N_7485);
or UO_908 (O_908,N_9751,N_9246);
nand UO_909 (O_909,N_8094,N_8302);
and UO_910 (O_910,N_7105,N_9884);
nand UO_911 (O_911,N_9311,N_6752);
nand UO_912 (O_912,N_5862,N_7130);
nor UO_913 (O_913,N_8307,N_7221);
nand UO_914 (O_914,N_7589,N_9366);
or UO_915 (O_915,N_9845,N_7600);
or UO_916 (O_916,N_5164,N_8234);
nand UO_917 (O_917,N_9130,N_7864);
and UO_918 (O_918,N_9591,N_5541);
or UO_919 (O_919,N_6805,N_7168);
nand UO_920 (O_920,N_9828,N_8727);
nand UO_921 (O_921,N_9346,N_9148);
xnor UO_922 (O_922,N_8000,N_5552);
nor UO_923 (O_923,N_7985,N_9479);
nor UO_924 (O_924,N_9515,N_7303);
xnor UO_925 (O_925,N_5685,N_7413);
or UO_926 (O_926,N_6913,N_8194);
or UO_927 (O_927,N_9566,N_8908);
nand UO_928 (O_928,N_5631,N_7016);
or UO_929 (O_929,N_9851,N_6341);
or UO_930 (O_930,N_8732,N_8585);
or UO_931 (O_931,N_6024,N_7700);
nand UO_932 (O_932,N_8757,N_6973);
nand UO_933 (O_933,N_8041,N_5225);
nor UO_934 (O_934,N_8630,N_6828);
nand UO_935 (O_935,N_9561,N_6096);
nor UO_936 (O_936,N_6465,N_8960);
or UO_937 (O_937,N_5547,N_8787);
nor UO_938 (O_938,N_9556,N_7567);
or UO_939 (O_939,N_5010,N_5865);
and UO_940 (O_940,N_6343,N_5224);
nor UO_941 (O_941,N_8176,N_8584);
and UO_942 (O_942,N_8865,N_9917);
xnor UO_943 (O_943,N_8085,N_5496);
nor UO_944 (O_944,N_5719,N_9219);
xnor UO_945 (O_945,N_7921,N_8433);
xor UO_946 (O_946,N_5699,N_8720);
xnor UO_947 (O_947,N_7483,N_9648);
nand UO_948 (O_948,N_8408,N_8679);
nor UO_949 (O_949,N_5652,N_7847);
or UO_950 (O_950,N_5400,N_5180);
xnor UO_951 (O_951,N_8565,N_6531);
xnor UO_952 (O_952,N_7922,N_8785);
or UO_953 (O_953,N_9652,N_7779);
nor UO_954 (O_954,N_8173,N_5958);
nand UO_955 (O_955,N_9234,N_6826);
and UO_956 (O_956,N_6768,N_7233);
and UO_957 (O_957,N_9596,N_7657);
or UO_958 (O_958,N_7418,N_6112);
or UO_959 (O_959,N_9829,N_5186);
or UO_960 (O_960,N_6617,N_8553);
nor UO_961 (O_961,N_9920,N_8827);
nor UO_962 (O_962,N_8416,N_9800);
and UO_963 (O_963,N_7124,N_7932);
and UO_964 (O_964,N_6743,N_9131);
xor UO_965 (O_965,N_7365,N_5306);
and UO_966 (O_966,N_9670,N_7370);
nor UO_967 (O_967,N_9964,N_7205);
xor UO_968 (O_968,N_9476,N_5617);
nand UO_969 (O_969,N_5412,N_5816);
nor UO_970 (O_970,N_6650,N_8477);
nand UO_971 (O_971,N_5242,N_5675);
and UO_972 (O_972,N_8921,N_8562);
or UO_973 (O_973,N_5797,N_8749);
or UO_974 (O_974,N_8961,N_7858);
nor UO_975 (O_975,N_7804,N_9637);
and UO_976 (O_976,N_8834,N_5850);
and UO_977 (O_977,N_6462,N_6797);
or UO_978 (O_978,N_8866,N_5248);
xor UO_979 (O_979,N_5125,N_8766);
nor UO_980 (O_980,N_8509,N_7026);
or UO_981 (O_981,N_5417,N_6853);
or UO_982 (O_982,N_5882,N_7195);
xor UO_983 (O_983,N_8351,N_7645);
nand UO_984 (O_984,N_8247,N_9643);
and UO_985 (O_985,N_9217,N_6389);
nor UO_986 (O_986,N_6305,N_7310);
xor UO_987 (O_987,N_5923,N_5822);
nor UO_988 (O_988,N_8987,N_5826);
nor UO_989 (O_989,N_9286,N_7144);
nand UO_990 (O_990,N_8318,N_8636);
nor UO_991 (O_991,N_8881,N_9744);
and UO_992 (O_992,N_6362,N_8239);
nor UO_993 (O_993,N_8673,N_8277);
and UO_994 (O_994,N_5044,N_6326);
or UO_995 (O_995,N_8686,N_6348);
and UO_996 (O_996,N_9024,N_5352);
or UO_997 (O_997,N_6854,N_5901);
xnor UO_998 (O_998,N_5466,N_8985);
nand UO_999 (O_999,N_7110,N_8049);
and UO_1000 (O_1000,N_9552,N_9806);
or UO_1001 (O_1001,N_8997,N_6084);
nand UO_1002 (O_1002,N_9358,N_7741);
nand UO_1003 (O_1003,N_5831,N_8070);
and UO_1004 (O_1004,N_7729,N_6514);
or UO_1005 (O_1005,N_7591,N_6202);
xnor UO_1006 (O_1006,N_6479,N_8331);
nand UO_1007 (O_1007,N_9657,N_5869);
nor UO_1008 (O_1008,N_6493,N_9820);
and UO_1009 (O_1009,N_9409,N_6604);
and UO_1010 (O_1010,N_9913,N_6792);
or UO_1011 (O_1011,N_5893,N_6000);
nand UO_1012 (O_1012,N_6153,N_8378);
nand UO_1013 (O_1013,N_9029,N_9462);
and UO_1014 (O_1014,N_5713,N_7734);
and UO_1015 (O_1015,N_9605,N_6118);
nor UO_1016 (O_1016,N_7718,N_8178);
xnor UO_1017 (O_1017,N_6648,N_7563);
and UO_1018 (O_1018,N_9624,N_9594);
nor UO_1019 (O_1019,N_5766,N_5369);
or UO_1020 (O_1020,N_8153,N_6015);
nor UO_1021 (O_1021,N_9157,N_7854);
or UO_1022 (O_1022,N_8892,N_8151);
nor UO_1023 (O_1023,N_9956,N_6618);
and UO_1024 (O_1024,N_6018,N_9050);
nand UO_1025 (O_1025,N_9095,N_6932);
nor UO_1026 (O_1026,N_8269,N_9925);
nor UO_1027 (O_1027,N_8904,N_5558);
xnor UO_1028 (O_1028,N_7620,N_5382);
nand UO_1029 (O_1029,N_6419,N_9192);
nand UO_1030 (O_1030,N_5880,N_9928);
or UO_1031 (O_1031,N_8221,N_7299);
xnor UO_1032 (O_1032,N_7346,N_9993);
nand UO_1033 (O_1033,N_5254,N_5096);
or UO_1034 (O_1034,N_5791,N_5297);
and UO_1035 (O_1035,N_8994,N_7406);
xor UO_1036 (O_1036,N_9048,N_9994);
nand UO_1037 (O_1037,N_5687,N_8589);
nand UO_1038 (O_1038,N_9440,N_5468);
nor UO_1039 (O_1039,N_6407,N_6564);
xnor UO_1040 (O_1040,N_5425,N_5634);
or UO_1041 (O_1041,N_5788,N_9027);
xnor UO_1042 (O_1042,N_7798,N_9573);
nand UO_1043 (O_1043,N_9966,N_8013);
and UO_1044 (O_1044,N_6885,N_5770);
xor UO_1045 (O_1045,N_6162,N_7457);
and UO_1046 (O_1046,N_5684,N_7651);
or UO_1047 (O_1047,N_7424,N_6549);
or UO_1048 (O_1048,N_9257,N_8767);
and UO_1049 (O_1049,N_6671,N_5994);
xnor UO_1050 (O_1050,N_6584,N_9417);
or UO_1051 (O_1051,N_9914,N_5863);
nand UO_1052 (O_1052,N_7832,N_9330);
or UO_1053 (O_1053,N_7676,N_9998);
xor UO_1054 (O_1054,N_7740,N_7643);
or UO_1055 (O_1055,N_8633,N_9238);
or UO_1056 (O_1056,N_8065,N_7333);
nand UO_1057 (O_1057,N_7215,N_5774);
xor UO_1058 (O_1058,N_5641,N_6614);
or UO_1059 (O_1059,N_6148,N_7880);
or UO_1060 (O_1060,N_7788,N_5087);
nand UO_1061 (O_1061,N_5679,N_5032);
nor UO_1062 (O_1062,N_6960,N_6071);
xor UO_1063 (O_1063,N_7052,N_6020);
and UO_1064 (O_1064,N_8798,N_5929);
nor UO_1065 (O_1065,N_7403,N_8913);
xnor UO_1066 (O_1066,N_9610,N_5773);
xor UO_1067 (O_1067,N_5733,N_7363);
or UO_1068 (O_1068,N_5976,N_7579);
and UO_1069 (O_1069,N_7863,N_5576);
nor UO_1070 (O_1070,N_6632,N_8110);
and UO_1071 (O_1071,N_7796,N_7448);
nand UO_1072 (O_1072,N_9819,N_7131);
nor UO_1073 (O_1073,N_5388,N_9530);
xor UO_1074 (O_1074,N_9651,N_5002);
or UO_1075 (O_1075,N_5602,N_6171);
xnor UO_1076 (O_1076,N_8588,N_7033);
nor UO_1077 (O_1077,N_8563,N_8469);
xor UO_1078 (O_1078,N_6457,N_7095);
nand UO_1079 (O_1079,N_5789,N_6998);
or UO_1080 (O_1080,N_8946,N_9076);
xnor UO_1081 (O_1081,N_6392,N_6437);
nand UO_1082 (O_1082,N_9018,N_6204);
and UO_1083 (O_1083,N_9629,N_5916);
or UO_1084 (O_1084,N_9857,N_8927);
nor UO_1085 (O_1085,N_6240,N_7782);
nand UO_1086 (O_1086,N_7129,N_8317);
nand UO_1087 (O_1087,N_6737,N_9967);
or UO_1088 (O_1088,N_9202,N_5814);
and UO_1089 (O_1089,N_5166,N_5839);
and UO_1090 (O_1090,N_9213,N_5158);
or UO_1091 (O_1091,N_9740,N_8492);
nand UO_1092 (O_1092,N_8032,N_5964);
nor UO_1093 (O_1093,N_9168,N_5321);
nor UO_1094 (O_1094,N_5025,N_5860);
xor UO_1095 (O_1095,N_6953,N_5508);
xor UO_1096 (O_1096,N_5449,N_8278);
xnor UO_1097 (O_1097,N_9789,N_7216);
xor UO_1098 (O_1098,N_8251,N_9434);
xnor UO_1099 (O_1099,N_6159,N_9179);
nor UO_1100 (O_1100,N_7356,N_9112);
nor UO_1101 (O_1101,N_8495,N_8644);
nor UO_1102 (O_1102,N_9379,N_5347);
and UO_1103 (O_1103,N_6782,N_9320);
nor UO_1104 (O_1104,N_5353,N_8694);
and UO_1105 (O_1105,N_5514,N_5018);
and UO_1106 (O_1106,N_5027,N_5209);
xnor UO_1107 (O_1107,N_5676,N_8159);
and UO_1108 (O_1108,N_5890,N_9516);
or UO_1109 (O_1109,N_6754,N_7008);
xnor UO_1110 (O_1110,N_6978,N_5006);
nand UO_1111 (O_1111,N_7584,N_6232);
xnor UO_1112 (O_1112,N_8754,N_5405);
nand UO_1113 (O_1113,N_9037,N_8189);
xnor UO_1114 (O_1114,N_8936,N_5757);
and UO_1115 (O_1115,N_7901,N_8360);
and UO_1116 (O_1116,N_7350,N_5694);
or UO_1117 (O_1117,N_7217,N_5709);
nor UO_1118 (O_1118,N_6622,N_7699);
and UO_1119 (O_1119,N_6715,N_7369);
nand UO_1120 (O_1120,N_7085,N_9971);
or UO_1121 (O_1121,N_6463,N_8661);
or UO_1122 (O_1122,N_9062,N_9924);
and UO_1123 (O_1123,N_9288,N_5611);
nor UO_1124 (O_1124,N_8958,N_7376);
or UO_1125 (O_1125,N_6090,N_5920);
and UO_1126 (O_1126,N_5706,N_9004);
nand UO_1127 (O_1127,N_9767,N_5304);
or UO_1128 (O_1128,N_8111,N_8771);
nand UO_1129 (O_1129,N_9526,N_8248);
xor UO_1130 (O_1130,N_8993,N_7086);
xnor UO_1131 (O_1131,N_8648,N_9072);
nor UO_1132 (O_1132,N_5776,N_9064);
or UO_1133 (O_1133,N_6794,N_6227);
nand UO_1134 (O_1134,N_7145,N_5835);
nand UO_1135 (O_1135,N_6106,N_5573);
nor UO_1136 (O_1136,N_7686,N_7561);
nand UO_1137 (O_1137,N_5753,N_6078);
nor UO_1138 (O_1138,N_8374,N_7001);
and UO_1139 (O_1139,N_8443,N_6021);
and UO_1140 (O_1140,N_7640,N_7575);
xnor UO_1141 (O_1141,N_5978,N_7739);
and UO_1142 (O_1142,N_9184,N_6467);
and UO_1143 (O_1143,N_7472,N_5245);
xor UO_1144 (O_1144,N_5536,N_8208);
xnor UO_1145 (O_1145,N_7154,N_5331);
nand UO_1146 (O_1146,N_9100,N_5362);
xnor UO_1147 (O_1147,N_5247,N_7383);
nor UO_1148 (O_1148,N_6489,N_6230);
or UO_1149 (O_1149,N_7913,N_6875);
xor UO_1150 (O_1150,N_7745,N_5214);
nor UO_1151 (O_1151,N_8769,N_6147);
nor UO_1152 (O_1152,N_7554,N_8804);
nand UO_1153 (O_1153,N_7826,N_5659);
nor UO_1154 (O_1154,N_8733,N_8973);
nand UO_1155 (O_1155,N_5965,N_6611);
or UO_1156 (O_1156,N_7597,N_5873);
and UO_1157 (O_1157,N_5343,N_6129);
and UO_1158 (O_1158,N_8594,N_9555);
xor UO_1159 (O_1159,N_7190,N_8004);
or UO_1160 (O_1160,N_9408,N_5234);
and UO_1161 (O_1161,N_8074,N_8478);
and UO_1162 (O_1162,N_9865,N_7495);
nand UO_1163 (O_1163,N_5848,N_8552);
and UO_1164 (O_1164,N_5453,N_7059);
nor UO_1165 (O_1165,N_6748,N_7155);
and UO_1166 (O_1166,N_8457,N_8344);
or UO_1167 (O_1167,N_9196,N_8482);
nor UO_1168 (O_1168,N_6043,N_9922);
nor UO_1169 (O_1169,N_6967,N_8717);
or UO_1170 (O_1170,N_7750,N_8885);
and UO_1171 (O_1171,N_9450,N_7879);
xor UO_1172 (O_1172,N_9714,N_9475);
xnor UO_1173 (O_1173,N_9162,N_6113);
xnor UO_1174 (O_1174,N_6025,N_6663);
xnor UO_1175 (O_1175,N_8256,N_7470);
nand UO_1176 (O_1176,N_8414,N_8306);
nor UO_1177 (O_1177,N_9918,N_5710);
xor UO_1178 (O_1178,N_9371,N_7023);
nand UO_1179 (O_1179,N_8772,N_6785);
xnor UO_1180 (O_1180,N_7997,N_7263);
or UO_1181 (O_1181,N_8522,N_6017);
nand UO_1182 (O_1182,N_8236,N_7693);
and UO_1183 (O_1183,N_8255,N_5195);
nor UO_1184 (O_1184,N_9768,N_7198);
or UO_1185 (O_1185,N_8951,N_6366);
nor UO_1186 (O_1186,N_9511,N_6901);
and UO_1187 (O_1187,N_7489,N_6986);
xnor UO_1188 (O_1188,N_6567,N_7063);
or UO_1189 (O_1189,N_5409,N_7404);
nor UO_1190 (O_1190,N_8133,N_7230);
or UO_1191 (O_1191,N_8828,N_6450);
nor UO_1192 (O_1192,N_8397,N_9031);
or UO_1193 (O_1193,N_6524,N_5787);
xnor UO_1194 (O_1194,N_6744,N_9622);
nor UO_1195 (O_1195,N_5840,N_5646);
or UO_1196 (O_1196,N_8688,N_9485);
xor UO_1197 (O_1197,N_5315,N_8704);
or UO_1198 (O_1198,N_5683,N_8794);
nor UO_1199 (O_1199,N_9523,N_6408);
xnor UO_1200 (O_1200,N_5760,N_7402);
xor UO_1201 (O_1201,N_6136,N_5498);
xnor UO_1202 (O_1202,N_6709,N_5843);
nor UO_1203 (O_1203,N_7269,N_5017);
xnor UO_1204 (O_1204,N_6183,N_7114);
xor UO_1205 (O_1205,N_7951,N_9310);
nand UO_1206 (O_1206,N_6174,N_6801);
or UO_1207 (O_1207,N_6662,N_6904);
xnor UO_1208 (O_1208,N_6238,N_6089);
xnor UO_1209 (O_1209,N_7092,N_6196);
and UO_1210 (O_1210,N_7169,N_8872);
and UO_1211 (O_1211,N_5613,N_9147);
or UO_1212 (O_1212,N_6087,N_6170);
xnor UO_1213 (O_1213,N_5336,N_7971);
and UO_1214 (O_1214,N_8328,N_6681);
or UO_1215 (O_1215,N_9837,N_8822);
nor UO_1216 (O_1216,N_6116,N_7342);
and UO_1217 (O_1217,N_7808,N_9718);
and UO_1218 (O_1218,N_9890,N_7361);
nor UO_1219 (O_1219,N_7093,N_8427);
and UO_1220 (O_1220,N_6428,N_9710);
or UO_1221 (O_1221,N_9604,N_8632);
xnor UO_1222 (O_1222,N_7242,N_6385);
nor UO_1223 (O_1223,N_6761,N_5564);
xor UO_1224 (O_1224,N_7702,N_6177);
nor UO_1225 (O_1225,N_9831,N_8831);
xor UO_1226 (O_1226,N_9888,N_9514);
nand UO_1227 (O_1227,N_7025,N_5299);
nand UO_1228 (O_1228,N_5698,N_9377);
nor UO_1229 (O_1229,N_5303,N_5866);
nor UO_1230 (O_1230,N_7982,N_5754);
or UO_1231 (O_1231,N_8057,N_9814);
nor UO_1232 (O_1232,N_8507,N_8003);
nand UO_1233 (O_1233,N_7519,N_5506);
xnor UO_1234 (O_1234,N_7637,N_9287);
xor UO_1235 (O_1235,N_7792,N_9588);
nand UO_1236 (O_1236,N_7218,N_8470);
nand UO_1237 (O_1237,N_6921,N_5666);
nor UO_1238 (O_1238,N_7884,N_9452);
nor UO_1239 (O_1239,N_9850,N_9954);
and UO_1240 (O_1240,N_6545,N_7776);
nor UO_1241 (O_1241,N_6337,N_5527);
xor UO_1242 (O_1242,N_8582,N_6114);
and UO_1243 (O_1243,N_7173,N_7207);
nor UO_1244 (O_1244,N_8442,N_8340);
and UO_1245 (O_1245,N_7943,N_7918);
or UO_1246 (O_1246,N_8380,N_5896);
and UO_1247 (O_1247,N_7975,N_5988);
or UO_1248 (O_1248,N_6026,N_8922);
nand UO_1249 (O_1249,N_6827,N_6286);
xnor UO_1250 (O_1250,N_7395,N_7705);
or UO_1251 (O_1251,N_6516,N_8339);
nor UO_1252 (O_1252,N_8491,N_5904);
xor UO_1253 (O_1253,N_5451,N_9712);
and UO_1254 (O_1254,N_5334,N_7298);
xnor UO_1255 (O_1255,N_5179,N_7163);
nor UO_1256 (O_1256,N_9818,N_5365);
nand UO_1257 (O_1257,N_7126,N_6249);
xnor UO_1258 (O_1258,N_7924,N_7048);
and UO_1259 (O_1259,N_6494,N_5307);
and UO_1260 (O_1260,N_9764,N_7486);
xor UO_1261 (O_1261,N_5742,N_8965);
nand UO_1262 (O_1262,N_5933,N_6319);
xnor UO_1263 (O_1263,N_9007,N_5170);
nand UO_1264 (O_1264,N_6912,N_7231);
and UO_1265 (O_1265,N_7353,N_7315);
nand UO_1266 (O_1266,N_6111,N_9703);
xor UO_1267 (O_1267,N_7044,N_6057);
nor UO_1268 (O_1268,N_9216,N_9500);
nand UO_1269 (O_1269,N_5118,N_7268);
and UO_1270 (O_1270,N_6512,N_9177);
or UO_1271 (O_1271,N_5159,N_7576);
or UO_1272 (O_1272,N_9333,N_7749);
and UO_1273 (O_1273,N_9435,N_9210);
nand UO_1274 (O_1274,N_6126,N_5664);
xor UO_1275 (O_1275,N_6426,N_6773);
nand UO_1276 (O_1276,N_7373,N_8229);
or UO_1277 (O_1277,N_5202,N_5047);
nand UO_1278 (O_1278,N_8950,N_6784);
nand UO_1279 (O_1279,N_8449,N_6987);
nor UO_1280 (O_1280,N_7887,N_9135);
xor UO_1281 (O_1281,N_8039,N_8789);
xnor UO_1282 (O_1282,N_5407,N_6762);
xor UO_1283 (O_1283,N_7194,N_9519);
nor UO_1284 (O_1284,N_8734,N_5806);
nor UO_1285 (O_1285,N_8453,N_8989);
xnor UO_1286 (O_1286,N_8690,N_5385);
and UO_1287 (O_1287,N_6447,N_7789);
nand UO_1288 (O_1288,N_7714,N_6624);
xor UO_1289 (O_1289,N_8924,N_8411);
and UO_1290 (O_1290,N_9391,N_7817);
nand UO_1291 (O_1291,N_8381,N_9164);
nand UO_1292 (O_1292,N_9681,N_8574);
nand UO_1293 (O_1293,N_6432,N_8230);
and UO_1294 (O_1294,N_8731,N_8611);
nor UO_1295 (O_1295,N_5313,N_6296);
and UO_1296 (O_1296,N_5290,N_5124);
xnor UO_1297 (O_1297,N_6358,N_5969);
and UO_1298 (O_1298,N_8366,N_7294);
or UO_1299 (O_1299,N_9198,N_9895);
and UO_1300 (O_1300,N_7021,N_6598);
or UO_1301 (O_1301,N_8116,N_5271);
or UO_1302 (O_1302,N_8525,N_7675);
xnor UO_1303 (O_1303,N_5357,N_9899);
and UO_1304 (O_1304,N_8903,N_8148);
nor UO_1305 (O_1305,N_5436,N_7067);
nor UO_1306 (O_1306,N_9755,N_6765);
or UO_1307 (O_1307,N_5250,N_6188);
nand UO_1308 (O_1308,N_9225,N_5572);
nor UO_1309 (O_1309,N_6237,N_9373);
nand UO_1310 (O_1310,N_6881,N_6474);
and UO_1311 (O_1311,N_8857,N_7777);
nand UO_1312 (O_1312,N_7892,N_5516);
nand UO_1313 (O_1313,N_8421,N_9240);
xnor UO_1314 (O_1314,N_9339,N_5847);
or UO_1315 (O_1315,N_5238,N_9142);
xor UO_1316 (O_1316,N_9874,N_8617);
and UO_1317 (O_1317,N_5909,N_6257);
xor UO_1318 (O_1318,N_8358,N_8975);
nand UO_1319 (O_1319,N_9119,N_6176);
and UO_1320 (O_1320,N_9756,N_7842);
nand UO_1321 (O_1321,N_9883,N_7452);
xnor UO_1322 (O_1322,N_6068,N_8285);
nand UO_1323 (O_1323,N_5974,N_5577);
xor UO_1324 (O_1324,N_5912,N_7417);
nand UO_1325 (O_1325,N_8257,N_5308);
or UO_1326 (O_1326,N_6544,N_6495);
and UO_1327 (O_1327,N_8832,N_6750);
xnor UO_1328 (O_1328,N_5895,N_9318);
xnor UO_1329 (O_1329,N_9351,N_5236);
or UO_1330 (O_1330,N_9389,N_9968);
or UO_1331 (O_1331,N_6969,N_5277);
and UO_1332 (O_1332,N_7926,N_6606);
or UO_1333 (O_1333,N_9793,N_9910);
nand UO_1334 (O_1334,N_7287,N_8077);
or UO_1335 (O_1335,N_9760,N_5183);
nor UO_1336 (O_1336,N_8150,N_9455);
and UO_1337 (O_1337,N_5042,N_9533);
or UO_1338 (O_1338,N_8912,N_6039);
and UO_1339 (O_1339,N_5148,N_5456);
nor UO_1340 (O_1340,N_5327,N_6991);
nand UO_1341 (O_1341,N_8698,N_7296);
and UO_1342 (O_1342,N_5778,N_9866);
nand UO_1343 (O_1343,N_9118,N_8742);
xnor UO_1344 (O_1344,N_5717,N_9886);
and UO_1345 (O_1345,N_8762,N_9267);
nor UO_1346 (O_1346,N_6215,N_6189);
xor UO_1347 (O_1347,N_7427,N_9779);
or UO_1348 (O_1348,N_6742,N_9732);
nor UO_1349 (O_1349,N_8559,N_7852);
nor UO_1350 (O_1350,N_6759,N_6402);
or UO_1351 (O_1351,N_6260,N_6298);
xor UO_1352 (O_1352,N_7302,N_8508);
or UO_1353 (O_1353,N_5593,N_8131);
nand UO_1354 (O_1354,N_9430,N_6370);
nand UO_1355 (O_1355,N_9181,N_7899);
and UO_1356 (O_1356,N_8167,N_9541);
or UO_1357 (O_1357,N_5491,N_8631);
nor UO_1358 (O_1358,N_8106,N_5342);
nor UO_1359 (O_1359,N_7335,N_7475);
xor UO_1360 (O_1360,N_6100,N_7358);
xor UO_1361 (O_1361,N_6434,N_8800);
and UO_1362 (O_1362,N_8657,N_5510);
nor UO_1363 (O_1363,N_5513,N_8710);
or UO_1364 (O_1364,N_5614,N_8445);
xnor UO_1365 (O_1365,N_6190,N_7399);
and UO_1366 (O_1366,N_5832,N_7953);
nand UO_1367 (O_1367,N_8967,N_7031);
or UO_1368 (O_1368,N_6303,N_6324);
or UO_1369 (O_1369,N_6627,N_8440);
xor UO_1370 (O_1370,N_5217,N_7873);
or UO_1371 (O_1371,N_8342,N_5872);
nor UO_1372 (O_1372,N_5021,N_6352);
nor UO_1373 (O_1373,N_8132,N_7478);
nand UO_1374 (O_1374,N_9896,N_6843);
xor UO_1375 (O_1375,N_6347,N_9795);
or UO_1376 (O_1376,N_8539,N_6694);
nor UO_1377 (O_1377,N_9722,N_6393);
nand UO_1378 (O_1378,N_7738,N_7164);
xnor UO_1379 (O_1379,N_6515,N_8693);
nor UO_1380 (O_1380,N_8984,N_8645);
or UO_1381 (O_1381,N_8870,N_8009);
or UO_1382 (O_1382,N_6830,N_6605);
or UO_1383 (O_1383,N_9846,N_7414);
and UO_1384 (O_1384,N_6806,N_5270);
nor UO_1385 (O_1385,N_9963,N_7608);
nor UO_1386 (O_1386,N_6935,N_9494);
and UO_1387 (O_1387,N_9079,N_5189);
xnor UO_1388 (O_1388,N_8308,N_6837);
and UO_1389 (O_1389,N_6589,N_7210);
and UO_1390 (O_1390,N_9644,N_9859);
nand UO_1391 (O_1391,N_9521,N_9912);
nand UO_1392 (O_1392,N_6812,N_7664);
xor UO_1393 (O_1393,N_9949,N_8086);
nor UO_1394 (O_1394,N_5692,N_5612);
xnor UO_1395 (O_1395,N_7135,N_8410);
and UO_1396 (O_1396,N_8521,N_6692);
xnor UO_1397 (O_1397,N_9864,N_5521);
and UO_1398 (O_1398,N_8020,N_9273);
nor UO_1399 (O_1399,N_9447,N_5607);
nand UO_1400 (O_1400,N_5165,N_5113);
nor UO_1401 (O_1401,N_5588,N_7336);
or UO_1402 (O_1402,N_6250,N_6563);
nor UO_1403 (O_1403,N_8549,N_5777);
nand UO_1404 (O_1404,N_6076,N_7165);
or UO_1405 (O_1405,N_7844,N_5187);
xnor UO_1406 (O_1406,N_5033,N_9567);
or UO_1407 (O_1407,N_5029,N_8336);
nand UO_1408 (O_1408,N_8267,N_8136);
xor UO_1409 (O_1409,N_7140,N_6321);
xor UO_1410 (O_1410,N_6842,N_6010);
nand UO_1411 (O_1411,N_9550,N_6984);
or UO_1412 (O_1412,N_9663,N_8012);
xor UO_1413 (O_1413,N_7411,N_8996);
nand UO_1414 (O_1414,N_8170,N_6513);
xnor UO_1415 (O_1415,N_7882,N_9153);
or UO_1416 (O_1416,N_9774,N_7079);
and UO_1417 (O_1417,N_5154,N_9065);
nand UO_1418 (O_1418,N_7622,N_7593);
xnor UO_1419 (O_1419,N_5755,N_9145);
nand UO_1420 (O_1420,N_7538,N_6019);
and UO_1421 (O_1421,N_6920,N_5444);
nor UO_1422 (O_1422,N_9620,N_5734);
and UO_1423 (O_1423,N_6657,N_8691);
or UO_1424 (O_1424,N_7009,N_9659);
and UO_1425 (O_1425,N_6441,N_8519);
xor UO_1426 (O_1426,N_5605,N_8982);
xnor UO_1427 (O_1427,N_5639,N_9364);
nand UO_1428 (O_1428,N_9180,N_7469);
nand UO_1429 (O_1429,N_9160,N_8527);
nand UO_1430 (O_1430,N_5437,N_9309);
xnor UO_1431 (O_1431,N_7490,N_7002);
xor UO_1432 (O_1432,N_6056,N_5497);
and UO_1433 (O_1433,N_8204,N_9284);
or UO_1434 (O_1434,N_5012,N_5169);
or UO_1435 (O_1435,N_9862,N_7274);
and UO_1436 (O_1436,N_8001,N_8319);
or UO_1437 (O_1437,N_8510,N_5337);
or UO_1438 (O_1438,N_9537,N_8227);
nand UO_1439 (O_1439,N_8299,N_9729);
or UO_1440 (O_1440,N_7908,N_7088);
nand UO_1441 (O_1441,N_8554,N_5447);
nor UO_1442 (O_1442,N_8909,N_7948);
nand UO_1443 (O_1443,N_7246,N_8054);
xor UO_1444 (O_1444,N_8524,N_8816);
or UO_1445 (O_1445,N_6277,N_9385);
xnor UO_1446 (O_1446,N_7770,N_7587);
and UO_1447 (O_1447,N_7843,N_8765);
xnor UO_1448 (O_1448,N_7569,N_6658);
and UO_1449 (O_1449,N_9336,N_9011);
or UO_1450 (O_1450,N_9094,N_8338);
nand UO_1451 (O_1451,N_8240,N_5739);
or UO_1452 (O_1452,N_7816,N_7822);
nor UO_1453 (O_1453,N_8046,N_6369);
xor UO_1454 (O_1454,N_5600,N_8860);
nand UO_1455 (O_1455,N_6836,N_5594);
xor UO_1456 (O_1456,N_7247,N_6670);
xor UO_1457 (O_1457,N_6573,N_6416);
xor UO_1458 (O_1458,N_6481,N_6091);
and UO_1459 (O_1459,N_9529,N_9290);
or UO_1460 (O_1460,N_6059,N_8406);
and UO_1461 (O_1461,N_9734,N_8160);
xor UO_1462 (O_1462,N_6433,N_7225);
nor UO_1463 (O_1463,N_9383,N_6254);
and UO_1464 (O_1464,N_7431,N_9741);
nand UO_1465 (O_1465,N_5889,N_6391);
nor UO_1466 (O_1466,N_7265,N_7379);
and UO_1467 (O_1467,N_5279,N_6834);
nor UO_1468 (O_1468,N_8107,N_7592);
nor UO_1469 (O_1469,N_6422,N_8683);
nor UO_1470 (O_1470,N_7338,N_7006);
nor UO_1471 (O_1471,N_8836,N_7896);
xnor UO_1472 (O_1472,N_6145,N_8472);
xnor UO_1473 (O_1473,N_8689,N_6265);
xnor UO_1474 (O_1474,N_6697,N_9174);
nor UO_1475 (O_1475,N_5747,N_7802);
xor UO_1476 (O_1476,N_8315,N_5549);
nor UO_1477 (O_1477,N_9036,N_9019);
nor UO_1478 (O_1478,N_9785,N_5702);
nand UO_1479 (O_1479,N_8392,N_5443);
nand UO_1480 (O_1480,N_5241,N_8649);
or UO_1481 (O_1481,N_8187,N_9256);
or UO_1482 (O_1482,N_6993,N_6473);
or UO_1483 (O_1483,N_9662,N_5043);
or UO_1484 (O_1484,N_9613,N_6947);
nor UO_1485 (O_1485,N_9674,N_7474);
nor UO_1486 (O_1486,N_6155,N_6874);
nor UO_1487 (O_1487,N_7098,N_7256);
and UO_1488 (O_1488,N_7018,N_5720);
and UO_1489 (O_1489,N_9220,N_7249);
nor UO_1490 (O_1490,N_8298,N_9684);
xnor UO_1491 (O_1491,N_6151,N_8621);
nor UO_1492 (O_1492,N_8667,N_6157);
or UO_1493 (O_1493,N_6306,N_5100);
and UO_1494 (O_1494,N_7568,N_7196);
xnor UO_1495 (O_1495,N_5162,N_9929);
and UO_1496 (O_1496,N_6997,N_7585);
and UO_1497 (O_1497,N_7004,N_6691);
nand UO_1498 (O_1498,N_9775,N_6082);
nand UO_1499 (O_1499,N_7382,N_9067);
endmodule