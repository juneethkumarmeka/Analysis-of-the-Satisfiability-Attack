module basic_2000_20000_2500_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1954,In_536);
nand U1 (N_1,In_186,In_943);
nor U2 (N_2,In_1799,In_1748);
or U3 (N_3,In_328,In_1559);
nor U4 (N_4,In_621,In_672);
or U5 (N_5,In_1042,In_1665);
nand U6 (N_6,In_1147,In_766);
or U7 (N_7,In_1103,In_155);
nand U8 (N_8,In_1771,In_729);
or U9 (N_9,In_708,In_930);
and U10 (N_10,In_739,In_1668);
or U11 (N_11,In_1045,In_1900);
xor U12 (N_12,In_1349,In_1208);
xnor U13 (N_13,In_234,In_427);
or U14 (N_14,In_128,In_1326);
nand U15 (N_15,In_99,In_480);
and U16 (N_16,In_515,In_1784);
and U17 (N_17,In_32,In_201);
xor U18 (N_18,In_1882,In_704);
nor U19 (N_19,In_1672,In_1416);
xnor U20 (N_20,In_1584,In_601);
nand U21 (N_21,In_1651,In_1593);
and U22 (N_22,In_1156,In_1294);
and U23 (N_23,In_1475,In_1544);
nor U24 (N_24,In_563,In_540);
nand U25 (N_25,In_1946,In_1090);
and U26 (N_26,In_1082,In_1387);
nand U27 (N_27,In_1497,In_486);
nor U28 (N_28,In_873,In_1253);
or U29 (N_29,In_221,In_583);
nor U30 (N_30,In_249,In_1749);
nor U31 (N_31,In_1774,In_1311);
nand U32 (N_32,In_240,In_1944);
nor U33 (N_33,In_1513,In_773);
and U34 (N_34,In_1605,In_403);
nand U35 (N_35,In_492,In_737);
nor U36 (N_36,In_503,In_317);
or U37 (N_37,In_830,In_1688);
or U38 (N_38,In_228,In_179);
nor U39 (N_39,In_1177,In_1409);
and U40 (N_40,In_802,In_40);
or U41 (N_41,In_588,In_612);
and U42 (N_42,In_1985,In_886);
and U43 (N_43,In_831,In_558);
xor U44 (N_44,In_1226,In_1747);
nand U45 (N_45,In_898,In_150);
nor U46 (N_46,In_1547,In_1967);
and U47 (N_47,In_1624,In_730);
nand U48 (N_48,In_1183,In_198);
nand U49 (N_49,In_557,In_523);
and U50 (N_50,In_33,In_1769);
and U51 (N_51,In_717,In_1172);
nand U52 (N_52,In_799,In_1104);
or U53 (N_53,In_1730,In_185);
nor U54 (N_54,In_241,In_8);
nand U55 (N_55,In_357,In_177);
and U56 (N_56,In_552,In_1667);
and U57 (N_57,In_531,In_767);
or U58 (N_58,In_291,In_67);
and U59 (N_59,In_1278,In_1427);
or U60 (N_60,In_209,In_1831);
xor U61 (N_61,In_751,In_821);
nand U62 (N_62,In_1167,In_1869);
or U63 (N_63,In_1453,In_1155);
nand U64 (N_64,In_1210,In_1468);
or U65 (N_65,In_215,In_891);
nand U66 (N_66,In_1778,In_297);
xnor U67 (N_67,In_1934,In_1603);
or U68 (N_68,In_1549,In_1890);
and U69 (N_69,In_1275,In_755);
or U70 (N_70,In_835,In_1928);
or U71 (N_71,In_1896,In_334);
and U72 (N_72,In_1841,In_624);
nor U73 (N_73,In_193,In_1578);
or U74 (N_74,In_347,In_736);
nand U75 (N_75,In_1775,In_725);
nor U76 (N_76,In_1997,In_1840);
nand U77 (N_77,In_928,In_1227);
nor U78 (N_78,In_1010,In_1884);
and U79 (N_79,In_1982,In_649);
and U80 (N_80,In_1408,In_1366);
nand U81 (N_81,In_1382,In_1198);
xnor U82 (N_82,In_1848,In_1063);
or U83 (N_83,In_1096,In_1034);
or U84 (N_84,In_1049,In_753);
nand U85 (N_85,In_1360,In_1650);
or U86 (N_86,In_1480,In_1136);
nand U87 (N_87,In_545,In_1850);
nor U88 (N_88,In_146,In_616);
nand U89 (N_89,In_1331,In_306);
nand U90 (N_90,In_1643,In_761);
xnor U91 (N_91,In_867,In_1361);
nand U92 (N_92,In_1510,In_1246);
and U93 (N_93,In_1597,In_996);
nand U94 (N_94,In_1904,In_532);
nor U95 (N_95,In_1916,In_775);
or U96 (N_96,In_527,In_166);
nor U97 (N_97,In_442,In_1680);
and U98 (N_98,In_230,In_1467);
and U99 (N_99,In_947,In_715);
nand U100 (N_100,In_436,In_1525);
and U101 (N_101,In_915,In_1715);
and U102 (N_102,In_394,In_1755);
nor U103 (N_103,In_932,In_1417);
nand U104 (N_104,In_52,In_1313);
or U105 (N_105,In_1125,In_571);
and U106 (N_106,In_686,In_1581);
xnor U107 (N_107,In_1239,In_541);
and U108 (N_108,In_814,In_103);
or U109 (N_109,In_220,In_1746);
nand U110 (N_110,In_1072,In_1364);
nand U111 (N_111,In_468,In_647);
and U112 (N_112,In_606,In_278);
or U113 (N_113,In_443,In_44);
or U114 (N_114,In_635,In_1835);
and U115 (N_115,In_1808,In_1907);
or U116 (N_116,In_1931,In_41);
or U117 (N_117,In_162,In_54);
xnor U118 (N_118,In_1441,In_1794);
nand U119 (N_119,In_256,In_1093);
nand U120 (N_120,In_1952,In_1545);
or U121 (N_121,In_1906,In_1724);
nor U122 (N_122,In_854,In_354);
nand U123 (N_123,In_254,In_1791);
nor U124 (N_124,In_859,In_543);
nand U125 (N_125,In_1685,In_1628);
and U126 (N_126,In_337,In_517);
nand U127 (N_127,In_794,In_1477);
or U128 (N_128,In_296,In_244);
and U129 (N_129,In_1401,In_1148);
and U130 (N_130,In_1599,In_1922);
or U131 (N_131,In_292,In_960);
or U132 (N_132,In_1918,In_630);
nor U133 (N_133,In_1518,In_1772);
or U134 (N_134,In_1436,In_1524);
xnor U135 (N_135,In_28,In_1109);
or U136 (N_136,In_1040,In_268);
or U137 (N_137,In_929,In_1654);
xor U138 (N_138,In_639,In_309);
or U139 (N_139,In_473,In_853);
or U140 (N_140,In_78,In_1369);
and U141 (N_141,In_1770,In_942);
or U142 (N_142,In_1254,In_1036);
and U143 (N_143,In_1189,In_1964);
xnor U144 (N_144,In_26,In_1265);
or U145 (N_145,In_1886,In_165);
nand U146 (N_146,In_661,In_242);
nor U147 (N_147,In_258,In_1532);
or U148 (N_148,In_1097,In_1065);
xnor U149 (N_149,In_1933,In_1975);
nand U150 (N_150,In_1872,In_1992);
and U151 (N_151,In_1833,In_1634);
nor U152 (N_152,In_1824,In_578);
or U153 (N_153,In_1892,In_625);
nor U154 (N_154,In_1702,In_1807);
xnor U155 (N_155,In_1785,In_1143);
and U156 (N_156,In_707,In_355);
nor U157 (N_157,In_210,In_567);
nor U158 (N_158,In_73,In_1590);
nand U159 (N_159,In_1368,In_95);
or U160 (N_160,In_243,In_48);
or U161 (N_161,In_1676,In_472);
nor U162 (N_162,In_702,In_343);
or U163 (N_163,In_559,In_627);
or U164 (N_164,In_1013,In_1009);
nor U165 (N_165,In_1212,In_1792);
nand U166 (N_166,In_20,In_433);
or U167 (N_167,In_1845,In_514);
nor U168 (N_168,In_581,In_314);
nor U169 (N_169,In_260,In_1767);
xnor U170 (N_170,In_812,In_1472);
or U171 (N_171,In_1819,In_984);
nor U172 (N_172,In_1397,In_594);
and U173 (N_173,In_811,In_1190);
nor U174 (N_174,In_883,In_1086);
nand U175 (N_175,In_677,In_250);
and U176 (N_176,In_275,In_18);
or U177 (N_177,In_922,In_1879);
and U178 (N_178,In_1973,In_1790);
nand U179 (N_179,In_1284,In_1849);
or U180 (N_180,In_1459,In_1078);
and U181 (N_181,In_408,In_213);
and U182 (N_182,In_1388,In_851);
or U183 (N_183,In_1255,In_281);
or U184 (N_184,In_1146,In_1337);
nor U185 (N_185,In_1744,In_323);
and U186 (N_186,In_1237,In_310);
nor U187 (N_187,In_776,In_1990);
nor U188 (N_188,In_266,In_1601);
and U189 (N_189,In_105,In_1057);
xnor U190 (N_190,In_998,In_642);
nor U191 (N_191,In_508,In_848);
nand U192 (N_192,In_36,In_758);
and U193 (N_193,In_1663,In_1410);
and U194 (N_194,In_1298,In_1202);
or U195 (N_195,In_195,In_1652);
nand U196 (N_196,In_1137,In_597);
nor U197 (N_197,In_450,In_456);
or U198 (N_198,In_1623,In_505);
nand U199 (N_199,In_844,In_1111);
and U200 (N_200,In_191,In_1699);
nor U201 (N_201,In_1897,In_1868);
nand U202 (N_202,In_1816,In_1956);
nor U203 (N_203,In_496,In_1540);
or U204 (N_204,In_290,In_1527);
or U205 (N_205,In_1421,In_101);
and U206 (N_206,In_1295,In_1693);
nor U207 (N_207,In_662,In_481);
nor U208 (N_208,In_817,In_1292);
or U209 (N_209,In_1708,In_1025);
and U210 (N_210,In_695,In_312);
nor U211 (N_211,In_828,In_705);
nor U212 (N_212,In_1741,In_1683);
nor U213 (N_213,In_490,In_1187);
nor U214 (N_214,In_1367,In_89);
nor U215 (N_215,In_1324,In_1562);
nand U216 (N_216,In_1998,In_787);
xor U217 (N_217,In_1535,In_1588);
nand U218 (N_218,In_425,In_1035);
or U219 (N_219,In_1616,In_464);
or U220 (N_220,In_93,In_1834);
nand U221 (N_221,In_172,In_1504);
nand U222 (N_222,In_1826,In_1076);
nor U223 (N_223,In_749,In_1804);
xnor U224 (N_224,In_1201,In_923);
or U225 (N_225,In_1555,In_113);
or U226 (N_226,In_525,In_1541);
nand U227 (N_227,In_1806,In_1640);
or U228 (N_228,In_1701,In_1285);
or U229 (N_229,In_196,In_587);
and U230 (N_230,In_1675,In_86);
nor U231 (N_231,In_723,In_1483);
xnor U232 (N_232,In_1249,In_229);
nor U233 (N_233,In_426,In_1739);
xnor U234 (N_234,In_735,In_114);
nand U235 (N_235,In_696,In_1768);
and U236 (N_236,In_768,In_1164);
and U237 (N_237,In_1589,In_1707);
xor U238 (N_238,In_987,In_1711);
xor U239 (N_239,In_1983,In_17);
nand U240 (N_240,In_964,In_423);
nor U241 (N_241,In_142,In_538);
nor U242 (N_242,In_1851,In_1805);
xnor U243 (N_243,In_1920,In_1620);
xor U244 (N_244,In_248,In_1705);
nand U245 (N_245,In_738,In_502);
nor U246 (N_246,In_1979,In_1948);
and U247 (N_247,In_367,In_15);
nand U248 (N_248,In_593,In_1487);
or U249 (N_249,In_1195,In_1902);
nand U250 (N_250,In_1080,In_1729);
nor U251 (N_251,In_907,In_1815);
and U252 (N_252,In_344,In_992);
nor U253 (N_253,In_25,In_1756);
or U254 (N_254,In_1371,In_1618);
xnor U255 (N_255,In_892,In_491);
nand U256 (N_256,In_152,In_219);
or U257 (N_257,In_833,In_1053);
nand U258 (N_258,In_1339,In_1585);
nand U259 (N_259,In_320,In_1012);
nand U260 (N_260,In_1994,In_719);
xor U261 (N_261,In_850,In_1558);
and U262 (N_262,In_34,In_805);
nand U263 (N_263,In_1971,In_1046);
or U264 (N_264,In_839,In_1128);
xnor U265 (N_265,In_373,In_660);
and U266 (N_266,In_346,In_1461);
and U267 (N_267,In_1129,In_1251);
and U268 (N_268,In_236,In_1241);
nand U269 (N_269,In_1084,In_1893);
or U270 (N_270,In_572,In_1611);
nor U271 (N_271,In_9,In_842);
xnor U272 (N_272,In_1393,In_447);
or U273 (N_273,In_1606,In_1801);
and U274 (N_274,In_1232,In_156);
and U275 (N_275,In_1029,In_762);
nand U276 (N_276,In_1380,In_1613);
nor U277 (N_277,In_111,In_398);
or U278 (N_278,In_1912,In_1288);
xor U279 (N_279,In_1553,In_1863);
nand U280 (N_280,In_77,In_382);
nor U281 (N_281,In_322,In_31);
nor U282 (N_282,In_1261,In_318);
nor U283 (N_283,In_670,In_862);
or U284 (N_284,In_743,In_1424);
and U285 (N_285,In_1580,In_1106);
and U286 (N_286,In_937,In_703);
and U287 (N_287,In_353,In_1016);
nor U288 (N_288,In_888,In_1466);
nand U289 (N_289,In_1793,In_1438);
xor U290 (N_290,In_1713,In_834);
nand U291 (N_291,In_1083,In_161);
and U292 (N_292,In_62,In_1965);
xor U293 (N_293,In_1556,In_108);
or U294 (N_294,In_1471,In_465);
nand U295 (N_295,In_1269,In_1276);
nor U296 (N_296,In_1852,In_498);
nor U297 (N_297,In_1329,In_1458);
nor U298 (N_298,In_1810,In_718);
nand U299 (N_299,In_1274,In_1529);
nand U300 (N_300,In_1318,In_1733);
or U301 (N_301,In_1308,In_1206);
or U302 (N_302,In_740,In_876);
or U303 (N_303,In_1655,In_1888);
and U304 (N_304,In_1714,In_712);
nor U305 (N_305,In_413,In_999);
xnor U306 (N_306,In_1330,In_965);
nor U307 (N_307,In_1531,In_956);
nor U308 (N_308,In_793,In_791);
and U309 (N_309,In_1684,In_1592);
and U310 (N_310,In_1864,In_1782);
or U311 (N_311,In_1719,In_225);
and U312 (N_312,In_852,In_1356);
nor U313 (N_313,In_507,In_485);
and U314 (N_314,In_895,In_832);
or U315 (N_315,In_1381,In_1345);
nand U316 (N_316,In_869,In_1048);
and U317 (N_317,In_253,In_1244);
or U318 (N_318,In_1950,In_1862);
nor U319 (N_319,In_282,In_381);
nor U320 (N_320,In_974,In_1386);
and U321 (N_321,In_1412,In_1018);
nor U322 (N_322,In_154,In_887);
nor U323 (N_323,In_1576,In_1697);
and U324 (N_324,In_1473,In_1234);
and U325 (N_325,In_1614,In_591);
or U326 (N_326,In_1115,In_1379);
nand U327 (N_327,In_1814,In_200);
xor U328 (N_328,In_1169,In_430);
and U329 (N_329,In_845,In_1822);
nor U330 (N_330,In_1250,In_1925);
nand U331 (N_331,In_1179,In_342);
nor U332 (N_332,In_1014,In_874);
and U333 (N_333,In_1823,In_400);
or U334 (N_334,In_1947,In_1674);
or U335 (N_335,In_157,In_1252);
nand U336 (N_336,In_837,In_1830);
nor U337 (N_337,In_872,In_1000);
nor U338 (N_338,In_726,In_1342);
nand U339 (N_339,In_1395,In_224);
or U340 (N_340,In_866,In_986);
nand U341 (N_341,In_1796,In_629);
nor U342 (N_342,In_1949,In_451);
xor U343 (N_343,In_1579,In_1268);
or U344 (N_344,In_145,In_378);
or U345 (N_345,In_1905,In_1629);
nand U346 (N_346,In_1737,In_170);
nand U347 (N_347,In_1060,In_1860);
nand U348 (N_348,In_214,In_1856);
or U349 (N_349,In_1131,In_962);
nor U350 (N_350,In_756,In_348);
nand U351 (N_351,In_904,In_72);
nand U352 (N_352,In_305,In_1493);
or U353 (N_353,In_388,In_879);
and U354 (N_354,In_1338,In_1530);
or U355 (N_355,In_1977,In_905);
and U356 (N_356,In_683,In_1134);
nand U357 (N_357,In_1445,In_1390);
nor U358 (N_358,In_1881,In_153);
or U359 (N_359,In_955,In_379);
or U360 (N_360,In_1575,In_1383);
and U361 (N_361,In_1871,In_1229);
nand U362 (N_362,In_1434,In_1891);
nand U363 (N_363,In_1516,In_1709);
nand U364 (N_364,In_1334,In_1070);
and U365 (N_365,In_246,In_434);
nand U366 (N_366,In_1068,In_1615);
nand U367 (N_367,In_1645,In_1821);
nor U368 (N_368,In_445,In_474);
nand U369 (N_369,In_372,In_56);
nor U370 (N_370,In_894,In_429);
nor U371 (N_371,In_422,In_110);
nor U372 (N_372,In_733,In_1866);
nand U373 (N_373,In_1112,In_97);
and U374 (N_374,In_900,In_1802);
xnor U375 (N_375,In_164,In_551);
or U376 (N_376,In_1763,In_1738);
and U377 (N_377,In_1075,In_1132);
or U378 (N_378,In_790,In_390);
nor U379 (N_379,In_147,In_1940);
nand U380 (N_380,In_1923,In_1293);
or U381 (N_381,In_204,In_395);
nand U382 (N_382,In_19,In_494);
and U383 (N_383,In_131,In_1264);
or U384 (N_384,In_1407,In_1362);
and U385 (N_385,In_526,In_35);
nor U386 (N_386,In_133,In_11);
nand U387 (N_387,In_1502,In_865);
and U388 (N_388,In_1139,In_1776);
xor U389 (N_389,In_617,In_226);
nor U390 (N_390,In_1612,In_264);
xor U391 (N_391,In_1761,In_1302);
and U392 (N_392,In_1566,In_1625);
xor U393 (N_393,In_1689,In_401);
nand U394 (N_394,In_51,In_1108);
or U395 (N_395,In_1536,In_1279);
and U396 (N_396,In_637,In_280);
and U397 (N_397,In_1809,In_1695);
or U398 (N_398,In_1153,In_972);
nor U399 (N_399,In_509,In_1389);
nand U400 (N_400,In_163,In_605);
and U401 (N_401,In_857,In_840);
xor U402 (N_402,In_410,In_1160);
nand U403 (N_403,In_1258,In_648);
nand U404 (N_404,In_175,In_1064);
and U405 (N_405,In_1474,In_329);
and U406 (N_406,In_1152,In_149);
xnor U407 (N_407,In_1631,In_469);
nor U408 (N_408,In_1211,In_553);
and U409 (N_409,In_467,In_420);
or U410 (N_410,In_385,In_950);
and U411 (N_411,In_293,In_697);
or U412 (N_412,In_80,In_1091);
nand U413 (N_413,In_138,In_364);
or U414 (N_414,In_979,In_1963);
nor U415 (N_415,In_369,In_16);
nand U416 (N_416,In_774,In_681);
nand U417 (N_417,In_1786,In_462);
and U418 (N_418,In_1098,In_518);
and U419 (N_419,In_1433,In_1089);
or U420 (N_420,In_838,In_92);
nand U421 (N_421,In_1908,In_1100);
xnor U422 (N_422,In_94,In_1681);
nor U423 (N_423,In_1519,In_1119);
nand U424 (N_424,In_1484,In_440);
and U425 (N_425,In_332,In_299);
and U426 (N_426,In_1154,In_554);
xor U427 (N_427,In_3,In_1765);
nand U428 (N_428,In_1133,In_819);
nor U429 (N_429,In_1828,In_1455);
or U430 (N_430,In_1602,In_1398);
nand U431 (N_431,In_565,In_1937);
nand U432 (N_432,In_1451,In_684);
xor U433 (N_433,In_1403,In_653);
and U434 (N_434,In_1846,In_1903);
nor U435 (N_435,In_788,In_1687);
and U436 (N_436,In_980,In_685);
nor U437 (N_437,In_846,In_547);
or U438 (N_438,In_1787,In_522);
and U439 (N_439,In_259,In_1743);
nor U440 (N_440,In_1610,In_1343);
and U441 (N_441,In_1520,In_623);
nor U442 (N_442,In_863,In_1149);
nor U443 (N_443,In_549,In_1372);
and U444 (N_444,In_815,In_598);
nand U445 (N_445,In_1439,In_303);
nand U446 (N_446,In_1120,In_1712);
and U447 (N_447,In_415,In_396);
and U448 (N_448,In_1759,In_217);
xor U449 (N_449,In_796,In_1353);
nand U450 (N_450,In_1151,In_409);
nor U451 (N_451,In_1686,In_1126);
nor U452 (N_452,In_1838,In_452);
nor U453 (N_453,In_1803,In_613);
and U454 (N_454,In_1054,In_669);
xor U455 (N_455,In_933,In_917);
and U456 (N_456,In_1500,In_1989);
nand U457 (N_457,In_1854,In_1305);
nor U458 (N_458,In_143,In_169);
and U459 (N_459,In_125,In_975);
nand U460 (N_460,In_1163,In_656);
or U461 (N_461,In_1314,In_1554);
nand U462 (N_462,In_1557,In_513);
nor U463 (N_463,In_363,In_1257);
xor U464 (N_464,In_804,In_14);
nor U465 (N_465,In_1193,In_1346);
xnor U466 (N_466,In_362,In_1619);
nor U467 (N_467,In_1030,In_1646);
and U468 (N_468,In_1171,In_1385);
and U469 (N_469,In_1736,In_1570);
nand U470 (N_470,In_1883,In_566);
nand U471 (N_471,In_1399,In_173);
and U472 (N_472,In_326,In_29);
and U473 (N_473,In_1262,In_1074);
and U474 (N_474,In_693,In_1569);
or U475 (N_475,In_664,In_1637);
and U476 (N_476,In_1716,In_528);
nand U477 (N_477,In_816,In_539);
or U478 (N_478,In_680,In_1501);
or U479 (N_479,In_941,In_1666);
nand U480 (N_480,In_688,In_978);
nand U481 (N_481,In_1396,In_550);
nor U482 (N_482,In_470,In_1943);
nand U483 (N_483,In_924,In_1114);
nor U484 (N_484,In_878,In_584);
and U485 (N_485,In_1205,In_1621);
nand U486 (N_486,In_1662,In_1374);
or U487 (N_487,In_849,In_1885);
and U488 (N_488,In_1411,In_1188);
nor U489 (N_489,In_759,In_1930);
nand U490 (N_490,In_1118,In_1017);
nor U491 (N_491,In_843,In_1066);
or U492 (N_492,In_564,In_1281);
xor U493 (N_493,In_1058,In_475);
or U494 (N_494,In_760,In_176);
nand U495 (N_495,In_809,In_626);
or U496 (N_496,In_1538,In_728);
or U497 (N_497,In_1568,In_981);
nor U498 (N_498,In_276,In_810);
or U499 (N_499,In_231,In_151);
nor U500 (N_500,In_417,In_1037);
or U501 (N_501,In_1225,In_534);
and U502 (N_502,In_1913,In_1222);
and U503 (N_503,In_1327,In_189);
nor U504 (N_504,In_1726,In_1085);
and U505 (N_505,In_1962,In_1951);
nand U506 (N_506,In_763,In_1218);
xor U507 (N_507,In_1450,In_1231);
and U508 (N_508,In_411,In_504);
and U509 (N_509,In_500,In_731);
nor U510 (N_510,In_595,In_269);
and U511 (N_511,In_1142,In_789);
nand U512 (N_512,In_238,In_1159);
or U513 (N_513,In_1981,In_60);
and U514 (N_514,In_1682,In_1499);
or U515 (N_515,In_335,In_694);
or U516 (N_516,In_1843,In_1968);
and U517 (N_517,In_948,In_199);
nor U518 (N_518,In_1742,In_1422);
or U519 (N_519,In_1464,In_1752);
or U520 (N_520,In_881,In_599);
nand U521 (N_521,In_646,In_1880);
or U522 (N_522,In_159,In_764);
nor U523 (N_523,In_1938,In_383);
nor U524 (N_524,In_1817,In_1443);
nand U525 (N_525,In_993,In_1875);
and U526 (N_526,In_1988,In_610);
or U527 (N_527,In_780,In_137);
and U528 (N_528,In_746,In_1463);
nor U529 (N_529,In_1573,In_1456);
or U530 (N_530,In_333,In_823);
nor U531 (N_531,In_1333,In_1429);
nor U532 (N_532,In_1052,In_1521);
or U533 (N_533,In_120,In_301);
nor U534 (N_534,In_1178,In_1757);
nand U535 (N_535,In_1043,In_813);
or U536 (N_536,In_945,In_577);
nor U537 (N_537,In_1297,In_107);
nand U538 (N_538,In_1384,In_1598);
nand U539 (N_539,In_903,In_1267);
and U540 (N_540,In_1495,In_446);
and U541 (N_541,In_245,In_600);
or U542 (N_542,In_1419,In_512);
xor U543 (N_543,In_1079,In_1336);
and U544 (N_544,In_1526,In_1431);
and U545 (N_545,In_529,In_1415);
nand U546 (N_546,In_666,In_934);
nand U547 (N_547,In_454,In_1023);
or U548 (N_548,In_1186,In_916);
and U549 (N_549,In_966,In_628);
nor U550 (N_550,In_340,In_1972);
xor U551 (N_551,In_1204,In_453);
and U552 (N_552,In_57,In_123);
or U553 (N_553,In_85,In_1350);
or U554 (N_554,In_130,In_1370);
and U555 (N_555,In_555,In_1543);
nand U556 (N_556,In_633,In_418);
nand U557 (N_557,In_701,In_1607);
xor U558 (N_558,In_1180,In_1363);
or U559 (N_559,In_847,In_414);
nor U560 (N_560,In_949,In_1375);
nand U561 (N_561,In_1223,In_1970);
or U562 (N_562,In_1323,In_1004);
xnor U563 (N_563,In_239,In_1319);
or U564 (N_564,In_1270,In_75);
and U565 (N_565,In_675,In_12);
nor U566 (N_566,In_1488,In_608);
nor U567 (N_567,In_463,In_573);
and U568 (N_568,In_586,In_1899);
nor U569 (N_569,In_122,In_1694);
nor U570 (N_570,In_882,In_1764);
and U571 (N_571,In_609,In_1031);
or U572 (N_572,In_1320,In_1812);
nand U573 (N_573,In_1773,In_82);
nand U574 (N_574,In_392,In_925);
xor U575 (N_575,In_255,In_1354);
nand U576 (N_576,In_1315,In_404);
or U577 (N_577,In_1406,In_1081);
nand U578 (N_578,In_1537,In_1196);
nor U579 (N_579,In_61,In_1827);
or U580 (N_580,In_754,In_216);
nor U581 (N_581,In_643,In_546);
or U582 (N_582,In_1498,In_1837);
or U583 (N_583,In_779,In_1976);
xor U584 (N_584,In_1021,In_477);
nor U585 (N_585,In_330,In_1955);
nor U586 (N_586,In_47,In_1656);
nor U587 (N_587,In_1865,In_596);
nand U588 (N_588,In_1428,In_1657);
nand U589 (N_589,In_1028,In_205);
or U590 (N_590,In_1287,In_927);
xnor U591 (N_591,In_771,In_1745);
nand U592 (N_592,In_1392,In_336);
nand U593 (N_593,In_285,In_1939);
or U594 (N_594,In_1507,In_1006);
and U595 (N_595,In_1373,In_1282);
or U596 (N_596,In_687,In_1648);
nand U597 (N_597,In_1564,In_274);
or U598 (N_598,In_1984,In_801);
or U599 (N_599,In_968,In_1780);
xnor U600 (N_600,In_233,In_1565);
nand U601 (N_601,In_188,In_1296);
nor U602 (N_602,In_1515,In_1877);
or U603 (N_603,In_897,In_1199);
nand U604 (N_604,In_339,In_1945);
and U605 (N_605,In_880,In_235);
nor U606 (N_606,In_747,In_289);
and U607 (N_607,In_619,In_1503);
and U608 (N_608,In_757,In_10);
and U609 (N_609,In_424,In_1910);
and U610 (N_610,In_218,In_1476);
or U611 (N_611,In_1095,In_2);
xnor U612 (N_612,In_158,In_1243);
and U613 (N_613,In_1238,In_769);
or U614 (N_614,In_308,In_98);
nor U615 (N_615,In_535,In_87);
xnor U616 (N_616,In_184,In_1460);
nand U617 (N_617,In_1056,In_1283);
nor U618 (N_618,In_1478,In_1);
nand U619 (N_619,In_1760,In_324);
or U620 (N_620,In_1444,In_1929);
or U621 (N_621,In_295,In_352);
nor U622 (N_622,In_83,In_1991);
nor U623 (N_623,In_104,In_1533);
xor U624 (N_624,In_431,In_1107);
nor U625 (N_625,In_338,In_1347);
and U626 (N_626,In_706,In_636);
nand U627 (N_627,In_437,In_1170);
and U628 (N_628,In_1486,In_1003);
nand U629 (N_629,In_674,In_875);
nand U630 (N_630,In_45,In_106);
nor U631 (N_631,In_168,In_1820);
nand U632 (N_632,In_720,In_1550);
and U633 (N_633,In_1266,In_350);
or U634 (N_634,In_926,In_1691);
or U635 (N_635,In_1247,In_722);
nand U636 (N_636,In_1832,In_1150);
nor U637 (N_637,In_615,In_1291);
nand U638 (N_638,In_1007,In_1754);
and U639 (N_639,In_399,In_896);
nor U640 (N_640,In_487,In_770);
or U641 (N_641,In_668,In_1608);
nand U642 (N_642,In_432,In_325);
xor U643 (N_643,In_1033,In_1121);
nor U644 (N_644,In_257,In_1914);
and U645 (N_645,In_112,In_1783);
and U646 (N_646,In_1332,In_806);
and U647 (N_647,In_570,In_313);
and U648 (N_648,In_1099,In_351);
nand U649 (N_649,In_476,In_1194);
and U650 (N_650,In_957,In_824);
nand U651 (N_651,In_752,In_920);
xnor U652 (N_652,In_1894,In_366);
nor U653 (N_653,In_911,In_88);
or U654 (N_654,In_1957,In_304);
xor U655 (N_655,In_969,In_797);
nor U656 (N_656,In_1290,In_117);
or U657 (N_657,In_1214,In_497);
nand U658 (N_658,In_913,In_808);
nor U659 (N_659,In_860,In_141);
xnor U660 (N_660,In_1703,In_709);
nor U661 (N_661,In_994,In_657);
nor U662 (N_662,In_1216,In_65);
or U663 (N_663,In_1174,In_1870);
and U664 (N_664,In_109,In_906);
nor U665 (N_665,In_321,In_341);
or U666 (N_666,In_64,In_1582);
or U667 (N_667,In_265,In_912);
nor U668 (N_668,In_1659,In_22);
and U669 (N_669,In_1122,In_1141);
nand U670 (N_670,In_1758,In_919);
nor U671 (N_671,In_1677,In_1876);
and U672 (N_672,In_1220,In_1465);
nor U673 (N_673,In_1024,In_1272);
nor U674 (N_674,In_1192,In_1996);
or U675 (N_675,In_1839,In_1426);
or U676 (N_676,In_901,In_1026);
nand U677 (N_677,In_1935,In_1479);
nor U678 (N_678,In_0,In_124);
or U679 (N_679,In_365,In_208);
or U680 (N_680,In_1795,In_673);
and U681 (N_681,In_319,In_864);
or U682 (N_682,In_1002,In_1001);
nand U683 (N_683,In_479,In_180);
and U684 (N_684,In_783,In_1440);
or U685 (N_685,In_421,In_84);
nor U686 (N_686,In_1932,In_579);
xnor U687 (N_687,In_777,In_100);
nor U688 (N_688,In_1574,In_102);
xor U689 (N_689,In_822,In_800);
and U690 (N_690,In_284,In_1609);
and U691 (N_691,In_732,In_841);
and U692 (N_692,In_1587,In_391);
and U693 (N_693,In_96,In_370);
and U694 (N_694,In_1489,In_1505);
and U695 (N_695,In_944,In_1145);
or U696 (N_696,In_772,In_1062);
and U697 (N_697,In_622,In_1514);
or U698 (N_698,In_533,In_1413);
nor U699 (N_699,In_1069,In_160);
and U700 (N_700,In_1539,In_1113);
nand U701 (N_701,In_1734,In_374);
nor U702 (N_702,In_345,In_368);
nor U703 (N_703,In_634,In_1067);
nor U704 (N_704,In_263,In_1797);
nor U705 (N_705,In_1140,In_1203);
nand U706 (N_706,In_1563,In_1509);
nor U707 (N_707,In_1221,In_1673);
or U708 (N_708,In_371,In_889);
or U709 (N_709,In_455,In_689);
xnor U710 (N_710,In_651,In_678);
or U711 (N_711,In_1470,In_510);
nor U712 (N_712,In_1061,In_252);
nand U713 (N_713,In_499,In_66);
nor U714 (N_714,In_288,In_1224);
nand U715 (N_715,In_69,In_1092);
or U716 (N_716,In_402,In_377);
nand U717 (N_717,In_985,In_663);
and U718 (N_718,In_1301,In_315);
nand U719 (N_719,In_271,In_270);
and U720 (N_720,In_1022,In_645);
and U721 (N_721,In_294,In_1995);
or U722 (N_722,In_1317,In_692);
or U723 (N_723,In_1546,In_1175);
and U724 (N_724,In_890,In_1316);
nor U725 (N_725,In_982,In_871);
xor U726 (N_726,In_607,In_361);
or U727 (N_727,In_713,In_990);
or U728 (N_728,In_1551,In_1661);
xor U729 (N_729,In_1176,In_439);
nand U730 (N_730,In_931,In_1874);
xnor U731 (N_731,In_190,In_76);
nand U732 (N_732,In_1829,In_1800);
nand U733 (N_733,In_46,In_300);
and U734 (N_734,In_575,In_1015);
or U735 (N_735,In_1191,In_38);
nand U736 (N_736,In_192,In_582);
or U737 (N_737,In_126,In_1032);
nor U738 (N_738,In_412,In_818);
xor U739 (N_739,In_1958,In_976);
or U740 (N_740,In_742,In_803);
or U741 (N_741,In_644,In_973);
nand U742 (N_742,In_995,In_416);
nor U743 (N_743,In_1777,In_1027);
nor U744 (N_744,In_397,In_1781);
nand U745 (N_745,In_283,In_602);
nand U746 (N_746,In_223,In_1242);
and U747 (N_747,In_699,In_428);
or U748 (N_748,In_1969,In_358);
and U749 (N_749,In_1858,In_1926);
nor U750 (N_750,In_1245,In_1130);
nand U751 (N_751,In_1999,In_1359);
and U752 (N_752,In_1647,In_187);
nand U753 (N_753,In_989,In_1304);
nand U754 (N_754,In_1405,In_1993);
and U755 (N_755,In_197,In_1173);
and U756 (N_756,In_716,In_1071);
and U757 (N_757,In_1248,In_466);
and U758 (N_758,In_1762,In_1873);
or U759 (N_759,In_1669,In_1117);
nand U760 (N_760,In_1867,In_936);
nand U761 (N_761,In_721,In_829);
nand U762 (N_762,In_521,In_1414);
nand U763 (N_763,In_1376,In_970);
nand U764 (N_764,In_983,In_542);
xor U765 (N_765,In_1391,In_893);
and U766 (N_766,In_1911,In_24);
nand U767 (N_767,In_1168,In_1485);
nand U768 (N_768,In_316,In_1184);
nand U769 (N_769,In_461,In_5);
or U770 (N_770,In_1209,In_665);
xnor U771 (N_771,In_181,In_222);
or U772 (N_772,In_140,In_1454);
and U773 (N_773,In_262,In_115);
or U774 (N_774,In_1679,In_227);
or U775 (N_775,In_1517,In_1452);
nor U776 (N_776,In_384,In_795);
xor U777 (N_777,In_1506,In_458);
or U778 (N_778,In_958,In_1735);
and U779 (N_779,In_885,In_183);
nand U780 (N_780,In_39,In_272);
nand U781 (N_781,In_1720,In_81);
nand U782 (N_782,In_129,In_785);
nand U783 (N_783,In_182,In_1731);
or U784 (N_784,In_202,In_1462);
nand U785 (N_785,In_1352,In_232);
and U786 (N_786,In_42,In_1124);
nand U787 (N_787,In_493,In_1560);
nand U788 (N_788,In_1627,In_1664);
nor U789 (N_789,In_1895,In_1289);
nand U790 (N_790,In_127,In_349);
or U791 (N_791,In_1901,In_1378);
nand U792 (N_792,In_389,In_727);
or U793 (N_793,In_1321,In_1260);
and U794 (N_794,In_952,In_91);
and U795 (N_795,In_909,In_441);
or U796 (N_796,In_714,In_641);
xor U797 (N_797,In_55,In_618);
and U798 (N_798,In_1200,In_1197);
nand U799 (N_799,In_1960,In_1548);
or U800 (N_800,In_908,In_506);
xnor U801 (N_801,In_1402,In_1528);
or U802 (N_802,In_1299,In_1087);
xor U803 (N_803,In_1335,In_1135);
or U804 (N_804,In_1425,In_899);
xnor U805 (N_805,In_495,In_1273);
nor U806 (N_806,In_511,In_1857);
xor U807 (N_807,In_1181,In_1889);
or U808 (N_808,In_516,In_1980);
or U809 (N_809,In_1365,In_386);
xor U810 (N_810,In_1811,In_174);
or U811 (N_811,In_1348,In_1309);
or U812 (N_812,In_484,In_1102);
nor U813 (N_813,In_638,In_116);
or U814 (N_814,In_1340,In_1959);
and U815 (N_815,In_311,In_1446);
nor U816 (N_816,In_1047,In_21);
nand U817 (N_817,In_1219,In_977);
and U818 (N_818,In_136,In_1358);
nand U819 (N_819,In_1966,In_1059);
and U820 (N_820,In_68,In_1447);
xor U821 (N_821,In_667,In_1482);
nand U822 (N_822,In_1670,In_483);
nand U823 (N_823,In_856,In_30);
or U824 (N_824,In_1011,In_375);
nor U825 (N_825,In_380,In_1432);
nand U826 (N_826,In_1855,In_1660);
or U827 (N_827,In_1740,In_741);
and U828 (N_828,In_1377,In_691);
and U829 (N_829,In_1721,In_1700);
or U830 (N_830,In_376,In_1942);
or U831 (N_831,In_1020,In_569);
and U832 (N_832,In_1228,In_1909);
and U833 (N_833,In_1617,In_1355);
or U834 (N_834,In_548,In_1496);
nand U835 (N_835,In_825,In_1158);
nor U836 (N_836,In_1718,In_1847);
nand U837 (N_837,In_682,In_614);
nor U838 (N_838,In_1921,In_951);
and U839 (N_839,In_870,In_459);
nor U840 (N_840,In_448,In_1723);
or U841 (N_841,In_918,In_700);
nor U842 (N_842,In_407,In_279);
nor U843 (N_843,In_1936,In_1658);
nand U844 (N_844,In_13,In_1577);
nand U845 (N_845,In_1161,In_267);
nor U846 (N_846,In_1307,In_4);
and U847 (N_847,In_734,In_940);
nand U848 (N_848,In_1898,In_1751);
or U849 (N_849,In_1642,In_576);
and U850 (N_850,In_939,In_1924);
or U851 (N_851,In_781,In_724);
or U852 (N_852,In_1127,In_1357);
and U853 (N_853,In_1050,In_778);
and U854 (N_854,In_1394,In_1110);
or U855 (N_855,In_273,In_659);
xor U856 (N_856,In_1511,In_1051);
and U857 (N_857,In_967,In_1696);
nand U858 (N_858,In_671,In_1138);
or U859 (N_859,In_1725,In_1271);
or U860 (N_860,In_1753,In_1987);
nand U861 (N_861,In_387,In_1600);
or U862 (N_862,In_1692,In_460);
xnor U863 (N_863,In_1344,In_1917);
and U864 (N_864,In_676,In_1986);
or U865 (N_865,In_855,In_1286);
nand U866 (N_866,In_1144,In_1280);
nor U867 (N_867,In_1005,In_1088);
nor U868 (N_868,In_482,In_560);
nand U869 (N_869,In_90,In_1312);
and U870 (N_870,In_1182,In_277);
nand U871 (N_871,In_1594,In_1449);
nand U872 (N_872,In_827,In_1878);
and U873 (N_873,In_1259,In_167);
nand U874 (N_874,In_963,In_203);
or U875 (N_875,In_58,In_524);
nand U876 (N_876,In_1861,In_1325);
and U877 (N_877,In_298,In_1094);
nor U878 (N_878,In_959,In_604);
nor U879 (N_879,In_121,In_1636);
nor U880 (N_880,In_938,In_603);
nor U881 (N_881,In_574,In_658);
and U882 (N_882,In_171,In_1256);
or U883 (N_883,In_331,In_1974);
or U884 (N_884,In_43,In_1233);
or U885 (N_885,In_1213,In_1039);
nor U886 (N_886,In_921,In_826);
and U887 (N_887,In_37,In_1105);
or U888 (N_888,In_632,In_1073);
or U889 (N_889,In_59,In_902);
nand U890 (N_890,In_946,In_419);
nor U891 (N_891,In_1277,In_1448);
and U892 (N_892,In_868,In_1322);
xnor U893 (N_893,In_1435,In_1633);
nor U894 (N_894,In_1710,In_1423);
or U895 (N_895,In_640,In_1185);
and U896 (N_896,In_1055,In_520);
or U897 (N_897,In_690,In_356);
or U898 (N_898,In_1722,In_261);
or U899 (N_899,In_1732,In_1166);
and U900 (N_900,In_562,In_654);
or U901 (N_901,In_580,In_1162);
and U902 (N_902,In_1583,In_1717);
and U903 (N_903,In_861,In_7);
or U904 (N_904,In_1491,In_119);
or U905 (N_905,In_1215,In_1798);
and U906 (N_906,In_820,In_53);
or U907 (N_907,In_1207,In_1306);
or U908 (N_908,In_997,In_744);
or U909 (N_909,In_592,In_1552);
nor U910 (N_910,In_1420,In_589);
or U911 (N_911,In_1690,In_70);
nand U912 (N_912,In_710,In_798);
nand U913 (N_913,In_1430,In_1915);
or U914 (N_914,In_1400,In_537);
nand U915 (N_915,In_1236,In_1927);
nor U916 (N_916,In_858,In_556);
nor U917 (N_917,In_1813,In_1508);
nor U918 (N_918,In_884,In_457);
nor U919 (N_919,In_1978,In_530);
or U920 (N_920,In_655,In_148);
or U921 (N_921,In_1853,In_118);
and U922 (N_922,In_954,In_1008);
nand U923 (N_923,In_1671,In_1019);
xor U924 (N_924,In_1789,In_782);
nor U925 (N_925,In_194,In_792);
xor U926 (N_926,In_489,In_1300);
or U927 (N_927,In_1263,In_71);
xor U928 (N_928,In_27,In_1635);
nor U929 (N_929,In_211,In_1457);
nor U930 (N_930,In_914,In_1572);
nor U931 (N_931,In_286,In_1240);
or U932 (N_932,In_135,In_953);
nor U933 (N_933,In_765,In_561);
nand U934 (N_934,In_1961,In_212);
nor U935 (N_935,In_1561,In_1571);
xnor U936 (N_936,In_1494,In_1678);
nor U937 (N_937,In_1591,In_23);
nor U938 (N_938,In_935,In_237);
nand U939 (N_939,In_488,In_1638);
nor U940 (N_940,In_438,In_784);
nor U941 (N_941,In_1230,In_1123);
nor U942 (N_942,In_444,In_544);
or U943 (N_943,In_1596,In_698);
and U944 (N_944,In_1941,In_585);
nand U945 (N_945,In_79,In_652);
and U946 (N_946,In_590,In_988);
or U947 (N_947,In_1630,In_247);
nor U948 (N_948,In_568,In_307);
xnor U949 (N_949,In_631,In_207);
nor U950 (N_950,In_1512,In_1626);
and U951 (N_951,In_1351,In_178);
xnor U952 (N_952,In_139,In_1844);
nor U953 (N_953,In_1750,In_405);
xor U954 (N_954,In_1157,In_63);
nor U955 (N_955,In_1859,In_519);
nand U956 (N_956,In_611,In_1727);
xor U957 (N_957,In_1522,In_1542);
nand U958 (N_958,In_501,In_1644);
nor U959 (N_959,In_206,In_1404);
xnor U960 (N_960,In_1641,In_1490);
and U961 (N_961,In_961,In_1706);
and U962 (N_962,In_1492,In_359);
nor U963 (N_963,In_134,In_1887);
or U964 (N_964,In_1632,In_1586);
or U965 (N_965,In_1165,In_1919);
nand U966 (N_966,In_1044,In_302);
xnor U967 (N_967,In_1328,In_786);
or U968 (N_968,In_1469,In_471);
and U969 (N_969,In_1649,In_1842);
or U970 (N_970,In_144,In_1534);
or U971 (N_971,In_1653,In_1341);
and U972 (N_972,In_287,In_1704);
or U973 (N_973,In_1217,In_1041);
and U974 (N_974,In_1604,In_836);
nand U975 (N_975,In_449,In_1310);
xor U976 (N_976,In_6,In_74);
and U977 (N_977,In_748,In_991);
nor U978 (N_978,In_1418,In_251);
nand U979 (N_979,In_50,In_877);
nand U980 (N_980,In_650,In_745);
nor U981 (N_981,In_132,In_1235);
or U982 (N_982,In_393,In_360);
nand U983 (N_983,In_971,In_1953);
and U984 (N_984,In_1766,In_1038);
nand U985 (N_985,In_1698,In_1818);
nor U986 (N_986,In_1567,In_1481);
and U987 (N_987,In_1303,In_910);
nor U988 (N_988,In_679,In_807);
nand U989 (N_989,In_1788,In_435);
nor U990 (N_990,In_1779,In_1077);
or U991 (N_991,In_49,In_1836);
xor U992 (N_992,In_1595,In_1825);
and U993 (N_993,In_750,In_1116);
or U994 (N_994,In_1728,In_1101);
or U995 (N_995,In_711,In_1639);
and U996 (N_996,In_620,In_478);
or U997 (N_997,In_1622,In_1523);
or U998 (N_998,In_1437,In_1442);
and U999 (N_999,In_406,In_327);
xnor U1000 (N_1000,In_818,In_1143);
and U1001 (N_1001,In_1926,In_1702);
nand U1002 (N_1002,In_179,In_1622);
nor U1003 (N_1003,In_431,In_675);
or U1004 (N_1004,In_798,In_624);
or U1005 (N_1005,In_900,In_139);
and U1006 (N_1006,In_665,In_1514);
nand U1007 (N_1007,In_571,In_1307);
nor U1008 (N_1008,In_473,In_1550);
xnor U1009 (N_1009,In_1612,In_403);
and U1010 (N_1010,In_335,In_1570);
nor U1011 (N_1011,In_182,In_256);
nand U1012 (N_1012,In_1815,In_1797);
nor U1013 (N_1013,In_178,In_1119);
and U1014 (N_1014,In_1807,In_1612);
or U1015 (N_1015,In_1920,In_147);
xnor U1016 (N_1016,In_124,In_1898);
nor U1017 (N_1017,In_888,In_1519);
nand U1018 (N_1018,In_1328,In_58);
nor U1019 (N_1019,In_1732,In_458);
or U1020 (N_1020,In_1853,In_479);
xor U1021 (N_1021,In_1801,In_617);
xor U1022 (N_1022,In_98,In_1787);
and U1023 (N_1023,In_689,In_1131);
or U1024 (N_1024,In_1596,In_1020);
nor U1025 (N_1025,In_868,In_1689);
nor U1026 (N_1026,In_33,In_37);
nand U1027 (N_1027,In_1949,In_751);
xnor U1028 (N_1028,In_232,In_24);
nand U1029 (N_1029,In_756,In_739);
nand U1030 (N_1030,In_1998,In_1446);
and U1031 (N_1031,In_1306,In_989);
nor U1032 (N_1032,In_1391,In_51);
nand U1033 (N_1033,In_667,In_202);
or U1034 (N_1034,In_1659,In_1105);
nor U1035 (N_1035,In_598,In_769);
xor U1036 (N_1036,In_1781,In_1281);
or U1037 (N_1037,In_1863,In_1133);
and U1038 (N_1038,In_1496,In_1773);
and U1039 (N_1039,In_1143,In_603);
or U1040 (N_1040,In_1828,In_801);
nand U1041 (N_1041,In_840,In_290);
nor U1042 (N_1042,In_200,In_816);
xnor U1043 (N_1043,In_1227,In_1498);
xor U1044 (N_1044,In_7,In_1814);
or U1045 (N_1045,In_259,In_467);
nor U1046 (N_1046,In_189,In_51);
or U1047 (N_1047,In_583,In_82);
or U1048 (N_1048,In_1398,In_199);
nor U1049 (N_1049,In_1019,In_24);
nand U1050 (N_1050,In_1690,In_1543);
xor U1051 (N_1051,In_367,In_27);
and U1052 (N_1052,In_460,In_1564);
or U1053 (N_1053,In_1217,In_1348);
nand U1054 (N_1054,In_1231,In_16);
xor U1055 (N_1055,In_598,In_874);
nand U1056 (N_1056,In_1777,In_1989);
or U1057 (N_1057,In_525,In_98);
nand U1058 (N_1058,In_1926,In_1852);
nand U1059 (N_1059,In_1648,In_1616);
and U1060 (N_1060,In_1465,In_59);
or U1061 (N_1061,In_1080,In_745);
or U1062 (N_1062,In_1778,In_119);
and U1063 (N_1063,In_1721,In_1846);
nor U1064 (N_1064,In_1024,In_1041);
and U1065 (N_1065,In_524,In_586);
nand U1066 (N_1066,In_774,In_357);
xor U1067 (N_1067,In_1480,In_1251);
nand U1068 (N_1068,In_1011,In_13);
xor U1069 (N_1069,In_1084,In_872);
or U1070 (N_1070,In_1088,In_1075);
and U1071 (N_1071,In_913,In_39);
nor U1072 (N_1072,In_188,In_1761);
and U1073 (N_1073,In_880,In_441);
or U1074 (N_1074,In_1508,In_220);
nor U1075 (N_1075,In_169,In_1374);
xnor U1076 (N_1076,In_863,In_1367);
nor U1077 (N_1077,In_1457,In_490);
xor U1078 (N_1078,In_1134,In_708);
nor U1079 (N_1079,In_1149,In_1346);
and U1080 (N_1080,In_1239,In_1136);
or U1081 (N_1081,In_504,In_1654);
or U1082 (N_1082,In_1841,In_1564);
nor U1083 (N_1083,In_1241,In_577);
or U1084 (N_1084,In_450,In_484);
nor U1085 (N_1085,In_1297,In_605);
xor U1086 (N_1086,In_1815,In_735);
nand U1087 (N_1087,In_1470,In_291);
nor U1088 (N_1088,In_1807,In_1390);
and U1089 (N_1089,In_1800,In_606);
or U1090 (N_1090,In_1020,In_31);
nand U1091 (N_1091,In_726,In_772);
or U1092 (N_1092,In_99,In_1288);
xnor U1093 (N_1093,In_898,In_1418);
and U1094 (N_1094,In_704,In_332);
or U1095 (N_1095,In_881,In_1828);
and U1096 (N_1096,In_217,In_9);
or U1097 (N_1097,In_1540,In_1515);
nand U1098 (N_1098,In_536,In_1749);
nor U1099 (N_1099,In_1486,In_118);
nand U1100 (N_1100,In_9,In_1957);
xnor U1101 (N_1101,In_1190,In_22);
nand U1102 (N_1102,In_1855,In_561);
nor U1103 (N_1103,In_1178,In_597);
nor U1104 (N_1104,In_1275,In_1524);
nor U1105 (N_1105,In_881,In_1802);
nand U1106 (N_1106,In_1615,In_1275);
and U1107 (N_1107,In_1219,In_1108);
nor U1108 (N_1108,In_1552,In_1748);
nor U1109 (N_1109,In_305,In_515);
or U1110 (N_1110,In_1051,In_1549);
xor U1111 (N_1111,In_1657,In_829);
and U1112 (N_1112,In_888,In_1048);
or U1113 (N_1113,In_1756,In_1339);
or U1114 (N_1114,In_747,In_1820);
or U1115 (N_1115,In_707,In_1815);
nor U1116 (N_1116,In_691,In_637);
nor U1117 (N_1117,In_82,In_1238);
nor U1118 (N_1118,In_1744,In_853);
xnor U1119 (N_1119,In_1779,In_1076);
or U1120 (N_1120,In_365,In_995);
nor U1121 (N_1121,In_1331,In_607);
and U1122 (N_1122,In_958,In_1676);
xnor U1123 (N_1123,In_433,In_1773);
and U1124 (N_1124,In_1877,In_1919);
and U1125 (N_1125,In_1580,In_119);
nor U1126 (N_1126,In_368,In_1306);
nor U1127 (N_1127,In_1221,In_1938);
or U1128 (N_1128,In_1544,In_1656);
or U1129 (N_1129,In_540,In_103);
nand U1130 (N_1130,In_1393,In_215);
nand U1131 (N_1131,In_1875,In_1623);
nand U1132 (N_1132,In_326,In_1026);
or U1133 (N_1133,In_1103,In_63);
nor U1134 (N_1134,In_620,In_364);
or U1135 (N_1135,In_1953,In_1538);
and U1136 (N_1136,In_140,In_424);
and U1137 (N_1137,In_1926,In_1915);
nor U1138 (N_1138,In_1731,In_1680);
nand U1139 (N_1139,In_1603,In_754);
and U1140 (N_1140,In_91,In_1526);
or U1141 (N_1141,In_34,In_1826);
or U1142 (N_1142,In_196,In_21);
nor U1143 (N_1143,In_936,In_1419);
nor U1144 (N_1144,In_1632,In_967);
and U1145 (N_1145,In_1001,In_1515);
xor U1146 (N_1146,In_47,In_1853);
nor U1147 (N_1147,In_1149,In_202);
nor U1148 (N_1148,In_1138,In_313);
or U1149 (N_1149,In_344,In_457);
nand U1150 (N_1150,In_931,In_1866);
xnor U1151 (N_1151,In_242,In_105);
or U1152 (N_1152,In_335,In_569);
and U1153 (N_1153,In_1561,In_492);
nor U1154 (N_1154,In_315,In_653);
nand U1155 (N_1155,In_1852,In_255);
nand U1156 (N_1156,In_661,In_688);
and U1157 (N_1157,In_1710,In_1363);
nand U1158 (N_1158,In_1775,In_1023);
xor U1159 (N_1159,In_324,In_751);
or U1160 (N_1160,In_1118,In_399);
or U1161 (N_1161,In_485,In_1744);
nor U1162 (N_1162,In_262,In_277);
xor U1163 (N_1163,In_1087,In_1047);
or U1164 (N_1164,In_192,In_1706);
or U1165 (N_1165,In_931,In_279);
xor U1166 (N_1166,In_949,In_456);
nor U1167 (N_1167,In_1429,In_292);
or U1168 (N_1168,In_505,In_367);
nand U1169 (N_1169,In_1326,In_1767);
nor U1170 (N_1170,In_548,In_1001);
or U1171 (N_1171,In_901,In_1652);
nand U1172 (N_1172,In_962,In_178);
and U1173 (N_1173,In_1829,In_1132);
nand U1174 (N_1174,In_334,In_338);
and U1175 (N_1175,In_1195,In_1506);
nor U1176 (N_1176,In_976,In_759);
and U1177 (N_1177,In_660,In_540);
or U1178 (N_1178,In_1670,In_1865);
nor U1179 (N_1179,In_1010,In_386);
nand U1180 (N_1180,In_1825,In_1070);
nand U1181 (N_1181,In_1179,In_963);
or U1182 (N_1182,In_18,In_465);
or U1183 (N_1183,In_237,In_1808);
or U1184 (N_1184,In_633,In_81);
xnor U1185 (N_1185,In_352,In_345);
nand U1186 (N_1186,In_118,In_964);
or U1187 (N_1187,In_1235,In_809);
and U1188 (N_1188,In_478,In_1443);
and U1189 (N_1189,In_1221,In_371);
or U1190 (N_1190,In_740,In_469);
or U1191 (N_1191,In_890,In_875);
and U1192 (N_1192,In_10,In_1120);
nor U1193 (N_1193,In_334,In_1834);
and U1194 (N_1194,In_972,In_1804);
or U1195 (N_1195,In_1470,In_1779);
nor U1196 (N_1196,In_1111,In_811);
nor U1197 (N_1197,In_979,In_373);
nand U1198 (N_1198,In_157,In_778);
or U1199 (N_1199,In_982,In_800);
or U1200 (N_1200,In_1637,In_517);
nor U1201 (N_1201,In_1625,In_47);
or U1202 (N_1202,In_1026,In_840);
nand U1203 (N_1203,In_285,In_1726);
nand U1204 (N_1204,In_979,In_0);
and U1205 (N_1205,In_16,In_225);
or U1206 (N_1206,In_889,In_1638);
and U1207 (N_1207,In_1438,In_773);
nand U1208 (N_1208,In_157,In_1541);
nor U1209 (N_1209,In_987,In_245);
or U1210 (N_1210,In_931,In_837);
or U1211 (N_1211,In_873,In_1288);
or U1212 (N_1212,In_1666,In_833);
or U1213 (N_1213,In_1700,In_593);
nand U1214 (N_1214,In_1546,In_1086);
and U1215 (N_1215,In_1602,In_1917);
and U1216 (N_1216,In_766,In_1393);
or U1217 (N_1217,In_457,In_906);
xnor U1218 (N_1218,In_892,In_1475);
nor U1219 (N_1219,In_251,In_62);
nor U1220 (N_1220,In_1382,In_157);
nor U1221 (N_1221,In_1278,In_955);
and U1222 (N_1222,In_568,In_240);
xnor U1223 (N_1223,In_1259,In_1127);
and U1224 (N_1224,In_1913,In_14);
and U1225 (N_1225,In_1114,In_378);
and U1226 (N_1226,In_1124,In_930);
or U1227 (N_1227,In_1953,In_719);
and U1228 (N_1228,In_786,In_624);
nand U1229 (N_1229,In_1424,In_1893);
or U1230 (N_1230,In_1477,In_1685);
nor U1231 (N_1231,In_137,In_1662);
nor U1232 (N_1232,In_393,In_373);
nand U1233 (N_1233,In_978,In_1723);
nor U1234 (N_1234,In_84,In_1338);
xnor U1235 (N_1235,In_631,In_811);
and U1236 (N_1236,In_1425,In_1488);
nor U1237 (N_1237,In_934,In_1640);
or U1238 (N_1238,In_951,In_760);
nand U1239 (N_1239,In_1407,In_736);
and U1240 (N_1240,In_1221,In_520);
or U1241 (N_1241,In_1465,In_1009);
nand U1242 (N_1242,In_1402,In_1275);
nand U1243 (N_1243,In_1810,In_1929);
and U1244 (N_1244,In_1893,In_701);
and U1245 (N_1245,In_449,In_371);
or U1246 (N_1246,In_976,In_389);
nand U1247 (N_1247,In_1264,In_1299);
or U1248 (N_1248,In_836,In_1246);
nor U1249 (N_1249,In_1897,In_1109);
xor U1250 (N_1250,In_1738,In_179);
xor U1251 (N_1251,In_709,In_1191);
nand U1252 (N_1252,In_1450,In_1012);
nor U1253 (N_1253,In_1496,In_1127);
nor U1254 (N_1254,In_1918,In_1415);
or U1255 (N_1255,In_71,In_45);
nor U1256 (N_1256,In_1025,In_888);
nor U1257 (N_1257,In_1448,In_561);
nor U1258 (N_1258,In_178,In_610);
or U1259 (N_1259,In_45,In_1220);
or U1260 (N_1260,In_1667,In_1377);
or U1261 (N_1261,In_1244,In_851);
nand U1262 (N_1262,In_984,In_1433);
or U1263 (N_1263,In_854,In_743);
nand U1264 (N_1264,In_1495,In_874);
nand U1265 (N_1265,In_1724,In_1829);
nor U1266 (N_1266,In_581,In_1705);
nor U1267 (N_1267,In_418,In_1918);
or U1268 (N_1268,In_1439,In_76);
nand U1269 (N_1269,In_30,In_330);
or U1270 (N_1270,In_1113,In_1845);
nand U1271 (N_1271,In_1911,In_157);
and U1272 (N_1272,In_413,In_1249);
and U1273 (N_1273,In_388,In_575);
nand U1274 (N_1274,In_1268,In_33);
nand U1275 (N_1275,In_1818,In_1820);
nor U1276 (N_1276,In_1978,In_1304);
and U1277 (N_1277,In_1341,In_883);
nand U1278 (N_1278,In_141,In_650);
nor U1279 (N_1279,In_1946,In_732);
nand U1280 (N_1280,In_1764,In_1318);
nor U1281 (N_1281,In_175,In_1662);
nand U1282 (N_1282,In_1729,In_1762);
and U1283 (N_1283,In_529,In_231);
nand U1284 (N_1284,In_1046,In_1461);
and U1285 (N_1285,In_745,In_1422);
or U1286 (N_1286,In_446,In_1748);
nand U1287 (N_1287,In_127,In_539);
and U1288 (N_1288,In_1523,In_1903);
nand U1289 (N_1289,In_953,In_1440);
nor U1290 (N_1290,In_1439,In_64);
nor U1291 (N_1291,In_679,In_398);
or U1292 (N_1292,In_1206,In_1279);
nor U1293 (N_1293,In_760,In_879);
and U1294 (N_1294,In_876,In_102);
nor U1295 (N_1295,In_809,In_1553);
and U1296 (N_1296,In_1438,In_37);
and U1297 (N_1297,In_1734,In_1569);
or U1298 (N_1298,In_1221,In_1005);
and U1299 (N_1299,In_415,In_972);
nor U1300 (N_1300,In_671,In_1657);
nand U1301 (N_1301,In_410,In_1029);
or U1302 (N_1302,In_376,In_1617);
and U1303 (N_1303,In_1081,In_72);
nor U1304 (N_1304,In_191,In_189);
nor U1305 (N_1305,In_532,In_678);
nand U1306 (N_1306,In_75,In_1677);
xor U1307 (N_1307,In_824,In_1208);
and U1308 (N_1308,In_304,In_868);
nand U1309 (N_1309,In_694,In_1791);
or U1310 (N_1310,In_1563,In_1273);
nand U1311 (N_1311,In_1454,In_90);
and U1312 (N_1312,In_483,In_1001);
or U1313 (N_1313,In_1896,In_1622);
nand U1314 (N_1314,In_1955,In_19);
or U1315 (N_1315,In_1313,In_983);
or U1316 (N_1316,In_694,In_1820);
nand U1317 (N_1317,In_1430,In_1663);
nor U1318 (N_1318,In_474,In_148);
and U1319 (N_1319,In_1040,In_1116);
nor U1320 (N_1320,In_791,In_774);
nor U1321 (N_1321,In_1628,In_1641);
xor U1322 (N_1322,In_638,In_114);
nand U1323 (N_1323,In_1897,In_654);
nand U1324 (N_1324,In_968,In_738);
nor U1325 (N_1325,In_340,In_1792);
or U1326 (N_1326,In_699,In_239);
and U1327 (N_1327,In_963,In_877);
nand U1328 (N_1328,In_127,In_403);
nor U1329 (N_1329,In_1111,In_964);
and U1330 (N_1330,In_616,In_898);
and U1331 (N_1331,In_1176,In_762);
xor U1332 (N_1332,In_499,In_24);
nand U1333 (N_1333,In_1367,In_390);
nand U1334 (N_1334,In_934,In_963);
nand U1335 (N_1335,In_1140,In_1601);
xor U1336 (N_1336,In_1201,In_151);
nor U1337 (N_1337,In_1230,In_385);
or U1338 (N_1338,In_1272,In_1759);
nor U1339 (N_1339,In_1202,In_847);
nor U1340 (N_1340,In_667,In_1065);
nand U1341 (N_1341,In_306,In_1801);
or U1342 (N_1342,In_377,In_1435);
nor U1343 (N_1343,In_161,In_547);
nor U1344 (N_1344,In_1727,In_932);
nand U1345 (N_1345,In_1211,In_812);
and U1346 (N_1346,In_1073,In_777);
or U1347 (N_1347,In_1632,In_1980);
or U1348 (N_1348,In_984,In_1114);
nand U1349 (N_1349,In_1008,In_504);
or U1350 (N_1350,In_277,In_1251);
or U1351 (N_1351,In_1513,In_230);
nand U1352 (N_1352,In_1259,In_352);
and U1353 (N_1353,In_15,In_435);
or U1354 (N_1354,In_678,In_754);
xnor U1355 (N_1355,In_1633,In_166);
nand U1356 (N_1356,In_484,In_210);
nor U1357 (N_1357,In_625,In_1759);
nand U1358 (N_1358,In_230,In_1006);
and U1359 (N_1359,In_645,In_496);
nor U1360 (N_1360,In_1234,In_1702);
and U1361 (N_1361,In_742,In_614);
or U1362 (N_1362,In_1689,In_1313);
and U1363 (N_1363,In_154,In_1970);
nand U1364 (N_1364,In_705,In_1365);
xor U1365 (N_1365,In_1549,In_848);
xnor U1366 (N_1366,In_1045,In_82);
xor U1367 (N_1367,In_1759,In_1161);
or U1368 (N_1368,In_1440,In_1750);
or U1369 (N_1369,In_411,In_260);
and U1370 (N_1370,In_1716,In_678);
or U1371 (N_1371,In_1645,In_1011);
nand U1372 (N_1372,In_112,In_412);
and U1373 (N_1373,In_714,In_81);
or U1374 (N_1374,In_17,In_1694);
or U1375 (N_1375,In_1339,In_1836);
and U1376 (N_1376,In_1513,In_784);
nand U1377 (N_1377,In_1572,In_678);
and U1378 (N_1378,In_1382,In_989);
nor U1379 (N_1379,In_613,In_1412);
and U1380 (N_1380,In_1624,In_1768);
or U1381 (N_1381,In_1897,In_614);
nand U1382 (N_1382,In_1892,In_117);
or U1383 (N_1383,In_1344,In_53);
nor U1384 (N_1384,In_1010,In_1348);
xor U1385 (N_1385,In_849,In_644);
nor U1386 (N_1386,In_1073,In_1417);
nand U1387 (N_1387,In_1570,In_1946);
nand U1388 (N_1388,In_885,In_609);
nor U1389 (N_1389,In_1113,In_876);
nor U1390 (N_1390,In_737,In_1102);
nor U1391 (N_1391,In_1279,In_196);
and U1392 (N_1392,In_157,In_549);
nor U1393 (N_1393,In_1476,In_916);
nor U1394 (N_1394,In_575,In_415);
or U1395 (N_1395,In_1111,In_821);
nand U1396 (N_1396,In_888,In_1470);
nand U1397 (N_1397,In_657,In_1524);
or U1398 (N_1398,In_545,In_495);
and U1399 (N_1399,In_562,In_1082);
nor U1400 (N_1400,In_1628,In_1501);
or U1401 (N_1401,In_93,In_1823);
and U1402 (N_1402,In_842,In_511);
nand U1403 (N_1403,In_1117,In_190);
nand U1404 (N_1404,In_656,In_897);
or U1405 (N_1405,In_1738,In_1906);
or U1406 (N_1406,In_1551,In_557);
nor U1407 (N_1407,In_1973,In_683);
or U1408 (N_1408,In_1141,In_1175);
xor U1409 (N_1409,In_1677,In_1674);
nor U1410 (N_1410,In_1752,In_947);
and U1411 (N_1411,In_1614,In_1382);
and U1412 (N_1412,In_177,In_644);
nand U1413 (N_1413,In_1196,In_357);
nor U1414 (N_1414,In_748,In_1832);
and U1415 (N_1415,In_1028,In_688);
nand U1416 (N_1416,In_772,In_1030);
nand U1417 (N_1417,In_1493,In_91);
nor U1418 (N_1418,In_725,In_1421);
and U1419 (N_1419,In_155,In_63);
or U1420 (N_1420,In_171,In_119);
nand U1421 (N_1421,In_542,In_1912);
or U1422 (N_1422,In_1667,In_507);
and U1423 (N_1423,In_1345,In_885);
nor U1424 (N_1424,In_1031,In_502);
nand U1425 (N_1425,In_1155,In_919);
xor U1426 (N_1426,In_515,In_723);
nor U1427 (N_1427,In_1392,In_557);
nor U1428 (N_1428,In_315,In_343);
or U1429 (N_1429,In_1846,In_480);
xnor U1430 (N_1430,In_256,In_1919);
and U1431 (N_1431,In_730,In_638);
nor U1432 (N_1432,In_1665,In_1713);
or U1433 (N_1433,In_339,In_249);
nor U1434 (N_1434,In_512,In_917);
and U1435 (N_1435,In_690,In_1840);
nor U1436 (N_1436,In_183,In_56);
or U1437 (N_1437,In_1767,In_1011);
nor U1438 (N_1438,In_378,In_1154);
nor U1439 (N_1439,In_1618,In_971);
or U1440 (N_1440,In_565,In_856);
nor U1441 (N_1441,In_1743,In_1751);
nand U1442 (N_1442,In_1985,In_491);
and U1443 (N_1443,In_1836,In_1459);
and U1444 (N_1444,In_1123,In_493);
xnor U1445 (N_1445,In_108,In_400);
and U1446 (N_1446,In_1430,In_713);
nor U1447 (N_1447,In_694,In_1571);
nor U1448 (N_1448,In_1564,In_1199);
nor U1449 (N_1449,In_1660,In_1455);
and U1450 (N_1450,In_966,In_1951);
nand U1451 (N_1451,In_1720,In_1310);
xnor U1452 (N_1452,In_774,In_1396);
and U1453 (N_1453,In_173,In_1720);
nand U1454 (N_1454,In_124,In_1968);
and U1455 (N_1455,In_1982,In_1135);
nor U1456 (N_1456,In_801,In_1526);
nor U1457 (N_1457,In_1974,In_121);
and U1458 (N_1458,In_273,In_777);
nand U1459 (N_1459,In_186,In_1356);
nand U1460 (N_1460,In_725,In_135);
or U1461 (N_1461,In_1895,In_591);
nor U1462 (N_1462,In_1605,In_963);
nor U1463 (N_1463,In_1869,In_1650);
or U1464 (N_1464,In_743,In_1789);
nand U1465 (N_1465,In_26,In_1900);
and U1466 (N_1466,In_892,In_303);
nor U1467 (N_1467,In_1340,In_1833);
or U1468 (N_1468,In_477,In_1537);
nand U1469 (N_1469,In_963,In_601);
nor U1470 (N_1470,In_432,In_577);
or U1471 (N_1471,In_1045,In_1556);
xnor U1472 (N_1472,In_224,In_1013);
and U1473 (N_1473,In_1073,In_732);
nor U1474 (N_1474,In_1431,In_212);
nor U1475 (N_1475,In_13,In_1926);
nand U1476 (N_1476,In_307,In_827);
or U1477 (N_1477,In_658,In_61);
nand U1478 (N_1478,In_1331,In_353);
nand U1479 (N_1479,In_1499,In_1188);
or U1480 (N_1480,In_14,In_543);
xor U1481 (N_1481,In_1620,In_1997);
and U1482 (N_1482,In_140,In_1411);
nor U1483 (N_1483,In_327,In_412);
xor U1484 (N_1484,In_364,In_1476);
or U1485 (N_1485,In_1311,In_1431);
and U1486 (N_1486,In_989,In_1383);
nor U1487 (N_1487,In_1699,In_219);
or U1488 (N_1488,In_1971,In_627);
nor U1489 (N_1489,In_179,In_9);
nor U1490 (N_1490,In_1434,In_58);
nand U1491 (N_1491,In_422,In_341);
or U1492 (N_1492,In_435,In_562);
or U1493 (N_1493,In_601,In_276);
and U1494 (N_1494,In_865,In_319);
or U1495 (N_1495,In_1704,In_1480);
xor U1496 (N_1496,In_1359,In_845);
xor U1497 (N_1497,In_48,In_478);
xnor U1498 (N_1498,In_1749,In_1435);
nor U1499 (N_1499,In_1055,In_1200);
nor U1500 (N_1500,In_44,In_1748);
nor U1501 (N_1501,In_616,In_685);
or U1502 (N_1502,In_68,In_1211);
nor U1503 (N_1503,In_1280,In_1218);
nand U1504 (N_1504,In_1126,In_1588);
or U1505 (N_1505,In_1833,In_1360);
xor U1506 (N_1506,In_1503,In_731);
nor U1507 (N_1507,In_1551,In_778);
nand U1508 (N_1508,In_524,In_1545);
nand U1509 (N_1509,In_1068,In_1705);
or U1510 (N_1510,In_1216,In_226);
and U1511 (N_1511,In_109,In_1479);
or U1512 (N_1512,In_1857,In_1126);
nor U1513 (N_1513,In_1471,In_1768);
and U1514 (N_1514,In_580,In_211);
and U1515 (N_1515,In_680,In_913);
or U1516 (N_1516,In_689,In_1640);
and U1517 (N_1517,In_412,In_179);
and U1518 (N_1518,In_1659,In_614);
nor U1519 (N_1519,In_74,In_1932);
or U1520 (N_1520,In_1039,In_1620);
or U1521 (N_1521,In_315,In_115);
nor U1522 (N_1522,In_1183,In_738);
nor U1523 (N_1523,In_1904,In_763);
and U1524 (N_1524,In_458,In_960);
nand U1525 (N_1525,In_922,In_604);
nor U1526 (N_1526,In_261,In_839);
or U1527 (N_1527,In_1391,In_1620);
nand U1528 (N_1528,In_124,In_1274);
nand U1529 (N_1529,In_963,In_847);
nor U1530 (N_1530,In_383,In_573);
nor U1531 (N_1531,In_480,In_395);
or U1532 (N_1532,In_1555,In_1481);
and U1533 (N_1533,In_693,In_310);
or U1534 (N_1534,In_279,In_1611);
or U1535 (N_1535,In_38,In_1153);
nand U1536 (N_1536,In_1986,In_211);
nor U1537 (N_1537,In_1546,In_1186);
nand U1538 (N_1538,In_1360,In_642);
and U1539 (N_1539,In_1882,In_1025);
nand U1540 (N_1540,In_468,In_1478);
nand U1541 (N_1541,In_1139,In_1801);
or U1542 (N_1542,In_851,In_1798);
xor U1543 (N_1543,In_1603,In_1333);
or U1544 (N_1544,In_1546,In_173);
and U1545 (N_1545,In_1936,In_436);
nor U1546 (N_1546,In_1200,In_356);
and U1547 (N_1547,In_477,In_837);
nand U1548 (N_1548,In_768,In_253);
nor U1549 (N_1549,In_493,In_196);
or U1550 (N_1550,In_1376,In_1681);
or U1551 (N_1551,In_932,In_270);
nand U1552 (N_1552,In_287,In_1915);
nand U1553 (N_1553,In_675,In_109);
nor U1554 (N_1554,In_616,In_150);
xnor U1555 (N_1555,In_777,In_1172);
nor U1556 (N_1556,In_22,In_913);
nand U1557 (N_1557,In_1822,In_1877);
nand U1558 (N_1558,In_462,In_407);
and U1559 (N_1559,In_62,In_1004);
nand U1560 (N_1560,In_1415,In_1649);
nor U1561 (N_1561,In_1529,In_1878);
and U1562 (N_1562,In_218,In_1096);
xnor U1563 (N_1563,In_228,In_1155);
or U1564 (N_1564,In_889,In_1142);
nand U1565 (N_1565,In_918,In_610);
nand U1566 (N_1566,In_996,In_1192);
and U1567 (N_1567,In_24,In_1076);
and U1568 (N_1568,In_230,In_1590);
and U1569 (N_1569,In_187,In_1676);
and U1570 (N_1570,In_1064,In_84);
nor U1571 (N_1571,In_1187,In_1918);
and U1572 (N_1572,In_467,In_1520);
nor U1573 (N_1573,In_802,In_253);
nand U1574 (N_1574,In_1652,In_1184);
nor U1575 (N_1575,In_1931,In_1925);
nor U1576 (N_1576,In_1197,In_1783);
nand U1577 (N_1577,In_1268,In_1563);
nand U1578 (N_1578,In_854,In_1503);
and U1579 (N_1579,In_1014,In_587);
or U1580 (N_1580,In_37,In_1567);
or U1581 (N_1581,In_1513,In_1398);
nor U1582 (N_1582,In_1207,In_722);
nand U1583 (N_1583,In_560,In_1442);
nor U1584 (N_1584,In_182,In_1016);
or U1585 (N_1585,In_1339,In_759);
nor U1586 (N_1586,In_1710,In_142);
xor U1587 (N_1587,In_1944,In_1868);
xnor U1588 (N_1588,In_49,In_68);
or U1589 (N_1589,In_340,In_1300);
nand U1590 (N_1590,In_1764,In_1397);
nand U1591 (N_1591,In_1043,In_507);
nand U1592 (N_1592,In_843,In_1785);
nor U1593 (N_1593,In_1967,In_904);
nand U1594 (N_1594,In_9,In_1595);
or U1595 (N_1595,In_593,In_303);
nand U1596 (N_1596,In_937,In_5);
nor U1597 (N_1597,In_317,In_615);
nand U1598 (N_1598,In_1214,In_635);
and U1599 (N_1599,In_964,In_1033);
xnor U1600 (N_1600,In_266,In_675);
or U1601 (N_1601,In_1589,In_435);
and U1602 (N_1602,In_945,In_826);
nand U1603 (N_1603,In_1922,In_698);
nor U1604 (N_1604,In_775,In_416);
nor U1605 (N_1605,In_349,In_9);
nor U1606 (N_1606,In_1169,In_783);
nand U1607 (N_1607,In_878,In_998);
or U1608 (N_1608,In_1383,In_712);
nand U1609 (N_1609,In_735,In_1077);
nand U1610 (N_1610,In_695,In_1979);
or U1611 (N_1611,In_1703,In_1454);
and U1612 (N_1612,In_590,In_1985);
nand U1613 (N_1613,In_1473,In_920);
nand U1614 (N_1614,In_192,In_1747);
xor U1615 (N_1615,In_108,In_1540);
nand U1616 (N_1616,In_1330,In_451);
or U1617 (N_1617,In_363,In_1239);
nand U1618 (N_1618,In_866,In_1971);
or U1619 (N_1619,In_1571,In_930);
or U1620 (N_1620,In_543,In_660);
nand U1621 (N_1621,In_199,In_1190);
and U1622 (N_1622,In_97,In_676);
nand U1623 (N_1623,In_516,In_870);
nand U1624 (N_1624,In_1470,In_279);
nand U1625 (N_1625,In_1682,In_851);
nor U1626 (N_1626,In_933,In_565);
and U1627 (N_1627,In_1147,In_1922);
xor U1628 (N_1628,In_255,In_706);
and U1629 (N_1629,In_1762,In_105);
nand U1630 (N_1630,In_12,In_912);
or U1631 (N_1631,In_1277,In_1590);
nand U1632 (N_1632,In_483,In_1442);
or U1633 (N_1633,In_1583,In_998);
nor U1634 (N_1634,In_986,In_819);
or U1635 (N_1635,In_1171,In_1529);
or U1636 (N_1636,In_187,In_246);
nand U1637 (N_1637,In_628,In_459);
nor U1638 (N_1638,In_372,In_1426);
nor U1639 (N_1639,In_1791,In_1905);
or U1640 (N_1640,In_1239,In_1870);
or U1641 (N_1641,In_685,In_443);
nand U1642 (N_1642,In_155,In_180);
xor U1643 (N_1643,In_841,In_1929);
nor U1644 (N_1644,In_404,In_73);
and U1645 (N_1645,In_1921,In_1897);
nor U1646 (N_1646,In_556,In_88);
nand U1647 (N_1647,In_1430,In_1497);
nand U1648 (N_1648,In_1033,In_217);
or U1649 (N_1649,In_1768,In_787);
nor U1650 (N_1650,In_1279,In_998);
or U1651 (N_1651,In_1362,In_621);
or U1652 (N_1652,In_1551,In_1378);
or U1653 (N_1653,In_1107,In_422);
and U1654 (N_1654,In_1222,In_413);
and U1655 (N_1655,In_1353,In_273);
and U1656 (N_1656,In_375,In_1157);
nor U1657 (N_1657,In_581,In_767);
nand U1658 (N_1658,In_1994,In_1775);
nand U1659 (N_1659,In_819,In_1573);
and U1660 (N_1660,In_1727,In_1185);
or U1661 (N_1661,In_1927,In_1877);
or U1662 (N_1662,In_1108,In_1387);
xor U1663 (N_1663,In_1010,In_327);
and U1664 (N_1664,In_389,In_503);
or U1665 (N_1665,In_1692,In_397);
or U1666 (N_1666,In_835,In_162);
nand U1667 (N_1667,In_1787,In_1007);
and U1668 (N_1668,In_1727,In_398);
nand U1669 (N_1669,In_1941,In_276);
and U1670 (N_1670,In_1458,In_495);
or U1671 (N_1671,In_1122,In_1145);
and U1672 (N_1672,In_1129,In_27);
or U1673 (N_1673,In_1609,In_1026);
and U1674 (N_1674,In_1094,In_1625);
nand U1675 (N_1675,In_68,In_1810);
xnor U1676 (N_1676,In_1170,In_1531);
or U1677 (N_1677,In_257,In_307);
nand U1678 (N_1678,In_1006,In_302);
and U1679 (N_1679,In_1818,In_1109);
nand U1680 (N_1680,In_769,In_445);
nor U1681 (N_1681,In_360,In_610);
and U1682 (N_1682,In_336,In_1390);
nand U1683 (N_1683,In_446,In_1018);
and U1684 (N_1684,In_1116,In_306);
and U1685 (N_1685,In_1327,In_1467);
and U1686 (N_1686,In_663,In_1390);
or U1687 (N_1687,In_992,In_870);
and U1688 (N_1688,In_232,In_1404);
nand U1689 (N_1689,In_1883,In_1724);
nor U1690 (N_1690,In_1916,In_1791);
xnor U1691 (N_1691,In_1662,In_1250);
and U1692 (N_1692,In_945,In_447);
nand U1693 (N_1693,In_511,In_891);
and U1694 (N_1694,In_1137,In_306);
nand U1695 (N_1695,In_1044,In_486);
or U1696 (N_1696,In_1330,In_1972);
or U1697 (N_1697,In_448,In_161);
nand U1698 (N_1698,In_1366,In_778);
and U1699 (N_1699,In_1351,In_51);
or U1700 (N_1700,In_1454,In_17);
and U1701 (N_1701,In_1586,In_1959);
nand U1702 (N_1702,In_1200,In_814);
nand U1703 (N_1703,In_1774,In_1408);
and U1704 (N_1704,In_775,In_415);
and U1705 (N_1705,In_447,In_810);
or U1706 (N_1706,In_26,In_1061);
nor U1707 (N_1707,In_1933,In_1887);
and U1708 (N_1708,In_1148,In_48);
and U1709 (N_1709,In_1600,In_1244);
or U1710 (N_1710,In_1477,In_64);
or U1711 (N_1711,In_1674,In_989);
nand U1712 (N_1712,In_126,In_1971);
xor U1713 (N_1713,In_351,In_1323);
and U1714 (N_1714,In_1765,In_65);
or U1715 (N_1715,In_1988,In_1927);
and U1716 (N_1716,In_1852,In_138);
or U1717 (N_1717,In_893,In_1368);
and U1718 (N_1718,In_1155,In_1181);
and U1719 (N_1719,In_112,In_1765);
nand U1720 (N_1720,In_1203,In_349);
or U1721 (N_1721,In_1378,In_1036);
nand U1722 (N_1722,In_1804,In_1359);
nand U1723 (N_1723,In_1809,In_1159);
nand U1724 (N_1724,In_217,In_577);
or U1725 (N_1725,In_1881,In_1291);
or U1726 (N_1726,In_1673,In_1740);
and U1727 (N_1727,In_222,In_1976);
nor U1728 (N_1728,In_1810,In_1031);
nand U1729 (N_1729,In_1387,In_1939);
or U1730 (N_1730,In_1410,In_1169);
and U1731 (N_1731,In_1458,In_1407);
nor U1732 (N_1732,In_1471,In_1117);
nand U1733 (N_1733,In_694,In_366);
or U1734 (N_1734,In_1745,In_622);
or U1735 (N_1735,In_1671,In_1906);
and U1736 (N_1736,In_258,In_845);
and U1737 (N_1737,In_1237,In_892);
nor U1738 (N_1738,In_1586,In_1625);
nand U1739 (N_1739,In_171,In_1552);
nor U1740 (N_1740,In_461,In_1687);
or U1741 (N_1741,In_987,In_222);
and U1742 (N_1742,In_785,In_905);
or U1743 (N_1743,In_768,In_475);
or U1744 (N_1744,In_1319,In_1962);
or U1745 (N_1745,In_1846,In_1895);
nand U1746 (N_1746,In_1334,In_38);
nand U1747 (N_1747,In_741,In_351);
and U1748 (N_1748,In_328,In_1406);
or U1749 (N_1749,In_574,In_297);
nor U1750 (N_1750,In_1044,In_1012);
nand U1751 (N_1751,In_1693,In_1689);
nor U1752 (N_1752,In_1169,In_718);
xnor U1753 (N_1753,In_1094,In_1112);
nand U1754 (N_1754,In_1161,In_1277);
or U1755 (N_1755,In_1445,In_1760);
and U1756 (N_1756,In_364,In_355);
nor U1757 (N_1757,In_1452,In_137);
nand U1758 (N_1758,In_298,In_1126);
nand U1759 (N_1759,In_1546,In_1911);
nor U1760 (N_1760,In_1371,In_416);
nand U1761 (N_1761,In_844,In_1113);
nand U1762 (N_1762,In_1245,In_321);
xnor U1763 (N_1763,In_1488,In_162);
or U1764 (N_1764,In_711,In_606);
or U1765 (N_1765,In_139,In_1975);
nor U1766 (N_1766,In_798,In_1164);
or U1767 (N_1767,In_1734,In_187);
or U1768 (N_1768,In_336,In_1514);
nand U1769 (N_1769,In_573,In_1281);
or U1770 (N_1770,In_1207,In_1350);
or U1771 (N_1771,In_2,In_1227);
or U1772 (N_1772,In_1360,In_1103);
or U1773 (N_1773,In_1129,In_1850);
or U1774 (N_1774,In_339,In_567);
nand U1775 (N_1775,In_30,In_522);
nand U1776 (N_1776,In_770,In_1944);
nand U1777 (N_1777,In_1677,In_142);
and U1778 (N_1778,In_1363,In_45);
and U1779 (N_1779,In_263,In_1270);
nor U1780 (N_1780,In_889,In_141);
or U1781 (N_1781,In_150,In_227);
nand U1782 (N_1782,In_706,In_1791);
xnor U1783 (N_1783,In_1075,In_661);
or U1784 (N_1784,In_1908,In_1982);
nand U1785 (N_1785,In_1053,In_334);
and U1786 (N_1786,In_619,In_347);
and U1787 (N_1787,In_1232,In_356);
nor U1788 (N_1788,In_1228,In_835);
and U1789 (N_1789,In_1220,In_328);
and U1790 (N_1790,In_1074,In_635);
xor U1791 (N_1791,In_1639,In_1897);
and U1792 (N_1792,In_290,In_236);
nor U1793 (N_1793,In_70,In_1674);
or U1794 (N_1794,In_938,In_1901);
nand U1795 (N_1795,In_1216,In_842);
or U1796 (N_1796,In_1658,In_614);
or U1797 (N_1797,In_866,In_1131);
nand U1798 (N_1798,In_1809,In_1324);
nand U1799 (N_1799,In_1296,In_1280);
nor U1800 (N_1800,In_1129,In_1872);
nor U1801 (N_1801,In_374,In_777);
and U1802 (N_1802,In_1864,In_148);
nand U1803 (N_1803,In_1451,In_538);
and U1804 (N_1804,In_1459,In_785);
or U1805 (N_1805,In_1977,In_104);
nor U1806 (N_1806,In_151,In_663);
nor U1807 (N_1807,In_1626,In_193);
or U1808 (N_1808,In_1695,In_1966);
nor U1809 (N_1809,In_1847,In_841);
and U1810 (N_1810,In_1194,In_827);
or U1811 (N_1811,In_1383,In_1428);
xor U1812 (N_1812,In_522,In_520);
or U1813 (N_1813,In_1566,In_426);
or U1814 (N_1814,In_1011,In_234);
nor U1815 (N_1815,In_894,In_395);
or U1816 (N_1816,In_1582,In_598);
or U1817 (N_1817,In_1918,In_1523);
or U1818 (N_1818,In_1824,In_1403);
nor U1819 (N_1819,In_1450,In_1027);
nor U1820 (N_1820,In_1578,In_1922);
nand U1821 (N_1821,In_803,In_882);
or U1822 (N_1822,In_1029,In_1429);
nor U1823 (N_1823,In_1435,In_1487);
or U1824 (N_1824,In_1338,In_600);
nor U1825 (N_1825,In_1123,In_1959);
nor U1826 (N_1826,In_720,In_1677);
or U1827 (N_1827,In_1989,In_765);
nor U1828 (N_1828,In_958,In_150);
or U1829 (N_1829,In_1643,In_122);
xor U1830 (N_1830,In_1434,In_1637);
or U1831 (N_1831,In_1962,In_752);
nand U1832 (N_1832,In_172,In_64);
or U1833 (N_1833,In_553,In_957);
nor U1834 (N_1834,In_380,In_203);
and U1835 (N_1835,In_508,In_399);
nand U1836 (N_1836,In_883,In_789);
nor U1837 (N_1837,In_1992,In_1339);
and U1838 (N_1838,In_76,In_550);
nor U1839 (N_1839,In_1843,In_1261);
or U1840 (N_1840,In_1466,In_824);
nand U1841 (N_1841,In_237,In_1521);
nor U1842 (N_1842,In_1890,In_682);
and U1843 (N_1843,In_520,In_494);
nand U1844 (N_1844,In_1338,In_1262);
nand U1845 (N_1845,In_1179,In_561);
xor U1846 (N_1846,In_1066,In_1931);
xor U1847 (N_1847,In_205,In_608);
and U1848 (N_1848,In_1855,In_254);
nand U1849 (N_1849,In_157,In_1626);
nor U1850 (N_1850,In_1139,In_38);
nand U1851 (N_1851,In_672,In_768);
or U1852 (N_1852,In_333,In_1378);
or U1853 (N_1853,In_1193,In_352);
nand U1854 (N_1854,In_1385,In_1011);
and U1855 (N_1855,In_1744,In_1776);
and U1856 (N_1856,In_1163,In_923);
and U1857 (N_1857,In_736,In_1029);
nand U1858 (N_1858,In_1042,In_1696);
nor U1859 (N_1859,In_1134,In_1250);
or U1860 (N_1860,In_1410,In_711);
nand U1861 (N_1861,In_1619,In_1068);
nor U1862 (N_1862,In_239,In_146);
and U1863 (N_1863,In_1141,In_1712);
nor U1864 (N_1864,In_198,In_1373);
nand U1865 (N_1865,In_1977,In_536);
and U1866 (N_1866,In_1460,In_1880);
nor U1867 (N_1867,In_1209,In_578);
nor U1868 (N_1868,In_236,In_1209);
nor U1869 (N_1869,In_1742,In_144);
nor U1870 (N_1870,In_1065,In_1295);
or U1871 (N_1871,In_943,In_1263);
and U1872 (N_1872,In_1027,In_1198);
nor U1873 (N_1873,In_1459,In_1406);
and U1874 (N_1874,In_1772,In_282);
or U1875 (N_1875,In_1176,In_943);
and U1876 (N_1876,In_1103,In_1532);
nand U1877 (N_1877,In_1493,In_794);
and U1878 (N_1878,In_1305,In_853);
or U1879 (N_1879,In_1678,In_1047);
xnor U1880 (N_1880,In_939,In_705);
nand U1881 (N_1881,In_197,In_1410);
and U1882 (N_1882,In_1410,In_462);
or U1883 (N_1883,In_1469,In_358);
nor U1884 (N_1884,In_89,In_656);
and U1885 (N_1885,In_190,In_1279);
or U1886 (N_1886,In_266,In_151);
or U1887 (N_1887,In_659,In_541);
nand U1888 (N_1888,In_869,In_652);
and U1889 (N_1889,In_1127,In_1440);
and U1890 (N_1890,In_1434,In_1980);
nor U1891 (N_1891,In_1153,In_172);
nand U1892 (N_1892,In_21,In_1059);
and U1893 (N_1893,In_1536,In_851);
nor U1894 (N_1894,In_1187,In_171);
nor U1895 (N_1895,In_1446,In_1801);
or U1896 (N_1896,In_29,In_773);
or U1897 (N_1897,In_1911,In_734);
and U1898 (N_1898,In_170,In_830);
nor U1899 (N_1899,In_1971,In_1248);
xor U1900 (N_1900,In_366,In_1369);
xor U1901 (N_1901,In_341,In_974);
or U1902 (N_1902,In_1133,In_451);
xor U1903 (N_1903,In_928,In_1839);
or U1904 (N_1904,In_1203,In_1811);
and U1905 (N_1905,In_1115,In_1043);
and U1906 (N_1906,In_1027,In_15);
nand U1907 (N_1907,In_1900,In_518);
or U1908 (N_1908,In_1184,In_462);
xnor U1909 (N_1909,In_803,In_1018);
or U1910 (N_1910,In_1058,In_664);
nand U1911 (N_1911,In_528,In_1340);
nor U1912 (N_1912,In_1146,In_1339);
and U1913 (N_1913,In_1683,In_1197);
or U1914 (N_1914,In_749,In_634);
nand U1915 (N_1915,In_136,In_355);
and U1916 (N_1916,In_776,In_895);
or U1917 (N_1917,In_1939,In_256);
xor U1918 (N_1918,In_1974,In_335);
nand U1919 (N_1919,In_353,In_1479);
nor U1920 (N_1920,In_674,In_218);
or U1921 (N_1921,In_1931,In_1892);
nor U1922 (N_1922,In_538,In_1514);
nand U1923 (N_1923,In_1798,In_1572);
or U1924 (N_1924,In_1225,In_610);
nor U1925 (N_1925,In_1487,In_690);
nor U1926 (N_1926,In_102,In_48);
and U1927 (N_1927,In_362,In_1456);
nand U1928 (N_1928,In_91,In_685);
and U1929 (N_1929,In_604,In_157);
nand U1930 (N_1930,In_655,In_1584);
or U1931 (N_1931,In_636,In_1183);
or U1932 (N_1932,In_165,In_119);
or U1933 (N_1933,In_356,In_1622);
and U1934 (N_1934,In_856,In_239);
nand U1935 (N_1935,In_1495,In_120);
nand U1936 (N_1936,In_1280,In_846);
and U1937 (N_1937,In_1613,In_1578);
or U1938 (N_1938,In_841,In_464);
and U1939 (N_1939,In_1333,In_724);
nor U1940 (N_1940,In_1731,In_310);
nand U1941 (N_1941,In_121,In_1199);
or U1942 (N_1942,In_1278,In_1740);
nand U1943 (N_1943,In_742,In_1191);
nor U1944 (N_1944,In_1615,In_14);
or U1945 (N_1945,In_1147,In_1921);
nand U1946 (N_1946,In_1884,In_750);
nor U1947 (N_1947,In_392,In_1269);
xor U1948 (N_1948,In_1467,In_1851);
nor U1949 (N_1949,In_134,In_668);
or U1950 (N_1950,In_471,In_1138);
nand U1951 (N_1951,In_902,In_421);
nand U1952 (N_1952,In_1980,In_1023);
and U1953 (N_1953,In_283,In_515);
nand U1954 (N_1954,In_1589,In_658);
nor U1955 (N_1955,In_1656,In_1076);
and U1956 (N_1956,In_1534,In_941);
nand U1957 (N_1957,In_602,In_441);
nor U1958 (N_1958,In_76,In_1259);
and U1959 (N_1959,In_1296,In_266);
and U1960 (N_1960,In_804,In_1011);
nor U1961 (N_1961,In_358,In_667);
and U1962 (N_1962,In_1093,In_1794);
or U1963 (N_1963,In_296,In_4);
or U1964 (N_1964,In_604,In_705);
or U1965 (N_1965,In_1099,In_1948);
or U1966 (N_1966,In_1153,In_1102);
or U1967 (N_1967,In_574,In_1541);
and U1968 (N_1968,In_1874,In_1899);
nor U1969 (N_1969,In_1830,In_753);
and U1970 (N_1970,In_1355,In_1299);
or U1971 (N_1971,In_1158,In_824);
and U1972 (N_1972,In_432,In_1017);
or U1973 (N_1973,In_104,In_555);
xor U1974 (N_1974,In_885,In_579);
nand U1975 (N_1975,In_1382,In_1339);
and U1976 (N_1976,In_741,In_924);
and U1977 (N_1977,In_238,In_1709);
nand U1978 (N_1978,In_1928,In_1620);
nor U1979 (N_1979,In_1776,In_986);
nor U1980 (N_1980,In_1748,In_634);
nand U1981 (N_1981,In_304,In_460);
or U1982 (N_1982,In_455,In_560);
nor U1983 (N_1983,In_170,In_1262);
xor U1984 (N_1984,In_1261,In_1615);
nor U1985 (N_1985,In_833,In_485);
or U1986 (N_1986,In_970,In_1769);
nand U1987 (N_1987,In_1037,In_358);
and U1988 (N_1988,In_781,In_737);
nand U1989 (N_1989,In_348,In_1928);
or U1990 (N_1990,In_85,In_1678);
nand U1991 (N_1991,In_50,In_371);
and U1992 (N_1992,In_1907,In_1759);
nand U1993 (N_1993,In_850,In_1880);
and U1994 (N_1994,In_334,In_1132);
nand U1995 (N_1995,In_1415,In_754);
nor U1996 (N_1996,In_1030,In_1141);
and U1997 (N_1997,In_588,In_419);
nor U1998 (N_1998,In_551,In_646);
or U1999 (N_1999,In_1440,In_1622);
nor U2000 (N_2000,In_1313,In_1033);
and U2001 (N_2001,In_215,In_122);
and U2002 (N_2002,In_201,In_1995);
or U2003 (N_2003,In_1304,In_1310);
nor U2004 (N_2004,In_1869,In_1376);
nand U2005 (N_2005,In_366,In_396);
xor U2006 (N_2006,In_974,In_1082);
and U2007 (N_2007,In_1525,In_905);
nand U2008 (N_2008,In_595,In_1675);
and U2009 (N_2009,In_1619,In_1925);
xnor U2010 (N_2010,In_1115,In_1289);
nand U2011 (N_2011,In_1397,In_1437);
nand U2012 (N_2012,In_1381,In_3);
or U2013 (N_2013,In_754,In_1558);
nor U2014 (N_2014,In_1129,In_376);
nand U2015 (N_2015,In_1216,In_259);
and U2016 (N_2016,In_1922,In_1593);
nor U2017 (N_2017,In_1893,In_978);
or U2018 (N_2018,In_1284,In_592);
nand U2019 (N_2019,In_1273,In_237);
nand U2020 (N_2020,In_462,In_1337);
nor U2021 (N_2021,In_621,In_1605);
nand U2022 (N_2022,In_1618,In_1344);
nand U2023 (N_2023,In_853,In_837);
nand U2024 (N_2024,In_1502,In_356);
nand U2025 (N_2025,In_1001,In_1954);
and U2026 (N_2026,In_184,In_1717);
or U2027 (N_2027,In_1968,In_1926);
xor U2028 (N_2028,In_721,In_84);
and U2029 (N_2029,In_964,In_1357);
nor U2030 (N_2030,In_50,In_1123);
xnor U2031 (N_2031,In_1631,In_792);
and U2032 (N_2032,In_455,In_736);
xor U2033 (N_2033,In_596,In_4);
or U2034 (N_2034,In_342,In_1656);
nor U2035 (N_2035,In_1447,In_896);
and U2036 (N_2036,In_180,In_442);
nor U2037 (N_2037,In_267,In_1074);
nand U2038 (N_2038,In_227,In_443);
or U2039 (N_2039,In_37,In_644);
nor U2040 (N_2040,In_1821,In_1867);
nor U2041 (N_2041,In_67,In_119);
nor U2042 (N_2042,In_592,In_807);
nand U2043 (N_2043,In_1915,In_1875);
nand U2044 (N_2044,In_1813,In_3);
nand U2045 (N_2045,In_333,In_1207);
nand U2046 (N_2046,In_1937,In_280);
or U2047 (N_2047,In_847,In_109);
or U2048 (N_2048,In_163,In_1078);
and U2049 (N_2049,In_1897,In_1359);
nand U2050 (N_2050,In_1464,In_271);
xnor U2051 (N_2051,In_50,In_1964);
nand U2052 (N_2052,In_185,In_1527);
xor U2053 (N_2053,In_1634,In_1);
nand U2054 (N_2054,In_292,In_1418);
nor U2055 (N_2055,In_151,In_95);
nand U2056 (N_2056,In_724,In_192);
and U2057 (N_2057,In_175,In_1375);
nand U2058 (N_2058,In_177,In_336);
and U2059 (N_2059,In_267,In_969);
and U2060 (N_2060,In_1040,In_345);
and U2061 (N_2061,In_12,In_762);
xnor U2062 (N_2062,In_826,In_1172);
nor U2063 (N_2063,In_1008,In_975);
or U2064 (N_2064,In_1982,In_1254);
or U2065 (N_2065,In_948,In_942);
or U2066 (N_2066,In_796,In_1336);
xor U2067 (N_2067,In_719,In_1043);
or U2068 (N_2068,In_1538,In_131);
xnor U2069 (N_2069,In_1138,In_711);
nor U2070 (N_2070,In_1296,In_1903);
nor U2071 (N_2071,In_1442,In_422);
and U2072 (N_2072,In_362,In_1252);
xor U2073 (N_2073,In_1118,In_1619);
nand U2074 (N_2074,In_1022,In_1537);
or U2075 (N_2075,In_656,In_337);
nor U2076 (N_2076,In_1309,In_91);
and U2077 (N_2077,In_1825,In_1091);
or U2078 (N_2078,In_140,In_1758);
or U2079 (N_2079,In_1154,In_1905);
or U2080 (N_2080,In_1091,In_309);
and U2081 (N_2081,In_1423,In_90);
nor U2082 (N_2082,In_1652,In_760);
nand U2083 (N_2083,In_47,In_1443);
nand U2084 (N_2084,In_331,In_607);
nor U2085 (N_2085,In_1110,In_1367);
and U2086 (N_2086,In_1906,In_1405);
or U2087 (N_2087,In_1380,In_173);
nor U2088 (N_2088,In_1199,In_945);
xnor U2089 (N_2089,In_1161,In_1188);
nor U2090 (N_2090,In_1940,In_1372);
nand U2091 (N_2091,In_1113,In_64);
nand U2092 (N_2092,In_1291,In_1675);
and U2093 (N_2093,In_74,In_1058);
nand U2094 (N_2094,In_383,In_1989);
and U2095 (N_2095,In_736,In_851);
or U2096 (N_2096,In_348,In_575);
nor U2097 (N_2097,In_1151,In_1054);
and U2098 (N_2098,In_1061,In_1420);
or U2099 (N_2099,In_220,In_1186);
nor U2100 (N_2100,In_301,In_452);
nor U2101 (N_2101,In_1892,In_1997);
or U2102 (N_2102,In_1981,In_1566);
and U2103 (N_2103,In_1992,In_1850);
nand U2104 (N_2104,In_119,In_74);
nor U2105 (N_2105,In_303,In_271);
or U2106 (N_2106,In_605,In_1131);
and U2107 (N_2107,In_1779,In_42);
nor U2108 (N_2108,In_388,In_1076);
or U2109 (N_2109,In_832,In_464);
xnor U2110 (N_2110,In_1903,In_76);
or U2111 (N_2111,In_950,In_719);
and U2112 (N_2112,In_664,In_1122);
nand U2113 (N_2113,In_404,In_256);
nor U2114 (N_2114,In_1839,In_183);
xnor U2115 (N_2115,In_362,In_427);
or U2116 (N_2116,In_916,In_871);
nor U2117 (N_2117,In_1356,In_1857);
nand U2118 (N_2118,In_250,In_1156);
nand U2119 (N_2119,In_237,In_1095);
nor U2120 (N_2120,In_1358,In_1294);
nor U2121 (N_2121,In_166,In_867);
nor U2122 (N_2122,In_1594,In_641);
and U2123 (N_2123,In_949,In_114);
nand U2124 (N_2124,In_1894,In_540);
and U2125 (N_2125,In_1161,In_367);
or U2126 (N_2126,In_677,In_995);
nand U2127 (N_2127,In_1347,In_1717);
nor U2128 (N_2128,In_1319,In_309);
or U2129 (N_2129,In_1743,In_289);
nor U2130 (N_2130,In_140,In_725);
nand U2131 (N_2131,In_922,In_1669);
or U2132 (N_2132,In_872,In_180);
or U2133 (N_2133,In_1984,In_1221);
nor U2134 (N_2134,In_1844,In_1957);
or U2135 (N_2135,In_1886,In_86);
or U2136 (N_2136,In_380,In_1349);
xnor U2137 (N_2137,In_1140,In_744);
or U2138 (N_2138,In_539,In_1953);
or U2139 (N_2139,In_1375,In_1921);
nor U2140 (N_2140,In_52,In_149);
nor U2141 (N_2141,In_1227,In_323);
nand U2142 (N_2142,In_127,In_766);
or U2143 (N_2143,In_1747,In_1850);
nand U2144 (N_2144,In_1901,In_274);
or U2145 (N_2145,In_1287,In_786);
nand U2146 (N_2146,In_635,In_946);
nor U2147 (N_2147,In_1368,In_1676);
nor U2148 (N_2148,In_592,In_1179);
nor U2149 (N_2149,In_1120,In_1971);
or U2150 (N_2150,In_950,In_412);
xor U2151 (N_2151,In_1293,In_19);
or U2152 (N_2152,In_1305,In_1765);
and U2153 (N_2153,In_1584,In_903);
nor U2154 (N_2154,In_529,In_118);
nor U2155 (N_2155,In_1896,In_1716);
or U2156 (N_2156,In_401,In_1044);
nor U2157 (N_2157,In_93,In_675);
nor U2158 (N_2158,In_866,In_148);
nor U2159 (N_2159,In_686,In_547);
and U2160 (N_2160,In_630,In_488);
nor U2161 (N_2161,In_1406,In_251);
or U2162 (N_2162,In_125,In_1892);
nand U2163 (N_2163,In_1938,In_663);
or U2164 (N_2164,In_608,In_108);
and U2165 (N_2165,In_5,In_1127);
nand U2166 (N_2166,In_364,In_600);
xnor U2167 (N_2167,In_396,In_1930);
and U2168 (N_2168,In_318,In_962);
or U2169 (N_2169,In_225,In_1663);
nor U2170 (N_2170,In_1612,In_1903);
or U2171 (N_2171,In_263,In_1183);
nor U2172 (N_2172,In_385,In_355);
nor U2173 (N_2173,In_1612,In_1166);
nor U2174 (N_2174,In_662,In_622);
or U2175 (N_2175,In_1962,In_371);
or U2176 (N_2176,In_428,In_1439);
nor U2177 (N_2177,In_31,In_326);
and U2178 (N_2178,In_1866,In_1080);
or U2179 (N_2179,In_560,In_1198);
nor U2180 (N_2180,In_1360,In_932);
nand U2181 (N_2181,In_1105,In_855);
nor U2182 (N_2182,In_926,In_1503);
xor U2183 (N_2183,In_870,In_1657);
or U2184 (N_2184,In_866,In_614);
or U2185 (N_2185,In_1658,In_168);
and U2186 (N_2186,In_1008,In_1382);
nor U2187 (N_2187,In_393,In_315);
nand U2188 (N_2188,In_943,In_405);
and U2189 (N_2189,In_159,In_1013);
nor U2190 (N_2190,In_1888,In_743);
nor U2191 (N_2191,In_608,In_1090);
xor U2192 (N_2192,In_1402,In_1750);
and U2193 (N_2193,In_932,In_1215);
or U2194 (N_2194,In_1599,In_444);
nand U2195 (N_2195,In_972,In_587);
or U2196 (N_2196,In_1443,In_611);
nand U2197 (N_2197,In_773,In_876);
and U2198 (N_2198,In_1266,In_439);
nor U2199 (N_2199,In_1998,In_1823);
and U2200 (N_2200,In_304,In_86);
and U2201 (N_2201,In_1742,In_877);
and U2202 (N_2202,In_21,In_660);
and U2203 (N_2203,In_1518,In_1893);
or U2204 (N_2204,In_374,In_799);
nor U2205 (N_2205,In_1103,In_1818);
and U2206 (N_2206,In_704,In_597);
nand U2207 (N_2207,In_1750,In_461);
nor U2208 (N_2208,In_985,In_431);
nor U2209 (N_2209,In_1959,In_744);
nand U2210 (N_2210,In_276,In_1303);
and U2211 (N_2211,In_1698,In_509);
or U2212 (N_2212,In_1930,In_1989);
and U2213 (N_2213,In_1008,In_659);
nand U2214 (N_2214,In_1078,In_1425);
nor U2215 (N_2215,In_24,In_1520);
and U2216 (N_2216,In_1642,In_1834);
xnor U2217 (N_2217,In_1060,In_320);
nand U2218 (N_2218,In_1553,In_1193);
nand U2219 (N_2219,In_1026,In_783);
and U2220 (N_2220,In_614,In_1354);
nor U2221 (N_2221,In_1207,In_329);
nor U2222 (N_2222,In_1017,In_926);
nor U2223 (N_2223,In_1599,In_1476);
nor U2224 (N_2224,In_1135,In_1851);
and U2225 (N_2225,In_1578,In_405);
or U2226 (N_2226,In_1105,In_595);
nand U2227 (N_2227,In_1436,In_1941);
and U2228 (N_2228,In_1775,In_862);
or U2229 (N_2229,In_1597,In_734);
or U2230 (N_2230,In_716,In_675);
or U2231 (N_2231,In_822,In_309);
nor U2232 (N_2232,In_1473,In_1413);
nand U2233 (N_2233,In_940,In_44);
and U2234 (N_2234,In_104,In_1006);
nor U2235 (N_2235,In_1129,In_944);
and U2236 (N_2236,In_985,In_1515);
nor U2237 (N_2237,In_1847,In_1095);
nand U2238 (N_2238,In_1805,In_1972);
nor U2239 (N_2239,In_206,In_752);
nor U2240 (N_2240,In_1042,In_257);
xnor U2241 (N_2241,In_1227,In_1534);
nor U2242 (N_2242,In_1377,In_800);
or U2243 (N_2243,In_1740,In_397);
and U2244 (N_2244,In_930,In_190);
and U2245 (N_2245,In_39,In_64);
or U2246 (N_2246,In_1011,In_470);
nand U2247 (N_2247,In_850,In_32);
nand U2248 (N_2248,In_1801,In_899);
nand U2249 (N_2249,In_157,In_1304);
and U2250 (N_2250,In_1231,In_849);
nor U2251 (N_2251,In_1696,In_13);
nor U2252 (N_2252,In_458,In_1130);
or U2253 (N_2253,In_1093,In_525);
nor U2254 (N_2254,In_1356,In_1940);
or U2255 (N_2255,In_702,In_330);
and U2256 (N_2256,In_627,In_1271);
or U2257 (N_2257,In_1299,In_1788);
and U2258 (N_2258,In_590,In_634);
and U2259 (N_2259,In_695,In_901);
nand U2260 (N_2260,In_1015,In_749);
nor U2261 (N_2261,In_1439,In_1376);
nand U2262 (N_2262,In_85,In_361);
nor U2263 (N_2263,In_1811,In_1167);
nor U2264 (N_2264,In_929,In_1683);
or U2265 (N_2265,In_1621,In_423);
nor U2266 (N_2266,In_911,In_1174);
and U2267 (N_2267,In_1228,In_534);
or U2268 (N_2268,In_1574,In_796);
xor U2269 (N_2269,In_1645,In_626);
nand U2270 (N_2270,In_98,In_1896);
nor U2271 (N_2271,In_1836,In_731);
and U2272 (N_2272,In_819,In_1789);
xor U2273 (N_2273,In_790,In_1823);
or U2274 (N_2274,In_738,In_1886);
nor U2275 (N_2275,In_277,In_325);
nor U2276 (N_2276,In_503,In_549);
nor U2277 (N_2277,In_27,In_900);
or U2278 (N_2278,In_1391,In_1894);
nand U2279 (N_2279,In_572,In_128);
nor U2280 (N_2280,In_1532,In_488);
nand U2281 (N_2281,In_241,In_1431);
or U2282 (N_2282,In_1014,In_1929);
and U2283 (N_2283,In_1713,In_594);
nor U2284 (N_2284,In_1415,In_608);
or U2285 (N_2285,In_708,In_1661);
and U2286 (N_2286,In_75,In_177);
nor U2287 (N_2287,In_618,In_250);
and U2288 (N_2288,In_1680,In_1453);
nand U2289 (N_2289,In_1171,In_1925);
nand U2290 (N_2290,In_1063,In_1461);
nor U2291 (N_2291,In_1203,In_792);
and U2292 (N_2292,In_311,In_1218);
nand U2293 (N_2293,In_254,In_134);
or U2294 (N_2294,In_1734,In_1521);
and U2295 (N_2295,In_1374,In_1714);
or U2296 (N_2296,In_1620,In_660);
nand U2297 (N_2297,In_1928,In_1419);
xor U2298 (N_2298,In_50,In_903);
and U2299 (N_2299,In_1087,In_1717);
or U2300 (N_2300,In_880,In_1472);
and U2301 (N_2301,In_1521,In_959);
nand U2302 (N_2302,In_242,In_1531);
nor U2303 (N_2303,In_1902,In_248);
nand U2304 (N_2304,In_1012,In_1840);
nand U2305 (N_2305,In_1156,In_966);
xnor U2306 (N_2306,In_495,In_478);
xnor U2307 (N_2307,In_1236,In_964);
nand U2308 (N_2308,In_554,In_1739);
nor U2309 (N_2309,In_1174,In_1555);
xnor U2310 (N_2310,In_1675,In_1142);
xnor U2311 (N_2311,In_652,In_1536);
or U2312 (N_2312,In_1826,In_903);
nand U2313 (N_2313,In_812,In_208);
and U2314 (N_2314,In_653,In_343);
nor U2315 (N_2315,In_1270,In_1972);
nor U2316 (N_2316,In_1239,In_1439);
nor U2317 (N_2317,In_604,In_238);
or U2318 (N_2318,In_1912,In_1527);
nor U2319 (N_2319,In_1611,In_746);
or U2320 (N_2320,In_1875,In_884);
and U2321 (N_2321,In_621,In_740);
or U2322 (N_2322,In_913,In_1882);
nand U2323 (N_2323,In_756,In_671);
nand U2324 (N_2324,In_1740,In_871);
nor U2325 (N_2325,In_178,In_1136);
or U2326 (N_2326,In_900,In_1467);
nand U2327 (N_2327,In_1883,In_1583);
or U2328 (N_2328,In_248,In_44);
nor U2329 (N_2329,In_546,In_679);
and U2330 (N_2330,In_1610,In_120);
and U2331 (N_2331,In_1643,In_709);
xor U2332 (N_2332,In_1592,In_400);
xnor U2333 (N_2333,In_910,In_1189);
nand U2334 (N_2334,In_1016,In_1744);
nand U2335 (N_2335,In_805,In_935);
nand U2336 (N_2336,In_76,In_1210);
nand U2337 (N_2337,In_1305,In_1984);
nand U2338 (N_2338,In_478,In_1694);
nand U2339 (N_2339,In_952,In_461);
and U2340 (N_2340,In_840,In_1916);
and U2341 (N_2341,In_1558,In_616);
nand U2342 (N_2342,In_114,In_1589);
nand U2343 (N_2343,In_1086,In_927);
xor U2344 (N_2344,In_1436,In_1619);
and U2345 (N_2345,In_591,In_848);
nor U2346 (N_2346,In_1826,In_1245);
nor U2347 (N_2347,In_1001,In_1814);
nand U2348 (N_2348,In_793,In_12);
and U2349 (N_2349,In_1566,In_536);
or U2350 (N_2350,In_1834,In_742);
nor U2351 (N_2351,In_1589,In_1416);
nor U2352 (N_2352,In_86,In_1493);
or U2353 (N_2353,In_212,In_654);
or U2354 (N_2354,In_1766,In_561);
nor U2355 (N_2355,In_265,In_717);
or U2356 (N_2356,In_1578,In_1809);
nand U2357 (N_2357,In_1354,In_162);
or U2358 (N_2358,In_204,In_1426);
and U2359 (N_2359,In_860,In_922);
nor U2360 (N_2360,In_1650,In_847);
and U2361 (N_2361,In_1474,In_1816);
nor U2362 (N_2362,In_1757,In_1546);
and U2363 (N_2363,In_1142,In_295);
or U2364 (N_2364,In_1537,In_1718);
nor U2365 (N_2365,In_1741,In_367);
nand U2366 (N_2366,In_254,In_302);
or U2367 (N_2367,In_355,In_916);
or U2368 (N_2368,In_1710,In_1590);
nand U2369 (N_2369,In_682,In_1387);
or U2370 (N_2370,In_1062,In_1601);
nand U2371 (N_2371,In_1214,In_74);
and U2372 (N_2372,In_1904,In_785);
nor U2373 (N_2373,In_1619,In_548);
nor U2374 (N_2374,In_1646,In_600);
nand U2375 (N_2375,In_996,In_1299);
xnor U2376 (N_2376,In_177,In_293);
nor U2377 (N_2377,In_1270,In_943);
or U2378 (N_2378,In_1090,In_1596);
nor U2379 (N_2379,In_1454,In_762);
nand U2380 (N_2380,In_1191,In_299);
or U2381 (N_2381,In_1286,In_332);
or U2382 (N_2382,In_1763,In_633);
nor U2383 (N_2383,In_652,In_153);
and U2384 (N_2384,In_1908,In_1291);
nor U2385 (N_2385,In_1973,In_1334);
and U2386 (N_2386,In_437,In_265);
or U2387 (N_2387,In_1712,In_1184);
or U2388 (N_2388,In_761,In_1539);
nand U2389 (N_2389,In_572,In_1050);
or U2390 (N_2390,In_1398,In_665);
and U2391 (N_2391,In_1462,In_29);
nand U2392 (N_2392,In_379,In_883);
nand U2393 (N_2393,In_842,In_1498);
and U2394 (N_2394,In_1678,In_306);
and U2395 (N_2395,In_241,In_1738);
or U2396 (N_2396,In_502,In_1963);
nand U2397 (N_2397,In_1943,In_515);
nor U2398 (N_2398,In_1246,In_1958);
nand U2399 (N_2399,In_1340,In_226);
nor U2400 (N_2400,In_1684,In_833);
and U2401 (N_2401,In_420,In_1595);
nand U2402 (N_2402,In_1481,In_1780);
or U2403 (N_2403,In_393,In_19);
and U2404 (N_2404,In_776,In_773);
and U2405 (N_2405,In_1425,In_1119);
and U2406 (N_2406,In_18,In_1058);
and U2407 (N_2407,In_1422,In_465);
or U2408 (N_2408,In_1997,In_292);
or U2409 (N_2409,In_787,In_1415);
nand U2410 (N_2410,In_1399,In_1712);
or U2411 (N_2411,In_93,In_884);
nand U2412 (N_2412,In_460,In_761);
nor U2413 (N_2413,In_664,In_575);
or U2414 (N_2414,In_922,In_874);
nor U2415 (N_2415,In_734,In_1341);
nand U2416 (N_2416,In_1023,In_1620);
and U2417 (N_2417,In_770,In_592);
nor U2418 (N_2418,In_1434,In_78);
nand U2419 (N_2419,In_1577,In_995);
nor U2420 (N_2420,In_1476,In_1889);
nor U2421 (N_2421,In_1902,In_1776);
nand U2422 (N_2422,In_32,In_704);
nor U2423 (N_2423,In_1260,In_1097);
nor U2424 (N_2424,In_1546,In_704);
and U2425 (N_2425,In_1973,In_1375);
nor U2426 (N_2426,In_1418,In_364);
or U2427 (N_2427,In_197,In_469);
nand U2428 (N_2428,In_1246,In_1569);
nand U2429 (N_2429,In_32,In_506);
or U2430 (N_2430,In_1363,In_1211);
or U2431 (N_2431,In_1644,In_1307);
and U2432 (N_2432,In_1590,In_477);
or U2433 (N_2433,In_1396,In_747);
nand U2434 (N_2434,In_459,In_789);
and U2435 (N_2435,In_1113,In_201);
nand U2436 (N_2436,In_939,In_1347);
nand U2437 (N_2437,In_1004,In_1795);
or U2438 (N_2438,In_918,In_1996);
or U2439 (N_2439,In_1820,In_1507);
and U2440 (N_2440,In_386,In_773);
or U2441 (N_2441,In_1819,In_154);
nor U2442 (N_2442,In_422,In_882);
xor U2443 (N_2443,In_73,In_626);
nor U2444 (N_2444,In_1124,In_1655);
and U2445 (N_2445,In_1253,In_134);
xor U2446 (N_2446,In_1661,In_465);
nor U2447 (N_2447,In_1456,In_1864);
and U2448 (N_2448,In_1792,In_688);
or U2449 (N_2449,In_894,In_1581);
nand U2450 (N_2450,In_641,In_334);
or U2451 (N_2451,In_829,In_329);
xnor U2452 (N_2452,In_1443,In_216);
nor U2453 (N_2453,In_1697,In_1863);
and U2454 (N_2454,In_641,In_11);
and U2455 (N_2455,In_984,In_460);
nand U2456 (N_2456,In_1979,In_1873);
nand U2457 (N_2457,In_1107,In_799);
or U2458 (N_2458,In_793,In_271);
and U2459 (N_2459,In_1904,In_943);
xnor U2460 (N_2460,In_663,In_302);
nor U2461 (N_2461,In_72,In_1078);
nand U2462 (N_2462,In_1168,In_1884);
and U2463 (N_2463,In_1319,In_729);
and U2464 (N_2464,In_604,In_1612);
and U2465 (N_2465,In_0,In_201);
or U2466 (N_2466,In_508,In_1856);
and U2467 (N_2467,In_300,In_807);
nand U2468 (N_2468,In_85,In_456);
nor U2469 (N_2469,In_663,In_72);
xor U2470 (N_2470,In_647,In_557);
and U2471 (N_2471,In_1904,In_1408);
or U2472 (N_2472,In_644,In_588);
or U2473 (N_2473,In_145,In_130);
nor U2474 (N_2474,In_1627,In_1934);
and U2475 (N_2475,In_1439,In_1002);
and U2476 (N_2476,In_473,In_1421);
nand U2477 (N_2477,In_116,In_862);
and U2478 (N_2478,In_96,In_934);
or U2479 (N_2479,In_893,In_1914);
or U2480 (N_2480,In_1044,In_43);
or U2481 (N_2481,In_1884,In_1361);
nor U2482 (N_2482,In_579,In_578);
nor U2483 (N_2483,In_1344,In_214);
xnor U2484 (N_2484,In_78,In_277);
and U2485 (N_2485,In_1919,In_564);
and U2486 (N_2486,In_1,In_1050);
nand U2487 (N_2487,In_1346,In_1231);
nor U2488 (N_2488,In_1056,In_1596);
and U2489 (N_2489,In_1522,In_1434);
and U2490 (N_2490,In_769,In_1425);
and U2491 (N_2491,In_3,In_161);
nand U2492 (N_2492,In_1740,In_1918);
nand U2493 (N_2493,In_857,In_492);
or U2494 (N_2494,In_294,In_638);
nor U2495 (N_2495,In_1468,In_605);
and U2496 (N_2496,In_1923,In_123);
nand U2497 (N_2497,In_1275,In_1629);
nor U2498 (N_2498,In_215,In_955);
or U2499 (N_2499,In_1732,In_1326);
nand U2500 (N_2500,In_1395,In_1943);
nand U2501 (N_2501,In_852,In_1597);
or U2502 (N_2502,In_1185,In_1407);
nand U2503 (N_2503,In_1190,In_782);
nand U2504 (N_2504,In_1192,In_928);
nor U2505 (N_2505,In_1118,In_654);
xor U2506 (N_2506,In_6,In_104);
nor U2507 (N_2507,In_155,In_1125);
nand U2508 (N_2508,In_395,In_1322);
and U2509 (N_2509,In_1287,In_1252);
nor U2510 (N_2510,In_1889,In_1606);
xor U2511 (N_2511,In_224,In_1682);
nand U2512 (N_2512,In_550,In_1266);
nor U2513 (N_2513,In_44,In_711);
or U2514 (N_2514,In_602,In_1275);
or U2515 (N_2515,In_1414,In_1705);
and U2516 (N_2516,In_429,In_208);
xor U2517 (N_2517,In_922,In_1960);
or U2518 (N_2518,In_314,In_782);
nor U2519 (N_2519,In_1081,In_1520);
nor U2520 (N_2520,In_1420,In_1092);
nor U2521 (N_2521,In_1369,In_622);
nor U2522 (N_2522,In_1709,In_574);
xor U2523 (N_2523,In_1467,In_459);
and U2524 (N_2524,In_1273,In_1167);
nand U2525 (N_2525,In_1391,In_1743);
nand U2526 (N_2526,In_719,In_709);
or U2527 (N_2527,In_531,In_1077);
and U2528 (N_2528,In_531,In_739);
and U2529 (N_2529,In_1168,In_712);
nand U2530 (N_2530,In_409,In_670);
nor U2531 (N_2531,In_402,In_1027);
nand U2532 (N_2532,In_870,In_295);
or U2533 (N_2533,In_565,In_99);
or U2534 (N_2534,In_1390,In_222);
and U2535 (N_2535,In_1418,In_401);
or U2536 (N_2536,In_1516,In_1087);
and U2537 (N_2537,In_112,In_1914);
nand U2538 (N_2538,In_1641,In_1123);
and U2539 (N_2539,In_781,In_991);
nor U2540 (N_2540,In_1693,In_1891);
nor U2541 (N_2541,In_177,In_1692);
and U2542 (N_2542,In_798,In_1358);
or U2543 (N_2543,In_50,In_1546);
nor U2544 (N_2544,In_875,In_1525);
nand U2545 (N_2545,In_749,In_1800);
nand U2546 (N_2546,In_692,In_384);
nor U2547 (N_2547,In_1481,In_1700);
and U2548 (N_2548,In_29,In_1275);
and U2549 (N_2549,In_569,In_1149);
or U2550 (N_2550,In_149,In_1310);
and U2551 (N_2551,In_1896,In_911);
nand U2552 (N_2552,In_1217,In_1660);
nand U2553 (N_2553,In_1790,In_1784);
and U2554 (N_2554,In_1981,In_211);
or U2555 (N_2555,In_1657,In_1010);
and U2556 (N_2556,In_97,In_1077);
and U2557 (N_2557,In_430,In_1795);
nor U2558 (N_2558,In_711,In_1553);
and U2559 (N_2559,In_773,In_1448);
nand U2560 (N_2560,In_337,In_1963);
nand U2561 (N_2561,In_1770,In_1071);
nor U2562 (N_2562,In_1093,In_1206);
xnor U2563 (N_2563,In_53,In_822);
nor U2564 (N_2564,In_733,In_291);
or U2565 (N_2565,In_1946,In_1702);
nor U2566 (N_2566,In_709,In_1425);
and U2567 (N_2567,In_431,In_119);
nand U2568 (N_2568,In_115,In_877);
xnor U2569 (N_2569,In_1216,In_1546);
nand U2570 (N_2570,In_878,In_1130);
or U2571 (N_2571,In_429,In_179);
nor U2572 (N_2572,In_60,In_1757);
nand U2573 (N_2573,In_44,In_1318);
nand U2574 (N_2574,In_1637,In_11);
or U2575 (N_2575,In_73,In_1033);
nor U2576 (N_2576,In_1384,In_1140);
nor U2577 (N_2577,In_396,In_506);
and U2578 (N_2578,In_505,In_1671);
nor U2579 (N_2579,In_1993,In_1472);
nand U2580 (N_2580,In_1963,In_1177);
nor U2581 (N_2581,In_784,In_621);
or U2582 (N_2582,In_401,In_257);
nor U2583 (N_2583,In_820,In_516);
xor U2584 (N_2584,In_531,In_584);
nand U2585 (N_2585,In_1297,In_1312);
and U2586 (N_2586,In_449,In_628);
nand U2587 (N_2587,In_286,In_191);
or U2588 (N_2588,In_1353,In_732);
nand U2589 (N_2589,In_557,In_68);
and U2590 (N_2590,In_1604,In_1916);
or U2591 (N_2591,In_32,In_886);
or U2592 (N_2592,In_295,In_1775);
and U2593 (N_2593,In_1683,In_1152);
and U2594 (N_2594,In_819,In_1521);
nand U2595 (N_2595,In_529,In_278);
nor U2596 (N_2596,In_425,In_646);
or U2597 (N_2597,In_117,In_797);
nand U2598 (N_2598,In_972,In_930);
or U2599 (N_2599,In_579,In_1686);
nand U2600 (N_2600,In_153,In_1592);
xor U2601 (N_2601,In_1583,In_229);
nor U2602 (N_2602,In_1782,In_325);
xnor U2603 (N_2603,In_64,In_1863);
nor U2604 (N_2604,In_1783,In_36);
and U2605 (N_2605,In_1707,In_1907);
or U2606 (N_2606,In_1116,In_681);
nor U2607 (N_2607,In_1082,In_547);
or U2608 (N_2608,In_87,In_1582);
and U2609 (N_2609,In_322,In_1747);
nand U2610 (N_2610,In_1043,In_773);
and U2611 (N_2611,In_20,In_1392);
and U2612 (N_2612,In_244,In_326);
or U2613 (N_2613,In_920,In_1923);
or U2614 (N_2614,In_1092,In_752);
and U2615 (N_2615,In_345,In_750);
nand U2616 (N_2616,In_827,In_1895);
nor U2617 (N_2617,In_1303,In_1227);
nor U2618 (N_2618,In_547,In_1551);
or U2619 (N_2619,In_1196,In_227);
nor U2620 (N_2620,In_1773,In_272);
and U2621 (N_2621,In_311,In_194);
nor U2622 (N_2622,In_1956,In_1225);
and U2623 (N_2623,In_1702,In_1743);
xor U2624 (N_2624,In_1289,In_1851);
and U2625 (N_2625,In_459,In_126);
nor U2626 (N_2626,In_598,In_1175);
and U2627 (N_2627,In_34,In_286);
or U2628 (N_2628,In_288,In_508);
nand U2629 (N_2629,In_207,In_1076);
and U2630 (N_2630,In_385,In_725);
nor U2631 (N_2631,In_1026,In_1663);
nand U2632 (N_2632,In_20,In_740);
nand U2633 (N_2633,In_49,In_486);
or U2634 (N_2634,In_752,In_628);
and U2635 (N_2635,In_1669,In_1200);
nor U2636 (N_2636,In_332,In_894);
and U2637 (N_2637,In_993,In_1644);
or U2638 (N_2638,In_1299,In_373);
and U2639 (N_2639,In_286,In_528);
nor U2640 (N_2640,In_991,In_1382);
nand U2641 (N_2641,In_116,In_1343);
nand U2642 (N_2642,In_1201,In_1689);
xnor U2643 (N_2643,In_409,In_802);
nor U2644 (N_2644,In_1462,In_1631);
or U2645 (N_2645,In_1074,In_1534);
or U2646 (N_2646,In_870,In_1449);
nor U2647 (N_2647,In_1144,In_1112);
nor U2648 (N_2648,In_158,In_1315);
and U2649 (N_2649,In_1507,In_802);
or U2650 (N_2650,In_1853,In_734);
and U2651 (N_2651,In_1231,In_1892);
and U2652 (N_2652,In_1323,In_155);
nand U2653 (N_2653,In_677,In_1113);
or U2654 (N_2654,In_1206,In_171);
or U2655 (N_2655,In_1042,In_1951);
and U2656 (N_2656,In_1635,In_1733);
or U2657 (N_2657,In_141,In_924);
nand U2658 (N_2658,In_1577,In_71);
nand U2659 (N_2659,In_930,In_1625);
or U2660 (N_2660,In_32,In_1239);
and U2661 (N_2661,In_1281,In_1173);
or U2662 (N_2662,In_1264,In_1260);
nand U2663 (N_2663,In_624,In_759);
xnor U2664 (N_2664,In_1327,In_1996);
nor U2665 (N_2665,In_1023,In_1524);
nor U2666 (N_2666,In_1973,In_343);
and U2667 (N_2667,In_1718,In_1433);
and U2668 (N_2668,In_751,In_364);
and U2669 (N_2669,In_447,In_1413);
and U2670 (N_2670,In_710,In_1903);
and U2671 (N_2671,In_1169,In_1750);
or U2672 (N_2672,In_139,In_1342);
nor U2673 (N_2673,In_1293,In_1381);
nand U2674 (N_2674,In_315,In_1546);
nor U2675 (N_2675,In_1057,In_1845);
nand U2676 (N_2676,In_102,In_984);
and U2677 (N_2677,In_806,In_450);
or U2678 (N_2678,In_625,In_430);
and U2679 (N_2679,In_1127,In_994);
and U2680 (N_2680,In_989,In_1690);
and U2681 (N_2681,In_1542,In_10);
nand U2682 (N_2682,In_239,In_659);
xor U2683 (N_2683,In_790,In_1613);
or U2684 (N_2684,In_883,In_880);
nor U2685 (N_2685,In_1911,In_750);
nand U2686 (N_2686,In_97,In_1386);
and U2687 (N_2687,In_153,In_193);
or U2688 (N_2688,In_1081,In_1485);
or U2689 (N_2689,In_189,In_1721);
nand U2690 (N_2690,In_1370,In_383);
and U2691 (N_2691,In_814,In_25);
or U2692 (N_2692,In_218,In_351);
nand U2693 (N_2693,In_1216,In_175);
or U2694 (N_2694,In_1590,In_939);
nor U2695 (N_2695,In_592,In_1059);
or U2696 (N_2696,In_701,In_773);
xor U2697 (N_2697,In_380,In_1700);
and U2698 (N_2698,In_1750,In_992);
or U2699 (N_2699,In_857,In_184);
nor U2700 (N_2700,In_1226,In_1425);
xnor U2701 (N_2701,In_1273,In_1383);
or U2702 (N_2702,In_1191,In_1826);
and U2703 (N_2703,In_427,In_766);
and U2704 (N_2704,In_1354,In_157);
and U2705 (N_2705,In_230,In_1369);
nor U2706 (N_2706,In_1407,In_692);
or U2707 (N_2707,In_1370,In_845);
nor U2708 (N_2708,In_1267,In_1166);
and U2709 (N_2709,In_436,In_1829);
nor U2710 (N_2710,In_1409,In_1424);
nand U2711 (N_2711,In_1175,In_1788);
nand U2712 (N_2712,In_1261,In_1310);
nand U2713 (N_2713,In_792,In_195);
or U2714 (N_2714,In_1306,In_1811);
xnor U2715 (N_2715,In_1892,In_999);
nand U2716 (N_2716,In_1929,In_1783);
nand U2717 (N_2717,In_1809,In_1813);
and U2718 (N_2718,In_724,In_1546);
nor U2719 (N_2719,In_528,In_372);
nor U2720 (N_2720,In_1293,In_244);
and U2721 (N_2721,In_1202,In_1786);
or U2722 (N_2722,In_880,In_450);
and U2723 (N_2723,In_1581,In_447);
nand U2724 (N_2724,In_387,In_517);
nor U2725 (N_2725,In_1136,In_1500);
and U2726 (N_2726,In_1184,In_1220);
or U2727 (N_2727,In_785,In_1866);
and U2728 (N_2728,In_1624,In_139);
xnor U2729 (N_2729,In_1626,In_131);
nor U2730 (N_2730,In_1566,In_1657);
and U2731 (N_2731,In_29,In_1050);
nor U2732 (N_2732,In_1364,In_656);
and U2733 (N_2733,In_1076,In_1106);
nor U2734 (N_2734,In_1274,In_1726);
and U2735 (N_2735,In_960,In_288);
nor U2736 (N_2736,In_1237,In_304);
and U2737 (N_2737,In_867,In_275);
nand U2738 (N_2738,In_1257,In_963);
and U2739 (N_2739,In_910,In_267);
nand U2740 (N_2740,In_1043,In_1208);
nor U2741 (N_2741,In_428,In_759);
nand U2742 (N_2742,In_759,In_1244);
nand U2743 (N_2743,In_41,In_1267);
nor U2744 (N_2744,In_1952,In_1518);
nand U2745 (N_2745,In_1209,In_1625);
and U2746 (N_2746,In_140,In_129);
or U2747 (N_2747,In_263,In_1305);
and U2748 (N_2748,In_31,In_187);
and U2749 (N_2749,In_1334,In_1484);
nor U2750 (N_2750,In_1929,In_1188);
nor U2751 (N_2751,In_313,In_714);
xnor U2752 (N_2752,In_1526,In_787);
or U2753 (N_2753,In_173,In_521);
nor U2754 (N_2754,In_1039,In_166);
and U2755 (N_2755,In_501,In_1089);
xnor U2756 (N_2756,In_1737,In_410);
xor U2757 (N_2757,In_718,In_197);
nor U2758 (N_2758,In_1894,In_884);
nor U2759 (N_2759,In_930,In_1200);
xnor U2760 (N_2760,In_1926,In_138);
xor U2761 (N_2761,In_221,In_338);
and U2762 (N_2762,In_840,In_1281);
nand U2763 (N_2763,In_143,In_1750);
or U2764 (N_2764,In_1634,In_1211);
xor U2765 (N_2765,In_622,In_837);
nor U2766 (N_2766,In_1865,In_1600);
or U2767 (N_2767,In_1040,In_336);
or U2768 (N_2768,In_1547,In_1077);
nand U2769 (N_2769,In_480,In_64);
and U2770 (N_2770,In_1412,In_1125);
and U2771 (N_2771,In_978,In_1626);
xor U2772 (N_2772,In_1109,In_886);
nor U2773 (N_2773,In_1095,In_986);
nor U2774 (N_2774,In_1999,In_1262);
nor U2775 (N_2775,In_1087,In_1095);
nand U2776 (N_2776,In_164,In_507);
nand U2777 (N_2777,In_381,In_1709);
nor U2778 (N_2778,In_1858,In_181);
nand U2779 (N_2779,In_375,In_1748);
or U2780 (N_2780,In_730,In_1227);
nand U2781 (N_2781,In_1237,In_1959);
nand U2782 (N_2782,In_1188,In_413);
and U2783 (N_2783,In_485,In_798);
nand U2784 (N_2784,In_1785,In_1739);
or U2785 (N_2785,In_1457,In_903);
and U2786 (N_2786,In_943,In_1099);
and U2787 (N_2787,In_1452,In_448);
and U2788 (N_2788,In_1349,In_1744);
and U2789 (N_2789,In_110,In_656);
and U2790 (N_2790,In_427,In_1816);
nor U2791 (N_2791,In_986,In_836);
nor U2792 (N_2792,In_402,In_1342);
or U2793 (N_2793,In_425,In_592);
nand U2794 (N_2794,In_659,In_665);
nand U2795 (N_2795,In_1280,In_174);
nor U2796 (N_2796,In_22,In_749);
and U2797 (N_2797,In_993,In_767);
nand U2798 (N_2798,In_1504,In_661);
or U2799 (N_2799,In_1688,In_705);
nor U2800 (N_2800,In_794,In_756);
and U2801 (N_2801,In_521,In_1300);
nor U2802 (N_2802,In_1613,In_1906);
or U2803 (N_2803,In_236,In_1155);
nor U2804 (N_2804,In_1512,In_1774);
nor U2805 (N_2805,In_1738,In_143);
and U2806 (N_2806,In_1484,In_729);
xor U2807 (N_2807,In_154,In_265);
or U2808 (N_2808,In_56,In_472);
nand U2809 (N_2809,In_142,In_717);
nor U2810 (N_2810,In_1047,In_677);
nor U2811 (N_2811,In_179,In_775);
or U2812 (N_2812,In_921,In_1952);
nor U2813 (N_2813,In_954,In_524);
nand U2814 (N_2814,In_1366,In_417);
nor U2815 (N_2815,In_1395,In_252);
or U2816 (N_2816,In_1694,In_333);
nor U2817 (N_2817,In_1361,In_1074);
or U2818 (N_2818,In_858,In_404);
and U2819 (N_2819,In_1177,In_1094);
and U2820 (N_2820,In_655,In_788);
or U2821 (N_2821,In_398,In_372);
xnor U2822 (N_2822,In_506,In_1903);
or U2823 (N_2823,In_1444,In_91);
nor U2824 (N_2824,In_306,In_1990);
nor U2825 (N_2825,In_288,In_271);
nand U2826 (N_2826,In_784,In_245);
or U2827 (N_2827,In_1792,In_1441);
and U2828 (N_2828,In_217,In_1412);
and U2829 (N_2829,In_588,In_32);
nand U2830 (N_2830,In_1723,In_1239);
nand U2831 (N_2831,In_1827,In_50);
xnor U2832 (N_2832,In_903,In_1759);
and U2833 (N_2833,In_515,In_548);
or U2834 (N_2834,In_860,In_1313);
and U2835 (N_2835,In_1979,In_1813);
nand U2836 (N_2836,In_1725,In_700);
or U2837 (N_2837,In_1191,In_156);
and U2838 (N_2838,In_946,In_1414);
and U2839 (N_2839,In_1437,In_1951);
nor U2840 (N_2840,In_594,In_1642);
or U2841 (N_2841,In_634,In_1693);
and U2842 (N_2842,In_100,In_1409);
nand U2843 (N_2843,In_1863,In_1329);
nand U2844 (N_2844,In_719,In_1528);
nand U2845 (N_2845,In_426,In_1268);
or U2846 (N_2846,In_1673,In_645);
and U2847 (N_2847,In_1039,In_1624);
nor U2848 (N_2848,In_1607,In_780);
nand U2849 (N_2849,In_741,In_1610);
nor U2850 (N_2850,In_829,In_1294);
nor U2851 (N_2851,In_330,In_1908);
or U2852 (N_2852,In_1171,In_504);
nor U2853 (N_2853,In_1582,In_909);
and U2854 (N_2854,In_1045,In_517);
and U2855 (N_2855,In_281,In_151);
xor U2856 (N_2856,In_1520,In_1304);
nand U2857 (N_2857,In_1041,In_1882);
and U2858 (N_2858,In_608,In_1469);
and U2859 (N_2859,In_1330,In_1877);
and U2860 (N_2860,In_1512,In_1167);
nand U2861 (N_2861,In_1075,In_1368);
and U2862 (N_2862,In_1236,In_918);
and U2863 (N_2863,In_147,In_1657);
nand U2864 (N_2864,In_1259,In_159);
and U2865 (N_2865,In_495,In_268);
nand U2866 (N_2866,In_978,In_1842);
nand U2867 (N_2867,In_1330,In_1204);
nor U2868 (N_2868,In_563,In_1613);
and U2869 (N_2869,In_1118,In_1001);
nand U2870 (N_2870,In_495,In_696);
nor U2871 (N_2871,In_1599,In_805);
nand U2872 (N_2872,In_22,In_497);
nand U2873 (N_2873,In_223,In_642);
and U2874 (N_2874,In_1162,In_759);
and U2875 (N_2875,In_352,In_342);
and U2876 (N_2876,In_908,In_689);
or U2877 (N_2877,In_1418,In_369);
nand U2878 (N_2878,In_281,In_1996);
nor U2879 (N_2879,In_406,In_1079);
nor U2880 (N_2880,In_158,In_1028);
nor U2881 (N_2881,In_1194,In_1701);
xnor U2882 (N_2882,In_1081,In_189);
nor U2883 (N_2883,In_1327,In_1631);
and U2884 (N_2884,In_1000,In_1825);
nor U2885 (N_2885,In_1570,In_1727);
nand U2886 (N_2886,In_783,In_501);
or U2887 (N_2887,In_519,In_597);
nor U2888 (N_2888,In_691,In_1883);
or U2889 (N_2889,In_1368,In_736);
nand U2890 (N_2890,In_170,In_1709);
nand U2891 (N_2891,In_302,In_157);
nand U2892 (N_2892,In_1698,In_190);
and U2893 (N_2893,In_883,In_471);
or U2894 (N_2894,In_1957,In_671);
or U2895 (N_2895,In_1408,In_797);
nand U2896 (N_2896,In_1452,In_1436);
nand U2897 (N_2897,In_992,In_1815);
and U2898 (N_2898,In_1054,In_985);
nand U2899 (N_2899,In_34,In_1507);
or U2900 (N_2900,In_435,In_53);
nand U2901 (N_2901,In_559,In_855);
nor U2902 (N_2902,In_1038,In_1556);
nor U2903 (N_2903,In_1773,In_241);
nor U2904 (N_2904,In_1908,In_36);
nand U2905 (N_2905,In_448,In_1218);
xor U2906 (N_2906,In_1918,In_1513);
xnor U2907 (N_2907,In_7,In_416);
nand U2908 (N_2908,In_290,In_1265);
and U2909 (N_2909,In_786,In_1449);
or U2910 (N_2910,In_1849,In_1150);
or U2911 (N_2911,In_1758,In_577);
nand U2912 (N_2912,In_1273,In_748);
nand U2913 (N_2913,In_47,In_1628);
nand U2914 (N_2914,In_380,In_1336);
nor U2915 (N_2915,In_827,In_1271);
xor U2916 (N_2916,In_1521,In_1126);
and U2917 (N_2917,In_97,In_222);
nor U2918 (N_2918,In_368,In_894);
nor U2919 (N_2919,In_1305,In_1022);
nor U2920 (N_2920,In_33,In_1534);
nor U2921 (N_2921,In_1205,In_1472);
and U2922 (N_2922,In_655,In_658);
xor U2923 (N_2923,In_760,In_1480);
nor U2924 (N_2924,In_168,In_243);
and U2925 (N_2925,In_1162,In_898);
and U2926 (N_2926,In_607,In_1560);
or U2927 (N_2927,In_84,In_1607);
or U2928 (N_2928,In_825,In_741);
nor U2929 (N_2929,In_420,In_1743);
or U2930 (N_2930,In_210,In_121);
xor U2931 (N_2931,In_1515,In_722);
and U2932 (N_2932,In_108,In_867);
or U2933 (N_2933,In_689,In_1659);
nand U2934 (N_2934,In_1888,In_1954);
xnor U2935 (N_2935,In_296,In_1905);
nand U2936 (N_2936,In_1733,In_1410);
xor U2937 (N_2937,In_290,In_1904);
and U2938 (N_2938,In_854,In_1583);
xnor U2939 (N_2939,In_770,In_570);
nor U2940 (N_2940,In_103,In_262);
nand U2941 (N_2941,In_1947,In_1834);
xor U2942 (N_2942,In_800,In_1570);
xnor U2943 (N_2943,In_120,In_28);
and U2944 (N_2944,In_1140,In_795);
nor U2945 (N_2945,In_1518,In_397);
xnor U2946 (N_2946,In_662,In_1376);
and U2947 (N_2947,In_1177,In_434);
nor U2948 (N_2948,In_595,In_1708);
or U2949 (N_2949,In_1438,In_1989);
or U2950 (N_2950,In_1923,In_179);
and U2951 (N_2951,In_1498,In_1946);
nor U2952 (N_2952,In_1988,In_1091);
nor U2953 (N_2953,In_215,In_1939);
nor U2954 (N_2954,In_853,In_1549);
nor U2955 (N_2955,In_994,In_47);
nor U2956 (N_2956,In_1034,In_915);
xor U2957 (N_2957,In_1858,In_393);
nand U2958 (N_2958,In_533,In_1972);
and U2959 (N_2959,In_1431,In_1066);
or U2960 (N_2960,In_1063,In_1502);
and U2961 (N_2961,In_1532,In_1260);
and U2962 (N_2962,In_1808,In_1080);
xnor U2963 (N_2963,In_1143,In_1279);
or U2964 (N_2964,In_698,In_138);
nand U2965 (N_2965,In_1064,In_1676);
nand U2966 (N_2966,In_1310,In_1015);
and U2967 (N_2967,In_1848,In_1497);
xnor U2968 (N_2968,In_835,In_1491);
and U2969 (N_2969,In_1754,In_1953);
or U2970 (N_2970,In_1349,In_1544);
nor U2971 (N_2971,In_939,In_324);
nor U2972 (N_2972,In_718,In_1686);
and U2973 (N_2973,In_1122,In_1359);
nand U2974 (N_2974,In_148,In_1860);
xor U2975 (N_2975,In_958,In_1023);
nor U2976 (N_2976,In_1803,In_1977);
nor U2977 (N_2977,In_1683,In_29);
and U2978 (N_2978,In_542,In_289);
nand U2979 (N_2979,In_454,In_668);
nand U2980 (N_2980,In_1826,In_401);
xnor U2981 (N_2981,In_47,In_1608);
or U2982 (N_2982,In_965,In_990);
nand U2983 (N_2983,In_1943,In_36);
xor U2984 (N_2984,In_370,In_907);
nand U2985 (N_2985,In_1444,In_1942);
nor U2986 (N_2986,In_570,In_1445);
nand U2987 (N_2987,In_1740,In_660);
xnor U2988 (N_2988,In_389,In_1117);
nor U2989 (N_2989,In_1042,In_428);
nand U2990 (N_2990,In_1930,In_768);
and U2991 (N_2991,In_1721,In_848);
nor U2992 (N_2992,In_1114,In_1536);
nand U2993 (N_2993,In_1277,In_1177);
or U2994 (N_2994,In_309,In_1732);
nand U2995 (N_2995,In_603,In_1763);
and U2996 (N_2996,In_769,In_1249);
nand U2997 (N_2997,In_857,In_912);
or U2998 (N_2998,In_1293,In_301);
or U2999 (N_2999,In_1863,In_41);
and U3000 (N_3000,In_519,In_180);
and U3001 (N_3001,In_1114,In_1988);
xor U3002 (N_3002,In_1544,In_15);
and U3003 (N_3003,In_1212,In_1137);
or U3004 (N_3004,In_1619,In_135);
or U3005 (N_3005,In_1389,In_1001);
nand U3006 (N_3006,In_932,In_282);
nor U3007 (N_3007,In_300,In_1891);
and U3008 (N_3008,In_1386,In_1850);
nor U3009 (N_3009,In_799,In_1923);
or U3010 (N_3010,In_1718,In_169);
nor U3011 (N_3011,In_594,In_245);
or U3012 (N_3012,In_266,In_227);
nand U3013 (N_3013,In_1498,In_944);
nor U3014 (N_3014,In_246,In_625);
nand U3015 (N_3015,In_1483,In_171);
and U3016 (N_3016,In_1918,In_392);
and U3017 (N_3017,In_1368,In_624);
and U3018 (N_3018,In_1508,In_345);
nand U3019 (N_3019,In_674,In_1221);
nor U3020 (N_3020,In_247,In_1656);
nor U3021 (N_3021,In_1062,In_515);
nor U3022 (N_3022,In_928,In_1713);
or U3023 (N_3023,In_1821,In_1519);
or U3024 (N_3024,In_1935,In_494);
nand U3025 (N_3025,In_1690,In_1126);
or U3026 (N_3026,In_1470,In_1613);
nand U3027 (N_3027,In_1631,In_360);
nand U3028 (N_3028,In_409,In_512);
nor U3029 (N_3029,In_1259,In_1310);
or U3030 (N_3030,In_1813,In_377);
or U3031 (N_3031,In_448,In_1858);
and U3032 (N_3032,In_909,In_1205);
and U3033 (N_3033,In_467,In_1594);
and U3034 (N_3034,In_1827,In_49);
and U3035 (N_3035,In_243,In_1869);
nor U3036 (N_3036,In_1402,In_637);
nor U3037 (N_3037,In_1828,In_67);
nor U3038 (N_3038,In_45,In_1731);
nor U3039 (N_3039,In_1549,In_1490);
or U3040 (N_3040,In_974,In_196);
xnor U3041 (N_3041,In_1174,In_131);
xor U3042 (N_3042,In_842,In_990);
xor U3043 (N_3043,In_1969,In_949);
and U3044 (N_3044,In_1210,In_1140);
and U3045 (N_3045,In_1759,In_1903);
or U3046 (N_3046,In_215,In_606);
and U3047 (N_3047,In_171,In_1395);
nor U3048 (N_3048,In_1202,In_1361);
nand U3049 (N_3049,In_196,In_1974);
nor U3050 (N_3050,In_1360,In_38);
nor U3051 (N_3051,In_393,In_205);
nand U3052 (N_3052,In_1770,In_1709);
or U3053 (N_3053,In_249,In_1616);
or U3054 (N_3054,In_425,In_1202);
and U3055 (N_3055,In_718,In_1433);
nor U3056 (N_3056,In_179,In_395);
nor U3057 (N_3057,In_26,In_61);
nand U3058 (N_3058,In_1967,In_813);
and U3059 (N_3059,In_1309,In_1106);
nand U3060 (N_3060,In_1681,In_375);
xor U3061 (N_3061,In_1088,In_526);
nor U3062 (N_3062,In_1928,In_1508);
nand U3063 (N_3063,In_1326,In_272);
or U3064 (N_3064,In_116,In_1347);
xor U3065 (N_3065,In_70,In_1499);
nand U3066 (N_3066,In_219,In_1159);
and U3067 (N_3067,In_1077,In_1549);
and U3068 (N_3068,In_1812,In_738);
nor U3069 (N_3069,In_428,In_895);
and U3070 (N_3070,In_642,In_236);
and U3071 (N_3071,In_1577,In_1508);
and U3072 (N_3072,In_1892,In_1550);
nor U3073 (N_3073,In_1661,In_578);
nor U3074 (N_3074,In_525,In_721);
xor U3075 (N_3075,In_1679,In_916);
xor U3076 (N_3076,In_1560,In_360);
xor U3077 (N_3077,In_385,In_338);
nor U3078 (N_3078,In_1730,In_28);
nor U3079 (N_3079,In_1231,In_425);
and U3080 (N_3080,In_1575,In_842);
nor U3081 (N_3081,In_744,In_1055);
xnor U3082 (N_3082,In_963,In_683);
xnor U3083 (N_3083,In_1252,In_1672);
nand U3084 (N_3084,In_1687,In_1677);
nand U3085 (N_3085,In_1576,In_1858);
nand U3086 (N_3086,In_130,In_1244);
xnor U3087 (N_3087,In_1635,In_504);
xnor U3088 (N_3088,In_1166,In_906);
or U3089 (N_3089,In_655,In_88);
nand U3090 (N_3090,In_1909,In_48);
or U3091 (N_3091,In_507,In_1727);
nand U3092 (N_3092,In_117,In_780);
and U3093 (N_3093,In_988,In_588);
and U3094 (N_3094,In_1350,In_865);
nand U3095 (N_3095,In_1836,In_638);
and U3096 (N_3096,In_1435,In_344);
nor U3097 (N_3097,In_1445,In_1133);
nand U3098 (N_3098,In_374,In_1002);
nand U3099 (N_3099,In_231,In_286);
or U3100 (N_3100,In_379,In_785);
and U3101 (N_3101,In_1522,In_1344);
nor U3102 (N_3102,In_573,In_1325);
xor U3103 (N_3103,In_1467,In_229);
nand U3104 (N_3104,In_537,In_1970);
and U3105 (N_3105,In_1120,In_1138);
nor U3106 (N_3106,In_766,In_1332);
or U3107 (N_3107,In_699,In_1751);
nand U3108 (N_3108,In_759,In_58);
and U3109 (N_3109,In_687,In_1460);
nand U3110 (N_3110,In_1853,In_1250);
nor U3111 (N_3111,In_1187,In_172);
nor U3112 (N_3112,In_258,In_1602);
nor U3113 (N_3113,In_1079,In_1262);
nor U3114 (N_3114,In_1167,In_1471);
nor U3115 (N_3115,In_1036,In_860);
and U3116 (N_3116,In_990,In_1139);
nand U3117 (N_3117,In_1830,In_1096);
xor U3118 (N_3118,In_777,In_318);
and U3119 (N_3119,In_1586,In_67);
nor U3120 (N_3120,In_1529,In_320);
nor U3121 (N_3121,In_1416,In_1660);
and U3122 (N_3122,In_348,In_849);
nor U3123 (N_3123,In_390,In_505);
nand U3124 (N_3124,In_1151,In_907);
or U3125 (N_3125,In_1361,In_1081);
and U3126 (N_3126,In_1791,In_874);
nor U3127 (N_3127,In_1384,In_698);
nor U3128 (N_3128,In_1377,In_1261);
nor U3129 (N_3129,In_1344,In_1438);
nand U3130 (N_3130,In_606,In_602);
or U3131 (N_3131,In_1015,In_27);
or U3132 (N_3132,In_1604,In_595);
nor U3133 (N_3133,In_970,In_56);
or U3134 (N_3134,In_1957,In_1128);
or U3135 (N_3135,In_1110,In_239);
nand U3136 (N_3136,In_552,In_1628);
nand U3137 (N_3137,In_1917,In_0);
xnor U3138 (N_3138,In_1663,In_1399);
or U3139 (N_3139,In_1189,In_492);
nor U3140 (N_3140,In_1166,In_858);
nand U3141 (N_3141,In_646,In_927);
nor U3142 (N_3142,In_335,In_561);
or U3143 (N_3143,In_1285,In_145);
and U3144 (N_3144,In_378,In_382);
or U3145 (N_3145,In_1064,In_227);
nand U3146 (N_3146,In_1918,In_534);
xor U3147 (N_3147,In_49,In_97);
nand U3148 (N_3148,In_866,In_1027);
or U3149 (N_3149,In_120,In_1958);
or U3150 (N_3150,In_1991,In_2);
nand U3151 (N_3151,In_759,In_1571);
or U3152 (N_3152,In_66,In_771);
xnor U3153 (N_3153,In_183,In_1568);
and U3154 (N_3154,In_1397,In_1148);
xor U3155 (N_3155,In_1705,In_1062);
nor U3156 (N_3156,In_373,In_204);
or U3157 (N_3157,In_312,In_1210);
nor U3158 (N_3158,In_813,In_719);
and U3159 (N_3159,In_423,In_1233);
or U3160 (N_3160,In_134,In_388);
nor U3161 (N_3161,In_1957,In_429);
or U3162 (N_3162,In_1871,In_343);
nor U3163 (N_3163,In_1658,In_1564);
nand U3164 (N_3164,In_1879,In_559);
nor U3165 (N_3165,In_1675,In_1370);
nand U3166 (N_3166,In_808,In_1012);
nor U3167 (N_3167,In_856,In_776);
xnor U3168 (N_3168,In_479,In_607);
nor U3169 (N_3169,In_269,In_42);
and U3170 (N_3170,In_138,In_854);
or U3171 (N_3171,In_1066,In_955);
nor U3172 (N_3172,In_1399,In_426);
nor U3173 (N_3173,In_275,In_1179);
nand U3174 (N_3174,In_683,In_1821);
nand U3175 (N_3175,In_1819,In_1984);
nor U3176 (N_3176,In_415,In_1461);
or U3177 (N_3177,In_1011,In_1244);
and U3178 (N_3178,In_523,In_1064);
and U3179 (N_3179,In_1171,In_870);
xnor U3180 (N_3180,In_496,In_1568);
nand U3181 (N_3181,In_1341,In_1158);
nand U3182 (N_3182,In_298,In_23);
xnor U3183 (N_3183,In_786,In_876);
nand U3184 (N_3184,In_296,In_202);
nor U3185 (N_3185,In_328,In_830);
or U3186 (N_3186,In_1702,In_805);
and U3187 (N_3187,In_816,In_652);
or U3188 (N_3188,In_151,In_758);
or U3189 (N_3189,In_1992,In_231);
nand U3190 (N_3190,In_1921,In_629);
nor U3191 (N_3191,In_481,In_142);
xor U3192 (N_3192,In_1100,In_72);
xnor U3193 (N_3193,In_568,In_547);
and U3194 (N_3194,In_1824,In_1380);
and U3195 (N_3195,In_1067,In_1924);
nand U3196 (N_3196,In_536,In_689);
nand U3197 (N_3197,In_141,In_1497);
or U3198 (N_3198,In_1217,In_78);
or U3199 (N_3199,In_828,In_1609);
or U3200 (N_3200,In_494,In_1576);
nand U3201 (N_3201,In_1767,In_1577);
and U3202 (N_3202,In_519,In_1793);
nor U3203 (N_3203,In_1581,In_440);
or U3204 (N_3204,In_542,In_591);
xor U3205 (N_3205,In_1485,In_767);
nand U3206 (N_3206,In_803,In_582);
and U3207 (N_3207,In_569,In_127);
nand U3208 (N_3208,In_1286,In_1051);
and U3209 (N_3209,In_1312,In_1221);
and U3210 (N_3210,In_483,In_333);
nor U3211 (N_3211,In_1341,In_849);
and U3212 (N_3212,In_974,In_582);
nor U3213 (N_3213,In_1369,In_1969);
nand U3214 (N_3214,In_1745,In_639);
nand U3215 (N_3215,In_935,In_1069);
or U3216 (N_3216,In_1507,In_1415);
xnor U3217 (N_3217,In_1741,In_1255);
nand U3218 (N_3218,In_20,In_528);
nor U3219 (N_3219,In_1979,In_1550);
nand U3220 (N_3220,In_276,In_987);
or U3221 (N_3221,In_1775,In_1899);
nand U3222 (N_3222,In_640,In_668);
nor U3223 (N_3223,In_848,In_284);
nor U3224 (N_3224,In_1379,In_1076);
nor U3225 (N_3225,In_1627,In_310);
nor U3226 (N_3226,In_716,In_1329);
xor U3227 (N_3227,In_1988,In_1713);
and U3228 (N_3228,In_273,In_812);
or U3229 (N_3229,In_1897,In_1333);
nor U3230 (N_3230,In_1778,In_1706);
or U3231 (N_3231,In_1761,In_529);
or U3232 (N_3232,In_337,In_163);
and U3233 (N_3233,In_1533,In_1407);
nor U3234 (N_3234,In_1483,In_330);
or U3235 (N_3235,In_866,In_234);
nand U3236 (N_3236,In_1753,In_1570);
and U3237 (N_3237,In_444,In_1849);
nor U3238 (N_3238,In_156,In_453);
and U3239 (N_3239,In_1844,In_406);
xnor U3240 (N_3240,In_485,In_1677);
nor U3241 (N_3241,In_1026,In_1288);
and U3242 (N_3242,In_1747,In_1158);
nand U3243 (N_3243,In_651,In_935);
nor U3244 (N_3244,In_665,In_392);
nand U3245 (N_3245,In_435,In_1946);
or U3246 (N_3246,In_235,In_1287);
nand U3247 (N_3247,In_1619,In_933);
or U3248 (N_3248,In_1108,In_1836);
or U3249 (N_3249,In_1148,In_1125);
and U3250 (N_3250,In_811,In_1018);
nand U3251 (N_3251,In_1644,In_1612);
and U3252 (N_3252,In_1699,In_346);
nand U3253 (N_3253,In_1460,In_132);
or U3254 (N_3254,In_1715,In_27);
and U3255 (N_3255,In_656,In_1537);
nand U3256 (N_3256,In_1052,In_139);
and U3257 (N_3257,In_269,In_1574);
nor U3258 (N_3258,In_853,In_189);
xnor U3259 (N_3259,In_1179,In_1823);
and U3260 (N_3260,In_311,In_263);
nor U3261 (N_3261,In_397,In_1373);
nand U3262 (N_3262,In_632,In_44);
or U3263 (N_3263,In_1067,In_1792);
xnor U3264 (N_3264,In_1290,In_912);
nand U3265 (N_3265,In_1629,In_1769);
nor U3266 (N_3266,In_1613,In_203);
and U3267 (N_3267,In_1255,In_431);
and U3268 (N_3268,In_435,In_1256);
nand U3269 (N_3269,In_205,In_1489);
or U3270 (N_3270,In_366,In_1740);
nor U3271 (N_3271,In_1386,In_829);
nor U3272 (N_3272,In_1757,In_1213);
nor U3273 (N_3273,In_1837,In_562);
or U3274 (N_3274,In_1873,In_1577);
or U3275 (N_3275,In_1247,In_450);
and U3276 (N_3276,In_195,In_1034);
and U3277 (N_3277,In_1310,In_1424);
xnor U3278 (N_3278,In_1100,In_275);
nor U3279 (N_3279,In_591,In_76);
nand U3280 (N_3280,In_1639,In_1521);
and U3281 (N_3281,In_1719,In_1222);
or U3282 (N_3282,In_1384,In_1055);
or U3283 (N_3283,In_1876,In_1871);
xor U3284 (N_3284,In_1128,In_655);
nor U3285 (N_3285,In_1426,In_1449);
xor U3286 (N_3286,In_1060,In_1039);
nand U3287 (N_3287,In_532,In_991);
nor U3288 (N_3288,In_1289,In_1061);
nand U3289 (N_3289,In_0,In_1814);
nand U3290 (N_3290,In_1280,In_1019);
nand U3291 (N_3291,In_1755,In_1880);
nor U3292 (N_3292,In_595,In_756);
and U3293 (N_3293,In_1174,In_1781);
nor U3294 (N_3294,In_229,In_608);
nor U3295 (N_3295,In_577,In_1630);
nand U3296 (N_3296,In_1479,In_1810);
or U3297 (N_3297,In_1797,In_1547);
xor U3298 (N_3298,In_1869,In_1928);
nor U3299 (N_3299,In_606,In_402);
nor U3300 (N_3300,In_1836,In_885);
and U3301 (N_3301,In_1711,In_1357);
nand U3302 (N_3302,In_1279,In_482);
or U3303 (N_3303,In_1189,In_883);
and U3304 (N_3304,In_27,In_297);
nor U3305 (N_3305,In_1983,In_1917);
and U3306 (N_3306,In_1376,In_492);
xnor U3307 (N_3307,In_666,In_221);
nand U3308 (N_3308,In_928,In_839);
xnor U3309 (N_3309,In_169,In_1965);
nand U3310 (N_3310,In_1994,In_1107);
or U3311 (N_3311,In_1052,In_145);
nand U3312 (N_3312,In_790,In_197);
and U3313 (N_3313,In_133,In_827);
nor U3314 (N_3314,In_854,In_639);
nand U3315 (N_3315,In_1552,In_1998);
nor U3316 (N_3316,In_239,In_1779);
xnor U3317 (N_3317,In_817,In_677);
and U3318 (N_3318,In_838,In_1359);
nor U3319 (N_3319,In_1638,In_973);
or U3320 (N_3320,In_1131,In_276);
nor U3321 (N_3321,In_704,In_1675);
and U3322 (N_3322,In_699,In_1117);
xor U3323 (N_3323,In_734,In_1740);
or U3324 (N_3324,In_804,In_226);
and U3325 (N_3325,In_1686,In_1692);
and U3326 (N_3326,In_638,In_1694);
nand U3327 (N_3327,In_521,In_184);
and U3328 (N_3328,In_500,In_852);
or U3329 (N_3329,In_1115,In_630);
nand U3330 (N_3330,In_569,In_1400);
or U3331 (N_3331,In_57,In_1577);
and U3332 (N_3332,In_1722,In_1030);
or U3333 (N_3333,In_1284,In_1736);
nand U3334 (N_3334,In_245,In_1989);
or U3335 (N_3335,In_1521,In_612);
xnor U3336 (N_3336,In_1041,In_1188);
nor U3337 (N_3337,In_780,In_69);
and U3338 (N_3338,In_347,In_782);
or U3339 (N_3339,In_759,In_1777);
nand U3340 (N_3340,In_1430,In_1101);
and U3341 (N_3341,In_1283,In_276);
nor U3342 (N_3342,In_1000,In_671);
nand U3343 (N_3343,In_1963,In_1356);
xnor U3344 (N_3344,In_213,In_15);
nor U3345 (N_3345,In_1680,In_1971);
and U3346 (N_3346,In_1672,In_203);
nor U3347 (N_3347,In_431,In_1547);
nand U3348 (N_3348,In_950,In_1702);
xor U3349 (N_3349,In_1112,In_1109);
or U3350 (N_3350,In_1334,In_1317);
nand U3351 (N_3351,In_328,In_1185);
or U3352 (N_3352,In_793,In_1214);
nor U3353 (N_3353,In_1412,In_442);
nand U3354 (N_3354,In_1378,In_1379);
and U3355 (N_3355,In_358,In_1585);
nand U3356 (N_3356,In_743,In_165);
or U3357 (N_3357,In_111,In_677);
nor U3358 (N_3358,In_1769,In_1233);
nor U3359 (N_3359,In_251,In_287);
or U3360 (N_3360,In_229,In_749);
nand U3361 (N_3361,In_512,In_1633);
nor U3362 (N_3362,In_1007,In_1212);
xnor U3363 (N_3363,In_49,In_694);
nand U3364 (N_3364,In_1840,In_515);
nor U3365 (N_3365,In_1002,In_779);
and U3366 (N_3366,In_992,In_193);
nor U3367 (N_3367,In_1375,In_1864);
nor U3368 (N_3368,In_1124,In_1463);
and U3369 (N_3369,In_1050,In_1600);
nand U3370 (N_3370,In_1004,In_17);
nand U3371 (N_3371,In_705,In_1058);
or U3372 (N_3372,In_1617,In_386);
and U3373 (N_3373,In_999,In_1356);
or U3374 (N_3374,In_317,In_751);
and U3375 (N_3375,In_945,In_1673);
nor U3376 (N_3376,In_1960,In_182);
nor U3377 (N_3377,In_1272,In_1907);
xor U3378 (N_3378,In_860,In_1040);
or U3379 (N_3379,In_1028,In_499);
or U3380 (N_3380,In_1474,In_457);
or U3381 (N_3381,In_1485,In_1397);
nand U3382 (N_3382,In_588,In_1971);
or U3383 (N_3383,In_131,In_963);
nand U3384 (N_3384,In_437,In_658);
nand U3385 (N_3385,In_488,In_1873);
and U3386 (N_3386,In_1044,In_798);
nor U3387 (N_3387,In_1368,In_1613);
nor U3388 (N_3388,In_1401,In_1942);
nand U3389 (N_3389,In_1765,In_949);
or U3390 (N_3390,In_1021,In_961);
nand U3391 (N_3391,In_373,In_1911);
or U3392 (N_3392,In_512,In_253);
nor U3393 (N_3393,In_1711,In_1507);
nor U3394 (N_3394,In_310,In_894);
or U3395 (N_3395,In_265,In_417);
or U3396 (N_3396,In_468,In_791);
nor U3397 (N_3397,In_951,In_1409);
nand U3398 (N_3398,In_1115,In_334);
nor U3399 (N_3399,In_1997,In_1943);
nand U3400 (N_3400,In_154,In_1764);
nand U3401 (N_3401,In_1934,In_1696);
and U3402 (N_3402,In_1862,In_1905);
and U3403 (N_3403,In_1518,In_1651);
nand U3404 (N_3404,In_92,In_1332);
and U3405 (N_3405,In_643,In_1748);
xnor U3406 (N_3406,In_80,In_1797);
and U3407 (N_3407,In_1996,In_1621);
and U3408 (N_3408,In_1251,In_257);
or U3409 (N_3409,In_46,In_953);
xnor U3410 (N_3410,In_1589,In_931);
or U3411 (N_3411,In_1211,In_801);
or U3412 (N_3412,In_987,In_285);
nor U3413 (N_3413,In_1311,In_1890);
nor U3414 (N_3414,In_1150,In_1089);
and U3415 (N_3415,In_128,In_515);
or U3416 (N_3416,In_60,In_14);
xor U3417 (N_3417,In_392,In_594);
or U3418 (N_3418,In_20,In_1414);
nor U3419 (N_3419,In_1011,In_1703);
nor U3420 (N_3420,In_279,In_1932);
nand U3421 (N_3421,In_1149,In_1100);
nor U3422 (N_3422,In_327,In_370);
nand U3423 (N_3423,In_823,In_361);
xor U3424 (N_3424,In_162,In_163);
nand U3425 (N_3425,In_1772,In_1599);
or U3426 (N_3426,In_1552,In_346);
nor U3427 (N_3427,In_644,In_1866);
nand U3428 (N_3428,In_287,In_1950);
nor U3429 (N_3429,In_1498,In_1138);
and U3430 (N_3430,In_1635,In_584);
nor U3431 (N_3431,In_1902,In_1768);
and U3432 (N_3432,In_596,In_1142);
and U3433 (N_3433,In_1652,In_1281);
nand U3434 (N_3434,In_810,In_1903);
or U3435 (N_3435,In_1291,In_622);
xor U3436 (N_3436,In_359,In_48);
xor U3437 (N_3437,In_1077,In_704);
nor U3438 (N_3438,In_109,In_1686);
and U3439 (N_3439,In_0,In_1458);
or U3440 (N_3440,In_1799,In_430);
nor U3441 (N_3441,In_1873,In_1333);
and U3442 (N_3442,In_1472,In_1468);
or U3443 (N_3443,In_147,In_532);
or U3444 (N_3444,In_1092,In_509);
xor U3445 (N_3445,In_699,In_736);
nor U3446 (N_3446,In_240,In_1104);
and U3447 (N_3447,In_1280,In_823);
or U3448 (N_3448,In_1798,In_342);
nor U3449 (N_3449,In_1188,In_1329);
nor U3450 (N_3450,In_245,In_1811);
and U3451 (N_3451,In_1462,In_719);
nand U3452 (N_3452,In_1443,In_1916);
xor U3453 (N_3453,In_1084,In_849);
or U3454 (N_3454,In_452,In_729);
and U3455 (N_3455,In_1996,In_1377);
and U3456 (N_3456,In_997,In_1588);
xor U3457 (N_3457,In_801,In_1638);
or U3458 (N_3458,In_35,In_873);
nor U3459 (N_3459,In_405,In_442);
nor U3460 (N_3460,In_989,In_1354);
or U3461 (N_3461,In_1331,In_1086);
nand U3462 (N_3462,In_187,In_289);
or U3463 (N_3463,In_1237,In_423);
and U3464 (N_3464,In_211,In_894);
and U3465 (N_3465,In_1067,In_1101);
nor U3466 (N_3466,In_778,In_1741);
nor U3467 (N_3467,In_237,In_1487);
nor U3468 (N_3468,In_1582,In_62);
and U3469 (N_3469,In_1398,In_76);
nor U3470 (N_3470,In_1200,In_635);
or U3471 (N_3471,In_1211,In_1084);
nor U3472 (N_3472,In_644,In_407);
and U3473 (N_3473,In_1702,In_706);
nor U3474 (N_3474,In_1781,In_38);
nor U3475 (N_3475,In_236,In_1840);
nor U3476 (N_3476,In_1989,In_72);
and U3477 (N_3477,In_113,In_1756);
nand U3478 (N_3478,In_981,In_1436);
nor U3479 (N_3479,In_669,In_1582);
nand U3480 (N_3480,In_1622,In_831);
nand U3481 (N_3481,In_1988,In_790);
nor U3482 (N_3482,In_781,In_387);
nor U3483 (N_3483,In_332,In_888);
or U3484 (N_3484,In_1599,In_1480);
xnor U3485 (N_3485,In_85,In_1387);
and U3486 (N_3486,In_664,In_1905);
and U3487 (N_3487,In_830,In_1558);
nand U3488 (N_3488,In_1974,In_1434);
and U3489 (N_3489,In_760,In_913);
nor U3490 (N_3490,In_1668,In_686);
nand U3491 (N_3491,In_1679,In_1210);
nand U3492 (N_3492,In_1008,In_1541);
nand U3493 (N_3493,In_1251,In_1473);
nor U3494 (N_3494,In_1184,In_718);
nand U3495 (N_3495,In_300,In_836);
or U3496 (N_3496,In_1171,In_1800);
or U3497 (N_3497,In_1313,In_1140);
and U3498 (N_3498,In_1334,In_351);
nand U3499 (N_3499,In_482,In_65);
nor U3500 (N_3500,In_750,In_1368);
and U3501 (N_3501,In_1321,In_1074);
or U3502 (N_3502,In_635,In_927);
and U3503 (N_3503,In_1602,In_900);
nand U3504 (N_3504,In_1835,In_1575);
or U3505 (N_3505,In_918,In_4);
and U3506 (N_3506,In_1710,In_1612);
nor U3507 (N_3507,In_379,In_1557);
nor U3508 (N_3508,In_1596,In_1373);
and U3509 (N_3509,In_1693,In_306);
or U3510 (N_3510,In_682,In_515);
xnor U3511 (N_3511,In_31,In_919);
nand U3512 (N_3512,In_1443,In_1356);
nand U3513 (N_3513,In_1769,In_866);
or U3514 (N_3514,In_759,In_1256);
nand U3515 (N_3515,In_1933,In_1323);
and U3516 (N_3516,In_1063,In_1910);
xor U3517 (N_3517,In_1384,In_203);
nor U3518 (N_3518,In_1572,In_746);
nor U3519 (N_3519,In_626,In_780);
nor U3520 (N_3520,In_963,In_1298);
nand U3521 (N_3521,In_637,In_1162);
nand U3522 (N_3522,In_618,In_423);
nor U3523 (N_3523,In_988,In_1217);
or U3524 (N_3524,In_819,In_348);
or U3525 (N_3525,In_386,In_952);
and U3526 (N_3526,In_1054,In_684);
or U3527 (N_3527,In_226,In_450);
xnor U3528 (N_3528,In_280,In_1735);
nor U3529 (N_3529,In_905,In_1889);
or U3530 (N_3530,In_1196,In_844);
and U3531 (N_3531,In_1973,In_241);
xor U3532 (N_3532,In_779,In_213);
nor U3533 (N_3533,In_1694,In_1936);
nand U3534 (N_3534,In_586,In_1958);
nand U3535 (N_3535,In_369,In_1495);
and U3536 (N_3536,In_493,In_1579);
and U3537 (N_3537,In_161,In_1956);
or U3538 (N_3538,In_1919,In_1392);
and U3539 (N_3539,In_1013,In_1624);
and U3540 (N_3540,In_473,In_1416);
nor U3541 (N_3541,In_397,In_1897);
and U3542 (N_3542,In_1122,In_1111);
xnor U3543 (N_3543,In_1197,In_1231);
nand U3544 (N_3544,In_1538,In_756);
and U3545 (N_3545,In_1580,In_1237);
and U3546 (N_3546,In_1719,In_1226);
nand U3547 (N_3547,In_109,In_1903);
nand U3548 (N_3548,In_116,In_734);
or U3549 (N_3549,In_1694,In_111);
and U3550 (N_3550,In_1437,In_891);
and U3551 (N_3551,In_842,In_1026);
and U3552 (N_3552,In_674,In_1924);
and U3553 (N_3553,In_1958,In_1674);
xnor U3554 (N_3554,In_184,In_760);
or U3555 (N_3555,In_1392,In_585);
nor U3556 (N_3556,In_238,In_1113);
or U3557 (N_3557,In_1483,In_1400);
xnor U3558 (N_3558,In_788,In_679);
nor U3559 (N_3559,In_491,In_1394);
and U3560 (N_3560,In_576,In_1342);
or U3561 (N_3561,In_1459,In_1466);
nand U3562 (N_3562,In_1698,In_1255);
and U3563 (N_3563,In_141,In_797);
or U3564 (N_3564,In_1180,In_1408);
nor U3565 (N_3565,In_1273,In_22);
nand U3566 (N_3566,In_1157,In_220);
nand U3567 (N_3567,In_458,In_1578);
nor U3568 (N_3568,In_1740,In_1328);
nor U3569 (N_3569,In_1286,In_1211);
or U3570 (N_3570,In_230,In_1271);
and U3571 (N_3571,In_1507,In_1425);
and U3572 (N_3572,In_999,In_849);
nand U3573 (N_3573,In_1356,In_1319);
nor U3574 (N_3574,In_1104,In_698);
nand U3575 (N_3575,In_951,In_751);
and U3576 (N_3576,In_1975,In_36);
and U3577 (N_3577,In_1440,In_1301);
nor U3578 (N_3578,In_1286,In_220);
or U3579 (N_3579,In_1624,In_436);
nor U3580 (N_3580,In_462,In_1143);
and U3581 (N_3581,In_1332,In_1759);
or U3582 (N_3582,In_1099,In_537);
xor U3583 (N_3583,In_646,In_898);
and U3584 (N_3584,In_605,In_114);
nand U3585 (N_3585,In_607,In_1090);
xnor U3586 (N_3586,In_1442,In_881);
nor U3587 (N_3587,In_1324,In_617);
or U3588 (N_3588,In_224,In_1831);
or U3589 (N_3589,In_719,In_104);
nor U3590 (N_3590,In_696,In_1332);
or U3591 (N_3591,In_1905,In_1853);
and U3592 (N_3592,In_133,In_749);
nor U3593 (N_3593,In_1382,In_1763);
xnor U3594 (N_3594,In_191,In_271);
or U3595 (N_3595,In_1728,In_583);
nand U3596 (N_3596,In_1136,In_753);
nand U3597 (N_3597,In_1051,In_522);
or U3598 (N_3598,In_706,In_858);
nor U3599 (N_3599,In_907,In_325);
xor U3600 (N_3600,In_334,In_969);
nand U3601 (N_3601,In_1364,In_297);
and U3602 (N_3602,In_1110,In_1062);
and U3603 (N_3603,In_736,In_334);
nand U3604 (N_3604,In_237,In_574);
or U3605 (N_3605,In_559,In_62);
nor U3606 (N_3606,In_1229,In_1104);
and U3607 (N_3607,In_369,In_867);
nor U3608 (N_3608,In_1553,In_1354);
or U3609 (N_3609,In_391,In_260);
or U3610 (N_3610,In_959,In_1583);
nand U3611 (N_3611,In_585,In_516);
nand U3612 (N_3612,In_1559,In_517);
nand U3613 (N_3613,In_1480,In_1412);
nand U3614 (N_3614,In_1422,In_249);
and U3615 (N_3615,In_838,In_805);
nand U3616 (N_3616,In_183,In_1979);
and U3617 (N_3617,In_616,In_369);
nand U3618 (N_3618,In_1401,In_1192);
and U3619 (N_3619,In_1660,In_1827);
nand U3620 (N_3620,In_1414,In_1286);
and U3621 (N_3621,In_691,In_1933);
nand U3622 (N_3622,In_1447,In_367);
xor U3623 (N_3623,In_98,In_816);
nor U3624 (N_3624,In_437,In_1349);
and U3625 (N_3625,In_1447,In_908);
nor U3626 (N_3626,In_50,In_954);
and U3627 (N_3627,In_363,In_1702);
nor U3628 (N_3628,In_43,In_345);
nand U3629 (N_3629,In_178,In_235);
nor U3630 (N_3630,In_1112,In_385);
nand U3631 (N_3631,In_1076,In_1369);
nand U3632 (N_3632,In_588,In_1601);
nor U3633 (N_3633,In_703,In_1869);
or U3634 (N_3634,In_1639,In_1349);
or U3635 (N_3635,In_90,In_750);
nor U3636 (N_3636,In_1806,In_1849);
nand U3637 (N_3637,In_252,In_30);
xnor U3638 (N_3638,In_1465,In_1450);
and U3639 (N_3639,In_654,In_1159);
nand U3640 (N_3640,In_1533,In_1441);
nor U3641 (N_3641,In_877,In_296);
or U3642 (N_3642,In_1447,In_1083);
and U3643 (N_3643,In_98,In_1943);
or U3644 (N_3644,In_1801,In_1917);
xor U3645 (N_3645,In_420,In_1439);
or U3646 (N_3646,In_1415,In_1057);
and U3647 (N_3647,In_434,In_128);
nor U3648 (N_3648,In_1840,In_50);
and U3649 (N_3649,In_1194,In_1905);
xor U3650 (N_3650,In_617,In_1535);
nand U3651 (N_3651,In_424,In_1842);
nand U3652 (N_3652,In_650,In_733);
nor U3653 (N_3653,In_1127,In_1585);
or U3654 (N_3654,In_630,In_235);
nand U3655 (N_3655,In_1543,In_79);
nand U3656 (N_3656,In_1007,In_1093);
and U3657 (N_3657,In_1279,In_1157);
and U3658 (N_3658,In_1886,In_480);
and U3659 (N_3659,In_20,In_791);
and U3660 (N_3660,In_649,In_1610);
or U3661 (N_3661,In_1169,In_153);
or U3662 (N_3662,In_1813,In_1049);
or U3663 (N_3663,In_1155,In_1201);
nor U3664 (N_3664,In_1265,In_1700);
nand U3665 (N_3665,In_1749,In_1655);
xor U3666 (N_3666,In_513,In_309);
nand U3667 (N_3667,In_930,In_346);
and U3668 (N_3668,In_818,In_1725);
nor U3669 (N_3669,In_1258,In_984);
nor U3670 (N_3670,In_1797,In_1320);
or U3671 (N_3671,In_1734,In_1740);
and U3672 (N_3672,In_532,In_275);
and U3673 (N_3673,In_1167,In_1538);
nor U3674 (N_3674,In_899,In_957);
and U3675 (N_3675,In_855,In_516);
nand U3676 (N_3676,In_1594,In_1346);
and U3677 (N_3677,In_1270,In_1960);
nand U3678 (N_3678,In_1088,In_987);
nand U3679 (N_3679,In_292,In_1337);
nor U3680 (N_3680,In_202,In_1392);
or U3681 (N_3681,In_617,In_1340);
nor U3682 (N_3682,In_1075,In_911);
nand U3683 (N_3683,In_1782,In_730);
nand U3684 (N_3684,In_253,In_448);
or U3685 (N_3685,In_1417,In_1890);
or U3686 (N_3686,In_917,In_1373);
and U3687 (N_3687,In_1758,In_551);
nor U3688 (N_3688,In_890,In_1116);
and U3689 (N_3689,In_518,In_534);
and U3690 (N_3690,In_1878,In_823);
nand U3691 (N_3691,In_1619,In_517);
nand U3692 (N_3692,In_357,In_1986);
nand U3693 (N_3693,In_1383,In_1754);
or U3694 (N_3694,In_752,In_168);
nand U3695 (N_3695,In_701,In_627);
nand U3696 (N_3696,In_1640,In_1015);
nor U3697 (N_3697,In_1695,In_1158);
nand U3698 (N_3698,In_679,In_43);
xor U3699 (N_3699,In_1978,In_1019);
or U3700 (N_3700,In_1168,In_1327);
and U3701 (N_3701,In_1274,In_831);
and U3702 (N_3702,In_1756,In_920);
and U3703 (N_3703,In_467,In_1736);
nand U3704 (N_3704,In_131,In_1517);
nand U3705 (N_3705,In_225,In_1042);
and U3706 (N_3706,In_883,In_321);
or U3707 (N_3707,In_1023,In_1161);
or U3708 (N_3708,In_1173,In_403);
or U3709 (N_3709,In_988,In_940);
nand U3710 (N_3710,In_1115,In_398);
or U3711 (N_3711,In_501,In_1736);
nor U3712 (N_3712,In_62,In_281);
or U3713 (N_3713,In_1386,In_1330);
xnor U3714 (N_3714,In_916,In_488);
nand U3715 (N_3715,In_1138,In_542);
nand U3716 (N_3716,In_674,In_1441);
xnor U3717 (N_3717,In_535,In_1512);
nand U3718 (N_3718,In_1557,In_231);
nand U3719 (N_3719,In_965,In_932);
or U3720 (N_3720,In_114,In_798);
and U3721 (N_3721,In_1397,In_1635);
nand U3722 (N_3722,In_634,In_1945);
or U3723 (N_3723,In_1796,In_1771);
or U3724 (N_3724,In_1402,In_903);
xnor U3725 (N_3725,In_1210,In_1459);
or U3726 (N_3726,In_149,In_1388);
nor U3727 (N_3727,In_593,In_293);
xor U3728 (N_3728,In_335,In_1941);
and U3729 (N_3729,In_1236,In_642);
nor U3730 (N_3730,In_1571,In_914);
nor U3731 (N_3731,In_1256,In_66);
nand U3732 (N_3732,In_1307,In_554);
and U3733 (N_3733,In_1940,In_238);
nor U3734 (N_3734,In_1947,In_765);
nor U3735 (N_3735,In_1859,In_1641);
nand U3736 (N_3736,In_785,In_1103);
nand U3737 (N_3737,In_1899,In_1694);
nor U3738 (N_3738,In_1789,In_1948);
or U3739 (N_3739,In_19,In_1534);
nor U3740 (N_3740,In_1221,In_1023);
or U3741 (N_3741,In_1150,In_330);
xnor U3742 (N_3742,In_183,In_488);
nand U3743 (N_3743,In_1192,In_311);
or U3744 (N_3744,In_225,In_873);
or U3745 (N_3745,In_1618,In_1685);
nand U3746 (N_3746,In_1628,In_1538);
or U3747 (N_3747,In_615,In_881);
nor U3748 (N_3748,In_1784,In_30);
or U3749 (N_3749,In_64,In_1159);
and U3750 (N_3750,In_1013,In_1834);
xnor U3751 (N_3751,In_23,In_125);
and U3752 (N_3752,In_148,In_1776);
or U3753 (N_3753,In_1491,In_782);
nor U3754 (N_3754,In_468,In_109);
xor U3755 (N_3755,In_1646,In_373);
or U3756 (N_3756,In_197,In_386);
and U3757 (N_3757,In_1369,In_1356);
and U3758 (N_3758,In_870,In_602);
xor U3759 (N_3759,In_1923,In_411);
or U3760 (N_3760,In_190,In_1325);
or U3761 (N_3761,In_765,In_703);
or U3762 (N_3762,In_890,In_764);
nand U3763 (N_3763,In_800,In_1027);
nand U3764 (N_3764,In_798,In_340);
xor U3765 (N_3765,In_614,In_637);
nand U3766 (N_3766,In_890,In_569);
and U3767 (N_3767,In_515,In_1405);
nand U3768 (N_3768,In_1386,In_910);
xnor U3769 (N_3769,In_1412,In_389);
nand U3770 (N_3770,In_464,In_967);
nand U3771 (N_3771,In_1283,In_1857);
or U3772 (N_3772,In_1525,In_813);
or U3773 (N_3773,In_159,In_1241);
or U3774 (N_3774,In_741,In_1915);
nand U3775 (N_3775,In_338,In_704);
nand U3776 (N_3776,In_475,In_1237);
xnor U3777 (N_3777,In_95,In_402);
nand U3778 (N_3778,In_1332,In_902);
and U3779 (N_3779,In_1460,In_180);
nor U3780 (N_3780,In_1036,In_51);
or U3781 (N_3781,In_282,In_422);
or U3782 (N_3782,In_1654,In_1988);
or U3783 (N_3783,In_1433,In_1100);
nor U3784 (N_3784,In_194,In_1088);
nor U3785 (N_3785,In_1255,In_266);
and U3786 (N_3786,In_832,In_613);
and U3787 (N_3787,In_1664,In_1685);
nor U3788 (N_3788,In_737,In_1722);
nor U3789 (N_3789,In_21,In_1205);
or U3790 (N_3790,In_1905,In_853);
and U3791 (N_3791,In_1751,In_1455);
and U3792 (N_3792,In_1471,In_1737);
xnor U3793 (N_3793,In_464,In_1764);
and U3794 (N_3794,In_915,In_239);
xnor U3795 (N_3795,In_1187,In_967);
nand U3796 (N_3796,In_523,In_1117);
nand U3797 (N_3797,In_1904,In_1136);
and U3798 (N_3798,In_367,In_7);
and U3799 (N_3799,In_425,In_942);
or U3800 (N_3800,In_372,In_600);
xnor U3801 (N_3801,In_162,In_1701);
nand U3802 (N_3802,In_627,In_1986);
nor U3803 (N_3803,In_54,In_588);
nand U3804 (N_3804,In_1511,In_1486);
and U3805 (N_3805,In_647,In_226);
and U3806 (N_3806,In_652,In_719);
nand U3807 (N_3807,In_595,In_131);
xor U3808 (N_3808,In_1932,In_1695);
nand U3809 (N_3809,In_1955,In_955);
nor U3810 (N_3810,In_738,In_1071);
or U3811 (N_3811,In_383,In_2);
and U3812 (N_3812,In_772,In_571);
and U3813 (N_3813,In_1202,In_580);
or U3814 (N_3814,In_1282,In_86);
nor U3815 (N_3815,In_765,In_1458);
and U3816 (N_3816,In_56,In_93);
nand U3817 (N_3817,In_214,In_396);
xnor U3818 (N_3818,In_1903,In_990);
or U3819 (N_3819,In_595,In_1876);
or U3820 (N_3820,In_375,In_1220);
nand U3821 (N_3821,In_858,In_570);
nor U3822 (N_3822,In_982,In_1864);
nand U3823 (N_3823,In_204,In_1231);
nand U3824 (N_3824,In_791,In_604);
or U3825 (N_3825,In_1298,In_494);
nor U3826 (N_3826,In_546,In_764);
or U3827 (N_3827,In_129,In_104);
and U3828 (N_3828,In_112,In_1235);
nor U3829 (N_3829,In_1320,In_626);
and U3830 (N_3830,In_1743,In_1957);
nor U3831 (N_3831,In_1669,In_1356);
and U3832 (N_3832,In_580,In_1057);
nor U3833 (N_3833,In_452,In_697);
and U3834 (N_3834,In_1532,In_1023);
nor U3835 (N_3835,In_850,In_379);
nor U3836 (N_3836,In_733,In_1201);
or U3837 (N_3837,In_1994,In_272);
nand U3838 (N_3838,In_1542,In_957);
or U3839 (N_3839,In_1815,In_1596);
and U3840 (N_3840,In_263,In_711);
or U3841 (N_3841,In_1182,In_1266);
nand U3842 (N_3842,In_1280,In_25);
or U3843 (N_3843,In_1936,In_1871);
xnor U3844 (N_3844,In_364,In_390);
nor U3845 (N_3845,In_1882,In_773);
nor U3846 (N_3846,In_1250,In_1388);
nand U3847 (N_3847,In_930,In_925);
nor U3848 (N_3848,In_958,In_1496);
nor U3849 (N_3849,In_1488,In_1391);
nand U3850 (N_3850,In_356,In_1172);
or U3851 (N_3851,In_1535,In_1956);
and U3852 (N_3852,In_996,In_334);
or U3853 (N_3853,In_921,In_776);
nor U3854 (N_3854,In_1820,In_357);
nor U3855 (N_3855,In_499,In_484);
and U3856 (N_3856,In_1891,In_1987);
and U3857 (N_3857,In_1580,In_1754);
xnor U3858 (N_3858,In_159,In_441);
xnor U3859 (N_3859,In_1797,In_47);
xor U3860 (N_3860,In_1784,In_381);
nor U3861 (N_3861,In_1395,In_1222);
and U3862 (N_3862,In_1407,In_112);
and U3863 (N_3863,In_1297,In_439);
and U3864 (N_3864,In_990,In_336);
and U3865 (N_3865,In_1975,In_839);
or U3866 (N_3866,In_1926,In_1039);
or U3867 (N_3867,In_108,In_639);
or U3868 (N_3868,In_174,In_328);
or U3869 (N_3869,In_1771,In_1815);
and U3870 (N_3870,In_1807,In_1842);
and U3871 (N_3871,In_201,In_1624);
nand U3872 (N_3872,In_746,In_75);
nand U3873 (N_3873,In_1634,In_161);
nand U3874 (N_3874,In_83,In_1557);
and U3875 (N_3875,In_903,In_1061);
or U3876 (N_3876,In_1653,In_896);
nand U3877 (N_3877,In_452,In_1335);
or U3878 (N_3878,In_971,In_220);
and U3879 (N_3879,In_321,In_1840);
nand U3880 (N_3880,In_1396,In_252);
nor U3881 (N_3881,In_1405,In_1728);
nor U3882 (N_3882,In_1040,In_265);
or U3883 (N_3883,In_132,In_936);
xnor U3884 (N_3884,In_1343,In_243);
nor U3885 (N_3885,In_771,In_1649);
and U3886 (N_3886,In_41,In_1297);
or U3887 (N_3887,In_1664,In_1766);
nand U3888 (N_3888,In_1107,In_1511);
nor U3889 (N_3889,In_250,In_1343);
or U3890 (N_3890,In_350,In_1018);
and U3891 (N_3891,In_1665,In_923);
and U3892 (N_3892,In_1627,In_29);
nor U3893 (N_3893,In_417,In_812);
nor U3894 (N_3894,In_49,In_285);
nor U3895 (N_3895,In_1601,In_1560);
nor U3896 (N_3896,In_1980,In_1517);
or U3897 (N_3897,In_1042,In_1103);
nand U3898 (N_3898,In_1855,In_1714);
and U3899 (N_3899,In_1946,In_1947);
nor U3900 (N_3900,In_786,In_736);
nor U3901 (N_3901,In_1756,In_966);
nor U3902 (N_3902,In_1319,In_1431);
nor U3903 (N_3903,In_385,In_464);
xnor U3904 (N_3904,In_1083,In_165);
nand U3905 (N_3905,In_1897,In_972);
and U3906 (N_3906,In_1675,In_177);
and U3907 (N_3907,In_875,In_957);
or U3908 (N_3908,In_1707,In_1964);
and U3909 (N_3909,In_362,In_1419);
or U3910 (N_3910,In_742,In_497);
nand U3911 (N_3911,In_1532,In_291);
xnor U3912 (N_3912,In_704,In_1948);
and U3913 (N_3913,In_193,In_187);
or U3914 (N_3914,In_204,In_1566);
or U3915 (N_3915,In_810,In_140);
nand U3916 (N_3916,In_1461,In_596);
nor U3917 (N_3917,In_387,In_896);
and U3918 (N_3918,In_228,In_351);
and U3919 (N_3919,In_239,In_1667);
nor U3920 (N_3920,In_13,In_1049);
nor U3921 (N_3921,In_571,In_973);
nor U3922 (N_3922,In_88,In_1147);
or U3923 (N_3923,In_1431,In_465);
nor U3924 (N_3924,In_287,In_963);
or U3925 (N_3925,In_1231,In_1115);
or U3926 (N_3926,In_1418,In_1255);
or U3927 (N_3927,In_655,In_1613);
nor U3928 (N_3928,In_1325,In_771);
xor U3929 (N_3929,In_1938,In_1374);
nor U3930 (N_3930,In_1223,In_1367);
nor U3931 (N_3931,In_1797,In_1399);
nor U3932 (N_3932,In_1747,In_642);
and U3933 (N_3933,In_805,In_1898);
nand U3934 (N_3934,In_1318,In_465);
and U3935 (N_3935,In_404,In_753);
and U3936 (N_3936,In_738,In_1387);
xnor U3937 (N_3937,In_1108,In_1211);
and U3938 (N_3938,In_272,In_1747);
and U3939 (N_3939,In_1613,In_609);
and U3940 (N_3940,In_1074,In_1729);
nor U3941 (N_3941,In_872,In_262);
or U3942 (N_3942,In_690,In_1528);
or U3943 (N_3943,In_1987,In_1983);
nand U3944 (N_3944,In_1244,In_1243);
or U3945 (N_3945,In_310,In_1058);
nor U3946 (N_3946,In_762,In_73);
or U3947 (N_3947,In_157,In_392);
or U3948 (N_3948,In_1157,In_1076);
or U3949 (N_3949,In_527,In_1455);
and U3950 (N_3950,In_153,In_948);
nor U3951 (N_3951,In_453,In_394);
and U3952 (N_3952,In_890,In_243);
nand U3953 (N_3953,In_42,In_1167);
nor U3954 (N_3954,In_157,In_1403);
nand U3955 (N_3955,In_1792,In_1814);
nor U3956 (N_3956,In_1724,In_1020);
or U3957 (N_3957,In_413,In_1102);
nand U3958 (N_3958,In_1234,In_6);
nor U3959 (N_3959,In_118,In_1464);
or U3960 (N_3960,In_578,In_966);
and U3961 (N_3961,In_334,In_645);
nor U3962 (N_3962,In_50,In_804);
or U3963 (N_3963,In_29,In_340);
xor U3964 (N_3964,In_1154,In_1070);
nand U3965 (N_3965,In_459,In_1595);
or U3966 (N_3966,In_1410,In_1804);
xnor U3967 (N_3967,In_30,In_625);
xor U3968 (N_3968,In_538,In_1507);
nand U3969 (N_3969,In_593,In_874);
or U3970 (N_3970,In_1282,In_1261);
or U3971 (N_3971,In_1890,In_593);
and U3972 (N_3972,In_917,In_1173);
nand U3973 (N_3973,In_1638,In_1597);
and U3974 (N_3974,In_1607,In_252);
nor U3975 (N_3975,In_1335,In_36);
and U3976 (N_3976,In_343,In_98);
nor U3977 (N_3977,In_31,In_371);
nand U3978 (N_3978,In_193,In_1042);
or U3979 (N_3979,In_1449,In_199);
or U3980 (N_3980,In_1099,In_1347);
nand U3981 (N_3981,In_1334,In_1976);
and U3982 (N_3982,In_1448,In_1274);
nor U3983 (N_3983,In_1876,In_55);
nand U3984 (N_3984,In_174,In_623);
or U3985 (N_3985,In_4,In_694);
or U3986 (N_3986,In_430,In_182);
and U3987 (N_3987,In_1707,In_1192);
nor U3988 (N_3988,In_98,In_344);
nor U3989 (N_3989,In_589,In_1863);
and U3990 (N_3990,In_1952,In_1800);
nand U3991 (N_3991,In_1411,In_1842);
and U3992 (N_3992,In_1904,In_430);
and U3993 (N_3993,In_133,In_774);
or U3994 (N_3994,In_164,In_1410);
nand U3995 (N_3995,In_760,In_1095);
nor U3996 (N_3996,In_506,In_242);
or U3997 (N_3997,In_1903,In_171);
nand U3998 (N_3998,In_82,In_1930);
nand U3999 (N_3999,In_329,In_55);
or U4000 (N_4000,N_2675,N_974);
and U4001 (N_4001,N_2205,N_256);
nor U4002 (N_4002,N_78,N_1072);
nand U4003 (N_4003,N_1907,N_3126);
and U4004 (N_4004,N_3076,N_2645);
nor U4005 (N_4005,N_647,N_1972);
nor U4006 (N_4006,N_956,N_2619);
nor U4007 (N_4007,N_818,N_2056);
and U4008 (N_4008,N_369,N_1420);
and U4009 (N_4009,N_3254,N_2281);
or U4010 (N_4010,N_3532,N_1180);
nand U4011 (N_4011,N_3342,N_2431);
or U4012 (N_4012,N_2865,N_3110);
nor U4013 (N_4013,N_532,N_465);
xnor U4014 (N_4014,N_1755,N_1964);
or U4015 (N_4015,N_1871,N_559);
and U4016 (N_4016,N_49,N_594);
nand U4017 (N_4017,N_1024,N_1930);
nand U4018 (N_4018,N_1874,N_3673);
or U4019 (N_4019,N_3138,N_148);
nand U4020 (N_4020,N_2122,N_255);
and U4021 (N_4021,N_2459,N_1778);
or U4022 (N_4022,N_2683,N_3423);
or U4023 (N_4023,N_3063,N_3435);
or U4024 (N_4024,N_1571,N_2694);
nand U4025 (N_4025,N_2048,N_928);
and U4026 (N_4026,N_1173,N_1667);
nand U4027 (N_4027,N_3225,N_3051);
nor U4028 (N_4028,N_1139,N_247);
and U4029 (N_4029,N_2939,N_3330);
nor U4030 (N_4030,N_1982,N_19);
nor U4031 (N_4031,N_3128,N_3460);
nand U4032 (N_4032,N_3405,N_1376);
and U4033 (N_4033,N_2700,N_413);
or U4034 (N_4034,N_1606,N_2495);
nor U4035 (N_4035,N_1225,N_2266);
nor U4036 (N_4036,N_3355,N_519);
xnor U4037 (N_4037,N_3518,N_374);
nor U4038 (N_4038,N_1888,N_3359);
and U4039 (N_4039,N_2913,N_625);
and U4040 (N_4040,N_870,N_2077);
nand U4041 (N_4041,N_3323,N_1639);
nor U4042 (N_4042,N_2852,N_1697);
and U4043 (N_4043,N_30,N_2279);
xnor U4044 (N_4044,N_2305,N_3736);
nand U4045 (N_4045,N_2170,N_3089);
or U4046 (N_4046,N_1104,N_2859);
nand U4047 (N_4047,N_3226,N_3374);
nand U4048 (N_4048,N_2467,N_3615);
or U4049 (N_4049,N_3776,N_1545);
or U4050 (N_4050,N_2349,N_498);
or U4051 (N_4051,N_2214,N_1273);
or U4052 (N_4052,N_280,N_3061);
and U4053 (N_4053,N_2656,N_1719);
nor U4054 (N_4054,N_527,N_3838);
nor U4055 (N_4055,N_2709,N_3772);
nand U4056 (N_4056,N_2481,N_584);
nor U4057 (N_4057,N_2401,N_1211);
or U4058 (N_4058,N_1891,N_3340);
or U4059 (N_4059,N_3073,N_529);
nand U4060 (N_4060,N_2784,N_1241);
nor U4061 (N_4061,N_556,N_1412);
or U4062 (N_4062,N_1352,N_3955);
nand U4063 (N_4063,N_267,N_3792);
xnor U4064 (N_4064,N_3317,N_3723);
and U4065 (N_4065,N_1620,N_521);
and U4066 (N_4066,N_210,N_3148);
nand U4067 (N_4067,N_1353,N_874);
and U4068 (N_4068,N_1044,N_1265);
xnor U4069 (N_4069,N_848,N_2771);
and U4070 (N_4070,N_2502,N_1365);
nor U4071 (N_4071,N_2354,N_3593);
nand U4072 (N_4072,N_1762,N_2107);
and U4073 (N_4073,N_2579,N_2673);
and U4074 (N_4074,N_442,N_1790);
nor U4075 (N_4075,N_2958,N_1860);
or U4076 (N_4076,N_1708,N_2345);
nor U4077 (N_4077,N_2057,N_1506);
or U4078 (N_4078,N_3559,N_544);
nand U4079 (N_4079,N_1853,N_1730);
or U4080 (N_4080,N_2216,N_293);
nor U4081 (N_4081,N_2612,N_3490);
xnor U4082 (N_4082,N_2867,N_2571);
xnor U4083 (N_4083,N_543,N_2231);
and U4084 (N_4084,N_3217,N_2275);
and U4085 (N_4085,N_1390,N_3818);
and U4086 (N_4086,N_35,N_95);
nand U4087 (N_4087,N_2693,N_2319);
nor U4088 (N_4088,N_3788,N_3098);
and U4089 (N_4089,N_997,N_551);
nand U4090 (N_4090,N_645,N_3806);
xnor U4091 (N_4091,N_2485,N_3961);
or U4092 (N_4092,N_274,N_2026);
nand U4093 (N_4093,N_1187,N_3678);
nand U4094 (N_4094,N_2080,N_1880);
nand U4095 (N_4095,N_1430,N_3492);
nor U4096 (N_4096,N_3781,N_745);
nor U4097 (N_4097,N_545,N_3557);
nor U4098 (N_4098,N_2994,N_2154);
or U4099 (N_4099,N_422,N_2920);
nand U4100 (N_4100,N_1338,N_2220);
or U4101 (N_4101,N_3214,N_299);
and U4102 (N_4102,N_2510,N_445);
nor U4103 (N_4103,N_1734,N_2777);
and U4104 (N_4104,N_740,N_671);
nand U4105 (N_4105,N_1889,N_2418);
and U4106 (N_4106,N_2559,N_3988);
or U4107 (N_4107,N_2373,N_638);
and U4108 (N_4108,N_2261,N_3605);
or U4109 (N_4109,N_1236,N_124);
nor U4110 (N_4110,N_3270,N_2443);
nor U4111 (N_4111,N_3426,N_475);
nor U4112 (N_4112,N_2534,N_1086);
nand U4113 (N_4113,N_1100,N_1903);
nor U4114 (N_4114,N_1451,N_1392);
or U4115 (N_4115,N_3048,N_739);
nand U4116 (N_4116,N_2166,N_1824);
nand U4117 (N_4117,N_151,N_2762);
nand U4118 (N_4118,N_1154,N_1910);
nor U4119 (N_4119,N_1562,N_325);
xnor U4120 (N_4120,N_322,N_718);
or U4121 (N_4121,N_2049,N_2325);
or U4122 (N_4122,N_3994,N_765);
and U4123 (N_4123,N_2455,N_2397);
and U4124 (N_4124,N_3619,N_1028);
or U4125 (N_4125,N_636,N_3672);
or U4126 (N_4126,N_411,N_2490);
and U4127 (N_4127,N_224,N_3923);
nand U4128 (N_4128,N_1996,N_3630);
nor U4129 (N_4129,N_3863,N_2696);
and U4130 (N_4130,N_1660,N_3985);
or U4131 (N_4131,N_473,N_2248);
and U4132 (N_4132,N_3815,N_1497);
nor U4133 (N_4133,N_2361,N_811);
nand U4134 (N_4134,N_3978,N_2246);
and U4135 (N_4135,N_238,N_1189);
xor U4136 (N_4136,N_2607,N_3050);
nor U4137 (N_4137,N_1320,N_3348);
nor U4138 (N_4138,N_755,N_706);
and U4139 (N_4139,N_574,N_2989);
xnor U4140 (N_4140,N_3521,N_966);
nand U4141 (N_4141,N_2640,N_2488);
and U4142 (N_4142,N_441,N_3765);
or U4143 (N_4143,N_2189,N_3307);
and U4144 (N_4144,N_90,N_1752);
nor U4145 (N_4145,N_3041,N_1630);
or U4146 (N_4146,N_171,N_2536);
nand U4147 (N_4147,N_847,N_3925);
or U4148 (N_4148,N_1738,N_1635);
and U4149 (N_4149,N_2505,N_3478);
xor U4150 (N_4150,N_1707,N_2066);
and U4151 (N_4151,N_3387,N_3866);
nand U4152 (N_4152,N_1544,N_2429);
or U4153 (N_4153,N_2428,N_2394);
and U4154 (N_4154,N_3780,N_1686);
and U4155 (N_4155,N_589,N_3417);
xnor U4156 (N_4156,N_1629,N_3240);
xor U4157 (N_4157,N_468,N_2099);
nor U4158 (N_4158,N_2921,N_3439);
nor U4159 (N_4159,N_1372,N_885);
nand U4160 (N_4160,N_728,N_2366);
and U4161 (N_4161,N_526,N_142);
and U4162 (N_4162,N_2774,N_2837);
nand U4163 (N_4163,N_1572,N_1602);
nor U4164 (N_4164,N_3596,N_125);
or U4165 (N_4165,N_1049,N_2123);
and U4166 (N_4166,N_3173,N_3831);
or U4167 (N_4167,N_3802,N_994);
or U4168 (N_4168,N_1117,N_1048);
nand U4169 (N_4169,N_714,N_2436);
and U4170 (N_4170,N_1835,N_2672);
nand U4171 (N_4171,N_3113,N_1410);
nand U4172 (N_4172,N_2069,N_1865);
or U4173 (N_4173,N_2702,N_531);
or U4174 (N_4174,N_387,N_3789);
nand U4175 (N_4175,N_1956,N_752);
and U4176 (N_4176,N_3336,N_3652);
xor U4177 (N_4177,N_2503,N_723);
xor U4178 (N_4178,N_3731,N_784);
and U4179 (N_4179,N_3300,N_3305);
nor U4180 (N_4180,N_3064,N_738);
nor U4181 (N_4181,N_1401,N_2509);
or U4182 (N_4182,N_347,N_1302);
and U4183 (N_4183,N_1375,N_2890);
and U4184 (N_4184,N_3143,N_1632);
or U4185 (N_4185,N_1673,N_2937);
or U4186 (N_4186,N_2406,N_2295);
nand U4187 (N_4187,N_1033,N_3436);
and U4188 (N_4188,N_1188,N_695);
xnor U4189 (N_4189,N_2857,N_3140);
nand U4190 (N_4190,N_432,N_455);
and U4191 (N_4191,N_1128,N_702);
nor U4192 (N_4192,N_1423,N_993);
and U4193 (N_4193,N_65,N_1524);
nor U4194 (N_4194,N_3510,N_1022);
and U4195 (N_4195,N_169,N_1834);
nand U4196 (N_4196,N_1715,N_2622);
nor U4197 (N_4197,N_2601,N_1841);
nor U4198 (N_4198,N_190,N_3211);
nand U4199 (N_4199,N_2810,N_2054);
or U4200 (N_4200,N_1050,N_1201);
nand U4201 (N_4201,N_1567,N_93);
nor U4202 (N_4202,N_2750,N_458);
nor U4203 (N_4203,N_331,N_1504);
xnor U4204 (N_4204,N_1789,N_1368);
nand U4205 (N_4205,N_3090,N_1323);
or U4206 (N_4206,N_3389,N_1788);
or U4207 (N_4207,N_562,N_1809);
nand U4208 (N_4208,N_1592,N_3493);
nand U4209 (N_4209,N_2803,N_1733);
nor U4210 (N_4210,N_1175,N_2965);
nor U4211 (N_4211,N_836,N_2746);
and U4212 (N_4212,N_3095,N_2323);
nor U4213 (N_4213,N_878,N_3667);
or U4214 (N_4214,N_87,N_1194);
or U4215 (N_4215,N_2222,N_364);
and U4216 (N_4216,N_3738,N_121);
and U4217 (N_4217,N_1543,N_3103);
or U4218 (N_4218,N_217,N_2003);
or U4219 (N_4219,N_3564,N_1280);
or U4220 (N_4220,N_3413,N_1313);
and U4221 (N_4221,N_3695,N_2200);
nor U4222 (N_4222,N_769,N_292);
nand U4223 (N_4223,N_2703,N_3071);
nor U4224 (N_4224,N_1884,N_1713);
nand U4225 (N_4225,N_656,N_1291);
and U4226 (N_4226,N_491,N_2263);
or U4227 (N_4227,N_1052,N_3019);
or U4228 (N_4228,N_1932,N_2882);
nor U4229 (N_4229,N_3266,N_3821);
or U4230 (N_4230,N_1445,N_856);
and U4231 (N_4231,N_2941,N_338);
nand U4232 (N_4232,N_2648,N_3219);
nand U4233 (N_4233,N_1138,N_2800);
nor U4234 (N_4234,N_3373,N_3507);
nand U4235 (N_4235,N_1811,N_3491);
nand U4236 (N_4236,N_1108,N_1517);
or U4237 (N_4237,N_158,N_2821);
nor U4238 (N_4238,N_2741,N_972);
and U4239 (N_4239,N_620,N_1794);
or U4240 (N_4240,N_308,N_3085);
and U4241 (N_4241,N_1388,N_1627);
or U4242 (N_4242,N_2899,N_3385);
or U4243 (N_4243,N_1604,N_2024);
nand U4244 (N_4244,N_350,N_3749);
xnor U4245 (N_4245,N_1906,N_3252);
or U4246 (N_4246,N_3269,N_832);
or U4247 (N_4247,N_1127,N_3508);
nand U4248 (N_4248,N_297,N_1818);
or U4249 (N_4249,N_3798,N_1181);
and U4250 (N_4250,N_2868,N_1383);
or U4251 (N_4251,N_3598,N_3123);
and U4252 (N_4252,N_760,N_417);
xnor U4253 (N_4253,N_580,N_2288);
nand U4254 (N_4254,N_385,N_3794);
and U4255 (N_4255,N_1787,N_3752);
nand U4256 (N_4256,N_881,N_1478);
and U4257 (N_4257,N_1526,N_363);
nor U4258 (N_4258,N_3465,N_91);
nand U4259 (N_4259,N_3446,N_866);
xor U4260 (N_4260,N_687,N_1057);
and U4261 (N_4261,N_1021,N_3718);
xor U4262 (N_4262,N_52,N_3916);
or U4263 (N_4263,N_407,N_989);
nand U4264 (N_4264,N_2299,N_2738);
nand U4265 (N_4265,N_1147,N_2008);
nor U4266 (N_4266,N_2438,N_2637);
nand U4267 (N_4267,N_1110,N_237);
or U4268 (N_4268,N_2863,N_1118);
nor U4269 (N_4269,N_869,N_3993);
and U4270 (N_4270,N_362,N_1255);
and U4271 (N_4271,N_2864,N_2155);
and U4272 (N_4272,N_3227,N_606);
nor U4273 (N_4273,N_2846,N_2101);
and U4274 (N_4274,N_2789,N_3918);
nand U4275 (N_4275,N_1184,N_2258);
nor U4276 (N_4276,N_955,N_1271);
and U4277 (N_4277,N_3498,N_2879);
xor U4278 (N_4278,N_2290,N_2807);
xor U4279 (N_4279,N_1799,N_2063);
nor U4280 (N_4280,N_2479,N_516);
nand U4281 (N_4281,N_1547,N_2924);
and U4282 (N_4282,N_141,N_3854);
or U4283 (N_4283,N_1123,N_2360);
nand U4284 (N_4284,N_2194,N_1266);
nand U4285 (N_4285,N_1174,N_86);
or U4286 (N_4286,N_1665,N_2707);
nand U4287 (N_4287,N_3722,N_2188);
and U4288 (N_4288,N_1391,N_3475);
nand U4289 (N_4289,N_2966,N_787);
nand U4290 (N_4290,N_1825,N_3778);
and U4291 (N_4291,N_1908,N_826);
and U4292 (N_4292,N_2790,N_2710);
and U4293 (N_4293,N_2954,N_1074);
nor U4294 (N_4294,N_1309,N_412);
and U4295 (N_4295,N_2969,N_429);
nand U4296 (N_4296,N_1166,N_3182);
or U4297 (N_4297,N_3274,N_3972);
nand U4298 (N_4298,N_1239,N_286);
and U4299 (N_4299,N_2778,N_244);
or U4300 (N_4300,N_145,N_2179);
nor U4301 (N_4301,N_2620,N_3977);
and U4302 (N_4302,N_1092,N_737);
nand U4303 (N_4303,N_954,N_3281);
nor U4304 (N_4304,N_2595,N_3105);
or U4305 (N_4305,N_3891,N_2357);
nand U4306 (N_4306,N_754,N_2473);
or U4307 (N_4307,N_243,N_1505);
and U4308 (N_4308,N_3030,N_2313);
nand U4309 (N_4309,N_3263,N_508);
nor U4310 (N_4310,N_1863,N_3602);
and U4311 (N_4311,N_2486,N_174);
nand U4312 (N_4312,N_3017,N_3430);
nor U4313 (N_4313,N_3398,N_2819);
nor U4314 (N_4314,N_5,N_2096);
and U4315 (N_4315,N_996,N_3685);
nand U4316 (N_4316,N_3273,N_630);
nor U4317 (N_4317,N_2767,N_164);
nor U4318 (N_4318,N_613,N_3494);
nand U4319 (N_4319,N_253,N_821);
xnor U4320 (N_4320,N_1061,N_2644);
and U4321 (N_4321,N_1000,N_3660);
xor U4322 (N_4322,N_1915,N_40);
and U4323 (N_4323,N_733,N_709);
and U4324 (N_4324,N_712,N_1396);
and U4325 (N_4325,N_55,N_942);
nand U4326 (N_4326,N_1124,N_639);
nor U4327 (N_4327,N_2042,N_2755);
xor U4328 (N_4328,N_116,N_524);
and U4329 (N_4329,N_2392,N_3839);
nand U4330 (N_4330,N_260,N_3216);
nand U4331 (N_4331,N_214,N_1528);
nor U4332 (N_4332,N_1398,N_3309);
or U4333 (N_4333,N_2199,N_2591);
nand U4334 (N_4334,N_713,N_3989);
or U4335 (N_4335,N_367,N_2037);
and U4336 (N_4336,N_1218,N_3107);
or U4337 (N_4337,N_981,N_2991);
xor U4338 (N_4338,N_3466,N_397);
nand U4339 (N_4339,N_3449,N_1014);
nor U4340 (N_4340,N_3109,N_2453);
xnor U4341 (N_4341,N_2456,N_2267);
nand U4342 (N_4342,N_3811,N_3919);
or U4343 (N_4343,N_2412,N_2289);
or U4344 (N_4344,N_1862,N_2109);
nor U4345 (N_4345,N_2573,N_3774);
nor U4346 (N_4346,N_2368,N_3661);
or U4347 (N_4347,N_992,N_2927);
and U4348 (N_4348,N_1753,N_1917);
xor U4349 (N_4349,N_3577,N_1263);
or U4350 (N_4350,N_3745,N_219);
and U4351 (N_4351,N_1859,N_2827);
and U4352 (N_4352,N_747,N_941);
nor U4353 (N_4353,N_2236,N_1857);
and U4354 (N_4354,N_564,N_3618);
and U4355 (N_4355,N_1510,N_640);
and U4356 (N_4356,N_1955,N_1705);
nor U4357 (N_4357,N_2972,N_600);
and U4358 (N_4358,N_1991,N_3246);
xnor U4359 (N_4359,N_798,N_1395);
nor U4360 (N_4360,N_1468,N_225);
or U4361 (N_4361,N_2580,N_701);
and U4362 (N_4362,N_2282,N_3057);
nor U4363 (N_4363,N_2963,N_3550);
nand U4364 (N_4364,N_3820,N_150);
or U4365 (N_4365,N_3195,N_3529);
nand U4366 (N_4366,N_2105,N_3911);
and U4367 (N_4367,N_3683,N_1113);
and U4368 (N_4368,N_1570,N_3908);
nand U4369 (N_4369,N_262,N_398);
and U4370 (N_4370,N_857,N_227);
and U4371 (N_4371,N_2535,N_276);
xor U4372 (N_4372,N_665,N_1951);
xnor U4373 (N_4373,N_2022,N_2134);
nand U4374 (N_4374,N_915,N_690);
and U4375 (N_4375,N_2265,N_2785);
or U4376 (N_4376,N_2225,N_1680);
and U4377 (N_4377,N_3548,N_2206);
or U4378 (N_4378,N_2276,N_3689);
nor U4379 (N_4379,N_1591,N_1931);
xor U4380 (N_4380,N_1551,N_2217);
or U4381 (N_4381,N_3999,N_3003);
nand U4382 (N_4382,N_1011,N_3347);
or U4383 (N_4383,N_1696,N_3295);
nand U4384 (N_4384,N_1658,N_538);
or U4385 (N_4385,N_2404,N_3710);
and U4386 (N_4386,N_3310,N_1176);
xor U4387 (N_4387,N_3083,N_1831);
or U4388 (N_4388,N_390,N_321);
and U4389 (N_4389,N_812,N_2445);
or U4390 (N_4390,N_1162,N_753);
xor U4391 (N_4391,N_3023,N_456);
xnor U4392 (N_4392,N_1989,N_619);
nor U4393 (N_4393,N_3910,N_2984);
and U4394 (N_4394,N_2437,N_2760);
nor U4395 (N_4395,N_1923,N_3768);
or U4396 (N_4396,N_2666,N_2849);
nor U4397 (N_4397,N_3333,N_684);
xor U4398 (N_4398,N_83,N_1227);
or U4399 (N_4399,N_352,N_2469);
nand U4400 (N_4400,N_3280,N_1995);
nor U4401 (N_4401,N_88,N_791);
nor U4402 (N_4402,N_3422,N_2605);
nand U4403 (N_4403,N_1204,N_1852);
nand U4404 (N_4404,N_222,N_1185);
and U4405 (N_4405,N_3982,N_3517);
and U4406 (N_4406,N_978,N_1942);
nand U4407 (N_4407,N_2507,N_336);
and U4408 (N_4408,N_3489,N_780);
and U4409 (N_4409,N_136,N_1643);
and U4410 (N_4410,N_2321,N_2961);
nand U4411 (N_4411,N_2089,N_940);
or U4412 (N_4412,N_2938,N_552);
and U4413 (N_4413,N_3210,N_2748);
nor U4414 (N_4414,N_1858,N_2087);
or U4415 (N_4415,N_3975,N_1508);
xor U4416 (N_4416,N_3706,N_3328);
nor U4417 (N_4417,N_1533,N_187);
nand U4418 (N_4418,N_2341,N_2326);
and U4419 (N_4419,N_1896,N_1483);
nor U4420 (N_4420,N_616,N_1358);
nor U4421 (N_4421,N_3884,N_1749);
or U4422 (N_4422,N_1436,N_970);
nand U4423 (N_4423,N_3651,N_2862);
nor U4424 (N_4424,N_601,N_2268);
xnor U4425 (N_4425,N_1464,N_1971);
or U4426 (N_4426,N_2468,N_3862);
xor U4427 (N_4427,N_17,N_28);
and U4428 (N_4428,N_2190,N_511);
and U4429 (N_4429,N_3187,N_2235);
and U4430 (N_4430,N_3159,N_1812);
or U4431 (N_4431,N_1679,N_1531);
or U4432 (N_4432,N_1764,N_918);
xnor U4433 (N_4433,N_3202,N_2690);
or U4434 (N_4434,N_1652,N_3203);
nand U4435 (N_4435,N_1424,N_820);
nor U4436 (N_4436,N_1219,N_2739);
xnor U4437 (N_4437,N_1550,N_3647);
nand U4438 (N_4438,N_3860,N_3573);
nor U4439 (N_4439,N_111,N_2461);
nand U4440 (N_4440,N_1136,N_1672);
and U4441 (N_4441,N_114,N_3484);
nor U4442 (N_4442,N_2772,N_1288);
and U4443 (N_4443,N_3571,N_2157);
xnor U4444 (N_4444,N_208,N_1586);
nand U4445 (N_4445,N_1037,N_1380);
xnor U4446 (N_4446,N_3816,N_775);
nor U4447 (N_4447,N_368,N_688);
xor U4448 (N_4448,N_74,N_1894);
nand U4449 (N_4449,N_1690,N_2284);
or U4450 (N_4450,N_2387,N_3597);
nor U4451 (N_4451,N_802,N_2421);
and U4452 (N_4452,N_968,N_3523);
or U4453 (N_4453,N_3964,N_50);
nor U4454 (N_4454,N_2130,N_2917);
nor U4455 (N_4455,N_2722,N_2204);
nand U4456 (N_4456,N_3877,N_696);
nor U4457 (N_4457,N_319,N_2527);
or U4458 (N_4458,N_707,N_1004);
nand U4459 (N_4459,N_653,N_2530);
nor U4460 (N_4460,N_697,N_77);
nand U4461 (N_4461,N_2414,N_575);
nand U4462 (N_4462,N_1344,N_2337);
or U4463 (N_4463,N_501,N_1234);
xnor U4464 (N_4464,N_767,N_1196);
or U4465 (N_4465,N_514,N_1984);
nor U4466 (N_4466,N_359,N_3165);
or U4467 (N_4467,N_3200,N_2953);
nor U4468 (N_4468,N_1419,N_1112);
nor U4469 (N_4469,N_3933,N_2148);
nor U4470 (N_4470,N_2797,N_2174);
nand U4471 (N_4471,N_599,N_1521);
nor U4472 (N_4472,N_1286,N_3147);
nand U4473 (N_4473,N_3118,N_1992);
and U4474 (N_4474,N_353,N_3766);
nand U4475 (N_4475,N_1578,N_2355);
nand U4476 (N_4476,N_1961,N_2480);
nor U4477 (N_4477,N_1151,N_590);
nand U4478 (N_4478,N_877,N_633);
nand U4479 (N_4479,N_1704,N_3429);
xor U4480 (N_4480,N_1966,N_2805);
and U4481 (N_4481,N_2344,N_415);
and U4482 (N_4482,N_3189,N_1921);
and U4483 (N_4483,N_3760,N_2993);
nand U4484 (N_4484,N_104,N_340);
and U4485 (N_4485,N_3360,N_2845);
nor U4486 (N_4486,N_2798,N_3611);
nor U4487 (N_4487,N_3817,N_785);
nor U4488 (N_4488,N_3101,N_1457);
nor U4489 (N_4489,N_2730,N_2517);
or U4490 (N_4490,N_2499,N_1523);
nand U4491 (N_4491,N_795,N_641);
and U4492 (N_4492,N_546,N_3962);
or U4493 (N_4493,N_98,N_534);
and U4494 (N_4494,N_15,N_2896);
or U4495 (N_4495,N_3500,N_2833);
nand U4496 (N_4496,N_175,N_568);
xor U4497 (N_4497,N_1786,N_1290);
xnor U4498 (N_4498,N_1070,N_1935);
or U4499 (N_4499,N_3579,N_1922);
and U4500 (N_4500,N_366,N_2985);
nand U4501 (N_4501,N_3241,N_2259);
nand U4502 (N_4502,N_605,N_2408);
nor U4503 (N_4503,N_853,N_3743);
nand U4504 (N_4504,N_2129,N_1010);
xnor U4505 (N_4505,N_1878,N_2604);
nand U4506 (N_4506,N_2639,N_2271);
nor U4507 (N_4507,N_1316,N_1111);
nand U4508 (N_4508,N_1411,N_1295);
or U4509 (N_4509,N_3552,N_2877);
and U4510 (N_4510,N_1229,N_3437);
and U4511 (N_4511,N_3022,N_24);
nor U4512 (N_4512,N_3799,N_1663);
and U4513 (N_4513,N_3275,N_3594);
and U4514 (N_4514,N_797,N_2094);
or U4515 (N_4515,N_3822,N_3031);
nor U4516 (N_4516,N_2609,N_1429);
nor U4517 (N_4517,N_3129,N_1840);
nor U4518 (N_4518,N_3,N_427);
or U4519 (N_4519,N_2788,N_405);
or U4520 (N_4520,N_3453,N_2968);
nand U4521 (N_4521,N_3830,N_312);
nand U4522 (N_4522,N_1826,N_2475);
nor U4523 (N_4523,N_1492,N_2230);
nor U4524 (N_4524,N_320,N_744);
xnor U4525 (N_4525,N_2770,N_2407);
xor U4526 (N_4526,N_3306,N_3869);
or U4527 (N_4527,N_2234,N_976);
or U4528 (N_4528,N_3056,N_446);
or U4529 (N_4529,N_2679,N_827);
xor U4530 (N_4530,N_245,N_1195);
nand U4531 (N_4531,N_889,N_2146);
or U4532 (N_4532,N_683,N_2983);
nor U4533 (N_4533,N_3852,N_1698);
nor U4534 (N_4534,N_482,N_717);
and U4535 (N_4535,N_563,N_1087);
nand U4536 (N_4536,N_1300,N_2661);
or U4537 (N_4537,N_2599,N_2470);
and U4538 (N_4538,N_3991,N_608);
nand U4539 (N_4539,N_3928,N_2830);
nor U4540 (N_4540,N_2775,N_2203);
or U4541 (N_4541,N_3135,N_2708);
or U4542 (N_4542,N_3154,N_3134);
and U4543 (N_4543,N_3314,N_1747);
and U4544 (N_4544,N_1744,N_2110);
or U4545 (N_4545,N_3979,N_1702);
nand U4546 (N_4546,N_2568,N_3221);
nor U4547 (N_4547,N_3763,N_2655);
or U4548 (N_4548,N_1539,N_301);
or U4549 (N_4549,N_1555,N_579);
nor U4550 (N_4550,N_1846,N_127);
nand U4551 (N_4551,N_1573,N_3851);
and U4552 (N_4552,N_3716,N_1977);
nand U4553 (N_4553,N_2618,N_2844);
or U4554 (N_4554,N_1437,N_2494);
or U4555 (N_4555,N_1335,N_3692);
xor U4556 (N_4556,N_2250,N_1488);
xnor U4557 (N_4557,N_3929,N_3132);
nand U4558 (N_4558,N_2159,N_2633);
and U4559 (N_4559,N_3883,N_910);
or U4560 (N_4560,N_1221,N_1902);
and U4561 (N_4561,N_958,N_1305);
nor U4562 (N_4562,N_2177,N_3539);
nand U4563 (N_4563,N_1047,N_3617);
xor U4564 (N_4564,N_1797,N_2272);
and U4565 (N_4565,N_3020,N_1403);
nand U4566 (N_4566,N_1129,N_880);
and U4567 (N_4567,N_3009,N_883);
xor U4568 (N_4568,N_3704,N_107);
and U4569 (N_4569,N_3461,N_3682);
nand U4570 (N_4570,N_945,N_2782);
or U4571 (N_4571,N_1647,N_1250);
nor U4572 (N_4572,N_271,N_2163);
and U4573 (N_4573,N_1222,N_1621);
or U4574 (N_4574,N_657,N_2575);
nor U4575 (N_4575,N_1023,N_300);
xor U4576 (N_4576,N_834,N_2826);
xor U4577 (N_4577,N_3904,N_1125);
or U4578 (N_4578,N_1043,N_317);
and U4579 (N_4579,N_835,N_1245);
xor U4580 (N_4580,N_264,N_3921);
nor U4581 (N_4581,N_3304,N_566);
nand U4582 (N_4582,N_3474,N_2229);
or U4583 (N_4583,N_447,N_558);
or U4584 (N_4584,N_2902,N_1292);
or U4585 (N_4585,N_3321,N_2237);
nand U4586 (N_4586,N_3728,N_1267);
and U4587 (N_4587,N_3741,N_953);
or U4588 (N_4588,N_2944,N_1285);
or U4589 (N_4589,N_2413,N_3455);
nand U4590 (N_4590,N_3264,N_2120);
nand U4591 (N_4591,N_134,N_3338);
nor U4592 (N_4592,N_648,N_3758);
and U4593 (N_4593,N_34,N_2957);
xor U4594 (N_4594,N_3106,N_100);
and U4595 (N_4595,N_3234,N_1249);
or U4596 (N_4596,N_1182,N_3291);
or U4597 (N_4597,N_1359,N_2245);
nor U4598 (N_4598,N_916,N_1066);
xnor U4599 (N_4599,N_1008,N_275);
and U4600 (N_4600,N_3835,N_1721);
and U4601 (N_4601,N_2140,N_3286);
xnor U4602 (N_4602,N_1120,N_2370);
xnor U4603 (N_4603,N_1065,N_2081);
and U4604 (N_4604,N_1371,N_3250);
and U4605 (N_4605,N_2815,N_2874);
or U4606 (N_4606,N_2038,N_1183);
and U4607 (N_4607,N_192,N_2253);
nand U4608 (N_4608,N_2251,N_1805);
nor U4609 (N_4609,N_1477,N_303);
and U4610 (N_4610,N_3292,N_3703);
or U4611 (N_4611,N_3551,N_2238);
nand U4612 (N_4612,N_3356,N_1475);
and U4613 (N_4613,N_1981,N_2426);
nor U4614 (N_4614,N_3424,N_1198);
and U4615 (N_4615,N_3881,N_3319);
or U4616 (N_4616,N_1283,N_1963);
or U4617 (N_4617,N_864,N_43);
nor U4618 (N_4618,N_133,N_1060);
nor U4619 (N_4619,N_1106,N_850);
nor U4620 (N_4620,N_1815,N_1881);
xnor U4621 (N_4621,N_3664,N_44);
nor U4622 (N_4622,N_3035,N_907);
or U4623 (N_4623,N_3344,N_1449);
nand U4624 (N_4624,N_3945,N_3960);
or U4625 (N_4625,N_2342,N_2015);
nor U4626 (N_4626,N_3104,N_3206);
nand U4627 (N_4627,N_1589,N_3764);
or U4628 (N_4628,N_746,N_705);
nor U4629 (N_4629,N_89,N_844);
nor U4630 (N_4630,N_1406,N_3021);
nand U4631 (N_4631,N_3421,N_2553);
or U4632 (N_4632,N_2854,N_1970);
or U4633 (N_4633,N_894,N_163);
and U4634 (N_4634,N_3638,N_206);
or U4635 (N_4635,N_2940,N_2383);
and U4636 (N_4636,N_3235,N_815);
nand U4637 (N_4637,N_1399,N_1593);
nor U4638 (N_4638,N_1405,N_81);
or U4639 (N_4639,N_2549,N_1202);
nor U4640 (N_4640,N_3707,N_3072);
or U4641 (N_4641,N_1083,N_3913);
and U4642 (N_4642,N_1934,N_862);
nand U4643 (N_4643,N_2012,N_3562);
nor U4644 (N_4644,N_919,N_3995);
nand U4645 (N_4645,N_1417,N_2736);
nand U4646 (N_4646,N_2884,N_103);
and U4647 (N_4647,N_1232,N_509);
or U4648 (N_4648,N_1224,N_1001);
nand U4649 (N_4649,N_3511,N_2044);
and U4650 (N_4650,N_2933,N_2137);
nand U4651 (N_4651,N_2753,N_908);
and U4652 (N_4652,N_663,N_3582);
nand U4653 (N_4653,N_2995,N_2999);
nor U4654 (N_4654,N_2531,N_750);
nor U4655 (N_4655,N_3740,N_3971);
nand U4656 (N_4656,N_3448,N_2976);
nor U4657 (N_4657,N_440,N_1287);
nor U4658 (N_4658,N_3859,N_376);
nand U4659 (N_4659,N_831,N_3892);
or U4660 (N_4660,N_2386,N_2176);
nand U4661 (N_4661,N_182,N_1763);
nor U4662 (N_4662,N_2079,N_1714);
or U4663 (N_4663,N_1472,N_1748);
nor U4664 (N_4664,N_305,N_1743);
or U4665 (N_4665,N_2196,N_2754);
and U4666 (N_4666,N_1904,N_1520);
nor U4667 (N_4667,N_1909,N_2331);
nor U4668 (N_4668,N_3033,N_3600);
and U4669 (N_4669,N_3686,N_1203);
nor U4670 (N_4670,N_2812,N_2851);
or U4671 (N_4671,N_2380,N_959);
nor U4672 (N_4672,N_1051,N_3058);
nor U4673 (N_4673,N_1434,N_2317);
or U4674 (N_4674,N_3542,N_1121);
or U4675 (N_4675,N_2131,N_1452);
or U4676 (N_4676,N_863,N_2346);
and U4677 (N_4677,N_2033,N_1675);
or U4678 (N_4678,N_2243,N_3032);
xnor U4679 (N_4679,N_1564,N_31);
xnor U4680 (N_4680,N_1190,N_1017);
nand U4681 (N_4681,N_3379,N_3524);
nand U4682 (N_4682,N_1700,N_3145);
and U4683 (N_4683,N_2818,N_3992);
or U4684 (N_4684,N_2153,N_2787);
and U4685 (N_4685,N_1501,N_990);
nand U4686 (N_4686,N_3808,N_2018);
or U4687 (N_4687,N_1013,N_3352);
and U4688 (N_4688,N_800,N_2610);
and U4689 (N_4689,N_3067,N_1150);
and U4690 (N_4690,N_939,N_1446);
or U4691 (N_4691,N_3412,N_2513);
nand U4692 (N_4692,N_249,N_3847);
and U4693 (N_4693,N_586,N_3185);
nor U4694 (N_4694,N_1256,N_1042);
xnor U4695 (N_4695,N_704,N_887);
xnor U4696 (N_4696,N_3644,N_1427);
and U4697 (N_4697,N_2090,N_318);
and U4698 (N_4698,N_3897,N_3452);
xnor U4699 (N_4699,N_1711,N_2285);
nand U4700 (N_4700,N_3864,N_3233);
nand U4701 (N_4701,N_1078,N_1979);
nor U4702 (N_4702,N_1960,N_1775);
nor U4703 (N_4703,N_185,N_2577);
and U4704 (N_4704,N_1170,N_792);
nor U4705 (N_4705,N_1275,N_790);
xnor U4706 (N_4706,N_3658,N_3717);
xnor U4707 (N_4707,N_2444,N_66);
and U4708 (N_4708,N_2318,N_3823);
or U4709 (N_4709,N_596,N_2520);
or U4710 (N_4710,N_3888,N_634);
nand U4711 (N_4711,N_735,N_3657);
or U4712 (N_4712,N_3383,N_80);
nand U4713 (N_4713,N_3471,N_1616);
nand U4714 (N_4714,N_1029,N_463);
nor U4715 (N_4715,N_1095,N_2970);
and U4716 (N_4716,N_1827,N_345);
or U4717 (N_4717,N_1530,N_1240);
nand U4718 (N_4718,N_3549,N_1298);
xnor U4719 (N_4719,N_724,N_829);
xnor U4720 (N_4720,N_3077,N_2195);
nor U4721 (N_4721,N_1823,N_2356);
and U4722 (N_4722,N_2014,N_1068);
and U4723 (N_4723,N_2964,N_1389);
or U4724 (N_4724,N_1347,N_3797);
and U4725 (N_4725,N_2866,N_824);
and U4726 (N_4726,N_2689,N_2458);
nor U4727 (N_4727,N_2562,N_3257);
xnor U4728 (N_4728,N_1740,N_1093);
nor U4729 (N_4729,N_2297,N_1798);
and U4730 (N_4730,N_1557,N_2027);
nand U4731 (N_4731,N_3409,N_386);
and U4732 (N_4732,N_2791,N_39);
nor U4733 (N_4733,N_1959,N_3912);
nor U4734 (N_4734,N_3433,N_3362);
nor U4735 (N_4735,N_1756,N_3974);
nand U4736 (N_4736,N_1079,N_3935);
or U4737 (N_4737,N_3509,N_3622);
or U4738 (N_4738,N_494,N_3166);
and U4739 (N_4739,N_230,N_2910);
nor U4740 (N_4740,N_807,N_1949);
nand U4741 (N_4741,N_3874,N_1345);
or U4742 (N_4742,N_2202,N_1467);
or U4743 (N_4743,N_1333,N_698);
or U4744 (N_4744,N_3188,N_1974);
xor U4745 (N_4745,N_61,N_3807);
xor U4746 (N_4746,N_223,N_3953);
nand U4747 (N_4747,N_1480,N_1096);
nand U4748 (N_4748,N_868,N_3393);
and U4749 (N_4749,N_2662,N_3496);
nand U4750 (N_4750,N_2743,N_2312);
xnor U4751 (N_4751,N_146,N_1435);
or U4752 (N_4752,N_3633,N_162);
xnor U4753 (N_4753,N_3149,N_3287);
nand U4754 (N_4754,N_382,N_583);
or U4755 (N_4755,N_920,N_1107);
nand U4756 (N_4756,N_1025,N_2975);
nor U4757 (N_4757,N_2165,N_2029);
nor U4758 (N_4758,N_3793,N_542);
nand U4759 (N_4759,N_3194,N_884);
or U4760 (N_4760,N_1622,N_26);
and U4761 (N_4761,N_391,N_629);
nor U4762 (N_4762,N_3243,N_130);
nor U4763 (N_4763,N_513,N_3080);
xor U4764 (N_4764,N_2021,N_2095);
nand U4765 (N_4765,N_1695,N_1007);
and U4766 (N_4766,N_2124,N_1542);
xor U4767 (N_4767,N_2808,N_3091);
nor U4768 (N_4768,N_1363,N_2635);
xor U4769 (N_4769,N_743,N_147);
xnor U4770 (N_4770,N_1637,N_10);
nor U4771 (N_4771,N_492,N_156);
nand U4772 (N_4772,N_1936,N_1807);
or U4773 (N_4773,N_3849,N_2210);
and U4774 (N_4774,N_252,N_2982);
nand U4775 (N_4775,N_2758,N_932);
nand U4776 (N_4776,N_1820,N_1444);
and U4777 (N_4777,N_1546,N_3044);
or U4778 (N_4778,N_3231,N_3207);
nor U4779 (N_4779,N_1832,N_2657);
nand U4780 (N_4780,N_3762,N_3370);
or U4781 (N_4781,N_2555,N_3898);
or U4782 (N_4782,N_2339,N_708);
nand U4783 (N_4783,N_304,N_3761);
or U4784 (N_4784,N_2761,N_3164);
or U4785 (N_4785,N_1975,N_2483);
or U4786 (N_4786,N_2416,N_2405);
nand U4787 (N_4787,N_3015,N_334);
nor U4788 (N_4788,N_3920,N_2928);
xnor U4789 (N_4789,N_3540,N_2856);
nor U4790 (N_4790,N_241,N_609);
nand U4791 (N_4791,N_2492,N_944);
nor U4792 (N_4792,N_3606,N_2634);
nor U4793 (N_4793,N_3809,N_131);
nor U4794 (N_4794,N_1677,N_69);
and U4795 (N_4795,N_1882,N_1678);
xnor U4796 (N_4796,N_1685,N_3846);
nor U4797 (N_4797,N_1328,N_3008);
and U4798 (N_4798,N_218,N_3583);
nor U4799 (N_4799,N_772,N_1770);
nand U4800 (N_4800,N_2074,N_68);
nand U4801 (N_4801,N_161,N_3959);
and U4802 (N_4802,N_1152,N_233);
and U4803 (N_4803,N_2590,N_2085);
nand U4804 (N_4804,N_7,N_1682);
or U4805 (N_4805,N_1782,N_1965);
nand U4806 (N_4806,N_1303,N_2543);
and U4807 (N_4807,N_2072,N_2873);
nand U4808 (N_4808,N_1600,N_503);
or U4809 (N_4809,N_126,N_1839);
nor U4810 (N_4810,N_3066,N_330);
or U4811 (N_4811,N_2836,N_1193);
or U4812 (N_4812,N_1617,N_2705);
or U4813 (N_4813,N_1145,N_3715);
and U4814 (N_4814,N_1772,N_1274);
xnor U4815 (N_4815,N_2850,N_1200);
nand U4816 (N_4816,N_1646,N_2883);
and U4817 (N_4817,N_3720,N_1409);
nand U4818 (N_4818,N_3153,N_1990);
nand U4819 (N_4819,N_3896,N_2255);
nor U4820 (N_4820,N_1097,N_3251);
nand U4821 (N_4821,N_3609,N_1718);
nand U4822 (N_4822,N_782,N_3222);
nor U4823 (N_4823,N_2228,N_2516);
or U4824 (N_4824,N_3001,N_995);
nor U4825 (N_4825,N_2112,N_882);
nand U4826 (N_4826,N_14,N_3441);
xnor U4827 (N_4827,N_3842,N_2462);
and U4828 (N_4828,N_1413,N_2127);
nor U4829 (N_4829,N_2422,N_3932);
or U4830 (N_4830,N_3312,N_489);
nor U4831 (N_4831,N_2632,N_2544);
xor U4832 (N_4832,N_37,N_1536);
or U4833 (N_4833,N_3016,N_631);
nand U4834 (N_4834,N_828,N_2000);
nand U4835 (N_4835,N_3527,N_1493);
nand U4836 (N_4836,N_3709,N_2450);
or U4837 (N_4837,N_1893,N_1370);
nand U4838 (N_4838,N_553,N_1741);
or U4839 (N_4839,N_184,N_3258);
nand U4840 (N_4840,N_1062,N_1845);
and U4841 (N_4841,N_2665,N_1374);
nor U4842 (N_4842,N_484,N_2558);
nand U4843 (N_4843,N_3394,N_1294);
or U4844 (N_4844,N_1130,N_1890);
xnor U4845 (N_4845,N_3538,N_3369);
nand U4846 (N_4846,N_404,N_2065);
nand U4847 (N_4847,N_2861,N_3980);
or U4848 (N_4848,N_438,N_2840);
nand U4849 (N_4849,N_3501,N_181);
or U4850 (N_4850,N_3927,N_1465);
and U4851 (N_4851,N_1251,N_1209);
nor U4852 (N_4852,N_200,N_1507);
or U4853 (N_4853,N_115,N_861);
and U4854 (N_4854,N_189,N_2365);
xnor U4855 (N_4855,N_1433,N_2872);
nor U4856 (N_4856,N_2515,N_982);
nand U4857 (N_4857,N_1541,N_2327);
or U4858 (N_4858,N_3151,N_3614);
and U4859 (N_4859,N_3900,N_36);
and U4860 (N_4860,N_3419,N_1378);
nand U4861 (N_4861,N_3584,N_1373);
nor U4862 (N_4862,N_3120,N_2688);
or U4863 (N_4863,N_680,N_302);
or U4864 (N_4864,N_3748,N_1441);
or U4865 (N_4865,N_2699,N_517);
and U4866 (N_4866,N_2,N_1973);
nand U4867 (N_4867,N_3976,N_2541);
nor U4868 (N_4868,N_1785,N_1261);
and U4869 (N_4869,N_1819,N_3176);
or U4870 (N_4870,N_3366,N_400);
nor U4871 (N_4871,N_2454,N_1674);
nor U4872 (N_4872,N_2180,N_1944);
xnor U4873 (N_4873,N_1279,N_1559);
and U4874 (N_4874,N_3669,N_1766);
nor U4875 (N_4875,N_2254,N_1676);
nand U4876 (N_4876,N_591,N_2786);
xnor U4877 (N_4877,N_58,N_1284);
xnor U4878 (N_4878,N_3733,N_3005);
nor U4879 (N_4879,N_3495,N_1816);
and U4880 (N_4880,N_2198,N_437);
or U4881 (N_4881,N_2651,N_1431);
and U4882 (N_4882,N_2747,N_3037);
nor U4883 (N_4883,N_3302,N_2410);
nor U4884 (N_4884,N_1168,N_220);
or U4885 (N_4885,N_3677,N_2400);
xnor U4886 (N_4886,N_3784,N_120);
nor U4887 (N_4887,N_2367,N_3681);
nor U4888 (N_4888,N_3087,N_343);
or U4889 (N_4889,N_485,N_967);
or U4890 (N_4890,N_2053,N_2537);
or U4891 (N_4891,N_2839,N_2169);
xnor U4892 (N_4892,N_615,N_3161);
or U4893 (N_4893,N_3192,N_3142);
nand U4894 (N_4894,N_2625,N_1503);
xnor U4895 (N_4895,N_3322,N_3464);
and U4896 (N_4896,N_973,N_3486);
nand U4897 (N_4897,N_459,N_2519);
and U4898 (N_4898,N_3432,N_2403);
and U4899 (N_4899,N_2338,N_666);
nor U4900 (N_4900,N_3029,N_2930);
and U4901 (N_4901,N_1059,N_1327);
xor U4902 (N_4902,N_984,N_2592);
or U4903 (N_4903,N_1849,N_3367);
and U4904 (N_4904,N_2997,N_430);
and U4905 (N_4905,N_664,N_540);
nand U4906 (N_4906,N_2630,N_2145);
nor U4907 (N_4907,N_259,N_112);
or U4908 (N_4908,N_3390,N_2201);
xnor U4909 (N_4909,N_361,N_1308);
and U4910 (N_4910,N_3544,N_2734);
or U4911 (N_4911,N_617,N_1692);
or U4912 (N_4912,N_3515,N_1159);
and U4913 (N_4913,N_3480,N_3785);
nand U4914 (N_4914,N_2498,N_1610);
nor U4915 (N_4915,N_495,N_510);
nor U4916 (N_4916,N_423,N_3676);
xnor U4917 (N_4917,N_395,N_2653);
or U4918 (N_4918,N_3783,N_3069);
or U4919 (N_4919,N_3901,N_1115);
and U4920 (N_4920,N_3800,N_3742);
or U4921 (N_4921,N_849,N_646);
nand U4922 (N_4922,N_879,N_1489);
nand U4923 (N_4923,N_128,N_3476);
nand U4924 (N_4924,N_3485,N_326);
and U4925 (N_4925,N_3934,N_2820);
or U4926 (N_4926,N_1760,N_1806);
nand U4927 (N_4927,N_356,N_3805);
xor U4928 (N_4928,N_2314,N_1511);
xor U4929 (N_4929,N_1897,N_2681);
and U4930 (N_4930,N_3554,N_2304);
nand U4931 (N_4931,N_346,N_3649);
and U4932 (N_4932,N_3174,N_593);
nor U4933 (N_4933,N_1077,N_3873);
nand U4934 (N_4934,N_1045,N_3632);
nor U4935 (N_4935,N_3942,N_38);
and U4936 (N_4936,N_2035,N_2114);
xnor U4937 (N_4937,N_235,N_1257);
xnor U4938 (N_4938,N_3621,N_2019);
or U4939 (N_4939,N_2020,N_290);
nand U4940 (N_4940,N_3675,N_3702);
or U4941 (N_4941,N_1828,N_2946);
nor U4942 (N_4942,N_2627,N_1205);
nand U4943 (N_4943,N_3699,N_3984);
and U4944 (N_4944,N_3026,N_1529);
and U4945 (N_4945,N_3725,N_1099);
and U4946 (N_4946,N_2551,N_277);
and U4947 (N_4947,N_1213,N_357);
nand U4948 (N_4948,N_1933,N_418);
and U4949 (N_4949,N_3368,N_947);
or U4950 (N_4950,N_3042,N_1015);
nor U4951 (N_4951,N_1615,N_1197);
and U4952 (N_4952,N_1277,N_2643);
nor U4953 (N_4953,N_3481,N_3968);
nand U4954 (N_4954,N_1311,N_1058);
or U4955 (N_4955,N_3112,N_3329);
nor U4956 (N_4956,N_1038,N_3525);
nor U4957 (N_4957,N_2719,N_203);
nand U4958 (N_4958,N_2649,N_964);
xnor U4959 (N_4959,N_1343,N_1206);
nor U4960 (N_4960,N_2955,N_1149);
and U4961 (N_4961,N_3711,N_3420);
nor U4962 (N_4962,N_384,N_2676);
and U4963 (N_4963,N_2291,N_3770);
and U4964 (N_4964,N_727,N_1153);
nand U4965 (N_4965,N_2336,N_2581);
nand U4966 (N_4966,N_2103,N_1422);
nor U4967 (N_4967,N_2034,N_469);
nor U4968 (N_4968,N_922,N_449);
xnor U4969 (N_4969,N_3825,N_1098);
nand U4970 (N_4970,N_3914,N_1727);
or U4971 (N_4971,N_2504,N_2411);
or U4972 (N_4972,N_3353,N_1848);
and U4973 (N_4973,N_270,N_2925);
nand U4974 (N_4974,N_651,N_1898);
and U4975 (N_4975,N_2546,N_3408);
nand U4976 (N_4976,N_11,N_999);
and U4977 (N_4977,N_3271,N_1950);
nand U4978 (N_4978,N_2589,N_1779);
nor U4979 (N_4979,N_1582,N_581);
nor U4980 (N_4980,N_3556,N_2278);
and U4981 (N_4981,N_2766,N_2472);
nor U4982 (N_4982,N_3803,N_2463);
nand U4983 (N_4983,N_2374,N_3753);
and U4984 (N_4984,N_2838,N_2831);
and U4985 (N_4985,N_16,N_1724);
and U4986 (N_4986,N_3248,N_621);
and U4987 (N_4987,N_2685,N_557);
nor U4988 (N_4988,N_2002,N_2036);
or U4989 (N_4989,N_1746,N_388);
nor U4990 (N_4990,N_1924,N_3684);
or U4991 (N_4991,N_897,N_3220);
or U4992 (N_4992,N_314,N_3285);
nor U4993 (N_4993,N_3790,N_3909);
xnor U4994 (N_4994,N_1341,N_1525);
or U4995 (N_4995,N_207,N_1470);
and U4996 (N_4996,N_1122,N_1916);
nor U4997 (N_4997,N_3012,N_1712);
nand U4998 (N_4998,N_2506,N_1914);
nor U4999 (N_4999,N_426,N_846);
and U5000 (N_5000,N_1597,N_1494);
or U5001 (N_5001,N_2098,N_679);
and U5002 (N_5002,N_2888,N_3879);
xnor U5003 (N_5003,N_1540,N_1595);
nor U5004 (N_5004,N_2769,N_2732);
nor U5005 (N_5005,N_2184,N_3443);
xor U5006 (N_5006,N_1299,N_2629);
and U5007 (N_5007,N_3530,N_1318);
nor U5008 (N_5008,N_2919,N_3459);
nand U5009 (N_5009,N_3727,N_471);
nand U5010 (N_5010,N_281,N_1585);
nor U5011 (N_5011,N_3462,N_751);
or U5012 (N_5012,N_3957,N_2756);
or U5013 (N_5013,N_2007,N_777);
nand U5014 (N_5014,N_1817,N_3516);
nand U5015 (N_5015,N_805,N_3956);
and U5016 (N_5016,N_722,N_3973);
and U5017 (N_5017,N_2726,N_3371);
xor U5018 (N_5018,N_3049,N_71);
or U5019 (N_5019,N_3046,N_522);
or U5020 (N_5020,N_2929,N_3841);
or U5021 (N_5021,N_3671,N_1443);
xnor U5022 (N_5022,N_2740,N_3086);
or U5023 (N_5023,N_2102,N_3819);
nor U5024 (N_5024,N_2825,N_781);
nand U5025 (N_5025,N_3533,N_3010);
nand U5026 (N_5026,N_748,N_2733);
and U5027 (N_5027,N_1230,N_421);
or U5028 (N_5028,N_1515,N_2759);
and U5029 (N_5029,N_2564,N_840);
and U5030 (N_5030,N_3757,N_2650);
nor U5031 (N_5031,N_3479,N_3346);
xor U5032 (N_5032,N_1020,N_1688);
nor U5033 (N_5033,N_154,N_588);
or U5034 (N_5034,N_2731,N_1653);
and U5035 (N_5035,N_2152,N_443);
nand U5036 (N_5036,N_1268,N_2466);
nand U5037 (N_5037,N_1664,N_3378);
and U5038 (N_5038,N_488,N_560);
nand U5039 (N_5039,N_2617,N_1500);
and U5040 (N_5040,N_3027,N_3303);
nand U5041 (N_5041,N_3193,N_756);
nand U5042 (N_5042,N_226,N_3936);
xnor U5043 (N_5043,N_1119,N_1360);
nand U5044 (N_5044,N_2092,N_3585);
nor U5045 (N_5045,N_188,N_3771);
or U5046 (N_5046,N_3966,N_2136);
or U5047 (N_5047,N_3245,N_436);
nor U5048 (N_5048,N_3648,N_2842);
nor U5049 (N_5049,N_766,N_3836);
nand U5050 (N_5050,N_2947,N_2691);
nand U5051 (N_5051,N_3034,N_3670);
and U5052 (N_5052,N_1379,N_3713);
or U5053 (N_5053,N_3229,N_204);
nand U5054 (N_5054,N_1920,N_1306);
xnor U5055 (N_5055,N_2452,N_3382);
and U5056 (N_5056,N_3653,N_628);
xor U5057 (N_5057,N_3737,N_3028);
and U5058 (N_5058,N_180,N_2050);
or U5059 (N_5059,N_402,N_451);
or U5060 (N_5060,N_1178,N_3198);
or U5061 (N_5061,N_2322,N_2193);
nor U5062 (N_5062,N_1400,N_1297);
nor U5063 (N_5063,N_2636,N_2567);
or U5064 (N_5064,N_3004,N_983);
or U5065 (N_5065,N_1366,N_2721);
nor U5066 (N_5066,N_9,N_938);
and U5067 (N_5067,N_2809,N_2916);
or U5068 (N_5068,N_1324,N_1340);
nor U5069 (N_5069,N_416,N_160);
and U5070 (N_5070,N_567,N_2795);
nor U5071 (N_5071,N_3320,N_1016);
and U5072 (N_5072,N_2308,N_1997);
or U5073 (N_5073,N_793,N_859);
and U5074 (N_5074,N_3543,N_1607);
xnor U5075 (N_5075,N_1046,N_1063);
xnor U5076 (N_5076,N_550,N_2427);
xnor U5077 (N_5077,N_3327,N_865);
or U5078 (N_5078,N_3867,N_1735);
nor U5079 (N_5079,N_1228,N_1425);
and U5080 (N_5080,N_961,N_2745);
nand U5081 (N_5081,N_2257,N_3963);
nor U5082 (N_5082,N_2315,N_3581);
or U5083 (N_5083,N_2943,N_1650);
and U5084 (N_5084,N_1210,N_2959);
nor U5085 (N_5085,N_1282,N_3375);
nand U5086 (N_5086,N_2951,N_2556);
xor U5087 (N_5087,N_2442,N_2260);
or U5088 (N_5088,N_3191,N_2560);
or U5089 (N_5089,N_1783,N_1238);
nor U5090 (N_5090,N_505,N_569);
and U5091 (N_5091,N_809,N_3082);
nor U5092 (N_5092,N_149,N_731);
and U5093 (N_5093,N_2806,N_193);
or U5094 (N_5094,N_2792,N_725);
nor U5095 (N_5095,N_3247,N_57);
or U5096 (N_5096,N_2880,N_117);
nor U5097 (N_5097,N_1537,N_2654);
nor U5098 (N_5098,N_2871,N_2425);
and U5099 (N_5099,N_783,N_3998);
nor U5100 (N_5100,N_231,N_3418);
or U5101 (N_5101,N_1781,N_1885);
or U5102 (N_5102,N_2757,N_576);
and U5103 (N_5103,N_2684,N_2070);
nor U5104 (N_5104,N_927,N_1);
or U5105 (N_5105,N_1315,N_3483);
or U5106 (N_5106,N_1109,N_2926);
and U5107 (N_5107,N_3700,N_265);
or U5108 (N_5108,N_3339,N_3599);
nand U5109 (N_5109,N_1448,N_234);
and U5110 (N_5110,N_344,N_1590);
nand U5111 (N_5111,N_1945,N_773);
nand U5112 (N_5112,N_435,N_3236);
nor U5113 (N_5113,N_960,N_1618);
nor U5114 (N_5114,N_2041,N_1792);
nand U5115 (N_5115,N_3712,N_2051);
xnor U5116 (N_5116,N_825,N_172);
nand U5117 (N_5117,N_732,N_3078);
and U5118 (N_5118,N_2389,N_3117);
nor U5119 (N_5119,N_1771,N_3981);
nor U5120 (N_5120,N_2765,N_1773);
nand U5121 (N_5121,N_1883,N_3514);
nor U5122 (N_5122,N_3223,N_2139);
or U5123 (N_5123,N_1160,N_1259);
nor U5124 (N_5124,N_3279,N_3326);
or U5125 (N_5125,N_2897,N_502);
or U5126 (N_5126,N_12,N_2742);
nor U5127 (N_5127,N_1101,N_213);
nand U5128 (N_5128,N_1645,N_3810);
nor U5129 (N_5129,N_1460,N_1158);
or U5130 (N_5130,N_3613,N_1728);
nand U5131 (N_5131,N_3578,N_1040);
nand U5132 (N_5132,N_518,N_998);
and U5133 (N_5133,N_1793,N_626);
and U5134 (N_5134,N_183,N_452);
or U5135 (N_5135,N_1968,N_2891);
nand U5136 (N_5136,N_3635,N_623);
or U5137 (N_5137,N_2300,N_434);
nor U5138 (N_5138,N_1640,N_1887);
and U5139 (N_5139,N_2329,N_2009);
xor U5140 (N_5140,N_2542,N_3201);
nor U5141 (N_5141,N_335,N_143);
nand U5142 (N_5142,N_221,N_138);
nor U5143 (N_5143,N_694,N_2518);
or U5144 (N_5144,N_3946,N_3038);
nand U5145 (N_5145,N_537,N_3434);
nor U5146 (N_5146,N_3858,N_2448);
or U5147 (N_5147,N_539,N_649);
and U5148 (N_5148,N_3468,N_3801);
or U5149 (N_5149,N_3576,N_1745);
nand U5150 (N_5150,N_3175,N_394);
or U5151 (N_5151,N_3497,N_3944);
and U5152 (N_5152,N_92,N_2593);
and U5153 (N_5153,N_803,N_1084);
nand U5154 (N_5154,N_3546,N_1499);
and U5155 (N_5155,N_1469,N_3893);
nor U5156 (N_5156,N_1867,N_3197);
and U5157 (N_5157,N_1978,N_1247);
xnor U5158 (N_5158,N_500,N_2611);
nor U5159 (N_5159,N_2583,N_660);
nor U5160 (N_5160,N_1587,N_3467);
nand U5161 (N_5161,N_177,N_1408);
nor U5162 (N_5162,N_2923,N_1377);
and U5163 (N_5163,N_3400,N_2172);
nand U5164 (N_5164,N_2749,N_1220);
xnor U5165 (N_5165,N_1208,N_261);
xnor U5166 (N_5166,N_1357,N_3487);
or U5167 (N_5167,N_2482,N_1012);
nand U5168 (N_5168,N_914,N_2040);
and U5169 (N_5169,N_3397,N_3526);
and U5170 (N_5170,N_2606,N_327);
nor U5171 (N_5171,N_2981,N_460);
nand U5172 (N_5172,N_2887,N_2432);
nand U5173 (N_5173,N_3139,N_2538);
and U5174 (N_5174,N_82,N_3666);
xnor U5175 (N_5175,N_3253,N_1648);
xnor U5176 (N_5176,N_1054,N_1192);
or U5177 (N_5177,N_3624,N_3156);
and U5178 (N_5178,N_1082,N_1421);
nor U5179 (N_5179,N_2240,N_2460);
nor U5180 (N_5180,N_1143,N_1495);
and U5181 (N_5181,N_572,N_2280);
nor U5182 (N_5182,N_2465,N_3000);
and U5183 (N_5183,N_822,N_1387);
xor U5184 (N_5184,N_3623,N_768);
and U5185 (N_5185,N_2415,N_483);
nor U5186 (N_5186,N_470,N_2269);
xnor U5187 (N_5187,N_1631,N_3121);
nor U5188 (N_5188,N_1307,N_2185);
nand U5189 (N_5189,N_18,N_3654);
nor U5190 (N_5190,N_3399,N_3045);
nand U5191 (N_5191,N_2804,N_1666);
xnor U5192 (N_5192,N_624,N_3734);
and U5193 (N_5193,N_3092,N_3404);
nor U5194 (N_5194,N_3767,N_1346);
or U5195 (N_5195,N_1233,N_3561);
nand U5196 (N_5196,N_3332,N_2714);
nor U5197 (N_5197,N_1076,N_2908);
nand U5198 (N_5198,N_2376,N_333);
or U5199 (N_5199,N_2055,N_2435);
or U5200 (N_5200,N_3096,N_291);
and U5201 (N_5201,N_3213,N_2076);
xor U5202 (N_5202,N_611,N_1895);
or U5203 (N_5203,N_1683,N_668);
and U5204 (N_5204,N_3199,N_2603);
or U5205 (N_5205,N_2449,N_179);
nor U5206 (N_5206,N_3482,N_1006);
nor U5207 (N_5207,N_1654,N_1394);
nor U5208 (N_5208,N_659,N_2173);
or U5209 (N_5209,N_952,N_2717);
nand U5210 (N_5210,N_1351,N_1094);
nand U5211 (N_5211,N_2728,N_2487);
or U5212 (N_5212,N_3260,N_1829);
nand U5213 (N_5213,N_2680,N_1179);
or U5214 (N_5214,N_2439,N_2889);
nand U5215 (N_5215,N_900,N_3708);
or U5216 (N_5216,N_1362,N_3567);
nand U5217 (N_5217,N_1720,N_497);
or U5218 (N_5218,N_2224,N_2552);
nor U5219 (N_5219,N_1693,N_1568);
nand U5220 (N_5220,N_1837,N_571);
nand U5221 (N_5221,N_1382,N_2780);
and U5222 (N_5222,N_1670,N_3181);
nand U5223 (N_5223,N_2652,N_1056);
and U5224 (N_5224,N_1795,N_1943);
and U5225 (N_5225,N_987,N_872);
nand U5226 (N_5226,N_166,N_60);
xnor U5227 (N_5227,N_3081,N_94);
or U5228 (N_5228,N_2794,N_3833);
xor U5229 (N_5229,N_295,N_1750);
and U5230 (N_5230,N_1641,N_1553);
or U5231 (N_5231,N_2430,N_1432);
and U5232 (N_5232,N_2324,N_2330);
or U5233 (N_5233,N_2996,N_2006);
nand U5234 (N_5234,N_2569,N_3065);
nand U5235 (N_5235,N_3428,N_2161);
nand U5236 (N_5236,N_852,N_2351);
nor U5237 (N_5237,N_1613,N_1314);
xor U5238 (N_5238,N_2417,N_3636);
nand U5239 (N_5239,N_3631,N_2334);
xnor U5240 (N_5240,N_499,N_905);
or U5241 (N_5241,N_132,N_3204);
nor U5242 (N_5242,N_1998,N_2967);
nand U5243 (N_5243,N_2835,N_896);
or U5244 (N_5244,N_2574,N_1466);
xnor U5245 (N_5245,N_925,N_268);
and U5246 (N_5246,N_54,N_1132);
or U5247 (N_5247,N_2441,N_898);
and U5248 (N_5248,N_3099,N_2613);
nor U5249 (N_5249,N_1439,N_512);
xor U5250 (N_5250,N_329,N_3060);
or U5251 (N_5251,N_1716,N_425);
xnor U5252 (N_5252,N_3537,N_2215);
or U5253 (N_5253,N_949,N_2779);
nor U5254 (N_5254,N_3906,N_2382);
nor U5255 (N_5255,N_794,N_2545);
nor U5256 (N_5256,N_2440,N_2359);
or U5257 (N_5257,N_3505,N_478);
or U5258 (N_5258,N_1580,N_3473);
or U5259 (N_5259,N_1729,N_1918);
nor U5260 (N_5260,N_1331,N_3124);
nand U5261 (N_5261,N_3746,N_2064);
and U5262 (N_5262,N_3650,N_1800);
nand U5263 (N_5263,N_288,N_1235);
or U5264 (N_5264,N_3102,N_2273);
and U5265 (N_5265,N_1926,N_4);
or U5266 (N_5266,N_3938,N_1671);
and U5267 (N_5267,N_2262,N_890);
or U5268 (N_5268,N_3002,N_3674);
nor U5269 (N_5269,N_3853,N_3013);
xnor U5270 (N_5270,N_2097,N_1842);
and U5271 (N_5271,N_3642,N_549);
nor U5272 (N_5272,N_3940,N_757);
nand U5273 (N_5273,N_196,N_2175);
and U5274 (N_5274,N_3868,N_3889);
or U5275 (N_5275,N_1064,N_3043);
nor U5276 (N_5276,N_109,N_246);
nand U5277 (N_5277,N_1710,N_1258);
nor U5278 (N_5278,N_3416,N_1911);
xor U5279 (N_5279,N_1326,N_410);
nor U5280 (N_5280,N_1223,N_2420);
and U5281 (N_5281,N_298,N_2371);
nand U5282 (N_5282,N_139,N_2578);
nor U5283 (N_5283,N_1260,N_595);
nand U5284 (N_5284,N_1032,N_311);
and U5285 (N_5285,N_1003,N_1565);
nor U5286 (N_5286,N_1005,N_1325);
or U5287 (N_5287,N_2847,N_2992);
nor U5288 (N_5288,N_685,N_3931);
nor U5289 (N_5289,N_3769,N_1776);
nor U5290 (N_5290,N_3870,N_45);
nor U5291 (N_5291,N_3915,N_1796);
nor U5292 (N_5292,N_476,N_2474);
and U5293 (N_5293,N_3392,N_858);
and U5294 (N_5294,N_2311,N_3351);
or U5295 (N_5295,N_2071,N_2572);
nor U5296 (N_5296,N_3890,N_48);
nor U5297 (N_5297,N_585,N_1215);
xor U5298 (N_5298,N_1742,N_2108);
and U5299 (N_5299,N_3574,N_3997);
or U5300 (N_5300,N_2164,N_392);
or U5301 (N_5301,N_2848,N_699);
nand U5302 (N_5302,N_3948,N_2023);
nor U5303 (N_5303,N_1689,N_3744);
nor U5304 (N_5304,N_979,N_2457);
nand U5305 (N_5305,N_3939,N_2011);
or U5306 (N_5306,N_1784,N_1993);
nand U5307 (N_5307,N_1877,N_1659);
nand U5308 (N_5308,N_1694,N_3130);
and U5309 (N_5309,N_2141,N_1554);
and U5310 (N_5310,N_2802,N_2333);
xnor U5311 (N_5311,N_711,N_909);
or U5312 (N_5312,N_1278,N_1967);
or U5313 (N_5313,N_1361,N_2211);
nand U5314 (N_5314,N_3857,N_1731);
and U5315 (N_5315,N_3284,N_627);
and U5316 (N_5316,N_73,N_2364);
and U5317 (N_5317,N_2698,N_1701);
and U5318 (N_5318,N_3580,N_3052);
or U5319 (N_5319,N_2823,N_250);
and U5320 (N_5320,N_3531,N_240);
nand U5321 (N_5321,N_144,N_935);
nand U5322 (N_5322,N_2302,N_3572);
and U5323 (N_5323,N_3903,N_3230);
xnor U5324 (N_5324,N_2004,N_2093);
nand U5325 (N_5325,N_375,N_273);
nor U5326 (N_5326,N_1381,N_209);
and U5327 (N_5327,N_528,N_3812);
xnor U5328 (N_5328,N_2162,N_810);
xor U5329 (N_5329,N_3288,N_1985);
nor U5330 (N_5330,N_3410,N_2046);
and U5331 (N_5331,N_2464,N_2191);
nand U5332 (N_5332,N_3345,N_2307);
xor U5333 (N_5333,N_380,N_2424);
xnor U5334 (N_5334,N_3450,N_3656);
and U5335 (N_5335,N_2587,N_3519);
nand U5336 (N_5336,N_342,N_2608);
xor U5337 (N_5337,N_316,N_3545);
nor U5338 (N_5338,N_3331,N_1177);
or U5339 (N_5339,N_186,N_2977);
and U5340 (N_5340,N_1019,N_3047);
xnor U5341 (N_5341,N_2768,N_3589);
xor U5342 (N_5342,N_3882,N_2974);
nand U5343 (N_5343,N_3179,N_3298);
or U5344 (N_5344,N_2942,N_79);
and U5345 (N_5345,N_59,N_1036);
or U5346 (N_5346,N_2725,N_1035);
or U5347 (N_5347,N_332,N_2646);
nor U5348 (N_5348,N_2532,N_2841);
and U5349 (N_5349,N_2433,N_3131);
xor U5350 (N_5350,N_2901,N_2621);
nor U5351 (N_5351,N_902,N_1684);
xnor U5352 (N_5352,N_720,N_873);
nor U5353 (N_5353,N_837,N_2016);
nand U5354 (N_5354,N_3777,N_2212);
nor U5355 (N_5355,N_3411,N_101);
xor U5356 (N_5356,N_176,N_3255);
nand U5357 (N_5357,N_1780,N_3983);
and U5358 (N_5358,N_2398,N_1091);
or U5359 (N_5359,N_3171,N_673);
and U5360 (N_5360,N_22,N_1134);
nor U5361 (N_5361,N_1563,N_650);
and U5362 (N_5362,N_931,N_106);
nor U5363 (N_5363,N_1474,N_3391);
and U5364 (N_5364,N_3054,N_2695);
nor U5365 (N_5365,N_1481,N_839);
nand U5366 (N_5366,N_2316,N_1723);
nand U5367 (N_5367,N_675,N_3141);
and U5368 (N_5368,N_3951,N_903);
and U5369 (N_5369,N_3895,N_2686);
and U5370 (N_5370,N_480,N_1732);
nand U5371 (N_5371,N_3947,N_2286);
xor U5372 (N_5372,N_477,N_1165);
or U5373 (N_5373,N_561,N_3698);
or U5374 (N_5374,N_1810,N_1767);
nand U5375 (N_5375,N_3536,N_3730);
and U5376 (N_5376,N_1765,N_3645);
and U5377 (N_5377,N_943,N_3205);
nand U5378 (N_5378,N_1081,N_2121);
xnor U5379 (N_5379,N_2602,N_632);
xor U5380 (N_5380,N_1262,N_279);
or U5381 (N_5381,N_1928,N_1337);
nor U5382 (N_5382,N_1404,N_2869);
or U5383 (N_5383,N_691,N_1513);
nand U5384 (N_5384,N_3528,N_2934);
nand U5385 (N_5385,N_3659,N_1581);
and U5386 (N_5386,N_2570,N_730);
nand U5387 (N_5387,N_2616,N_2659);
or U5388 (N_5388,N_1644,N_2528);
or U5389 (N_5389,N_294,N_2539);
nor U5390 (N_5390,N_1656,N_2393);
nor U5391 (N_5391,N_2801,N_3775);
and U5392 (N_5392,N_2523,N_2834);
nand U5393 (N_5393,N_3641,N_3856);
nand U5394 (N_5394,N_2735,N_1994);
or U5395 (N_5395,N_2001,N_3726);
or U5396 (N_5396,N_84,N_786);
nor U5397 (N_5397,N_2171,N_2082);
xor U5398 (N_5398,N_667,N_875);
nand U5399 (N_5399,N_3791,N_2720);
and U5400 (N_5400,N_3024,N_2907);
and U5401 (N_5401,N_3018,N_372);
or U5402 (N_5402,N_3457,N_3184);
xnor U5403 (N_5403,N_191,N_1514);
nor U5404 (N_5404,N_1957,N_2030);
nand U5405 (N_5405,N_3357,N_3469);
or U5406 (N_5406,N_654,N_2362);
and U5407 (N_5407,N_1114,N_358);
nand U5408 (N_5408,N_1393,N_2143);
xor U5409 (N_5409,N_1186,N_1876);
nor U5410 (N_5410,N_851,N_23);
nand U5411 (N_5411,N_472,N_1758);
or U5412 (N_5412,N_3335,N_1244);
or U5413 (N_5413,N_72,N_1039);
nand U5414 (N_5414,N_1067,N_2521);
or U5415 (N_5415,N_1397,N_3244);
nor U5416 (N_5416,N_2692,N_1461);
xor U5417 (N_5417,N_2751,N_1649);
or U5418 (N_5418,N_1668,N_3062);
and U5419 (N_5419,N_1703,N_3425);
nor U5420 (N_5420,N_6,N_2178);
or U5421 (N_5421,N_1498,N_710);
nand U5422 (N_5422,N_194,N_3267);
or U5423 (N_5423,N_2894,N_3827);
nand U5424 (N_5424,N_860,N_396);
nand U5425 (N_5425,N_1140,N_2068);
and U5426 (N_5426,N_450,N_2729);
and U5427 (N_5427,N_2493,N_1941);
and U5428 (N_5428,N_2547,N_371);
and U5429 (N_5429,N_2060,N_578);
nor U5430 (N_5430,N_2875,N_3750);
nand U5431 (N_5431,N_1569,N_3954);
or U5432 (N_5432,N_1217,N_3157);
and U5433 (N_5433,N_985,N_2274);
nand U5434 (N_5434,N_2682,N_2781);
and U5435 (N_5435,N_1558,N_1428);
nor U5436 (N_5436,N_29,N_457);
nor U5437 (N_5437,N_3277,N_3170);
or U5438 (N_5438,N_2032,N_1509);
nand U5439 (N_5439,N_51,N_3655);
nor U5440 (N_5440,N_3381,N_788);
nand U5441 (N_5441,N_1055,N_2514);
nor U5442 (N_5442,N_1661,N_2358);
and U5443 (N_5443,N_3924,N_2219);
or U5444 (N_5444,N_813,N_2687);
nor U5445 (N_5445,N_3238,N_401);
and U5446 (N_5446,N_762,N_1691);
and U5447 (N_5447,N_548,N_1577);
xor U5448 (N_5448,N_3885,N_307);
or U5449 (N_5449,N_354,N_1736);
and U5450 (N_5450,N_3691,N_236);
xor U5451 (N_5451,N_2116,N_778);
xnor U5452 (N_5452,N_2168,N_1655);
nand U5453 (N_5453,N_2017,N_1135);
or U5454 (N_5454,N_202,N_3315);
or U5455 (N_5455,N_2776,N_2664);
nand U5456 (N_5456,N_3569,N_3444);
nand U5457 (N_5457,N_2233,N_2117);
nand U5458 (N_5458,N_3845,N_2881);
nor U5459 (N_5459,N_867,N_1491);
nor U5460 (N_5460,N_838,N_2496);
and U5461 (N_5461,N_2043,N_801);
and U5462 (N_5462,N_2724,N_1836);
nand U5463 (N_5463,N_239,N_2508);
nor U5464 (N_5464,N_2716,N_736);
or U5465 (N_5465,N_258,N_266);
or U5466 (N_5466,N_159,N_808);
or U5467 (N_5467,N_2149,N_855);
and U5468 (N_5468,N_2588,N_3512);
nand U5469 (N_5469,N_603,N_2384);
xor U5470 (N_5470,N_2713,N_3440);
and U5471 (N_5471,N_2945,N_110);
nand U5472 (N_5472,N_3905,N_817);
xnor U5473 (N_5473,N_2151,N_1142);
nand U5474 (N_5474,N_1583,N_3297);
or U5475 (N_5475,N_816,N_2582);
nor U5476 (N_5476,N_3759,N_913);
and U5477 (N_5477,N_3843,N_3786);
nand U5478 (N_5478,N_1348,N_1538);
xor U5479 (N_5479,N_2218,N_3969);
and U5480 (N_5480,N_2706,N_1270);
or U5481 (N_5481,N_1161,N_3668);
nand U5482 (N_5482,N_1612,N_655);
or U5483 (N_5483,N_406,N_2086);
or U5484 (N_5484,N_3337,N_716);
xor U5485 (N_5485,N_3735,N_2912);
and U5486 (N_5486,N_1463,N_2987);
nor U5487 (N_5487,N_108,N_152);
nand U5488 (N_5488,N_3122,N_309);
nor U5489 (N_5489,N_3011,N_76);
nor U5490 (N_5490,N_1440,N_2104);
nand U5491 (N_5491,N_2025,N_1133);
nand U5492 (N_5492,N_2343,N_2208);
nor U5493 (N_5493,N_643,N_3917);
or U5494 (N_5494,N_3261,N_3970);
or U5495 (N_5495,N_3376,N_3014);
nand U5496 (N_5496,N_1085,N_2678);
nand U5497 (N_5497,N_2347,N_3779);
or U5498 (N_5498,N_2091,N_242);
nor U5499 (N_5499,N_3278,N_3059);
nand U5500 (N_5500,N_598,N_1455);
nand U5501 (N_5501,N_1416,N_2221);
nor U5502 (N_5502,N_670,N_2962);
nand U5503 (N_5503,N_3456,N_962);
and U5504 (N_5504,N_2239,N_2614);
nand U5505 (N_5505,N_20,N_662);
nand U5506 (N_5506,N_3504,N_2584);
and U5507 (N_5507,N_2209,N_3363);
nand U5508 (N_5508,N_1490,N_1938);
and U5509 (N_5509,N_377,N_951);
and U5510 (N_5510,N_306,N_2799);
or U5511 (N_5511,N_841,N_3127);
or U5512 (N_5512,N_310,N_313);
or U5513 (N_5513,N_3070,N_1556);
nand U5514 (N_5514,N_3754,N_1980);
and U5515 (N_5515,N_3325,N_3855);
and U5516 (N_5516,N_8,N_153);
xor U5517 (N_5517,N_3079,N_2348);
and U5518 (N_5518,N_3125,N_2369);
xnor U5519 (N_5519,N_1484,N_2477);
and U5520 (N_5520,N_2668,N_2903);
or U5521 (N_5521,N_3364,N_1321);
and U5522 (N_5522,N_2566,N_282);
or U5523 (N_5523,N_2712,N_216);
nand U5524 (N_5524,N_2501,N_2563);
or U5525 (N_5525,N_3380,N_3053);
and U5526 (N_5526,N_3445,N_2270);
nor U5527 (N_5527,N_1699,N_565);
nand U5528 (N_5528,N_2980,N_2817);
and U5529 (N_5529,N_3503,N_97);
nand U5530 (N_5530,N_2484,N_3705);
or U5531 (N_5531,N_3150,N_2158);
nor U5532 (N_5532,N_47,N_3167);
nand U5533 (N_5533,N_2576,N_272);
or U5534 (N_5534,N_1216,N_496);
and U5535 (N_5535,N_741,N_3629);
nor U5536 (N_5536,N_635,N_1002);
nand U5537 (N_5537,N_3276,N_3697);
and U5538 (N_5538,N_506,N_554);
nor U5539 (N_5539,N_1739,N_2100);
nand U5540 (N_5540,N_1866,N_936);
nand U5541 (N_5541,N_676,N_464);
nor U5542 (N_5542,N_1169,N_1276);
or U5543 (N_5543,N_3458,N_614);
and U5544 (N_5544,N_2377,N_2067);
xor U5545 (N_5545,N_693,N_2378);
and U5546 (N_5546,N_2895,N_924);
or U5547 (N_5547,N_3178,N_2886);
or U5548 (N_5548,N_3837,N_2375);
xor U5549 (N_5549,N_3115,N_2062);
or U5550 (N_5550,N_3177,N_2332);
nand U5551 (N_5551,N_3283,N_481);
or U5552 (N_5552,N_1669,N_1126);
and U5553 (N_5553,N_3813,N_1080);
nor U5554 (N_5554,N_2832,N_349);
xnor U5555 (N_5555,N_2829,N_2396);
and U5556 (N_5556,N_102,N_454);
nand U5557 (N_5557,N_1619,N_198);
and U5558 (N_5558,N_1289,N_2814);
nor U5559 (N_5559,N_370,N_1901);
xor U5560 (N_5560,N_758,N_1532);
or U5561 (N_5561,N_3922,N_2352);
or U5562 (N_5562,N_1415,N_3055);
or U5563 (N_5563,N_917,N_3407);
or U5564 (N_5564,N_1642,N_3249);
nor U5565 (N_5565,N_911,N_3447);
nor U5566 (N_5566,N_3262,N_3756);
nor U5567 (N_5567,N_348,N_3996);
and U5568 (N_5568,N_612,N_3878);
nand U5569 (N_5569,N_2669,N_3442);
nand U5570 (N_5570,N_3987,N_486);
nand U5571 (N_5571,N_2905,N_3144);
or U5572 (N_5572,N_3829,N_248);
xnor U5573 (N_5573,N_1171,N_2303);
nand U5574 (N_5574,N_3795,N_845);
or U5575 (N_5575,N_3136,N_283);
or U5576 (N_5576,N_3871,N_2533);
or U5577 (N_5577,N_2283,N_796);
nor U5578 (N_5578,N_2816,N_804);
and U5579 (N_5579,N_2293,N_2783);
nor U5580 (N_5580,N_1304,N_1269);
nand U5581 (N_5581,N_2870,N_1754);
and U5582 (N_5582,N_2247,N_2950);
or U5583 (N_5583,N_2952,N_1243);
and U5584 (N_5584,N_2497,N_3212);
and U5585 (N_5585,N_46,N_3590);
nand U5586 (N_5586,N_3172,N_2256);
or U5587 (N_5587,N_1633,N_2372);
nor U5588 (N_5588,N_3209,N_2047);
or U5589 (N_5589,N_1737,N_2111);
or U5590 (N_5590,N_1041,N_2594);
and U5591 (N_5591,N_2419,N_946);
or U5592 (N_5592,N_3751,N_2677);
xnor U5593 (N_5593,N_1148,N_672);
nand U5594 (N_5594,N_2249,N_63);
nand U5595 (N_5595,N_3620,N_618);
or U5596 (N_5596,N_3074,N_779);
or U5597 (N_5597,N_1207,N_3941);
or U5598 (N_5598,N_763,N_1594);
and U5599 (N_5599,N_948,N_3814);
nand U5600 (N_5600,N_3755,N_466);
nor U5601 (N_5601,N_700,N_1986);
xnor U5602 (N_5602,N_2294,N_3040);
and U5603 (N_5603,N_1237,N_2213);
nor U5604 (N_5604,N_2125,N_965);
nor U5605 (N_5605,N_1625,N_637);
nor U5606 (N_5606,N_1706,N_1349);
xnor U5607 (N_5607,N_977,N_622);
and U5608 (N_5608,N_3272,N_1948);
nor U5609 (N_5609,N_3427,N_2658);
nor U5610 (N_5610,N_3990,N_893);
nor U5611 (N_5611,N_1053,N_3937);
nor U5612 (N_5612,N_597,N_1605);
or U5613 (N_5613,N_3907,N_2252);
nor U5614 (N_5614,N_2381,N_3094);
nand U5615 (N_5615,N_3558,N_891);
or U5616 (N_5616,N_1937,N_1962);
and U5617 (N_5617,N_2565,N_1027);
nor U5618 (N_5618,N_3958,N_1814);
nand U5619 (N_5619,N_1608,N_3451);
nand U5620 (N_5620,N_3796,N_774);
nor U5621 (N_5621,N_168,N_3553);
nand U5622 (N_5622,N_27,N_1496);
xnor U5623 (N_5623,N_1579,N_1769);
xor U5624 (N_5624,N_1777,N_2860);
nand U5625 (N_5625,N_3663,N_888);
and U5626 (N_5626,N_971,N_439);
nor U5627 (N_5627,N_3522,N_3570);
nand U5628 (N_5628,N_1940,N_3116);
nor U5629 (N_5629,N_604,N_2641);
nor U5630 (N_5630,N_424,N_3499);
and U5631 (N_5631,N_3488,N_2764);
or U5632 (N_5632,N_3626,N_1833);
xor U5633 (N_5633,N_926,N_2187);
nor U5634 (N_5634,N_573,N_3242);
nand U5635 (N_5635,N_1473,N_1925);
xnor U5636 (N_5636,N_1875,N_284);
and U5637 (N_5637,N_1791,N_355);
nor U5638 (N_5638,N_381,N_1872);
and U5639 (N_5639,N_682,N_2512);
nand U5640 (N_5640,N_674,N_403);
nand U5641 (N_5641,N_3119,N_3601);
nand U5642 (N_5642,N_980,N_1861);
or U5643 (N_5643,N_2671,N_3850);
or U5644 (N_5644,N_658,N_2718);
xnor U5645 (N_5645,N_3886,N_2013);
nand U5646 (N_5646,N_3158,N_1574);
or U5647 (N_5647,N_167,N_393);
nand U5648 (N_5648,N_1623,N_2986);
or U5649 (N_5649,N_1596,N_830);
nor U5650 (N_5650,N_2737,N_1726);
or U5651 (N_5651,N_3872,N_383);
nor U5652 (N_5652,N_3844,N_895);
and U5653 (N_5653,N_2113,N_2320);
and U5654 (N_5654,N_669,N_1634);
xnor U5655 (N_5655,N_2540,N_1447);
nor U5656 (N_5656,N_3361,N_25);
or U5657 (N_5657,N_1969,N_1813);
nor U5658 (N_5658,N_2932,N_3603);
and U5659 (N_5659,N_2119,N_3186);
or U5660 (N_5660,N_2915,N_1167);
and U5661 (N_5661,N_799,N_715);
nor U5662 (N_5662,N_3294,N_1102);
xor U5663 (N_5663,N_462,N_3721);
nand U5664 (N_5664,N_2853,N_2390);
nor U5665 (N_5665,N_892,N_3108);
or U5666 (N_5666,N_3680,N_2600);
or U5667 (N_5667,N_2522,N_1355);
xor U5668 (N_5668,N_2813,N_67);
and U5669 (N_5669,N_3520,N_3075);
xor U5670 (N_5670,N_2822,N_533);
nand U5671 (N_5671,N_3848,N_1453);
nand U5672 (N_5672,N_2971,N_2723);
nand U5673 (N_5673,N_3804,N_3265);
and U5674 (N_5674,N_2892,N_1146);
xnor U5675 (N_5675,N_2147,N_3343);
xnor U5676 (N_5676,N_1332,N_3324);
or U5677 (N_5677,N_3218,N_3826);
xor U5678 (N_5678,N_490,N_2133);
and U5679 (N_5679,N_1456,N_32);
and U5680 (N_5680,N_1761,N_173);
nor U5681 (N_5681,N_1485,N_1459);
nand U5682 (N_5682,N_2548,N_681);
nor U5683 (N_5683,N_3719,N_2727);
xnor U5684 (N_5684,N_2192,N_3604);
nand U5685 (N_5685,N_988,N_1725);
and U5686 (N_5686,N_1069,N_3190);
or U5687 (N_5687,N_507,N_3967);
or U5688 (N_5688,N_1929,N_570);
and U5689 (N_5689,N_1364,N_2909);
xor U5690 (N_5690,N_1681,N_2715);
and U5691 (N_5691,N_1899,N_433);
or U5692 (N_5692,N_431,N_661);
nor U5693 (N_5693,N_2554,N_2631);
or U5694 (N_5694,N_1636,N_3431);
and U5695 (N_5695,N_1317,N_2642);
nor U5696 (N_5696,N_991,N_53);
and U5697 (N_5697,N_2858,N_1768);
or U5698 (N_5698,N_195,N_2763);
and U5699 (N_5699,N_2144,N_1822);
and U5700 (N_5700,N_2855,N_3093);
or U5701 (N_5701,N_3341,N_3643);
nand U5702 (N_5702,N_3290,N_577);
or U5703 (N_5703,N_205,N_165);
nor U5704 (N_5704,N_1426,N_3386);
nor U5705 (N_5705,N_278,N_1651);
or U5706 (N_5706,N_2118,N_3299);
or U5707 (N_5707,N_155,N_3696);
nand U5708 (N_5708,N_2385,N_1518);
xnor U5709 (N_5709,N_1855,N_2052);
and U5710 (N_5710,N_3506,N_2142);
nor U5711 (N_5711,N_1339,N_2597);
xor U5712 (N_5712,N_771,N_3662);
nor U5713 (N_5713,N_1844,N_1369);
nor U5714 (N_5714,N_2167,N_1628);
or U5715 (N_5715,N_2391,N_3773);
nand U5716 (N_5716,N_1912,N_3036);
nor U5717 (N_5717,N_123,N_409);
and U5718 (N_5718,N_3986,N_592);
nor U5719 (N_5719,N_1900,N_3950);
and U5720 (N_5720,N_937,N_1141);
xnor U5721 (N_5721,N_1873,N_1163);
nand U5722 (N_5722,N_3358,N_1803);
and U5723 (N_5723,N_899,N_2674);
nand U5724 (N_5724,N_1144,N_287);
or U5725 (N_5725,N_2126,N_1987);
nor U5726 (N_5726,N_3586,N_761);
or U5727 (N_5727,N_118,N_2893);
nand U5728 (N_5728,N_2031,N_1603);
nand U5729 (N_5729,N_2447,N_3311);
nor U5730 (N_5730,N_33,N_1522);
nand U5731 (N_5731,N_1598,N_1105);
nor U5732 (N_5732,N_1264,N_296);
or U5733 (N_5733,N_2287,N_912);
or U5734 (N_5734,N_3563,N_62);
nor U5735 (N_5735,N_677,N_1248);
nand U5736 (N_5736,N_2906,N_3088);
xnor U5737 (N_5737,N_1026,N_3133);
and U5738 (N_5738,N_3824,N_3401);
xor U5739 (N_5739,N_3701,N_1527);
and U5740 (N_5740,N_1034,N_3535);
xor U5741 (N_5741,N_2150,N_975);
nor U5742 (N_5742,N_3232,N_1864);
xnor U5743 (N_5743,N_75,N_3415);
or U5744 (N_5744,N_1759,N_1757);
and U5745 (N_5745,N_2328,N_1293);
nand U5746 (N_5746,N_3162,N_1164);
and U5747 (N_5747,N_199,N_351);
nor U5748 (N_5748,N_3296,N_3687);
or U5749 (N_5749,N_3224,N_2045);
and U5750 (N_5750,N_3097,N_3215);
or U5751 (N_5751,N_929,N_2931);
or U5752 (N_5752,N_2811,N_1722);
and U5753 (N_5753,N_1954,N_1838);
or U5754 (N_5754,N_1709,N_1384);
and U5755 (N_5755,N_2132,N_3628);
nor U5756 (N_5756,N_1599,N_2335);
or U5757 (N_5757,N_3566,N_3832);
xor U5758 (N_5758,N_3902,N_2667);
xnor U5759 (N_5759,N_3665,N_2561);
and U5760 (N_5760,N_1089,N_1356);
nor U5761 (N_5761,N_257,N_692);
nor U5762 (N_5762,N_1919,N_901);
nand U5763 (N_5763,N_1566,N_1407);
nand U5764 (N_5764,N_986,N_2135);
or U5765 (N_5765,N_3625,N_13);
xor U5766 (N_5766,N_3943,N_2028);
or U5767 (N_5767,N_1952,N_211);
xnor U5768 (N_5768,N_1988,N_3541);
nor U5769 (N_5769,N_2615,N_3595);
nor U5770 (N_5770,N_1905,N_3477);
nor U5771 (N_5771,N_2936,N_1386);
or U5772 (N_5772,N_1471,N_3627);
and U5773 (N_5773,N_535,N_1502);
nor U5774 (N_5774,N_1843,N_3388);
xnor U5775 (N_5775,N_2623,N_2156);
nor U5776 (N_5776,N_2446,N_379);
and U5777 (N_5777,N_1774,N_1519);
and U5778 (N_5778,N_2904,N_2586);
nor U5779 (N_5779,N_1330,N_2596);
nor U5780 (N_5780,N_2301,N_2379);
and U5781 (N_5781,N_3114,N_3316);
and U5782 (N_5782,N_759,N_776);
or U5783 (N_5783,N_3350,N_448);
and U5784 (N_5784,N_1611,N_3894);
nor U5785 (N_5785,N_3268,N_1131);
and U5786 (N_5786,N_2914,N_289);
and U5787 (N_5787,N_461,N_1088);
nor U5788 (N_5788,N_135,N_360);
nor U5789 (N_5789,N_467,N_934);
nor U5790 (N_5790,N_1329,N_99);
nand U5791 (N_5791,N_232,N_3152);
or U5792 (N_5792,N_3926,N_3100);
nand U5793 (N_5793,N_408,N_2298);
nand U5794 (N_5794,N_2949,N_2296);
or U5795 (N_5795,N_1172,N_3610);
nand U5796 (N_5796,N_2828,N_21);
or U5797 (N_5797,N_1030,N_2524);
nand U5798 (N_5798,N_678,N_1999);
nand U5799 (N_5799,N_541,N_2039);
or U5800 (N_5800,N_2711,N_122);
or U5801 (N_5801,N_1454,N_2138);
nand U5802 (N_5802,N_2478,N_1856);
nor U5803 (N_5803,N_3616,N_2638);
and U5804 (N_5804,N_2701,N_2353);
and U5805 (N_5805,N_3513,N_721);
nand U5806 (N_5806,N_1851,N_1624);
xnor U5807 (N_5807,N_378,N_3168);
xnor U5808 (N_5808,N_819,N_2402);
or U5809 (N_5809,N_0,N_1018);
nor U5810 (N_5810,N_2647,N_328);
or U5811 (N_5811,N_3834,N_1231);
nand U5812 (N_5812,N_2395,N_3693);
nor U5813 (N_5813,N_2988,N_1662);
nor U5814 (N_5814,N_2363,N_3714);
nor U5815 (N_5815,N_1312,N_1009);
nand U5816 (N_5816,N_1334,N_2843);
or U5817 (N_5817,N_2900,N_228);
xnor U5818 (N_5818,N_729,N_1402);
and U5819 (N_5819,N_2010,N_555);
or U5820 (N_5820,N_2244,N_2911);
or U5821 (N_5821,N_642,N_2978);
or U5822 (N_5822,N_70,N_1516);
or U5823 (N_5823,N_842,N_3313);
nand U5824 (N_5824,N_419,N_3575);
nand U5825 (N_5825,N_3377,N_833);
and U5826 (N_5826,N_2585,N_2083);
nor U5827 (N_5827,N_1103,N_789);
nor U5828 (N_5828,N_2598,N_2197);
nor U5829 (N_5829,N_742,N_2948);
and U5830 (N_5830,N_1336,N_1246);
xnor U5831 (N_5831,N_644,N_479);
nor U5832 (N_5832,N_1534,N_1157);
or U5833 (N_5833,N_2626,N_3607);
nor U5834 (N_5834,N_1854,N_602);
or U5835 (N_5835,N_3289,N_3395);
nor U5836 (N_5836,N_843,N_2922);
and U5837 (N_5837,N_41,N_814);
or U5838 (N_5838,N_2476,N_2309);
and U5839 (N_5839,N_1116,N_428);
nand U5840 (N_5840,N_2752,N_1886);
nand U5841 (N_5841,N_3256,N_1342);
or U5842 (N_5842,N_2183,N_607);
nand U5843 (N_5843,N_2998,N_950);
or U5844 (N_5844,N_341,N_2973);
nor U5845 (N_5845,N_2182,N_3591);
nor U5846 (N_5846,N_3470,N_1801);
xnor U5847 (N_5847,N_212,N_444);
nand U5848 (N_5848,N_1354,N_337);
and U5849 (N_5849,N_2491,N_2181);
or U5850 (N_5850,N_547,N_806);
nand U5851 (N_5851,N_1350,N_178);
nor U5852 (N_5852,N_2898,N_2885);
and U5853 (N_5853,N_2557,N_3463);
nor U5854 (N_5854,N_3293,N_504);
nand U5855 (N_5855,N_3160,N_1584);
nand U5856 (N_5856,N_2451,N_113);
xnor U5857 (N_5857,N_3612,N_3865);
and U5858 (N_5858,N_157,N_1367);
nand U5859 (N_5859,N_339,N_1155);
and U5860 (N_5860,N_2292,N_1442);
nand U5861 (N_5861,N_2242,N_3568);
nor U5862 (N_5862,N_1156,N_1476);
and U5863 (N_5863,N_1717,N_487);
and U5864 (N_5864,N_1802,N_876);
nand U5865 (N_5865,N_3208,N_2960);
nor U5866 (N_5866,N_2824,N_3840);
nor U5867 (N_5867,N_315,N_3472);
xnor U5868 (N_5868,N_2876,N_3137);
nor U5869 (N_5869,N_42,N_2990);
and U5870 (N_5870,N_414,N_886);
and U5871 (N_5871,N_170,N_3180);
nor U5872 (N_5872,N_1751,N_3025);
and U5873 (N_5873,N_2073,N_2388);
nor U5874 (N_5874,N_3694,N_3587);
nor U5875 (N_5875,N_3639,N_1137);
nand U5876 (N_5876,N_1808,N_587);
and U5877 (N_5877,N_1458,N_3196);
xor U5878 (N_5878,N_1601,N_105);
nand U5879 (N_5879,N_3183,N_3282);
and U5880 (N_5880,N_365,N_2277);
nand U5881 (N_5881,N_2500,N_3679);
nor U5882 (N_5882,N_582,N_3547);
and U5883 (N_5883,N_1252,N_129);
and U5884 (N_5884,N_3454,N_923);
nor U5885 (N_5885,N_686,N_3588);
nor U5886 (N_5886,N_1958,N_1281);
and U5887 (N_5887,N_3007,N_137);
nand U5888 (N_5888,N_2399,N_1588);
or U5889 (N_5889,N_1804,N_1535);
and U5890 (N_5890,N_3403,N_1560);
nor U5891 (N_5891,N_921,N_3555);
nand U5892 (N_5892,N_323,N_1322);
nand U5893 (N_5893,N_3608,N_523);
nor U5894 (N_5894,N_3634,N_689);
nor U5895 (N_5895,N_373,N_215);
and U5896 (N_5896,N_930,N_3646);
nor U5897 (N_5897,N_2061,N_269);
or U5898 (N_5898,N_2525,N_3406);
or U5899 (N_5899,N_1253,N_2471);
nor U5900 (N_5900,N_2223,N_933);
or U5901 (N_5901,N_2059,N_2128);
xnor U5902 (N_5902,N_2550,N_399);
nand U5903 (N_5903,N_1869,N_3228);
or U5904 (N_5904,N_871,N_2744);
nand U5905 (N_5905,N_2084,N_3402);
nand U5906 (N_5906,N_2660,N_2511);
or U5907 (N_5907,N_3899,N_2793);
and U5908 (N_5908,N_3163,N_2434);
and U5909 (N_5909,N_1214,N_1850);
nor U5910 (N_5910,N_3365,N_2115);
or U5911 (N_5911,N_1226,N_3372);
and U5912 (N_5912,N_3876,N_96);
nor U5913 (N_5913,N_2340,N_1939);
nor U5914 (N_5914,N_969,N_3640);
and U5915 (N_5915,N_1548,N_1191);
nand U5916 (N_5916,N_719,N_3414);
nor U5917 (N_5917,N_3502,N_263);
nand U5918 (N_5918,N_1576,N_56);
or U5919 (N_5919,N_1983,N_1609);
nand U5920 (N_5920,N_1414,N_2160);
and U5921 (N_5921,N_2624,N_1549);
nand U5922 (N_5922,N_1073,N_3787);
and U5923 (N_5923,N_1614,N_2526);
or U5924 (N_5924,N_324,N_1552);
or U5925 (N_5925,N_3875,N_2956);
xor U5926 (N_5926,N_703,N_3729);
or U5927 (N_5927,N_1561,N_1927);
and U5928 (N_5928,N_520,N_64);
nor U5929 (N_5929,N_2226,N_2075);
and U5930 (N_5930,N_2796,N_1450);
nand U5931 (N_5931,N_3334,N_3949);
or U5932 (N_5932,N_2005,N_1847);
and U5933 (N_5933,N_1947,N_1687);
and U5934 (N_5934,N_1976,N_2628);
xnor U5935 (N_5935,N_1296,N_201);
and U5936 (N_5936,N_515,N_2227);
or U5937 (N_5937,N_2935,N_3861);
or U5938 (N_5938,N_770,N_1821);
nor U5939 (N_5939,N_2704,N_734);
and U5940 (N_5940,N_3349,N_906);
xnor U5941 (N_5941,N_140,N_957);
nor U5942 (N_5942,N_3690,N_3565);
nor U5943 (N_5943,N_389,N_3237);
nand U5944 (N_5944,N_1879,N_251);
xor U5945 (N_5945,N_823,N_2078);
nor U5946 (N_5946,N_3887,N_3952);
or U5947 (N_5947,N_3965,N_3308);
nand U5948 (N_5948,N_530,N_3239);
nor U5949 (N_5949,N_3724,N_2350);
or U5950 (N_5950,N_2232,N_420);
or U5951 (N_5951,N_2979,N_1913);
nor U5952 (N_5952,N_3155,N_1953);
nand U5953 (N_5953,N_2409,N_2529);
nand U5954 (N_5954,N_3688,N_2918);
nor U5955 (N_5955,N_1385,N_2773);
and U5956 (N_5956,N_3068,N_3039);
nand U5957 (N_5957,N_726,N_3384);
or U5958 (N_5958,N_1319,N_1830);
nand U5959 (N_5959,N_2423,N_1482);
nand U5960 (N_5960,N_3782,N_3318);
nand U5961 (N_5961,N_3084,N_2663);
or U5962 (N_5962,N_2310,N_1892);
and U5963 (N_5963,N_3637,N_854);
and U5964 (N_5964,N_2489,N_493);
and U5965 (N_5965,N_2058,N_3169);
or U5966 (N_5966,N_2264,N_1071);
nor U5967 (N_5967,N_1031,N_1657);
nand U5968 (N_5968,N_2186,N_2306);
or U5969 (N_5969,N_1301,N_610);
and U5970 (N_5970,N_749,N_904);
nand U5971 (N_5971,N_3747,N_3259);
nor U5972 (N_5972,N_1272,N_536);
xnor U5973 (N_5973,N_3438,N_3732);
nand U5974 (N_5974,N_3396,N_1868);
nand U5975 (N_5975,N_474,N_3111);
nand U5976 (N_5976,N_1870,N_85);
nor U5977 (N_5977,N_229,N_3354);
nand U5978 (N_5978,N_3930,N_2241);
xnor U5979 (N_5979,N_1479,N_2088);
or U5980 (N_5980,N_1638,N_1310);
nor U5981 (N_5981,N_3828,N_963);
or U5982 (N_5982,N_2106,N_1462);
nor U5983 (N_5983,N_652,N_2878);
or U5984 (N_5984,N_3880,N_3146);
nand U5985 (N_5985,N_1212,N_2207);
or U5986 (N_5986,N_254,N_2697);
and U5987 (N_5987,N_525,N_764);
nand U5988 (N_5988,N_3560,N_1242);
or U5989 (N_5989,N_1438,N_1487);
or U5990 (N_5990,N_197,N_1090);
nand U5991 (N_5991,N_285,N_1486);
or U5992 (N_5992,N_1075,N_3534);
and U5993 (N_5993,N_1418,N_1512);
and U5994 (N_5994,N_1575,N_119);
nor U5995 (N_5995,N_3301,N_3006);
nand U5996 (N_5996,N_1626,N_3592);
nand U5997 (N_5997,N_3739,N_1199);
nand U5998 (N_5998,N_453,N_1254);
and U5999 (N_5999,N_1946,N_2670);
or U6000 (N_6000,N_1816,N_271);
or U6001 (N_6001,N_3601,N_2531);
xnor U6002 (N_6002,N_2920,N_1932);
nand U6003 (N_6003,N_258,N_950);
nand U6004 (N_6004,N_2328,N_3811);
or U6005 (N_6005,N_3096,N_3156);
nor U6006 (N_6006,N_2786,N_2326);
nand U6007 (N_6007,N_3389,N_1796);
or U6008 (N_6008,N_1264,N_866);
nor U6009 (N_6009,N_3879,N_2303);
nand U6010 (N_6010,N_2405,N_170);
nor U6011 (N_6011,N_708,N_1395);
or U6012 (N_6012,N_3060,N_2020);
and U6013 (N_6013,N_3578,N_2646);
or U6014 (N_6014,N_2347,N_3431);
xnor U6015 (N_6015,N_1470,N_993);
or U6016 (N_6016,N_3773,N_209);
and U6017 (N_6017,N_2908,N_797);
and U6018 (N_6018,N_436,N_3478);
xnor U6019 (N_6019,N_3902,N_3470);
nor U6020 (N_6020,N_3551,N_3930);
nand U6021 (N_6021,N_1371,N_48);
nor U6022 (N_6022,N_240,N_2333);
nand U6023 (N_6023,N_256,N_357);
and U6024 (N_6024,N_125,N_3687);
nand U6025 (N_6025,N_1266,N_3442);
or U6026 (N_6026,N_3710,N_1464);
or U6027 (N_6027,N_1257,N_1881);
and U6028 (N_6028,N_3876,N_2630);
or U6029 (N_6029,N_693,N_2493);
or U6030 (N_6030,N_391,N_2807);
or U6031 (N_6031,N_2631,N_690);
nand U6032 (N_6032,N_3957,N_1784);
and U6033 (N_6033,N_545,N_2961);
xor U6034 (N_6034,N_2153,N_1319);
and U6035 (N_6035,N_908,N_2743);
nand U6036 (N_6036,N_2860,N_449);
or U6037 (N_6037,N_1492,N_3499);
and U6038 (N_6038,N_3025,N_2089);
nand U6039 (N_6039,N_2893,N_676);
nand U6040 (N_6040,N_297,N_716);
or U6041 (N_6041,N_1703,N_609);
and U6042 (N_6042,N_1298,N_2307);
and U6043 (N_6043,N_3690,N_284);
nor U6044 (N_6044,N_652,N_1885);
nand U6045 (N_6045,N_2851,N_643);
nor U6046 (N_6046,N_1688,N_878);
or U6047 (N_6047,N_3863,N_3926);
nand U6048 (N_6048,N_1509,N_751);
and U6049 (N_6049,N_1171,N_2781);
xor U6050 (N_6050,N_1974,N_1266);
nor U6051 (N_6051,N_2641,N_1705);
or U6052 (N_6052,N_311,N_737);
nand U6053 (N_6053,N_727,N_3056);
or U6054 (N_6054,N_1302,N_3165);
or U6055 (N_6055,N_2661,N_2018);
or U6056 (N_6056,N_3535,N_857);
and U6057 (N_6057,N_119,N_1152);
nand U6058 (N_6058,N_940,N_1371);
nand U6059 (N_6059,N_3966,N_1861);
and U6060 (N_6060,N_722,N_631);
nand U6061 (N_6061,N_1114,N_2296);
xor U6062 (N_6062,N_3152,N_2749);
nand U6063 (N_6063,N_2870,N_2047);
nand U6064 (N_6064,N_3949,N_1927);
or U6065 (N_6065,N_807,N_1447);
xnor U6066 (N_6066,N_910,N_195);
xnor U6067 (N_6067,N_2079,N_2284);
and U6068 (N_6068,N_1074,N_3900);
nor U6069 (N_6069,N_1649,N_457);
or U6070 (N_6070,N_2956,N_1524);
and U6071 (N_6071,N_3652,N_817);
nor U6072 (N_6072,N_1322,N_436);
and U6073 (N_6073,N_2174,N_1818);
and U6074 (N_6074,N_3277,N_2836);
nand U6075 (N_6075,N_1785,N_685);
nand U6076 (N_6076,N_2967,N_552);
xor U6077 (N_6077,N_3857,N_2473);
or U6078 (N_6078,N_223,N_3898);
nand U6079 (N_6079,N_651,N_1553);
nand U6080 (N_6080,N_721,N_3676);
or U6081 (N_6081,N_1836,N_928);
or U6082 (N_6082,N_177,N_678);
or U6083 (N_6083,N_389,N_820);
and U6084 (N_6084,N_3061,N_2511);
and U6085 (N_6085,N_656,N_2980);
nor U6086 (N_6086,N_1063,N_2561);
nor U6087 (N_6087,N_694,N_2850);
or U6088 (N_6088,N_2691,N_2515);
and U6089 (N_6089,N_2668,N_3391);
xor U6090 (N_6090,N_2014,N_2362);
nand U6091 (N_6091,N_3470,N_362);
or U6092 (N_6092,N_439,N_3863);
and U6093 (N_6093,N_1652,N_2585);
nor U6094 (N_6094,N_941,N_3324);
nor U6095 (N_6095,N_2871,N_2457);
nand U6096 (N_6096,N_3077,N_3862);
or U6097 (N_6097,N_1279,N_1209);
xnor U6098 (N_6098,N_1137,N_996);
and U6099 (N_6099,N_1915,N_3506);
and U6100 (N_6100,N_3568,N_2292);
nand U6101 (N_6101,N_1418,N_960);
nor U6102 (N_6102,N_2122,N_1465);
and U6103 (N_6103,N_300,N_1053);
nor U6104 (N_6104,N_1681,N_696);
and U6105 (N_6105,N_524,N_537);
or U6106 (N_6106,N_3003,N_1655);
nor U6107 (N_6107,N_3608,N_1332);
and U6108 (N_6108,N_3067,N_3470);
nor U6109 (N_6109,N_1663,N_2117);
or U6110 (N_6110,N_69,N_297);
and U6111 (N_6111,N_3826,N_2305);
or U6112 (N_6112,N_463,N_2722);
or U6113 (N_6113,N_3311,N_911);
nor U6114 (N_6114,N_2735,N_121);
nor U6115 (N_6115,N_241,N_922);
or U6116 (N_6116,N_2744,N_3599);
nor U6117 (N_6117,N_732,N_3428);
nand U6118 (N_6118,N_2533,N_555);
or U6119 (N_6119,N_630,N_2610);
nor U6120 (N_6120,N_1917,N_3237);
and U6121 (N_6121,N_2364,N_3807);
nor U6122 (N_6122,N_2183,N_3567);
or U6123 (N_6123,N_411,N_2696);
and U6124 (N_6124,N_1115,N_3537);
nand U6125 (N_6125,N_767,N_3733);
nor U6126 (N_6126,N_51,N_626);
xnor U6127 (N_6127,N_580,N_3451);
and U6128 (N_6128,N_346,N_352);
xor U6129 (N_6129,N_704,N_84);
nand U6130 (N_6130,N_458,N_2660);
xnor U6131 (N_6131,N_287,N_1187);
and U6132 (N_6132,N_2618,N_1309);
and U6133 (N_6133,N_111,N_2463);
or U6134 (N_6134,N_1648,N_457);
and U6135 (N_6135,N_1003,N_1062);
nand U6136 (N_6136,N_3843,N_1231);
nor U6137 (N_6137,N_1164,N_1012);
or U6138 (N_6138,N_2318,N_3671);
nand U6139 (N_6139,N_1868,N_813);
or U6140 (N_6140,N_3321,N_2179);
nand U6141 (N_6141,N_3094,N_2698);
nand U6142 (N_6142,N_1646,N_2455);
xor U6143 (N_6143,N_3031,N_1032);
nand U6144 (N_6144,N_3884,N_2710);
or U6145 (N_6145,N_2552,N_3249);
and U6146 (N_6146,N_48,N_2096);
xnor U6147 (N_6147,N_1344,N_1631);
and U6148 (N_6148,N_723,N_1775);
nor U6149 (N_6149,N_2943,N_2735);
nand U6150 (N_6150,N_3109,N_2993);
and U6151 (N_6151,N_3835,N_177);
or U6152 (N_6152,N_633,N_2634);
and U6153 (N_6153,N_1813,N_697);
nor U6154 (N_6154,N_2924,N_191);
and U6155 (N_6155,N_1614,N_2624);
or U6156 (N_6156,N_2199,N_2923);
nor U6157 (N_6157,N_520,N_3232);
or U6158 (N_6158,N_1727,N_1853);
nor U6159 (N_6159,N_2027,N_3685);
or U6160 (N_6160,N_2574,N_1756);
nand U6161 (N_6161,N_3553,N_3641);
and U6162 (N_6162,N_306,N_2557);
nand U6163 (N_6163,N_2411,N_914);
nor U6164 (N_6164,N_236,N_3940);
nand U6165 (N_6165,N_1894,N_3328);
or U6166 (N_6166,N_3665,N_408);
and U6167 (N_6167,N_2481,N_3320);
xnor U6168 (N_6168,N_1589,N_396);
or U6169 (N_6169,N_1198,N_1804);
and U6170 (N_6170,N_1262,N_1249);
nand U6171 (N_6171,N_896,N_2310);
nand U6172 (N_6172,N_3093,N_3922);
and U6173 (N_6173,N_3571,N_1110);
nor U6174 (N_6174,N_176,N_1504);
nor U6175 (N_6175,N_1813,N_789);
and U6176 (N_6176,N_3500,N_785);
or U6177 (N_6177,N_2428,N_3598);
and U6178 (N_6178,N_1188,N_3724);
nand U6179 (N_6179,N_1464,N_672);
and U6180 (N_6180,N_3015,N_3313);
or U6181 (N_6181,N_1903,N_1959);
or U6182 (N_6182,N_2944,N_3095);
nand U6183 (N_6183,N_3135,N_2980);
or U6184 (N_6184,N_3616,N_993);
xnor U6185 (N_6185,N_635,N_3138);
or U6186 (N_6186,N_1686,N_1696);
and U6187 (N_6187,N_2392,N_2662);
nand U6188 (N_6188,N_611,N_1257);
and U6189 (N_6189,N_621,N_138);
xor U6190 (N_6190,N_333,N_1165);
nor U6191 (N_6191,N_3936,N_864);
nand U6192 (N_6192,N_3390,N_2859);
nor U6193 (N_6193,N_2065,N_2186);
nor U6194 (N_6194,N_2042,N_2198);
nor U6195 (N_6195,N_3271,N_3074);
or U6196 (N_6196,N_2368,N_2042);
nand U6197 (N_6197,N_1520,N_1127);
nor U6198 (N_6198,N_2355,N_3705);
nor U6199 (N_6199,N_1100,N_3743);
xor U6200 (N_6200,N_3027,N_2594);
and U6201 (N_6201,N_2459,N_770);
or U6202 (N_6202,N_1735,N_442);
nand U6203 (N_6203,N_3201,N_1779);
nor U6204 (N_6204,N_1658,N_3484);
nor U6205 (N_6205,N_1057,N_543);
or U6206 (N_6206,N_3509,N_1847);
or U6207 (N_6207,N_3999,N_3325);
and U6208 (N_6208,N_2853,N_713);
nor U6209 (N_6209,N_1269,N_2378);
or U6210 (N_6210,N_662,N_929);
and U6211 (N_6211,N_1283,N_3460);
nor U6212 (N_6212,N_2418,N_3853);
nor U6213 (N_6213,N_1054,N_3602);
nor U6214 (N_6214,N_3098,N_2758);
or U6215 (N_6215,N_2458,N_1751);
and U6216 (N_6216,N_2481,N_590);
or U6217 (N_6217,N_1799,N_453);
nor U6218 (N_6218,N_665,N_1815);
nor U6219 (N_6219,N_3993,N_1960);
nor U6220 (N_6220,N_2418,N_1528);
xnor U6221 (N_6221,N_2079,N_691);
xor U6222 (N_6222,N_766,N_416);
nor U6223 (N_6223,N_2566,N_1229);
and U6224 (N_6224,N_1895,N_1200);
or U6225 (N_6225,N_512,N_1198);
xor U6226 (N_6226,N_1914,N_2520);
nand U6227 (N_6227,N_2480,N_834);
or U6228 (N_6228,N_2322,N_1673);
or U6229 (N_6229,N_3055,N_1716);
xnor U6230 (N_6230,N_2275,N_777);
nand U6231 (N_6231,N_3843,N_2848);
or U6232 (N_6232,N_2062,N_1138);
and U6233 (N_6233,N_2626,N_1319);
nor U6234 (N_6234,N_3420,N_2789);
or U6235 (N_6235,N_2722,N_3171);
nor U6236 (N_6236,N_158,N_405);
xnor U6237 (N_6237,N_2035,N_260);
and U6238 (N_6238,N_2234,N_1049);
and U6239 (N_6239,N_1827,N_1703);
or U6240 (N_6240,N_569,N_2751);
or U6241 (N_6241,N_1036,N_2216);
nand U6242 (N_6242,N_3539,N_3287);
nor U6243 (N_6243,N_937,N_1848);
nor U6244 (N_6244,N_2169,N_3262);
nor U6245 (N_6245,N_1543,N_2315);
or U6246 (N_6246,N_2928,N_68);
and U6247 (N_6247,N_3434,N_2376);
and U6248 (N_6248,N_1962,N_1058);
nor U6249 (N_6249,N_1422,N_67);
nand U6250 (N_6250,N_1876,N_3816);
and U6251 (N_6251,N_2211,N_1637);
or U6252 (N_6252,N_2165,N_254);
or U6253 (N_6253,N_3545,N_38);
or U6254 (N_6254,N_524,N_3319);
or U6255 (N_6255,N_1209,N_2737);
or U6256 (N_6256,N_1443,N_3690);
xnor U6257 (N_6257,N_1616,N_6);
nor U6258 (N_6258,N_3565,N_1864);
or U6259 (N_6259,N_2116,N_817);
and U6260 (N_6260,N_1055,N_1083);
and U6261 (N_6261,N_970,N_2082);
and U6262 (N_6262,N_3981,N_3967);
and U6263 (N_6263,N_3541,N_3756);
nand U6264 (N_6264,N_2940,N_2923);
nor U6265 (N_6265,N_2090,N_2713);
nand U6266 (N_6266,N_3471,N_1046);
or U6267 (N_6267,N_749,N_629);
nor U6268 (N_6268,N_3545,N_506);
and U6269 (N_6269,N_1611,N_684);
and U6270 (N_6270,N_2685,N_2606);
nor U6271 (N_6271,N_86,N_2500);
nor U6272 (N_6272,N_3504,N_2049);
or U6273 (N_6273,N_3527,N_1607);
or U6274 (N_6274,N_762,N_3599);
or U6275 (N_6275,N_2289,N_2944);
xor U6276 (N_6276,N_1899,N_2592);
or U6277 (N_6277,N_279,N_1662);
nand U6278 (N_6278,N_3040,N_3580);
and U6279 (N_6279,N_1188,N_1457);
xor U6280 (N_6280,N_3539,N_3006);
or U6281 (N_6281,N_3471,N_868);
and U6282 (N_6282,N_1695,N_2136);
xnor U6283 (N_6283,N_3117,N_1203);
or U6284 (N_6284,N_693,N_919);
nor U6285 (N_6285,N_2461,N_3739);
nand U6286 (N_6286,N_1161,N_542);
or U6287 (N_6287,N_309,N_3088);
or U6288 (N_6288,N_200,N_1360);
xor U6289 (N_6289,N_730,N_259);
nor U6290 (N_6290,N_3889,N_3634);
nand U6291 (N_6291,N_3718,N_2259);
and U6292 (N_6292,N_600,N_2927);
or U6293 (N_6293,N_3312,N_1775);
and U6294 (N_6294,N_2580,N_1100);
or U6295 (N_6295,N_1725,N_1761);
nand U6296 (N_6296,N_565,N_3850);
or U6297 (N_6297,N_2829,N_3418);
or U6298 (N_6298,N_1468,N_1945);
nand U6299 (N_6299,N_2035,N_3906);
and U6300 (N_6300,N_1632,N_3959);
nand U6301 (N_6301,N_1950,N_2581);
or U6302 (N_6302,N_2940,N_1785);
xnor U6303 (N_6303,N_556,N_1468);
nand U6304 (N_6304,N_1258,N_446);
or U6305 (N_6305,N_2675,N_3434);
and U6306 (N_6306,N_2831,N_2745);
and U6307 (N_6307,N_1380,N_3426);
and U6308 (N_6308,N_2030,N_3375);
and U6309 (N_6309,N_1103,N_3027);
xnor U6310 (N_6310,N_2399,N_2829);
nor U6311 (N_6311,N_2564,N_3380);
nand U6312 (N_6312,N_241,N_2997);
nor U6313 (N_6313,N_343,N_943);
and U6314 (N_6314,N_1609,N_166);
nor U6315 (N_6315,N_1899,N_879);
or U6316 (N_6316,N_3716,N_3837);
or U6317 (N_6317,N_1987,N_969);
and U6318 (N_6318,N_1007,N_3416);
nand U6319 (N_6319,N_2505,N_3356);
and U6320 (N_6320,N_3697,N_2021);
nand U6321 (N_6321,N_3336,N_2313);
and U6322 (N_6322,N_750,N_2288);
or U6323 (N_6323,N_1682,N_370);
and U6324 (N_6324,N_799,N_27);
and U6325 (N_6325,N_3573,N_3758);
nand U6326 (N_6326,N_439,N_3786);
nand U6327 (N_6327,N_3673,N_3217);
nor U6328 (N_6328,N_1363,N_2374);
and U6329 (N_6329,N_1886,N_124);
and U6330 (N_6330,N_3712,N_270);
nand U6331 (N_6331,N_629,N_2914);
nor U6332 (N_6332,N_3138,N_2535);
or U6333 (N_6333,N_3177,N_575);
and U6334 (N_6334,N_2296,N_2881);
and U6335 (N_6335,N_1838,N_871);
nand U6336 (N_6336,N_1198,N_2418);
nor U6337 (N_6337,N_18,N_1020);
xnor U6338 (N_6338,N_2783,N_2460);
and U6339 (N_6339,N_1221,N_2747);
and U6340 (N_6340,N_3,N_31);
nor U6341 (N_6341,N_2252,N_1704);
and U6342 (N_6342,N_3989,N_1986);
and U6343 (N_6343,N_310,N_670);
nand U6344 (N_6344,N_1678,N_975);
or U6345 (N_6345,N_2324,N_820);
nor U6346 (N_6346,N_2791,N_1542);
and U6347 (N_6347,N_2388,N_3232);
nor U6348 (N_6348,N_3862,N_2355);
xor U6349 (N_6349,N_1208,N_2054);
xor U6350 (N_6350,N_3062,N_1303);
and U6351 (N_6351,N_2907,N_1040);
nor U6352 (N_6352,N_492,N_3311);
nand U6353 (N_6353,N_3153,N_1231);
or U6354 (N_6354,N_143,N_2291);
and U6355 (N_6355,N_3448,N_3890);
and U6356 (N_6356,N_3047,N_1535);
or U6357 (N_6357,N_3823,N_2431);
nor U6358 (N_6358,N_3717,N_2912);
nand U6359 (N_6359,N_1162,N_2225);
nor U6360 (N_6360,N_2600,N_2011);
or U6361 (N_6361,N_445,N_2140);
nand U6362 (N_6362,N_121,N_766);
or U6363 (N_6363,N_3021,N_1258);
nor U6364 (N_6364,N_1193,N_183);
or U6365 (N_6365,N_1021,N_2376);
or U6366 (N_6366,N_588,N_862);
and U6367 (N_6367,N_2650,N_186);
or U6368 (N_6368,N_192,N_1688);
and U6369 (N_6369,N_293,N_2161);
nor U6370 (N_6370,N_3568,N_369);
nor U6371 (N_6371,N_1164,N_443);
or U6372 (N_6372,N_2714,N_1518);
or U6373 (N_6373,N_1918,N_2202);
nor U6374 (N_6374,N_3175,N_2177);
xnor U6375 (N_6375,N_2710,N_2870);
and U6376 (N_6376,N_1015,N_646);
nor U6377 (N_6377,N_1067,N_2610);
and U6378 (N_6378,N_1167,N_3400);
and U6379 (N_6379,N_199,N_3565);
xnor U6380 (N_6380,N_3221,N_3932);
xor U6381 (N_6381,N_2329,N_85);
xor U6382 (N_6382,N_2811,N_2600);
or U6383 (N_6383,N_571,N_2287);
nand U6384 (N_6384,N_1920,N_1632);
and U6385 (N_6385,N_2755,N_2002);
and U6386 (N_6386,N_337,N_3898);
nor U6387 (N_6387,N_2342,N_1280);
nor U6388 (N_6388,N_2206,N_3414);
and U6389 (N_6389,N_3094,N_3596);
or U6390 (N_6390,N_3133,N_3723);
nand U6391 (N_6391,N_3084,N_2975);
or U6392 (N_6392,N_1881,N_2185);
nor U6393 (N_6393,N_490,N_749);
nor U6394 (N_6394,N_1327,N_1139);
and U6395 (N_6395,N_3376,N_540);
or U6396 (N_6396,N_1527,N_2592);
nor U6397 (N_6397,N_3404,N_3562);
or U6398 (N_6398,N_1854,N_537);
or U6399 (N_6399,N_1652,N_822);
nand U6400 (N_6400,N_1206,N_1135);
nor U6401 (N_6401,N_2338,N_3423);
nand U6402 (N_6402,N_2376,N_3562);
nand U6403 (N_6403,N_2509,N_2846);
and U6404 (N_6404,N_1715,N_2026);
or U6405 (N_6405,N_839,N_1728);
nand U6406 (N_6406,N_3893,N_3787);
nor U6407 (N_6407,N_3259,N_3830);
nor U6408 (N_6408,N_3262,N_1522);
or U6409 (N_6409,N_1419,N_2250);
and U6410 (N_6410,N_3769,N_2556);
nand U6411 (N_6411,N_2594,N_240);
nor U6412 (N_6412,N_3994,N_433);
or U6413 (N_6413,N_3946,N_1350);
nand U6414 (N_6414,N_2859,N_3670);
and U6415 (N_6415,N_3410,N_277);
xor U6416 (N_6416,N_2144,N_3066);
and U6417 (N_6417,N_3075,N_3101);
xnor U6418 (N_6418,N_1030,N_2354);
and U6419 (N_6419,N_2066,N_3728);
and U6420 (N_6420,N_2533,N_1007);
or U6421 (N_6421,N_3479,N_2740);
or U6422 (N_6422,N_1335,N_2043);
and U6423 (N_6423,N_294,N_2773);
nor U6424 (N_6424,N_2663,N_284);
and U6425 (N_6425,N_3102,N_2320);
nand U6426 (N_6426,N_3952,N_3420);
and U6427 (N_6427,N_2279,N_1382);
nand U6428 (N_6428,N_3354,N_3939);
or U6429 (N_6429,N_1672,N_1210);
or U6430 (N_6430,N_1578,N_611);
and U6431 (N_6431,N_186,N_3458);
or U6432 (N_6432,N_897,N_652);
or U6433 (N_6433,N_1545,N_2249);
nor U6434 (N_6434,N_2439,N_2610);
or U6435 (N_6435,N_110,N_3161);
and U6436 (N_6436,N_2596,N_3556);
nand U6437 (N_6437,N_552,N_252);
or U6438 (N_6438,N_177,N_3426);
and U6439 (N_6439,N_3909,N_3618);
nor U6440 (N_6440,N_1824,N_1415);
nand U6441 (N_6441,N_812,N_2797);
and U6442 (N_6442,N_1276,N_2078);
or U6443 (N_6443,N_3349,N_1075);
nand U6444 (N_6444,N_3678,N_1523);
or U6445 (N_6445,N_1664,N_58);
nand U6446 (N_6446,N_66,N_578);
and U6447 (N_6447,N_1058,N_3429);
nor U6448 (N_6448,N_77,N_2450);
xor U6449 (N_6449,N_3594,N_3063);
and U6450 (N_6450,N_2182,N_457);
and U6451 (N_6451,N_2221,N_661);
and U6452 (N_6452,N_2675,N_536);
xnor U6453 (N_6453,N_1600,N_1184);
nand U6454 (N_6454,N_1155,N_3489);
nand U6455 (N_6455,N_665,N_2618);
nand U6456 (N_6456,N_3132,N_2521);
and U6457 (N_6457,N_2738,N_2307);
and U6458 (N_6458,N_3836,N_3628);
nor U6459 (N_6459,N_3093,N_3554);
nor U6460 (N_6460,N_3789,N_3947);
nor U6461 (N_6461,N_3850,N_2649);
nand U6462 (N_6462,N_565,N_3393);
nor U6463 (N_6463,N_3822,N_1255);
and U6464 (N_6464,N_3419,N_2067);
nor U6465 (N_6465,N_2135,N_2782);
or U6466 (N_6466,N_557,N_3004);
nor U6467 (N_6467,N_869,N_2420);
and U6468 (N_6468,N_1449,N_3449);
nand U6469 (N_6469,N_1203,N_239);
nor U6470 (N_6470,N_558,N_2796);
nor U6471 (N_6471,N_1834,N_3469);
or U6472 (N_6472,N_1899,N_3600);
xor U6473 (N_6473,N_2768,N_1455);
and U6474 (N_6474,N_1971,N_949);
xnor U6475 (N_6475,N_3756,N_3278);
nand U6476 (N_6476,N_982,N_1094);
nor U6477 (N_6477,N_1501,N_3333);
nand U6478 (N_6478,N_2604,N_1030);
nor U6479 (N_6479,N_2972,N_3937);
or U6480 (N_6480,N_2073,N_3591);
or U6481 (N_6481,N_1019,N_3020);
xor U6482 (N_6482,N_2469,N_1553);
nor U6483 (N_6483,N_419,N_2628);
or U6484 (N_6484,N_3036,N_1683);
nor U6485 (N_6485,N_1045,N_224);
nand U6486 (N_6486,N_1208,N_1175);
nand U6487 (N_6487,N_3472,N_2649);
nand U6488 (N_6488,N_199,N_555);
and U6489 (N_6489,N_1031,N_891);
xor U6490 (N_6490,N_3651,N_2274);
nand U6491 (N_6491,N_3888,N_3853);
or U6492 (N_6492,N_3560,N_1763);
or U6493 (N_6493,N_1220,N_176);
nand U6494 (N_6494,N_3687,N_3505);
xnor U6495 (N_6495,N_1184,N_1890);
nor U6496 (N_6496,N_1301,N_2923);
and U6497 (N_6497,N_708,N_3667);
or U6498 (N_6498,N_3296,N_3616);
nor U6499 (N_6499,N_2843,N_2059);
and U6500 (N_6500,N_90,N_2215);
nand U6501 (N_6501,N_418,N_533);
and U6502 (N_6502,N_2579,N_2792);
nor U6503 (N_6503,N_2472,N_1853);
or U6504 (N_6504,N_688,N_2506);
nor U6505 (N_6505,N_504,N_3174);
nor U6506 (N_6506,N_3865,N_3014);
or U6507 (N_6507,N_1439,N_2412);
nand U6508 (N_6508,N_3735,N_2445);
xnor U6509 (N_6509,N_1922,N_2056);
nor U6510 (N_6510,N_3689,N_1802);
and U6511 (N_6511,N_3341,N_2522);
nand U6512 (N_6512,N_2401,N_138);
and U6513 (N_6513,N_553,N_1821);
nor U6514 (N_6514,N_108,N_3927);
or U6515 (N_6515,N_1356,N_372);
nor U6516 (N_6516,N_189,N_1089);
nor U6517 (N_6517,N_1990,N_1853);
and U6518 (N_6518,N_533,N_967);
or U6519 (N_6519,N_652,N_1456);
nand U6520 (N_6520,N_2668,N_2223);
nand U6521 (N_6521,N_47,N_1788);
or U6522 (N_6522,N_2092,N_1020);
nor U6523 (N_6523,N_2544,N_3148);
or U6524 (N_6524,N_3125,N_126);
nor U6525 (N_6525,N_3361,N_3534);
and U6526 (N_6526,N_125,N_115);
and U6527 (N_6527,N_3130,N_2211);
nor U6528 (N_6528,N_262,N_2092);
nand U6529 (N_6529,N_40,N_1706);
nor U6530 (N_6530,N_1861,N_997);
xor U6531 (N_6531,N_2677,N_1416);
and U6532 (N_6532,N_3812,N_520);
and U6533 (N_6533,N_2010,N_1991);
xnor U6534 (N_6534,N_3215,N_154);
and U6535 (N_6535,N_3517,N_1977);
nor U6536 (N_6536,N_2724,N_1045);
or U6537 (N_6537,N_3061,N_1276);
nor U6538 (N_6538,N_2448,N_2643);
xor U6539 (N_6539,N_1182,N_1528);
nand U6540 (N_6540,N_3117,N_470);
nand U6541 (N_6541,N_786,N_3258);
or U6542 (N_6542,N_872,N_694);
nor U6543 (N_6543,N_353,N_636);
and U6544 (N_6544,N_1501,N_1704);
nand U6545 (N_6545,N_2712,N_2556);
nand U6546 (N_6546,N_605,N_1133);
and U6547 (N_6547,N_3525,N_1808);
or U6548 (N_6548,N_3134,N_347);
nand U6549 (N_6549,N_3795,N_2675);
nor U6550 (N_6550,N_1534,N_2864);
nand U6551 (N_6551,N_3846,N_2278);
nor U6552 (N_6552,N_2137,N_620);
or U6553 (N_6553,N_992,N_619);
or U6554 (N_6554,N_688,N_3768);
nand U6555 (N_6555,N_2389,N_966);
and U6556 (N_6556,N_3435,N_2130);
nor U6557 (N_6557,N_3069,N_471);
nand U6558 (N_6558,N_692,N_1814);
nor U6559 (N_6559,N_712,N_2863);
nor U6560 (N_6560,N_2865,N_2827);
and U6561 (N_6561,N_1442,N_56);
nand U6562 (N_6562,N_1281,N_3632);
or U6563 (N_6563,N_2410,N_1849);
nor U6564 (N_6564,N_2156,N_250);
nand U6565 (N_6565,N_2757,N_2573);
and U6566 (N_6566,N_3881,N_2341);
nand U6567 (N_6567,N_3343,N_138);
nor U6568 (N_6568,N_1310,N_2050);
nor U6569 (N_6569,N_2061,N_1271);
xor U6570 (N_6570,N_1271,N_3535);
nand U6571 (N_6571,N_1407,N_154);
nand U6572 (N_6572,N_1801,N_1966);
and U6573 (N_6573,N_2201,N_288);
nor U6574 (N_6574,N_1899,N_3378);
and U6575 (N_6575,N_2848,N_1601);
or U6576 (N_6576,N_311,N_3868);
or U6577 (N_6577,N_387,N_1446);
nand U6578 (N_6578,N_2365,N_1312);
or U6579 (N_6579,N_459,N_3930);
and U6580 (N_6580,N_3701,N_757);
and U6581 (N_6581,N_3770,N_1549);
nand U6582 (N_6582,N_3925,N_3173);
or U6583 (N_6583,N_1648,N_565);
nor U6584 (N_6584,N_1387,N_135);
or U6585 (N_6585,N_577,N_178);
nor U6586 (N_6586,N_1144,N_1197);
nor U6587 (N_6587,N_1408,N_379);
nor U6588 (N_6588,N_2747,N_1640);
nand U6589 (N_6589,N_3927,N_469);
nor U6590 (N_6590,N_3747,N_861);
nor U6591 (N_6591,N_651,N_1887);
nor U6592 (N_6592,N_1941,N_3931);
or U6593 (N_6593,N_3901,N_3538);
and U6594 (N_6594,N_2207,N_1857);
nor U6595 (N_6595,N_2574,N_3485);
nor U6596 (N_6596,N_3820,N_2114);
and U6597 (N_6597,N_401,N_1629);
nor U6598 (N_6598,N_1164,N_1047);
nor U6599 (N_6599,N_3272,N_3729);
xor U6600 (N_6600,N_1369,N_3464);
nand U6601 (N_6601,N_2045,N_385);
or U6602 (N_6602,N_412,N_3162);
and U6603 (N_6603,N_3661,N_1525);
and U6604 (N_6604,N_398,N_1806);
nor U6605 (N_6605,N_2918,N_1558);
xor U6606 (N_6606,N_3468,N_1412);
nand U6607 (N_6607,N_2448,N_695);
and U6608 (N_6608,N_3545,N_3622);
nand U6609 (N_6609,N_2681,N_1387);
and U6610 (N_6610,N_3930,N_2111);
nand U6611 (N_6611,N_3251,N_423);
or U6612 (N_6612,N_1268,N_1607);
and U6613 (N_6613,N_1941,N_610);
and U6614 (N_6614,N_3237,N_2129);
or U6615 (N_6615,N_3260,N_1303);
or U6616 (N_6616,N_1314,N_790);
or U6617 (N_6617,N_652,N_2171);
and U6618 (N_6618,N_918,N_3886);
or U6619 (N_6619,N_1040,N_2717);
xor U6620 (N_6620,N_483,N_2094);
nand U6621 (N_6621,N_232,N_3444);
xnor U6622 (N_6622,N_2892,N_2543);
nor U6623 (N_6623,N_870,N_3168);
or U6624 (N_6624,N_2607,N_2688);
and U6625 (N_6625,N_3915,N_340);
nor U6626 (N_6626,N_1549,N_588);
or U6627 (N_6627,N_1718,N_3675);
nor U6628 (N_6628,N_1305,N_1169);
xor U6629 (N_6629,N_316,N_2618);
nor U6630 (N_6630,N_1697,N_1262);
or U6631 (N_6631,N_1956,N_934);
xor U6632 (N_6632,N_2167,N_2481);
or U6633 (N_6633,N_1078,N_1638);
xnor U6634 (N_6634,N_2951,N_3616);
nor U6635 (N_6635,N_1769,N_3411);
nor U6636 (N_6636,N_1660,N_2079);
nand U6637 (N_6637,N_3243,N_872);
or U6638 (N_6638,N_2890,N_307);
nor U6639 (N_6639,N_2980,N_1474);
xnor U6640 (N_6640,N_3462,N_1048);
or U6641 (N_6641,N_886,N_818);
xnor U6642 (N_6642,N_3349,N_2891);
nor U6643 (N_6643,N_3794,N_2557);
nand U6644 (N_6644,N_2093,N_3668);
and U6645 (N_6645,N_263,N_18);
nand U6646 (N_6646,N_303,N_3871);
nor U6647 (N_6647,N_1195,N_2390);
or U6648 (N_6648,N_3016,N_2125);
nand U6649 (N_6649,N_3584,N_1026);
and U6650 (N_6650,N_1826,N_3350);
or U6651 (N_6651,N_1437,N_3530);
nor U6652 (N_6652,N_3193,N_357);
or U6653 (N_6653,N_850,N_2101);
and U6654 (N_6654,N_2547,N_2544);
nand U6655 (N_6655,N_3308,N_594);
and U6656 (N_6656,N_3265,N_203);
xnor U6657 (N_6657,N_1837,N_1896);
and U6658 (N_6658,N_625,N_404);
nor U6659 (N_6659,N_1149,N_139);
nand U6660 (N_6660,N_3488,N_2702);
and U6661 (N_6661,N_2006,N_1742);
nor U6662 (N_6662,N_2103,N_1682);
xor U6663 (N_6663,N_2376,N_263);
nand U6664 (N_6664,N_961,N_2141);
or U6665 (N_6665,N_3720,N_532);
nor U6666 (N_6666,N_3759,N_2484);
nand U6667 (N_6667,N_2377,N_70);
or U6668 (N_6668,N_3083,N_560);
and U6669 (N_6669,N_3259,N_2496);
or U6670 (N_6670,N_1728,N_1872);
nand U6671 (N_6671,N_3397,N_117);
nand U6672 (N_6672,N_1591,N_187);
nand U6673 (N_6673,N_2682,N_349);
nand U6674 (N_6674,N_2686,N_3105);
nand U6675 (N_6675,N_2210,N_1675);
and U6676 (N_6676,N_3655,N_1562);
nand U6677 (N_6677,N_2721,N_2529);
or U6678 (N_6678,N_3242,N_3347);
and U6679 (N_6679,N_2109,N_124);
nor U6680 (N_6680,N_350,N_2557);
or U6681 (N_6681,N_2566,N_485);
and U6682 (N_6682,N_1862,N_3378);
or U6683 (N_6683,N_195,N_1153);
xnor U6684 (N_6684,N_1138,N_2898);
nor U6685 (N_6685,N_3324,N_3692);
nor U6686 (N_6686,N_2299,N_756);
and U6687 (N_6687,N_2592,N_1776);
nand U6688 (N_6688,N_617,N_808);
xor U6689 (N_6689,N_811,N_2885);
nand U6690 (N_6690,N_1827,N_865);
or U6691 (N_6691,N_3373,N_1953);
and U6692 (N_6692,N_1343,N_1996);
and U6693 (N_6693,N_3739,N_345);
nor U6694 (N_6694,N_1142,N_542);
nand U6695 (N_6695,N_1427,N_2055);
or U6696 (N_6696,N_3101,N_2162);
and U6697 (N_6697,N_1360,N_845);
nand U6698 (N_6698,N_1663,N_3593);
nand U6699 (N_6699,N_2602,N_1481);
xor U6700 (N_6700,N_2317,N_279);
nor U6701 (N_6701,N_83,N_1872);
nor U6702 (N_6702,N_2256,N_1337);
or U6703 (N_6703,N_183,N_3668);
and U6704 (N_6704,N_2901,N_1795);
or U6705 (N_6705,N_979,N_834);
or U6706 (N_6706,N_1829,N_1062);
nor U6707 (N_6707,N_1408,N_3138);
nand U6708 (N_6708,N_3009,N_1488);
nor U6709 (N_6709,N_3831,N_1899);
nand U6710 (N_6710,N_2226,N_877);
nand U6711 (N_6711,N_2801,N_392);
or U6712 (N_6712,N_3491,N_2291);
xnor U6713 (N_6713,N_1642,N_927);
or U6714 (N_6714,N_1333,N_473);
nand U6715 (N_6715,N_1280,N_1270);
xnor U6716 (N_6716,N_910,N_3110);
nand U6717 (N_6717,N_2478,N_916);
or U6718 (N_6718,N_2984,N_2714);
nor U6719 (N_6719,N_1828,N_584);
nor U6720 (N_6720,N_1177,N_914);
nor U6721 (N_6721,N_529,N_3199);
and U6722 (N_6722,N_909,N_743);
nor U6723 (N_6723,N_486,N_3105);
nor U6724 (N_6724,N_1489,N_35);
nor U6725 (N_6725,N_2831,N_734);
nor U6726 (N_6726,N_2974,N_3252);
or U6727 (N_6727,N_3359,N_699);
or U6728 (N_6728,N_327,N_1030);
nand U6729 (N_6729,N_3935,N_3356);
and U6730 (N_6730,N_1956,N_2314);
nor U6731 (N_6731,N_2807,N_899);
or U6732 (N_6732,N_1853,N_3508);
xnor U6733 (N_6733,N_1478,N_172);
nor U6734 (N_6734,N_816,N_1372);
nor U6735 (N_6735,N_3346,N_691);
nor U6736 (N_6736,N_60,N_1778);
and U6737 (N_6737,N_2778,N_691);
or U6738 (N_6738,N_1783,N_360);
xor U6739 (N_6739,N_1570,N_2227);
and U6740 (N_6740,N_2826,N_2565);
or U6741 (N_6741,N_2631,N_498);
and U6742 (N_6742,N_2312,N_3484);
nor U6743 (N_6743,N_2204,N_3602);
nand U6744 (N_6744,N_1183,N_3220);
nand U6745 (N_6745,N_3065,N_3357);
nand U6746 (N_6746,N_3194,N_2062);
nand U6747 (N_6747,N_2647,N_2970);
nor U6748 (N_6748,N_1199,N_2598);
or U6749 (N_6749,N_538,N_3422);
nand U6750 (N_6750,N_2822,N_812);
nor U6751 (N_6751,N_846,N_1923);
or U6752 (N_6752,N_539,N_1181);
and U6753 (N_6753,N_1797,N_2660);
nand U6754 (N_6754,N_2288,N_2032);
xor U6755 (N_6755,N_428,N_2682);
nand U6756 (N_6756,N_3930,N_1642);
nor U6757 (N_6757,N_1132,N_104);
or U6758 (N_6758,N_3233,N_783);
or U6759 (N_6759,N_3453,N_1586);
nand U6760 (N_6760,N_292,N_1980);
nand U6761 (N_6761,N_1396,N_3512);
or U6762 (N_6762,N_3380,N_304);
nand U6763 (N_6763,N_970,N_2364);
xor U6764 (N_6764,N_3430,N_2815);
xnor U6765 (N_6765,N_3811,N_3889);
or U6766 (N_6766,N_451,N_838);
xor U6767 (N_6767,N_3939,N_119);
or U6768 (N_6768,N_2277,N_2140);
and U6769 (N_6769,N_1966,N_672);
nor U6770 (N_6770,N_2803,N_450);
or U6771 (N_6771,N_3601,N_2243);
or U6772 (N_6772,N_2196,N_892);
nor U6773 (N_6773,N_1883,N_845);
nand U6774 (N_6774,N_1143,N_2362);
nor U6775 (N_6775,N_2160,N_2549);
nand U6776 (N_6776,N_1704,N_3878);
nand U6777 (N_6777,N_1226,N_2090);
or U6778 (N_6778,N_3403,N_58);
nor U6779 (N_6779,N_2589,N_3469);
or U6780 (N_6780,N_493,N_1572);
or U6781 (N_6781,N_2796,N_1603);
or U6782 (N_6782,N_1253,N_1436);
xnor U6783 (N_6783,N_3404,N_3682);
xnor U6784 (N_6784,N_3621,N_3873);
or U6785 (N_6785,N_2804,N_2311);
nand U6786 (N_6786,N_766,N_480);
nor U6787 (N_6787,N_1212,N_3936);
or U6788 (N_6788,N_3570,N_1030);
nor U6789 (N_6789,N_89,N_139);
and U6790 (N_6790,N_3736,N_3300);
or U6791 (N_6791,N_2291,N_79);
and U6792 (N_6792,N_2994,N_3586);
xnor U6793 (N_6793,N_417,N_179);
nor U6794 (N_6794,N_1767,N_475);
nand U6795 (N_6795,N_1056,N_3294);
or U6796 (N_6796,N_2878,N_3062);
nor U6797 (N_6797,N_951,N_3210);
or U6798 (N_6798,N_3761,N_1677);
nor U6799 (N_6799,N_3325,N_3475);
and U6800 (N_6800,N_3925,N_2313);
nand U6801 (N_6801,N_3241,N_553);
or U6802 (N_6802,N_2196,N_2773);
nor U6803 (N_6803,N_2007,N_3164);
and U6804 (N_6804,N_1104,N_3945);
nor U6805 (N_6805,N_2612,N_121);
and U6806 (N_6806,N_2692,N_3237);
or U6807 (N_6807,N_551,N_270);
and U6808 (N_6808,N_714,N_3391);
nor U6809 (N_6809,N_1848,N_2494);
nor U6810 (N_6810,N_2313,N_3558);
or U6811 (N_6811,N_1536,N_1773);
nand U6812 (N_6812,N_1999,N_876);
or U6813 (N_6813,N_1606,N_1532);
nand U6814 (N_6814,N_3790,N_111);
and U6815 (N_6815,N_2985,N_3236);
nor U6816 (N_6816,N_1942,N_605);
or U6817 (N_6817,N_624,N_330);
and U6818 (N_6818,N_3229,N_2887);
nand U6819 (N_6819,N_1663,N_1080);
and U6820 (N_6820,N_432,N_921);
and U6821 (N_6821,N_428,N_2624);
or U6822 (N_6822,N_2446,N_924);
nor U6823 (N_6823,N_3869,N_674);
nand U6824 (N_6824,N_981,N_380);
nor U6825 (N_6825,N_3904,N_3886);
and U6826 (N_6826,N_1225,N_3494);
nand U6827 (N_6827,N_3002,N_2712);
xor U6828 (N_6828,N_1433,N_2425);
nand U6829 (N_6829,N_2862,N_3718);
xnor U6830 (N_6830,N_2518,N_3960);
xor U6831 (N_6831,N_3288,N_2186);
nand U6832 (N_6832,N_414,N_725);
or U6833 (N_6833,N_1779,N_2994);
and U6834 (N_6834,N_1036,N_2800);
nor U6835 (N_6835,N_273,N_3022);
nor U6836 (N_6836,N_2484,N_3981);
and U6837 (N_6837,N_100,N_421);
or U6838 (N_6838,N_162,N_2627);
or U6839 (N_6839,N_3641,N_1804);
and U6840 (N_6840,N_469,N_3521);
nor U6841 (N_6841,N_125,N_1212);
xor U6842 (N_6842,N_1387,N_3207);
and U6843 (N_6843,N_3577,N_597);
or U6844 (N_6844,N_1388,N_3756);
and U6845 (N_6845,N_3019,N_936);
and U6846 (N_6846,N_2522,N_2478);
nor U6847 (N_6847,N_1573,N_953);
nor U6848 (N_6848,N_2681,N_1781);
or U6849 (N_6849,N_962,N_1052);
nor U6850 (N_6850,N_1181,N_808);
xnor U6851 (N_6851,N_314,N_3219);
nor U6852 (N_6852,N_3740,N_2335);
and U6853 (N_6853,N_1576,N_1442);
nand U6854 (N_6854,N_769,N_2681);
nor U6855 (N_6855,N_3989,N_342);
and U6856 (N_6856,N_831,N_1580);
nand U6857 (N_6857,N_3755,N_1407);
and U6858 (N_6858,N_2405,N_3704);
and U6859 (N_6859,N_3670,N_2140);
xor U6860 (N_6860,N_2254,N_1098);
nor U6861 (N_6861,N_3179,N_2097);
xnor U6862 (N_6862,N_2124,N_3701);
or U6863 (N_6863,N_2652,N_1264);
and U6864 (N_6864,N_1124,N_2539);
and U6865 (N_6865,N_1355,N_2058);
or U6866 (N_6866,N_975,N_3589);
or U6867 (N_6867,N_2490,N_117);
and U6868 (N_6868,N_143,N_15);
nand U6869 (N_6869,N_2375,N_1857);
nand U6870 (N_6870,N_673,N_1699);
or U6871 (N_6871,N_1728,N_374);
nor U6872 (N_6872,N_3640,N_1860);
nand U6873 (N_6873,N_3333,N_2015);
nor U6874 (N_6874,N_2537,N_2488);
or U6875 (N_6875,N_361,N_3583);
nand U6876 (N_6876,N_162,N_1870);
nor U6877 (N_6877,N_1178,N_3055);
nor U6878 (N_6878,N_3465,N_2072);
nor U6879 (N_6879,N_2029,N_3948);
xor U6880 (N_6880,N_3612,N_2401);
nor U6881 (N_6881,N_1980,N_1683);
or U6882 (N_6882,N_3694,N_2501);
nand U6883 (N_6883,N_3107,N_2397);
nor U6884 (N_6884,N_3291,N_1388);
nand U6885 (N_6885,N_3062,N_2897);
or U6886 (N_6886,N_2160,N_1617);
nand U6887 (N_6887,N_644,N_3072);
and U6888 (N_6888,N_2620,N_2110);
nand U6889 (N_6889,N_3867,N_2617);
or U6890 (N_6890,N_2953,N_1832);
and U6891 (N_6891,N_1325,N_338);
and U6892 (N_6892,N_256,N_1958);
and U6893 (N_6893,N_986,N_904);
nor U6894 (N_6894,N_3429,N_158);
or U6895 (N_6895,N_1544,N_1586);
xor U6896 (N_6896,N_2450,N_3791);
xor U6897 (N_6897,N_2253,N_3342);
and U6898 (N_6898,N_3079,N_324);
nand U6899 (N_6899,N_930,N_1986);
nand U6900 (N_6900,N_742,N_2627);
xnor U6901 (N_6901,N_3871,N_3005);
nor U6902 (N_6902,N_1791,N_809);
or U6903 (N_6903,N_3795,N_1512);
or U6904 (N_6904,N_3876,N_3997);
and U6905 (N_6905,N_2,N_2882);
nor U6906 (N_6906,N_1354,N_99);
nor U6907 (N_6907,N_2409,N_3848);
nand U6908 (N_6908,N_2239,N_3375);
or U6909 (N_6909,N_1576,N_1506);
and U6910 (N_6910,N_1304,N_751);
nor U6911 (N_6911,N_901,N_1546);
and U6912 (N_6912,N_3657,N_407);
or U6913 (N_6913,N_2941,N_1519);
xnor U6914 (N_6914,N_936,N_3925);
xor U6915 (N_6915,N_1180,N_1155);
nand U6916 (N_6916,N_2778,N_557);
xor U6917 (N_6917,N_1687,N_2576);
or U6918 (N_6918,N_967,N_131);
nand U6919 (N_6919,N_3844,N_230);
or U6920 (N_6920,N_1053,N_1435);
nor U6921 (N_6921,N_920,N_464);
nor U6922 (N_6922,N_2010,N_2122);
and U6923 (N_6923,N_807,N_1688);
nor U6924 (N_6924,N_2353,N_1792);
or U6925 (N_6925,N_3197,N_1237);
nand U6926 (N_6926,N_3527,N_189);
or U6927 (N_6927,N_2833,N_2747);
and U6928 (N_6928,N_2530,N_3298);
or U6929 (N_6929,N_830,N_2937);
nand U6930 (N_6930,N_917,N_2273);
xor U6931 (N_6931,N_423,N_2848);
xor U6932 (N_6932,N_2725,N_2463);
and U6933 (N_6933,N_2711,N_548);
nand U6934 (N_6934,N_1358,N_2017);
nand U6935 (N_6935,N_1523,N_358);
nor U6936 (N_6936,N_3807,N_889);
nor U6937 (N_6937,N_785,N_2422);
nand U6938 (N_6938,N_1715,N_949);
nor U6939 (N_6939,N_3240,N_444);
and U6940 (N_6940,N_2043,N_1226);
or U6941 (N_6941,N_1439,N_1072);
nor U6942 (N_6942,N_2664,N_1827);
and U6943 (N_6943,N_3540,N_3674);
nand U6944 (N_6944,N_1159,N_35);
or U6945 (N_6945,N_2220,N_3943);
nand U6946 (N_6946,N_2750,N_680);
and U6947 (N_6947,N_2817,N_2985);
nand U6948 (N_6948,N_2624,N_817);
and U6949 (N_6949,N_3435,N_2117);
nand U6950 (N_6950,N_774,N_2273);
nand U6951 (N_6951,N_777,N_1901);
nor U6952 (N_6952,N_3637,N_813);
and U6953 (N_6953,N_1451,N_1310);
and U6954 (N_6954,N_312,N_2102);
xor U6955 (N_6955,N_2370,N_244);
or U6956 (N_6956,N_2309,N_1130);
and U6957 (N_6957,N_841,N_744);
nor U6958 (N_6958,N_2921,N_1951);
nand U6959 (N_6959,N_2701,N_2665);
nand U6960 (N_6960,N_1160,N_3202);
or U6961 (N_6961,N_3459,N_2259);
or U6962 (N_6962,N_1701,N_2961);
and U6963 (N_6963,N_1693,N_3018);
nand U6964 (N_6964,N_2180,N_3666);
and U6965 (N_6965,N_3098,N_3396);
nand U6966 (N_6966,N_25,N_1359);
xnor U6967 (N_6967,N_310,N_913);
or U6968 (N_6968,N_2179,N_394);
and U6969 (N_6969,N_3092,N_821);
nor U6970 (N_6970,N_3322,N_587);
and U6971 (N_6971,N_2437,N_3379);
nor U6972 (N_6972,N_2709,N_2183);
xor U6973 (N_6973,N_1571,N_2642);
nand U6974 (N_6974,N_2293,N_1074);
xnor U6975 (N_6975,N_757,N_1338);
or U6976 (N_6976,N_3817,N_625);
nor U6977 (N_6977,N_2657,N_3633);
and U6978 (N_6978,N_2813,N_727);
or U6979 (N_6979,N_3101,N_3354);
or U6980 (N_6980,N_1782,N_1644);
nor U6981 (N_6981,N_1451,N_3482);
and U6982 (N_6982,N_51,N_1106);
and U6983 (N_6983,N_1396,N_2986);
or U6984 (N_6984,N_609,N_3586);
nand U6985 (N_6985,N_3498,N_1423);
and U6986 (N_6986,N_1249,N_79);
or U6987 (N_6987,N_149,N_2501);
or U6988 (N_6988,N_1514,N_2642);
nand U6989 (N_6989,N_3845,N_1558);
nand U6990 (N_6990,N_2528,N_2788);
or U6991 (N_6991,N_3305,N_3817);
and U6992 (N_6992,N_2642,N_3503);
xnor U6993 (N_6993,N_1318,N_237);
nor U6994 (N_6994,N_2540,N_1901);
xor U6995 (N_6995,N_3714,N_3846);
or U6996 (N_6996,N_3636,N_1849);
nor U6997 (N_6997,N_3208,N_2806);
nor U6998 (N_6998,N_1032,N_246);
nand U6999 (N_6999,N_2429,N_673);
nand U7000 (N_7000,N_843,N_1178);
or U7001 (N_7001,N_713,N_2708);
and U7002 (N_7002,N_2361,N_3363);
nand U7003 (N_7003,N_1939,N_193);
nor U7004 (N_7004,N_3478,N_3110);
and U7005 (N_7005,N_182,N_2593);
and U7006 (N_7006,N_405,N_3666);
and U7007 (N_7007,N_3701,N_2040);
nand U7008 (N_7008,N_3070,N_3104);
or U7009 (N_7009,N_3269,N_2403);
and U7010 (N_7010,N_1280,N_2446);
nand U7011 (N_7011,N_2221,N_810);
nand U7012 (N_7012,N_1999,N_3656);
xor U7013 (N_7013,N_176,N_605);
or U7014 (N_7014,N_2777,N_1452);
nand U7015 (N_7015,N_1682,N_3257);
and U7016 (N_7016,N_1242,N_1375);
xor U7017 (N_7017,N_3233,N_713);
nand U7018 (N_7018,N_1814,N_2411);
nor U7019 (N_7019,N_2010,N_1407);
or U7020 (N_7020,N_1904,N_3604);
nor U7021 (N_7021,N_252,N_326);
and U7022 (N_7022,N_1342,N_2399);
and U7023 (N_7023,N_2743,N_2032);
nand U7024 (N_7024,N_79,N_2636);
nand U7025 (N_7025,N_3247,N_3939);
nor U7026 (N_7026,N_93,N_2720);
nor U7027 (N_7027,N_3602,N_2665);
nor U7028 (N_7028,N_3222,N_3124);
and U7029 (N_7029,N_2782,N_3432);
nor U7030 (N_7030,N_1334,N_355);
xnor U7031 (N_7031,N_2308,N_2486);
and U7032 (N_7032,N_1976,N_3973);
and U7033 (N_7033,N_334,N_620);
or U7034 (N_7034,N_1766,N_2622);
or U7035 (N_7035,N_2606,N_2056);
nor U7036 (N_7036,N_945,N_922);
or U7037 (N_7037,N_2920,N_2064);
nand U7038 (N_7038,N_2323,N_105);
xnor U7039 (N_7039,N_3735,N_2421);
nand U7040 (N_7040,N_837,N_3094);
and U7041 (N_7041,N_3832,N_2874);
nand U7042 (N_7042,N_1064,N_1583);
nand U7043 (N_7043,N_245,N_835);
nor U7044 (N_7044,N_968,N_1543);
and U7045 (N_7045,N_836,N_2303);
nor U7046 (N_7046,N_679,N_2389);
and U7047 (N_7047,N_2861,N_117);
and U7048 (N_7048,N_2097,N_1170);
or U7049 (N_7049,N_1849,N_1216);
or U7050 (N_7050,N_768,N_3394);
or U7051 (N_7051,N_1915,N_1132);
nor U7052 (N_7052,N_2119,N_1007);
xor U7053 (N_7053,N_126,N_2871);
and U7054 (N_7054,N_2755,N_2952);
nand U7055 (N_7055,N_1057,N_1209);
and U7056 (N_7056,N_3389,N_3172);
or U7057 (N_7057,N_1097,N_1942);
or U7058 (N_7058,N_854,N_2621);
nand U7059 (N_7059,N_2767,N_1340);
nand U7060 (N_7060,N_4,N_3330);
nor U7061 (N_7061,N_230,N_2526);
or U7062 (N_7062,N_2768,N_3388);
nand U7063 (N_7063,N_3833,N_3412);
nand U7064 (N_7064,N_19,N_3576);
nand U7065 (N_7065,N_2217,N_3330);
or U7066 (N_7066,N_359,N_3775);
and U7067 (N_7067,N_2491,N_2309);
nor U7068 (N_7068,N_1993,N_3599);
nor U7069 (N_7069,N_107,N_2588);
nor U7070 (N_7070,N_449,N_3565);
nand U7071 (N_7071,N_1884,N_2710);
or U7072 (N_7072,N_1481,N_3998);
and U7073 (N_7073,N_1005,N_260);
nand U7074 (N_7074,N_2215,N_825);
nand U7075 (N_7075,N_1467,N_1996);
or U7076 (N_7076,N_3412,N_478);
nor U7077 (N_7077,N_483,N_2624);
and U7078 (N_7078,N_2927,N_3991);
nor U7079 (N_7079,N_3739,N_2437);
nand U7080 (N_7080,N_1186,N_2761);
nand U7081 (N_7081,N_3062,N_722);
and U7082 (N_7082,N_3363,N_2498);
or U7083 (N_7083,N_3397,N_2844);
or U7084 (N_7084,N_1130,N_86);
xor U7085 (N_7085,N_522,N_3135);
xnor U7086 (N_7086,N_2924,N_1896);
nor U7087 (N_7087,N_2858,N_968);
or U7088 (N_7088,N_514,N_2751);
xnor U7089 (N_7089,N_226,N_1950);
nand U7090 (N_7090,N_2534,N_49);
xnor U7091 (N_7091,N_633,N_431);
and U7092 (N_7092,N_3346,N_1043);
nand U7093 (N_7093,N_529,N_2438);
nor U7094 (N_7094,N_945,N_3958);
nand U7095 (N_7095,N_684,N_3050);
or U7096 (N_7096,N_1426,N_1005);
or U7097 (N_7097,N_1562,N_671);
or U7098 (N_7098,N_779,N_410);
nor U7099 (N_7099,N_1875,N_2579);
xnor U7100 (N_7100,N_760,N_113);
or U7101 (N_7101,N_3597,N_855);
or U7102 (N_7102,N_167,N_2666);
nand U7103 (N_7103,N_3720,N_2640);
nor U7104 (N_7104,N_635,N_837);
nor U7105 (N_7105,N_2941,N_2199);
nor U7106 (N_7106,N_1572,N_657);
or U7107 (N_7107,N_1028,N_714);
xor U7108 (N_7108,N_1615,N_2181);
nand U7109 (N_7109,N_3350,N_2748);
and U7110 (N_7110,N_1101,N_1661);
nand U7111 (N_7111,N_3384,N_1490);
nor U7112 (N_7112,N_347,N_337);
nand U7113 (N_7113,N_2583,N_761);
nor U7114 (N_7114,N_3946,N_3075);
nor U7115 (N_7115,N_1777,N_2709);
nand U7116 (N_7116,N_2069,N_3898);
nand U7117 (N_7117,N_2694,N_2599);
nand U7118 (N_7118,N_3223,N_3894);
xor U7119 (N_7119,N_1651,N_3446);
nor U7120 (N_7120,N_2762,N_1936);
nand U7121 (N_7121,N_2255,N_3319);
xnor U7122 (N_7122,N_29,N_1514);
nor U7123 (N_7123,N_3373,N_2785);
or U7124 (N_7124,N_2125,N_3955);
nand U7125 (N_7125,N_1616,N_3877);
or U7126 (N_7126,N_1636,N_1457);
nor U7127 (N_7127,N_2759,N_1415);
or U7128 (N_7128,N_1548,N_428);
nor U7129 (N_7129,N_2674,N_748);
nand U7130 (N_7130,N_1964,N_983);
xor U7131 (N_7131,N_294,N_1238);
nor U7132 (N_7132,N_3579,N_3390);
and U7133 (N_7133,N_691,N_3639);
nor U7134 (N_7134,N_1488,N_2219);
and U7135 (N_7135,N_1581,N_3059);
nand U7136 (N_7136,N_96,N_2625);
nor U7137 (N_7137,N_3167,N_1119);
xnor U7138 (N_7138,N_851,N_1214);
nor U7139 (N_7139,N_3639,N_2294);
nor U7140 (N_7140,N_535,N_2016);
xnor U7141 (N_7141,N_2940,N_2477);
and U7142 (N_7142,N_171,N_666);
or U7143 (N_7143,N_1990,N_2428);
or U7144 (N_7144,N_1890,N_1609);
nand U7145 (N_7145,N_1031,N_3612);
xnor U7146 (N_7146,N_2632,N_3028);
nand U7147 (N_7147,N_3219,N_141);
or U7148 (N_7148,N_1424,N_1405);
or U7149 (N_7149,N_3830,N_3442);
nand U7150 (N_7150,N_1260,N_3037);
nand U7151 (N_7151,N_2624,N_2770);
or U7152 (N_7152,N_2649,N_627);
or U7153 (N_7153,N_556,N_1986);
nand U7154 (N_7154,N_1706,N_1370);
or U7155 (N_7155,N_57,N_1756);
nor U7156 (N_7156,N_1834,N_2662);
nand U7157 (N_7157,N_1022,N_1246);
nand U7158 (N_7158,N_2324,N_1893);
nor U7159 (N_7159,N_2143,N_1054);
nand U7160 (N_7160,N_2854,N_2908);
nor U7161 (N_7161,N_3760,N_2896);
nor U7162 (N_7162,N_1650,N_3432);
nor U7163 (N_7163,N_121,N_1817);
and U7164 (N_7164,N_1833,N_3712);
or U7165 (N_7165,N_368,N_1467);
or U7166 (N_7166,N_3303,N_2753);
or U7167 (N_7167,N_2107,N_2470);
nand U7168 (N_7168,N_3149,N_3030);
and U7169 (N_7169,N_3564,N_1874);
nand U7170 (N_7170,N_1285,N_1298);
or U7171 (N_7171,N_822,N_1479);
and U7172 (N_7172,N_3006,N_2711);
and U7173 (N_7173,N_2735,N_3656);
nor U7174 (N_7174,N_2973,N_1630);
or U7175 (N_7175,N_3533,N_1650);
nand U7176 (N_7176,N_3334,N_3579);
and U7177 (N_7177,N_1114,N_3518);
and U7178 (N_7178,N_2792,N_1780);
nand U7179 (N_7179,N_1867,N_1761);
or U7180 (N_7180,N_2374,N_2625);
and U7181 (N_7181,N_1663,N_2649);
or U7182 (N_7182,N_755,N_3287);
and U7183 (N_7183,N_12,N_1049);
nand U7184 (N_7184,N_1615,N_2767);
nor U7185 (N_7185,N_2148,N_2168);
xor U7186 (N_7186,N_3128,N_2368);
and U7187 (N_7187,N_275,N_1913);
xnor U7188 (N_7188,N_3826,N_296);
nand U7189 (N_7189,N_2559,N_3261);
and U7190 (N_7190,N_2367,N_2951);
nand U7191 (N_7191,N_2194,N_2284);
and U7192 (N_7192,N_2967,N_490);
or U7193 (N_7193,N_986,N_2406);
and U7194 (N_7194,N_1202,N_893);
nor U7195 (N_7195,N_1175,N_3867);
nor U7196 (N_7196,N_3157,N_2468);
and U7197 (N_7197,N_281,N_2844);
nor U7198 (N_7198,N_1320,N_1548);
or U7199 (N_7199,N_872,N_3152);
and U7200 (N_7200,N_3245,N_3126);
xor U7201 (N_7201,N_2721,N_1517);
or U7202 (N_7202,N_640,N_2643);
and U7203 (N_7203,N_3799,N_2219);
nand U7204 (N_7204,N_2703,N_3371);
nor U7205 (N_7205,N_2244,N_1776);
and U7206 (N_7206,N_2743,N_2467);
nor U7207 (N_7207,N_2409,N_2084);
nor U7208 (N_7208,N_2476,N_2504);
nor U7209 (N_7209,N_3228,N_2189);
xor U7210 (N_7210,N_2887,N_3121);
or U7211 (N_7211,N_2977,N_379);
nor U7212 (N_7212,N_56,N_1308);
or U7213 (N_7213,N_759,N_1887);
nand U7214 (N_7214,N_2953,N_3014);
nand U7215 (N_7215,N_317,N_3618);
or U7216 (N_7216,N_2,N_917);
and U7217 (N_7217,N_3447,N_2603);
or U7218 (N_7218,N_48,N_2651);
xor U7219 (N_7219,N_299,N_1653);
nor U7220 (N_7220,N_1439,N_2433);
nor U7221 (N_7221,N_3523,N_3957);
nand U7222 (N_7222,N_849,N_3215);
nand U7223 (N_7223,N_3948,N_793);
xnor U7224 (N_7224,N_3285,N_370);
and U7225 (N_7225,N_2181,N_3292);
or U7226 (N_7226,N_3733,N_1606);
or U7227 (N_7227,N_1125,N_1531);
and U7228 (N_7228,N_3275,N_1325);
nor U7229 (N_7229,N_2336,N_401);
or U7230 (N_7230,N_758,N_807);
or U7231 (N_7231,N_992,N_1756);
nand U7232 (N_7232,N_469,N_3998);
xnor U7233 (N_7233,N_876,N_1011);
and U7234 (N_7234,N_502,N_1714);
xnor U7235 (N_7235,N_2801,N_239);
or U7236 (N_7236,N_94,N_1533);
nand U7237 (N_7237,N_2665,N_1184);
nor U7238 (N_7238,N_325,N_2594);
nand U7239 (N_7239,N_2311,N_1279);
or U7240 (N_7240,N_3856,N_250);
and U7241 (N_7241,N_742,N_192);
nor U7242 (N_7242,N_1060,N_3988);
xor U7243 (N_7243,N_3034,N_1005);
and U7244 (N_7244,N_1758,N_2306);
nand U7245 (N_7245,N_1445,N_3065);
and U7246 (N_7246,N_580,N_612);
nand U7247 (N_7247,N_3133,N_1159);
or U7248 (N_7248,N_899,N_3675);
nand U7249 (N_7249,N_2218,N_3110);
nor U7250 (N_7250,N_3894,N_1576);
or U7251 (N_7251,N_148,N_2818);
nor U7252 (N_7252,N_636,N_408);
xor U7253 (N_7253,N_2107,N_1855);
and U7254 (N_7254,N_2361,N_1250);
or U7255 (N_7255,N_3078,N_2871);
or U7256 (N_7256,N_3422,N_1320);
and U7257 (N_7257,N_2509,N_165);
nor U7258 (N_7258,N_2979,N_1456);
nand U7259 (N_7259,N_3849,N_1385);
and U7260 (N_7260,N_2181,N_1463);
nand U7261 (N_7261,N_999,N_1650);
nor U7262 (N_7262,N_1599,N_3175);
or U7263 (N_7263,N_3450,N_3389);
nor U7264 (N_7264,N_3697,N_1103);
and U7265 (N_7265,N_102,N_671);
xnor U7266 (N_7266,N_3930,N_3039);
nor U7267 (N_7267,N_3335,N_285);
and U7268 (N_7268,N_1363,N_3158);
nand U7269 (N_7269,N_432,N_1524);
xor U7270 (N_7270,N_1379,N_127);
or U7271 (N_7271,N_2756,N_472);
and U7272 (N_7272,N_1042,N_573);
and U7273 (N_7273,N_1661,N_3688);
nand U7274 (N_7274,N_894,N_521);
nand U7275 (N_7275,N_2719,N_3214);
nor U7276 (N_7276,N_1470,N_3871);
nor U7277 (N_7277,N_3793,N_681);
or U7278 (N_7278,N_2745,N_3145);
and U7279 (N_7279,N_559,N_2948);
nor U7280 (N_7280,N_3591,N_2980);
and U7281 (N_7281,N_3009,N_2681);
or U7282 (N_7282,N_2025,N_3578);
and U7283 (N_7283,N_68,N_2803);
nor U7284 (N_7284,N_1327,N_2021);
nor U7285 (N_7285,N_2864,N_793);
nand U7286 (N_7286,N_1603,N_1180);
nor U7287 (N_7287,N_3138,N_2446);
nor U7288 (N_7288,N_300,N_2798);
xor U7289 (N_7289,N_2688,N_1827);
nor U7290 (N_7290,N_1175,N_2005);
and U7291 (N_7291,N_1392,N_1963);
nor U7292 (N_7292,N_779,N_1436);
xnor U7293 (N_7293,N_1241,N_3514);
nor U7294 (N_7294,N_836,N_1968);
xor U7295 (N_7295,N_3387,N_2114);
and U7296 (N_7296,N_3530,N_2729);
or U7297 (N_7297,N_3971,N_1126);
nand U7298 (N_7298,N_3865,N_1423);
nand U7299 (N_7299,N_1716,N_2848);
or U7300 (N_7300,N_2301,N_1916);
nor U7301 (N_7301,N_1894,N_3539);
and U7302 (N_7302,N_228,N_1122);
nand U7303 (N_7303,N_602,N_971);
xor U7304 (N_7304,N_788,N_1217);
or U7305 (N_7305,N_1558,N_1210);
nand U7306 (N_7306,N_3564,N_589);
nor U7307 (N_7307,N_512,N_3052);
or U7308 (N_7308,N_121,N_3820);
xor U7309 (N_7309,N_2355,N_2284);
nand U7310 (N_7310,N_66,N_3912);
xor U7311 (N_7311,N_1643,N_2665);
nand U7312 (N_7312,N_3303,N_609);
nor U7313 (N_7313,N_1628,N_1987);
nand U7314 (N_7314,N_834,N_2360);
and U7315 (N_7315,N_128,N_1045);
or U7316 (N_7316,N_3338,N_3165);
or U7317 (N_7317,N_2904,N_3707);
or U7318 (N_7318,N_1695,N_3706);
nor U7319 (N_7319,N_2493,N_1111);
or U7320 (N_7320,N_2914,N_378);
xnor U7321 (N_7321,N_3100,N_1668);
or U7322 (N_7322,N_2814,N_3788);
nand U7323 (N_7323,N_3718,N_262);
or U7324 (N_7324,N_3725,N_3770);
or U7325 (N_7325,N_985,N_3560);
nor U7326 (N_7326,N_1334,N_1971);
or U7327 (N_7327,N_2566,N_2300);
nand U7328 (N_7328,N_1074,N_552);
or U7329 (N_7329,N_1300,N_1340);
or U7330 (N_7330,N_1763,N_2199);
nand U7331 (N_7331,N_3055,N_2915);
nand U7332 (N_7332,N_479,N_1117);
nor U7333 (N_7333,N_1872,N_1655);
and U7334 (N_7334,N_3558,N_2762);
xor U7335 (N_7335,N_3691,N_2239);
nor U7336 (N_7336,N_2897,N_202);
or U7337 (N_7337,N_2011,N_2078);
nand U7338 (N_7338,N_816,N_729);
nand U7339 (N_7339,N_2277,N_3848);
nand U7340 (N_7340,N_2726,N_1208);
nand U7341 (N_7341,N_135,N_3669);
or U7342 (N_7342,N_3027,N_556);
nor U7343 (N_7343,N_2191,N_3548);
and U7344 (N_7344,N_3780,N_15);
and U7345 (N_7345,N_1421,N_499);
and U7346 (N_7346,N_51,N_3894);
or U7347 (N_7347,N_3587,N_2853);
nand U7348 (N_7348,N_1015,N_2122);
nand U7349 (N_7349,N_2198,N_3579);
nor U7350 (N_7350,N_1249,N_1851);
nand U7351 (N_7351,N_1527,N_1214);
xnor U7352 (N_7352,N_2041,N_3552);
nor U7353 (N_7353,N_2277,N_1102);
nand U7354 (N_7354,N_1335,N_2506);
and U7355 (N_7355,N_1562,N_236);
xor U7356 (N_7356,N_2929,N_1549);
nor U7357 (N_7357,N_3748,N_3891);
nand U7358 (N_7358,N_2900,N_3223);
or U7359 (N_7359,N_1831,N_2193);
nand U7360 (N_7360,N_2514,N_1653);
or U7361 (N_7361,N_3626,N_302);
nand U7362 (N_7362,N_908,N_3506);
or U7363 (N_7363,N_2404,N_3316);
and U7364 (N_7364,N_3677,N_3620);
or U7365 (N_7365,N_2004,N_441);
and U7366 (N_7366,N_777,N_313);
or U7367 (N_7367,N_1670,N_1771);
or U7368 (N_7368,N_3828,N_3063);
and U7369 (N_7369,N_1418,N_2490);
or U7370 (N_7370,N_3900,N_3824);
nor U7371 (N_7371,N_2198,N_3036);
and U7372 (N_7372,N_115,N_559);
nand U7373 (N_7373,N_1441,N_3874);
or U7374 (N_7374,N_5,N_3435);
and U7375 (N_7375,N_2851,N_2574);
or U7376 (N_7376,N_2917,N_999);
nor U7377 (N_7377,N_2112,N_3778);
nor U7378 (N_7378,N_1951,N_174);
and U7379 (N_7379,N_2203,N_3559);
nor U7380 (N_7380,N_705,N_2105);
nand U7381 (N_7381,N_2222,N_783);
or U7382 (N_7382,N_3387,N_1187);
nor U7383 (N_7383,N_1617,N_1016);
nor U7384 (N_7384,N_1909,N_283);
nand U7385 (N_7385,N_1212,N_1079);
nor U7386 (N_7386,N_1018,N_1589);
and U7387 (N_7387,N_1485,N_328);
and U7388 (N_7388,N_308,N_3479);
or U7389 (N_7389,N_2359,N_1630);
xor U7390 (N_7390,N_1616,N_2992);
xor U7391 (N_7391,N_2154,N_291);
and U7392 (N_7392,N_3146,N_448);
and U7393 (N_7393,N_2579,N_2298);
and U7394 (N_7394,N_1289,N_1077);
or U7395 (N_7395,N_3080,N_97);
xnor U7396 (N_7396,N_838,N_1450);
and U7397 (N_7397,N_2693,N_301);
nand U7398 (N_7398,N_2657,N_3171);
nor U7399 (N_7399,N_3219,N_601);
nor U7400 (N_7400,N_3351,N_1376);
and U7401 (N_7401,N_3540,N_2185);
or U7402 (N_7402,N_1292,N_2248);
or U7403 (N_7403,N_2327,N_611);
nand U7404 (N_7404,N_320,N_3659);
or U7405 (N_7405,N_3004,N_3913);
and U7406 (N_7406,N_2058,N_409);
nand U7407 (N_7407,N_284,N_1201);
nor U7408 (N_7408,N_2090,N_3306);
nand U7409 (N_7409,N_602,N_287);
or U7410 (N_7410,N_3182,N_1490);
or U7411 (N_7411,N_2325,N_2765);
nand U7412 (N_7412,N_2025,N_3666);
nor U7413 (N_7413,N_3591,N_2413);
or U7414 (N_7414,N_626,N_1318);
nand U7415 (N_7415,N_292,N_2436);
and U7416 (N_7416,N_3035,N_916);
or U7417 (N_7417,N_2503,N_424);
or U7418 (N_7418,N_377,N_2630);
xnor U7419 (N_7419,N_1292,N_3761);
nand U7420 (N_7420,N_20,N_1589);
nor U7421 (N_7421,N_3789,N_3421);
nand U7422 (N_7422,N_139,N_3261);
and U7423 (N_7423,N_2719,N_812);
nand U7424 (N_7424,N_3317,N_2626);
xnor U7425 (N_7425,N_3530,N_3549);
and U7426 (N_7426,N_3241,N_2740);
nand U7427 (N_7427,N_564,N_194);
nor U7428 (N_7428,N_2831,N_1864);
xnor U7429 (N_7429,N_2231,N_237);
xnor U7430 (N_7430,N_2663,N_2932);
or U7431 (N_7431,N_916,N_2177);
xnor U7432 (N_7432,N_441,N_2610);
or U7433 (N_7433,N_954,N_2471);
or U7434 (N_7434,N_2120,N_3382);
nor U7435 (N_7435,N_2995,N_1075);
nor U7436 (N_7436,N_2708,N_3886);
nand U7437 (N_7437,N_2953,N_348);
and U7438 (N_7438,N_2395,N_3048);
xor U7439 (N_7439,N_1490,N_2492);
and U7440 (N_7440,N_1626,N_1392);
nor U7441 (N_7441,N_82,N_2054);
xor U7442 (N_7442,N_2022,N_3663);
nand U7443 (N_7443,N_763,N_1298);
nor U7444 (N_7444,N_1425,N_939);
and U7445 (N_7445,N_3134,N_843);
nor U7446 (N_7446,N_3729,N_96);
or U7447 (N_7447,N_610,N_3435);
nand U7448 (N_7448,N_491,N_2959);
and U7449 (N_7449,N_2860,N_1703);
or U7450 (N_7450,N_1973,N_1247);
or U7451 (N_7451,N_287,N_2012);
and U7452 (N_7452,N_1107,N_3243);
nor U7453 (N_7453,N_1889,N_3819);
and U7454 (N_7454,N_3362,N_2262);
or U7455 (N_7455,N_2645,N_1512);
nand U7456 (N_7456,N_2634,N_22);
nor U7457 (N_7457,N_2596,N_1798);
or U7458 (N_7458,N_2156,N_57);
and U7459 (N_7459,N_2336,N_2992);
nor U7460 (N_7460,N_3290,N_2074);
or U7461 (N_7461,N_3418,N_1654);
and U7462 (N_7462,N_3129,N_2792);
or U7463 (N_7463,N_1188,N_782);
nand U7464 (N_7464,N_340,N_939);
nor U7465 (N_7465,N_870,N_3333);
nand U7466 (N_7466,N_1347,N_3829);
and U7467 (N_7467,N_2312,N_2004);
nor U7468 (N_7468,N_3512,N_3994);
xnor U7469 (N_7469,N_3147,N_954);
or U7470 (N_7470,N_106,N_717);
nand U7471 (N_7471,N_3063,N_3199);
xnor U7472 (N_7472,N_3737,N_1871);
and U7473 (N_7473,N_1377,N_3106);
or U7474 (N_7474,N_1775,N_2836);
or U7475 (N_7475,N_3975,N_36);
nand U7476 (N_7476,N_1273,N_414);
and U7477 (N_7477,N_429,N_3204);
nand U7478 (N_7478,N_72,N_2852);
xor U7479 (N_7479,N_3174,N_1055);
nor U7480 (N_7480,N_3226,N_3557);
nor U7481 (N_7481,N_3526,N_2382);
xor U7482 (N_7482,N_1518,N_1262);
nand U7483 (N_7483,N_3204,N_2959);
nor U7484 (N_7484,N_430,N_1286);
nor U7485 (N_7485,N_2800,N_2519);
nand U7486 (N_7486,N_1614,N_1559);
nor U7487 (N_7487,N_3119,N_1949);
or U7488 (N_7488,N_2619,N_3672);
nand U7489 (N_7489,N_3521,N_2187);
nor U7490 (N_7490,N_1763,N_1628);
or U7491 (N_7491,N_704,N_1274);
nor U7492 (N_7492,N_2568,N_3044);
nor U7493 (N_7493,N_2757,N_267);
or U7494 (N_7494,N_639,N_3943);
nor U7495 (N_7495,N_1507,N_1164);
nand U7496 (N_7496,N_1154,N_3357);
or U7497 (N_7497,N_3292,N_2838);
xor U7498 (N_7498,N_3987,N_64);
nor U7499 (N_7499,N_1060,N_297);
and U7500 (N_7500,N_899,N_2042);
nor U7501 (N_7501,N_126,N_1984);
or U7502 (N_7502,N_1898,N_790);
and U7503 (N_7503,N_771,N_1631);
nand U7504 (N_7504,N_893,N_3799);
or U7505 (N_7505,N_3218,N_2976);
nor U7506 (N_7506,N_3868,N_407);
or U7507 (N_7507,N_3521,N_3568);
or U7508 (N_7508,N_2451,N_2820);
and U7509 (N_7509,N_803,N_2070);
xor U7510 (N_7510,N_203,N_2090);
or U7511 (N_7511,N_1113,N_526);
xnor U7512 (N_7512,N_3983,N_264);
nand U7513 (N_7513,N_554,N_1343);
nor U7514 (N_7514,N_2487,N_3425);
nor U7515 (N_7515,N_3448,N_344);
and U7516 (N_7516,N_2075,N_1772);
and U7517 (N_7517,N_2228,N_1283);
and U7518 (N_7518,N_1611,N_1933);
or U7519 (N_7519,N_1073,N_172);
or U7520 (N_7520,N_3898,N_3255);
nand U7521 (N_7521,N_861,N_3660);
and U7522 (N_7522,N_3240,N_2557);
and U7523 (N_7523,N_578,N_1371);
and U7524 (N_7524,N_781,N_1169);
nand U7525 (N_7525,N_1805,N_3116);
or U7526 (N_7526,N_955,N_3591);
xor U7527 (N_7527,N_3937,N_2411);
nand U7528 (N_7528,N_703,N_884);
nor U7529 (N_7529,N_2855,N_3261);
and U7530 (N_7530,N_3917,N_2211);
xor U7531 (N_7531,N_1058,N_2176);
and U7532 (N_7532,N_79,N_735);
nand U7533 (N_7533,N_1297,N_769);
or U7534 (N_7534,N_1454,N_2672);
or U7535 (N_7535,N_1365,N_935);
and U7536 (N_7536,N_1753,N_1707);
nor U7537 (N_7537,N_87,N_3644);
and U7538 (N_7538,N_3273,N_1424);
and U7539 (N_7539,N_1179,N_672);
or U7540 (N_7540,N_2012,N_3282);
and U7541 (N_7541,N_2884,N_2820);
nand U7542 (N_7542,N_2740,N_2547);
nor U7543 (N_7543,N_2650,N_1383);
nand U7544 (N_7544,N_3594,N_2444);
nor U7545 (N_7545,N_679,N_2925);
nand U7546 (N_7546,N_2850,N_1591);
and U7547 (N_7547,N_567,N_3050);
nor U7548 (N_7548,N_2048,N_2005);
nor U7549 (N_7549,N_173,N_3388);
nand U7550 (N_7550,N_448,N_3552);
nand U7551 (N_7551,N_3562,N_1817);
and U7552 (N_7552,N_44,N_3762);
nand U7553 (N_7553,N_137,N_3785);
and U7554 (N_7554,N_2614,N_741);
nor U7555 (N_7555,N_3030,N_2518);
and U7556 (N_7556,N_310,N_2835);
xor U7557 (N_7557,N_928,N_2080);
nor U7558 (N_7558,N_1191,N_255);
and U7559 (N_7559,N_3869,N_2001);
and U7560 (N_7560,N_3866,N_1865);
and U7561 (N_7561,N_1939,N_3921);
nor U7562 (N_7562,N_1471,N_2695);
and U7563 (N_7563,N_1061,N_3270);
xnor U7564 (N_7564,N_1813,N_1585);
nand U7565 (N_7565,N_993,N_2358);
nor U7566 (N_7566,N_1520,N_3285);
or U7567 (N_7567,N_3025,N_2771);
nand U7568 (N_7568,N_2110,N_2106);
xnor U7569 (N_7569,N_254,N_3899);
nand U7570 (N_7570,N_3419,N_1418);
xor U7571 (N_7571,N_562,N_3934);
and U7572 (N_7572,N_581,N_136);
and U7573 (N_7573,N_3885,N_726);
or U7574 (N_7574,N_3771,N_1910);
and U7575 (N_7575,N_2605,N_758);
nor U7576 (N_7576,N_3829,N_834);
and U7577 (N_7577,N_1167,N_3181);
and U7578 (N_7578,N_2292,N_2579);
nand U7579 (N_7579,N_1459,N_990);
nand U7580 (N_7580,N_918,N_1917);
xor U7581 (N_7581,N_3327,N_3474);
nor U7582 (N_7582,N_1410,N_3516);
or U7583 (N_7583,N_1885,N_2344);
or U7584 (N_7584,N_3033,N_2078);
or U7585 (N_7585,N_3958,N_768);
and U7586 (N_7586,N_3713,N_1277);
or U7587 (N_7587,N_2463,N_3472);
and U7588 (N_7588,N_232,N_241);
or U7589 (N_7589,N_2182,N_616);
nor U7590 (N_7590,N_695,N_3924);
nand U7591 (N_7591,N_144,N_713);
and U7592 (N_7592,N_693,N_2874);
xor U7593 (N_7593,N_1542,N_1596);
or U7594 (N_7594,N_2302,N_3457);
nand U7595 (N_7595,N_2668,N_951);
and U7596 (N_7596,N_2679,N_1277);
and U7597 (N_7597,N_1096,N_1289);
and U7598 (N_7598,N_691,N_2293);
nand U7599 (N_7599,N_656,N_316);
nor U7600 (N_7600,N_2433,N_575);
or U7601 (N_7601,N_3039,N_342);
nand U7602 (N_7602,N_2048,N_3998);
or U7603 (N_7603,N_1772,N_1349);
nand U7604 (N_7604,N_338,N_144);
or U7605 (N_7605,N_1246,N_3019);
nor U7606 (N_7606,N_359,N_529);
and U7607 (N_7607,N_1603,N_3021);
nor U7608 (N_7608,N_1183,N_229);
and U7609 (N_7609,N_2579,N_1217);
nor U7610 (N_7610,N_3117,N_1320);
or U7611 (N_7611,N_2528,N_766);
xnor U7612 (N_7612,N_2507,N_3722);
or U7613 (N_7613,N_529,N_488);
and U7614 (N_7614,N_3459,N_60);
nor U7615 (N_7615,N_1360,N_2916);
xnor U7616 (N_7616,N_1767,N_2914);
nand U7617 (N_7617,N_3925,N_92);
nor U7618 (N_7618,N_11,N_1422);
and U7619 (N_7619,N_2075,N_1505);
nand U7620 (N_7620,N_43,N_3450);
nand U7621 (N_7621,N_1679,N_1221);
nor U7622 (N_7622,N_2920,N_1668);
or U7623 (N_7623,N_67,N_213);
or U7624 (N_7624,N_2116,N_2107);
nor U7625 (N_7625,N_2608,N_2996);
and U7626 (N_7626,N_1700,N_863);
xnor U7627 (N_7627,N_3067,N_513);
nand U7628 (N_7628,N_1429,N_1861);
or U7629 (N_7629,N_3957,N_1956);
and U7630 (N_7630,N_3716,N_1946);
and U7631 (N_7631,N_1088,N_3397);
nand U7632 (N_7632,N_3459,N_2530);
and U7633 (N_7633,N_3479,N_3674);
or U7634 (N_7634,N_2240,N_2289);
and U7635 (N_7635,N_3888,N_1876);
and U7636 (N_7636,N_1421,N_625);
xnor U7637 (N_7637,N_486,N_1141);
and U7638 (N_7638,N_164,N_2118);
and U7639 (N_7639,N_2511,N_1490);
nand U7640 (N_7640,N_3190,N_2909);
and U7641 (N_7641,N_3836,N_3661);
nor U7642 (N_7642,N_2701,N_2084);
or U7643 (N_7643,N_1109,N_3586);
or U7644 (N_7644,N_133,N_3515);
xor U7645 (N_7645,N_722,N_1136);
nor U7646 (N_7646,N_3152,N_1819);
nor U7647 (N_7647,N_713,N_965);
xnor U7648 (N_7648,N_3083,N_2980);
or U7649 (N_7649,N_2144,N_10);
nor U7650 (N_7650,N_3741,N_2137);
and U7651 (N_7651,N_1629,N_2096);
nand U7652 (N_7652,N_32,N_1356);
nand U7653 (N_7653,N_2821,N_2608);
and U7654 (N_7654,N_2580,N_2285);
xor U7655 (N_7655,N_467,N_637);
nor U7656 (N_7656,N_2420,N_849);
or U7657 (N_7657,N_3728,N_3493);
and U7658 (N_7658,N_3389,N_1697);
or U7659 (N_7659,N_122,N_3276);
and U7660 (N_7660,N_1912,N_684);
or U7661 (N_7661,N_3030,N_3453);
nor U7662 (N_7662,N_531,N_2447);
or U7663 (N_7663,N_63,N_2485);
nand U7664 (N_7664,N_842,N_686);
nor U7665 (N_7665,N_2676,N_261);
and U7666 (N_7666,N_1261,N_1816);
nor U7667 (N_7667,N_1330,N_1519);
xnor U7668 (N_7668,N_9,N_2675);
nor U7669 (N_7669,N_2351,N_3142);
nor U7670 (N_7670,N_1229,N_2208);
or U7671 (N_7671,N_2243,N_393);
and U7672 (N_7672,N_1915,N_287);
nand U7673 (N_7673,N_2769,N_326);
nor U7674 (N_7674,N_2318,N_2974);
or U7675 (N_7675,N_3302,N_1425);
nand U7676 (N_7676,N_3106,N_3939);
and U7677 (N_7677,N_2168,N_3719);
and U7678 (N_7678,N_1095,N_1015);
nand U7679 (N_7679,N_2476,N_3333);
nor U7680 (N_7680,N_503,N_2718);
nor U7681 (N_7681,N_2262,N_1619);
nand U7682 (N_7682,N_186,N_935);
nor U7683 (N_7683,N_995,N_252);
or U7684 (N_7684,N_1157,N_1041);
and U7685 (N_7685,N_3432,N_715);
and U7686 (N_7686,N_1629,N_3616);
nand U7687 (N_7687,N_2686,N_2846);
and U7688 (N_7688,N_2373,N_73);
and U7689 (N_7689,N_718,N_3062);
and U7690 (N_7690,N_1072,N_344);
xor U7691 (N_7691,N_3383,N_1656);
and U7692 (N_7692,N_445,N_135);
or U7693 (N_7693,N_227,N_3303);
nor U7694 (N_7694,N_277,N_1243);
and U7695 (N_7695,N_3121,N_2845);
nor U7696 (N_7696,N_1086,N_12);
nor U7697 (N_7697,N_94,N_2283);
or U7698 (N_7698,N_3643,N_3216);
and U7699 (N_7699,N_3584,N_3017);
or U7700 (N_7700,N_3859,N_2633);
and U7701 (N_7701,N_492,N_1736);
nor U7702 (N_7702,N_1716,N_1568);
nor U7703 (N_7703,N_2186,N_877);
nor U7704 (N_7704,N_3579,N_2526);
and U7705 (N_7705,N_3555,N_1932);
nand U7706 (N_7706,N_2511,N_133);
or U7707 (N_7707,N_2085,N_2605);
nand U7708 (N_7708,N_924,N_2913);
nor U7709 (N_7709,N_1017,N_20);
or U7710 (N_7710,N_1024,N_1307);
and U7711 (N_7711,N_3406,N_110);
or U7712 (N_7712,N_2677,N_2529);
and U7713 (N_7713,N_2384,N_671);
nor U7714 (N_7714,N_1771,N_1130);
or U7715 (N_7715,N_3828,N_3794);
xor U7716 (N_7716,N_1452,N_149);
nand U7717 (N_7717,N_3703,N_777);
and U7718 (N_7718,N_3834,N_3455);
or U7719 (N_7719,N_3813,N_3495);
and U7720 (N_7720,N_1099,N_3625);
or U7721 (N_7721,N_1434,N_1256);
nor U7722 (N_7722,N_2963,N_530);
or U7723 (N_7723,N_3938,N_3944);
nor U7724 (N_7724,N_1303,N_3802);
nand U7725 (N_7725,N_453,N_484);
xor U7726 (N_7726,N_1728,N_2960);
and U7727 (N_7727,N_1938,N_304);
and U7728 (N_7728,N_145,N_2394);
or U7729 (N_7729,N_3221,N_1324);
or U7730 (N_7730,N_1000,N_2417);
nand U7731 (N_7731,N_3095,N_1449);
nand U7732 (N_7732,N_1140,N_1289);
nor U7733 (N_7733,N_2314,N_995);
or U7734 (N_7734,N_1909,N_2936);
xnor U7735 (N_7735,N_382,N_1079);
nand U7736 (N_7736,N_925,N_3715);
and U7737 (N_7737,N_615,N_440);
xor U7738 (N_7738,N_3500,N_3192);
nor U7739 (N_7739,N_918,N_908);
nor U7740 (N_7740,N_384,N_3416);
nand U7741 (N_7741,N_2571,N_3232);
or U7742 (N_7742,N_3235,N_314);
xnor U7743 (N_7743,N_3061,N_1710);
or U7744 (N_7744,N_1376,N_3557);
and U7745 (N_7745,N_2862,N_514);
or U7746 (N_7746,N_542,N_1542);
nor U7747 (N_7747,N_2999,N_1517);
nor U7748 (N_7748,N_2837,N_2590);
nor U7749 (N_7749,N_55,N_467);
nand U7750 (N_7750,N_1308,N_2643);
and U7751 (N_7751,N_1947,N_1928);
and U7752 (N_7752,N_2007,N_2561);
and U7753 (N_7753,N_812,N_2290);
or U7754 (N_7754,N_2206,N_1404);
or U7755 (N_7755,N_2436,N_1105);
nor U7756 (N_7756,N_3005,N_3604);
xnor U7757 (N_7757,N_1473,N_3326);
nor U7758 (N_7758,N_1429,N_1641);
nand U7759 (N_7759,N_3088,N_1153);
and U7760 (N_7760,N_2929,N_3204);
nor U7761 (N_7761,N_3719,N_873);
or U7762 (N_7762,N_3835,N_2382);
nor U7763 (N_7763,N_250,N_1734);
and U7764 (N_7764,N_494,N_3264);
nand U7765 (N_7765,N_1213,N_3219);
nor U7766 (N_7766,N_145,N_2308);
nand U7767 (N_7767,N_1729,N_3054);
nand U7768 (N_7768,N_2700,N_2303);
and U7769 (N_7769,N_1204,N_3095);
nor U7770 (N_7770,N_375,N_1150);
nor U7771 (N_7771,N_3591,N_2902);
nor U7772 (N_7772,N_3480,N_1591);
nand U7773 (N_7773,N_1352,N_556);
nand U7774 (N_7774,N_184,N_3690);
nor U7775 (N_7775,N_675,N_2872);
xnor U7776 (N_7776,N_226,N_2077);
nor U7777 (N_7777,N_74,N_2999);
and U7778 (N_7778,N_965,N_3016);
or U7779 (N_7779,N_1818,N_2128);
nand U7780 (N_7780,N_2453,N_410);
or U7781 (N_7781,N_1034,N_829);
nand U7782 (N_7782,N_3936,N_2467);
or U7783 (N_7783,N_3094,N_3985);
xor U7784 (N_7784,N_3901,N_1878);
or U7785 (N_7785,N_659,N_1903);
nor U7786 (N_7786,N_654,N_1636);
nor U7787 (N_7787,N_3791,N_3140);
and U7788 (N_7788,N_584,N_2202);
or U7789 (N_7789,N_507,N_461);
or U7790 (N_7790,N_1799,N_1290);
xor U7791 (N_7791,N_3798,N_1596);
xnor U7792 (N_7792,N_1899,N_1206);
and U7793 (N_7793,N_347,N_818);
or U7794 (N_7794,N_2673,N_3481);
nor U7795 (N_7795,N_20,N_3352);
or U7796 (N_7796,N_1061,N_169);
or U7797 (N_7797,N_3343,N_1211);
and U7798 (N_7798,N_1040,N_3445);
nand U7799 (N_7799,N_584,N_3742);
nor U7800 (N_7800,N_1151,N_1725);
and U7801 (N_7801,N_773,N_474);
and U7802 (N_7802,N_3706,N_1454);
nand U7803 (N_7803,N_3992,N_3635);
or U7804 (N_7804,N_1640,N_2484);
nand U7805 (N_7805,N_1090,N_789);
xor U7806 (N_7806,N_3592,N_3508);
and U7807 (N_7807,N_2879,N_3820);
nand U7808 (N_7808,N_3273,N_3096);
and U7809 (N_7809,N_599,N_3480);
nor U7810 (N_7810,N_489,N_1852);
nand U7811 (N_7811,N_1409,N_2063);
nand U7812 (N_7812,N_3830,N_3606);
or U7813 (N_7813,N_1508,N_1133);
nor U7814 (N_7814,N_1702,N_1386);
nand U7815 (N_7815,N_2439,N_1420);
nand U7816 (N_7816,N_2280,N_2208);
nor U7817 (N_7817,N_2645,N_3092);
and U7818 (N_7818,N_1442,N_2332);
nor U7819 (N_7819,N_657,N_1926);
nor U7820 (N_7820,N_2873,N_1551);
or U7821 (N_7821,N_2265,N_916);
or U7822 (N_7822,N_2460,N_305);
and U7823 (N_7823,N_1876,N_342);
nor U7824 (N_7824,N_747,N_252);
nor U7825 (N_7825,N_1257,N_3104);
nand U7826 (N_7826,N_3167,N_2364);
nand U7827 (N_7827,N_2489,N_480);
nor U7828 (N_7828,N_1069,N_1079);
and U7829 (N_7829,N_55,N_1437);
and U7830 (N_7830,N_910,N_3018);
xor U7831 (N_7831,N_1446,N_597);
nand U7832 (N_7832,N_3554,N_2726);
nor U7833 (N_7833,N_1748,N_3882);
nor U7834 (N_7834,N_3558,N_137);
nand U7835 (N_7835,N_908,N_284);
nor U7836 (N_7836,N_2012,N_3946);
nand U7837 (N_7837,N_2291,N_1446);
or U7838 (N_7838,N_1288,N_1866);
or U7839 (N_7839,N_2401,N_143);
and U7840 (N_7840,N_2594,N_1333);
xor U7841 (N_7841,N_3755,N_1186);
and U7842 (N_7842,N_3309,N_180);
nor U7843 (N_7843,N_2007,N_2179);
and U7844 (N_7844,N_2483,N_3317);
nor U7845 (N_7845,N_3257,N_759);
nand U7846 (N_7846,N_3650,N_2715);
nor U7847 (N_7847,N_69,N_2168);
or U7848 (N_7848,N_1312,N_3114);
or U7849 (N_7849,N_3008,N_1974);
and U7850 (N_7850,N_398,N_965);
xnor U7851 (N_7851,N_2074,N_2940);
nand U7852 (N_7852,N_1475,N_1917);
nand U7853 (N_7853,N_3750,N_402);
nor U7854 (N_7854,N_1636,N_3254);
nand U7855 (N_7855,N_1691,N_2544);
or U7856 (N_7856,N_2615,N_140);
nor U7857 (N_7857,N_38,N_2953);
nand U7858 (N_7858,N_3010,N_231);
or U7859 (N_7859,N_3359,N_2349);
and U7860 (N_7860,N_728,N_1317);
and U7861 (N_7861,N_3414,N_2711);
xor U7862 (N_7862,N_1042,N_2433);
nor U7863 (N_7863,N_2693,N_794);
nand U7864 (N_7864,N_235,N_2608);
or U7865 (N_7865,N_1370,N_3869);
nand U7866 (N_7866,N_3004,N_442);
or U7867 (N_7867,N_2631,N_2613);
nor U7868 (N_7868,N_3521,N_1568);
and U7869 (N_7869,N_302,N_1910);
or U7870 (N_7870,N_2456,N_1219);
or U7871 (N_7871,N_564,N_2690);
or U7872 (N_7872,N_2655,N_3121);
xnor U7873 (N_7873,N_1603,N_1218);
xor U7874 (N_7874,N_1975,N_3737);
nor U7875 (N_7875,N_401,N_2927);
xnor U7876 (N_7876,N_76,N_701);
xor U7877 (N_7877,N_884,N_3791);
or U7878 (N_7878,N_3832,N_2982);
nand U7879 (N_7879,N_1820,N_203);
nor U7880 (N_7880,N_1186,N_2901);
nor U7881 (N_7881,N_3039,N_3101);
or U7882 (N_7882,N_2463,N_341);
or U7883 (N_7883,N_3461,N_1804);
nor U7884 (N_7884,N_3251,N_3000);
or U7885 (N_7885,N_119,N_2626);
or U7886 (N_7886,N_3580,N_125);
nand U7887 (N_7887,N_1336,N_3522);
nand U7888 (N_7888,N_2986,N_2504);
xor U7889 (N_7889,N_1502,N_1133);
and U7890 (N_7890,N_1458,N_2206);
nor U7891 (N_7891,N_3133,N_1867);
or U7892 (N_7892,N_125,N_3304);
and U7893 (N_7893,N_2181,N_3898);
nor U7894 (N_7894,N_620,N_3510);
nand U7895 (N_7895,N_833,N_2380);
and U7896 (N_7896,N_3166,N_3085);
and U7897 (N_7897,N_2172,N_1886);
or U7898 (N_7898,N_1944,N_2951);
and U7899 (N_7899,N_3835,N_1130);
nand U7900 (N_7900,N_598,N_1275);
nand U7901 (N_7901,N_1876,N_2505);
xnor U7902 (N_7902,N_3596,N_1457);
nand U7903 (N_7903,N_1762,N_3952);
nor U7904 (N_7904,N_3857,N_2700);
nand U7905 (N_7905,N_1263,N_715);
and U7906 (N_7906,N_2086,N_3014);
or U7907 (N_7907,N_3526,N_1780);
nor U7908 (N_7908,N_3392,N_3956);
nor U7909 (N_7909,N_819,N_1730);
nand U7910 (N_7910,N_3124,N_2002);
nand U7911 (N_7911,N_172,N_2638);
xor U7912 (N_7912,N_2165,N_862);
xnor U7913 (N_7913,N_2268,N_2815);
nor U7914 (N_7914,N_2227,N_249);
nand U7915 (N_7915,N_2511,N_433);
nor U7916 (N_7916,N_3010,N_2602);
or U7917 (N_7917,N_2530,N_3103);
or U7918 (N_7918,N_2952,N_503);
nand U7919 (N_7919,N_594,N_2543);
nor U7920 (N_7920,N_2390,N_3210);
xnor U7921 (N_7921,N_3745,N_3840);
nand U7922 (N_7922,N_3390,N_3062);
or U7923 (N_7923,N_3234,N_321);
or U7924 (N_7924,N_139,N_3370);
or U7925 (N_7925,N_3671,N_2026);
nor U7926 (N_7926,N_1155,N_2477);
and U7927 (N_7927,N_1033,N_3443);
nand U7928 (N_7928,N_1633,N_1291);
and U7929 (N_7929,N_1064,N_3940);
or U7930 (N_7930,N_3353,N_2873);
and U7931 (N_7931,N_1466,N_1258);
and U7932 (N_7932,N_1380,N_2622);
and U7933 (N_7933,N_1341,N_2136);
nand U7934 (N_7934,N_1063,N_2562);
nor U7935 (N_7935,N_601,N_3696);
nand U7936 (N_7936,N_2527,N_3182);
and U7937 (N_7937,N_1928,N_850);
or U7938 (N_7938,N_794,N_2908);
xnor U7939 (N_7939,N_3314,N_844);
nor U7940 (N_7940,N_1848,N_1942);
xor U7941 (N_7941,N_790,N_2241);
nor U7942 (N_7942,N_2537,N_1393);
nor U7943 (N_7943,N_581,N_1265);
or U7944 (N_7944,N_1224,N_2190);
nor U7945 (N_7945,N_570,N_2930);
nand U7946 (N_7946,N_3464,N_1659);
and U7947 (N_7947,N_3128,N_3249);
nor U7948 (N_7948,N_2103,N_921);
and U7949 (N_7949,N_3961,N_1003);
nand U7950 (N_7950,N_544,N_278);
or U7951 (N_7951,N_979,N_2472);
and U7952 (N_7952,N_1632,N_2488);
nand U7953 (N_7953,N_792,N_1035);
nand U7954 (N_7954,N_1174,N_1081);
or U7955 (N_7955,N_1121,N_2081);
and U7956 (N_7956,N_1411,N_1025);
nor U7957 (N_7957,N_1793,N_819);
or U7958 (N_7958,N_2899,N_1321);
nand U7959 (N_7959,N_1864,N_575);
nor U7960 (N_7960,N_3100,N_2028);
nand U7961 (N_7961,N_3280,N_3271);
nor U7962 (N_7962,N_417,N_3575);
xnor U7963 (N_7963,N_2297,N_1087);
nand U7964 (N_7964,N_3039,N_3079);
or U7965 (N_7965,N_215,N_1195);
xor U7966 (N_7966,N_483,N_1760);
nor U7967 (N_7967,N_1925,N_716);
or U7968 (N_7968,N_1644,N_1477);
nand U7969 (N_7969,N_2030,N_2663);
xnor U7970 (N_7970,N_2523,N_3003);
or U7971 (N_7971,N_2542,N_3580);
nor U7972 (N_7972,N_3842,N_705);
nand U7973 (N_7973,N_2841,N_2743);
and U7974 (N_7974,N_1478,N_1538);
nand U7975 (N_7975,N_563,N_797);
or U7976 (N_7976,N_522,N_1442);
and U7977 (N_7977,N_544,N_1844);
or U7978 (N_7978,N_3733,N_3985);
xnor U7979 (N_7979,N_2912,N_3483);
nand U7980 (N_7980,N_1561,N_1650);
xor U7981 (N_7981,N_966,N_3809);
nand U7982 (N_7982,N_3220,N_1254);
and U7983 (N_7983,N_3296,N_1369);
or U7984 (N_7984,N_3970,N_790);
or U7985 (N_7985,N_13,N_582);
nand U7986 (N_7986,N_873,N_2126);
xnor U7987 (N_7987,N_3240,N_756);
or U7988 (N_7988,N_1269,N_2481);
or U7989 (N_7989,N_2329,N_3586);
or U7990 (N_7990,N_2696,N_1970);
and U7991 (N_7991,N_1045,N_2001);
xor U7992 (N_7992,N_3232,N_3956);
nand U7993 (N_7993,N_2732,N_1635);
nor U7994 (N_7994,N_3105,N_2128);
or U7995 (N_7995,N_3236,N_2206);
nor U7996 (N_7996,N_2253,N_2063);
and U7997 (N_7997,N_2063,N_741);
or U7998 (N_7998,N_3778,N_1918);
nand U7999 (N_7999,N_3521,N_3393);
nor U8000 (N_8000,N_5329,N_4817);
nand U8001 (N_8001,N_7881,N_4282);
or U8002 (N_8002,N_4091,N_5830);
and U8003 (N_8003,N_6548,N_7762);
nor U8004 (N_8004,N_4059,N_6794);
or U8005 (N_8005,N_7134,N_7900);
and U8006 (N_8006,N_4149,N_5735);
or U8007 (N_8007,N_4766,N_4217);
or U8008 (N_8008,N_4662,N_5376);
nand U8009 (N_8009,N_7676,N_5310);
xor U8010 (N_8010,N_7383,N_7897);
nand U8011 (N_8011,N_4487,N_5425);
or U8012 (N_8012,N_5980,N_4209);
or U8013 (N_8013,N_7585,N_7004);
xor U8014 (N_8014,N_4201,N_5570);
and U8015 (N_8015,N_5098,N_7410);
or U8016 (N_8016,N_5985,N_4014);
xor U8017 (N_8017,N_4734,N_6469);
or U8018 (N_8018,N_6370,N_6598);
nand U8019 (N_8019,N_6079,N_5208);
nor U8020 (N_8020,N_7871,N_5911);
and U8021 (N_8021,N_6204,N_5486);
and U8022 (N_8022,N_7747,N_5280);
nor U8023 (N_8023,N_7925,N_7673);
or U8024 (N_8024,N_6703,N_5439);
or U8025 (N_8025,N_7868,N_4844);
nand U8026 (N_8026,N_6217,N_6261);
nor U8027 (N_8027,N_7649,N_5424);
or U8028 (N_8028,N_7041,N_4576);
nand U8029 (N_8029,N_7519,N_7730);
and U8030 (N_8030,N_6190,N_7083);
and U8031 (N_8031,N_6872,N_7243);
nor U8032 (N_8032,N_4741,N_4211);
or U8033 (N_8033,N_6048,N_4926);
nor U8034 (N_8034,N_5034,N_5727);
nor U8035 (N_8035,N_7005,N_4649);
nor U8036 (N_8036,N_7028,N_4053);
nand U8037 (N_8037,N_4917,N_4041);
and U8038 (N_8038,N_5437,N_5451);
nand U8039 (N_8039,N_7547,N_6206);
and U8040 (N_8040,N_6482,N_6455);
and U8041 (N_8041,N_6222,N_7505);
and U8042 (N_8042,N_4461,N_5742);
nor U8043 (N_8043,N_6827,N_5772);
and U8044 (N_8044,N_7801,N_6139);
or U8045 (N_8045,N_6306,N_4336);
and U8046 (N_8046,N_4160,N_5796);
and U8047 (N_8047,N_6467,N_7159);
and U8048 (N_8048,N_5074,N_5102);
and U8049 (N_8049,N_6937,N_4470);
nand U8050 (N_8050,N_5542,N_4774);
xor U8051 (N_8051,N_7259,N_5131);
nor U8052 (N_8052,N_6849,N_7589);
or U8053 (N_8053,N_5674,N_4704);
and U8054 (N_8054,N_7966,N_5651);
or U8055 (N_8055,N_5505,N_5368);
nand U8056 (N_8056,N_5285,N_4909);
and U8057 (N_8057,N_7012,N_7638);
and U8058 (N_8058,N_6444,N_6241);
or U8059 (N_8059,N_6745,N_5309);
and U8060 (N_8060,N_7232,N_7467);
nor U8061 (N_8061,N_6046,N_7114);
and U8062 (N_8062,N_7604,N_5400);
or U8063 (N_8063,N_5002,N_6078);
and U8064 (N_8064,N_5971,N_4192);
nand U8065 (N_8065,N_6213,N_5264);
and U8066 (N_8066,N_7003,N_4578);
nor U8067 (N_8067,N_6552,N_5766);
xnor U8068 (N_8068,N_6972,N_7408);
xor U8069 (N_8069,N_4165,N_4894);
and U8070 (N_8070,N_6502,N_4496);
nand U8071 (N_8071,N_4150,N_5601);
xor U8072 (N_8072,N_6735,N_7937);
nand U8073 (N_8073,N_4017,N_5898);
nor U8074 (N_8074,N_5687,N_6181);
nor U8075 (N_8075,N_6295,N_5691);
xor U8076 (N_8076,N_6615,N_7392);
nand U8077 (N_8077,N_7888,N_7054);
nor U8078 (N_8078,N_5694,N_6596);
nand U8079 (N_8079,N_6808,N_6219);
xnor U8080 (N_8080,N_5224,N_4412);
or U8081 (N_8081,N_5793,N_5759);
xor U8082 (N_8082,N_5914,N_4686);
nand U8083 (N_8083,N_4982,N_6053);
nor U8084 (N_8084,N_7065,N_6129);
nor U8085 (N_8085,N_4203,N_5352);
or U8086 (N_8086,N_6947,N_5315);
or U8087 (N_8087,N_5711,N_7636);
or U8088 (N_8088,N_6863,N_4543);
nand U8089 (N_8089,N_6030,N_4376);
and U8090 (N_8090,N_6700,N_4589);
nand U8091 (N_8091,N_5036,N_7103);
nor U8092 (N_8092,N_6413,N_5426);
xnor U8093 (N_8093,N_4719,N_7430);
or U8094 (N_8094,N_7353,N_4657);
and U8095 (N_8095,N_7279,N_7541);
or U8096 (N_8096,N_5108,N_4436);
xor U8097 (N_8097,N_7149,N_4912);
nor U8098 (N_8098,N_7434,N_7387);
xnor U8099 (N_8099,N_4285,N_6893);
and U8100 (N_8100,N_4433,N_5498);
or U8101 (N_8101,N_5397,N_6476);
or U8102 (N_8102,N_7714,N_6066);
and U8103 (N_8103,N_6389,N_7729);
or U8104 (N_8104,N_4667,N_4904);
nor U8105 (N_8105,N_5761,N_5910);
xor U8106 (N_8106,N_6511,N_7153);
and U8107 (N_8107,N_7380,N_7095);
nand U8108 (N_8108,N_6242,N_4821);
and U8109 (N_8109,N_4976,N_4652);
xnor U8110 (N_8110,N_7664,N_6970);
or U8111 (N_8111,N_5567,N_7652);
and U8112 (N_8112,N_7704,N_4930);
nor U8113 (N_8113,N_7378,N_5341);
nand U8114 (N_8114,N_4591,N_6178);
nand U8115 (N_8115,N_6299,N_6918);
nand U8116 (N_8116,N_6479,N_4881);
nor U8117 (N_8117,N_4590,N_4730);
nor U8118 (N_8118,N_4922,N_5681);
nand U8119 (N_8119,N_7366,N_7337);
or U8120 (N_8120,N_5475,N_7677);
xnor U8121 (N_8121,N_6080,N_5906);
xnor U8122 (N_8122,N_4274,N_6378);
nand U8123 (N_8123,N_6730,N_6161);
nand U8124 (N_8124,N_5948,N_4480);
xnor U8125 (N_8125,N_5398,N_5013);
or U8126 (N_8126,N_4036,N_6009);
or U8127 (N_8127,N_5062,N_4365);
nor U8128 (N_8128,N_7863,N_5647);
or U8129 (N_8129,N_5859,N_5555);
nand U8130 (N_8130,N_5808,N_6957);
xnor U8131 (N_8131,N_6949,N_4573);
or U8132 (N_8132,N_6092,N_7835);
nand U8133 (N_8133,N_7064,N_6198);
or U8134 (N_8134,N_7039,N_4987);
xor U8135 (N_8135,N_6977,N_5695);
and U8136 (N_8136,N_7423,N_4527);
nor U8137 (N_8137,N_6857,N_5129);
and U8138 (N_8138,N_6096,N_5493);
xnor U8139 (N_8139,N_5938,N_6240);
and U8140 (N_8140,N_6343,N_4561);
or U8141 (N_8141,N_7424,N_6047);
nor U8142 (N_8142,N_4369,N_6706);
and U8143 (N_8143,N_4549,N_5223);
nand U8144 (N_8144,N_6817,N_7379);
and U8145 (N_8145,N_7246,N_4528);
nor U8146 (N_8146,N_4236,N_6400);
nor U8147 (N_8147,N_6226,N_4373);
or U8148 (N_8148,N_5130,N_5693);
and U8149 (N_8149,N_6074,N_4843);
or U8150 (N_8150,N_5631,N_4037);
nand U8151 (N_8151,N_5125,N_6811);
and U8152 (N_8152,N_7557,N_7503);
nor U8153 (N_8153,N_5239,N_4532);
or U8154 (N_8154,N_7463,N_6787);
nand U8155 (N_8155,N_6646,N_6355);
or U8156 (N_8156,N_5586,N_5629);
nand U8157 (N_8157,N_4749,N_4378);
nand U8158 (N_8158,N_4009,N_6890);
nor U8159 (N_8159,N_5816,N_4712);
nor U8160 (N_8160,N_4295,N_6589);
and U8161 (N_8161,N_4700,N_7139);
nand U8162 (N_8162,N_4238,N_5669);
nor U8163 (N_8163,N_5620,N_4032);
or U8164 (N_8164,N_4568,N_7110);
and U8165 (N_8165,N_7174,N_4331);
nand U8166 (N_8166,N_4050,N_4610);
nor U8167 (N_8167,N_6256,N_4880);
nor U8168 (N_8168,N_7521,N_6326);
nand U8169 (N_8169,N_4232,N_6799);
or U8170 (N_8170,N_6304,N_6889);
or U8171 (N_8171,N_4316,N_5641);
or U8172 (N_8172,N_7293,N_4212);
nand U8173 (N_8173,N_7875,N_7726);
or U8174 (N_8174,N_4015,N_5010);
or U8175 (N_8175,N_5724,N_5583);
nor U8176 (N_8176,N_5824,N_6776);
nor U8177 (N_8177,N_4494,N_6016);
xnor U8178 (N_8178,N_4191,N_4193);
or U8179 (N_8179,N_5085,N_4508);
nand U8180 (N_8180,N_4617,N_7450);
or U8181 (N_8181,N_6702,N_7839);
nand U8182 (N_8182,N_5494,N_4321);
and U8183 (N_8183,N_5446,N_4335);
or U8184 (N_8184,N_5399,N_5061);
or U8185 (N_8185,N_6900,N_4435);
and U8186 (N_8186,N_6394,N_5119);
and U8187 (N_8187,N_7694,N_6607);
or U8188 (N_8188,N_6846,N_4409);
or U8189 (N_8189,N_5872,N_4577);
or U8190 (N_8190,N_4554,N_6273);
xnor U8191 (N_8191,N_6250,N_4586);
nor U8192 (N_8192,N_4304,N_5060);
xor U8193 (N_8193,N_6435,N_5053);
nand U8194 (N_8194,N_7831,N_7775);
nor U8195 (N_8195,N_7693,N_5884);
and U8196 (N_8196,N_7926,N_5750);
nand U8197 (N_8197,N_7143,N_5500);
nand U8198 (N_8198,N_7513,N_7502);
nand U8199 (N_8199,N_6969,N_5541);
nand U8200 (N_8200,N_4825,N_5605);
nand U8201 (N_8201,N_4449,N_5522);
nand U8202 (N_8202,N_6715,N_4600);
and U8203 (N_8203,N_7335,N_7540);
nor U8204 (N_8204,N_4608,N_7130);
and U8205 (N_8205,N_4643,N_6763);
or U8206 (N_8206,N_6524,N_5762);
and U8207 (N_8207,N_4557,N_5679);
xnor U8208 (N_8208,N_5178,N_5283);
or U8209 (N_8209,N_4640,N_4934);
nor U8210 (N_8210,N_7940,N_7556);
and U8211 (N_8211,N_6627,N_6556);
nand U8212 (N_8212,N_7523,N_4445);
or U8213 (N_8213,N_4563,N_5623);
nand U8214 (N_8214,N_7852,N_4382);
nor U8215 (N_8215,N_7218,N_5805);
and U8216 (N_8216,N_5997,N_6574);
nand U8217 (N_8217,N_4984,N_5508);
nand U8218 (N_8218,N_5933,N_7033);
nand U8219 (N_8219,N_7975,N_7819);
and U8220 (N_8220,N_7894,N_7080);
and U8221 (N_8221,N_5875,N_6968);
and U8222 (N_8222,N_4312,N_5356);
and U8223 (N_8223,N_5524,N_7111);
or U8224 (N_8224,N_4899,N_5466);
nand U8225 (N_8225,N_6837,N_7272);
xor U8226 (N_8226,N_5704,N_7990);
or U8227 (N_8227,N_5913,N_4935);
xor U8228 (N_8228,N_7422,N_5552);
nor U8229 (N_8229,N_5929,N_4883);
and U8230 (N_8230,N_5496,N_6407);
and U8231 (N_8231,N_7885,N_5050);
or U8232 (N_8232,N_4342,N_6403);
and U8233 (N_8233,N_5252,N_5560);
and U8234 (N_8234,N_5431,N_5245);
and U8235 (N_8235,N_7264,N_5801);
nor U8236 (N_8236,N_6585,N_6527);
nand U8237 (N_8237,N_5253,N_7340);
and U8238 (N_8238,N_7498,N_7622);
nor U8239 (N_8239,N_7344,N_6934);
nand U8240 (N_8240,N_7689,N_5829);
nand U8241 (N_8241,N_6133,N_7312);
nor U8242 (N_8242,N_7367,N_5767);
or U8243 (N_8243,N_7560,N_6429);
xor U8244 (N_8244,N_4943,N_4673);
and U8245 (N_8245,N_6713,N_4659);
or U8246 (N_8246,N_7125,N_5465);
nor U8247 (N_8247,N_7466,N_6886);
nand U8248 (N_8248,N_5249,N_6603);
nor U8249 (N_8249,N_6822,N_7240);
and U8250 (N_8250,N_7323,N_5456);
nor U8251 (N_8251,N_5643,N_7511);
nor U8252 (N_8252,N_6657,N_6835);
nand U8253 (N_8253,N_7811,N_4020);
nand U8254 (N_8254,N_7286,N_4101);
xor U8255 (N_8255,N_4395,N_4126);
nor U8256 (N_8256,N_6126,N_4998);
nor U8257 (N_8257,N_6392,N_4961);
xnor U8258 (N_8258,N_6123,N_5683);
nand U8259 (N_8259,N_7461,N_7950);
or U8260 (N_8260,N_5656,N_7550);
and U8261 (N_8261,N_7883,N_6506);
nand U8262 (N_8262,N_5891,N_6254);
and U8263 (N_8263,N_5530,N_6543);
nand U8264 (N_8264,N_4245,N_5210);
and U8265 (N_8265,N_7204,N_4383);
nand U8266 (N_8266,N_6354,N_4227);
nand U8267 (N_8267,N_5383,N_4744);
nor U8268 (N_8268,N_6288,N_7128);
nor U8269 (N_8269,N_4776,N_6493);
xnor U8270 (N_8270,N_5680,N_4098);
xnor U8271 (N_8271,N_5395,N_5696);
or U8272 (N_8272,N_7766,N_6866);
or U8273 (N_8273,N_4251,N_6922);
xnor U8274 (N_8274,N_5030,N_5168);
and U8275 (N_8275,N_5489,N_4672);
and U8276 (N_8276,N_4742,N_7668);
or U8277 (N_8277,N_4629,N_6581);
or U8278 (N_8278,N_6514,N_5518);
and U8279 (N_8279,N_4911,N_5664);
or U8280 (N_8280,N_4124,N_4398);
nand U8281 (N_8281,N_7138,N_5423);
nor U8282 (N_8282,N_5877,N_7632);
nand U8283 (N_8283,N_5177,N_6002);
nand U8284 (N_8284,N_7749,N_6451);
nand U8285 (N_8285,N_5271,N_4340);
and U8286 (N_8286,N_7119,N_4454);
nand U8287 (N_8287,N_5499,N_4186);
or U8288 (N_8288,N_6914,N_5721);
nor U8289 (N_8289,N_7844,N_7317);
or U8290 (N_8290,N_4856,N_7180);
or U8291 (N_8291,N_4018,N_6928);
nor U8292 (N_8292,N_5257,N_5749);
and U8293 (N_8293,N_5051,N_5211);
nand U8294 (N_8294,N_6069,N_5783);
or U8295 (N_8295,N_4003,N_5026);
nor U8296 (N_8296,N_7024,N_6879);
nand U8297 (N_8297,N_4136,N_7186);
and U8298 (N_8298,N_7815,N_4641);
and U8299 (N_8299,N_4351,N_5232);
nand U8300 (N_8300,N_5983,N_7440);
nor U8301 (N_8301,N_5764,N_7332);
xnor U8302 (N_8302,N_7501,N_4143);
and U8303 (N_8303,N_6829,N_4684);
nand U8304 (N_8304,N_5106,N_6120);
or U8305 (N_8305,N_6437,N_4394);
nand U8306 (N_8306,N_6194,N_6619);
and U8307 (N_8307,N_4424,N_5588);
xnor U8308 (N_8308,N_7938,N_6741);
nand U8309 (N_8309,N_6023,N_4613);
or U8310 (N_8310,N_7362,N_5012);
or U8311 (N_8311,N_7961,N_6117);
or U8312 (N_8312,N_7487,N_6932);
nor U8313 (N_8313,N_7862,N_5305);
and U8314 (N_8314,N_4747,N_6712);
nand U8315 (N_8315,N_7132,N_6399);
nor U8316 (N_8316,N_6082,N_5219);
nor U8317 (N_8317,N_4208,N_5327);
and U8318 (N_8318,N_5752,N_7027);
or U8319 (N_8319,N_5460,N_7697);
or U8320 (N_8320,N_6224,N_5375);
nand U8321 (N_8321,N_6854,N_4927);
nand U8322 (N_8322,N_7349,N_6992);
nor U8323 (N_8323,N_4172,N_4220);
nand U8324 (N_8324,N_6523,N_7731);
nand U8325 (N_8325,N_6460,N_4465);
nor U8326 (N_8326,N_7623,N_7405);
or U8327 (N_8327,N_4016,N_6107);
nand U8328 (N_8328,N_5369,N_6771);
and U8329 (N_8329,N_7529,N_6954);
or U8330 (N_8330,N_6953,N_5093);
and U8331 (N_8331,N_5322,N_6233);
nand U8332 (N_8332,N_7816,N_6522);
nor U8333 (N_8333,N_4829,N_4145);
and U8334 (N_8334,N_7545,N_4088);
or U8335 (N_8335,N_7266,N_4469);
or U8336 (N_8336,N_7055,N_5353);
xnor U8337 (N_8337,N_6601,N_4345);
nor U8338 (N_8338,N_6475,N_4417);
and U8339 (N_8339,N_6363,N_6673);
or U8340 (N_8340,N_7842,N_5844);
xnor U8341 (N_8341,N_4127,N_5422);
nor U8342 (N_8342,N_7220,N_4505);
or U8343 (N_8343,N_5385,N_5066);
and U8344 (N_8344,N_5506,N_5896);
and U8345 (N_8345,N_5757,N_5078);
nand U8346 (N_8346,N_7479,N_7754);
or U8347 (N_8347,N_7600,N_4552);
nor U8348 (N_8348,N_7867,N_4773);
nor U8349 (N_8349,N_7203,N_7887);
nor U8350 (N_8350,N_7102,N_4807);
xor U8351 (N_8351,N_7850,N_4390);
or U8352 (N_8352,N_6832,N_5531);
and U8353 (N_8353,N_6518,N_6975);
or U8354 (N_8354,N_5421,N_4711);
and U8355 (N_8355,N_7206,N_6892);
nor U8356 (N_8356,N_7598,N_7963);
or U8357 (N_8357,N_7251,N_7849);
or U8358 (N_8358,N_4462,N_5165);
or U8359 (N_8359,N_5449,N_6590);
nand U8360 (N_8360,N_5418,N_7445);
nand U8361 (N_8361,N_5110,N_5254);
xor U8362 (N_8362,N_4778,N_4913);
and U8363 (N_8363,N_4428,N_4655);
or U8364 (N_8364,N_4426,N_4787);
nor U8365 (N_8365,N_4518,N_7592);
or U8366 (N_8366,N_5458,N_7346);
nor U8367 (N_8367,N_6788,N_5912);
nand U8368 (N_8368,N_7280,N_6999);
nor U8369 (N_8369,N_7235,N_4474);
or U8370 (N_8370,N_5337,N_6350);
nor U8371 (N_8371,N_6247,N_5135);
and U8372 (N_8372,N_4703,N_6510);
and U8373 (N_8373,N_7277,N_5049);
and U8374 (N_8374,N_6790,N_4099);
nor U8375 (N_8375,N_5908,N_4109);
or U8376 (N_8376,N_4955,N_7091);
nor U8377 (N_8377,N_4890,N_5540);
xor U8378 (N_8378,N_5788,N_4258);
nor U8379 (N_8379,N_5291,N_4010);
nand U8380 (N_8380,N_7735,N_7696);
nand U8381 (N_8381,N_5006,N_7603);
and U8382 (N_8382,N_5768,N_7207);
or U8383 (N_8383,N_7921,N_6798);
nor U8384 (N_8384,N_4420,N_4653);
nor U8385 (N_8385,N_5846,N_5441);
or U8386 (N_8386,N_7758,N_4607);
and U8387 (N_8387,N_5199,N_5529);
xor U8388 (N_8388,N_5220,N_6061);
xnor U8389 (N_8389,N_7258,N_7588);
and U8390 (N_8390,N_4560,N_6236);
and U8391 (N_8391,N_6653,N_7916);
nor U8392 (N_8392,N_7167,N_4254);
or U8393 (N_8393,N_4635,N_6157);
nand U8394 (N_8394,N_6809,N_6324);
nand U8395 (N_8395,N_5577,N_7559);
nor U8396 (N_8396,N_7645,N_4519);
nand U8397 (N_8397,N_5833,N_7106);
nor U8398 (N_8398,N_5765,N_5373);
nand U8399 (N_8399,N_7173,N_7384);
xnor U8400 (N_8400,N_4928,N_6752);
or U8401 (N_8401,N_6642,N_4111);
nor U8402 (N_8402,N_6680,N_6780);
xor U8403 (N_8403,N_6985,N_6500);
and U8404 (N_8404,N_5642,N_4938);
and U8405 (N_8405,N_7049,N_4065);
nor U8406 (N_8406,N_6310,N_6095);
or U8407 (N_8407,N_5281,N_5532);
and U8408 (N_8408,N_6372,N_6320);
xnor U8409 (N_8409,N_7647,N_5430);
nor U8410 (N_8410,N_5951,N_6568);
or U8411 (N_8411,N_4141,N_5815);
and U8412 (N_8412,N_5706,N_6628);
nand U8413 (N_8413,N_4688,N_6472);
xnor U8414 (N_8414,N_6176,N_7909);
nand U8415 (N_8415,N_4805,N_4030);
or U8416 (N_8416,N_5472,N_6941);
xnor U8417 (N_8417,N_4968,N_7767);
nand U8418 (N_8418,N_5622,N_4860);
nand U8419 (N_8419,N_7542,N_7152);
and U8420 (N_8420,N_7789,N_5650);
or U8421 (N_8421,N_7584,N_7047);
and U8422 (N_8422,N_4222,N_7299);
nor U8423 (N_8423,N_7752,N_6575);
nor U8424 (N_8424,N_5289,N_4503);
nand U8425 (N_8425,N_7462,N_7241);
nor U8426 (N_8426,N_4797,N_5247);
nand U8427 (N_8427,N_7575,N_4991);
or U8428 (N_8428,N_7973,N_4978);
nand U8429 (N_8429,N_4658,N_6498);
nor U8430 (N_8430,N_4178,N_5412);
xor U8431 (N_8431,N_6022,N_6132);
nor U8432 (N_8432,N_6387,N_4895);
xnor U8433 (N_8433,N_4246,N_4966);
or U8434 (N_8434,N_7201,N_7341);
nor U8435 (N_8435,N_6051,N_6263);
nand U8436 (N_8436,N_5056,N_4089);
nand U8437 (N_8437,N_4674,N_4215);
xnor U8438 (N_8438,N_5151,N_6731);
or U8439 (N_8439,N_7653,N_4651);
nand U8440 (N_8440,N_6396,N_7998);
and U8441 (N_8441,N_4034,N_5660);
or U8442 (N_8442,N_7528,N_4451);
xor U8443 (N_8443,N_5944,N_4497);
and U8444 (N_8444,N_4319,N_4594);
xnor U8445 (N_8445,N_4828,N_5081);
and U8446 (N_8446,N_7724,N_6077);
and U8447 (N_8447,N_6447,N_6150);
xor U8448 (N_8448,N_5578,N_6920);
nor U8449 (N_8449,N_4213,N_4931);
and U8450 (N_8450,N_7316,N_5616);
or U8451 (N_8451,N_7932,N_6216);
nor U8452 (N_8452,N_4153,N_4870);
and U8453 (N_8453,N_7891,N_5744);
and U8454 (N_8454,N_5909,N_6828);
nor U8455 (N_8455,N_5094,N_5539);
nor U8456 (N_8456,N_4087,N_6988);
nor U8457 (N_8457,N_6774,N_7869);
nor U8458 (N_8458,N_4423,N_4252);
or U8459 (N_8459,N_4362,N_5045);
nor U8460 (N_8460,N_5420,N_5836);
and U8461 (N_8461,N_5003,N_6245);
nor U8462 (N_8462,N_5546,N_5668);
nand U8463 (N_8463,N_7935,N_4743);
nand U8464 (N_8464,N_5890,N_7942);
or U8465 (N_8465,N_6909,N_5100);
nand U8466 (N_8466,N_6595,N_6088);
and U8467 (N_8467,N_6979,N_4079);
xor U8468 (N_8468,N_6094,N_7746);
nor U8469 (N_8469,N_4598,N_4841);
nor U8470 (N_8470,N_5038,N_4415);
or U8471 (N_8471,N_5134,N_7976);
nand U8472 (N_8472,N_7886,N_6667);
nor U8473 (N_8473,N_5477,N_4767);
nand U8474 (N_8474,N_5543,N_6661);
xnor U8475 (N_8475,N_7859,N_7309);
and U8476 (N_8476,N_4393,N_4775);
xor U8477 (N_8477,N_4863,N_4366);
nand U8478 (N_8478,N_7401,N_6772);
or U8479 (N_8479,N_4156,N_7257);
nand U8480 (N_8480,N_7491,N_5454);
xnor U8481 (N_8481,N_7856,N_5720);
xor U8482 (N_8482,N_5996,N_5348);
nand U8483 (N_8483,N_5854,N_4375);
and U8484 (N_8484,N_6065,N_5812);
and U8485 (N_8485,N_5777,N_7101);
or U8486 (N_8486,N_7113,N_6470);
nand U8487 (N_8487,N_5473,N_7913);
or U8488 (N_8488,N_5517,N_6209);
and U8489 (N_8489,N_5480,N_7597);
nand U8490 (N_8490,N_4846,N_4592);
nand U8491 (N_8491,N_6411,N_7342);
and U8492 (N_8492,N_5228,N_5099);
and U8493 (N_8493,N_6335,N_6692);
xor U8494 (N_8494,N_4388,N_5046);
and U8495 (N_8495,N_7711,N_4901);
nor U8496 (N_8496,N_4777,N_5994);
nand U8497 (N_8497,N_6235,N_6744);
and U8498 (N_8498,N_7345,N_5700);
and U8499 (N_8499,N_6687,N_4758);
and U8500 (N_8500,N_4862,N_4510);
and U8501 (N_8501,N_6786,N_4471);
and U8502 (N_8502,N_4823,N_4768);
and U8503 (N_8503,N_7605,N_5654);
or U8504 (N_8504,N_4495,N_7046);
or U8505 (N_8505,N_6982,N_4701);
and U8506 (N_8506,N_5163,N_4513);
or U8507 (N_8507,N_7716,N_4897);
or U8508 (N_8508,N_4407,N_6616);
nand U8509 (N_8509,N_4678,N_4332);
nand U8510 (N_8510,N_7452,N_6873);
nor U8511 (N_8511,N_7199,N_5826);
xnor U8512 (N_8512,N_5079,N_6381);
and U8513 (N_8513,N_6751,N_7060);
and U8514 (N_8514,N_5780,N_4205);
nand U8515 (N_8515,N_5853,N_7912);
nand U8516 (N_8516,N_6877,N_7248);
or U8517 (N_8517,N_7732,N_6385);
xnor U8518 (N_8518,N_7594,N_5435);
nand U8519 (N_8519,N_4400,N_7195);
nand U8520 (N_8520,N_7695,N_6175);
nor U8521 (N_8521,N_6946,N_7780);
and U8522 (N_8522,N_7265,N_5296);
xor U8523 (N_8523,N_4764,N_7442);
xnor U8524 (N_8524,N_5428,N_7514);
or U8525 (N_8525,N_4818,N_4371);
nor U8526 (N_8526,N_5784,N_6218);
nor U8527 (N_8527,N_6898,N_6845);
or U8528 (N_8528,N_6212,N_6309);
nand U8529 (N_8529,N_5267,N_4317);
nor U8530 (N_8530,N_7122,N_7037);
and U8531 (N_8531,N_4380,N_6773);
or U8532 (N_8532,N_4174,N_5141);
xor U8533 (N_8533,N_7062,N_6336);
nand U8534 (N_8534,N_5284,N_6609);
nor U8535 (N_8535,N_6365,N_7267);
nor U8536 (N_8536,N_4190,N_7873);
nor U8537 (N_8537,N_5405,N_4602);
nor U8538 (N_8538,N_6622,N_7712);
and U8539 (N_8539,N_6592,N_5029);
nand U8540 (N_8540,N_6227,N_7097);
or U8541 (N_8541,N_7161,N_7786);
nor U8542 (N_8542,N_5071,N_7682);
nor U8543 (N_8543,N_5886,N_6197);
and U8544 (N_8544,N_6101,N_5483);
or U8545 (N_8545,N_5670,N_7978);
nand U8546 (N_8546,N_4798,N_7829);
and U8547 (N_8547,N_4035,N_6529);
nand U8548 (N_8548,N_5262,N_6586);
nand U8549 (N_8549,N_4612,N_4437);
or U8550 (N_8550,N_5297,N_6294);
nor U8551 (N_8551,N_7076,N_6929);
xor U8552 (N_8552,N_7669,N_5171);
xor U8553 (N_8553,N_5946,N_7031);
nor U8554 (N_8554,N_4261,N_4484);
nand U8555 (N_8555,N_7244,N_6602);
xor U8556 (N_8556,N_7373,N_5001);
and U8557 (N_8557,N_6698,N_4240);
and U8558 (N_8558,N_7607,N_6901);
or U8559 (N_8559,N_5024,N_6029);
or U8560 (N_8560,N_4438,N_5653);
or U8561 (N_8561,N_4924,N_7793);
and U8562 (N_8562,N_7471,N_5527);
nand U8563 (N_8563,N_5378,N_7216);
and U8564 (N_8564,N_6073,N_7804);
nand U8565 (N_8565,N_4754,N_5644);
nor U8566 (N_8566,N_5236,N_6050);
nand U8567 (N_8567,N_7959,N_4326);
nand U8568 (N_8568,N_5242,N_6160);
nor U8569 (N_8569,N_6011,N_7838);
and U8570 (N_8570,N_5572,N_6352);
nor U8571 (N_8571,N_5626,N_6419);
or U8572 (N_8572,N_5673,N_4460);
and U8573 (N_8573,N_7782,N_6784);
or U8574 (N_8574,N_5155,N_5039);
nand U8575 (N_8575,N_6265,N_7534);
nor U8576 (N_8576,N_6423,N_5562);
nand U8577 (N_8577,N_5956,N_4442);
and U8578 (N_8578,N_5820,N_4654);
or U8579 (N_8579,N_4827,N_4682);
xnor U8580 (N_8580,N_6923,N_7713);
nor U8581 (N_8581,N_4851,N_5292);
nand U8582 (N_8582,N_7419,N_5963);
nor U8583 (N_8583,N_6944,N_7544);
or U8584 (N_8584,N_4681,N_6055);
or U8585 (N_8585,N_7002,N_6359);
and U8586 (N_8586,N_6689,N_4785);
nor U8587 (N_8587,N_7233,N_5382);
nand U8588 (N_8588,N_4656,N_5959);
nor U8589 (N_8589,N_7360,N_6572);
or U8590 (N_8590,N_5717,N_7517);
nand U8591 (N_8591,N_4338,N_4914);
xor U8592 (N_8592,N_6577,N_4889);
nand U8593 (N_8593,N_5625,N_5528);
and U8594 (N_8594,N_4865,N_7256);
and U8595 (N_8595,N_5358,N_5665);
or U8596 (N_8596,N_4339,N_6571);
xor U8597 (N_8597,N_7198,N_5014);
and U8598 (N_8598,N_5127,N_6777);
nor U8599 (N_8599,N_4314,N_7032);
and U8600 (N_8600,N_7438,N_6438);
xor U8601 (N_8601,N_7146,N_5710);
nand U8602 (N_8602,N_7627,N_4562);
nand U8603 (N_8603,N_5878,N_4452);
and U8604 (N_8604,N_5175,N_4679);
and U8605 (N_8605,N_4206,N_4918);
nor U8606 (N_8606,N_7289,N_7977);
nand U8607 (N_8607,N_7795,N_7160);
nor U8608 (N_8608,N_7563,N_7347);
and U8609 (N_8609,N_6532,N_7577);
or U8610 (N_8610,N_4980,N_5697);
or U8611 (N_8611,N_6733,N_5748);
or U8612 (N_8612,N_5390,N_7035);
and U8613 (N_8613,N_7176,N_5104);
and U8614 (N_8614,N_4490,N_5417);
or U8615 (N_8615,N_6885,N_5408);
or U8616 (N_8616,N_7680,N_6664);
or U8617 (N_8617,N_4642,N_6495);
nand U8618 (N_8618,N_5955,N_7967);
xor U8619 (N_8619,N_7791,N_6349);
or U8620 (N_8620,N_7325,N_4886);
nand U8621 (N_8621,N_5429,N_5241);
nor U8622 (N_8622,N_7276,N_7929);
nand U8623 (N_8623,N_4275,N_7812);
nand U8624 (N_8624,N_4139,N_6563);
or U8625 (N_8625,N_7659,N_5666);
nand U8626 (N_8626,N_6880,N_6547);
xor U8627 (N_8627,N_6329,N_6168);
and U8628 (N_8628,N_6277,N_4107);
and U8629 (N_8629,N_6305,N_5709);
nand U8630 (N_8630,N_5350,N_4812);
nor U8631 (N_8631,N_5927,N_5040);
and U8632 (N_8632,N_4757,N_5713);
xnor U8633 (N_8633,N_4293,N_4855);
nor U8634 (N_8634,N_7701,N_6405);
xnor U8635 (N_8635,N_6478,N_4905);
xor U8636 (N_8636,N_6545,N_4128);
nor U8637 (N_8637,N_7639,N_6450);
or U8638 (N_8638,N_6537,N_7372);
nand U8639 (N_8639,N_5025,N_6155);
and U8640 (N_8640,N_7483,N_7288);
or U8641 (N_8641,N_4604,N_7982);
nor U8642 (N_8642,N_7320,N_5302);
or U8643 (N_8643,N_6318,N_4915);
xor U8644 (N_8644,N_4108,N_4811);
or U8645 (N_8645,N_7104,N_5101);
nor U8646 (N_8646,N_7770,N_4921);
nand U8647 (N_8647,N_6116,N_6754);
nand U8648 (N_8648,N_4695,N_5004);
and U8649 (N_8649,N_5502,N_7756);
nand U8650 (N_8650,N_7089,N_5781);
xnor U8651 (N_8651,N_5244,N_7561);
nor U8652 (N_8652,N_7426,N_6666);
xnor U8653 (N_8653,N_7646,N_4761);
or U8654 (N_8654,N_5640,N_6587);
nand U8655 (N_8655,N_4832,N_5326);
nor U8656 (N_8656,N_7136,N_7084);
and U8657 (N_8657,N_4992,N_6508);
or U8658 (N_8658,N_7036,N_5892);
or U8659 (N_8659,N_4368,N_4944);
nand U8660 (N_8660,N_7406,N_5162);
and U8661 (N_8661,N_4802,N_7882);
or U8662 (N_8662,N_4511,N_7040);
xnor U8663 (N_8663,N_7115,N_4012);
or U8664 (N_8664,N_6442,N_4029);
nand U8665 (N_8665,N_5196,N_7070);
and U8666 (N_8666,N_4218,N_4949);
nand U8667 (N_8667,N_5690,N_6743);
xnor U8668 (N_8668,N_5834,N_6823);
nand U8669 (N_8669,N_6330,N_7352);
or U8670 (N_8670,N_7229,N_7494);
nor U8671 (N_8671,N_7404,N_5814);
nor U8672 (N_8672,N_5054,N_6704);
nor U8673 (N_8673,N_4733,N_5514);
nor U8674 (N_8674,N_7700,N_5159);
xor U8675 (N_8675,N_4675,N_5516);
nor U8676 (N_8676,N_7889,N_7007);
nand U8677 (N_8677,N_4180,N_5342);
nor U8678 (N_8678,N_6497,N_5952);
and U8679 (N_8679,N_4699,N_5467);
nor U8680 (N_8680,N_5627,N_6007);
nand U8681 (N_8681,N_5675,N_7145);
or U8682 (N_8682,N_5649,N_6404);
nor U8683 (N_8683,N_6183,N_6542);
nand U8684 (N_8684,N_7364,N_6262);
or U8685 (N_8685,N_5158,N_4707);
nand U8686 (N_8686,N_7063,N_7045);
nand U8687 (N_8687,N_4241,N_7823);
nor U8688 (N_8688,N_4066,N_7310);
xor U8689 (N_8689,N_6331,N_6477);
and U8690 (N_8690,N_4748,N_6274);
nand U8691 (N_8691,N_7000,N_4396);
or U8692 (N_8692,N_6848,N_7492);
and U8693 (N_8693,N_6010,N_4455);
nor U8694 (N_8694,N_5027,N_5188);
nor U8695 (N_8695,N_7088,N_6709);
or U8696 (N_8696,N_6913,N_4788);
and U8697 (N_8697,N_7361,N_5402);
and U8698 (N_8698,N_6054,N_4830);
nor U8699 (N_8699,N_4873,N_7595);
or U8700 (N_8700,N_5538,N_4164);
nor U8701 (N_8701,N_6149,N_5987);
and U8702 (N_8702,N_5970,N_5549);
and U8703 (N_8703,N_4584,N_5258);
nor U8704 (N_8704,N_5133,N_7774);
nor U8705 (N_8705,N_7722,N_4305);
xnor U8706 (N_8706,N_7910,N_7393);
nor U8707 (N_8707,N_7641,N_5981);
nor U8708 (N_8708,N_4406,N_4683);
xor U8709 (N_8709,N_5116,N_4159);
nand U8710 (N_8710,N_5655,N_7635);
or U8711 (N_8711,N_7314,N_6067);
and U8712 (N_8712,N_5563,N_5589);
and U8713 (N_8713,N_4962,N_7470);
or U8714 (N_8714,N_4936,N_6630);
xnor U8715 (N_8715,N_5734,N_4954);
nand U8716 (N_8716,N_5120,N_4131);
xor U8717 (N_8717,N_5894,N_5349);
nand U8718 (N_8718,N_6087,N_6440);
or U8719 (N_8719,N_7565,N_7099);
nor U8720 (N_8720,N_4611,N_4708);
or U8721 (N_8721,N_6279,N_7650);
or U8722 (N_8722,N_4199,N_7141);
and U8723 (N_8723,N_4387,N_7611);
xnor U8724 (N_8724,N_6422,N_5556);
nor U8725 (N_8725,N_6426,N_4637);
nor U8726 (N_8726,N_4509,N_6764);
or U8727 (N_8727,N_7262,N_6638);
or U8728 (N_8728,N_5052,N_7144);
nand U8729 (N_8729,N_4219,N_5550);
or U8730 (N_8730,N_4411,N_5364);
nand U8731 (N_8731,N_6807,N_6593);
nand U8732 (N_8732,N_6028,N_6463);
or U8733 (N_8733,N_5969,N_6639);
nand U8734 (N_8734,N_4808,N_4374);
and U8735 (N_8735,N_6099,N_6468);
nor U8736 (N_8736,N_7023,N_7992);
nor U8737 (N_8737,N_6834,N_4660);
nor U8738 (N_8738,N_7609,N_6674);
xnor U8739 (N_8739,N_5278,N_5090);
nand U8740 (N_8740,N_4166,N_4049);
xnor U8741 (N_8741,N_6555,N_4771);
or U8742 (N_8742,N_4148,N_6041);
and U8743 (N_8743,N_5314,N_6814);
xor U8744 (N_8744,N_7158,N_6738);
and U8745 (N_8745,N_6042,N_7796);
xnor U8746 (N_8746,N_5712,N_6496);
nand U8747 (N_8747,N_7954,N_7918);
or U8748 (N_8748,N_4363,N_6933);
nand U8749 (N_8749,N_7516,N_7817);
nand U8750 (N_8750,N_7411,N_5198);
and U8751 (N_8751,N_6690,N_4323);
xor U8752 (N_8752,N_6714,N_5126);
and U8753 (N_8753,N_6635,N_5229);
nand U8754 (N_8754,N_5624,N_6912);
and U8755 (N_8755,N_6152,N_7902);
and U8756 (N_8756,N_5063,N_6253);
nand U8757 (N_8757,N_5065,N_4671);
nor U8758 (N_8758,N_6662,N_4155);
and U8759 (N_8759,N_7029,N_6271);
xor U8760 (N_8760,N_7338,N_4489);
nand U8761 (N_8761,N_5822,N_4281);
nand U8762 (N_8762,N_7318,N_7348);
and U8763 (N_8763,N_5485,N_6064);
nand U8764 (N_8764,N_6297,N_4072);
nor U8765 (N_8765,N_5708,N_7798);
and U8766 (N_8766,N_5637,N_4443);
xor U8767 (N_8767,N_6998,N_6724);
xor U8768 (N_8768,N_5918,N_7285);
and U8769 (N_8769,N_6225,N_6943);
nand U8770 (N_8770,N_7717,N_7779);
and U8771 (N_8771,N_4769,N_4491);
nor U8772 (N_8772,N_5411,N_6765);
nor U8773 (N_8773,N_7090,N_7539);
xor U8774 (N_8774,N_6565,N_5379);
xnor U8775 (N_8775,N_5355,N_6539);
nor U8776 (N_8776,N_6756,N_7154);
or U8777 (N_8777,N_4981,N_6516);
nor U8778 (N_8778,N_4432,N_5321);
nor U8779 (N_8779,N_7326,N_4260);
or U8780 (N_8780,N_7305,N_4103);
or U8781 (N_8781,N_5190,N_4106);
or U8782 (N_8782,N_4539,N_6815);
or U8783 (N_8783,N_4439,N_7803);
xnor U8784 (N_8784,N_6075,N_7018);
xor U8785 (N_8785,N_6221,N_4063);
xor U8786 (N_8786,N_6201,N_7200);
or U8787 (N_8787,N_4350,N_5835);
nor U8788 (N_8788,N_4669,N_4188);
or U8789 (N_8789,N_6110,N_7489);
and U8790 (N_8790,N_6140,N_7184);
and U8791 (N_8791,N_6312,N_6973);
and U8792 (N_8792,N_5924,N_5943);
and U8793 (N_8793,N_6237,N_5887);
and U8794 (N_8794,N_4882,N_7828);
and U8795 (N_8795,N_4698,N_4551);
or U8796 (N_8796,N_4603,N_4054);
nor U8797 (N_8797,N_4132,N_4919);
nor U8798 (N_8798,N_6801,N_6749);
and U8799 (N_8799,N_4043,N_6471);
nor U8800 (N_8800,N_6736,N_4402);
nor U8801 (N_8801,N_4548,N_6800);
and U8802 (N_8802,N_6321,N_7656);
nand U8803 (N_8803,N_7327,N_4318);
nand U8804 (N_8804,N_5621,N_6169);
or U8805 (N_8805,N_4879,N_5202);
or U8806 (N_8806,N_4125,N_4997);
nand U8807 (N_8807,N_4303,N_5414);
and U8808 (N_8808,N_4075,N_6384);
or U8809 (N_8809,N_4685,N_7371);
or U8810 (N_8810,N_6416,N_4750);
nor U8811 (N_8811,N_6353,N_7269);
and U8812 (N_8812,N_4421,N_4225);
nor U8813 (N_8813,N_6259,N_5212);
or U8814 (N_8814,N_5317,N_6308);
nand U8815 (N_8815,N_6833,N_5299);
and U8816 (N_8816,N_6582,N_7051);
or U8817 (N_8817,N_7117,N_7147);
and U8818 (N_8818,N_5839,N_5023);
nand U8819 (N_8819,N_4114,N_4320);
nor U8820 (N_8820,N_6856,N_7193);
nor U8821 (N_8821,N_7832,N_4440);
nor U8822 (N_8822,N_5070,N_4392);
and U8823 (N_8823,N_6255,N_4173);
xnor U8824 (N_8824,N_7596,N_5343);
nand U8825 (N_8825,N_4204,N_7997);
nor U8826 (N_8826,N_7944,N_4477);
nor U8827 (N_8827,N_7127,N_6813);
xnor U8828 (N_8828,N_7126,N_5607);
or U8829 (N_8829,N_5686,N_6040);
nor U8830 (N_8830,N_6436,N_6474);
nor U8831 (N_8831,N_5722,N_6171);
and U8832 (N_8832,N_6177,N_6382);
and U8833 (N_8833,N_7930,N_5707);
and U8834 (N_8834,N_7190,N_7183);
nand U8835 (N_8835,N_4697,N_4187);
nand U8836 (N_8836,N_6351,N_4910);
xnor U8837 (N_8837,N_4078,N_6927);
and U8838 (N_8838,N_7939,N_7415);
xnor U8839 (N_8839,N_7417,N_7537);
xnor U8840 (N_8840,N_7602,N_4547);
and U8841 (N_8841,N_4906,N_6819);
xor U8842 (N_8842,N_6904,N_6043);
nor U8843 (N_8843,N_6559,N_6488);
or U8844 (N_8844,N_4024,N_4616);
nand U8845 (N_8845,N_4121,N_5658);
and U8846 (N_8846,N_7441,N_6267);
or U8847 (N_8847,N_6825,N_7994);
or U8848 (N_8848,N_4171,N_5057);
nand U8849 (N_8849,N_4272,N_6348);
and U8850 (N_8850,N_7249,N_5497);
xnor U8851 (N_8851,N_5684,N_6513);
nand U8852 (N_8852,N_4524,N_7608);
nor U8853 (N_8853,N_5756,N_6186);
and U8854 (N_8854,N_6643,N_5786);
nor U8855 (N_8855,N_6390,N_7311);
xor U8856 (N_8856,N_4207,N_7618);
nand U8857 (N_8857,N_5215,N_6368);
or U8858 (N_8858,N_7014,N_5097);
nand U8859 (N_8859,N_5581,N_5410);
nand U8860 (N_8860,N_4986,N_5774);
or U8861 (N_8861,N_7790,N_5048);
and U8862 (N_8862,N_7477,N_6280);
and U8863 (N_8863,N_4278,N_4718);
nand U8864 (N_8864,N_4263,N_5170);
and U8865 (N_8865,N_7788,N_6930);
nor U8866 (N_8866,N_5525,N_7368);
xnor U8867 (N_8867,N_6211,N_7086);
nand U8868 (N_8868,N_6239,N_5718);
nand U8869 (N_8869,N_4623,N_5316);
nor U8870 (N_8870,N_4687,N_7543);
nor U8871 (N_8871,N_6882,N_5347);
nand U8872 (N_8872,N_7739,N_7020);
and U8873 (N_8873,N_7826,N_4115);
or U8874 (N_8874,N_5359,N_6311);
and U8875 (N_8875,N_5633,N_6141);
nand U8876 (N_8876,N_7861,N_7237);
nand U8877 (N_8877,N_4322,N_4792);
or U8878 (N_8878,N_6371,N_4858);
xor U8879 (N_8879,N_5501,N_7599);
nand U8880 (N_8880,N_6705,N_5973);
and U8881 (N_8881,N_5180,N_5300);
and U8882 (N_8882,N_6089,N_6098);
nand U8883 (N_8883,N_6505,N_5982);
and U8884 (N_8884,N_7753,N_4726);
xor U8885 (N_8885,N_5282,N_5088);
and U8886 (N_8886,N_5445,N_5075);
nand U8887 (N_8887,N_4110,N_5448);
nor U8888 (N_8888,N_7586,N_4550);
nor U8889 (N_8889,N_7333,N_7112);
and U8890 (N_8890,N_7987,N_7116);
nand U8891 (N_8891,N_6701,N_5810);
nor U8892 (N_8892,N_5798,N_7294);
or U8893 (N_8893,N_7252,N_7999);
xor U8894 (N_8894,N_5068,N_4826);
and U8895 (N_8895,N_6081,N_5672);
nand U8896 (N_8896,N_4796,N_5251);
nor U8897 (N_8897,N_7633,N_5789);
nand U8898 (N_8898,N_5139,N_7551);
nand U8899 (N_8899,N_7566,N_7369);
and U8900 (N_8900,N_6483,N_5406);
nor U8901 (N_8901,N_5009,N_7740);
and U8902 (N_8902,N_6249,N_5827);
or U8903 (N_8903,N_7443,N_7074);
or U8904 (N_8904,N_4973,N_6675);
and U8905 (N_8905,N_5962,N_4933);
nand U8906 (N_8906,N_4294,N_6446);
xor U8907 (N_8907,N_6401,N_6884);
nand U8908 (N_8908,N_7260,N_5802);
or U8909 (N_8909,N_5746,N_5113);
xor U8910 (N_8910,N_7324,N_5263);
nand U8911 (N_8911,N_6182,N_5866);
and U8912 (N_8912,N_5974,N_7934);
and U8913 (N_8913,N_5725,N_6991);
or U8914 (N_8914,N_5964,N_4940);
nor U8915 (N_8915,N_7956,N_5832);
and U8916 (N_8916,N_5033,N_6301);
nand U8917 (N_8917,N_5124,N_4062);
nor U8918 (N_8918,N_4725,N_6049);
nor U8919 (N_8919,N_6534,N_7580);
or U8920 (N_8920,N_7382,N_4896);
and U8921 (N_8921,N_6012,N_5519);
or U8922 (N_8922,N_5216,N_7957);
or U8923 (N_8923,N_6269,N_6230);
and U8924 (N_8924,N_7759,N_4290);
xor U8925 (N_8925,N_4908,N_7071);
nor U8926 (N_8926,N_5462,N_5311);
xor U8927 (N_8927,N_7162,N_6597);
and U8928 (N_8928,N_7077,N_5520);
xor U8929 (N_8929,N_7359,N_5574);
or U8930 (N_8930,N_4946,N_4138);
nor U8931 (N_8931,N_4569,N_5977);
and U8932 (N_8932,N_6020,N_7751);
and U8933 (N_8933,N_7810,N_7865);
or U8934 (N_8934,N_5064,N_5966);
and U8935 (N_8935,N_5225,N_5233);
nor U8936 (N_8936,N_4472,N_5059);
nor U8937 (N_8937,N_7847,N_5504);
nand U8938 (N_8938,N_7512,N_7892);
nor U8939 (N_8939,N_5008,N_4994);
nor U8940 (N_8940,N_5357,N_4958);
xor U8941 (N_8941,N_6214,N_5367);
or U8942 (N_8942,N_4264,N_6716);
or U8943 (N_8943,N_4850,N_6660);
or U8944 (N_8944,N_7044,N_6298);
xor U8945 (N_8945,N_7570,N_6083);
and U8946 (N_8946,N_4327,N_5595);
nor U8947 (N_8947,N_4404,N_4056);
nand U8948 (N_8948,N_7273,N_4957);
nor U8949 (N_8949,N_5547,N_6266);
and U8950 (N_8950,N_7674,N_7376);
nor U8951 (N_8951,N_7818,N_6003);
and U8952 (N_8952,N_7402,N_7178);
or U8953 (N_8953,N_6950,N_4296);
nor U8954 (N_8954,N_6490,N_4133);
and U8955 (N_8955,N_5862,N_4343);
nor U8956 (N_8956,N_6432,N_7806);
and U8957 (N_8957,N_6645,N_4975);
xor U8958 (N_8958,N_4869,N_6462);
and U8959 (N_8959,N_6393,N_7834);
nor U8960 (N_8960,N_4073,N_7610);
and U8961 (N_8961,N_4270,N_7313);
or U8962 (N_8962,N_7617,N_5389);
nor U8963 (N_8963,N_4546,N_4479);
or U8964 (N_8964,N_6533,N_5523);
nor U8965 (N_8965,N_6013,N_6789);
and U8966 (N_8966,N_5845,N_7469);
nand U8967 (N_8967,N_4384,N_7073);
nor U8968 (N_8968,N_4529,N_7705);
and U8969 (N_8969,N_6452,N_7590);
nand U8970 (N_8970,N_6441,N_6364);
or U8971 (N_8971,N_4058,N_6388);
or U8972 (N_8972,N_7454,N_5391);
nand U8973 (N_8973,N_4228,N_7969);
nand U8974 (N_8974,N_4130,N_4226);
nor U8975 (N_8975,N_5787,N_5852);
and U8976 (N_8976,N_6418,N_5331);
and U8977 (N_8977,N_7660,N_7807);
and U8978 (N_8978,N_6056,N_6959);
nand U8979 (N_8979,N_6967,N_7958);
nand U8980 (N_8980,N_5603,N_6068);
and U8981 (N_8981,N_7263,N_4330);
and U8982 (N_8982,N_7435,N_6290);
and U8983 (N_8983,N_7508,N_5194);
xor U8984 (N_8984,N_5265,N_6448);
or U8985 (N_8985,N_6844,N_7860);
and U8986 (N_8986,N_6747,N_6838);
nand U8987 (N_8987,N_4837,N_4875);
and U8988 (N_8988,N_4646,N_4670);
nor U8989 (N_8989,N_7890,N_4732);
or U8990 (N_8990,N_6728,N_4372);
and U8991 (N_8991,N_7163,N_7459);
and U8992 (N_8992,N_6688,N_6158);
nor U8993 (N_8993,N_5965,N_4288);
or U8994 (N_8994,N_7093,N_4781);
nand U8995 (N_8995,N_7196,N_6729);
and U8996 (N_8996,N_6640,N_4300);
xor U8997 (N_8997,N_4000,N_4177);
and U8998 (N_8998,N_4647,N_4142);
and U8999 (N_8999,N_6187,N_7460);
nor U9000 (N_9000,N_6865,N_7194);
and U9001 (N_9001,N_6361,N_5899);
nor U9002 (N_9002,N_5580,N_5091);
or U9003 (N_9003,N_6143,N_4990);
and U9004 (N_9004,N_6579,N_4633);
xnor U9005 (N_9005,N_7388,N_7416);
nand U9006 (N_9006,N_6864,N_6449);
nor U9007 (N_9007,N_4620,N_4988);
xor U9008 (N_9008,N_7568,N_5140);
or U9009 (N_9009,N_6578,N_6566);
xor U9010 (N_9010,N_6179,N_4301);
or U9011 (N_9011,N_4729,N_4892);
nand U9012 (N_9012,N_4512,N_6135);
nand U9013 (N_9013,N_6916,N_6208);
or U9014 (N_9014,N_7703,N_7983);
and U9015 (N_9015,N_7583,N_4434);
and U9016 (N_9016,N_6993,N_6238);
xnor U9017 (N_9017,N_6232,N_4483);
nor U9018 (N_9018,N_6895,N_4722);
nor U9019 (N_9019,N_4939,N_5189);
nand U9020 (N_9020,N_4202,N_5867);
nor U9021 (N_9021,N_7308,N_7662);
xnor U9022 (N_9022,N_4069,N_5037);
nand U9023 (N_9023,N_5167,N_6990);
nor U9024 (N_9024,N_6707,N_4614);
xor U9025 (N_9025,N_6272,N_7398);
xor U9026 (N_9026,N_6659,N_5432);
nand U9027 (N_9027,N_4429,N_4249);
or U9028 (N_9028,N_4419,N_7777);
nand U9029 (N_9029,N_7825,N_7157);
xor U9030 (N_9030,N_5998,N_7558);
and U9031 (N_9031,N_7209,N_4266);
nor U9032 (N_9032,N_4622,N_6683);
nor U9033 (N_9033,N_7016,N_6070);
or U9034 (N_9034,N_5841,N_4283);
nor U9035 (N_9035,N_5676,N_4287);
or U9036 (N_9036,N_6782,N_5112);
and U9037 (N_9037,N_7554,N_6205);
xor U9038 (N_9038,N_4714,N_5851);
nand U9039 (N_9039,N_4334,N_4243);
nor U9040 (N_9040,N_7458,N_4255);
nor U9041 (N_9041,N_6397,N_5031);
nor U9042 (N_9042,N_6322,N_4247);
and U9043 (N_9043,N_4628,N_5490);
nor U9044 (N_9044,N_5920,N_5598);
and U9045 (N_9045,N_4152,N_7197);
nor U9046 (N_9046,N_5293,N_5295);
nor U9047 (N_9047,N_7108,N_7291);
or U9048 (N_9048,N_5035,N_6956);
nand U9049 (N_9049,N_7336,N_4575);
nor U9050 (N_9050,N_5646,N_4259);
nand U9051 (N_9051,N_4650,N_5403);
or U9052 (N_9052,N_7737,N_7429);
nor U9053 (N_9053,N_5145,N_4783);
or U9054 (N_9054,N_6021,N_5775);
and U9055 (N_9055,N_4488,N_6357);
nand U9056 (N_9056,N_5021,N_6319);
nand U9057 (N_9057,N_6793,N_6919);
nand U9058 (N_9058,N_7778,N_4353);
and U9059 (N_9059,N_7386,N_4721);
and U9060 (N_9060,N_5677,N_5482);
nand U9061 (N_9061,N_6737,N_6491);
or U9062 (N_9062,N_5464,N_4956);
or U9063 (N_9063,N_6484,N_4057);
and U9064 (N_9064,N_7226,N_6538);
nor U9065 (N_9065,N_6633,N_4195);
nor U9066 (N_9066,N_6130,N_6406);
and U9067 (N_9067,N_6626,N_6052);
and U9068 (N_9068,N_5087,N_6750);
and U9069 (N_9069,N_7945,N_4746);
nand U9070 (N_9070,N_7931,N_4297);
nor U9071 (N_9071,N_5632,N_6026);
nand U9072 (N_9072,N_6410,N_4840);
nand U9073 (N_9073,N_5156,N_4638);
nand U9074 (N_9074,N_4644,N_7268);
nand U9075 (N_9075,N_7001,N_4467);
nand U9076 (N_9076,N_5967,N_5339);
and U9077 (N_9077,N_6869,N_6681);
xnor U9078 (N_9078,N_6734,N_4416);
and U9079 (N_9079,N_5526,N_6034);
and U9080 (N_9080,N_6767,N_6758);
and U9081 (N_9081,N_5602,N_4702);
xnor U9082 (N_9082,N_7688,N_4200);
and U9083 (N_9083,N_4418,N_6521);
or U9084 (N_9084,N_4094,N_7920);
nand U9085 (N_9085,N_6373,N_4540);
xnor U9086 (N_9086,N_5256,N_5157);
xor U9087 (N_9087,N_7391,N_5613);
and U9088 (N_9088,N_7972,N_5457);
nand U9089 (N_9089,N_7480,N_4042);
or U9090 (N_9090,N_5384,N_6118);
nor U9091 (N_9091,N_5888,N_6672);
nor U9092 (N_9092,N_5863,N_5077);
nor U9093 (N_9093,N_6344,N_4515);
and U9094 (N_9094,N_5286,N_4129);
xnor U9095 (N_9095,N_5931,N_7827);
or U9096 (N_9096,N_6826,N_7667);
nand U9097 (N_9097,N_6917,N_5484);
or U9098 (N_9098,N_4803,N_5330);
and U9099 (N_9099,N_4499,N_5273);
or U9100 (N_9100,N_5121,N_6494);
nor U9101 (N_9101,N_6678,N_6485);
xnor U9102 (N_9102,N_5470,N_6443);
and U9103 (N_9103,N_6125,N_4341);
nand U9104 (N_9104,N_5442,N_4349);
nand U9105 (N_9105,N_4780,N_5755);
nand U9106 (N_9106,N_7905,N_7307);
and U9107 (N_9107,N_4408,N_4061);
or U9108 (N_9108,N_7179,N_7390);
nand U9109 (N_9109,N_7606,N_7300);
nor U9110 (N_9110,N_6896,N_7334);
nand U9111 (N_9111,N_5227,N_5396);
nor U9112 (N_9112,N_6173,N_6374);
or U9113 (N_9113,N_5261,N_4964);
or U9114 (N_9114,N_7864,N_7582);
and U9115 (N_9115,N_7971,N_5771);
and U9116 (N_9116,N_4347,N_5246);
and U9117 (N_9117,N_7437,N_5307);
or U9118 (N_9118,N_6268,N_6608);
and U9119 (N_9119,N_6540,N_7072);
nor U9120 (N_9120,N_7851,N_7675);
or U9121 (N_9121,N_5366,N_5136);
nand U9122 (N_9122,N_7988,N_6337);
or U9123 (N_9123,N_7042,N_7270);
nand U9124 (N_9124,N_6940,N_6573);
or U9125 (N_9125,N_4267,N_5758);
xor U9126 (N_9126,N_6517,N_6180);
nor U9127 (N_9127,N_5922,N_6408);
or U9128 (N_9128,N_5444,N_7524);
and U9129 (N_9129,N_4898,N_7156);
xor U9130 (N_9130,N_5011,N_4070);
nand U9131 (N_9131,N_7876,N_7302);
or U9132 (N_9132,N_5989,N_7275);
or U9133 (N_9133,N_6260,N_6339);
nand U9134 (N_9134,N_4520,N_5657);
or U9135 (N_9135,N_6199,N_5270);
nor U9136 (N_9136,N_5365,N_7750);
or U9137 (N_9137,N_5268,N_5274);
and U9138 (N_9138,N_5984,N_6024);
nor U9139 (N_9139,N_6612,N_5409);
nand U9140 (N_9140,N_7837,N_6748);
or U9141 (N_9141,N_7499,N_7238);
nor U9142 (N_9142,N_4310,N_7734);
or U9143 (N_9143,N_4738,N_6617);
nand U9144 (N_9144,N_5153,N_5453);
nand U9145 (N_9145,N_4478,N_5635);
nor U9146 (N_9146,N_4972,N_7525);
nand U9147 (N_9147,N_4648,N_6334);
nor U9148 (N_9148,N_4158,N_4444);
nor U9149 (N_9149,N_6341,N_5503);
and U9150 (N_9150,N_4531,N_6473);
and U9151 (N_9151,N_7792,N_4526);
and U9152 (N_9152,N_7719,N_5821);
nor U9153 (N_9153,N_5469,N_6759);
nand U9154 (N_9154,N_4605,N_7495);
nor U9155 (N_9155,N_5146,N_4903);
and U9156 (N_9156,N_7781,N_4344);
or U9157 (N_9157,N_5047,N_7616);
or U9158 (N_9158,N_4558,N_6580);
xnor U9159 (N_9159,N_7447,N_7212);
nor U9160 (N_9160,N_7637,N_6902);
xnor U9161 (N_9161,N_6154,N_6345);
nor U9162 (N_9162,N_7884,N_5320);
and U9163 (N_9163,N_6842,N_5923);
xnor U9164 (N_9164,N_5471,N_4838);
and U9165 (N_9165,N_6018,N_4427);
nand U9166 (N_9166,N_7800,N_6431);
nor U9167 (N_9167,N_6721,N_5161);
and U9168 (N_9168,N_4693,N_5195);
and U9169 (N_9169,N_7947,N_5804);
nand U9170 (N_9170,N_5201,N_6859);
or U9171 (N_9171,N_6417,N_4666);
or U9172 (N_9172,N_5702,N_4950);
nor U9173 (N_9173,N_6562,N_7518);
or U9174 (N_9174,N_7968,N_6525);
and U9175 (N_9175,N_5338,N_4816);
and U9176 (N_9176,N_7034,N_7321);
nor U9177 (N_9177,N_5128,N_6509);
and U9178 (N_9178,N_6203,N_6631);
and U9179 (N_9179,N_4356,N_7879);
nand U9180 (N_9180,N_4085,N_7011);
or U9181 (N_9181,N_6504,N_7911);
nor U9182 (N_9182,N_5298,N_7170);
nand U9183 (N_9183,N_6317,N_5611);
nor U9184 (N_9184,N_4848,N_6600);
nor U9185 (N_9185,N_5173,N_7621);
nand U9186 (N_9186,N_7061,N_5132);
nor U9187 (N_9187,N_7593,N_7142);
nor U9188 (N_9188,N_5207,N_4680);
nor U9189 (N_9189,N_6284,N_7820);
nand U9190 (N_9190,N_7109,N_5976);
nor U9191 (N_9191,N_7684,N_6192);
or U9192 (N_9192,N_7399,N_5986);
or U9193 (N_9193,N_4403,N_4298);
or U9194 (N_9194,N_4737,N_7651);
nand U9195 (N_9195,N_7808,N_4689);
or U9196 (N_9196,N_4234,N_4248);
xnor U9197 (N_9197,N_6651,N_5018);
and U9198 (N_9198,N_6894,N_5645);
xnor U9199 (N_9199,N_5544,N_5606);
and U9200 (N_9200,N_5181,N_5639);
nor U9201 (N_9201,N_5975,N_7799);
or U9202 (N_9202,N_6006,N_4845);
xnor U9203 (N_9203,N_5733,N_6624);
or U9204 (N_9204,N_7188,N_5176);
nor U9205 (N_9205,N_5172,N_4095);
or U9206 (N_9206,N_7473,N_6433);
nand U9207 (N_9207,N_6015,N_7358);
nand U9208 (N_9208,N_6936,N_5080);
or U9209 (N_9209,N_6876,N_4502);
or U9210 (N_9210,N_7628,N_5945);
or U9211 (N_9211,N_7571,N_6720);
or U9212 (N_9212,N_5779,N_5897);
nor U9213 (N_9213,N_4596,N_4337);
or U9214 (N_9214,N_6549,N_4216);
xnor U9215 (N_9215,N_6342,N_7624);
nor U9216 (N_9216,N_5566,N_7591);
and U9217 (N_9217,N_7644,N_6456);
and U9218 (N_9218,N_4618,N_7096);
or U9219 (N_9219,N_4084,N_4360);
and U9220 (N_9220,N_4566,N_5941);
nor U9221 (N_9221,N_7761,N_5813);
nor U9222 (N_9222,N_7057,N_6383);
nand U9223 (N_9223,N_4151,N_6004);
nor U9224 (N_9224,N_4464,N_7710);
nor U9225 (N_9225,N_5535,N_7414);
or U9226 (N_9226,N_5388,N_6719);
xor U9227 (N_9227,N_5105,N_6727);
nand U9228 (N_9228,N_7374,N_7397);
nor U9229 (N_9229,N_7629,N_6193);
nor U9230 (N_9230,N_6694,N_6281);
nand U9231 (N_9231,N_7094,N_4579);
nand U9232 (N_9232,N_7017,N_7802);
and U9233 (N_9233,N_4665,N_4786);
or U9234 (N_9234,N_4871,N_6063);
nor U9235 (N_9235,N_6114,N_5991);
nor U9236 (N_9236,N_7182,N_5255);
nor U9237 (N_9237,N_6584,N_6327);
nand U9238 (N_9238,N_6091,N_7960);
nand U9239 (N_9239,N_5488,N_5510);
nor U9240 (N_9240,N_4799,N_5248);
and U9241 (N_9241,N_7365,N_7663);
xnor U9242 (N_9242,N_4031,N_6122);
nand U9243 (N_9243,N_5571,N_4824);
nand U9244 (N_9244,N_5928,N_4256);
xnor U9245 (N_9245,N_5803,N_4717);
or U9246 (N_9246,N_6036,N_7067);
nor U9247 (N_9247,N_4224,N_7841);
nor U9248 (N_9248,N_6648,N_7683);
xor U9249 (N_9249,N_7230,N_5868);
or U9250 (N_9250,N_5370,N_4117);
nand U9251 (N_9251,N_6287,N_7857);
nand U9252 (N_9252,N_7043,N_7282);
and U9253 (N_9253,N_4876,N_4516);
or U9254 (N_9254,N_6380,N_5323);
nor U9255 (N_9255,N_7702,N_4636);
xnor U9256 (N_9256,N_5723,N_7211);
nor U9257 (N_9257,N_7250,N_4082);
and U9258 (N_9258,N_4025,N_6821);
nand U9259 (N_9259,N_5193,N_4273);
nor U9260 (N_9260,N_4710,N_4815);
nor U9261 (N_9261,N_6830,N_4706);
nand U9262 (N_9262,N_5260,N_5739);
nand U9263 (N_9263,N_7381,N_6915);
nor U9264 (N_9264,N_6519,N_7687);
nor U9265 (N_9265,N_5143,N_6402);
nand U9266 (N_9266,N_4716,N_7486);
or U9267 (N_9267,N_4971,N_5277);
and U9268 (N_9268,N_7075,N_4583);
or U9269 (N_9269,N_6766,N_7215);
nand U9270 (N_9270,N_4096,N_5688);
nand U9271 (N_9271,N_7504,N_4081);
nand U9272 (N_9272,N_6952,N_6315);
nand U9273 (N_9273,N_7822,N_6852);
nor U9274 (N_9274,N_6093,N_6770);
nor U9275 (N_9275,N_7613,N_5492);
nor U9276 (N_9276,N_7564,N_7050);
and U9277 (N_9277,N_4715,N_5185);
and U9278 (N_9278,N_4292,N_4866);
or U9279 (N_9279,N_7771,N_6427);
and U9280 (N_9280,N_4040,N_6156);
or U9281 (N_9281,N_6948,N_7527);
nor U9282 (N_9282,N_4198,N_5903);
and U9283 (N_9283,N_7476,N_7085);
or U9284 (N_9284,N_5328,N_5837);
or U9285 (N_9285,N_6458,N_4157);
or U9286 (N_9286,N_4804,N_6019);
and U9287 (N_9287,N_6665,N_4280);
or U9288 (N_9288,N_6185,N_7202);
and U9289 (N_9289,N_6039,N_5782);
nand U9290 (N_9290,N_7239,N_7187);
nor U9291 (N_9291,N_7224,N_5096);
or U9292 (N_9292,N_7805,N_4916);
and U9293 (N_9293,N_5393,N_4522);
nor U9294 (N_9294,N_5461,N_5776);
nor U9295 (N_9295,N_7692,N_4284);
nand U9296 (N_9296,N_5164,N_6655);
xor U9297 (N_9297,N_7532,N_4028);
nor U9298 (N_9298,N_6647,N_6843);
or U9299 (N_9299,N_4959,N_7484);
and U9300 (N_9300,N_4077,N_7965);
nand U9301 (N_9301,N_7744,N_4759);
nor U9302 (N_9302,N_7941,N_6434);
xnor U9303 (N_9303,N_5069,N_5685);
nor U9304 (N_9304,N_7757,N_7898);
or U9305 (N_9305,N_7631,N_5509);
or U9306 (N_9306,N_7214,N_6338);
and U9307 (N_9307,N_5619,N_6550);
nand U9308 (N_9308,N_6760,N_4357);
or U9309 (N_9309,N_4621,N_4002);
nor U9310 (N_9310,N_6296,N_7553);
and U9311 (N_9311,N_5917,N_6162);
nand U9312 (N_9312,N_4800,N_4276);
and U9313 (N_9313,N_4571,N_5850);
nand U9314 (N_9314,N_5294,N_6119);
or U9315 (N_9315,N_6925,N_5819);
nor U9316 (N_9316,N_4517,N_6938);
or U9317 (N_9317,N_7363,N_4311);
and U9318 (N_9318,N_7107,N_6409);
or U9319 (N_9319,N_7574,N_4606);
nor U9320 (N_9320,N_5152,N_4250);
xor U9321 (N_9321,N_5015,N_4535);
and U9322 (N_9322,N_4482,N_4230);
nand U9323 (N_9323,N_4038,N_6072);
nor U9324 (N_9324,N_5032,N_5092);
xnor U9325 (N_9325,N_7234,N_7895);
xnor U9326 (N_9326,N_7451,N_7538);
or U9327 (N_9327,N_6980,N_6105);
and U9328 (N_9328,N_7872,N_7848);
or U9329 (N_9329,N_4952,N_4731);
or U9330 (N_9330,N_6057,N_6644);
nand U9331 (N_9331,N_4262,N_6414);
nor U9332 (N_9332,N_5575,N_4457);
and U9333 (N_9333,N_7995,N_7283);
nor U9334 (N_9334,N_7903,N_6769);
or U9335 (N_9335,N_6718,N_7720);
and U9336 (N_9336,N_4819,N_7520);
or U9337 (N_9337,N_6897,N_4709);
nand U9338 (N_9338,N_7685,N_4308);
nand U9339 (N_9339,N_7843,N_5147);
nor U9340 (N_9340,N_6697,N_7172);
nor U9341 (N_9341,N_4235,N_7723);
or U9342 (N_9342,N_7824,N_4884);
xnor U9343 (N_9343,N_6862,N_5275);
or U9344 (N_9344,N_5579,N_6961);
and U9345 (N_9345,N_4466,N_7485);
or U9346 (N_9346,N_4597,N_4306);
nand U9347 (N_9347,N_4888,N_6641);
xor U9348 (N_9348,N_7794,N_6569);
nor U9349 (N_9349,N_4868,N_4328);
nand U9350 (N_9350,N_5778,N_6480);
or U9351 (N_9351,N_4370,N_7736);
nand U9352 (N_9352,N_4967,N_5536);
nor U9353 (N_9353,N_4632,N_5847);
nand U9354 (N_9354,N_7919,N_4795);
nand U9355 (N_9355,N_5067,N_7783);
nor U9356 (N_9356,N_5183,N_5476);
or U9357 (N_9357,N_5968,N_4182);
and U9358 (N_9358,N_4486,N_5557);
or U9359 (N_9359,N_5907,N_4631);
or U9360 (N_9360,N_5729,N_6286);
nor U9361 (N_9361,N_4953,N_6172);
nor U9362 (N_9362,N_5205,N_6252);
nand U9363 (N_9363,N_7691,N_4385);
nor U9364 (N_9364,N_6963,N_4253);
nand U9365 (N_9365,N_6060,N_5169);
nand U9366 (N_9366,N_4277,N_5741);
xor U9367 (N_9367,N_5447,N_7412);
nand U9368 (N_9368,N_4664,N_5682);
or U9369 (N_9369,N_7620,N_6196);
and U9370 (N_9370,N_6086,N_6858);
nor U9371 (N_9371,N_4555,N_7576);
and U9372 (N_9372,N_7168,N_5790);
or U9373 (N_9373,N_7634,N_7409);
or U9374 (N_9374,N_7355,N_4144);
xor U9375 (N_9375,N_6333,N_5594);
or U9376 (N_9376,N_6486,N_7809);
nand U9377 (N_9377,N_4315,N_6632);
xor U9378 (N_9378,N_6464,N_7343);
nand U9379 (N_9379,N_4377,N_7247);
or U9380 (N_9380,N_5043,N_4770);
nor U9381 (N_9381,N_4537,N_7059);
nand U9382 (N_9382,N_6875,N_5287);
and U9383 (N_9383,N_6561,N_6652);
and U9384 (N_9384,N_7672,N_7679);
nand U9385 (N_9385,N_4740,N_7933);
and U9386 (N_9386,N_7081,N_7375);
nor U9387 (N_9387,N_7436,N_5214);
nor U9388 (N_9388,N_7488,N_6332);
or U9389 (N_9389,N_7213,N_5187);
and U9390 (N_9390,N_5900,N_5306);
and U9391 (N_9391,N_5363,N_5312);
nand U9392 (N_9392,N_5919,N_6551);
xnor U9393 (N_9393,N_5209,N_5336);
xnor U9394 (N_9394,N_6210,N_7052);
nor U9395 (N_9395,N_6163,N_7866);
nor U9396 (N_9396,N_7830,N_4189);
nor U9397 (N_9397,N_5380,N_4137);
xor U9398 (N_9398,N_4092,N_4122);
nand U9399 (N_9399,N_7261,N_4877);
or U9400 (N_9400,N_6685,N_5433);
nand U9401 (N_9401,N_7948,N_5017);
or U9402 (N_9402,N_7403,N_5879);
and U9403 (N_9403,N_7465,N_7906);
nand U9404 (N_9404,N_4346,N_7413);
xnor U9405 (N_9405,N_4231,N_7708);
nand U9406 (N_9406,N_6375,N_4854);
xor U9407 (N_9407,N_6905,N_7019);
nor U9408 (N_9408,N_4047,N_4727);
nor U9409 (N_9409,N_5354,N_6314);
xor U9410 (N_9410,N_4005,N_7225);
xnor U9411 (N_9411,N_5269,N_4359);
nand U9412 (N_9412,N_5401,N_7171);
xnor U9413 (N_9413,N_6243,N_4023);
or U9414 (N_9414,N_6313,N_4167);
and U9415 (N_9415,N_7255,N_6958);
or U9416 (N_9416,N_5427,N_6995);
and U9417 (N_9417,N_4161,N_4942);
xnor U9418 (N_9418,N_6663,N_4541);
nand U9419 (N_9419,N_5817,N_7022);
xnor U9420 (N_9420,N_7468,N_5372);
nand U9421 (N_9421,N_4463,N_7100);
and U9422 (N_9422,N_7227,N_6420);
nor U9423 (N_9423,N_4784,N_7331);
and U9424 (N_9424,N_5377,N_5590);
nand U9425 (N_9425,N_5610,N_6997);
nor U9426 (N_9426,N_4696,N_5182);
or U9427 (N_9427,N_5860,N_5537);
and U9428 (N_9428,N_5558,N_5507);
nor U9429 (N_9429,N_4313,N_4422);
nor U9430 (N_9430,N_6128,N_4694);
or U9431 (N_9431,N_5568,N_5266);
xor U9432 (N_9432,N_7254,N_5166);
nor U9433 (N_9433,N_7914,N_4175);
xnor U9434 (N_9434,N_6604,N_6487);
nand U9435 (N_9435,N_7304,N_4162);
and U9436 (N_9436,N_5800,N_7105);
nand U9437 (N_9437,N_7038,N_6127);
and U9438 (N_9438,N_5332,N_5811);
nand U9439 (N_9439,N_4364,N_6445);
or U9440 (N_9440,N_4060,N_6033);
nand U9441 (N_9441,N_4405,N_5073);
nand U9442 (N_9442,N_4112,N_4945);
or U9443 (N_9443,N_7880,N_6289);
and U9444 (N_9444,N_5351,N_4834);
and U9445 (N_9445,N_5743,N_7082);
nor U9446 (N_9446,N_5731,N_6184);
xnor U9447 (N_9447,N_4076,N_7297);
and U9448 (N_9448,N_5769,N_5217);
xnor U9449 (N_9449,N_7625,N_6677);
or U9450 (N_9450,N_6907,N_7745);
or U9451 (N_9451,N_7510,N_7658);
or U9452 (N_9452,N_6693,N_7133);
and U9453 (N_9453,N_7131,N_4229);
or U9454 (N_9454,N_7665,N_5926);
or U9455 (N_9455,N_6285,N_6636);
xnor U9456 (N_9456,N_6535,N_6564);
nor U9457 (N_9457,N_4572,N_7015);
or U9458 (N_9458,N_6428,N_5243);
or U9459 (N_9459,N_4989,N_4504);
nand U9460 (N_9460,N_4333,N_6796);
nor U9461 (N_9461,N_5889,N_6810);
nand U9462 (N_9462,N_4564,N_4925);
xnor U9463 (N_9463,N_7339,N_6797);
nor U9464 (N_9464,N_5979,N_7768);
nor U9465 (N_9465,N_6466,N_6623);
nor U9466 (N_9466,N_5434,N_4999);
or U9467 (N_9467,N_6650,N_7904);
and U9468 (N_9468,N_5692,N_5745);
or U9469 (N_9469,N_7013,N_7555);
nand U9470 (N_9470,N_5871,N_4233);
or U9471 (N_9471,N_7191,N_4763);
xor U9472 (N_9472,N_5392,N_6293);
nor U9473 (N_9473,N_6939,N_7507);
and U9474 (N_9474,N_5937,N_6740);
and U9475 (N_9475,N_7129,N_5111);
and U9476 (N_9476,N_7917,N_6989);
nand U9477 (N_9477,N_4239,N_6142);
nand U9478 (N_9478,N_6328,N_6167);
or U9479 (N_9479,N_6994,N_4468);
nand U9480 (N_9480,N_4677,N_7581);
xor U9481 (N_9481,N_5007,N_7301);
nor U9482 (N_9482,N_4752,N_7548);
nor U9483 (N_9483,N_6851,N_5478);
nor U9484 (N_9484,N_4728,N_7278);
nor U9485 (N_9485,N_4120,N_5324);
nand U9486 (N_9486,N_4279,N_7330);
or U9487 (N_9487,N_5443,N_6000);
nor U9488 (N_9488,N_4289,N_4619);
or U9489 (N_9489,N_4013,N_6860);
and U9490 (N_9490,N_6783,N_4974);
or U9491 (N_9491,N_4521,N_5599);
nand U9492 (N_9492,N_6870,N_6145);
and U9493 (N_9493,N_6931,N_6366);
and U9494 (N_9494,N_5000,N_7432);
xor U9495 (N_9495,N_6251,N_5072);
nor U9496 (N_9496,N_6911,N_5699);
xor U9497 (N_9497,N_5122,N_6005);
and U9498 (N_9498,N_7923,N_6553);
xor U9499 (N_9499,N_7177,N_4736);
or U9500 (N_9500,N_6044,N_4430);
nor U9501 (N_9501,N_6606,N_6520);
nor U9502 (N_9502,N_5565,N_4324);
xnor U9503 (N_9503,N_5319,N_5234);
xor U9504 (N_9504,N_4105,N_5362);
nand U9505 (N_9505,N_6725,N_6062);
or U9506 (N_9506,N_5513,N_6231);
xnor U9507 (N_9507,N_6228,N_6908);
xnor U9508 (N_9508,N_5512,N_7315);
nor U9509 (N_9509,N_6453,N_6820);
nand U9510 (N_9510,N_6391,N_4545);
and U9511 (N_9511,N_4154,N_5585);
nor U9512 (N_9512,N_5874,N_6229);
nand U9513 (N_9513,N_7400,N_6732);
and U9514 (N_9514,N_6100,N_6935);
or U9515 (N_9515,N_5592,N_4476);
and U9516 (N_9516,N_4271,N_5569);
nand U9517 (N_9517,N_5953,N_4756);
or U9518 (N_9518,N_6951,N_7845);
nand U9519 (N_9519,N_5474,N_5842);
nand U9520 (N_9520,N_6695,N_4431);
nor U9521 (N_9521,N_6085,N_5957);
nor U9522 (N_9522,N_5992,N_5612);
nand U9523 (N_9523,N_7008,N_6115);
nor U9524 (N_9524,N_4574,N_6246);
or U9525 (N_9525,N_4627,N_7951);
nand U9526 (N_9526,N_5144,N_7552);
xnor U9527 (N_9527,N_5455,N_5416);
nor U9528 (N_9528,N_6151,N_5022);
and U9529 (N_9529,N_5736,N_4661);
or U9530 (N_9530,N_4634,N_7431);
or U9531 (N_9531,N_7223,N_4948);
or U9532 (N_9532,N_7078,N_7877);
nand U9533 (N_9533,N_4588,N_5028);
nor U9534 (N_9534,N_7185,N_7630);
or U9535 (N_9535,N_4307,N_4822);
nand U9536 (N_9536,N_7874,N_7840);
xor U9537 (N_9537,N_4448,N_7626);
or U9538 (N_9538,N_5222,N_5876);
and U9539 (N_9539,N_6188,N_6686);
or U9540 (N_9540,N_4302,N_7893);
xnor U9541 (N_9541,N_5436,N_7418);
nor U9542 (N_9542,N_6816,N_5753);
nand U9543 (N_9543,N_7765,N_7446);
and U9544 (N_9544,N_6325,N_4498);
nand U9545 (N_9545,N_7615,N_6984);
and U9546 (N_9546,N_7899,N_7472);
nor U9547 (N_9547,N_4663,N_5118);
nand U9548 (N_9548,N_7421,N_7175);
and U9549 (N_9549,N_4609,N_4864);
nand U9550 (N_9550,N_7118,N_7764);
nor U9551 (N_9551,N_5335,N_7797);
xor U9552 (N_9552,N_6501,N_6112);
xnor U9553 (N_9553,N_7056,N_5084);
or U9554 (N_9554,N_4399,N_7738);
and U9555 (N_9555,N_7922,N_5604);
nand U9556 (N_9556,N_4147,N_5662);
nor U9557 (N_9557,N_6671,N_4051);
nor U9558 (N_9558,N_4459,N_7079);
and U9559 (N_9559,N_7166,N_7836);
nand U9560 (N_9560,N_6726,N_4048);
and U9561 (N_9561,N_4453,N_4493);
and U9562 (N_9562,N_7709,N_4836);
nand U9563 (N_9563,N_6439,N_5148);
and U9564 (N_9564,N_7457,N_6891);
xor U9565 (N_9565,N_6303,N_7351);
and U9566 (N_9566,N_5290,N_5840);
and U9567 (N_9567,N_4810,N_7755);
or U9568 (N_9568,N_4210,N_6113);
nand U9569 (N_9569,N_4567,N_7763);
nor U9570 (N_9570,N_7087,N_7562);
nand U9571 (N_9571,N_5600,N_6679);
xnor U9572 (N_9572,N_6200,N_4080);
xnor U9573 (N_9573,N_4391,N_5559);
nor U9574 (N_9574,N_7991,N_7670);
and U9575 (N_9575,N_7908,N_6964);
or U9576 (N_9576,N_6195,N_4269);
or U9577 (N_9577,N_5419,N_5730);
and U9578 (N_9578,N_6855,N_4947);
nor U9579 (N_9579,N_6102,N_5371);
nand U9580 (N_9580,N_6307,N_6379);
nand U9581 (N_9581,N_7453,N_4960);
nand U9582 (N_9582,N_6536,N_7707);
or U9583 (N_9583,N_7009,N_7303);
and U9584 (N_9584,N_7357,N_7522);
nand U9585 (N_9585,N_5521,N_7533);
nand U9586 (N_9586,N_4553,N_5463);
xnor U9587 (N_9587,N_6136,N_4325);
nand U9588 (N_9588,N_5740,N_4533);
and U9589 (N_9589,N_6109,N_6346);
and U9590 (N_9590,N_6926,N_6699);
nor U9591 (N_9591,N_6558,N_6282);
nand U9592 (N_9592,N_6489,N_6711);
and U9593 (N_9593,N_6144,N_5553);
or U9594 (N_9594,N_5648,N_6722);
nand U9595 (N_9595,N_6108,N_4645);
nand U9596 (N_9596,N_4286,N_4839);
nand U9597 (N_9597,N_4176,N_5881);
or U9598 (N_9598,N_5573,N_4626);
xnor U9599 (N_9599,N_4760,N_7949);
or U9600 (N_9600,N_4849,N_4951);
nand U9601 (N_9601,N_7356,N_4413);
nand U9602 (N_9602,N_5394,N_5942);
nor U9603 (N_9603,N_7661,N_4753);
or U9604 (N_9604,N_6276,N_7526);
and U9605 (N_9605,N_5218,N_5638);
or U9606 (N_9606,N_4983,N_6059);
or U9607 (N_9607,N_6275,N_5719);
nand U9608 (N_9608,N_6377,N_4559);
or U9609 (N_9609,N_7284,N_7058);
nor U9610 (N_9610,N_4996,N_6369);
nor U9611 (N_9611,N_6739,N_7165);
nand U9612 (N_9612,N_6691,N_7986);
or U9613 (N_9613,N_7936,N_4872);
and U9614 (N_9614,N_4506,N_4299);
and U9615 (N_9615,N_5828,N_7328);
or U9616 (N_9616,N_4242,N_4414);
or U9617 (N_9617,N_4690,N_5904);
nor U9618 (N_9618,N_6874,N_6753);
or U9619 (N_9619,N_7567,N_5806);
nand U9620 (N_9620,N_6621,N_4580);
nor U9621 (N_9621,N_6528,N_4071);
nand U9622 (N_9622,N_6499,N_4842);
nor U9623 (N_9623,N_6658,N_7979);
and U9624 (N_9624,N_7535,N_4309);
or U9625 (N_9625,N_5479,N_6785);
nand U9626 (N_9626,N_4993,N_5117);
nand U9627 (N_9627,N_5935,N_6316);
and U9628 (N_9628,N_7271,N_5179);
and U9629 (N_9629,N_7718,N_5197);
and U9630 (N_9630,N_7943,N_4907);
or U9631 (N_9631,N_5318,N_4534);
nor U9632 (N_9632,N_4223,N_6146);
and U9633 (N_9633,N_5936,N_5491);
xnor U9634 (N_9634,N_7878,N_4790);
nand U9635 (N_9635,N_4542,N_4995);
nand U9636 (N_9636,N_5760,N_4113);
nand U9637 (N_9637,N_5671,N_4902);
or U9638 (N_9638,N_5947,N_7546);
or U9639 (N_9639,N_4814,N_5381);
or U9640 (N_9640,N_5652,N_5041);
nand U9641 (N_9641,N_5333,N_5107);
nor U9642 (N_9642,N_7776,N_4055);
and U9643 (N_9643,N_6111,N_6778);
or U9644 (N_9644,N_6850,N_4361);
nand U9645 (N_9645,N_7120,N_5703);
or U9646 (N_9646,N_6356,N_7121);
or U9647 (N_9647,N_6588,N_6270);
nor U9648 (N_9648,N_5481,N_7814);
nand U9649 (N_9649,N_5301,N_5576);
and U9650 (N_9650,N_6839,N_7985);
and U9651 (N_9651,N_6625,N_4979);
nor U9652 (N_9652,N_7785,N_4887);
nand U9653 (N_9653,N_5340,N_4893);
nand U9654 (N_9654,N_7464,N_5184);
or U9655 (N_9655,N_7855,N_7870);
and U9656 (N_9656,N_4852,N_4525);
or U9657 (N_9657,N_6804,N_5192);
or U9658 (N_9658,N_5993,N_5667);
nand U9659 (N_9659,N_6921,N_7192);
or U9660 (N_9660,N_7927,N_6097);
nand U9661 (N_9661,N_4772,N_5407);
nand U9662 (N_9662,N_5855,N_6966);
xnor U9663 (N_9663,N_4367,N_5873);
and U9664 (N_9664,N_5515,N_4507);
nor U9665 (N_9665,N_6037,N_6567);
nand U9666 (N_9666,N_6058,N_7228);
and U9667 (N_9667,N_7698,N_7989);
and U9668 (N_9668,N_5773,N_4724);
xnor U9669 (N_9669,N_4458,N_4813);
nor U9670 (N_9670,N_6424,N_7427);
nor U9671 (N_9671,N_6557,N_6425);
and U9672 (N_9672,N_7306,N_5921);
nor U9673 (N_9673,N_4183,N_7281);
nand U9674 (N_9674,N_4615,N_5231);
and U9675 (N_9675,N_7536,N_5089);
nor U9676 (N_9676,N_6910,N_6795);
nand U9677 (N_9677,N_4885,N_5916);
or U9678 (N_9678,N_6996,N_5103);
and U9679 (N_9679,N_6976,N_5334);
nand U9680 (N_9680,N_5689,N_6220);
and U9681 (N_9681,N_6983,N_7242);
nand U9682 (N_9682,N_7549,N_6215);
or U9683 (N_9683,N_7640,N_5770);
nand U9684 (N_9684,N_6878,N_4859);
nand U9685 (N_9685,N_4093,N_5858);
xor U9686 (N_9686,N_7151,N_4134);
nor U9687 (N_9687,N_5596,N_4593);
and U9688 (N_9688,N_7657,N_4920);
xnor U9689 (N_9689,N_5902,N_4544);
or U9690 (N_9690,N_4352,N_4941);
xor U9691 (N_9691,N_5240,N_6398);
xnor U9692 (N_9692,N_7482,N_7573);
nand U9693 (N_9693,N_6867,N_5511);
or U9694 (N_9694,N_6818,N_6454);
and U9695 (N_9695,N_7428,N_6806);
or U9696 (N_9696,N_5925,N_4185);
nor U9697 (N_9697,N_6526,N_7396);
or U9698 (N_9698,N_7727,N_6001);
and U9699 (N_9699,N_5934,N_4450);
and U9700 (N_9700,N_6038,N_5988);
xor U9701 (N_9701,N_5150,N_6831);
or U9702 (N_9702,N_6035,N_5272);
nor U9703 (N_9703,N_4692,N_7506);
nand U9704 (N_9704,N_6257,N_6888);
nor U9705 (N_9705,N_5082,N_4570);
nand U9706 (N_9706,N_6515,N_4720);
or U9707 (N_9707,N_6613,N_6792);
and U9708 (N_9708,N_7497,N_4765);
nor U9709 (N_9709,N_5901,N_7448);
nand U9710 (N_9710,N_7896,N_7612);
nor U9711 (N_9711,N_5698,N_6761);
xor U9712 (N_9712,N_4179,N_5848);
and U9713 (N_9713,N_6594,N_4196);
nand U9714 (N_9714,N_7955,N_4581);
or U9715 (N_9715,N_6757,N_6605);
or U9716 (N_9716,N_7728,N_5279);
xor U9717 (N_9717,N_5949,N_5807);
nor U9718 (N_9718,N_5701,N_4257);
nor U9719 (N_9719,N_5387,N_5230);
nand U9720 (N_9720,N_5468,N_4044);
nand U9721 (N_9721,N_5732,N_7614);
nor U9722 (N_9722,N_4676,N_4083);
nand U9723 (N_9723,N_5288,N_6903);
nor U9724 (N_9724,N_5972,N_6924);
and U9725 (N_9725,N_5200,N_5785);
nor U9726 (N_9726,N_6362,N_7901);
xnor U9727 (N_9727,N_5303,N_4045);
or U9728 (N_9728,N_7123,N_6164);
nor U9729 (N_9729,N_6779,N_4977);
nor U9730 (N_9730,N_4565,N_6071);
nor U9731 (N_9731,N_7350,N_5259);
or U9732 (N_9732,N_6025,N_7296);
nand U9733 (N_9733,N_7389,N_6302);
nand U9734 (N_9734,N_6376,N_7509);
nor U9735 (N_9735,N_5593,N_7205);
or U9736 (N_9736,N_6191,N_4475);
nand U9737 (N_9737,N_7021,N_7821);
nand U9738 (N_9738,N_6159,N_6412);
and U9739 (N_9739,N_7715,N_6530);
nor U9740 (N_9740,N_5346,N_6576);
or U9741 (N_9741,N_6836,N_4046);
nand U9742 (N_9742,N_7493,N_4723);
or U9743 (N_9743,N_5345,N_7980);
nand U9744 (N_9744,N_5915,N_6684);
and U9745 (N_9745,N_7006,N_7066);
nor U9746 (N_9746,N_7769,N_6134);
xnor U9747 (N_9747,N_7456,N_6570);
or U9748 (N_9748,N_6708,N_4007);
and U9749 (N_9749,N_6649,N_4538);
and U9750 (N_9750,N_7743,N_5614);
nor U9751 (N_9751,N_4481,N_6868);
and U9752 (N_9752,N_5636,N_4168);
nor U9753 (N_9753,N_4456,N_6871);
xor U9754 (N_9754,N_6682,N_5791);
or U9755 (N_9755,N_7354,N_4867);
and U9756 (N_9756,N_6987,N_6965);
and U9757 (N_9757,N_7169,N_5809);
or U9758 (N_9758,N_7219,N_6762);
and U9759 (N_9759,N_7846,N_5716);
nor U9760 (N_9760,N_5990,N_4791);
nand U9761 (N_9761,N_5628,N_7295);
nand U9762 (N_9762,N_7329,N_6386);
nor U9763 (N_9763,N_5533,N_6812);
nor U9764 (N_9764,N_6234,N_7962);
nand U9765 (N_9765,N_4801,N_7455);
and U9766 (N_9766,N_6723,N_5095);
or U9767 (N_9767,N_5932,N_7572);
nor U9768 (N_9768,N_5582,N_6742);
nand U9769 (N_9769,N_6084,N_5221);
and U9770 (N_9770,N_7231,N_6668);
nor U9771 (N_9771,N_4853,N_7772);
or U9772 (N_9772,N_6360,N_7787);
or U9773 (N_9773,N_7964,N_6103);
or U9774 (N_9774,N_5799,N_4762);
and U9775 (N_9775,N_4861,N_4789);
and U9776 (N_9776,N_6347,N_5825);
nand U9777 (N_9777,N_7010,N_4485);
nand U9778 (N_9778,N_5308,N_6244);
nor U9779 (N_9779,N_5895,N_5142);
and U9780 (N_9780,N_7439,N_5276);
nand U9781 (N_9781,N_6027,N_5857);
xor U9782 (N_9782,N_5415,N_6367);
and U9783 (N_9783,N_4713,N_5325);
nand U9784 (N_9784,N_6781,N_5055);
and U9785 (N_9785,N_5797,N_7742);
and U9786 (N_9786,N_6017,N_6841);
nand U9787 (N_9787,N_5883,N_5083);
nor U9788 (N_9788,N_4135,N_6358);
and U9789 (N_9789,N_5795,N_6746);
and U9790 (N_9790,N_5763,N_5191);
xnor U9791 (N_9791,N_4146,N_6768);
nor U9792 (N_9792,N_5659,N_4501);
or U9793 (N_9793,N_6802,N_4500);
and U9794 (N_9794,N_4170,N_6090);
or U9795 (N_9795,N_5404,N_4739);
nor U9796 (N_9796,N_5864,N_4809);
nor U9797 (N_9797,N_7681,N_7655);
and U9798 (N_9798,N_7760,N_7377);
and U9799 (N_9799,N_5869,N_6291);
and U9800 (N_9800,N_6670,N_7907);
nor U9801 (N_9801,N_6899,N_4194);
nand U9802 (N_9802,N_7395,N_4473);
and U9803 (N_9803,N_6153,N_5754);
nor U9804 (N_9804,N_7500,N_4001);
or U9805 (N_9805,N_5313,N_6032);
or U9806 (N_9806,N_5016,N_7773);
nand U9807 (N_9807,N_7407,N_4857);
nand U9808 (N_9808,N_7733,N_4329);
and U9809 (N_9809,N_7394,N_5856);
and U9810 (N_9810,N_6710,N_5728);
and U9811 (N_9811,N_4755,N_4265);
xnor U9812 (N_9812,N_5114,N_7854);
nand U9813 (N_9813,N_6676,N_4595);
nor U9814 (N_9814,N_6283,N_6981);
and U9815 (N_9815,N_5138,N_5905);
nand U9816 (N_9816,N_6942,N_4965);
and U9817 (N_9817,N_4006,N_4523);
xor U9818 (N_9818,N_4181,N_7490);
and U9819 (N_9819,N_4530,N_4052);
nor U9820 (N_9820,N_6654,N_4097);
or U9821 (N_9821,N_7578,N_7601);
xor U9822 (N_9822,N_4184,N_7236);
xor U9823 (N_9823,N_7292,N_4963);
nand U9824 (N_9824,N_7654,N_6945);
or U9825 (N_9825,N_5237,N_5213);
xor U9826 (N_9826,N_7092,N_6503);
nor U9827 (N_9827,N_6248,N_4745);
nand U9828 (N_9828,N_7030,N_5861);
or U9829 (N_9829,N_7433,N_6791);
nand U9830 (N_9830,N_7666,N_7210);
or U9831 (N_9831,N_7981,N_5450);
nand U9832 (N_9832,N_4601,N_6805);
xor U9833 (N_9833,N_7648,N_5109);
nand U9834 (N_9834,N_4074,N_7274);
nor U9835 (N_9835,N_4639,N_6106);
nand U9836 (N_9836,N_4348,N_6031);
nand U9837 (N_9837,N_5534,N_6395);
or U9838 (N_9838,N_6223,N_4004);
nand U9839 (N_9839,N_6840,N_7245);
and U9840 (N_9840,N_4358,N_5738);
and U9841 (N_9841,N_6461,N_5374);
and U9842 (N_9842,N_5360,N_5019);
or U9843 (N_9843,N_6614,N_6008);
and U9844 (N_9844,N_4625,N_6883);
and U9845 (N_9845,N_4064,N_7150);
nor U9846 (N_9846,N_7217,N_4806);
xor U9847 (N_9847,N_4794,N_5961);
or U9848 (N_9848,N_5823,N_4237);
nand U9849 (N_9849,N_5587,N_4782);
nand U9850 (N_9850,N_6104,N_4379);
or U9851 (N_9851,N_7587,N_7721);
or U9852 (N_9852,N_5235,N_5849);
or U9853 (N_9853,N_7699,N_6656);
nand U9854 (N_9854,N_4140,N_7853);
or U9855 (N_9855,N_7053,N_5818);
nor U9856 (N_9856,N_7953,N_5591);
nor U9857 (N_9857,N_5747,N_6853);
or U9858 (N_9858,N_5226,N_6459);
xor U9859 (N_9859,N_4355,N_7290);
and U9860 (N_9860,N_5880,N_7784);
and U9861 (N_9861,N_6189,N_6962);
nand U9862 (N_9862,N_5160,N_6775);
and U9863 (N_9863,N_5882,N_5058);
nand U9864 (N_9864,N_6637,N_4244);
and U9865 (N_9865,N_5149,N_4891);
or U9866 (N_9866,N_5792,N_6803);
or U9867 (N_9867,N_7741,N_7952);
nand U9868 (N_9868,N_7569,N_4831);
nor U9869 (N_9869,N_6544,N_6634);
nor U9870 (N_9870,N_6492,N_4779);
and U9871 (N_9871,N_6599,N_7706);
nand U9872 (N_9872,N_7993,N_6124);
nand U9873 (N_9873,N_6457,N_5617);
nor U9874 (N_9874,N_5361,N_4985);
and U9875 (N_9875,N_6166,N_7221);
nor U9876 (N_9876,N_5930,N_4067);
nor U9877 (N_9877,N_5663,N_4587);
xnor U9878 (N_9878,N_7098,N_4221);
or U9879 (N_9879,N_5005,N_5584);
and U9880 (N_9880,N_4026,N_7481);
nand U9881 (N_9881,N_5634,N_4027);
nand U9882 (N_9882,N_7208,N_4214);
nor U9883 (N_9883,N_4039,N_7690);
nor U9884 (N_9884,N_6847,N_7449);
nand U9885 (N_9885,N_7475,N_7164);
and U9886 (N_9886,N_6340,N_6174);
nor U9887 (N_9887,N_6546,N_4446);
nor U9888 (N_9888,N_6755,N_4878);
nor U9889 (N_9889,N_7189,N_6618);
or U9890 (N_9890,N_7619,N_4291);
nand U9891 (N_9891,N_7140,N_4104);
nand U9892 (N_9892,N_6512,N_6202);
xnor U9893 (N_9893,N_6960,N_5487);
nor U9894 (N_9894,N_5995,N_5154);
xnor U9895 (N_9895,N_5440,N_5344);
and U9896 (N_9896,N_6978,N_4397);
and U9897 (N_9897,N_6421,N_5413);
xor U9898 (N_9898,N_7996,N_4008);
nor U9899 (N_9899,N_5618,N_4630);
or U9900 (N_9900,N_5838,N_4100);
and U9901 (N_9901,N_5186,N_5885);
nor U9902 (N_9902,N_7643,N_4021);
nand U9903 (N_9903,N_7530,N_5950);
nand U9904 (N_9904,N_6881,N_4624);
nor U9905 (N_9905,N_5042,N_4268);
xnor U9906 (N_9906,N_7813,N_7444);
or U9907 (N_9907,N_5661,N_6278);
nor U9908 (N_9908,N_5615,N_4536);
and U9909 (N_9909,N_4923,N_7319);
or U9910 (N_9910,N_5386,N_7385);
xnor U9911 (N_9911,N_6481,N_6955);
or U9912 (N_9912,N_4102,N_7924);
and U9913 (N_9913,N_6906,N_6138);
or U9914 (N_9914,N_7474,N_4425);
and U9915 (N_9915,N_6974,N_5608);
xor U9916 (N_9916,N_6717,N_5609);
nand U9917 (N_9917,N_4381,N_4033);
nor U9918 (N_9918,N_6170,N_4585);
nor U9919 (N_9919,N_4969,N_6465);
xnor U9920 (N_9920,N_6165,N_7026);
nor U9921 (N_9921,N_7068,N_5554);
nor U9922 (N_9922,N_4556,N_6696);
nor U9923 (N_9923,N_6583,N_7025);
and U9924 (N_9924,N_5960,N_6430);
or U9925 (N_9925,N_4735,N_6121);
and U9926 (N_9926,N_5076,N_5954);
and U9927 (N_9927,N_7420,N_4929);
and U9928 (N_9928,N_6620,N_5203);
nor U9929 (N_9929,N_7642,N_4900);
or U9930 (N_9930,N_6264,N_5714);
or U9931 (N_9931,N_5044,N_5174);
or U9932 (N_9932,N_4441,N_7984);
nor U9933 (N_9933,N_4011,N_4118);
nand U9934 (N_9934,N_7124,N_5459);
or U9935 (N_9935,N_5865,N_5870);
nor U9936 (N_9936,N_5438,N_6131);
or U9937 (N_9937,N_4163,N_4874);
or U9938 (N_9938,N_7135,N_5020);
xor U9939 (N_9939,N_5726,N_5939);
nor U9940 (N_9940,N_5551,N_7858);
nand U9941 (N_9941,N_4090,N_6554);
or U9942 (N_9942,N_4386,N_4820);
and U9943 (N_9943,N_4582,N_4833);
or U9944 (N_9944,N_7671,N_7725);
or U9945 (N_9945,N_7915,N_4599);
and U9946 (N_9946,N_4086,N_7370);
and U9947 (N_9947,N_6610,N_6971);
nand U9948 (N_9948,N_5250,N_4022);
or U9949 (N_9949,N_6415,N_4751);
or U9950 (N_9950,N_7748,N_5086);
xor U9951 (N_9951,N_6323,N_5751);
nor U9952 (N_9952,N_7155,N_5705);
or U9953 (N_9953,N_5630,N_4389);
and U9954 (N_9954,N_6147,N_5794);
xor U9955 (N_9955,N_7148,N_5495);
or U9956 (N_9956,N_4119,N_4847);
or U9957 (N_9957,N_7531,N_4835);
or U9958 (N_9958,N_6045,N_4354);
nand U9959 (N_9959,N_7974,N_6258);
or U9960 (N_9960,N_4793,N_6591);
nor U9961 (N_9961,N_5978,N_5137);
nor U9962 (N_9962,N_5831,N_4514);
and U9963 (N_9963,N_6148,N_7181);
nor U9964 (N_9964,N_4169,N_5893);
nor U9965 (N_9965,N_4068,N_4116);
or U9966 (N_9966,N_4970,N_7425);
xnor U9967 (N_9967,N_6629,N_5958);
nand U9968 (N_9968,N_6207,N_5715);
or U9969 (N_9969,N_4691,N_5999);
xor U9970 (N_9970,N_4123,N_5597);
or U9971 (N_9971,N_7496,N_5304);
and U9972 (N_9972,N_5115,N_5940);
nand U9973 (N_9973,N_5238,N_6137);
nand U9974 (N_9974,N_5564,N_5204);
nor U9975 (N_9975,N_7322,N_6541);
or U9976 (N_9976,N_7928,N_4410);
nand U9977 (N_9977,N_6531,N_5678);
nand U9978 (N_9978,N_6507,N_4937);
nor U9979 (N_9979,N_6560,N_7579);
nand U9980 (N_9980,N_4705,N_4447);
and U9981 (N_9981,N_7833,N_6986);
nor U9982 (N_9982,N_6669,N_7678);
or U9983 (N_9983,N_7515,N_6076);
xnor U9984 (N_9984,N_7287,N_5452);
nand U9985 (N_9985,N_5548,N_7222);
nand U9986 (N_9986,N_7137,N_7686);
nor U9987 (N_9987,N_6861,N_6292);
nand U9988 (N_9988,N_6300,N_5843);
nand U9989 (N_9989,N_7970,N_6014);
nand U9990 (N_9990,N_4019,N_5561);
nand U9991 (N_9991,N_5206,N_7298);
nor U9992 (N_9992,N_7048,N_5545);
nand U9993 (N_9993,N_6611,N_7478);
nand U9994 (N_9994,N_4932,N_7946);
nand U9995 (N_9995,N_4492,N_7069);
and U9996 (N_9996,N_6824,N_4401);
nand U9997 (N_9997,N_6887,N_5737);
or U9998 (N_9998,N_4668,N_5123);
xnor U9999 (N_9999,N_4197,N_7253);
nor U10000 (N_10000,N_7221,N_6834);
nand U10001 (N_10001,N_4471,N_6016);
nor U10002 (N_10002,N_6919,N_6037);
nor U10003 (N_10003,N_4224,N_6575);
nor U10004 (N_10004,N_7434,N_5243);
and U10005 (N_10005,N_5795,N_5545);
nand U10006 (N_10006,N_7736,N_7728);
nand U10007 (N_10007,N_6714,N_4611);
and U10008 (N_10008,N_7209,N_5695);
xnor U10009 (N_10009,N_5664,N_6752);
nor U10010 (N_10010,N_4196,N_7883);
or U10011 (N_10011,N_4011,N_6464);
or U10012 (N_10012,N_5842,N_4768);
nand U10013 (N_10013,N_7668,N_7594);
nor U10014 (N_10014,N_7192,N_6320);
and U10015 (N_10015,N_4345,N_4783);
xnor U10016 (N_10016,N_6502,N_7345);
and U10017 (N_10017,N_5902,N_4319);
xor U10018 (N_10018,N_7548,N_7260);
nor U10019 (N_10019,N_4507,N_6632);
and U10020 (N_10020,N_7880,N_7422);
nand U10021 (N_10021,N_4838,N_5446);
and U10022 (N_10022,N_4189,N_7809);
xor U10023 (N_10023,N_6853,N_6541);
or U10024 (N_10024,N_4550,N_4385);
or U10025 (N_10025,N_7288,N_6634);
nor U10026 (N_10026,N_7726,N_7386);
and U10027 (N_10027,N_5240,N_6404);
and U10028 (N_10028,N_7599,N_4921);
or U10029 (N_10029,N_4465,N_7666);
or U10030 (N_10030,N_7725,N_5704);
xnor U10031 (N_10031,N_7370,N_6611);
nand U10032 (N_10032,N_7066,N_4661);
and U10033 (N_10033,N_7908,N_6292);
nand U10034 (N_10034,N_5533,N_4115);
or U10035 (N_10035,N_6515,N_4639);
nand U10036 (N_10036,N_6265,N_4952);
nor U10037 (N_10037,N_6990,N_4877);
or U10038 (N_10038,N_7506,N_6511);
nor U10039 (N_10039,N_4287,N_6557);
nand U10040 (N_10040,N_4431,N_7059);
xor U10041 (N_10041,N_5276,N_6345);
or U10042 (N_10042,N_5394,N_7940);
nor U10043 (N_10043,N_5490,N_7595);
xor U10044 (N_10044,N_5825,N_4283);
nor U10045 (N_10045,N_4158,N_6160);
and U10046 (N_10046,N_6890,N_5223);
nor U10047 (N_10047,N_7363,N_6950);
and U10048 (N_10048,N_5196,N_5180);
nand U10049 (N_10049,N_4662,N_6948);
nand U10050 (N_10050,N_5011,N_4330);
nor U10051 (N_10051,N_7636,N_7127);
or U10052 (N_10052,N_6358,N_7053);
nand U10053 (N_10053,N_5016,N_7838);
nand U10054 (N_10054,N_5472,N_7027);
nand U10055 (N_10055,N_4817,N_7769);
nor U10056 (N_10056,N_5533,N_4722);
nor U10057 (N_10057,N_4886,N_6479);
nand U10058 (N_10058,N_7233,N_7355);
or U10059 (N_10059,N_5591,N_6722);
nand U10060 (N_10060,N_7031,N_5831);
nand U10061 (N_10061,N_4997,N_4721);
and U10062 (N_10062,N_5643,N_4835);
and U10063 (N_10063,N_6409,N_6431);
nand U10064 (N_10064,N_5062,N_4798);
and U10065 (N_10065,N_4709,N_5548);
or U10066 (N_10066,N_4148,N_4365);
or U10067 (N_10067,N_7923,N_4084);
nor U10068 (N_10068,N_4504,N_6198);
nor U10069 (N_10069,N_7308,N_7136);
nand U10070 (N_10070,N_6624,N_6014);
nor U10071 (N_10071,N_7790,N_5877);
or U10072 (N_10072,N_5483,N_6210);
or U10073 (N_10073,N_7296,N_4890);
nand U10074 (N_10074,N_7140,N_4343);
or U10075 (N_10075,N_7884,N_4840);
xnor U10076 (N_10076,N_5022,N_7221);
or U10077 (N_10077,N_5619,N_7387);
or U10078 (N_10078,N_4039,N_6257);
nor U10079 (N_10079,N_7000,N_6450);
nor U10080 (N_10080,N_7759,N_5895);
nor U10081 (N_10081,N_6880,N_4381);
nor U10082 (N_10082,N_7065,N_6812);
and U10083 (N_10083,N_4741,N_4405);
nor U10084 (N_10084,N_5691,N_7249);
nor U10085 (N_10085,N_6485,N_6626);
and U10086 (N_10086,N_5460,N_5122);
or U10087 (N_10087,N_4711,N_6776);
and U10088 (N_10088,N_6427,N_4014);
nand U10089 (N_10089,N_4908,N_7179);
nor U10090 (N_10090,N_4694,N_7172);
or U10091 (N_10091,N_7130,N_7694);
and U10092 (N_10092,N_7224,N_4059);
nand U10093 (N_10093,N_7345,N_6449);
and U10094 (N_10094,N_4049,N_7242);
nand U10095 (N_10095,N_6043,N_5583);
nand U10096 (N_10096,N_5532,N_4847);
xnor U10097 (N_10097,N_4028,N_4253);
or U10098 (N_10098,N_5410,N_7708);
or U10099 (N_10099,N_4545,N_5978);
and U10100 (N_10100,N_4017,N_5046);
nor U10101 (N_10101,N_5058,N_4267);
and U10102 (N_10102,N_4130,N_4626);
or U10103 (N_10103,N_6000,N_7049);
nor U10104 (N_10104,N_4334,N_7515);
and U10105 (N_10105,N_7512,N_5049);
xor U10106 (N_10106,N_4740,N_4961);
nor U10107 (N_10107,N_6683,N_4767);
and U10108 (N_10108,N_4830,N_7356);
nor U10109 (N_10109,N_5288,N_5133);
or U10110 (N_10110,N_4851,N_5902);
or U10111 (N_10111,N_5081,N_5995);
or U10112 (N_10112,N_7619,N_4951);
or U10113 (N_10113,N_5458,N_6192);
xor U10114 (N_10114,N_6386,N_6029);
and U10115 (N_10115,N_6506,N_6736);
and U10116 (N_10116,N_7675,N_7751);
nor U10117 (N_10117,N_5427,N_5947);
nor U10118 (N_10118,N_7042,N_4302);
nand U10119 (N_10119,N_4922,N_5364);
xor U10120 (N_10120,N_5542,N_7623);
nor U10121 (N_10121,N_7491,N_4917);
nor U10122 (N_10122,N_7069,N_5235);
or U10123 (N_10123,N_5253,N_4451);
or U10124 (N_10124,N_5116,N_7594);
and U10125 (N_10125,N_6931,N_4397);
nand U10126 (N_10126,N_4749,N_6596);
and U10127 (N_10127,N_7328,N_7099);
or U10128 (N_10128,N_4683,N_5771);
or U10129 (N_10129,N_5054,N_6484);
nand U10130 (N_10130,N_5307,N_7819);
nand U10131 (N_10131,N_7958,N_7720);
or U10132 (N_10132,N_6866,N_6414);
or U10133 (N_10133,N_5768,N_5432);
and U10134 (N_10134,N_5339,N_6530);
nand U10135 (N_10135,N_5006,N_5916);
and U10136 (N_10136,N_4353,N_7385);
and U10137 (N_10137,N_4788,N_4437);
nand U10138 (N_10138,N_6269,N_5914);
nor U10139 (N_10139,N_6819,N_7737);
nor U10140 (N_10140,N_6639,N_5821);
or U10141 (N_10141,N_7938,N_5244);
and U10142 (N_10142,N_6149,N_7473);
or U10143 (N_10143,N_6449,N_7447);
nand U10144 (N_10144,N_6598,N_7346);
or U10145 (N_10145,N_6278,N_4392);
and U10146 (N_10146,N_7565,N_7609);
or U10147 (N_10147,N_6295,N_5609);
or U10148 (N_10148,N_6081,N_4040);
nand U10149 (N_10149,N_4221,N_4602);
and U10150 (N_10150,N_6003,N_6452);
and U10151 (N_10151,N_5893,N_6714);
or U10152 (N_10152,N_4681,N_6792);
xor U10153 (N_10153,N_7968,N_6269);
nand U10154 (N_10154,N_5266,N_7019);
nand U10155 (N_10155,N_5793,N_4473);
nand U10156 (N_10156,N_6877,N_5431);
and U10157 (N_10157,N_5521,N_5269);
and U10158 (N_10158,N_5222,N_6716);
nand U10159 (N_10159,N_7193,N_4835);
or U10160 (N_10160,N_7585,N_4641);
nor U10161 (N_10161,N_7470,N_4796);
or U10162 (N_10162,N_6837,N_5373);
or U10163 (N_10163,N_7424,N_4593);
xor U10164 (N_10164,N_5912,N_4309);
or U10165 (N_10165,N_5541,N_6758);
and U10166 (N_10166,N_5456,N_7941);
nor U10167 (N_10167,N_6268,N_6234);
and U10168 (N_10168,N_5620,N_4842);
and U10169 (N_10169,N_5642,N_5073);
nor U10170 (N_10170,N_5719,N_5800);
and U10171 (N_10171,N_4978,N_5112);
and U10172 (N_10172,N_7512,N_4894);
and U10173 (N_10173,N_6669,N_7316);
xnor U10174 (N_10174,N_7744,N_7526);
nor U10175 (N_10175,N_7590,N_6607);
or U10176 (N_10176,N_4809,N_7507);
or U10177 (N_10177,N_7832,N_7913);
nand U10178 (N_10178,N_6430,N_6414);
nand U10179 (N_10179,N_6226,N_6642);
or U10180 (N_10180,N_6166,N_5250);
and U10181 (N_10181,N_4811,N_6414);
or U10182 (N_10182,N_4823,N_6834);
or U10183 (N_10183,N_5855,N_7796);
nand U10184 (N_10184,N_7834,N_4535);
and U10185 (N_10185,N_4003,N_7661);
or U10186 (N_10186,N_6720,N_7469);
and U10187 (N_10187,N_5042,N_5447);
nor U10188 (N_10188,N_4482,N_4312);
or U10189 (N_10189,N_4032,N_4243);
nor U10190 (N_10190,N_6650,N_7894);
or U10191 (N_10191,N_7820,N_5289);
xnor U10192 (N_10192,N_4435,N_6547);
xor U10193 (N_10193,N_6346,N_5248);
and U10194 (N_10194,N_6171,N_5645);
and U10195 (N_10195,N_4012,N_5538);
and U10196 (N_10196,N_4335,N_4336);
nor U10197 (N_10197,N_5210,N_4078);
or U10198 (N_10198,N_7431,N_5230);
nor U10199 (N_10199,N_7666,N_5327);
xor U10200 (N_10200,N_6940,N_4417);
and U10201 (N_10201,N_7603,N_4408);
nor U10202 (N_10202,N_7911,N_6814);
xor U10203 (N_10203,N_7798,N_4162);
xnor U10204 (N_10204,N_7808,N_7103);
and U10205 (N_10205,N_5349,N_7156);
and U10206 (N_10206,N_6377,N_6881);
nand U10207 (N_10207,N_6877,N_5858);
nand U10208 (N_10208,N_4612,N_7273);
nor U10209 (N_10209,N_4534,N_5593);
nand U10210 (N_10210,N_4340,N_5449);
xor U10211 (N_10211,N_6088,N_5017);
nor U10212 (N_10212,N_5611,N_6411);
or U10213 (N_10213,N_5068,N_6064);
nand U10214 (N_10214,N_6801,N_5443);
or U10215 (N_10215,N_7941,N_5574);
or U10216 (N_10216,N_5008,N_5241);
or U10217 (N_10217,N_7323,N_6435);
nor U10218 (N_10218,N_5354,N_6784);
or U10219 (N_10219,N_4732,N_5039);
or U10220 (N_10220,N_4606,N_4840);
nor U10221 (N_10221,N_7676,N_5495);
nand U10222 (N_10222,N_7426,N_6021);
nand U10223 (N_10223,N_4687,N_6358);
nor U10224 (N_10224,N_4711,N_6567);
nor U10225 (N_10225,N_7266,N_5687);
nor U10226 (N_10226,N_6489,N_7311);
nand U10227 (N_10227,N_4163,N_7768);
and U10228 (N_10228,N_5338,N_5736);
nor U10229 (N_10229,N_4889,N_7803);
xor U10230 (N_10230,N_6423,N_5684);
nor U10231 (N_10231,N_5517,N_4429);
and U10232 (N_10232,N_5914,N_6787);
and U10233 (N_10233,N_5758,N_7064);
xor U10234 (N_10234,N_6344,N_6846);
nand U10235 (N_10235,N_4783,N_5436);
nand U10236 (N_10236,N_5158,N_7103);
xor U10237 (N_10237,N_5825,N_7359);
xor U10238 (N_10238,N_4508,N_7885);
nor U10239 (N_10239,N_6614,N_5188);
or U10240 (N_10240,N_5146,N_7039);
and U10241 (N_10241,N_4742,N_6905);
xnor U10242 (N_10242,N_5869,N_6611);
nand U10243 (N_10243,N_5089,N_6023);
nand U10244 (N_10244,N_7648,N_4380);
or U10245 (N_10245,N_5121,N_4861);
and U10246 (N_10246,N_4050,N_7074);
or U10247 (N_10247,N_6160,N_6900);
nand U10248 (N_10248,N_5767,N_6006);
nand U10249 (N_10249,N_7253,N_4080);
nand U10250 (N_10250,N_6506,N_5866);
nand U10251 (N_10251,N_4886,N_4508);
nand U10252 (N_10252,N_4780,N_6551);
and U10253 (N_10253,N_7421,N_4508);
and U10254 (N_10254,N_5905,N_4859);
or U10255 (N_10255,N_5678,N_7657);
and U10256 (N_10256,N_5611,N_7647);
or U10257 (N_10257,N_6746,N_7342);
nand U10258 (N_10258,N_5939,N_4557);
and U10259 (N_10259,N_7687,N_6647);
nor U10260 (N_10260,N_5297,N_6717);
xnor U10261 (N_10261,N_6090,N_4663);
nor U10262 (N_10262,N_7914,N_4327);
or U10263 (N_10263,N_7622,N_4732);
and U10264 (N_10264,N_5948,N_7628);
nor U10265 (N_10265,N_7870,N_6844);
xnor U10266 (N_10266,N_4296,N_4695);
nand U10267 (N_10267,N_7799,N_4092);
or U10268 (N_10268,N_6782,N_6670);
nand U10269 (N_10269,N_4028,N_6910);
xor U10270 (N_10270,N_4566,N_6148);
and U10271 (N_10271,N_7311,N_5385);
nand U10272 (N_10272,N_7116,N_7684);
nand U10273 (N_10273,N_7715,N_4292);
and U10274 (N_10274,N_5843,N_7392);
nor U10275 (N_10275,N_5635,N_4917);
nor U10276 (N_10276,N_7838,N_7110);
nor U10277 (N_10277,N_4698,N_7233);
and U10278 (N_10278,N_4201,N_4678);
nand U10279 (N_10279,N_6423,N_7617);
nor U10280 (N_10280,N_6778,N_5792);
xnor U10281 (N_10281,N_4076,N_5624);
and U10282 (N_10282,N_5511,N_6594);
or U10283 (N_10283,N_7983,N_5393);
nand U10284 (N_10284,N_5769,N_7646);
nand U10285 (N_10285,N_6698,N_7270);
or U10286 (N_10286,N_6261,N_4728);
xnor U10287 (N_10287,N_4004,N_6088);
and U10288 (N_10288,N_4875,N_5373);
and U10289 (N_10289,N_7988,N_5649);
xnor U10290 (N_10290,N_5712,N_4636);
nor U10291 (N_10291,N_5142,N_7125);
xor U10292 (N_10292,N_7376,N_7712);
or U10293 (N_10293,N_5067,N_5803);
and U10294 (N_10294,N_4945,N_6717);
and U10295 (N_10295,N_7713,N_6211);
and U10296 (N_10296,N_5744,N_5495);
and U10297 (N_10297,N_4176,N_6535);
nand U10298 (N_10298,N_6434,N_5302);
and U10299 (N_10299,N_7221,N_5008);
xnor U10300 (N_10300,N_7456,N_7136);
nor U10301 (N_10301,N_6490,N_4618);
nand U10302 (N_10302,N_6414,N_7934);
nand U10303 (N_10303,N_5541,N_7103);
nor U10304 (N_10304,N_4868,N_7539);
nor U10305 (N_10305,N_6506,N_5903);
and U10306 (N_10306,N_5904,N_7746);
nand U10307 (N_10307,N_6186,N_6420);
nor U10308 (N_10308,N_5490,N_5119);
nor U10309 (N_10309,N_4760,N_4647);
or U10310 (N_10310,N_6755,N_4921);
xnor U10311 (N_10311,N_7199,N_6264);
nor U10312 (N_10312,N_4965,N_4748);
nor U10313 (N_10313,N_4548,N_6674);
xor U10314 (N_10314,N_7218,N_4440);
xor U10315 (N_10315,N_5146,N_4956);
or U10316 (N_10316,N_4740,N_4105);
and U10317 (N_10317,N_5861,N_4222);
xor U10318 (N_10318,N_4043,N_4489);
and U10319 (N_10319,N_7038,N_4941);
nand U10320 (N_10320,N_4403,N_7774);
and U10321 (N_10321,N_7257,N_6544);
and U10322 (N_10322,N_5049,N_6544);
and U10323 (N_10323,N_4036,N_6856);
and U10324 (N_10324,N_4020,N_6486);
nand U10325 (N_10325,N_6831,N_5970);
nand U10326 (N_10326,N_7633,N_5642);
and U10327 (N_10327,N_6500,N_5423);
or U10328 (N_10328,N_5639,N_5501);
or U10329 (N_10329,N_6890,N_4108);
or U10330 (N_10330,N_5839,N_4669);
nand U10331 (N_10331,N_5097,N_6859);
nor U10332 (N_10332,N_7139,N_6069);
and U10333 (N_10333,N_5410,N_4413);
nor U10334 (N_10334,N_5367,N_4283);
or U10335 (N_10335,N_4982,N_6430);
nor U10336 (N_10336,N_5128,N_4465);
nand U10337 (N_10337,N_4383,N_6756);
or U10338 (N_10338,N_5422,N_5211);
nand U10339 (N_10339,N_4910,N_4956);
and U10340 (N_10340,N_5120,N_7376);
and U10341 (N_10341,N_7064,N_5439);
nor U10342 (N_10342,N_6491,N_5144);
and U10343 (N_10343,N_4031,N_7909);
and U10344 (N_10344,N_6424,N_5160);
and U10345 (N_10345,N_6502,N_6057);
nor U10346 (N_10346,N_7915,N_6213);
or U10347 (N_10347,N_5400,N_7134);
nand U10348 (N_10348,N_4546,N_7796);
nand U10349 (N_10349,N_7510,N_6607);
and U10350 (N_10350,N_5871,N_5066);
and U10351 (N_10351,N_7587,N_4806);
nand U10352 (N_10352,N_4530,N_6185);
nand U10353 (N_10353,N_6501,N_5498);
nor U10354 (N_10354,N_5336,N_4861);
nor U10355 (N_10355,N_5975,N_5768);
and U10356 (N_10356,N_4568,N_7782);
nand U10357 (N_10357,N_4110,N_4951);
nand U10358 (N_10358,N_4923,N_6305);
or U10359 (N_10359,N_4120,N_6066);
nor U10360 (N_10360,N_4067,N_6332);
nand U10361 (N_10361,N_5799,N_7577);
and U10362 (N_10362,N_4240,N_4096);
nor U10363 (N_10363,N_7086,N_4788);
nor U10364 (N_10364,N_6290,N_7876);
or U10365 (N_10365,N_5984,N_6635);
nand U10366 (N_10366,N_4608,N_7333);
nand U10367 (N_10367,N_5807,N_4079);
or U10368 (N_10368,N_5376,N_7041);
nor U10369 (N_10369,N_7795,N_6339);
or U10370 (N_10370,N_6938,N_6623);
nand U10371 (N_10371,N_4465,N_7359);
and U10372 (N_10372,N_4286,N_6140);
or U10373 (N_10373,N_7216,N_5808);
nand U10374 (N_10374,N_7146,N_7004);
nor U10375 (N_10375,N_4845,N_5969);
and U10376 (N_10376,N_6036,N_6763);
nand U10377 (N_10377,N_5113,N_5846);
or U10378 (N_10378,N_4258,N_5376);
nor U10379 (N_10379,N_7933,N_5154);
and U10380 (N_10380,N_5547,N_6018);
or U10381 (N_10381,N_6041,N_5987);
or U10382 (N_10382,N_5562,N_7584);
nor U10383 (N_10383,N_6958,N_5258);
and U10384 (N_10384,N_5036,N_7558);
nand U10385 (N_10385,N_6121,N_5587);
nand U10386 (N_10386,N_5145,N_5883);
nand U10387 (N_10387,N_5269,N_6544);
and U10388 (N_10388,N_5153,N_6326);
or U10389 (N_10389,N_7574,N_4013);
or U10390 (N_10390,N_5493,N_4636);
nand U10391 (N_10391,N_6816,N_5848);
xor U10392 (N_10392,N_7249,N_7514);
nor U10393 (N_10393,N_6227,N_7715);
or U10394 (N_10394,N_6003,N_5139);
and U10395 (N_10395,N_5437,N_5898);
and U10396 (N_10396,N_6138,N_4731);
nand U10397 (N_10397,N_5495,N_5208);
nand U10398 (N_10398,N_7995,N_7843);
nand U10399 (N_10399,N_6186,N_5206);
nor U10400 (N_10400,N_7785,N_6284);
nand U10401 (N_10401,N_5708,N_4832);
xnor U10402 (N_10402,N_6208,N_5702);
nor U10403 (N_10403,N_7820,N_5789);
nand U10404 (N_10404,N_5152,N_7176);
and U10405 (N_10405,N_4188,N_4393);
and U10406 (N_10406,N_4031,N_6442);
nor U10407 (N_10407,N_7823,N_7253);
nor U10408 (N_10408,N_7072,N_4992);
nand U10409 (N_10409,N_7988,N_4174);
and U10410 (N_10410,N_4501,N_6184);
nor U10411 (N_10411,N_4876,N_7271);
nor U10412 (N_10412,N_6073,N_4774);
nand U10413 (N_10413,N_7746,N_4128);
and U10414 (N_10414,N_7749,N_7908);
nand U10415 (N_10415,N_7709,N_5402);
and U10416 (N_10416,N_7896,N_6865);
nand U10417 (N_10417,N_7244,N_6178);
and U10418 (N_10418,N_6298,N_4870);
nor U10419 (N_10419,N_4232,N_4872);
xor U10420 (N_10420,N_5625,N_5313);
and U10421 (N_10421,N_5238,N_4371);
nand U10422 (N_10422,N_5137,N_5844);
nor U10423 (N_10423,N_7917,N_4897);
and U10424 (N_10424,N_6135,N_4845);
or U10425 (N_10425,N_4273,N_4994);
and U10426 (N_10426,N_4225,N_7275);
xnor U10427 (N_10427,N_5580,N_5759);
or U10428 (N_10428,N_6459,N_5858);
nand U10429 (N_10429,N_4236,N_6642);
nor U10430 (N_10430,N_4528,N_5273);
or U10431 (N_10431,N_6577,N_6124);
nor U10432 (N_10432,N_6263,N_5413);
nor U10433 (N_10433,N_7940,N_7300);
nand U10434 (N_10434,N_6937,N_7647);
nand U10435 (N_10435,N_5467,N_4341);
and U10436 (N_10436,N_7146,N_7650);
xnor U10437 (N_10437,N_4120,N_4464);
and U10438 (N_10438,N_4130,N_5604);
nand U10439 (N_10439,N_5583,N_7403);
nor U10440 (N_10440,N_5057,N_6510);
and U10441 (N_10441,N_4722,N_7514);
nand U10442 (N_10442,N_5413,N_5804);
nor U10443 (N_10443,N_6130,N_7647);
or U10444 (N_10444,N_4512,N_6226);
xnor U10445 (N_10445,N_5177,N_6757);
nand U10446 (N_10446,N_6047,N_4149);
nand U10447 (N_10447,N_4362,N_6021);
nor U10448 (N_10448,N_7051,N_7689);
or U10449 (N_10449,N_4855,N_5412);
nor U10450 (N_10450,N_7992,N_5654);
or U10451 (N_10451,N_7527,N_4432);
and U10452 (N_10452,N_4315,N_5564);
xor U10453 (N_10453,N_6266,N_7676);
nor U10454 (N_10454,N_6059,N_6868);
and U10455 (N_10455,N_5866,N_6203);
nand U10456 (N_10456,N_5464,N_4569);
nor U10457 (N_10457,N_7688,N_6016);
nand U10458 (N_10458,N_6574,N_5448);
and U10459 (N_10459,N_6395,N_7155);
or U10460 (N_10460,N_4217,N_7289);
and U10461 (N_10461,N_7953,N_4228);
or U10462 (N_10462,N_7711,N_5104);
nand U10463 (N_10463,N_7666,N_6142);
and U10464 (N_10464,N_7028,N_6182);
and U10465 (N_10465,N_6812,N_4120);
and U10466 (N_10466,N_6627,N_5808);
or U10467 (N_10467,N_6262,N_7353);
nand U10468 (N_10468,N_7152,N_6592);
and U10469 (N_10469,N_6050,N_6997);
nand U10470 (N_10470,N_5663,N_4670);
or U10471 (N_10471,N_6615,N_4179);
nor U10472 (N_10472,N_5730,N_7479);
or U10473 (N_10473,N_5882,N_6242);
and U10474 (N_10474,N_5966,N_7066);
nor U10475 (N_10475,N_4125,N_6663);
and U10476 (N_10476,N_7577,N_4707);
or U10477 (N_10477,N_6261,N_5290);
nor U10478 (N_10478,N_4063,N_6515);
xor U10479 (N_10479,N_7164,N_6709);
nand U10480 (N_10480,N_7348,N_4801);
nor U10481 (N_10481,N_7019,N_7353);
nor U10482 (N_10482,N_6723,N_4654);
or U10483 (N_10483,N_5009,N_7695);
nor U10484 (N_10484,N_5093,N_5601);
or U10485 (N_10485,N_4934,N_5173);
nand U10486 (N_10486,N_7967,N_5719);
xor U10487 (N_10487,N_4619,N_7215);
and U10488 (N_10488,N_6273,N_6568);
or U10489 (N_10489,N_4312,N_4121);
and U10490 (N_10490,N_6952,N_6433);
nand U10491 (N_10491,N_6455,N_5730);
nand U10492 (N_10492,N_6043,N_7709);
nor U10493 (N_10493,N_4751,N_7879);
and U10494 (N_10494,N_6174,N_5550);
nand U10495 (N_10495,N_6613,N_5783);
or U10496 (N_10496,N_4696,N_7395);
or U10497 (N_10497,N_7726,N_5650);
and U10498 (N_10498,N_4674,N_6204);
nand U10499 (N_10499,N_4320,N_7410);
nor U10500 (N_10500,N_6358,N_5543);
or U10501 (N_10501,N_5238,N_4785);
nor U10502 (N_10502,N_4800,N_7616);
and U10503 (N_10503,N_4918,N_5708);
and U10504 (N_10504,N_7904,N_6199);
and U10505 (N_10505,N_5000,N_5822);
nor U10506 (N_10506,N_6295,N_5493);
nor U10507 (N_10507,N_7801,N_5182);
nor U10508 (N_10508,N_5686,N_5798);
xor U10509 (N_10509,N_4082,N_6630);
or U10510 (N_10510,N_5215,N_4038);
and U10511 (N_10511,N_4683,N_7624);
and U10512 (N_10512,N_6731,N_4168);
and U10513 (N_10513,N_5932,N_7556);
xnor U10514 (N_10514,N_5175,N_4644);
nand U10515 (N_10515,N_5250,N_4435);
and U10516 (N_10516,N_7182,N_5449);
nor U10517 (N_10517,N_4766,N_6892);
or U10518 (N_10518,N_7724,N_7180);
nor U10519 (N_10519,N_4264,N_6672);
or U10520 (N_10520,N_7042,N_5313);
nor U10521 (N_10521,N_5848,N_6720);
nor U10522 (N_10522,N_5389,N_7804);
or U10523 (N_10523,N_4240,N_5047);
or U10524 (N_10524,N_4752,N_4250);
nand U10525 (N_10525,N_5539,N_6752);
nand U10526 (N_10526,N_7001,N_7724);
and U10527 (N_10527,N_5560,N_4582);
nor U10528 (N_10528,N_7142,N_7805);
and U10529 (N_10529,N_7288,N_4333);
nand U10530 (N_10530,N_4639,N_4860);
nand U10531 (N_10531,N_7018,N_6234);
or U10532 (N_10532,N_6983,N_4416);
or U10533 (N_10533,N_5496,N_4191);
nand U10534 (N_10534,N_7189,N_5591);
nand U10535 (N_10535,N_5221,N_7840);
or U10536 (N_10536,N_5075,N_5320);
nor U10537 (N_10537,N_5269,N_6168);
or U10538 (N_10538,N_7594,N_4895);
and U10539 (N_10539,N_5771,N_6496);
and U10540 (N_10540,N_4009,N_7544);
or U10541 (N_10541,N_7241,N_7957);
nor U10542 (N_10542,N_4484,N_6974);
and U10543 (N_10543,N_4471,N_5660);
nor U10544 (N_10544,N_6805,N_5781);
or U10545 (N_10545,N_7261,N_4662);
and U10546 (N_10546,N_5732,N_4002);
nor U10547 (N_10547,N_6663,N_6559);
and U10548 (N_10548,N_5918,N_4403);
nand U10549 (N_10549,N_6557,N_4124);
nand U10550 (N_10550,N_6142,N_7814);
or U10551 (N_10551,N_4143,N_7836);
or U10552 (N_10552,N_4465,N_6963);
nor U10553 (N_10553,N_5675,N_6515);
and U10554 (N_10554,N_4292,N_4471);
and U10555 (N_10555,N_7660,N_5990);
and U10556 (N_10556,N_5046,N_7640);
and U10557 (N_10557,N_5508,N_7143);
or U10558 (N_10558,N_6941,N_4702);
nand U10559 (N_10559,N_6283,N_7375);
and U10560 (N_10560,N_5054,N_4060);
nor U10561 (N_10561,N_7803,N_5168);
and U10562 (N_10562,N_5036,N_7355);
xnor U10563 (N_10563,N_5730,N_5960);
nand U10564 (N_10564,N_7224,N_4475);
nand U10565 (N_10565,N_4889,N_7724);
and U10566 (N_10566,N_5033,N_4616);
or U10567 (N_10567,N_4297,N_6997);
nand U10568 (N_10568,N_7349,N_4452);
and U10569 (N_10569,N_5524,N_6073);
nand U10570 (N_10570,N_4554,N_6705);
nand U10571 (N_10571,N_4447,N_7940);
nand U10572 (N_10572,N_6430,N_5395);
nand U10573 (N_10573,N_5763,N_7257);
nand U10574 (N_10574,N_6137,N_7273);
and U10575 (N_10575,N_4068,N_5987);
and U10576 (N_10576,N_5330,N_7235);
nor U10577 (N_10577,N_4632,N_7023);
nor U10578 (N_10578,N_5877,N_5532);
nand U10579 (N_10579,N_5596,N_4936);
xor U10580 (N_10580,N_4494,N_5050);
nand U10581 (N_10581,N_7334,N_4745);
or U10582 (N_10582,N_5113,N_4498);
and U10583 (N_10583,N_6515,N_7458);
nand U10584 (N_10584,N_6100,N_6650);
and U10585 (N_10585,N_4544,N_6140);
and U10586 (N_10586,N_7046,N_6107);
nor U10587 (N_10587,N_4801,N_6140);
nand U10588 (N_10588,N_4188,N_6508);
nand U10589 (N_10589,N_5616,N_4402);
and U10590 (N_10590,N_7535,N_7191);
and U10591 (N_10591,N_7731,N_7781);
nor U10592 (N_10592,N_6136,N_5478);
nor U10593 (N_10593,N_4130,N_4109);
nor U10594 (N_10594,N_7453,N_7535);
nand U10595 (N_10595,N_7430,N_7336);
xnor U10596 (N_10596,N_5853,N_6361);
and U10597 (N_10597,N_6926,N_5611);
and U10598 (N_10598,N_6479,N_6060);
nand U10599 (N_10599,N_6291,N_4520);
or U10600 (N_10600,N_6014,N_6073);
or U10601 (N_10601,N_7551,N_5720);
or U10602 (N_10602,N_4858,N_4361);
nand U10603 (N_10603,N_5982,N_6080);
xnor U10604 (N_10604,N_5962,N_5798);
nor U10605 (N_10605,N_5356,N_7881);
xnor U10606 (N_10606,N_6128,N_6192);
nand U10607 (N_10607,N_6715,N_6893);
nand U10608 (N_10608,N_5024,N_6951);
and U10609 (N_10609,N_5017,N_5449);
and U10610 (N_10610,N_7968,N_7929);
nand U10611 (N_10611,N_7243,N_6255);
nand U10612 (N_10612,N_6648,N_5994);
or U10613 (N_10613,N_5105,N_4763);
nand U10614 (N_10614,N_5599,N_7529);
and U10615 (N_10615,N_7952,N_7502);
nand U10616 (N_10616,N_7254,N_5132);
nand U10617 (N_10617,N_7379,N_6850);
and U10618 (N_10618,N_7283,N_5167);
and U10619 (N_10619,N_6117,N_4964);
or U10620 (N_10620,N_5466,N_7556);
nand U10621 (N_10621,N_4588,N_7251);
nand U10622 (N_10622,N_7850,N_4268);
or U10623 (N_10623,N_6301,N_5206);
and U10624 (N_10624,N_4942,N_6427);
xor U10625 (N_10625,N_5838,N_5366);
and U10626 (N_10626,N_4034,N_5980);
or U10627 (N_10627,N_5157,N_6309);
nor U10628 (N_10628,N_6073,N_4052);
nor U10629 (N_10629,N_4821,N_5628);
nor U10630 (N_10630,N_6151,N_4558);
nand U10631 (N_10631,N_7069,N_5296);
nor U10632 (N_10632,N_5814,N_4498);
or U10633 (N_10633,N_4623,N_7295);
and U10634 (N_10634,N_6636,N_4570);
xor U10635 (N_10635,N_7306,N_5785);
and U10636 (N_10636,N_6452,N_7819);
or U10637 (N_10637,N_4942,N_4524);
nand U10638 (N_10638,N_4389,N_6116);
or U10639 (N_10639,N_6229,N_5636);
nor U10640 (N_10640,N_7861,N_6714);
nor U10641 (N_10641,N_4676,N_4041);
and U10642 (N_10642,N_5677,N_7689);
nor U10643 (N_10643,N_4887,N_7044);
nor U10644 (N_10644,N_7568,N_7541);
or U10645 (N_10645,N_6491,N_5671);
nor U10646 (N_10646,N_6792,N_5635);
nor U10647 (N_10647,N_6125,N_5310);
and U10648 (N_10648,N_4843,N_5334);
nand U10649 (N_10649,N_6253,N_7136);
or U10650 (N_10650,N_5905,N_7051);
and U10651 (N_10651,N_4960,N_5886);
and U10652 (N_10652,N_5731,N_5273);
xor U10653 (N_10653,N_5635,N_4294);
or U10654 (N_10654,N_5416,N_7137);
or U10655 (N_10655,N_7384,N_6159);
or U10656 (N_10656,N_4128,N_7277);
nor U10657 (N_10657,N_6503,N_6459);
xnor U10658 (N_10658,N_7722,N_6178);
and U10659 (N_10659,N_4337,N_5669);
nor U10660 (N_10660,N_5469,N_5494);
nor U10661 (N_10661,N_7456,N_5411);
xnor U10662 (N_10662,N_5188,N_4389);
nand U10663 (N_10663,N_4779,N_7623);
nor U10664 (N_10664,N_7572,N_5465);
or U10665 (N_10665,N_5090,N_7402);
and U10666 (N_10666,N_7609,N_4346);
nand U10667 (N_10667,N_4333,N_7286);
or U10668 (N_10668,N_7019,N_5505);
and U10669 (N_10669,N_6697,N_5714);
nand U10670 (N_10670,N_7252,N_6727);
xor U10671 (N_10671,N_7752,N_5775);
and U10672 (N_10672,N_5058,N_4576);
and U10673 (N_10673,N_7789,N_5922);
nor U10674 (N_10674,N_6088,N_5161);
and U10675 (N_10675,N_7555,N_4139);
and U10676 (N_10676,N_5496,N_5804);
nand U10677 (N_10677,N_5059,N_6149);
and U10678 (N_10678,N_7631,N_7669);
or U10679 (N_10679,N_4693,N_5949);
nand U10680 (N_10680,N_7120,N_4757);
nor U10681 (N_10681,N_5851,N_5063);
nor U10682 (N_10682,N_6503,N_5288);
xor U10683 (N_10683,N_6889,N_5586);
xnor U10684 (N_10684,N_5715,N_5424);
nand U10685 (N_10685,N_6753,N_5945);
nor U10686 (N_10686,N_6641,N_7344);
xnor U10687 (N_10687,N_6548,N_5214);
xor U10688 (N_10688,N_4122,N_7476);
nand U10689 (N_10689,N_5637,N_6303);
nand U10690 (N_10690,N_6469,N_6131);
xor U10691 (N_10691,N_5707,N_5840);
or U10692 (N_10692,N_4893,N_5058);
or U10693 (N_10693,N_7711,N_4690);
nor U10694 (N_10694,N_7448,N_4120);
nor U10695 (N_10695,N_4433,N_6647);
and U10696 (N_10696,N_5526,N_7488);
xnor U10697 (N_10697,N_7062,N_5218);
and U10698 (N_10698,N_5187,N_4046);
xor U10699 (N_10699,N_5829,N_6240);
nand U10700 (N_10700,N_4150,N_4069);
nand U10701 (N_10701,N_6686,N_5832);
nor U10702 (N_10702,N_5393,N_4117);
nand U10703 (N_10703,N_5817,N_5582);
and U10704 (N_10704,N_5679,N_6254);
or U10705 (N_10705,N_6093,N_5518);
nor U10706 (N_10706,N_7536,N_7756);
nor U10707 (N_10707,N_4202,N_5217);
and U10708 (N_10708,N_4916,N_7372);
nor U10709 (N_10709,N_5515,N_5170);
and U10710 (N_10710,N_7492,N_6305);
or U10711 (N_10711,N_6290,N_5595);
and U10712 (N_10712,N_6706,N_5408);
and U10713 (N_10713,N_7145,N_5941);
and U10714 (N_10714,N_7888,N_5635);
nor U10715 (N_10715,N_6998,N_5598);
nor U10716 (N_10716,N_4090,N_5391);
xor U10717 (N_10717,N_7510,N_4264);
nor U10718 (N_10718,N_7109,N_4359);
nand U10719 (N_10719,N_7171,N_6199);
and U10720 (N_10720,N_4440,N_7256);
xnor U10721 (N_10721,N_7363,N_7669);
or U10722 (N_10722,N_7203,N_6623);
nor U10723 (N_10723,N_5151,N_6454);
and U10724 (N_10724,N_5353,N_6549);
nor U10725 (N_10725,N_5559,N_6676);
and U10726 (N_10726,N_6680,N_7168);
nand U10727 (N_10727,N_7368,N_4276);
or U10728 (N_10728,N_4480,N_6004);
nand U10729 (N_10729,N_5615,N_5267);
nand U10730 (N_10730,N_7065,N_5782);
nor U10731 (N_10731,N_7689,N_5455);
nand U10732 (N_10732,N_4724,N_6446);
nand U10733 (N_10733,N_5778,N_5357);
nand U10734 (N_10734,N_5015,N_6759);
or U10735 (N_10735,N_4383,N_4413);
and U10736 (N_10736,N_5957,N_7549);
nor U10737 (N_10737,N_6884,N_6080);
or U10738 (N_10738,N_7607,N_5219);
and U10739 (N_10739,N_4962,N_4652);
and U10740 (N_10740,N_6515,N_7574);
nand U10741 (N_10741,N_6930,N_4208);
nor U10742 (N_10742,N_7329,N_7123);
nand U10743 (N_10743,N_4999,N_5231);
xnor U10744 (N_10744,N_5649,N_5781);
and U10745 (N_10745,N_7513,N_4677);
nand U10746 (N_10746,N_4357,N_4651);
or U10747 (N_10747,N_7703,N_5674);
nand U10748 (N_10748,N_6152,N_4335);
nor U10749 (N_10749,N_5501,N_4912);
or U10750 (N_10750,N_6941,N_4732);
and U10751 (N_10751,N_5591,N_5038);
nor U10752 (N_10752,N_5192,N_7591);
and U10753 (N_10753,N_6298,N_6402);
nand U10754 (N_10754,N_5370,N_6004);
or U10755 (N_10755,N_5656,N_6059);
xor U10756 (N_10756,N_4912,N_6952);
nor U10757 (N_10757,N_4497,N_6840);
nand U10758 (N_10758,N_6413,N_7146);
nor U10759 (N_10759,N_5309,N_6280);
nand U10760 (N_10760,N_7061,N_5802);
and U10761 (N_10761,N_7191,N_4515);
and U10762 (N_10762,N_6991,N_7108);
nor U10763 (N_10763,N_5317,N_4863);
nor U10764 (N_10764,N_5254,N_6730);
and U10765 (N_10765,N_7540,N_7351);
or U10766 (N_10766,N_5013,N_4204);
and U10767 (N_10767,N_5375,N_6877);
nor U10768 (N_10768,N_4953,N_4296);
nor U10769 (N_10769,N_4294,N_7346);
and U10770 (N_10770,N_7982,N_5457);
nand U10771 (N_10771,N_7216,N_6675);
or U10772 (N_10772,N_4601,N_7710);
or U10773 (N_10773,N_7638,N_4332);
and U10774 (N_10774,N_4891,N_4810);
xor U10775 (N_10775,N_4619,N_4365);
or U10776 (N_10776,N_5278,N_5631);
and U10777 (N_10777,N_5086,N_4103);
and U10778 (N_10778,N_7356,N_7185);
or U10779 (N_10779,N_5404,N_4047);
and U10780 (N_10780,N_7811,N_6282);
and U10781 (N_10781,N_6009,N_5980);
xnor U10782 (N_10782,N_5405,N_5742);
nor U10783 (N_10783,N_6017,N_4967);
and U10784 (N_10784,N_4632,N_5127);
and U10785 (N_10785,N_4179,N_5159);
nor U10786 (N_10786,N_6924,N_4508);
nor U10787 (N_10787,N_6785,N_5537);
nor U10788 (N_10788,N_4043,N_6448);
and U10789 (N_10789,N_5286,N_6912);
nor U10790 (N_10790,N_6892,N_4490);
or U10791 (N_10791,N_6648,N_5766);
and U10792 (N_10792,N_5356,N_4044);
nand U10793 (N_10793,N_6003,N_5962);
or U10794 (N_10794,N_5430,N_5577);
or U10795 (N_10795,N_4725,N_7309);
and U10796 (N_10796,N_4011,N_7312);
and U10797 (N_10797,N_5138,N_4628);
and U10798 (N_10798,N_4486,N_4752);
nand U10799 (N_10799,N_6491,N_6971);
nor U10800 (N_10800,N_5660,N_7436);
nand U10801 (N_10801,N_7681,N_6137);
xnor U10802 (N_10802,N_4575,N_7496);
xor U10803 (N_10803,N_4257,N_4876);
and U10804 (N_10804,N_4114,N_7863);
or U10805 (N_10805,N_7226,N_7246);
nand U10806 (N_10806,N_7382,N_5586);
xnor U10807 (N_10807,N_4006,N_7426);
nand U10808 (N_10808,N_4664,N_7672);
nand U10809 (N_10809,N_4320,N_7255);
nor U10810 (N_10810,N_7680,N_4692);
nand U10811 (N_10811,N_5056,N_4582);
or U10812 (N_10812,N_4586,N_4546);
nand U10813 (N_10813,N_4578,N_4851);
nand U10814 (N_10814,N_4756,N_6533);
or U10815 (N_10815,N_7139,N_4111);
nor U10816 (N_10816,N_5964,N_6943);
or U10817 (N_10817,N_6031,N_7914);
nand U10818 (N_10818,N_5937,N_7462);
nand U10819 (N_10819,N_4566,N_4439);
and U10820 (N_10820,N_7270,N_5056);
and U10821 (N_10821,N_7913,N_7581);
xor U10822 (N_10822,N_5633,N_7271);
nand U10823 (N_10823,N_7417,N_7948);
nor U10824 (N_10824,N_7109,N_6796);
or U10825 (N_10825,N_6738,N_4736);
and U10826 (N_10826,N_5023,N_4569);
or U10827 (N_10827,N_5364,N_4323);
and U10828 (N_10828,N_5323,N_4676);
xnor U10829 (N_10829,N_6892,N_7478);
and U10830 (N_10830,N_7932,N_5601);
or U10831 (N_10831,N_4074,N_4065);
or U10832 (N_10832,N_6506,N_4762);
nand U10833 (N_10833,N_7790,N_6217);
nand U10834 (N_10834,N_4460,N_4818);
nor U10835 (N_10835,N_7132,N_7735);
nand U10836 (N_10836,N_7541,N_7708);
nand U10837 (N_10837,N_4083,N_4088);
nand U10838 (N_10838,N_6740,N_7407);
or U10839 (N_10839,N_6915,N_7722);
or U10840 (N_10840,N_6254,N_7492);
xor U10841 (N_10841,N_6555,N_4340);
and U10842 (N_10842,N_4868,N_5123);
or U10843 (N_10843,N_5939,N_4867);
nand U10844 (N_10844,N_6160,N_7895);
nor U10845 (N_10845,N_4437,N_4466);
nor U10846 (N_10846,N_4292,N_6373);
nor U10847 (N_10847,N_5034,N_7142);
nand U10848 (N_10848,N_5595,N_5440);
xor U10849 (N_10849,N_4779,N_4458);
or U10850 (N_10850,N_5512,N_5097);
nor U10851 (N_10851,N_4373,N_4770);
and U10852 (N_10852,N_7096,N_7727);
nor U10853 (N_10853,N_6487,N_7566);
or U10854 (N_10854,N_4335,N_7277);
or U10855 (N_10855,N_5230,N_4076);
or U10856 (N_10856,N_7395,N_5515);
and U10857 (N_10857,N_7749,N_5093);
or U10858 (N_10858,N_6689,N_4096);
nor U10859 (N_10859,N_7343,N_6077);
and U10860 (N_10860,N_6369,N_4320);
and U10861 (N_10861,N_7459,N_6953);
or U10862 (N_10862,N_5675,N_4282);
nand U10863 (N_10863,N_7847,N_6973);
xor U10864 (N_10864,N_4536,N_7017);
or U10865 (N_10865,N_5306,N_4938);
nor U10866 (N_10866,N_5696,N_6493);
and U10867 (N_10867,N_7658,N_6145);
and U10868 (N_10868,N_4308,N_5830);
nor U10869 (N_10869,N_5628,N_5188);
and U10870 (N_10870,N_6526,N_4297);
nor U10871 (N_10871,N_4371,N_4948);
and U10872 (N_10872,N_4204,N_4309);
and U10873 (N_10873,N_7778,N_6884);
xor U10874 (N_10874,N_5346,N_5067);
or U10875 (N_10875,N_4059,N_5509);
and U10876 (N_10876,N_7732,N_7776);
xnor U10877 (N_10877,N_4284,N_7730);
and U10878 (N_10878,N_6678,N_4742);
and U10879 (N_10879,N_7422,N_7955);
or U10880 (N_10880,N_6568,N_4141);
nand U10881 (N_10881,N_4890,N_4697);
nor U10882 (N_10882,N_7147,N_4448);
or U10883 (N_10883,N_7750,N_7864);
nand U10884 (N_10884,N_7145,N_6960);
and U10885 (N_10885,N_5397,N_7813);
xor U10886 (N_10886,N_5756,N_4661);
nor U10887 (N_10887,N_6965,N_5375);
nand U10888 (N_10888,N_7718,N_6213);
and U10889 (N_10889,N_5516,N_6043);
nor U10890 (N_10890,N_6963,N_6598);
nor U10891 (N_10891,N_6130,N_6293);
nor U10892 (N_10892,N_7972,N_6465);
xnor U10893 (N_10893,N_4810,N_7207);
xor U10894 (N_10894,N_4290,N_6745);
nand U10895 (N_10895,N_4331,N_7084);
xor U10896 (N_10896,N_4541,N_6065);
nand U10897 (N_10897,N_6775,N_6788);
or U10898 (N_10898,N_5255,N_5562);
xnor U10899 (N_10899,N_5949,N_6856);
and U10900 (N_10900,N_4658,N_4643);
nand U10901 (N_10901,N_6415,N_7712);
or U10902 (N_10902,N_7852,N_5789);
nand U10903 (N_10903,N_7291,N_4706);
or U10904 (N_10904,N_7305,N_4716);
or U10905 (N_10905,N_4971,N_4359);
and U10906 (N_10906,N_7766,N_6664);
nor U10907 (N_10907,N_5130,N_5545);
and U10908 (N_10908,N_6900,N_4932);
or U10909 (N_10909,N_6657,N_7380);
nand U10910 (N_10910,N_4645,N_7293);
nor U10911 (N_10911,N_4723,N_4362);
xor U10912 (N_10912,N_7405,N_6419);
and U10913 (N_10913,N_4963,N_6850);
and U10914 (N_10914,N_6608,N_7683);
nor U10915 (N_10915,N_7462,N_5268);
and U10916 (N_10916,N_7147,N_6914);
or U10917 (N_10917,N_4362,N_6706);
nand U10918 (N_10918,N_4182,N_4590);
nand U10919 (N_10919,N_7999,N_5568);
nor U10920 (N_10920,N_6075,N_7230);
nor U10921 (N_10921,N_6983,N_7789);
and U10922 (N_10922,N_5779,N_4728);
nand U10923 (N_10923,N_4155,N_6075);
nand U10924 (N_10924,N_6293,N_7115);
or U10925 (N_10925,N_7270,N_7848);
or U10926 (N_10926,N_7710,N_5627);
and U10927 (N_10927,N_4237,N_4876);
nand U10928 (N_10928,N_7716,N_4397);
xor U10929 (N_10929,N_4034,N_7665);
and U10930 (N_10930,N_6442,N_4241);
and U10931 (N_10931,N_6402,N_7014);
and U10932 (N_10932,N_4951,N_4973);
or U10933 (N_10933,N_6597,N_4781);
or U10934 (N_10934,N_5977,N_4481);
and U10935 (N_10935,N_5847,N_6934);
nand U10936 (N_10936,N_5278,N_4747);
or U10937 (N_10937,N_6795,N_5393);
xnor U10938 (N_10938,N_4308,N_6040);
nor U10939 (N_10939,N_7576,N_5014);
and U10940 (N_10940,N_4494,N_4846);
nand U10941 (N_10941,N_5127,N_4094);
or U10942 (N_10942,N_5845,N_5620);
and U10943 (N_10943,N_5656,N_5541);
and U10944 (N_10944,N_5084,N_6089);
or U10945 (N_10945,N_6400,N_6656);
nor U10946 (N_10946,N_6255,N_6317);
nor U10947 (N_10947,N_5097,N_4746);
and U10948 (N_10948,N_4394,N_4674);
xnor U10949 (N_10949,N_6724,N_6265);
or U10950 (N_10950,N_6419,N_4221);
and U10951 (N_10951,N_5040,N_5586);
nor U10952 (N_10952,N_4107,N_7970);
and U10953 (N_10953,N_6857,N_6678);
and U10954 (N_10954,N_5714,N_5776);
or U10955 (N_10955,N_7978,N_4281);
nand U10956 (N_10956,N_4349,N_6525);
and U10957 (N_10957,N_5560,N_6183);
and U10958 (N_10958,N_7068,N_4992);
nor U10959 (N_10959,N_4136,N_5427);
and U10960 (N_10960,N_6245,N_5697);
nand U10961 (N_10961,N_4508,N_7648);
nand U10962 (N_10962,N_6720,N_4067);
or U10963 (N_10963,N_7403,N_4289);
or U10964 (N_10964,N_6934,N_5412);
nor U10965 (N_10965,N_6261,N_7982);
nor U10966 (N_10966,N_6830,N_7871);
xor U10967 (N_10967,N_4063,N_5629);
nand U10968 (N_10968,N_6222,N_4747);
or U10969 (N_10969,N_5100,N_4762);
or U10970 (N_10970,N_6936,N_6413);
nand U10971 (N_10971,N_6563,N_6384);
or U10972 (N_10972,N_5745,N_4027);
and U10973 (N_10973,N_5410,N_7305);
or U10974 (N_10974,N_6647,N_7964);
or U10975 (N_10975,N_7112,N_7380);
and U10976 (N_10976,N_5606,N_6507);
nor U10977 (N_10977,N_7174,N_7617);
nand U10978 (N_10978,N_4605,N_4233);
nand U10979 (N_10979,N_7667,N_4978);
nor U10980 (N_10980,N_4139,N_5230);
and U10981 (N_10981,N_7897,N_5641);
or U10982 (N_10982,N_6578,N_5425);
and U10983 (N_10983,N_7432,N_5957);
xnor U10984 (N_10984,N_6546,N_6605);
and U10985 (N_10985,N_6050,N_7421);
nand U10986 (N_10986,N_4368,N_4941);
nor U10987 (N_10987,N_6051,N_5047);
xor U10988 (N_10988,N_4918,N_5577);
nand U10989 (N_10989,N_4583,N_6560);
xor U10990 (N_10990,N_4861,N_7028);
xnor U10991 (N_10991,N_7450,N_4678);
or U10992 (N_10992,N_6708,N_4015);
nor U10993 (N_10993,N_5540,N_4784);
and U10994 (N_10994,N_7568,N_6004);
nand U10995 (N_10995,N_7494,N_4803);
and U10996 (N_10996,N_6114,N_6011);
nand U10997 (N_10997,N_6148,N_7337);
nor U10998 (N_10998,N_5584,N_4974);
or U10999 (N_10999,N_4362,N_6415);
or U11000 (N_11000,N_4240,N_7432);
and U11001 (N_11001,N_4468,N_5386);
nor U11002 (N_11002,N_5041,N_7691);
and U11003 (N_11003,N_5142,N_6562);
nor U11004 (N_11004,N_7300,N_7343);
nor U11005 (N_11005,N_5557,N_6220);
and U11006 (N_11006,N_7839,N_7298);
nor U11007 (N_11007,N_4951,N_6371);
nand U11008 (N_11008,N_4456,N_7753);
and U11009 (N_11009,N_7123,N_5609);
nand U11010 (N_11010,N_4491,N_4421);
nand U11011 (N_11011,N_4623,N_4634);
and U11012 (N_11012,N_6350,N_5205);
and U11013 (N_11013,N_5582,N_4236);
nand U11014 (N_11014,N_6107,N_4493);
or U11015 (N_11015,N_4261,N_5610);
and U11016 (N_11016,N_6274,N_5789);
or U11017 (N_11017,N_7247,N_5994);
nand U11018 (N_11018,N_6055,N_5914);
nor U11019 (N_11019,N_4945,N_5089);
nor U11020 (N_11020,N_6780,N_4077);
nand U11021 (N_11021,N_5016,N_5488);
nor U11022 (N_11022,N_6534,N_7361);
nand U11023 (N_11023,N_5368,N_5645);
nor U11024 (N_11024,N_4262,N_6538);
xnor U11025 (N_11025,N_7288,N_5447);
and U11026 (N_11026,N_5307,N_7422);
nor U11027 (N_11027,N_6914,N_7593);
and U11028 (N_11028,N_6594,N_4238);
nor U11029 (N_11029,N_6488,N_4778);
nor U11030 (N_11030,N_4085,N_4418);
or U11031 (N_11031,N_5472,N_6495);
nand U11032 (N_11032,N_5060,N_4791);
and U11033 (N_11033,N_7569,N_6833);
and U11034 (N_11034,N_7136,N_6494);
nand U11035 (N_11035,N_5649,N_5349);
and U11036 (N_11036,N_6871,N_6231);
and U11037 (N_11037,N_7131,N_5079);
nand U11038 (N_11038,N_7458,N_7015);
nor U11039 (N_11039,N_7356,N_7066);
nand U11040 (N_11040,N_6849,N_7991);
nor U11041 (N_11041,N_7212,N_6113);
or U11042 (N_11042,N_6932,N_7262);
nand U11043 (N_11043,N_4165,N_4357);
nand U11044 (N_11044,N_7091,N_6837);
nor U11045 (N_11045,N_6009,N_4874);
or U11046 (N_11046,N_7359,N_4363);
xor U11047 (N_11047,N_4489,N_4032);
nand U11048 (N_11048,N_6933,N_7357);
xnor U11049 (N_11049,N_7582,N_6603);
nand U11050 (N_11050,N_5305,N_6675);
or U11051 (N_11051,N_4896,N_5301);
nand U11052 (N_11052,N_7394,N_4804);
nor U11053 (N_11053,N_5838,N_6664);
xnor U11054 (N_11054,N_4506,N_7318);
and U11055 (N_11055,N_6492,N_5074);
nand U11056 (N_11056,N_4773,N_6212);
or U11057 (N_11057,N_6681,N_6934);
nor U11058 (N_11058,N_6752,N_4320);
xor U11059 (N_11059,N_6004,N_7649);
and U11060 (N_11060,N_5441,N_7681);
or U11061 (N_11061,N_4880,N_5993);
or U11062 (N_11062,N_7435,N_4865);
nor U11063 (N_11063,N_4002,N_5055);
or U11064 (N_11064,N_7872,N_7032);
nor U11065 (N_11065,N_5486,N_6980);
and U11066 (N_11066,N_6345,N_6874);
nand U11067 (N_11067,N_6257,N_7503);
and U11068 (N_11068,N_5524,N_5822);
or U11069 (N_11069,N_4831,N_5388);
nand U11070 (N_11070,N_7155,N_5445);
nor U11071 (N_11071,N_6698,N_7010);
xnor U11072 (N_11072,N_7623,N_7977);
or U11073 (N_11073,N_4762,N_5439);
or U11074 (N_11074,N_5946,N_5869);
nor U11075 (N_11075,N_7226,N_5592);
nand U11076 (N_11076,N_4268,N_5114);
or U11077 (N_11077,N_4119,N_5003);
nor U11078 (N_11078,N_5141,N_6769);
nor U11079 (N_11079,N_4364,N_6335);
and U11080 (N_11080,N_5419,N_7422);
nor U11081 (N_11081,N_7382,N_4810);
and U11082 (N_11082,N_4334,N_7107);
or U11083 (N_11083,N_6070,N_6729);
or U11084 (N_11084,N_5449,N_7924);
xor U11085 (N_11085,N_7104,N_6066);
or U11086 (N_11086,N_5347,N_4268);
or U11087 (N_11087,N_4271,N_5657);
nor U11088 (N_11088,N_4463,N_4115);
and U11089 (N_11089,N_4668,N_4399);
or U11090 (N_11090,N_4803,N_5032);
nor U11091 (N_11091,N_5033,N_6555);
nor U11092 (N_11092,N_6291,N_6411);
and U11093 (N_11093,N_4975,N_6244);
nor U11094 (N_11094,N_7827,N_7913);
nand U11095 (N_11095,N_6863,N_7962);
nor U11096 (N_11096,N_5876,N_4227);
nand U11097 (N_11097,N_6648,N_7041);
nor U11098 (N_11098,N_7208,N_7968);
or U11099 (N_11099,N_4090,N_7625);
nand U11100 (N_11100,N_7578,N_6624);
or U11101 (N_11101,N_4030,N_6100);
nor U11102 (N_11102,N_7004,N_4065);
nor U11103 (N_11103,N_5179,N_4961);
nand U11104 (N_11104,N_4338,N_5779);
or U11105 (N_11105,N_6137,N_6176);
or U11106 (N_11106,N_4224,N_6078);
and U11107 (N_11107,N_5290,N_6801);
or U11108 (N_11108,N_6277,N_6827);
and U11109 (N_11109,N_4155,N_5831);
or U11110 (N_11110,N_4867,N_4468);
xnor U11111 (N_11111,N_4943,N_6680);
nor U11112 (N_11112,N_5389,N_6426);
or U11113 (N_11113,N_6850,N_6966);
or U11114 (N_11114,N_5093,N_6837);
nand U11115 (N_11115,N_4186,N_6153);
nand U11116 (N_11116,N_5857,N_6526);
and U11117 (N_11117,N_4804,N_6339);
or U11118 (N_11118,N_4669,N_5451);
nor U11119 (N_11119,N_4043,N_4443);
and U11120 (N_11120,N_4285,N_5051);
or U11121 (N_11121,N_6141,N_6219);
and U11122 (N_11122,N_4618,N_7332);
and U11123 (N_11123,N_6414,N_7647);
nand U11124 (N_11124,N_5524,N_7380);
nand U11125 (N_11125,N_5793,N_6519);
and U11126 (N_11126,N_5113,N_5440);
or U11127 (N_11127,N_5278,N_4685);
nor U11128 (N_11128,N_7763,N_4748);
nand U11129 (N_11129,N_4077,N_6881);
and U11130 (N_11130,N_7549,N_6902);
xor U11131 (N_11131,N_6220,N_4426);
nor U11132 (N_11132,N_6152,N_7580);
xnor U11133 (N_11133,N_7406,N_4828);
xnor U11134 (N_11134,N_7385,N_7817);
or U11135 (N_11135,N_6849,N_4578);
or U11136 (N_11136,N_7248,N_4142);
xor U11137 (N_11137,N_5726,N_7621);
and U11138 (N_11138,N_5006,N_5853);
nor U11139 (N_11139,N_5189,N_4737);
nor U11140 (N_11140,N_5941,N_5082);
and U11141 (N_11141,N_6213,N_5888);
and U11142 (N_11142,N_5076,N_6289);
xnor U11143 (N_11143,N_6208,N_4882);
nand U11144 (N_11144,N_5668,N_7270);
or U11145 (N_11145,N_7967,N_6989);
or U11146 (N_11146,N_4054,N_7042);
xor U11147 (N_11147,N_4686,N_7170);
nor U11148 (N_11148,N_4876,N_4297);
or U11149 (N_11149,N_5882,N_5432);
nand U11150 (N_11150,N_6354,N_7644);
nor U11151 (N_11151,N_6055,N_7257);
xnor U11152 (N_11152,N_5558,N_4324);
xor U11153 (N_11153,N_5064,N_6204);
nand U11154 (N_11154,N_5510,N_5052);
nor U11155 (N_11155,N_4998,N_6970);
and U11156 (N_11156,N_5201,N_5497);
or U11157 (N_11157,N_7783,N_7167);
and U11158 (N_11158,N_5005,N_5779);
nand U11159 (N_11159,N_7232,N_4215);
nor U11160 (N_11160,N_4545,N_4620);
nand U11161 (N_11161,N_5773,N_7927);
and U11162 (N_11162,N_7194,N_4080);
nand U11163 (N_11163,N_7125,N_6464);
xnor U11164 (N_11164,N_4993,N_4499);
xnor U11165 (N_11165,N_4521,N_5701);
and U11166 (N_11166,N_7723,N_7192);
nand U11167 (N_11167,N_5294,N_5929);
and U11168 (N_11168,N_5148,N_5008);
and U11169 (N_11169,N_4122,N_4333);
or U11170 (N_11170,N_6308,N_4875);
nand U11171 (N_11171,N_4547,N_4886);
nor U11172 (N_11172,N_4110,N_6403);
xor U11173 (N_11173,N_4349,N_6539);
or U11174 (N_11174,N_6684,N_7327);
and U11175 (N_11175,N_4307,N_4375);
nor U11176 (N_11176,N_5653,N_7344);
and U11177 (N_11177,N_6387,N_7885);
nand U11178 (N_11178,N_5370,N_4712);
xnor U11179 (N_11179,N_7374,N_4144);
nor U11180 (N_11180,N_4475,N_6754);
and U11181 (N_11181,N_4771,N_7639);
nand U11182 (N_11182,N_5022,N_4300);
nor U11183 (N_11183,N_7754,N_6867);
nand U11184 (N_11184,N_4353,N_4164);
nand U11185 (N_11185,N_5106,N_7768);
nand U11186 (N_11186,N_5206,N_4329);
and U11187 (N_11187,N_7499,N_5937);
or U11188 (N_11188,N_5174,N_6125);
nand U11189 (N_11189,N_6735,N_5417);
or U11190 (N_11190,N_4488,N_4980);
nand U11191 (N_11191,N_6634,N_7078);
or U11192 (N_11192,N_7938,N_7078);
or U11193 (N_11193,N_6009,N_7665);
nor U11194 (N_11194,N_7040,N_4650);
and U11195 (N_11195,N_4045,N_6632);
and U11196 (N_11196,N_6733,N_6778);
nor U11197 (N_11197,N_6088,N_5330);
and U11198 (N_11198,N_5688,N_5016);
nor U11199 (N_11199,N_7087,N_7190);
and U11200 (N_11200,N_6612,N_5825);
nand U11201 (N_11201,N_5773,N_4768);
and U11202 (N_11202,N_7568,N_4236);
and U11203 (N_11203,N_7925,N_4800);
xor U11204 (N_11204,N_4426,N_6043);
nand U11205 (N_11205,N_7154,N_6254);
xor U11206 (N_11206,N_7953,N_5055);
nor U11207 (N_11207,N_5852,N_4325);
nor U11208 (N_11208,N_4765,N_6544);
nand U11209 (N_11209,N_7353,N_6702);
nor U11210 (N_11210,N_7970,N_5043);
nor U11211 (N_11211,N_4894,N_4295);
or U11212 (N_11212,N_5111,N_6904);
and U11213 (N_11213,N_5816,N_6471);
and U11214 (N_11214,N_5130,N_4974);
nor U11215 (N_11215,N_4682,N_5011);
nand U11216 (N_11216,N_4635,N_5986);
xor U11217 (N_11217,N_4555,N_4934);
nand U11218 (N_11218,N_5108,N_5781);
or U11219 (N_11219,N_6268,N_7033);
xor U11220 (N_11220,N_6691,N_4004);
nor U11221 (N_11221,N_7477,N_7603);
nand U11222 (N_11222,N_6372,N_5912);
xor U11223 (N_11223,N_4124,N_4456);
or U11224 (N_11224,N_6307,N_5461);
or U11225 (N_11225,N_4318,N_5317);
nor U11226 (N_11226,N_4722,N_6999);
or U11227 (N_11227,N_6570,N_6332);
nand U11228 (N_11228,N_5927,N_6801);
xor U11229 (N_11229,N_5376,N_7236);
nand U11230 (N_11230,N_5355,N_4840);
xnor U11231 (N_11231,N_7917,N_6491);
nor U11232 (N_11232,N_6436,N_5152);
and U11233 (N_11233,N_6692,N_4040);
nand U11234 (N_11234,N_6990,N_4101);
and U11235 (N_11235,N_4279,N_6978);
or U11236 (N_11236,N_7066,N_5909);
xnor U11237 (N_11237,N_6938,N_5923);
or U11238 (N_11238,N_4959,N_6287);
and U11239 (N_11239,N_5760,N_7668);
nor U11240 (N_11240,N_7732,N_7701);
and U11241 (N_11241,N_4251,N_7338);
nand U11242 (N_11242,N_7379,N_7923);
or U11243 (N_11243,N_4627,N_6056);
nor U11244 (N_11244,N_6931,N_5465);
or U11245 (N_11245,N_6944,N_6404);
nor U11246 (N_11246,N_4258,N_5162);
nand U11247 (N_11247,N_6546,N_7624);
nand U11248 (N_11248,N_5224,N_5598);
and U11249 (N_11249,N_6368,N_7481);
xnor U11250 (N_11250,N_6941,N_6368);
nor U11251 (N_11251,N_4151,N_4550);
and U11252 (N_11252,N_6297,N_6534);
nand U11253 (N_11253,N_5827,N_4463);
nor U11254 (N_11254,N_4771,N_7311);
or U11255 (N_11255,N_5331,N_7419);
nand U11256 (N_11256,N_5104,N_5549);
nor U11257 (N_11257,N_6118,N_5476);
and U11258 (N_11258,N_4096,N_7341);
or U11259 (N_11259,N_5900,N_5975);
nor U11260 (N_11260,N_4749,N_5965);
or U11261 (N_11261,N_6463,N_5504);
or U11262 (N_11262,N_4336,N_7651);
nor U11263 (N_11263,N_4950,N_4795);
nand U11264 (N_11264,N_5439,N_5434);
or U11265 (N_11265,N_6301,N_5084);
or U11266 (N_11266,N_4880,N_4672);
nand U11267 (N_11267,N_4614,N_7951);
nand U11268 (N_11268,N_7500,N_5991);
or U11269 (N_11269,N_4659,N_5362);
nand U11270 (N_11270,N_5040,N_6738);
nand U11271 (N_11271,N_5292,N_5538);
and U11272 (N_11272,N_6422,N_7814);
nor U11273 (N_11273,N_5958,N_7540);
nand U11274 (N_11274,N_4575,N_6904);
nor U11275 (N_11275,N_4444,N_5760);
or U11276 (N_11276,N_4817,N_6017);
and U11277 (N_11277,N_4716,N_5587);
and U11278 (N_11278,N_4172,N_7085);
nor U11279 (N_11279,N_7951,N_6509);
nand U11280 (N_11280,N_5652,N_5622);
or U11281 (N_11281,N_4124,N_4107);
nor U11282 (N_11282,N_6366,N_7922);
xor U11283 (N_11283,N_7788,N_4097);
or U11284 (N_11284,N_7308,N_6637);
nand U11285 (N_11285,N_4572,N_5131);
nand U11286 (N_11286,N_6315,N_5051);
or U11287 (N_11287,N_7979,N_6793);
or U11288 (N_11288,N_5677,N_5176);
xor U11289 (N_11289,N_6532,N_6013);
or U11290 (N_11290,N_4279,N_5919);
nand U11291 (N_11291,N_5454,N_5356);
nor U11292 (N_11292,N_4115,N_5227);
nor U11293 (N_11293,N_4277,N_6244);
and U11294 (N_11294,N_4155,N_4434);
nand U11295 (N_11295,N_6174,N_6203);
or U11296 (N_11296,N_7338,N_4576);
or U11297 (N_11297,N_6737,N_6568);
nor U11298 (N_11298,N_6399,N_7622);
nand U11299 (N_11299,N_5088,N_7244);
nand U11300 (N_11300,N_7078,N_6347);
nand U11301 (N_11301,N_6114,N_7258);
and U11302 (N_11302,N_6825,N_7583);
and U11303 (N_11303,N_4855,N_4968);
nand U11304 (N_11304,N_6930,N_6201);
nand U11305 (N_11305,N_5016,N_4921);
or U11306 (N_11306,N_4115,N_7307);
nand U11307 (N_11307,N_5888,N_5640);
nor U11308 (N_11308,N_6174,N_7576);
and U11309 (N_11309,N_5553,N_7668);
nor U11310 (N_11310,N_5456,N_7200);
and U11311 (N_11311,N_5411,N_7681);
and U11312 (N_11312,N_6505,N_5487);
and U11313 (N_11313,N_5979,N_7033);
nand U11314 (N_11314,N_6071,N_6507);
nand U11315 (N_11315,N_7546,N_7396);
nor U11316 (N_11316,N_6522,N_6899);
nor U11317 (N_11317,N_5744,N_7793);
or U11318 (N_11318,N_5125,N_7733);
nor U11319 (N_11319,N_5698,N_7905);
and U11320 (N_11320,N_5068,N_5780);
nand U11321 (N_11321,N_7363,N_4074);
or U11322 (N_11322,N_7549,N_6419);
xor U11323 (N_11323,N_7110,N_4328);
nor U11324 (N_11324,N_6322,N_7397);
nand U11325 (N_11325,N_7471,N_4398);
and U11326 (N_11326,N_7213,N_7927);
and U11327 (N_11327,N_4376,N_7425);
or U11328 (N_11328,N_7477,N_6581);
and U11329 (N_11329,N_7063,N_7896);
nand U11330 (N_11330,N_5243,N_6852);
and U11331 (N_11331,N_7696,N_4933);
or U11332 (N_11332,N_5846,N_5602);
nand U11333 (N_11333,N_6493,N_7362);
nand U11334 (N_11334,N_5468,N_5162);
and U11335 (N_11335,N_5241,N_4825);
nor U11336 (N_11336,N_5752,N_4607);
nor U11337 (N_11337,N_7582,N_7572);
and U11338 (N_11338,N_5004,N_5557);
nor U11339 (N_11339,N_4311,N_7094);
nand U11340 (N_11340,N_7844,N_4197);
nor U11341 (N_11341,N_5442,N_7176);
and U11342 (N_11342,N_4956,N_6081);
and U11343 (N_11343,N_4264,N_7805);
nand U11344 (N_11344,N_6026,N_5150);
nor U11345 (N_11345,N_6088,N_7341);
and U11346 (N_11346,N_5235,N_6545);
nor U11347 (N_11347,N_6724,N_4937);
nor U11348 (N_11348,N_6369,N_5979);
and U11349 (N_11349,N_6728,N_5196);
nor U11350 (N_11350,N_6601,N_7658);
nor U11351 (N_11351,N_7649,N_5736);
and U11352 (N_11352,N_7091,N_4697);
nand U11353 (N_11353,N_5792,N_5206);
nand U11354 (N_11354,N_7726,N_6395);
and U11355 (N_11355,N_7000,N_7001);
nand U11356 (N_11356,N_5698,N_7524);
and U11357 (N_11357,N_5731,N_5320);
or U11358 (N_11358,N_7438,N_6113);
nand U11359 (N_11359,N_4630,N_6656);
nor U11360 (N_11360,N_5178,N_7228);
or U11361 (N_11361,N_6979,N_6392);
or U11362 (N_11362,N_5842,N_4230);
or U11363 (N_11363,N_5933,N_5618);
xnor U11364 (N_11364,N_7717,N_6110);
nor U11365 (N_11365,N_6997,N_4322);
or U11366 (N_11366,N_6682,N_5503);
nor U11367 (N_11367,N_7622,N_7332);
nor U11368 (N_11368,N_6848,N_6390);
xnor U11369 (N_11369,N_6629,N_5578);
nor U11370 (N_11370,N_7956,N_6565);
or U11371 (N_11371,N_4569,N_4105);
nor U11372 (N_11372,N_5182,N_7399);
nand U11373 (N_11373,N_5103,N_4260);
nor U11374 (N_11374,N_7781,N_7923);
or U11375 (N_11375,N_7485,N_4191);
nand U11376 (N_11376,N_6345,N_6500);
and U11377 (N_11377,N_4530,N_7983);
or U11378 (N_11378,N_6177,N_5166);
and U11379 (N_11379,N_5427,N_6334);
or U11380 (N_11380,N_7549,N_5697);
and U11381 (N_11381,N_6159,N_4319);
nor U11382 (N_11382,N_6456,N_7697);
or U11383 (N_11383,N_7885,N_5597);
or U11384 (N_11384,N_5823,N_4115);
and U11385 (N_11385,N_4871,N_6271);
and U11386 (N_11386,N_7091,N_7256);
nor U11387 (N_11387,N_5797,N_7668);
or U11388 (N_11388,N_7483,N_7413);
or U11389 (N_11389,N_6550,N_4630);
nand U11390 (N_11390,N_4121,N_4169);
nor U11391 (N_11391,N_7561,N_7839);
or U11392 (N_11392,N_7771,N_4868);
nor U11393 (N_11393,N_6634,N_4556);
nand U11394 (N_11394,N_7064,N_4263);
nand U11395 (N_11395,N_7251,N_5864);
and U11396 (N_11396,N_6688,N_7387);
xor U11397 (N_11397,N_5624,N_5320);
and U11398 (N_11398,N_4206,N_7600);
or U11399 (N_11399,N_7704,N_6852);
or U11400 (N_11400,N_4525,N_6872);
nor U11401 (N_11401,N_6673,N_5651);
or U11402 (N_11402,N_6967,N_6958);
or U11403 (N_11403,N_6169,N_7647);
or U11404 (N_11404,N_6679,N_4864);
or U11405 (N_11405,N_4827,N_5513);
nor U11406 (N_11406,N_7343,N_6645);
xnor U11407 (N_11407,N_5113,N_7629);
nor U11408 (N_11408,N_7585,N_6601);
or U11409 (N_11409,N_7725,N_4783);
and U11410 (N_11410,N_5949,N_5512);
or U11411 (N_11411,N_6743,N_4012);
nand U11412 (N_11412,N_7834,N_7556);
nand U11413 (N_11413,N_5280,N_7896);
or U11414 (N_11414,N_4587,N_4808);
nor U11415 (N_11415,N_6845,N_6751);
nand U11416 (N_11416,N_6367,N_6704);
and U11417 (N_11417,N_7590,N_5177);
nor U11418 (N_11418,N_7317,N_6195);
nand U11419 (N_11419,N_6744,N_5870);
nand U11420 (N_11420,N_4092,N_5690);
or U11421 (N_11421,N_5458,N_7872);
nand U11422 (N_11422,N_6045,N_7953);
nor U11423 (N_11423,N_7139,N_5510);
and U11424 (N_11424,N_4939,N_7718);
or U11425 (N_11425,N_6158,N_5260);
nand U11426 (N_11426,N_7350,N_4837);
nor U11427 (N_11427,N_5468,N_4947);
nand U11428 (N_11428,N_7313,N_6219);
and U11429 (N_11429,N_4562,N_7502);
and U11430 (N_11430,N_5366,N_7843);
or U11431 (N_11431,N_6657,N_6211);
and U11432 (N_11432,N_7313,N_6925);
or U11433 (N_11433,N_6205,N_4964);
or U11434 (N_11434,N_5108,N_6596);
xor U11435 (N_11435,N_4528,N_5516);
nand U11436 (N_11436,N_5703,N_5809);
xnor U11437 (N_11437,N_4817,N_7258);
nand U11438 (N_11438,N_7068,N_5325);
nand U11439 (N_11439,N_5659,N_6676);
or U11440 (N_11440,N_4555,N_7146);
or U11441 (N_11441,N_6013,N_4544);
nor U11442 (N_11442,N_4303,N_7751);
or U11443 (N_11443,N_4828,N_7931);
or U11444 (N_11444,N_6713,N_4326);
nor U11445 (N_11445,N_5969,N_7773);
and U11446 (N_11446,N_5975,N_4301);
nand U11447 (N_11447,N_7932,N_4362);
xnor U11448 (N_11448,N_5295,N_6713);
or U11449 (N_11449,N_7247,N_4400);
nor U11450 (N_11450,N_4394,N_6690);
or U11451 (N_11451,N_7016,N_7389);
xnor U11452 (N_11452,N_7379,N_4091);
or U11453 (N_11453,N_4486,N_4366);
and U11454 (N_11454,N_5734,N_6715);
or U11455 (N_11455,N_4337,N_7284);
nand U11456 (N_11456,N_5783,N_4331);
nand U11457 (N_11457,N_6292,N_7732);
and U11458 (N_11458,N_6264,N_6200);
or U11459 (N_11459,N_5296,N_4274);
nand U11460 (N_11460,N_7806,N_5206);
or U11461 (N_11461,N_7446,N_5932);
and U11462 (N_11462,N_7716,N_7865);
or U11463 (N_11463,N_5128,N_6940);
and U11464 (N_11464,N_7122,N_4340);
nand U11465 (N_11465,N_4997,N_6555);
nand U11466 (N_11466,N_6178,N_7861);
and U11467 (N_11467,N_7729,N_5168);
nor U11468 (N_11468,N_6513,N_4440);
nor U11469 (N_11469,N_4922,N_7536);
and U11470 (N_11470,N_6923,N_6266);
and U11471 (N_11471,N_6332,N_6281);
nand U11472 (N_11472,N_6618,N_4114);
nor U11473 (N_11473,N_7477,N_7400);
or U11474 (N_11474,N_7357,N_7576);
nand U11475 (N_11475,N_7777,N_4737);
or U11476 (N_11476,N_4273,N_7035);
or U11477 (N_11477,N_7988,N_7182);
and U11478 (N_11478,N_5663,N_7528);
or U11479 (N_11479,N_5510,N_5755);
nor U11480 (N_11480,N_5579,N_6180);
and U11481 (N_11481,N_6109,N_7423);
nor U11482 (N_11482,N_4538,N_4584);
nor U11483 (N_11483,N_4515,N_4421);
nor U11484 (N_11484,N_5942,N_5389);
nand U11485 (N_11485,N_7240,N_5382);
nor U11486 (N_11486,N_5466,N_7128);
nor U11487 (N_11487,N_7041,N_6347);
nor U11488 (N_11488,N_7099,N_5022);
or U11489 (N_11489,N_7691,N_4602);
and U11490 (N_11490,N_5125,N_5620);
nor U11491 (N_11491,N_6380,N_6572);
nand U11492 (N_11492,N_6537,N_6639);
or U11493 (N_11493,N_5307,N_6876);
nor U11494 (N_11494,N_7013,N_5546);
or U11495 (N_11495,N_4436,N_5960);
and U11496 (N_11496,N_5383,N_5246);
nor U11497 (N_11497,N_6723,N_5354);
nand U11498 (N_11498,N_6913,N_5484);
nand U11499 (N_11499,N_5581,N_7767);
nor U11500 (N_11500,N_4466,N_4282);
nand U11501 (N_11501,N_7643,N_5092);
or U11502 (N_11502,N_5054,N_6109);
and U11503 (N_11503,N_6405,N_7166);
xor U11504 (N_11504,N_5191,N_6333);
nor U11505 (N_11505,N_5239,N_7351);
and U11506 (N_11506,N_6580,N_5613);
nor U11507 (N_11507,N_7656,N_7395);
nand U11508 (N_11508,N_4855,N_4154);
nand U11509 (N_11509,N_4393,N_7714);
or U11510 (N_11510,N_4396,N_6959);
and U11511 (N_11511,N_6370,N_4604);
nor U11512 (N_11512,N_5503,N_4496);
or U11513 (N_11513,N_7226,N_6983);
nand U11514 (N_11514,N_7874,N_5046);
or U11515 (N_11515,N_7847,N_5561);
and U11516 (N_11516,N_7650,N_4743);
or U11517 (N_11517,N_7277,N_4018);
or U11518 (N_11518,N_4798,N_7080);
or U11519 (N_11519,N_7646,N_4564);
or U11520 (N_11520,N_7710,N_6834);
nor U11521 (N_11521,N_5204,N_6928);
nand U11522 (N_11522,N_6778,N_6527);
or U11523 (N_11523,N_7578,N_5325);
nand U11524 (N_11524,N_6061,N_6846);
and U11525 (N_11525,N_6482,N_5766);
nand U11526 (N_11526,N_7930,N_4378);
or U11527 (N_11527,N_4177,N_7506);
nand U11528 (N_11528,N_5863,N_5956);
nand U11529 (N_11529,N_4513,N_6462);
nand U11530 (N_11530,N_7083,N_6801);
and U11531 (N_11531,N_4327,N_4358);
xor U11532 (N_11532,N_7236,N_5420);
and U11533 (N_11533,N_5772,N_5620);
xnor U11534 (N_11534,N_5100,N_6598);
nand U11535 (N_11535,N_4139,N_6311);
and U11536 (N_11536,N_4585,N_6003);
nand U11537 (N_11537,N_7783,N_6721);
or U11538 (N_11538,N_6163,N_4303);
nand U11539 (N_11539,N_6883,N_7276);
nand U11540 (N_11540,N_4789,N_4615);
and U11541 (N_11541,N_4926,N_5325);
nor U11542 (N_11542,N_7715,N_4190);
nand U11543 (N_11543,N_7999,N_4601);
and U11544 (N_11544,N_6103,N_4908);
nor U11545 (N_11545,N_7150,N_6436);
nor U11546 (N_11546,N_4260,N_4850);
or U11547 (N_11547,N_7081,N_7634);
and U11548 (N_11548,N_7841,N_4756);
nor U11549 (N_11549,N_7147,N_6368);
and U11550 (N_11550,N_6617,N_6115);
or U11551 (N_11551,N_4355,N_7794);
or U11552 (N_11552,N_4045,N_6906);
and U11553 (N_11553,N_7313,N_7141);
xnor U11554 (N_11554,N_7602,N_5367);
and U11555 (N_11555,N_7618,N_4046);
and U11556 (N_11556,N_4124,N_6659);
and U11557 (N_11557,N_5518,N_6933);
nand U11558 (N_11558,N_7209,N_7275);
or U11559 (N_11559,N_5748,N_7132);
nor U11560 (N_11560,N_5468,N_7294);
nand U11561 (N_11561,N_6008,N_5734);
or U11562 (N_11562,N_7349,N_5499);
or U11563 (N_11563,N_4209,N_7675);
nor U11564 (N_11564,N_4180,N_6493);
or U11565 (N_11565,N_7605,N_6157);
nor U11566 (N_11566,N_5492,N_5087);
or U11567 (N_11567,N_5928,N_5300);
nand U11568 (N_11568,N_4686,N_4284);
nor U11569 (N_11569,N_6030,N_4159);
xor U11570 (N_11570,N_7279,N_4378);
nor U11571 (N_11571,N_6073,N_7901);
and U11572 (N_11572,N_4952,N_6099);
nor U11573 (N_11573,N_5959,N_7739);
nand U11574 (N_11574,N_7540,N_6328);
or U11575 (N_11575,N_7103,N_5690);
nor U11576 (N_11576,N_7502,N_6108);
nor U11577 (N_11577,N_7841,N_4017);
or U11578 (N_11578,N_4924,N_4748);
nand U11579 (N_11579,N_7827,N_6111);
nor U11580 (N_11580,N_4668,N_7866);
nand U11581 (N_11581,N_5187,N_6357);
nor U11582 (N_11582,N_4021,N_6068);
nor U11583 (N_11583,N_7057,N_4977);
and U11584 (N_11584,N_5077,N_4189);
or U11585 (N_11585,N_6721,N_7063);
and U11586 (N_11586,N_7027,N_5401);
nor U11587 (N_11587,N_6881,N_4310);
or U11588 (N_11588,N_7689,N_7925);
xnor U11589 (N_11589,N_7843,N_7086);
and U11590 (N_11590,N_5856,N_6220);
or U11591 (N_11591,N_4754,N_4617);
nor U11592 (N_11592,N_5589,N_4176);
nand U11593 (N_11593,N_4696,N_7495);
xnor U11594 (N_11594,N_4812,N_5474);
xor U11595 (N_11595,N_5219,N_5124);
or U11596 (N_11596,N_7928,N_5188);
or U11597 (N_11597,N_7547,N_7781);
or U11598 (N_11598,N_7835,N_5932);
nor U11599 (N_11599,N_5576,N_6400);
nor U11600 (N_11600,N_6710,N_5575);
and U11601 (N_11601,N_7327,N_7478);
and U11602 (N_11602,N_5578,N_5834);
and U11603 (N_11603,N_7067,N_5841);
nor U11604 (N_11604,N_4929,N_4917);
nor U11605 (N_11605,N_5357,N_5350);
nor U11606 (N_11606,N_6628,N_6660);
or U11607 (N_11607,N_5716,N_4711);
nor U11608 (N_11608,N_6411,N_5860);
or U11609 (N_11609,N_6902,N_7400);
and U11610 (N_11610,N_5669,N_5631);
or U11611 (N_11611,N_5542,N_7659);
or U11612 (N_11612,N_7902,N_5086);
and U11613 (N_11613,N_7602,N_6684);
nor U11614 (N_11614,N_6598,N_6923);
nor U11615 (N_11615,N_7216,N_4697);
and U11616 (N_11616,N_7472,N_7791);
and U11617 (N_11617,N_6627,N_4925);
nand U11618 (N_11618,N_4900,N_6841);
nand U11619 (N_11619,N_5371,N_5663);
and U11620 (N_11620,N_7209,N_4857);
and U11621 (N_11621,N_7916,N_7882);
or U11622 (N_11622,N_4349,N_6936);
or U11623 (N_11623,N_6113,N_4952);
or U11624 (N_11624,N_5703,N_5143);
and U11625 (N_11625,N_7526,N_7089);
xor U11626 (N_11626,N_4379,N_4902);
xor U11627 (N_11627,N_4585,N_6422);
nor U11628 (N_11628,N_7793,N_7275);
nand U11629 (N_11629,N_4510,N_4315);
nand U11630 (N_11630,N_5951,N_7381);
and U11631 (N_11631,N_4508,N_6969);
nor U11632 (N_11632,N_4282,N_7071);
and U11633 (N_11633,N_6968,N_6577);
and U11634 (N_11634,N_7974,N_7906);
or U11635 (N_11635,N_4606,N_6685);
nor U11636 (N_11636,N_5582,N_4490);
or U11637 (N_11637,N_4985,N_4362);
nand U11638 (N_11638,N_6352,N_5790);
nor U11639 (N_11639,N_6862,N_7955);
or U11640 (N_11640,N_4300,N_4582);
nand U11641 (N_11641,N_6432,N_5834);
and U11642 (N_11642,N_6571,N_4174);
xnor U11643 (N_11643,N_6618,N_6258);
and U11644 (N_11644,N_6583,N_6989);
and U11645 (N_11645,N_7972,N_4950);
or U11646 (N_11646,N_5379,N_7044);
nor U11647 (N_11647,N_4138,N_7319);
xor U11648 (N_11648,N_7662,N_7190);
and U11649 (N_11649,N_4213,N_6150);
nor U11650 (N_11650,N_6413,N_4185);
nor U11651 (N_11651,N_4135,N_5034);
nor U11652 (N_11652,N_4887,N_4859);
and U11653 (N_11653,N_5235,N_6311);
and U11654 (N_11654,N_7547,N_5461);
nand U11655 (N_11655,N_4368,N_7550);
and U11656 (N_11656,N_7450,N_5679);
nand U11657 (N_11657,N_7472,N_5512);
and U11658 (N_11658,N_5999,N_6262);
nand U11659 (N_11659,N_4386,N_6135);
nor U11660 (N_11660,N_7309,N_7611);
nor U11661 (N_11661,N_4191,N_7454);
or U11662 (N_11662,N_6122,N_7518);
nor U11663 (N_11663,N_5092,N_7039);
nor U11664 (N_11664,N_6178,N_5997);
and U11665 (N_11665,N_5197,N_7451);
or U11666 (N_11666,N_5175,N_5276);
nor U11667 (N_11667,N_6978,N_7950);
nor U11668 (N_11668,N_6523,N_5941);
and U11669 (N_11669,N_4366,N_4202);
nand U11670 (N_11670,N_5941,N_4734);
and U11671 (N_11671,N_5268,N_6936);
nand U11672 (N_11672,N_6572,N_7258);
nor U11673 (N_11673,N_5638,N_7069);
nand U11674 (N_11674,N_5668,N_7717);
and U11675 (N_11675,N_7997,N_7559);
nand U11676 (N_11676,N_6417,N_7531);
xor U11677 (N_11677,N_6297,N_7363);
and U11678 (N_11678,N_6174,N_7584);
or U11679 (N_11679,N_6293,N_6096);
nand U11680 (N_11680,N_7581,N_5679);
nand U11681 (N_11681,N_4012,N_5593);
nor U11682 (N_11682,N_4773,N_6531);
and U11683 (N_11683,N_5558,N_7124);
or U11684 (N_11684,N_4171,N_6376);
nand U11685 (N_11685,N_6421,N_4012);
or U11686 (N_11686,N_4826,N_4397);
and U11687 (N_11687,N_6399,N_4185);
nand U11688 (N_11688,N_6259,N_5256);
xnor U11689 (N_11689,N_6573,N_7727);
and U11690 (N_11690,N_4563,N_6291);
and U11691 (N_11691,N_5342,N_4084);
nand U11692 (N_11692,N_5203,N_6572);
nand U11693 (N_11693,N_4059,N_5083);
nor U11694 (N_11694,N_7693,N_7045);
or U11695 (N_11695,N_7156,N_7424);
and U11696 (N_11696,N_4127,N_4569);
nand U11697 (N_11697,N_6598,N_4677);
and U11698 (N_11698,N_5581,N_6797);
nor U11699 (N_11699,N_5650,N_5611);
and U11700 (N_11700,N_4791,N_6511);
or U11701 (N_11701,N_5911,N_7956);
xor U11702 (N_11702,N_6296,N_6569);
or U11703 (N_11703,N_6399,N_6988);
nand U11704 (N_11704,N_6127,N_4105);
nand U11705 (N_11705,N_5170,N_4900);
nor U11706 (N_11706,N_4137,N_5679);
or U11707 (N_11707,N_4638,N_7228);
and U11708 (N_11708,N_5453,N_6822);
and U11709 (N_11709,N_5011,N_5436);
nor U11710 (N_11710,N_4847,N_6199);
or U11711 (N_11711,N_4523,N_6572);
nor U11712 (N_11712,N_7307,N_6385);
nor U11713 (N_11713,N_4699,N_5664);
nand U11714 (N_11714,N_5446,N_7327);
nand U11715 (N_11715,N_6613,N_7273);
and U11716 (N_11716,N_4931,N_6652);
or U11717 (N_11717,N_4239,N_5784);
and U11718 (N_11718,N_4306,N_7659);
or U11719 (N_11719,N_6366,N_7725);
nand U11720 (N_11720,N_4156,N_6634);
and U11721 (N_11721,N_6425,N_7768);
nor U11722 (N_11722,N_6275,N_7574);
nand U11723 (N_11723,N_7436,N_5583);
nor U11724 (N_11724,N_6977,N_6518);
nor U11725 (N_11725,N_7536,N_5449);
xor U11726 (N_11726,N_6764,N_4642);
nand U11727 (N_11727,N_5094,N_6161);
or U11728 (N_11728,N_6522,N_7426);
and U11729 (N_11729,N_7838,N_5621);
or U11730 (N_11730,N_5771,N_5660);
and U11731 (N_11731,N_6642,N_6821);
nand U11732 (N_11732,N_4098,N_5410);
or U11733 (N_11733,N_5095,N_6957);
or U11734 (N_11734,N_6841,N_7352);
xor U11735 (N_11735,N_7897,N_6942);
nand U11736 (N_11736,N_7441,N_7983);
nor U11737 (N_11737,N_4344,N_6185);
or U11738 (N_11738,N_6988,N_7406);
or U11739 (N_11739,N_7427,N_5583);
or U11740 (N_11740,N_4688,N_6400);
nand U11741 (N_11741,N_4950,N_6147);
xor U11742 (N_11742,N_5322,N_6583);
or U11743 (N_11743,N_7256,N_6185);
or U11744 (N_11744,N_5812,N_4275);
nand U11745 (N_11745,N_7640,N_6237);
nor U11746 (N_11746,N_5696,N_6021);
xor U11747 (N_11747,N_6134,N_7390);
nor U11748 (N_11748,N_5589,N_7201);
nor U11749 (N_11749,N_4513,N_5057);
xnor U11750 (N_11750,N_5539,N_5807);
nand U11751 (N_11751,N_7171,N_5585);
nand U11752 (N_11752,N_5627,N_4653);
or U11753 (N_11753,N_5714,N_6490);
or U11754 (N_11754,N_5685,N_4314);
xor U11755 (N_11755,N_6054,N_5913);
or U11756 (N_11756,N_4886,N_5411);
and U11757 (N_11757,N_4570,N_5310);
nand U11758 (N_11758,N_6249,N_6900);
nand U11759 (N_11759,N_4561,N_7321);
nand U11760 (N_11760,N_7273,N_4789);
nor U11761 (N_11761,N_4447,N_7959);
nand U11762 (N_11762,N_7920,N_5601);
nand U11763 (N_11763,N_5577,N_5023);
or U11764 (N_11764,N_7567,N_5662);
or U11765 (N_11765,N_6229,N_7864);
or U11766 (N_11766,N_4189,N_5118);
or U11767 (N_11767,N_5173,N_5297);
or U11768 (N_11768,N_4654,N_4635);
nand U11769 (N_11769,N_5303,N_6655);
and U11770 (N_11770,N_7859,N_7849);
and U11771 (N_11771,N_7874,N_4555);
or U11772 (N_11772,N_7096,N_4048);
nand U11773 (N_11773,N_4005,N_6635);
nor U11774 (N_11774,N_4361,N_5748);
and U11775 (N_11775,N_5536,N_7362);
nand U11776 (N_11776,N_7770,N_5569);
nand U11777 (N_11777,N_5899,N_4895);
nor U11778 (N_11778,N_7226,N_6008);
nand U11779 (N_11779,N_7820,N_7963);
xnor U11780 (N_11780,N_5348,N_5597);
or U11781 (N_11781,N_7591,N_5676);
and U11782 (N_11782,N_5733,N_5952);
and U11783 (N_11783,N_5764,N_7744);
and U11784 (N_11784,N_6735,N_6863);
nand U11785 (N_11785,N_6100,N_6653);
nand U11786 (N_11786,N_7261,N_4118);
nand U11787 (N_11787,N_5122,N_7300);
and U11788 (N_11788,N_6831,N_6902);
or U11789 (N_11789,N_7512,N_4506);
nand U11790 (N_11790,N_5697,N_4784);
nor U11791 (N_11791,N_6861,N_4960);
nor U11792 (N_11792,N_4889,N_4941);
and U11793 (N_11793,N_7348,N_5706);
nand U11794 (N_11794,N_7342,N_5372);
nor U11795 (N_11795,N_5922,N_7230);
and U11796 (N_11796,N_6210,N_5657);
and U11797 (N_11797,N_6581,N_4861);
nand U11798 (N_11798,N_6590,N_4869);
and U11799 (N_11799,N_4749,N_5663);
nor U11800 (N_11800,N_4589,N_6978);
nor U11801 (N_11801,N_4348,N_7946);
nand U11802 (N_11802,N_5722,N_7082);
nor U11803 (N_11803,N_6079,N_5481);
nand U11804 (N_11804,N_4093,N_6378);
and U11805 (N_11805,N_4441,N_5043);
nor U11806 (N_11806,N_7475,N_7939);
nor U11807 (N_11807,N_5634,N_5088);
nor U11808 (N_11808,N_6394,N_5964);
nor U11809 (N_11809,N_5255,N_6716);
xor U11810 (N_11810,N_7402,N_6848);
and U11811 (N_11811,N_4399,N_7949);
nor U11812 (N_11812,N_5760,N_7216);
or U11813 (N_11813,N_7142,N_5077);
and U11814 (N_11814,N_7453,N_6303);
nand U11815 (N_11815,N_7167,N_4180);
nand U11816 (N_11816,N_4720,N_7728);
or U11817 (N_11817,N_4148,N_5504);
or U11818 (N_11818,N_4600,N_4762);
and U11819 (N_11819,N_6661,N_6577);
nand U11820 (N_11820,N_6802,N_6340);
nand U11821 (N_11821,N_7702,N_5492);
and U11822 (N_11822,N_5217,N_4591);
and U11823 (N_11823,N_4153,N_7584);
nor U11824 (N_11824,N_4852,N_7098);
or U11825 (N_11825,N_5162,N_7569);
nand U11826 (N_11826,N_4716,N_4329);
and U11827 (N_11827,N_7759,N_7094);
or U11828 (N_11828,N_4533,N_6675);
or U11829 (N_11829,N_5250,N_7793);
nor U11830 (N_11830,N_6042,N_4019);
nor U11831 (N_11831,N_4444,N_5379);
or U11832 (N_11832,N_6640,N_7461);
nand U11833 (N_11833,N_5072,N_6548);
nor U11834 (N_11834,N_6576,N_6548);
or U11835 (N_11835,N_5319,N_5725);
or U11836 (N_11836,N_7520,N_4614);
and U11837 (N_11837,N_5603,N_7732);
and U11838 (N_11838,N_7304,N_6501);
and U11839 (N_11839,N_6857,N_5711);
or U11840 (N_11840,N_5529,N_4453);
nor U11841 (N_11841,N_7588,N_5242);
nand U11842 (N_11842,N_5474,N_4964);
nand U11843 (N_11843,N_6217,N_4894);
or U11844 (N_11844,N_4908,N_4252);
and U11845 (N_11845,N_6506,N_6347);
and U11846 (N_11846,N_4788,N_4298);
or U11847 (N_11847,N_5447,N_5788);
nor U11848 (N_11848,N_4118,N_4739);
nand U11849 (N_11849,N_6144,N_7082);
and U11850 (N_11850,N_5383,N_5015);
nand U11851 (N_11851,N_5061,N_4673);
nand U11852 (N_11852,N_7645,N_5774);
and U11853 (N_11853,N_5504,N_5176);
and U11854 (N_11854,N_4230,N_5864);
or U11855 (N_11855,N_5648,N_5466);
and U11856 (N_11856,N_7695,N_4989);
or U11857 (N_11857,N_4792,N_7354);
xor U11858 (N_11858,N_4241,N_5388);
or U11859 (N_11859,N_5534,N_6428);
and U11860 (N_11860,N_5813,N_6304);
or U11861 (N_11861,N_7015,N_6808);
and U11862 (N_11862,N_5052,N_6435);
nor U11863 (N_11863,N_5034,N_7937);
nor U11864 (N_11864,N_4315,N_7243);
or U11865 (N_11865,N_4549,N_5487);
or U11866 (N_11866,N_4657,N_4319);
nand U11867 (N_11867,N_6357,N_4655);
and U11868 (N_11868,N_5887,N_5759);
or U11869 (N_11869,N_5384,N_4198);
nor U11870 (N_11870,N_6415,N_5671);
or U11871 (N_11871,N_4226,N_4683);
and U11872 (N_11872,N_7722,N_5527);
and U11873 (N_11873,N_5156,N_6622);
nor U11874 (N_11874,N_5504,N_6788);
xnor U11875 (N_11875,N_5205,N_4873);
xor U11876 (N_11876,N_5600,N_6318);
nand U11877 (N_11877,N_5626,N_4660);
or U11878 (N_11878,N_7928,N_6096);
or U11879 (N_11879,N_6666,N_4049);
or U11880 (N_11880,N_7685,N_4668);
nand U11881 (N_11881,N_4663,N_4204);
nand U11882 (N_11882,N_7335,N_6434);
nor U11883 (N_11883,N_6204,N_4002);
or U11884 (N_11884,N_7472,N_6474);
and U11885 (N_11885,N_5956,N_7223);
nor U11886 (N_11886,N_7554,N_6616);
or U11887 (N_11887,N_6133,N_6990);
or U11888 (N_11888,N_4085,N_5374);
nand U11889 (N_11889,N_4448,N_6714);
xor U11890 (N_11890,N_6851,N_4189);
and U11891 (N_11891,N_5476,N_4612);
or U11892 (N_11892,N_5344,N_7273);
nor U11893 (N_11893,N_5283,N_7828);
nor U11894 (N_11894,N_7676,N_6946);
or U11895 (N_11895,N_7811,N_5921);
nor U11896 (N_11896,N_7198,N_6540);
or U11897 (N_11897,N_6553,N_4454);
or U11898 (N_11898,N_6035,N_7033);
xnor U11899 (N_11899,N_4880,N_6150);
nand U11900 (N_11900,N_7823,N_5810);
nor U11901 (N_11901,N_7030,N_4896);
nor U11902 (N_11902,N_4903,N_7397);
nand U11903 (N_11903,N_6727,N_4557);
or U11904 (N_11904,N_6256,N_5717);
nand U11905 (N_11905,N_4373,N_7840);
nor U11906 (N_11906,N_5108,N_6977);
nand U11907 (N_11907,N_4824,N_5747);
nor U11908 (N_11908,N_4336,N_5469);
nand U11909 (N_11909,N_4141,N_7939);
and U11910 (N_11910,N_7157,N_6661);
or U11911 (N_11911,N_5571,N_6929);
nand U11912 (N_11912,N_4078,N_4635);
nor U11913 (N_11913,N_4971,N_6656);
nor U11914 (N_11914,N_4948,N_5663);
nor U11915 (N_11915,N_4019,N_6614);
nor U11916 (N_11916,N_4308,N_6049);
nor U11917 (N_11917,N_7941,N_6250);
or U11918 (N_11918,N_6982,N_6518);
and U11919 (N_11919,N_7238,N_7664);
or U11920 (N_11920,N_7901,N_6330);
and U11921 (N_11921,N_4373,N_4271);
nand U11922 (N_11922,N_5591,N_6041);
and U11923 (N_11923,N_5594,N_5809);
or U11924 (N_11924,N_7545,N_7120);
and U11925 (N_11925,N_6199,N_4212);
or U11926 (N_11926,N_5146,N_4311);
nand U11927 (N_11927,N_5120,N_5136);
or U11928 (N_11928,N_6256,N_5682);
nand U11929 (N_11929,N_7198,N_5197);
xor U11930 (N_11930,N_7483,N_4906);
xor U11931 (N_11931,N_4843,N_4430);
nor U11932 (N_11932,N_6805,N_6166);
nand U11933 (N_11933,N_5299,N_5128);
and U11934 (N_11934,N_6344,N_4298);
nand U11935 (N_11935,N_4943,N_5815);
xnor U11936 (N_11936,N_6094,N_4748);
xor U11937 (N_11937,N_6106,N_5898);
and U11938 (N_11938,N_6089,N_4523);
nor U11939 (N_11939,N_7135,N_5331);
or U11940 (N_11940,N_5780,N_5113);
or U11941 (N_11941,N_4909,N_4866);
nor U11942 (N_11942,N_7547,N_6361);
nand U11943 (N_11943,N_4105,N_6835);
and U11944 (N_11944,N_7910,N_5249);
nor U11945 (N_11945,N_5388,N_5012);
nand U11946 (N_11946,N_5865,N_6370);
or U11947 (N_11947,N_5269,N_5212);
and U11948 (N_11948,N_7935,N_5030);
and U11949 (N_11949,N_7917,N_7434);
and U11950 (N_11950,N_5513,N_5164);
nor U11951 (N_11951,N_5956,N_6430);
nor U11952 (N_11952,N_5293,N_6789);
or U11953 (N_11953,N_7065,N_6339);
nor U11954 (N_11954,N_5945,N_6071);
or U11955 (N_11955,N_5124,N_4980);
nor U11956 (N_11956,N_7557,N_5567);
or U11957 (N_11957,N_6764,N_6805);
nor U11958 (N_11958,N_5191,N_6296);
or U11959 (N_11959,N_5521,N_6005);
nor U11960 (N_11960,N_7434,N_5838);
nor U11961 (N_11961,N_4776,N_4284);
nor U11962 (N_11962,N_4428,N_5015);
or U11963 (N_11963,N_6250,N_6412);
or U11964 (N_11964,N_4401,N_7767);
nand U11965 (N_11965,N_5253,N_5401);
or U11966 (N_11966,N_7794,N_5623);
nand U11967 (N_11967,N_6709,N_6414);
and U11968 (N_11968,N_7015,N_6593);
or U11969 (N_11969,N_6690,N_5951);
nand U11970 (N_11970,N_5610,N_6436);
nand U11971 (N_11971,N_7847,N_6745);
xnor U11972 (N_11972,N_7286,N_6210);
or U11973 (N_11973,N_6422,N_6599);
nor U11974 (N_11974,N_5404,N_6592);
nand U11975 (N_11975,N_7489,N_6961);
and U11976 (N_11976,N_4644,N_4652);
and U11977 (N_11977,N_6502,N_4047);
nor U11978 (N_11978,N_7341,N_5251);
and U11979 (N_11979,N_7565,N_5953);
nor U11980 (N_11980,N_7569,N_6472);
and U11981 (N_11981,N_5026,N_7627);
or U11982 (N_11982,N_4662,N_4811);
xor U11983 (N_11983,N_4543,N_7751);
nor U11984 (N_11984,N_7907,N_7859);
xor U11985 (N_11985,N_7812,N_7135);
nor U11986 (N_11986,N_5246,N_6648);
or U11987 (N_11987,N_5210,N_6291);
and U11988 (N_11988,N_7717,N_6321);
or U11989 (N_11989,N_6742,N_6641);
xnor U11990 (N_11990,N_6385,N_4696);
nor U11991 (N_11991,N_6211,N_5436);
or U11992 (N_11992,N_6052,N_7400);
nand U11993 (N_11993,N_4990,N_5008);
xnor U11994 (N_11994,N_4051,N_4746);
or U11995 (N_11995,N_6722,N_5337);
nand U11996 (N_11996,N_7221,N_4831);
nor U11997 (N_11997,N_4623,N_4565);
or U11998 (N_11998,N_5723,N_6661);
or U11999 (N_11999,N_4105,N_4347);
xor U12000 (N_12000,N_10897,N_11191);
or U12001 (N_12001,N_9710,N_9368);
xnor U12002 (N_12002,N_10328,N_9884);
and U12003 (N_12003,N_8613,N_8597);
or U12004 (N_12004,N_8161,N_10905);
nand U12005 (N_12005,N_11988,N_8453);
nand U12006 (N_12006,N_9495,N_11259);
nor U12007 (N_12007,N_9401,N_8858);
nor U12008 (N_12008,N_11593,N_11324);
or U12009 (N_12009,N_8745,N_9173);
nand U12010 (N_12010,N_11963,N_9905);
nand U12011 (N_12011,N_11475,N_11323);
and U12012 (N_12012,N_9068,N_10592);
xor U12013 (N_12013,N_8705,N_9136);
and U12014 (N_12014,N_8947,N_11087);
nand U12015 (N_12015,N_10194,N_10842);
nand U12016 (N_12016,N_10467,N_11747);
or U12017 (N_12017,N_8490,N_8267);
xor U12018 (N_12018,N_11535,N_8581);
xor U12019 (N_12019,N_8233,N_10498);
nor U12020 (N_12020,N_10189,N_11695);
or U12021 (N_12021,N_10646,N_11224);
and U12022 (N_12022,N_10811,N_9546);
or U12023 (N_12023,N_8016,N_9670);
nor U12024 (N_12024,N_9180,N_11041);
or U12025 (N_12025,N_11335,N_9825);
nand U12026 (N_12026,N_8528,N_11331);
nand U12027 (N_12027,N_11974,N_9599);
nor U12028 (N_12028,N_8417,N_9145);
xor U12029 (N_12029,N_11564,N_8555);
and U12030 (N_12030,N_11135,N_8454);
and U12031 (N_12031,N_10308,N_11295);
nor U12032 (N_12032,N_9780,N_9505);
or U12033 (N_12033,N_10003,N_9121);
or U12034 (N_12034,N_8551,N_8691);
or U12035 (N_12035,N_9523,N_10914);
and U12036 (N_12036,N_9773,N_8464);
xor U12037 (N_12037,N_10954,N_10044);
or U12038 (N_12038,N_10407,N_9272);
and U12039 (N_12039,N_8805,N_8870);
nand U12040 (N_12040,N_10276,N_9630);
or U12041 (N_12041,N_10443,N_9005);
and U12042 (N_12042,N_11557,N_8862);
or U12043 (N_12043,N_10840,N_11085);
or U12044 (N_12044,N_8494,N_10250);
xnor U12045 (N_12045,N_10806,N_8650);
nand U12046 (N_12046,N_8808,N_11687);
or U12047 (N_12047,N_8123,N_8635);
or U12048 (N_12048,N_10005,N_11029);
or U12049 (N_12049,N_8620,N_8220);
and U12050 (N_12050,N_9692,N_10444);
and U12051 (N_12051,N_11631,N_10882);
or U12052 (N_12052,N_8375,N_9685);
or U12053 (N_12053,N_9702,N_11171);
xor U12054 (N_12054,N_10666,N_8480);
or U12055 (N_12055,N_10945,N_11826);
xor U12056 (N_12056,N_9956,N_8859);
xnor U12057 (N_12057,N_10802,N_8582);
nand U12058 (N_12058,N_11227,N_10026);
and U12059 (N_12059,N_9922,N_8338);
nand U12060 (N_12060,N_11009,N_10637);
and U12061 (N_12061,N_11169,N_8628);
xor U12062 (N_12062,N_10821,N_8173);
nand U12063 (N_12063,N_8914,N_8769);
nor U12064 (N_12064,N_8910,N_11855);
or U12065 (N_12065,N_9726,N_10151);
nand U12066 (N_12066,N_10149,N_11678);
and U12067 (N_12067,N_8410,N_8368);
nor U12068 (N_12068,N_10014,N_8950);
xor U12069 (N_12069,N_9674,N_10318);
nand U12070 (N_12070,N_8242,N_8106);
nor U12071 (N_12071,N_9694,N_9170);
and U12072 (N_12072,N_10765,N_9298);
nand U12073 (N_12073,N_8204,N_11370);
and U12074 (N_12074,N_9854,N_8967);
or U12075 (N_12075,N_8447,N_11140);
nor U12076 (N_12076,N_8603,N_9991);
and U12077 (N_12077,N_8543,N_8191);
nor U12078 (N_12078,N_8920,N_9963);
nand U12079 (N_12079,N_9405,N_9666);
nand U12080 (N_12080,N_10873,N_9757);
xnor U12081 (N_12081,N_8339,N_11510);
nor U12082 (N_12082,N_8725,N_11483);
and U12083 (N_12083,N_8326,N_9116);
nor U12084 (N_12084,N_10936,N_11566);
and U12085 (N_12085,N_10346,N_11782);
or U12086 (N_12086,N_8423,N_8665);
or U12087 (N_12087,N_9192,N_9347);
or U12088 (N_12088,N_11646,N_9011);
nor U12089 (N_12089,N_8974,N_8975);
or U12090 (N_12090,N_11480,N_8116);
xnor U12091 (N_12091,N_10870,N_8824);
or U12092 (N_12092,N_11115,N_8874);
xnor U12093 (N_12093,N_9700,N_8653);
and U12094 (N_12094,N_9103,N_9101);
or U12095 (N_12095,N_11552,N_11292);
nand U12096 (N_12096,N_9339,N_10862);
xnor U12097 (N_12097,N_8068,N_8440);
or U12098 (N_12098,N_11351,N_9548);
and U12099 (N_12099,N_9578,N_10772);
nor U12100 (N_12100,N_8625,N_8751);
xnor U12101 (N_12101,N_11032,N_11147);
or U12102 (N_12102,N_10514,N_10174);
or U12103 (N_12103,N_11817,N_10199);
nor U12104 (N_12104,N_8159,N_11904);
and U12105 (N_12105,N_9438,N_9624);
nand U12106 (N_12106,N_11555,N_10904);
and U12107 (N_12107,N_9304,N_8228);
xor U12108 (N_12108,N_9734,N_10434);
nor U12109 (N_12109,N_11304,N_11313);
nand U12110 (N_12110,N_10272,N_9736);
or U12111 (N_12111,N_10283,N_10245);
and U12112 (N_12112,N_10559,N_11458);
nor U12113 (N_12113,N_9222,N_11922);
nand U12114 (N_12114,N_9319,N_9570);
nand U12115 (N_12115,N_9830,N_9099);
and U12116 (N_12116,N_10972,N_8885);
nor U12117 (N_12117,N_8479,N_8119);
or U12118 (N_12118,N_10799,N_9974);
or U12119 (N_12119,N_8046,N_8309);
nor U12120 (N_12120,N_8511,N_9018);
and U12121 (N_12121,N_9021,N_8747);
or U12122 (N_12122,N_11400,N_11494);
nor U12123 (N_12123,N_11832,N_10633);
nor U12124 (N_12124,N_8693,N_10169);
or U12125 (N_12125,N_8938,N_8349);
nand U12126 (N_12126,N_11488,N_10978);
nor U12127 (N_12127,N_8564,N_9445);
nand U12128 (N_12128,N_10251,N_11132);
nand U12129 (N_12129,N_8990,N_11769);
nand U12130 (N_12130,N_9318,N_11680);
or U12131 (N_12131,N_11444,N_8534);
and U12132 (N_12132,N_8413,N_8126);
nor U12133 (N_12133,N_8599,N_9329);
and U12134 (N_12134,N_9739,N_11257);
or U12135 (N_12135,N_11160,N_11692);
and U12136 (N_12136,N_9097,N_10947);
nand U12137 (N_12137,N_11675,N_10817);
or U12138 (N_12138,N_9331,N_8796);
xor U12139 (N_12139,N_11888,N_8029);
or U12140 (N_12140,N_8755,N_9254);
and U12141 (N_12141,N_9551,N_10848);
nor U12142 (N_12142,N_8571,N_8917);
nand U12143 (N_12143,N_9718,N_11317);
nor U12144 (N_12144,N_11641,N_10390);
or U12145 (N_12145,N_11078,N_8017);
nand U12146 (N_12146,N_8221,N_11875);
nor U12147 (N_12147,N_8579,N_9310);
nor U12148 (N_12148,N_8292,N_10565);
nand U12149 (N_12149,N_11663,N_9423);
nor U12150 (N_12150,N_9032,N_11544);
nand U12151 (N_12151,N_11780,N_10237);
nor U12152 (N_12152,N_11380,N_11155);
nand U12153 (N_12153,N_11126,N_9389);
nand U12154 (N_12154,N_8629,N_8592);
nand U12155 (N_12155,N_10773,N_11028);
nor U12156 (N_12156,N_9366,N_8499);
and U12157 (N_12157,N_8364,N_9038);
nor U12158 (N_12158,N_9260,N_8671);
and U12159 (N_12159,N_10373,N_8832);
xnor U12160 (N_12160,N_11397,N_9490);
nand U12161 (N_12161,N_10068,N_8295);
nor U12162 (N_12162,N_10400,N_8380);
nor U12163 (N_12163,N_10607,N_10710);
nor U12164 (N_12164,N_8127,N_9340);
or U12165 (N_12165,N_10542,N_11275);
nor U12166 (N_12166,N_10928,N_8425);
and U12167 (N_12167,N_11670,N_9615);
and U12168 (N_12168,N_10794,N_11860);
or U12169 (N_12169,N_11419,N_9746);
nand U12170 (N_12170,N_11993,N_9699);
and U12171 (N_12171,N_8647,N_8083);
nand U12172 (N_12172,N_11568,N_9189);
or U12173 (N_12173,N_8130,N_9436);
nor U12174 (N_12174,N_8759,N_10223);
nor U12175 (N_12175,N_10152,N_10437);
nor U12176 (N_12176,N_11610,N_9859);
and U12177 (N_12177,N_10035,N_8913);
or U12178 (N_12178,N_11497,N_9671);
or U12179 (N_12179,N_9029,N_8897);
nor U12180 (N_12180,N_11558,N_10186);
or U12181 (N_12181,N_9359,N_11866);
nand U12182 (N_12182,N_9497,N_10497);
nor U12183 (N_12183,N_10638,N_10389);
nor U12184 (N_12184,N_8426,N_11203);
and U12185 (N_12185,N_8789,N_8896);
or U12186 (N_12186,N_10563,N_9480);
or U12187 (N_12187,N_8929,N_10060);
nor U12188 (N_12188,N_11720,N_10111);
nor U12189 (N_12189,N_9634,N_10148);
or U12190 (N_12190,N_8246,N_9434);
and U12191 (N_12191,N_9278,N_11836);
and U12192 (N_12192,N_9918,N_8101);
and U12193 (N_12193,N_10012,N_9194);
nor U12194 (N_12194,N_9747,N_9727);
xor U12195 (N_12195,N_9462,N_8398);
or U12196 (N_12196,N_10341,N_8959);
nor U12197 (N_12197,N_10323,N_11967);
and U12198 (N_12198,N_11429,N_8794);
or U12199 (N_12199,N_8611,N_9297);
and U12200 (N_12200,N_10690,N_9288);
or U12201 (N_12201,N_10475,N_11586);
and U12202 (N_12202,N_11363,N_9186);
and U12203 (N_12203,N_8222,N_8421);
nor U12204 (N_12204,N_10949,N_9740);
and U12205 (N_12205,N_9646,N_9496);
nand U12206 (N_12206,N_11514,N_11759);
nor U12207 (N_12207,N_11755,N_11193);
xnor U12208 (N_12208,N_10360,N_8728);
nor U12209 (N_12209,N_8209,N_9123);
nand U12210 (N_12210,N_11660,N_10278);
and U12211 (N_12211,N_9152,N_9315);
nand U12212 (N_12212,N_9945,N_8873);
nor U12213 (N_12213,N_11760,N_9954);
nand U12214 (N_12214,N_11430,N_10380);
nand U12215 (N_12215,N_10224,N_11045);
or U12216 (N_12216,N_8644,N_9817);
nand U12217 (N_12217,N_11664,N_9861);
or U12218 (N_12218,N_11774,N_9172);
and U12219 (N_12219,N_10852,N_10711);
xnor U12220 (N_12220,N_11353,N_8090);
nor U12221 (N_12221,N_10422,N_8304);
nor U12222 (N_12222,N_8594,N_10062);
or U12223 (N_12223,N_11329,N_10619);
and U12224 (N_12224,N_8356,N_11212);
or U12225 (N_12225,N_8903,N_10902);
and U12226 (N_12226,N_9536,N_11445);
and U12227 (N_12227,N_11576,N_8335);
or U12228 (N_12228,N_10867,N_11813);
and U12229 (N_12229,N_9994,N_8215);
and U12230 (N_12230,N_11017,N_9291);
or U12231 (N_12231,N_11384,N_8631);
nor U12232 (N_12232,N_8855,N_10963);
or U12233 (N_12233,N_11615,N_9990);
nand U12234 (N_12234,N_9308,N_11862);
nor U12235 (N_12235,N_10512,N_11617);
nand U12236 (N_12236,N_10952,N_8839);
nand U12237 (N_12237,N_11473,N_11221);
and U12238 (N_12238,N_10034,N_9568);
and U12239 (N_12239,N_8496,N_9748);
nand U12240 (N_12240,N_9407,N_11044);
nand U12241 (N_12241,N_8030,N_10273);
nand U12242 (N_12242,N_10015,N_10307);
nand U12243 (N_12243,N_10898,N_8863);
nor U12244 (N_12244,N_11711,N_11625);
or U12245 (N_12245,N_9356,N_8009);
nor U12246 (N_12246,N_10743,N_10896);
nand U12247 (N_12247,N_11464,N_11255);
nand U12248 (N_12248,N_9768,N_8442);
or U12249 (N_12249,N_9124,N_9904);
or U12250 (N_12250,N_9062,N_8846);
nand U12251 (N_12251,N_11794,N_10625);
nor U12252 (N_12252,N_11381,N_11603);
and U12253 (N_12253,N_10139,N_10966);
or U12254 (N_12254,N_8879,N_11287);
nor U12255 (N_12255,N_9176,N_8732);
and U12256 (N_12256,N_9798,N_9362);
or U12257 (N_12257,N_9003,N_11966);
and U12258 (N_12258,N_9790,N_11269);
or U12259 (N_12259,N_11919,N_11604);
nor U12260 (N_12260,N_11549,N_8469);
or U12261 (N_12261,N_11097,N_11873);
nand U12262 (N_12262,N_9576,N_9522);
nand U12263 (N_12263,N_9167,N_8062);
or U12264 (N_12264,N_11674,N_9809);
or U12265 (N_12265,N_11136,N_9082);
xnor U12266 (N_12266,N_10198,N_8107);
nand U12267 (N_12267,N_11327,N_8214);
and U12268 (N_12268,N_9007,N_10145);
or U12269 (N_12269,N_10193,N_11242);
nand U12270 (N_12270,N_8450,N_11457);
nor U12271 (N_12271,N_11033,N_11143);
or U12272 (N_12272,N_11144,N_8231);
and U12273 (N_12273,N_10304,N_9885);
xnor U12274 (N_12274,N_11758,N_10819);
and U12275 (N_12275,N_9113,N_10924);
nor U12276 (N_12276,N_8901,N_8283);
nand U12277 (N_12277,N_10253,N_8925);
or U12278 (N_12278,N_9625,N_8580);
and U12279 (N_12279,N_10334,N_8485);
or U12280 (N_12280,N_10961,N_8663);
nor U12281 (N_12281,N_10236,N_11688);
or U12282 (N_12282,N_8767,N_10386);
or U12283 (N_12283,N_11827,N_9935);
nand U12284 (N_12284,N_10737,N_10418);
xor U12285 (N_12285,N_9418,N_10409);
and U12286 (N_12286,N_8097,N_8198);
nand U12287 (N_12287,N_9932,N_11262);
or U12288 (N_12288,N_9849,N_11312);
or U12289 (N_12289,N_8174,N_11086);
xnor U12290 (N_12290,N_11602,N_8666);
xnor U12291 (N_12291,N_10849,N_8812);
nor U12292 (N_12292,N_9792,N_11819);
or U12293 (N_12293,N_9088,N_10994);
xnor U12294 (N_12294,N_10775,N_10384);
and U12295 (N_12295,N_11089,N_10717);
xnor U12296 (N_12296,N_10287,N_8753);
nor U12297 (N_12297,N_10071,N_11180);
xor U12298 (N_12298,N_11772,N_11185);
xor U12299 (N_12299,N_8698,N_10540);
nand U12300 (N_12300,N_9358,N_8113);
nand U12301 (N_12301,N_9326,N_10172);
nor U12302 (N_12302,N_10571,N_8876);
and U12303 (N_12303,N_10326,N_8780);
xor U12304 (N_12304,N_11522,N_9332);
and U12305 (N_12305,N_10686,N_11249);
or U12306 (N_12306,N_10298,N_11525);
or U12307 (N_12307,N_11924,N_10433);
nor U12308 (N_12308,N_9075,N_9962);
nor U12309 (N_12309,N_9508,N_9510);
or U12310 (N_12310,N_11350,N_9870);
nand U12311 (N_12311,N_8646,N_8811);
or U12312 (N_12312,N_9487,N_9380);
or U12313 (N_12313,N_8763,N_10981);
and U12314 (N_12314,N_8752,N_10958);
xor U12315 (N_12315,N_9800,N_9451);
and U12316 (N_12316,N_10385,N_8371);
and U12317 (N_12317,N_10581,N_10312);
or U12318 (N_12318,N_8040,N_9774);
nor U12319 (N_12319,N_11077,N_11509);
or U12320 (N_12320,N_9512,N_8300);
or U12321 (N_12321,N_8537,N_11047);
xnor U12322 (N_12322,N_9146,N_10211);
nand U12323 (N_12323,N_8972,N_9268);
nor U12324 (N_12324,N_9061,N_10241);
or U12325 (N_12325,N_8164,N_8568);
and U12326 (N_12326,N_10510,N_9305);
and U12327 (N_12327,N_11960,N_11054);
nor U12328 (N_12328,N_11465,N_8719);
nand U12329 (N_12329,N_10899,N_9892);
nand U12330 (N_12330,N_9246,N_11513);
xnor U12331 (N_12331,N_9428,N_11561);
or U12332 (N_12332,N_8888,N_9584);
or U12333 (N_12333,N_8773,N_11981);
nor U12334 (N_12334,N_10869,N_10125);
or U12335 (N_12335,N_11986,N_8962);
nor U12336 (N_12336,N_9979,N_9066);
nand U12337 (N_12337,N_8617,N_8388);
nand U12338 (N_12338,N_9993,N_9858);
nand U12339 (N_12339,N_8206,N_8358);
nor U12340 (N_12340,N_11655,N_11040);
nor U12341 (N_12341,N_9472,N_8607);
nor U12342 (N_12342,N_11644,N_8328);
nand U12343 (N_12343,N_11744,N_11463);
nor U12344 (N_12344,N_11074,N_10365);
or U12345 (N_12345,N_9562,N_10080);
and U12346 (N_12346,N_9067,N_10347);
and U12347 (N_12347,N_9275,N_11202);
nand U12348 (N_12348,N_8183,N_8834);
xnor U12349 (N_12349,N_10461,N_9525);
nand U12350 (N_12350,N_11130,N_10118);
and U12351 (N_12351,N_10116,N_8932);
nand U12352 (N_12352,N_11002,N_8995);
or U12353 (N_12353,N_8530,N_11416);
or U12354 (N_12354,N_10160,N_10053);
nor U12355 (N_12355,N_9887,N_8149);
nand U12356 (N_12356,N_11057,N_11863);
or U12357 (N_12357,N_8632,N_10138);
nand U12358 (N_12358,N_11121,N_9683);
or U12359 (N_12359,N_10397,N_8217);
nand U12360 (N_12360,N_10881,N_9925);
or U12361 (N_12361,N_11689,N_11719);
nand U12362 (N_12362,N_11183,N_11196);
or U12363 (N_12363,N_11864,N_10621);
and U12364 (N_12364,N_11885,N_11244);
nand U12365 (N_12365,N_8155,N_10927);
nand U12366 (N_12366,N_9943,N_10156);
and U12367 (N_12367,N_10417,N_10931);
nor U12368 (N_12368,N_9691,N_8318);
or U12369 (N_12369,N_11069,N_10244);
and U12370 (N_12370,N_9144,N_8312);
nand U12371 (N_12371,N_8872,N_8487);
nand U12372 (N_12372,N_10526,N_9457);
and U12373 (N_12373,N_11709,N_8574);
nand U12374 (N_12374,N_8104,N_8777);
or U12375 (N_12375,N_9477,N_10701);
or U12376 (N_12376,N_8188,N_11530);
nor U12377 (N_12377,N_10515,N_11311);
or U12378 (N_12378,N_10212,N_10242);
nor U12379 (N_12379,N_10599,N_8906);
and U12380 (N_12380,N_11371,N_9784);
nand U12381 (N_12381,N_10886,N_11968);
nand U12382 (N_12382,N_8875,N_8782);
nor U12383 (N_12383,N_10089,N_9529);
and U12384 (N_12384,N_11891,N_8094);
nor U12385 (N_12385,N_9533,N_10132);
nand U12386 (N_12386,N_10504,N_8177);
nand U12387 (N_12387,N_8247,N_9530);
nand U12388 (N_12388,N_8802,N_10698);
nor U12389 (N_12389,N_10529,N_8238);
nand U12390 (N_12390,N_11146,N_8385);
and U12391 (N_12391,N_10591,N_11971);
nand U12392 (N_12392,N_11310,N_9470);
nor U12393 (N_12393,N_9009,N_8652);
nand U12394 (N_12394,N_10008,N_11868);
xor U12395 (N_12395,N_10973,N_11050);
nand U12396 (N_12396,N_11879,N_11936);
nand U12397 (N_12397,N_10162,N_11515);
or U12398 (N_12398,N_10336,N_8852);
or U12399 (N_12399,N_9204,N_8393);
and U12400 (N_12400,N_10548,N_11649);
nand U12401 (N_12401,N_9714,N_10471);
nand U12402 (N_12402,N_8694,N_11100);
nand U12403 (N_12403,N_8436,N_10718);
or U12404 (N_12404,N_10166,N_10104);
and U12405 (N_12405,N_10900,N_8189);
nand U12406 (N_12406,N_9862,N_11661);
nor U12407 (N_12407,N_10256,N_10496);
nand U12408 (N_12408,N_10078,N_9863);
nor U12409 (N_12409,N_8501,N_8912);
nor U12410 (N_12410,N_9958,N_9385);
and U12411 (N_12411,N_9988,N_8641);
xnor U12412 (N_12412,N_8791,N_8701);
nand U12413 (N_12413,N_10779,N_8036);
or U12414 (N_12414,N_8809,N_11949);
or U12415 (N_12415,N_11282,N_10480);
and U12416 (N_12416,N_9656,N_11189);
nor U12417 (N_12417,N_11601,N_10262);
nor U12418 (N_12418,N_10602,N_8010);
nor U12419 (N_12419,N_11460,N_9102);
and U12420 (N_12420,N_9803,N_11027);
xor U12421 (N_12421,N_11658,N_11810);
nand U12422 (N_12422,N_10195,N_9920);
nand U12423 (N_12423,N_10383,N_10922);
or U12424 (N_12424,N_11344,N_9968);
xnor U12425 (N_12425,N_9182,N_10431);
and U12426 (N_12426,N_8575,N_10029);
and U12427 (N_12427,N_11787,N_10865);
or U12428 (N_12428,N_10135,N_10031);
nand U12429 (N_12429,N_11975,N_8082);
nor U12430 (N_12430,N_8883,N_8122);
nor U12431 (N_12431,N_10688,N_9588);
nand U12432 (N_12432,N_10321,N_8352);
nor U12433 (N_12433,N_8365,N_11500);
or U12434 (N_12434,N_11293,N_11349);
nand U12435 (N_12435,N_11920,N_11336);
or U12436 (N_12436,N_11438,N_11538);
nand U12437 (N_12437,N_9054,N_10600);
nand U12438 (N_12438,N_9149,N_9360);
and U12439 (N_12439,N_11710,N_11957);
nor U12440 (N_12440,N_11874,N_9402);
nand U12441 (N_12441,N_11520,N_10345);
nand U12442 (N_12442,N_11788,N_11567);
or U12443 (N_12443,N_11783,N_9964);
nand U12444 (N_12444,N_11039,N_10700);
nand U12445 (N_12445,N_9722,N_9788);
or U12446 (N_12446,N_11036,N_10228);
nand U12447 (N_12447,N_8545,N_8979);
or U12448 (N_12448,N_10204,N_8011);
and U12449 (N_12449,N_11172,N_9680);
nor U12450 (N_12450,N_10042,N_10857);
or U12451 (N_12451,N_8379,N_10518);
or U12452 (N_12452,N_8853,N_8366);
or U12453 (N_12453,N_10640,N_11123);
nand U12454 (N_12454,N_9731,N_10609);
and U12455 (N_12455,N_9216,N_11360);
nand U12456 (N_12456,N_8721,N_8151);
nor U12457 (N_12457,N_9353,N_9447);
nor U12458 (N_12458,N_11281,N_9980);
and U12459 (N_12459,N_9491,N_10456);
nor U12460 (N_12460,N_9575,N_10239);
nand U12461 (N_12461,N_11210,N_10675);
nand U12462 (N_12462,N_11153,N_10916);
nand U12463 (N_12463,N_10301,N_10294);
or U12464 (N_12464,N_8656,N_10982);
or U12465 (N_12465,N_11003,N_9707);
nor U12466 (N_12466,N_11447,N_11439);
or U12467 (N_12467,N_11314,N_11048);
or U12468 (N_12468,N_9138,N_10335);
and U12469 (N_12469,N_10703,N_10416);
nand U12470 (N_12470,N_8133,N_9583);
or U12471 (N_12471,N_8648,N_10642);
xnor U12472 (N_12472,N_8482,N_9223);
nor U12473 (N_12473,N_8531,N_9791);
and U12474 (N_12474,N_10082,N_11732);
or U12475 (N_12475,N_8315,N_8240);
and U12476 (N_12476,N_10387,N_11569);
nand U12477 (N_12477,N_11635,N_8243);
nor U12478 (N_12478,N_10233,N_11944);
or U12479 (N_12479,N_11420,N_8195);
nand U12480 (N_12480,N_10179,N_8877);
and U12481 (N_12481,N_8978,N_9764);
or U12482 (N_12482,N_8076,N_10593);
nor U12483 (N_12483,N_10489,N_10750);
and U12484 (N_12484,N_10530,N_10910);
nand U12485 (N_12485,N_11532,N_10115);
xnor U12486 (N_12486,N_8096,N_10894);
and U12487 (N_12487,N_8184,N_11572);
nand U12488 (N_12488,N_8807,N_10788);
nand U12489 (N_12489,N_8958,N_10920);
nand U12490 (N_12490,N_11165,N_10850);
nand U12491 (N_12491,N_11927,N_8668);
nand U12492 (N_12492,N_9659,N_10129);
and U12493 (N_12493,N_11468,N_8712);
or U12494 (N_12494,N_9723,N_10316);
nor U12495 (N_12495,N_10127,N_11984);
nand U12496 (N_12496,N_8079,N_10620);
nor U12497 (N_12497,N_8835,N_9081);
nor U12498 (N_12498,N_11636,N_10230);
and U12499 (N_12499,N_10830,N_8977);
nand U12500 (N_12500,N_11913,N_11179);
and U12501 (N_12501,N_8045,N_11543);
or U12502 (N_12502,N_10369,N_10083);
and U12503 (N_12503,N_10415,N_8506);
nand U12504 (N_12504,N_11230,N_9585);
and U12505 (N_12505,N_10753,N_11706);
or U12506 (N_12506,N_8329,N_11776);
nor U12507 (N_12507,N_9341,N_10655);
nand U12508 (N_12508,N_10579,N_9134);
nand U12509 (N_12509,N_8542,N_9064);
nand U12510 (N_12510,N_8176,N_10259);
and U12511 (N_12511,N_8324,N_9433);
nand U12512 (N_12512,N_8291,N_11869);
nand U12513 (N_12513,N_10353,N_8614);
and U12514 (N_12514,N_8508,N_11516);
nor U12515 (N_12515,N_10742,N_9015);
nor U12516 (N_12516,N_9944,N_11723);
and U12517 (N_12517,N_8738,N_11847);
xor U12518 (N_12518,N_9055,N_10822);
or U12519 (N_12519,N_11200,N_9166);
nor U12520 (N_12520,N_9786,N_10613);
and U12521 (N_12521,N_9732,N_11433);
nor U12522 (N_12522,N_8071,N_10329);
nor U12523 (N_12523,N_8615,N_9865);
and U12524 (N_12524,N_10095,N_9716);
nor U12525 (N_12525,N_11948,N_10872);
nor U12526 (N_12526,N_8347,N_8355);
and U12527 (N_12527,N_11124,N_8952);
or U12528 (N_12528,N_8946,N_11995);
xnor U12529 (N_12529,N_11777,N_10673);
or U12530 (N_12530,N_10054,N_11990);
nand U12531 (N_12531,N_9388,N_9730);
and U12532 (N_12532,N_10634,N_10134);
and U12533 (N_12533,N_11778,N_11748);
nor U12534 (N_12534,N_9627,N_10511);
xor U12535 (N_12535,N_8092,N_9911);
or U12536 (N_12536,N_9663,N_8717);
and U12537 (N_12537,N_9902,N_11129);
nor U12538 (N_12538,N_8923,N_8658);
xnor U12539 (N_12539,N_9839,N_10785);
and U12540 (N_12540,N_9030,N_8192);
and U12541 (N_12541,N_9371,N_11091);
nand U12542 (N_12542,N_10909,N_9330);
or U12543 (N_12543,N_8667,N_11745);
or U12544 (N_12544,N_10495,N_10516);
and U12545 (N_12545,N_11846,N_11816);
or U12546 (N_12546,N_8443,N_11222);
nand U12547 (N_12547,N_11897,N_11682);
and U12548 (N_12548,N_11521,N_9745);
and U12549 (N_12549,N_11359,N_8716);
or U12550 (N_12550,N_8486,N_8218);
nor U12551 (N_12551,N_8004,N_8591);
and U12552 (N_12552,N_10689,N_11870);
nand U12553 (N_12553,N_11942,N_10841);
and U12554 (N_12554,N_10059,N_8241);
nor U12555 (N_12555,N_11440,N_10110);
or U12556 (N_12556,N_9787,N_9650);
or U12557 (N_12557,N_11935,N_10871);
and U12558 (N_12558,N_11321,N_11253);
and U12559 (N_12559,N_8919,N_9996);
nand U12560 (N_12560,N_11906,N_10331);
and U12561 (N_12561,N_10942,N_10731);
xnor U12562 (N_12562,N_11609,N_9468);
nor U12563 (N_12563,N_10953,N_10074);
or U12564 (N_12564,N_10378,N_9153);
or U12565 (N_12565,N_9531,N_9789);
or U12566 (N_12566,N_10680,N_11930);
or U12567 (N_12567,N_11952,N_11983);
nand U12568 (N_12568,N_9386,N_10541);
and U12569 (N_12569,N_8626,N_10804);
and U12570 (N_12570,N_9601,N_11411);
nor U12571 (N_12571,N_10838,N_10716);
and U12572 (N_12572,N_11111,N_9012);
nand U12573 (N_12573,N_11004,N_11241);
nor U12574 (N_12574,N_10793,N_10427);
and U12575 (N_12575,N_10258,N_11233);
and U12576 (N_12576,N_8232,N_8182);
or U12577 (N_12577,N_8168,N_8664);
or U12578 (N_12578,N_11037,N_10096);
and U12579 (N_12579,N_10975,N_9159);
xnor U12580 (N_12580,N_9724,N_11818);
nand U12581 (N_12581,N_10476,N_9024);
nor U12582 (N_12582,N_11341,N_8084);
nor U12583 (N_12583,N_11899,N_11587);
or U12584 (N_12584,N_8507,N_8609);
nand U12585 (N_12585,N_8181,N_10248);
and U12586 (N_12586,N_10812,N_8585);
and U12587 (N_12587,N_10315,N_8005);
or U12588 (N_12588,N_9795,N_11094);
and U12589 (N_12589,N_8019,N_9236);
and U12590 (N_12590,N_11734,N_11539);
and U12591 (N_12591,N_9987,N_11346);
nor U12592 (N_12592,N_8984,N_11795);
xnor U12593 (N_12593,N_11613,N_8089);
and U12594 (N_12594,N_8829,N_9377);
nand U12595 (N_12595,N_10574,N_10375);
nand U12596 (N_12596,N_11596,N_11340);
and U12597 (N_12597,N_8078,N_8899);
and U12598 (N_12598,N_8788,N_10807);
or U12599 (N_12599,N_10488,N_8223);
nand U12600 (N_12600,N_8560,N_10553);
and U12601 (N_12601,N_10800,N_11694);
or U12602 (N_12602,N_11628,N_9534);
nand U12603 (N_12603,N_10671,N_8774);
and U12604 (N_12604,N_11630,N_9429);
or U12605 (N_12605,N_11102,N_8341);
nor U12606 (N_12606,N_9453,N_11162);
nor U12607 (N_12607,N_10452,N_11965);
and U12608 (N_12608,N_11962,N_8766);
nor U12609 (N_12609,N_10482,N_11061);
and U12610 (N_12610,N_8120,N_11157);
and U12611 (N_12611,N_10568,N_9779);
nor U12612 (N_12612,N_8471,N_10877);
nand U12613 (N_12613,N_8602,N_10996);
and U12614 (N_12614,N_8025,N_10660);
nand U12615 (N_12615,N_8535,N_11398);
or U12616 (N_12616,N_10252,N_9290);
xor U12617 (N_12617,N_11900,N_10608);
or U12618 (N_12618,N_11797,N_8171);
xor U12619 (N_12619,N_11401,N_11226);
and U12620 (N_12620,N_11452,N_11629);
nand U12621 (N_12621,N_11092,N_11947);
or U12622 (N_12622,N_10458,N_9020);
or U12623 (N_12623,N_9617,N_9978);
nand U12624 (N_12624,N_11339,N_8420);
nand U12625 (N_12625,N_10943,N_9077);
or U12626 (N_12626,N_9203,N_11645);
or U12627 (N_12627,N_11347,N_8154);
and U12628 (N_12628,N_8115,N_9794);
nor U12629 (N_12629,N_10022,N_9889);
xnor U12630 (N_12630,N_10491,N_10967);
or U12631 (N_12631,N_11796,N_8836);
or U12632 (N_12632,N_11638,N_11206);
nor U12633 (N_12633,N_8605,N_8512);
nand U12634 (N_12634,N_11757,N_9215);
xor U12635 (N_12635,N_8230,N_8726);
nor U12636 (N_12636,N_10605,N_10687);
and U12637 (N_12637,N_8822,N_11838);
or U12638 (N_12638,N_9065,N_11978);
and U12639 (N_12639,N_8265,N_11182);
nor U12640 (N_12640,N_9394,N_10647);
or U12641 (N_12641,N_8271,N_8202);
or U12642 (N_12642,N_10645,N_11823);
and U12643 (N_12643,N_11698,N_11116);
and U12644 (N_12644,N_8996,N_11884);
or U12645 (N_12645,N_8953,N_9100);
and U12646 (N_12646,N_8418,N_10187);
xnor U12647 (N_12647,N_10837,N_10835);
or U12648 (N_12648,N_9831,N_11422);
or U12649 (N_12649,N_8199,N_11739);
or U12650 (N_12650,N_8757,N_9289);
nand U12651 (N_12651,N_11570,N_10843);
and U12652 (N_12652,N_10024,N_8044);
nor U12653 (N_12653,N_9752,N_10282);
or U12654 (N_12654,N_9384,N_11276);
nor U12655 (N_12655,N_11379,N_8890);
xor U12656 (N_12656,N_11937,N_9783);
nor U12657 (N_12657,N_9509,N_10159);
or U12658 (N_12658,N_8484,N_11098);
or U12659 (N_12659,N_8077,N_8103);
nor U12660 (N_12660,N_8032,N_9008);
xor U12661 (N_12661,N_9957,N_8927);
xnor U12662 (N_12662,N_8710,N_10618);
nor U12663 (N_12663,N_8998,N_8465);
xnor U12664 (N_12664,N_10858,N_10921);
nand U12665 (N_12665,N_9452,N_10623);
or U12666 (N_12666,N_9456,N_10522);
xnor U12667 (N_12667,N_11595,N_8724);
nor U12668 (N_12668,N_10445,N_10722);
and U12669 (N_12669,N_9619,N_10847);
nor U12670 (N_12670,N_8634,N_11681);
and U12671 (N_12671,N_8039,N_10930);
or U12672 (N_12672,N_11015,N_10006);
and U12673 (N_12673,N_10227,N_8124);
and U12674 (N_12674,N_8987,N_10465);
nor U12675 (N_12675,N_8298,N_8638);
nand U12676 (N_12676,N_8734,N_9390);
or U12677 (N_12677,N_9160,N_10057);
nor U12678 (N_12678,N_11671,N_10317);
nand U12679 (N_12679,N_8604,N_9237);
nor U12680 (N_12680,N_8640,N_11302);
or U12681 (N_12681,N_8532,N_8702);
and U12682 (N_12682,N_9177,N_9799);
or U12683 (N_12683,N_11970,N_8153);
or U12684 (N_12684,N_10485,N_10755);
or U12685 (N_12685,N_8053,N_10203);
nor U12686 (N_12686,N_8207,N_10154);
and U12687 (N_12687,N_9899,N_9728);
or U12688 (N_12688,N_8105,N_9912);
xnor U12689 (N_12689,N_9414,N_11656);
or U12690 (N_12690,N_10000,N_11926);
and U12691 (N_12691,N_10912,N_10697);
nand U12692 (N_12692,N_9374,N_10810);
and U12693 (N_12693,N_11955,N_11762);
nor U12694 (N_12694,N_9971,N_10192);
xnor U12695 (N_12695,N_9063,N_9191);
and U12696 (N_12696,N_10435,N_11134);
xnor U12697 (N_12697,N_9776,N_10049);
nand U12698 (N_12698,N_8973,N_8114);
or U12699 (N_12699,N_11600,N_10890);
or U12700 (N_12700,N_10826,N_11731);
and U12701 (N_12701,N_8048,N_8563);
nor U12702 (N_12702,N_9096,N_11043);
nor U12703 (N_12703,N_9179,N_10693);
nand U12704 (N_12704,N_10643,N_8966);
xnor U12705 (N_12705,N_9869,N_10560);
nor U12706 (N_12706,N_8956,N_8803);
and U12707 (N_12707,N_10342,N_11019);
and U12708 (N_12708,N_8612,N_10558);
nor U12709 (N_12709,N_11119,N_9301);
nor U12710 (N_12710,N_11857,N_10460);
and U12711 (N_12711,N_11145,N_10780);
nand U12712 (N_12712,N_11940,N_11889);
nand U12713 (N_12713,N_10064,N_10532);
nor U12714 (N_12714,N_8431,N_9547);
and U12715 (N_12715,N_9527,N_10293);
or U12716 (N_12716,N_9606,N_10932);
or U12717 (N_12717,N_8567,N_11607);
and U12718 (N_12718,N_8374,N_11770);
nand U12719 (N_12719,N_9110,N_8688);
nor U12720 (N_12720,N_11842,N_8302);
and U12721 (N_12721,N_11956,N_10338);
nand U12722 (N_12722,N_8708,N_11767);
and U12723 (N_12723,N_11163,N_10712);
or U12724 (N_12724,N_8529,N_8306);
and U12725 (N_12725,N_9367,N_10085);
xnor U12726 (N_12726,N_9621,N_8210);
nor U12727 (N_12727,N_11712,N_10100);
nor U12728 (N_12728,N_9439,N_10584);
nand U12729 (N_12729,N_10533,N_8110);
and U12730 (N_12730,N_11168,N_8143);
nor U12731 (N_12731,N_8284,N_10255);
nand U12732 (N_12732,N_8384,N_8842);
and U12733 (N_12733,N_11910,N_9594);
and U12734 (N_12734,N_11096,N_9306);
or U12735 (N_12735,N_8985,N_9992);
or U12736 (N_12736,N_9190,N_11699);
and U12737 (N_12737,N_8034,N_10575);
nand U12738 (N_12738,N_10449,N_9473);
or U12739 (N_12739,N_8438,N_8681);
nor U12740 (N_12740,N_8185,N_11672);
and U12741 (N_12741,N_11038,N_9195);
and U12742 (N_12742,N_8557,N_11443);
and U12743 (N_12743,N_11425,N_9856);
nor U12744 (N_12744,N_8804,N_10513);
nand U12745 (N_12745,N_9459,N_10521);
nor U12746 (N_12746,N_8226,N_9498);
xnor U12747 (N_12747,N_9913,N_8363);
xnor U12748 (N_12748,N_10137,N_10401);
and U12749 (N_12749,N_10539,N_11161);
and U12750 (N_12750,N_11159,N_11547);
or U12751 (N_12751,N_10839,N_10289);
nand U12752 (N_12752,N_10320,N_10564);
nand U12753 (N_12753,N_8488,N_9878);
and U12754 (N_12754,N_9766,N_11368);
or U12755 (N_12755,N_8986,N_10379);
or U12756 (N_12756,N_8093,N_9678);
nand U12757 (N_12757,N_9403,N_10457);
nor U12758 (N_12758,N_9285,N_9155);
nand U12759 (N_12759,N_10503,N_9515);
nor U12760 (N_12760,N_9567,N_9524);
nand U12761 (N_12761,N_9313,N_8150);
nor U12762 (N_12762,N_8406,N_11580);
and U12763 (N_12763,N_8273,N_11178);
nand U12764 (N_12764,N_8100,N_9711);
and U12765 (N_12765,N_10790,N_8997);
xor U12766 (N_12766,N_9091,N_9936);
and U12767 (N_12767,N_8935,N_11517);
and U12768 (N_12768,N_8274,N_8981);
nand U12769 (N_12769,N_9261,N_11352);
and U12770 (N_12770,N_11598,N_9112);
nand U12771 (N_12771,N_9541,N_11858);
nor U12772 (N_12772,N_8411,N_11238);
xnor U12773 (N_12773,N_10454,N_9597);
nor U12774 (N_12774,N_9408,N_9034);
nand U12775 (N_12775,N_10413,N_8718);
and U12776 (N_12776,N_10028,N_8012);
xor U12777 (N_12777,N_11691,N_10769);
nand U12778 (N_12778,N_10791,N_11199);
nor U12779 (N_12779,N_11477,N_9325);
and U12780 (N_12780,N_11454,N_10414);
or U12781 (N_12781,N_9645,N_10164);
and U12782 (N_12782,N_10598,N_11839);
nor U12783 (N_12783,N_10508,N_8636);
or U12784 (N_12784,N_9269,N_11492);
nor U12785 (N_12785,N_11373,N_11791);
nor U12786 (N_12786,N_9872,N_9629);
nor U12787 (N_12787,N_9516,N_10405);
or U12788 (N_12788,N_9983,N_10279);
and U12789 (N_12789,N_8419,N_8026);
nand U12790 (N_12790,N_9244,N_8166);
nand U12791 (N_12791,N_10709,N_11156);
nor U12792 (N_12792,N_9682,N_8387);
and U12793 (N_12793,N_11026,N_10831);
or U12794 (N_12794,N_10120,N_9975);
xor U12795 (N_12795,N_11343,N_8907);
or U12796 (N_12796,N_8275,N_10885);
and U12797 (N_12797,N_10167,N_8722);
nand U12798 (N_12798,N_8502,N_8942);
or U12799 (N_12799,N_11127,N_10299);
or U12800 (N_12800,N_10959,N_11456);
and U12801 (N_12801,N_8827,N_9908);
xnor U12802 (N_12802,N_9493,N_11807);
or U12803 (N_12803,N_9611,N_11081);
nor U12804 (N_12804,N_10190,N_10968);
xnor U12805 (N_12805,N_11118,N_8065);
or U12806 (N_12806,N_8186,N_10724);
and U12807 (N_12807,N_8483,N_8918);
nor U12808 (N_12808,N_11431,N_11441);
nor U12809 (N_12809,N_9098,N_8703);
and U12810 (N_12810,N_11845,N_9046);
or U12811 (N_12811,N_8964,N_10399);
and U12812 (N_12812,N_8939,N_9104);
nor U12813 (N_12813,N_8474,N_10941);
nor U12814 (N_12814,N_11991,N_8099);
or U12815 (N_12815,N_10573,N_9235);
or U12816 (N_12816,N_9848,N_11880);
nand U12817 (N_12817,N_9837,N_9295);
and U12818 (N_12818,N_8960,N_8407);
nor U12819 (N_12819,N_10538,N_10844);
nand U12820 (N_12820,N_10260,N_9614);
nand U12821 (N_12821,N_10184,N_9070);
xor U12822 (N_12822,N_11637,N_11432);
or U12823 (N_12823,N_10784,N_10892);
nand U12824 (N_12824,N_11388,N_9397);
and U12825 (N_12825,N_8331,N_11358);
or U12826 (N_12826,N_11284,N_10880);
nand U12827 (N_12827,N_10906,N_11740);
xor U12828 (N_12828,N_10663,N_9906);
and U12829 (N_12829,N_9782,N_9616);
and U12830 (N_12830,N_11274,N_10469);
nor U12831 (N_12831,N_8513,N_10216);
or U12832 (N_12832,N_11651,N_8672);
nand U12833 (N_12833,N_9517,N_9970);
nor U12834 (N_12834,N_10090,N_9379);
nand U12835 (N_12835,N_9805,N_10537);
and U12836 (N_12836,N_9760,N_9263);
and U12837 (N_12837,N_10310,N_11562);
and U12838 (N_12838,N_10578,N_9514);
nor U12839 (N_12839,N_10188,N_8768);
nor U12840 (N_12840,N_9874,N_8795);
and U12841 (N_12841,N_9336,N_10297);
and U12842 (N_12842,N_9639,N_8816);
and U12843 (N_12843,N_11484,N_10381);
and U12844 (N_12844,N_9701,N_11559);
or U12845 (N_12845,N_8608,N_9137);
and U12846 (N_12846,N_11065,N_11348);
nor U12847 (N_12847,N_8540,N_10550);
nand U12848 (N_12848,N_10453,N_8922);
or U12849 (N_12849,N_11451,N_8351);
and U12850 (N_12850,N_11149,N_9814);
nand U12851 (N_12851,N_8649,N_11726);
nand U12852 (N_12852,N_11020,N_8448);
and U12853 (N_12853,N_8313,N_11938);
and U12854 (N_12854,N_10410,N_11652);
nand U12855 (N_12855,N_9412,N_8424);
nor U12856 (N_12856,N_8258,N_11413);
or U12857 (N_12857,N_11526,N_8911);
or U12858 (N_12858,N_8301,N_11434);
nand U12859 (N_12859,N_10708,N_9506);
nor U12860 (N_12860,N_8337,N_11702);
xor U12861 (N_12861,N_8976,N_11152);
and U12862 (N_12862,N_8362,N_10756);
xnor U12863 (N_12863,N_8837,N_8539);
xnor U12864 (N_12864,N_11404,N_10639);
nor U12865 (N_12865,N_11542,N_8951);
nand U12866 (N_12866,N_11964,N_11414);
nor U12867 (N_12867,N_9672,N_10938);
nor U12868 (N_12868,N_10234,N_10730);
xnor U12869 (N_12869,N_10998,N_9049);
or U12870 (N_12870,N_9417,N_8790);
or U12871 (N_12871,N_8234,N_10684);
and U12872 (N_12872,N_8156,N_10977);
or U12873 (N_12873,N_10020,N_11333);
or U12874 (N_12874,N_9399,N_9109);
xnor U12875 (N_12875,N_9199,N_9579);
and U12876 (N_12876,N_9411,N_10238);
xnor U12877 (N_12877,N_9762,N_9572);
and U12878 (N_12878,N_8619,N_8038);
nand U12879 (N_12879,N_10834,N_11804);
nor U12880 (N_12880,N_11342,N_9258);
nor U12881 (N_12881,N_9382,N_9847);
and U12882 (N_12882,N_11392,N_8764);
nand U12883 (N_12883,N_8251,N_10144);
xor U12884 (N_12884,N_11793,N_9427);
and U12885 (N_12885,N_10527,N_9829);
xnor U12886 (N_12886,N_8261,N_11512);
nor U12887 (N_12887,N_8400,N_11328);
and U12888 (N_12888,N_8262,N_11953);
xnor U12889 (N_12889,N_9664,N_11268);
and U12890 (N_12890,N_8941,N_11270);
or U12891 (N_12891,N_9587,N_8125);
nor U12892 (N_12892,N_10051,N_9801);
xor U12893 (N_12893,N_10290,N_10845);
nor U12894 (N_12894,N_8422,N_9675);
nor U12895 (N_12895,N_8435,N_10685);
nand U12896 (N_12896,N_8509,N_8762);
nor U12897 (N_12897,N_11499,N_10783);
nor U12898 (N_12898,N_9824,N_11386);
or U12899 (N_12899,N_9165,N_11263);
or U12900 (N_12900,N_10787,N_10146);
nor U12901 (N_12901,N_10933,N_9120);
or U12902 (N_12902,N_10677,N_10551);
or U12903 (N_12903,N_11254,N_10324);
nor U12904 (N_12904,N_9549,N_8086);
and U12905 (N_12905,N_11738,N_9387);
nand U12906 (N_12906,N_8389,N_10221);
xnor U12907 (N_12907,N_9720,N_10396);
xnor U12908 (N_12908,N_10863,N_9058);
and U12909 (N_12909,N_11252,N_10747);
nor U12910 (N_12910,N_10665,N_9141);
xnor U12911 (N_12911,N_9053,N_8067);
and U12912 (N_12912,N_9941,N_11248);
and U12913 (N_12913,N_10364,N_11523);
and U12914 (N_12914,N_10235,N_11219);
xnor U12915 (N_12915,N_11361,N_8589);
or U12916 (N_12916,N_8735,N_10729);
and U12917 (N_12917,N_8416,N_9643);
xor U12918 (N_12918,N_10995,N_11223);
nor U12919 (N_12919,N_9396,N_10991);
nor U12920 (N_12920,N_9335,N_8924);
or U12921 (N_12921,N_10993,N_10268);
and U12922 (N_12922,N_10225,N_9933);
or U12923 (N_12923,N_10222,N_8750);
and U12924 (N_12924,N_8797,N_10987);
or U12925 (N_12925,N_10462,N_9600);
nor U12926 (N_12926,N_9641,N_11824);
nor U12927 (N_12927,N_10587,N_8272);
nand U12928 (N_12928,N_8264,N_11491);
nor U12929 (N_12929,N_11901,N_9322);
and U12930 (N_12930,N_9753,N_11378);
nand U12931 (N_12931,N_10554,N_10989);
or U12932 (N_12932,N_11148,N_10691);
and U12933 (N_12933,N_10887,N_10614);
nand U12934 (N_12934,N_10626,N_8345);
and U12935 (N_12935,N_8522,N_11052);
and U12936 (N_12936,N_10183,N_8819);
and U12937 (N_12937,N_8167,N_8908);
nand U12938 (N_12938,N_8405,N_9917);
and U12939 (N_12939,N_10818,N_8886);
nor U12940 (N_12940,N_11620,N_10801);
nand U12941 (N_12941,N_11218,N_10447);
nand U12942 (N_12942,N_9708,N_9907);
and U12943 (N_12943,N_10048,N_11614);
xor U12944 (N_12944,N_8378,N_9886);
nand U12945 (N_12945,N_11266,N_10948);
xnor U12946 (N_12946,N_11750,N_9264);
or U12947 (N_12947,N_10263,N_8659);
and U12948 (N_12948,N_8118,N_10073);
nand U12949 (N_12949,N_8622,N_9649);
or U12950 (N_12950,N_8201,N_11554);
or U12951 (N_12951,N_10855,N_11996);
nand U12952 (N_12952,N_10611,N_9855);
and U12953 (N_12953,N_10702,N_9901);
or U12954 (N_12954,N_10809,N_9454);
or U12955 (N_12955,N_9563,N_10500);
and U12956 (N_12956,N_11190,N_10630);
or U12957 (N_12957,N_9421,N_9777);
or U12958 (N_12958,N_10269,N_9577);
and U12959 (N_12959,N_11211,N_11461);
or U12960 (N_12960,N_8690,N_9521);
nand U12961 (N_12961,N_10247,N_10641);
xor U12962 (N_12962,N_10140,N_9276);
nor U12963 (N_12963,N_8135,N_8965);
and U12964 (N_12964,N_9657,N_11246);
and U12965 (N_12965,N_8821,N_10549);
nand U12966 (N_12966,N_9415,N_8255);
nand U12967 (N_12967,N_11385,N_8882);
and U12968 (N_12968,N_11486,N_8260);
and U12969 (N_12969,N_8623,N_11608);
and U12970 (N_12970,N_10013,N_9469);
or U12971 (N_12971,N_10650,N_10763);
nand U12972 (N_12972,N_9432,N_8572);
or U12973 (N_12973,N_10016,N_9618);
nor U12974 (N_12974,N_10767,N_11653);
xnor U12975 (N_12975,N_10990,N_9076);
xnor U12976 (N_12976,N_9224,N_8434);
nand U12977 (N_12977,N_8806,N_10828);
and U12978 (N_12978,N_9169,N_11415);
or U12979 (N_12979,N_9850,N_10829);
and U12980 (N_12980,N_9807,N_8720);
or U12981 (N_12981,N_10696,N_11945);
xnor U12982 (N_12982,N_9526,N_9888);
nor U12983 (N_12983,N_8128,N_10473);
or U12984 (N_12984,N_9590,N_10072);
nand U12985 (N_12985,N_8289,N_10295);
and U12986 (N_12986,N_8396,N_11068);
or U12987 (N_12987,N_10070,N_8570);
and U12988 (N_12988,N_11114,N_10102);
nand U12989 (N_12989,N_9311,N_8250);
or U12990 (N_12990,N_11994,N_10586);
and U12991 (N_12991,N_9317,N_8353);
nand U12992 (N_12992,N_9161,N_10267);
and U12993 (N_12993,N_8288,N_11657);
xor U12994 (N_12994,N_10986,N_9026);
nand U12995 (N_12995,N_11498,N_11410);
nand U12996 (N_12996,N_11648,N_10377);
nand U12997 (N_12997,N_10795,N_10210);
and U12998 (N_12998,N_11024,N_10032);
nor U12999 (N_12999,N_9107,N_11448);
or U13000 (N_13000,N_11877,N_11852);
or U13001 (N_13001,N_9875,N_11277);
nor U13002 (N_13002,N_9697,N_9323);
and U13003 (N_13003,N_10861,N_8968);
or U13004 (N_13004,N_8817,N_8013);
and U13005 (N_13005,N_10658,N_9406);
or U13006 (N_13006,N_10723,N_10594);
nor U13007 (N_13007,N_10911,N_10923);
and U13008 (N_13008,N_9574,N_9893);
nor U13009 (N_13009,N_11493,N_9181);
nand U13010 (N_13010,N_8680,N_8992);
or U13011 (N_13011,N_9342,N_8624);
and U13012 (N_13012,N_8014,N_9756);
and U13013 (N_13013,N_8041,N_10846);
nor U13014 (N_13014,N_9333,N_9087);
and U13015 (N_13015,N_10585,N_8970);
or U13016 (N_13016,N_11775,N_11354);
nand U13017 (N_13017,N_10033,N_10759);
and U13018 (N_13018,N_9934,N_9357);
or U13019 (N_13019,N_8775,N_11495);
or U13020 (N_13020,N_10757,N_11018);
or U13021 (N_13021,N_10935,N_11175);
and U13022 (N_13022,N_9898,N_11279);
nand U13023 (N_13023,N_8744,N_10340);
nand U13024 (N_13024,N_8944,N_11158);
nor U13025 (N_13025,N_10962,N_11703);
nor U13026 (N_13026,N_8460,N_10874);
or U13027 (N_13027,N_10372,N_9271);
and U13028 (N_13028,N_8098,N_9202);
nor U13029 (N_13029,N_11979,N_8146);
or U13030 (N_13030,N_8765,N_8249);
nand U13031 (N_13031,N_8340,N_9504);
or U13032 (N_13032,N_8342,N_8833);
and U13033 (N_13033,N_11583,N_10291);
nor U13034 (N_13034,N_10825,N_9834);
xor U13035 (N_13035,N_10741,N_9464);
or U13036 (N_13036,N_9245,N_11977);
nand U13037 (N_13037,N_9184,N_10107);
nor U13038 (N_13038,N_9564,N_10439);
nor U13039 (N_13039,N_11072,N_8317);
and U13040 (N_13040,N_11122,N_10442);
nor U13041 (N_13041,N_8051,N_10601);
nor U13042 (N_13042,N_9488,N_9212);
nand U13043 (N_13043,N_10728,N_8028);
or U13044 (N_13044,N_10337,N_9880);
and U13045 (N_13045,N_10974,N_8988);
nand U13046 (N_13046,N_9022,N_10789);
or U13047 (N_13047,N_9781,N_9811);
nand U13048 (N_13048,N_11364,N_9404);
or U13049 (N_13049,N_8139,N_10864);
and U13050 (N_13050,N_9183,N_11686);
and U13051 (N_13051,N_10371,N_9620);
and U13052 (N_13052,N_8140,N_8578);
or U13053 (N_13053,N_9845,N_8916);
xnor U13054 (N_13054,N_11943,N_9827);
xnor U13055 (N_13055,N_8670,N_9017);
or U13056 (N_13056,N_9455,N_8844);
or U13057 (N_13057,N_9595,N_11761);
or U13058 (N_13058,N_11075,N_9484);
or U13059 (N_13059,N_8798,N_11436);
or U13060 (N_13060,N_9543,N_8593);
or U13061 (N_13061,N_9303,N_9881);
and U13062 (N_13062,N_9717,N_8376);
and U13063 (N_13063,N_11487,N_10997);
and U13064 (N_13064,N_10751,N_10285);
and U13065 (N_13065,N_11280,N_10464);
and U13066 (N_13066,N_9334,N_11186);
and U13067 (N_13067,N_11768,N_11049);
nand U13068 (N_13068,N_9220,N_9292);
nor U13069 (N_13069,N_11565,N_8224);
and U13070 (N_13070,N_10004,N_9923);
and U13071 (N_13071,N_10388,N_9896);
nand U13072 (N_13072,N_10103,N_10836);
xnor U13073 (N_13073,N_9422,N_8963);
xor U13074 (N_13074,N_8826,N_8179);
nand U13075 (N_13075,N_8630,N_11225);
or U13076 (N_13076,N_8692,N_8781);
and U13077 (N_13077,N_10617,N_8305);
and U13078 (N_13078,N_10370,N_10499);
or U13079 (N_13079,N_8559,N_9345);
nand U13080 (N_13080,N_9363,N_10108);
and U13081 (N_13081,N_9640,N_10556);
xor U13082 (N_13082,N_10109,N_10854);
nand U13083 (N_13083,N_10069,N_11908);
nor U13084 (N_13084,N_9755,N_10984);
nand U13085 (N_13085,N_9483,N_10797);
nor U13086 (N_13086,N_9226,N_11064);
and U13087 (N_13087,N_9559,N_8117);
nand U13088 (N_13088,N_11939,N_9605);
nand U13089 (N_13089,N_9050,N_10055);
and U13090 (N_13090,N_9376,N_8457);
nor U13091 (N_13091,N_11545,N_9744);
nor U13092 (N_13092,N_11756,N_11551);
xnor U13093 (N_13093,N_10813,N_9693);
nand U13094 (N_13094,N_11622,N_9538);
nor U13095 (N_13095,N_9910,N_9622);
xnor U13096 (N_13096,N_11553,N_9277);
or U13097 (N_13097,N_8256,N_8006);
nand U13098 (N_13098,N_10352,N_10632);
xnor U13099 (N_13099,N_8814,N_8686);
and U13100 (N_13100,N_10058,N_11109);
or U13101 (N_13101,N_9059,N_9208);
nor U13102 (N_13102,N_8148,N_9677);
nor U13103 (N_13103,N_8554,N_10311);
and U13104 (N_13104,N_9150,N_11932);
nor U13105 (N_13105,N_11741,N_9431);
nand U13106 (N_13106,N_10883,N_11424);
or U13107 (N_13107,N_8510,N_8290);
and U13108 (N_13108,N_11941,N_8749);
nor U13109 (N_13109,N_8654,N_11031);
nor U13110 (N_13110,N_8727,N_10704);
nor U13111 (N_13111,N_8642,N_9952);
nor U13112 (N_13112,N_10520,N_9591);
nor U13113 (N_13113,N_10727,N_9686);
nor U13114 (N_13114,N_8144,N_10667);
nor U13115 (N_13115,N_10964,N_11666);
nor U13116 (N_13116,N_10976,N_10628);
nand U13117 (N_13117,N_10937,N_9255);
nand U13118 (N_13118,N_8779,N_10133);
nor U13119 (N_13119,N_8527,N_8689);
xor U13120 (N_13120,N_11917,N_8596);
nor U13121 (N_13121,N_8948,N_11812);
or U13122 (N_13122,N_10635,N_9919);
nand U13123 (N_13123,N_11239,N_10484);
and U13124 (N_13124,N_8491,N_10094);
nor U13125 (N_13125,N_9658,N_11231);
nor U13126 (N_13126,N_8895,N_11187);
and U13127 (N_13127,N_11865,N_8069);
nand U13128 (N_13128,N_9079,N_8394);
nand U13129 (N_13129,N_11056,N_9486);
nand U13130 (N_13130,N_11705,N_11742);
or U13131 (N_13131,N_8915,N_9461);
nor U13132 (N_13132,N_11008,N_9287);
and U13133 (N_13133,N_10175,N_8945);
nor U13134 (N_13134,N_11099,N_9684);
nor U13135 (N_13135,N_8756,N_8892);
nand U13136 (N_13136,N_11843,N_10343);
and U13137 (N_13137,N_10627,N_9909);
nor U13138 (N_13138,N_10173,N_8746);
or U13139 (N_13139,N_9891,N_8035);
and U13140 (N_13140,N_11844,N_9669);
or U13141 (N_13141,N_11201,N_11727);
or U13142 (N_13142,N_10206,N_10157);
nor U13143 (N_13143,N_10985,N_8845);
and U13144 (N_13144,N_11272,N_9262);
nor U13145 (N_13145,N_8055,N_9883);
or U13146 (N_13146,N_9320,N_11479);
nor U13147 (N_13147,N_8408,N_10168);
nor U13148 (N_13148,N_10674,N_8954);
or U13149 (N_13149,N_9307,N_8359);
xor U13150 (N_13150,N_11285,N_9539);
or U13151 (N_13151,N_9712,N_8088);
or U13152 (N_13152,N_8556,N_10535);
nand U13153 (N_13153,N_11264,N_11647);
nand U13154 (N_13154,N_9868,N_8683);
nand U13155 (N_13155,N_9193,N_11330);
nor U13156 (N_13156,N_8799,N_8020);
nand U13157 (N_13157,N_11773,N_11067);
or U13158 (N_13158,N_10395,N_9866);
nand U13159 (N_13159,N_10803,N_10277);
or U13160 (N_13160,N_11893,N_11496);
nand U13161 (N_13161,N_10725,N_11405);
nor U13162 (N_13162,N_8303,N_8141);
or U13163 (N_13163,N_9312,N_9324);
nand U13164 (N_13164,N_8245,N_8678);
nand U13165 (N_13165,N_10833,N_8452);
or U13166 (N_13166,N_9299,N_10087);
and U13167 (N_13167,N_11289,N_10670);
or U13168 (N_13168,N_10915,N_8569);
xnor U13169 (N_13169,N_9232,N_9706);
and U13170 (N_13170,N_9785,N_10629);
nand U13171 (N_13171,N_8921,N_9982);
nor U13172 (N_13172,N_8197,N_10092);
and U13173 (N_13173,N_10355,N_9164);
and U13174 (N_13174,N_9413,N_9843);
nor U13175 (N_13175,N_11639,N_8200);
nor U13176 (N_13176,N_8584,N_8856);
nor U13177 (N_13177,N_11108,N_8415);
xnor U13178 (N_13178,N_9001,N_10676);
nand U13179 (N_13179,N_9648,N_11076);
or U13180 (N_13180,N_11467,N_11391);
and U13181 (N_13181,N_8880,N_10274);
and U13182 (N_13182,N_11472,N_8180);
nor U13183 (N_13183,N_9949,N_11250);
nor U13184 (N_13184,N_11450,N_8713);
and U13185 (N_13185,N_11786,N_11716);
and U13186 (N_13186,N_10067,N_10740);
nand U13187 (N_13187,N_9989,N_11506);
and U13188 (N_13188,N_11338,N_8610);
or U13189 (N_13189,N_8377,N_9154);
or U13190 (N_13190,N_10093,N_8891);
nand U13191 (N_13191,N_9228,N_8461);
and U13192 (N_13192,N_10063,N_9890);
nor U13193 (N_13193,N_11504,N_8445);
nor U13194 (N_13194,N_11485,N_9441);
and U13195 (N_13195,N_8333,N_11131);
or U13196 (N_13196,N_8459,N_10403);
and U13197 (N_13197,N_10901,N_11912);
nand U13198 (N_13198,N_9004,N_8343);
nor U13199 (N_13199,N_8203,N_10672);
nand U13200 (N_13200,N_11406,N_9476);
or U13201 (N_13201,N_11550,N_9051);
nand U13202 (N_13202,N_9822,N_8134);
nor U13203 (N_13203,N_9002,N_11006);
xor U13204 (N_13204,N_8633,N_8282);
xnor U13205 (N_13205,N_11073,N_8244);
or U13206 (N_13206,N_10205,N_8136);
nor U13207 (N_13207,N_9175,N_11973);
nor U13208 (N_13208,N_10472,N_8573);
and U13209 (N_13209,N_10153,N_10649);
or U13210 (N_13210,N_8095,N_9953);
nand U13211 (N_13211,N_8332,N_8818);
nor U13212 (N_13212,N_9537,N_11320);
nand U13213 (N_13213,N_11455,N_9440);
or U13214 (N_13214,N_8676,N_11228);
xnor U13215 (N_13215,N_11478,N_10903);
or U13216 (N_13216,N_9984,N_8477);
nand U13217 (N_13217,N_9240,N_11105);
or U13218 (N_13218,N_10209,N_10202);
nand U13219 (N_13219,N_9581,N_8033);
nand U13220 (N_13220,N_8729,N_9209);
and U13221 (N_13221,N_10859,N_9463);
nand U13222 (N_13222,N_9344,N_9057);
and U13223 (N_13223,N_8286,N_9361);
or U13224 (N_13224,N_10119,N_11999);
or U13225 (N_13225,N_11799,N_10583);
and U13226 (N_13226,N_9838,N_9337);
nor U13227 (N_13227,N_11247,N_10219);
nand U13228 (N_13228,N_11390,N_8409);
or U13229 (N_13229,N_9095,N_11082);
or U13230 (N_13230,N_8058,N_8021);
nor U13231 (N_13231,N_11128,N_11998);
or U13232 (N_13232,N_11007,N_9900);
and U13233 (N_13233,N_9309,N_8449);
nand U13234 (N_13234,N_9751,N_8800);
or U13235 (N_13235,N_10275,N_10746);
nand U13236 (N_13236,N_10748,N_11717);
and U13237 (N_13237,N_10815,N_8687);
nor U13238 (N_13238,N_9040,N_9072);
and U13239 (N_13239,N_8257,N_10451);
and U13240 (N_13240,N_11325,N_9844);
or U13241 (N_13241,N_9284,N_9921);
nor U13242 (N_13242,N_8383,N_8949);
and U13243 (N_13243,N_11294,N_11579);
nor U13244 (N_13244,N_10257,N_10030);
nand U13245 (N_13245,N_9635,N_11177);
or U13246 (N_13246,N_10678,N_9867);
or U13247 (N_13247,N_9647,N_9143);
and U13248 (N_13248,N_8147,N_11592);
and U13249 (N_13249,N_9631,N_8538);
nand U13250 (N_13250,N_8521,N_11992);
or U13251 (N_13251,N_8517,N_10562);
or U13252 (N_13252,N_11511,N_9644);
nand U13253 (N_13253,N_9025,N_8699);
xor U13254 (N_13254,N_10597,N_9471);
nor U13255 (N_13255,N_9812,N_11989);
nor U13256 (N_13256,N_8064,N_8344);
and U13257 (N_13257,N_8704,N_11042);
xor U13258 (N_13258,N_11369,N_10734);
nand U13259 (N_13259,N_8533,N_9828);
nand U13260 (N_13260,N_9198,N_11724);
or U13261 (N_13261,N_9503,N_9039);
and U13262 (N_13262,N_8905,N_10182);
and U13263 (N_13263,N_11683,N_9327);
and U13264 (N_13264,N_8293,N_10122);
nand U13265 (N_13265,N_8002,N_10155);
nor U13266 (N_13266,N_10327,N_9879);
or U13267 (N_13267,N_9651,N_9628);
nor U13268 (N_13268,N_10424,N_10112);
and U13269 (N_13269,N_9930,N_9279);
nor U13270 (N_13270,N_8212,N_9765);
and U13271 (N_13271,N_8714,N_11290);
or U13272 (N_13272,N_9041,N_11790);
or U13273 (N_13273,N_10524,N_8281);
nor U13274 (N_13274,N_10523,N_9270);
and U13275 (N_13275,N_11714,N_8561);
nand U13276 (N_13276,N_10893,N_11881);
and U13277 (N_13277,N_9749,N_9129);
nand U13278 (N_13278,N_11969,N_8057);
or U13279 (N_13279,N_10459,N_10762);
nand U13280 (N_13280,N_9006,N_11871);
xnor U13281 (N_13281,N_11251,N_8576);
and U13282 (N_13282,N_8018,N_11300);
or U13283 (N_13283,N_9571,N_11976);
and U13284 (N_13284,N_9610,N_11850);
nor U13285 (N_13285,N_11150,N_9444);
or U13286 (N_13286,N_9219,N_9903);
and U13287 (N_13287,N_11446,N_10349);
or U13288 (N_13288,N_11859,N_8216);
nand U13289 (N_13289,N_10025,N_10944);
or U13290 (N_13290,N_11519,N_9586);
xor U13291 (N_13291,N_9373,N_10517);
nand U13292 (N_13292,N_11170,N_9705);
nand U13293 (N_13293,N_8730,N_10965);
nor U13294 (N_13294,N_10098,N_10735);
and U13295 (N_13295,N_8169,N_11151);
xor U13296 (N_13296,N_9250,N_11407);
and U13297 (N_13297,N_9200,N_10776);
nand U13298 (N_13298,N_11735,N_8937);
or U13299 (N_13299,N_9553,N_11267);
nand U13300 (N_13300,N_9841,N_9119);
and U13301 (N_13301,N_10777,N_8825);
nand U13302 (N_13302,N_10314,N_10313);
nand U13303 (N_13303,N_8553,N_10333);
nand U13304 (N_13304,N_10505,N_11382);
or U13305 (N_13305,N_11764,N_11437);
or U13306 (N_13306,N_10603,N_8813);
nand U13307 (N_13307,N_11332,N_8008);
or U13308 (N_13308,N_10045,N_8736);
nor U13309 (N_13309,N_10590,N_8793);
nand U13310 (N_13310,N_8129,N_11278);
nor U13311 (N_13311,N_10036,N_10778);
nor U13312 (N_13312,N_11366,N_11700);
or U13313 (N_13313,N_11902,N_9229);
nand U13314 (N_13314,N_10570,N_10165);
nor U13315 (N_13315,N_9518,N_11890);
or U13316 (N_13316,N_8225,N_9156);
xor U13317 (N_13317,N_9425,N_11403);
and U13318 (N_13318,N_8102,N_11389);
and U13319 (N_13319,N_9084,N_10231);
or U13320 (N_13320,N_11923,N_9467);
xor U13321 (N_13321,N_9703,N_8639);
nand U13322 (N_13322,N_8674,N_11582);
or U13323 (N_13323,N_10161,N_8468);
nor U13324 (N_13324,N_11584,N_8651);
nand U13325 (N_13325,N_10420,N_9609);
nor U13326 (N_13326,N_9725,N_8354);
nand U13327 (N_13327,N_9852,N_9481);
and U13328 (N_13328,N_11933,N_8621);
nand U13329 (N_13329,N_8001,N_9251);
nand U13330 (N_13330,N_9056,N_9819);
xor U13331 (N_13331,N_10483,N_11014);
nand U13332 (N_13332,N_9767,N_8601);
and U13333 (N_13333,N_8370,N_9448);
xor U13334 (N_13334,N_9348,N_9981);
and U13335 (N_13335,N_11872,N_11261);
and U13336 (N_13336,N_8175,N_10281);
nand U13337 (N_13337,N_10037,N_11626);
xnor U13338 (N_13338,N_8741,N_11110);
nor U13339 (N_13339,N_11905,N_11471);
or U13340 (N_13340,N_11887,N_9442);
and U13341 (N_13341,N_9151,N_8323);
and U13342 (N_13342,N_9833,N_10561);
and U13343 (N_13343,N_9213,N_8052);
xnor U13344 (N_13344,N_9171,N_8869);
nor U13345 (N_13345,N_9623,N_8007);
nand U13346 (N_13346,N_9552,N_9090);
nor U13347 (N_13347,N_8073,N_9761);
xnor U13348 (N_13348,N_9349,N_10745);
xnor U13349 (N_13349,N_10114,N_10478);
nand U13350 (N_13350,N_11528,N_10577);
or U13351 (N_13351,N_10185,N_11301);
nor U13352 (N_13352,N_11011,N_9499);
or U13353 (N_13353,N_11578,N_11435);
nor U13354 (N_13354,N_9023,N_11234);
or U13355 (N_13355,N_9369,N_8884);
nand U13356 (N_13356,N_9241,N_8675);
or U13357 (N_13357,N_11112,N_9607);
nor U13358 (N_13358,N_8142,N_10733);
or U13359 (N_13359,N_9071,N_11548);
xnor U13360 (N_13360,N_9293,N_9561);
nand U13361 (N_13361,N_9555,N_10428);
or U13362 (N_13362,N_9873,N_11573);
nand U13363 (N_13363,N_11080,N_11383);
xnor U13364 (N_13364,N_11642,N_10713);
nand U13365 (N_13365,N_10046,N_11217);
nand U13366 (N_13366,N_11805,N_11883);
xnor U13367 (N_13367,N_9960,N_10479);
xor U13368 (N_13368,N_11265,N_9687);
nor U13369 (N_13369,N_10506,N_8657);
or U13370 (N_13370,N_9392,N_11173);
and U13371 (N_13371,N_8163,N_9589);
nor U13372 (N_13372,N_8121,N_10201);
nand U13373 (N_13373,N_8091,N_9916);
or U13374 (N_13374,N_10325,N_9350);
and U13375 (N_13375,N_9815,N_9882);
nor U13376 (N_13376,N_11785,N_8145);
nand U13377 (N_13377,N_9048,N_10652);
and U13378 (N_13378,N_11529,N_10814);
or U13379 (N_13379,N_10393,N_9294);
or U13380 (N_13380,N_11107,N_11556);
nand U13381 (N_13381,N_10354,N_10761);
and U13382 (N_13382,N_10595,N_11387);
nor U13383 (N_13383,N_11574,N_11138);
nor U13384 (N_13384,N_8109,N_8085);
and U13385 (N_13385,N_10163,N_9383);
and U13386 (N_13386,N_9125,N_11154);
nand U13387 (N_13387,N_9083,N_11071);
or U13388 (N_13388,N_8904,N_8373);
and U13389 (N_13389,N_8861,N_8504);
and U13390 (N_13390,N_8866,N_10786);
and U13391 (N_13391,N_8760,N_10576);
nor U13392 (N_13392,N_8723,N_10432);
nor U13393 (N_13393,N_8566,N_9409);
and U13394 (N_13394,N_9474,N_11737);
or U13395 (N_13395,N_8235,N_11417);
or U13396 (N_13396,N_11779,N_8999);
nor U13397 (N_13397,N_9698,N_8194);
nand U13398 (N_13398,N_11305,N_9286);
nand U13399 (N_13399,N_10545,N_10760);
nor U13400 (N_13400,N_9060,N_8287);
and U13401 (N_13401,N_11022,N_10376);
xnor U13402 (N_13402,N_11205,N_10450);
nor U13403 (N_13403,N_9959,N_11541);
nand U13404 (N_13404,N_8280,N_10147);
or U13405 (N_13405,N_10305,N_10351);
nor U13406 (N_13406,N_10895,N_10421);
nand U13407 (N_13407,N_9094,N_11643);
nor U13408 (N_13408,N_11337,N_11825);
xnor U13409 (N_13409,N_11987,N_9598);
nor U13410 (N_13410,N_8598,N_10661);
xnor U13411 (N_13411,N_11800,N_9741);
and U13412 (N_13412,N_10411,N_9985);
or U13413 (N_13413,N_11213,N_8820);
nand U13414 (N_13414,N_9424,N_9804);
and U13415 (N_13415,N_8111,N_8492);
and U13416 (N_13416,N_9743,N_11536);
nand U13417 (N_13417,N_11393,N_11633);
nor U13418 (N_13418,N_10339,N_9205);
and U13419 (N_13419,N_9924,N_10178);
nand U13420 (N_13420,N_11640,N_8748);
and U13421 (N_13421,N_10879,N_9118);
and U13422 (N_13422,N_10612,N_9460);
nor U13423 (N_13423,N_8558,N_8433);
nor U13424 (N_13424,N_10429,N_11618);
and U13425 (N_13425,N_11659,N_11809);
nand U13426 (N_13426,N_9823,N_10382);
and U13427 (N_13427,N_9808,N_9033);
and U13428 (N_13428,N_10309,N_11442);
nand U13429 (N_13429,N_9679,N_11046);
nand U13430 (N_13430,N_10150,N_8520);
nor U13431 (N_13431,N_10366,N_10124);
or U13432 (N_13432,N_11751,N_11309);
nand U13433 (N_13433,N_8783,N_8213);
nor U13434 (N_13434,N_10368,N_8590);
nor U13435 (N_13435,N_8050,N_9652);
nand U13436 (N_13436,N_9069,N_8980);
nand U13437 (N_13437,N_8087,N_11286);
nand U13438 (N_13438,N_11188,N_11886);
or U13439 (N_13439,N_9961,N_9500);
nor U13440 (N_13440,N_9430,N_10509);
or U13441 (N_13441,N_11713,N_9929);
and U13442 (N_13442,N_9197,N_8583);
and U13443 (N_13443,N_9238,N_8404);
xor U13444 (N_13444,N_9818,N_9770);
nor U13445 (N_13445,N_8054,N_9938);
or U13446 (N_13446,N_11402,N_9370);
or U13447 (N_13447,N_9976,N_8437);
nand U13448 (N_13448,N_11408,N_11841);
nand U13449 (N_13449,N_8849,N_11374);
or U13450 (N_13450,N_10292,N_10960);
and U13451 (N_13451,N_11505,N_9256);
nand U13452 (N_13452,N_11828,N_11728);
and U13453 (N_13453,N_9147,N_11001);
or U13454 (N_13454,N_8933,N_8715);
or U13455 (N_13455,N_8152,N_10705);
and U13456 (N_13456,N_9400,N_9239);
and U13457 (N_13457,N_9826,N_10123);
or U13458 (N_13458,N_8229,N_11563);
nor U13459 (N_13459,N_9230,N_9328);
and U13460 (N_13460,N_9851,N_8268);
nor U13461 (N_13461,N_10436,N_8047);
or U13462 (N_13462,N_9168,N_11139);
nor U13463 (N_13463,N_10868,N_8172);
and U13464 (N_13464,N_10017,N_10284);
nand U13465 (N_13465,N_10644,N_11911);
or U13466 (N_13466,N_10502,N_9085);
nor U13467 (N_13467,N_11240,N_10394);
nor U13468 (N_13468,N_9950,N_9513);
and U13469 (N_13469,N_9895,N_8943);
and U13470 (N_13470,N_8865,N_10076);
or U13471 (N_13471,N_10572,N_11909);
and U13472 (N_13472,N_10653,N_11236);
xnor U13473 (N_13473,N_10764,N_10752);
nand U13474 (N_13474,N_11016,N_11950);
nor U13475 (N_13475,N_9633,N_11079);
and U13476 (N_13476,N_9010,N_8455);
nor U13477 (N_13477,N_9042,N_10955);
or U13478 (N_13478,N_11624,N_9864);
or U13479 (N_13479,N_11421,N_11502);
or U13480 (N_13480,N_8536,N_10348);
xor U13481 (N_13481,N_8931,N_8516);
and U13482 (N_13482,N_11113,N_8860);
nor U13483 (N_13483,N_8252,N_10271);
nor U13484 (N_13484,N_9554,N_8495);
xnor U13485 (N_13485,N_11581,N_10270);
nand U13486 (N_13486,N_9626,N_9446);
nor U13487 (N_13487,N_11849,N_8549);
nand U13488 (N_13488,N_9511,N_8957);
nor U13489 (N_13489,N_8489,N_10662);
or U13490 (N_13490,N_9940,N_8414);
and U13491 (N_13491,N_9259,N_9265);
nor U13492 (N_13492,N_8627,N_9972);
or U13493 (N_13493,N_11449,N_11166);
and U13494 (N_13494,N_10398,N_10980);
or U13495 (N_13495,N_11070,N_8546);
or U13496 (N_13496,N_11612,N_11619);
or U13497 (N_13497,N_10552,N_10939);
and U13498 (N_13498,N_10077,N_11101);
and U13499 (N_13499,N_8645,N_9000);
or U13500 (N_13500,N_9637,N_9796);
or U13501 (N_13501,N_8550,N_11821);
or U13502 (N_13502,N_10226,N_10088);
or U13503 (N_13503,N_9372,N_10027);
or U13504 (N_13504,N_10692,N_11103);
or U13505 (N_13505,N_8898,N_8801);
nand U13506 (N_13506,N_8707,N_11133);
nor U13507 (N_13507,N_11597,N_11198);
nand U13508 (N_13508,N_9045,N_11668);
xor U13509 (N_13509,N_11876,N_9653);
xor U13510 (N_13510,N_8673,N_11243);
nor U13511 (N_13511,N_9676,N_8586);
xnor U13512 (N_13512,N_9560,N_11306);
or U13513 (N_13513,N_8472,N_9836);
nor U13514 (N_13514,N_9225,N_10707);
nand U13515 (N_13515,N_10038,N_10041);
and U13516 (N_13516,N_8382,N_8138);
and U13517 (N_13517,N_9416,N_11399);
or U13518 (N_13518,N_10681,N_10261);
or U13519 (N_13519,N_8391,N_10934);
and U13520 (N_13520,N_10047,N_10726);
or U13521 (N_13521,N_11059,N_9998);
xor U13522 (N_13522,N_10636,N_8080);
nor U13523 (N_13523,N_9735,N_11811);
or U13524 (N_13524,N_10213,N_11141);
or U13525 (N_13525,N_9089,N_8254);
nand U13526 (N_13526,N_8024,N_10300);
nor U13527 (N_13527,N_11834,N_8439);
nor U13528 (N_13528,N_11084,N_11060);
nand U13529 (N_13529,N_10043,N_11453);
nor U13530 (N_13530,N_9520,N_9036);
nand U13531 (N_13531,N_8733,N_10771);
nor U13532 (N_13532,N_9528,N_9126);
or U13533 (N_13533,N_10117,N_8061);
and U13534 (N_13534,N_10232,N_10679);
or U13535 (N_13535,N_9681,N_11470);
nand U13536 (N_13536,N_8322,N_10555);
nand U13537 (N_13537,N_8498,N_10992);
and U13538 (N_13538,N_10531,N_11034);
nand U13539 (N_13539,N_11621,N_11972);
or U13540 (N_13540,N_10075,N_11466);
and U13541 (N_13541,N_9130,N_10507);
and U13542 (N_13542,N_8850,N_9558);
or U13543 (N_13543,N_10128,N_8056);
and U13544 (N_13544,N_10362,N_9750);
nand U13545 (N_13545,N_11801,N_8043);
and U13546 (N_13546,N_10659,N_8227);
nor U13547 (N_13547,N_10402,N_8237);
nor U13548 (N_13548,N_8679,N_9860);
nand U13549 (N_13549,N_11318,N_8060);
and U13550 (N_13550,N_10141,N_8541);
xnor U13551 (N_13551,N_9252,N_8696);
or U13552 (N_13552,N_9737,N_9206);
or U13553 (N_13553,N_11914,N_8178);
xnor U13554 (N_13554,N_8000,N_9174);
nor U13555 (N_13555,N_9569,N_10823);
nand U13556 (N_13556,N_11763,N_11229);
or U13557 (N_13557,N_10519,N_10501);
and U13558 (N_13558,N_11853,N_11104);
and U13559 (N_13559,N_9871,N_10715);
nor U13560 (N_13560,N_11892,N_9316);
and U13561 (N_13561,N_11854,N_9178);
nor U13562 (N_13562,N_10207,N_8059);
nor U13563 (N_13563,N_10891,N_10827);
nor U13564 (N_13564,N_10732,N_11985);
xor U13565 (N_13565,N_9769,N_11591);
or U13566 (N_13566,N_9654,N_10296);
nor U13567 (N_13567,N_9043,N_11476);
and U13568 (N_13568,N_8294,N_11375);
and U13569 (N_13569,N_11599,N_9267);
nor U13570 (N_13570,N_9690,N_8297);
nand U13571 (N_13571,N_10796,N_8160);
and U13572 (N_13572,N_8893,N_11083);
or U13573 (N_13573,N_9122,N_8259);
and U13574 (N_13574,N_11288,N_9937);
nor U13575 (N_13575,N_10229,N_11362);
nor U13576 (N_13576,N_8677,N_8372);
and U13577 (N_13577,N_8662,N_11167);
nand U13578 (N_13578,N_10546,N_9114);
nand U13579 (N_13579,N_9266,N_11503);
or U13580 (N_13580,N_10851,N_9364);
or U13581 (N_13581,N_9709,N_9507);
nor U13582 (N_13582,N_8412,N_11055);
and U13583 (N_13583,N_9636,N_9037);
nor U13584 (N_13584,N_10466,N_10214);
xor U13585 (N_13585,N_11679,N_11918);
xnor U13586 (N_13586,N_10052,N_11291);
and U13587 (N_13587,N_10940,N_9532);
or U13588 (N_13588,N_11667,N_10878);
and U13589 (N_13589,N_8761,N_11540);
xnor U13590 (N_13590,N_11307,N_9820);
nor U13591 (N_13591,N_9321,N_8466);
nor U13592 (N_13592,N_9201,N_11260);
or U13593 (N_13593,N_9475,N_10419);
or U13594 (N_13594,N_10200,N_9274);
and U13595 (N_13595,N_9052,N_11005);
nand U13596 (N_13596,N_8042,N_9108);
nor U13597 (N_13597,N_10477,N_11308);
and U13598 (N_13598,N_10136,N_11474);
or U13599 (N_13599,N_11125,N_9973);
and U13600 (N_13600,N_10455,N_10971);
nor U13601 (N_13601,N_9227,N_10425);
nand U13602 (N_13602,N_9044,N_11925);
nand U13603 (N_13603,N_9821,N_10950);
or U13604 (N_13604,N_8327,N_10668);
or U13605 (N_13605,N_11605,N_11428);
xnor U13606 (N_13606,N_10669,N_8307);
nor U13607 (N_13607,N_10097,N_11594);
and U13608 (N_13608,N_10739,N_8969);
or U13609 (N_13609,N_8700,N_9139);
or U13610 (N_13610,N_9758,N_8868);
or U13611 (N_13611,N_8190,N_11560);
and U13612 (N_13612,N_9302,N_11376);
xor U13613 (N_13613,N_8565,N_10866);
and U13614 (N_13614,N_8266,N_10181);
or U13615 (N_13615,N_11654,N_11409);
nand U13616 (N_13616,N_8022,N_9346);
or U13617 (N_13617,N_10081,N_8074);
xor U13618 (N_13618,N_9721,N_11685);
nand U13619 (N_13619,N_11575,N_10356);
nor U13620 (N_13620,N_9608,N_8740);
nor U13621 (N_13621,N_9667,N_8606);
or U13622 (N_13622,N_8196,N_10792);
xnor U13623 (N_13623,N_8514,N_8758);
and U13624 (N_13624,N_10582,N_9437);
or U13625 (N_13625,N_11822,N_8467);
or U13626 (N_13626,N_9966,N_10066);
or U13627 (N_13627,N_8269,N_9465);
and U13628 (N_13628,N_8618,N_9995);
nor U13629 (N_13629,N_10217,N_9592);
nor U13630 (N_13630,N_11830,N_10957);
or U13631 (N_13631,N_11837,N_11903);
or U13632 (N_13632,N_9566,N_11708);
or U13633 (N_13633,N_10091,N_11023);
or U13634 (N_13634,N_9967,N_11298);
and U13635 (N_13635,N_8463,N_9955);
or U13636 (N_13636,N_8325,N_11961);
or U13637 (N_13637,N_9638,N_10547);
and U13638 (N_13638,N_10758,N_9840);
xnor U13639 (N_13639,N_11606,N_9035);
xor U13640 (N_13640,N_9273,N_11894);
nor U13641 (N_13641,N_11537,N_10126);
or U13642 (N_13642,N_10404,N_11831);
and U13643 (N_13643,N_8428,N_10113);
nor U13644 (N_13644,N_8397,N_11481);
nor U13645 (N_13645,N_8193,N_9846);
or U13646 (N_13646,N_11216,N_8299);
and U13647 (N_13647,N_9115,N_9835);
nand U13648 (N_13648,N_10988,N_11798);
or U13649 (N_13649,N_8991,N_9162);
and U13650 (N_13650,N_10176,N_8742);
or U13651 (N_13651,N_8131,N_9857);
or U13652 (N_13652,N_8462,N_10426);
or U13653 (N_13653,N_8669,N_9398);
and U13654 (N_13654,N_8112,N_9778);
nand U13655 (N_13655,N_9031,N_9580);
or U13656 (N_13656,N_8205,N_10330);
or U13657 (N_13657,N_11524,N_9519);
or U13658 (N_13658,N_9314,N_11665);
nand U13659 (N_13659,N_10631,N_8075);
nor U13660 (N_13660,N_10374,N_9557);
and U13661 (N_13661,N_8132,N_11632);
or U13662 (N_13662,N_11367,N_8936);
nand U13663 (N_13663,N_8926,N_11299);
or U13664 (N_13664,N_9655,N_8684);
xnor U13665 (N_13665,N_8441,N_11697);
nor U13666 (N_13666,N_8847,N_9540);
nand U13667 (N_13667,N_11802,N_9243);
nor U13668 (N_13668,N_11907,N_10423);
nor U13669 (N_13669,N_11334,N_8170);
or U13670 (N_13670,N_8015,N_9105);
or U13671 (N_13671,N_8276,N_8518);
nand U13672 (N_13672,N_8208,N_9759);
and U13673 (N_13673,N_10011,N_10191);
xor U13674 (N_13674,N_9797,N_8600);
and U13675 (N_13675,N_8350,N_8685);
nand U13676 (N_13676,N_11676,N_10876);
and U13677 (N_13677,N_9131,N_8346);
or U13678 (N_13678,N_8031,N_9763);
xnor U13679 (N_13679,N_10280,N_11851);
nand U13680 (N_13680,N_11704,N_8595);
and U13681 (N_13681,N_11833,N_10002);
nand U13682 (N_13682,N_8211,N_11707);
xnor U13683 (N_13683,N_9965,N_11765);
nand U13684 (N_13684,N_8785,N_10243);
nand U13685 (N_13685,N_9668,N_10694);
and U13686 (N_13686,N_9997,N_10079);
or U13687 (N_13687,N_9300,N_10018);
or U13688 (N_13688,N_9593,N_10656);
nor U13689 (N_13689,N_8787,N_11753);
nand U13690 (N_13690,N_8427,N_10448);
or U13691 (N_13691,N_10884,N_8316);
nor U13692 (N_13692,N_8930,N_11546);
and U13693 (N_13693,N_11194,N_8253);
nand U13694 (N_13694,N_11736,N_10350);
or U13695 (N_13695,N_11195,N_11806);
and U13696 (N_13696,N_8239,N_9810);
nand U13697 (N_13697,N_10913,N_8776);
or U13698 (N_13698,N_11459,N_9582);
nand U13699 (N_13699,N_10856,N_9939);
nand U13700 (N_13700,N_8279,N_8451);
nor U13701 (N_13701,N_9914,N_10557);
nand U13702 (N_13702,N_9704,N_9802);
nor U13703 (N_13703,N_10999,N_8830);
nor U13704 (N_13704,N_9247,N_9352);
or U13705 (N_13705,N_10925,N_8386);
nand U13706 (N_13706,N_9338,N_10056);
and U13707 (N_13707,N_11303,N_10007);
nand U13708 (N_13708,N_8524,N_9946);
nand U13709 (N_13709,N_8854,N_9565);
nand U13710 (N_13710,N_11946,N_9969);
nand U13711 (N_13711,N_10738,N_10970);
nor U13712 (N_13712,N_11627,N_11896);
or U13713 (N_13713,N_10392,N_11508);
nor U13714 (N_13714,N_10105,N_9450);
xnor U13715 (N_13715,N_11577,N_8909);
or U13716 (N_13716,N_11035,N_10286);
and U13717 (N_13717,N_9354,N_11010);
nor U13718 (N_13718,N_10408,N_11589);
or U13719 (N_13719,N_10438,N_11784);
nand U13720 (N_13720,N_9813,N_8081);
nand U13721 (N_13721,N_8616,N_11106);
nor U13722 (N_13722,N_10208,N_11814);
xor U13723 (N_13723,N_9612,N_11090);
xnor U13724 (N_13724,N_9016,N_11345);
nand U13725 (N_13725,N_10177,N_8367);
nor U13726 (N_13726,N_9343,N_10615);
nand U13727 (N_13727,N_8587,N_10319);
and U13728 (N_13728,N_11394,N_8165);
xnor U13729 (N_13729,N_8319,N_10266);
nand U13730 (N_13730,N_11588,N_9013);
and U13731 (N_13731,N_8519,N_11518);
nand U13732 (N_13732,N_11063,N_10569);
and U13733 (N_13733,N_9948,N_11789);
and U13734 (N_13734,N_11256,N_11192);
nand U13735 (N_13735,N_9573,N_10306);
xor U13736 (N_13736,N_9218,N_11725);
and U13737 (N_13737,N_9999,N_9080);
or U13738 (N_13738,N_9092,N_8310);
and U13739 (N_13739,N_11051,N_9729);
or U13740 (N_13740,N_10358,N_10010);
or U13741 (N_13741,N_11209,N_11951);
xnor U13742 (N_13742,N_11982,N_11958);
nand U13743 (N_13743,N_9132,N_10699);
or U13744 (N_13744,N_9351,N_10580);
nor U13745 (N_13745,N_10853,N_9542);
nand U13746 (N_13746,N_10566,N_8525);
nand U13747 (N_13747,N_9501,N_9106);
nand U13748 (N_13748,N_8361,N_8458);
and U13749 (N_13749,N_11954,N_11696);
and U13750 (N_13750,N_9894,N_8894);
nor U13751 (N_13751,N_10106,N_8395);
or U13752 (N_13752,N_9793,N_11781);
nor U13753 (N_13753,N_10470,N_11590);
and U13754 (N_13754,N_11650,N_8660);
nand U13755 (N_13755,N_9458,N_11980);
nor U13756 (N_13756,N_10907,N_8296);
nor U13757 (N_13757,N_8066,N_9665);
or U13758 (N_13758,N_9435,N_10406);
nand U13759 (N_13759,N_9210,N_11534);
xnor U13760 (N_13760,N_11237,N_8476);
nand U13761 (N_13761,N_11053,N_11137);
nand U13762 (N_13762,N_11058,N_11215);
and U13763 (N_13763,N_8706,N_10158);
and U13764 (N_13764,N_10604,N_8399);
nor U13765 (N_13765,N_9381,N_8357);
nor U13766 (N_13766,N_11916,N_9603);
and U13767 (N_13767,N_8934,N_11808);
nor U13768 (N_13768,N_8444,N_9719);
and U13769 (N_13769,N_10050,N_10610);
nand U13770 (N_13770,N_9661,N_10361);
and U13771 (N_13771,N_9853,N_8792);
or U13772 (N_13772,N_8857,N_10131);
or U13773 (N_13773,N_8737,N_10926);
nor U13774 (N_13774,N_11718,N_10170);
nor U13775 (N_13775,N_10065,N_10683);
or U13776 (N_13776,N_8526,N_10624);
nand U13777 (N_13777,N_9876,N_9233);
xnor U13778 (N_13778,N_9111,N_11721);
and U13779 (N_13779,N_9550,N_8429);
nor U13780 (N_13780,N_11316,N_11427);
or U13781 (N_13781,N_11326,N_8336);
xor U13782 (N_13782,N_9196,N_9214);
or U13783 (N_13783,N_9257,N_11533);
nor U13784 (N_13784,N_8823,N_11025);
or U13785 (N_13785,N_8219,N_10363);
or U13786 (N_13786,N_8848,N_9660);
xnor U13787 (N_13787,N_11462,N_8505);
nand U13788 (N_13788,N_8277,N_8828);
and U13789 (N_13789,N_10749,N_8655);
or U13790 (N_13790,N_8330,N_10130);
or U13791 (N_13791,N_9897,N_8831);
nor U13792 (N_13792,N_9926,N_10860);
nor U13793 (N_13793,N_8864,N_8994);
and U13794 (N_13794,N_8739,N_9074);
nor U13795 (N_13795,N_8709,N_10009);
xor U13796 (N_13796,N_11164,N_9662);
nand U13797 (N_13797,N_8562,N_8392);
or U13798 (N_13798,N_10589,N_8320);
or U13799 (N_13799,N_9479,N_10536);
nand U13800 (N_13800,N_10766,N_10534);
nor U13801 (N_13801,N_11730,N_9248);
nand U13802 (N_13802,N_10824,N_9027);
and U13803 (N_13803,N_10969,N_10332);
and U13804 (N_13804,N_10917,N_9986);
nor U13805 (N_13805,N_8403,N_10908);
and U13806 (N_13806,N_10888,N_10021);
nor U13807 (N_13807,N_9128,N_10744);
and U13808 (N_13808,N_10616,N_10543);
nand U13809 (N_13809,N_8661,N_9604);
nor U13810 (N_13810,N_9738,N_9695);
xor U13811 (N_13811,N_8695,N_9296);
nand U13812 (N_13812,N_11673,N_11296);
nor U13813 (N_13813,N_8682,N_10588);
nand U13814 (N_13814,N_10215,N_9157);
and U13815 (N_13815,N_8961,N_10929);
or U13816 (N_13816,N_9775,N_9420);
nand U13817 (N_13817,N_10302,N_10754);
and U13818 (N_13818,N_8771,N_10019);
and U13819 (N_13819,N_11690,N_9142);
xor U13820 (N_13820,N_11715,N_11921);
nand U13821 (N_13821,N_8577,N_8390);
and U13822 (N_13822,N_8993,N_8900);
nor U13823 (N_13823,N_9093,N_10657);
or U13824 (N_13824,N_10468,N_9466);
xnor U13825 (N_13825,N_11733,N_11829);
and U13826 (N_13826,N_9535,N_11792);
or U13827 (N_13827,N_9133,N_11701);
xnor U13828 (N_13828,N_11882,N_11235);
nand U13829 (N_13829,N_8754,N_11245);
nor U13830 (N_13830,N_9019,N_9596);
or U13831 (N_13831,N_8955,N_10774);
and U13832 (N_13832,N_10322,N_11469);
or U13833 (N_13833,N_10918,N_10951);
or U13834 (N_13834,N_10101,N_11898);
xor U13835 (N_13835,N_11611,N_10487);
xnor U13836 (N_13836,N_8547,N_8878);
nand U13837 (N_13837,N_9489,N_8308);
nor U13838 (N_13838,N_10121,N_11297);
nor U13839 (N_13839,N_11030,N_11176);
xor U13840 (N_13840,N_11174,N_11365);
nand U13841 (N_13841,N_11867,N_8263);
nand U13842 (N_13842,N_9502,N_9613);
or U13843 (N_13843,N_8523,N_9951);
xnor U13844 (N_13844,N_8867,N_9545);
and U13845 (N_13845,N_9689,N_11283);
or U13846 (N_13846,N_10474,N_9253);
nor U13847 (N_13847,N_9231,N_8772);
or U13848 (N_13848,N_11571,N_10720);
or U13849 (N_13849,N_10919,N_8003);
nand U13850 (N_13850,N_10240,N_11771);
or U13851 (N_13851,N_8278,N_11752);
xor U13852 (N_13852,N_10490,N_10654);
xor U13853 (N_13853,N_9395,N_11915);
nor U13854 (N_13854,N_9754,N_11142);
and U13855 (N_13855,N_11319,N_10736);
nand U13856 (N_13856,N_11662,N_9355);
xnor U13857 (N_13857,N_9249,N_9078);
nand U13858 (N_13858,N_8473,N_8786);
and U13859 (N_13859,N_10492,N_10412);
or U13860 (N_13860,N_10648,N_8515);
xor U13861 (N_13861,N_10695,N_11000);
and U13862 (N_13862,N_10651,N_9816);
and U13863 (N_13863,N_11585,N_11489);
and U13864 (N_13864,N_10023,N_9073);
nand U13865 (N_13865,N_11396,N_8637);
nand U13866 (N_13866,N_10039,N_8871);
nor U13867 (N_13867,N_9772,N_9494);
nand U13868 (N_13868,N_8983,N_8743);
nand U13869 (N_13869,N_11490,N_11815);
or U13870 (N_13870,N_9158,N_8285);
and U13871 (N_13871,N_8049,N_8731);
or U13872 (N_13872,N_11315,N_8270);
and U13873 (N_13873,N_8940,N_9188);
or U13874 (N_13874,N_11207,N_9185);
nand U13875 (N_13875,N_9014,N_9485);
nand U13876 (N_13876,N_8456,N_11743);
nor U13877 (N_13877,N_10197,N_11062);
nand U13878 (N_13878,N_8158,N_11273);
xnor U13879 (N_13879,N_11861,N_8137);
nand U13880 (N_13880,N_10180,N_8348);
nor U13881 (N_13881,N_10061,N_11214);
nor U13882 (N_13882,N_11840,N_10606);
or U13883 (N_13883,N_8475,N_9632);
xnor U13884 (N_13884,N_11929,N_9642);
or U13885 (N_13885,N_8887,N_11395);
or U13886 (N_13886,N_10875,N_11412);
xor U13887 (N_13887,N_8548,N_11677);
nor U13888 (N_13888,N_9217,N_9771);
or U13889 (N_13889,N_9877,N_10254);
nor U13890 (N_13890,N_10816,N_10367);
or U13891 (N_13891,N_9556,N_11820);
and U13892 (N_13892,N_11848,N_10171);
nand U13893 (N_13893,N_10983,N_8810);
and U13894 (N_13894,N_8248,N_10721);
and U13895 (N_13895,N_10596,N_11803);
nand U13896 (N_13896,N_10099,N_11729);
and U13897 (N_13897,N_8072,N_10001);
or U13898 (N_13898,N_8478,N_10805);
nand U13899 (N_13899,N_11959,N_8023);
nand U13900 (N_13900,N_8430,N_10463);
and U13901 (N_13901,N_9140,N_11426);
or U13902 (N_13902,N_10303,N_11356);
or U13903 (N_13903,N_10494,N_8157);
nor U13904 (N_13904,N_9688,N_9410);
or U13905 (N_13905,N_9375,N_8401);
nor U13906 (N_13906,N_10979,N_11507);
nor U13907 (N_13907,N_9696,N_10719);
nor U13908 (N_13908,N_9282,N_8843);
nand U13909 (N_13909,N_10946,N_8314);
nand U13910 (N_13910,N_9927,N_11012);
or U13911 (N_13911,N_11634,N_11204);
nand U13912 (N_13912,N_8481,N_10567);
nand U13913 (N_13913,N_9806,N_9733);
or U13914 (N_13914,N_8360,N_9977);
and U13915 (N_13915,N_8711,N_11754);
xor U13916 (N_13916,N_10832,N_8971);
or U13917 (N_13917,N_9492,N_8236);
and U13918 (N_13918,N_11423,N_11934);
and U13919 (N_13919,N_11878,N_11835);
nand U13920 (N_13920,N_9419,N_8840);
nor U13921 (N_13921,N_8588,N_11271);
nor U13922 (N_13922,N_10682,N_10264);
nor U13923 (N_13923,N_10440,N_9715);
and U13924 (N_13924,N_10288,N_10344);
xor U13925 (N_13925,N_9187,N_8815);
xor U13926 (N_13926,N_9832,N_8187);
or U13927 (N_13927,N_9028,N_8446);
and U13928 (N_13928,N_10249,N_11258);
and U13929 (N_13929,N_11372,N_9393);
or U13930 (N_13930,N_11095,N_11093);
nand U13931 (N_13931,N_10218,N_10525);
nand U13932 (N_13932,N_10889,N_10770);
or U13933 (N_13933,N_11669,N_11722);
nand U13934 (N_13934,N_11021,N_11746);
nor U13935 (N_13935,N_9148,N_9842);
or U13936 (N_13936,N_10486,N_8037);
or U13937 (N_13937,N_8902,N_9443);
nor U13938 (N_13938,N_9234,N_10220);
nor U13939 (N_13939,N_8321,N_10430);
and U13940 (N_13940,N_9281,N_9283);
nand U13941 (N_13941,N_10441,N_9713);
nand U13942 (N_13942,N_10768,N_11013);
and U13943 (N_13943,N_8889,N_8311);
and U13944 (N_13944,N_8552,N_8470);
xnor U13945 (N_13945,N_11693,N_8851);
or U13946 (N_13946,N_11684,N_11856);
and U13947 (N_13947,N_10391,N_8643);
nor U13948 (N_13948,N_10493,N_10782);
nor U13949 (N_13949,N_11616,N_9365);
nand U13950 (N_13950,N_11527,N_9127);
nand U13951 (N_13951,N_8334,N_11117);
xor U13952 (N_13952,N_10246,N_11749);
nand U13953 (N_13953,N_8493,N_10265);
xnor U13954 (N_13954,N_8778,N_11322);
nand U13955 (N_13955,N_9163,N_10706);
or U13956 (N_13956,N_11928,N_9478);
or U13957 (N_13957,N_11377,N_11895);
and U13958 (N_13958,N_9426,N_9211);
or U13959 (N_13959,N_9207,N_11501);
nand U13960 (N_13960,N_10040,N_9391);
and U13961 (N_13961,N_10664,N_8027);
or U13962 (N_13962,N_11120,N_10357);
xnor U13963 (N_13963,N_8881,N_9931);
nand U13964 (N_13964,N_9482,N_8432);
nand U13965 (N_13965,N_8402,N_9135);
and U13966 (N_13966,N_11208,N_10084);
or U13967 (N_13967,N_10798,N_8070);
or U13968 (N_13968,N_10808,N_10481);
and U13969 (N_13969,N_11197,N_9928);
nand U13970 (N_13970,N_9221,N_10714);
nand U13971 (N_13971,N_9117,N_11220);
or U13972 (N_13972,N_9047,N_9602);
nor U13973 (N_13973,N_9915,N_10781);
and U13974 (N_13974,N_11181,N_10086);
nor U13975 (N_13975,N_8770,N_10143);
nand U13976 (N_13976,N_8381,N_9280);
or U13977 (N_13977,N_8544,N_8838);
and U13978 (N_13978,N_9942,N_11997);
nor U13979 (N_13979,N_9947,N_9544);
nand U13980 (N_13980,N_9449,N_11766);
and U13981 (N_13981,N_10528,N_9742);
or U13982 (N_13982,N_8841,N_11184);
nor U13983 (N_13983,N_10359,N_10956);
nor U13984 (N_13984,N_8369,N_8697);
nor U13985 (N_13985,N_8497,N_9242);
nand U13986 (N_13986,N_11355,N_11357);
or U13987 (N_13987,N_9378,N_10820);
nand U13988 (N_13988,N_8784,N_8063);
nand U13989 (N_13989,N_11232,N_11531);
or U13990 (N_13990,N_11418,N_10622);
and U13991 (N_13991,N_9086,N_8500);
and U13992 (N_13992,N_8503,N_11066);
or U13993 (N_13993,N_11931,N_11623);
or U13994 (N_13994,N_8162,N_9673);
and U13995 (N_13995,N_10446,N_8982);
nand U13996 (N_13996,N_11088,N_11482);
nor U13997 (N_13997,N_10142,N_8928);
and U13998 (N_13998,N_10196,N_8108);
nor U13999 (N_13999,N_8989,N_10544);
nor U14000 (N_14000,N_10699,N_9745);
nor U14001 (N_14001,N_9909,N_10105);
nor U14002 (N_14002,N_10075,N_10322);
or U14003 (N_14003,N_8830,N_8037);
and U14004 (N_14004,N_9403,N_9052);
nor U14005 (N_14005,N_8468,N_8643);
nand U14006 (N_14006,N_11828,N_10306);
and U14007 (N_14007,N_8509,N_8817);
xnor U14008 (N_14008,N_10818,N_9265);
xnor U14009 (N_14009,N_10300,N_9161);
or U14010 (N_14010,N_11925,N_9087);
nand U14011 (N_14011,N_9000,N_10435);
and U14012 (N_14012,N_8593,N_10424);
nor U14013 (N_14013,N_8451,N_8548);
or U14014 (N_14014,N_10653,N_10056);
nand U14015 (N_14015,N_9941,N_11155);
and U14016 (N_14016,N_11221,N_8253);
or U14017 (N_14017,N_9487,N_11135);
nor U14018 (N_14018,N_10132,N_10940);
or U14019 (N_14019,N_11496,N_11822);
or U14020 (N_14020,N_10057,N_8187);
nand U14021 (N_14021,N_10420,N_10011);
nor U14022 (N_14022,N_9689,N_8394);
xnor U14023 (N_14023,N_8530,N_8936);
nand U14024 (N_14024,N_10865,N_8742);
and U14025 (N_14025,N_9909,N_10068);
nor U14026 (N_14026,N_10137,N_10610);
xnor U14027 (N_14027,N_8774,N_8010);
or U14028 (N_14028,N_8662,N_9143);
nand U14029 (N_14029,N_10631,N_10336);
and U14030 (N_14030,N_8418,N_8217);
xnor U14031 (N_14031,N_8317,N_9589);
nand U14032 (N_14032,N_9775,N_10625);
xnor U14033 (N_14033,N_11823,N_11479);
or U14034 (N_14034,N_10091,N_9504);
and U14035 (N_14035,N_9407,N_11666);
nand U14036 (N_14036,N_11137,N_8319);
nor U14037 (N_14037,N_8565,N_8124);
nand U14038 (N_14038,N_11820,N_10916);
and U14039 (N_14039,N_10216,N_9887);
nor U14040 (N_14040,N_9491,N_9570);
and U14041 (N_14041,N_11481,N_10402);
nor U14042 (N_14042,N_10710,N_9858);
nor U14043 (N_14043,N_8096,N_10822);
and U14044 (N_14044,N_10185,N_9908);
nand U14045 (N_14045,N_10437,N_9182);
xor U14046 (N_14046,N_11886,N_11671);
and U14047 (N_14047,N_8520,N_10749);
or U14048 (N_14048,N_8312,N_10150);
xnor U14049 (N_14049,N_8782,N_11832);
or U14050 (N_14050,N_11012,N_10414);
and U14051 (N_14051,N_11647,N_11933);
nor U14052 (N_14052,N_10406,N_10942);
or U14053 (N_14053,N_11109,N_8623);
nor U14054 (N_14054,N_10716,N_11552);
xor U14055 (N_14055,N_10813,N_9034);
nor U14056 (N_14056,N_9513,N_8865);
or U14057 (N_14057,N_10887,N_8106);
and U14058 (N_14058,N_8985,N_9395);
nand U14059 (N_14059,N_8285,N_11310);
nand U14060 (N_14060,N_11633,N_11371);
and U14061 (N_14061,N_9062,N_10062);
nand U14062 (N_14062,N_8401,N_10597);
and U14063 (N_14063,N_10147,N_8900);
and U14064 (N_14064,N_10673,N_9606);
or U14065 (N_14065,N_11890,N_9799);
xnor U14066 (N_14066,N_11588,N_9165);
nand U14067 (N_14067,N_10288,N_8714);
and U14068 (N_14068,N_10458,N_8940);
nand U14069 (N_14069,N_10515,N_10149);
nand U14070 (N_14070,N_8705,N_8347);
or U14071 (N_14071,N_8986,N_8537);
nand U14072 (N_14072,N_9492,N_8928);
nor U14073 (N_14073,N_10324,N_11821);
xor U14074 (N_14074,N_9942,N_9457);
nand U14075 (N_14075,N_11746,N_9980);
nor U14076 (N_14076,N_8142,N_11837);
xnor U14077 (N_14077,N_9950,N_10731);
nor U14078 (N_14078,N_10616,N_8420);
or U14079 (N_14079,N_9173,N_10067);
nand U14080 (N_14080,N_10040,N_8618);
xnor U14081 (N_14081,N_8333,N_8390);
and U14082 (N_14082,N_11088,N_10261);
xor U14083 (N_14083,N_10310,N_9919);
nor U14084 (N_14084,N_9333,N_10029);
nand U14085 (N_14085,N_10324,N_10171);
nand U14086 (N_14086,N_9932,N_10273);
and U14087 (N_14087,N_11533,N_10655);
xnor U14088 (N_14088,N_11194,N_11378);
or U14089 (N_14089,N_8636,N_9156);
nor U14090 (N_14090,N_8687,N_9138);
and U14091 (N_14091,N_8973,N_10659);
and U14092 (N_14092,N_8706,N_9377);
and U14093 (N_14093,N_9709,N_9128);
and U14094 (N_14094,N_8684,N_9392);
nor U14095 (N_14095,N_11829,N_10435);
nand U14096 (N_14096,N_8516,N_9444);
and U14097 (N_14097,N_10797,N_9135);
and U14098 (N_14098,N_10271,N_8654);
nor U14099 (N_14099,N_10074,N_8257);
nor U14100 (N_14100,N_11499,N_8639);
nand U14101 (N_14101,N_8899,N_8529);
or U14102 (N_14102,N_8538,N_8142);
and U14103 (N_14103,N_9947,N_10068);
and U14104 (N_14104,N_11562,N_8089);
nand U14105 (N_14105,N_11646,N_11054);
nand U14106 (N_14106,N_11900,N_10114);
and U14107 (N_14107,N_11059,N_9977);
xnor U14108 (N_14108,N_8865,N_11558);
nand U14109 (N_14109,N_10229,N_11691);
nand U14110 (N_14110,N_10291,N_9896);
nand U14111 (N_14111,N_8334,N_10226);
nand U14112 (N_14112,N_9462,N_8786);
and U14113 (N_14113,N_8497,N_9218);
or U14114 (N_14114,N_10052,N_10943);
and U14115 (N_14115,N_8104,N_9633);
or U14116 (N_14116,N_8959,N_8939);
or U14117 (N_14117,N_9158,N_11577);
nand U14118 (N_14118,N_9991,N_8722);
nand U14119 (N_14119,N_9522,N_9871);
nand U14120 (N_14120,N_11078,N_8772);
nand U14121 (N_14121,N_9514,N_10905);
and U14122 (N_14122,N_10171,N_11833);
and U14123 (N_14123,N_11512,N_10892);
and U14124 (N_14124,N_8338,N_9613);
nor U14125 (N_14125,N_11210,N_10045);
nor U14126 (N_14126,N_11481,N_10011);
nand U14127 (N_14127,N_9042,N_9063);
or U14128 (N_14128,N_8899,N_9967);
and U14129 (N_14129,N_8368,N_10031);
nand U14130 (N_14130,N_9420,N_9048);
or U14131 (N_14131,N_11837,N_8312);
nor U14132 (N_14132,N_10323,N_11362);
xnor U14133 (N_14133,N_8066,N_11031);
and U14134 (N_14134,N_8276,N_8987);
nor U14135 (N_14135,N_11975,N_11998);
nand U14136 (N_14136,N_11154,N_10785);
and U14137 (N_14137,N_8506,N_11463);
and U14138 (N_14138,N_11722,N_10068);
nand U14139 (N_14139,N_11808,N_8702);
xnor U14140 (N_14140,N_10409,N_8778);
or U14141 (N_14141,N_10958,N_9016);
nand U14142 (N_14142,N_10654,N_10675);
nand U14143 (N_14143,N_9290,N_9821);
and U14144 (N_14144,N_11373,N_11996);
nand U14145 (N_14145,N_8609,N_10711);
xor U14146 (N_14146,N_11709,N_8478);
nand U14147 (N_14147,N_9145,N_10081);
nor U14148 (N_14148,N_10424,N_8665);
or U14149 (N_14149,N_9224,N_8696);
xnor U14150 (N_14150,N_8099,N_10884);
nand U14151 (N_14151,N_8874,N_11527);
nand U14152 (N_14152,N_10018,N_8293);
nor U14153 (N_14153,N_10489,N_9821);
nand U14154 (N_14154,N_11443,N_8224);
nor U14155 (N_14155,N_10279,N_10667);
nor U14156 (N_14156,N_10667,N_10523);
nand U14157 (N_14157,N_10669,N_8357);
and U14158 (N_14158,N_9180,N_9902);
and U14159 (N_14159,N_8261,N_8644);
nand U14160 (N_14160,N_9399,N_11224);
nor U14161 (N_14161,N_8628,N_8454);
and U14162 (N_14162,N_9781,N_8939);
or U14163 (N_14163,N_10428,N_8591);
nor U14164 (N_14164,N_9955,N_10786);
nand U14165 (N_14165,N_10656,N_11390);
nand U14166 (N_14166,N_10538,N_8632);
nor U14167 (N_14167,N_10913,N_8542);
nor U14168 (N_14168,N_9347,N_10818);
or U14169 (N_14169,N_10979,N_10419);
xor U14170 (N_14170,N_8778,N_10135);
xnor U14171 (N_14171,N_9276,N_10214);
nand U14172 (N_14172,N_10437,N_9223);
nand U14173 (N_14173,N_11953,N_9425);
or U14174 (N_14174,N_11510,N_10863);
or U14175 (N_14175,N_11609,N_9562);
nand U14176 (N_14176,N_8992,N_9568);
nor U14177 (N_14177,N_9420,N_11734);
or U14178 (N_14178,N_11971,N_10724);
and U14179 (N_14179,N_11161,N_10170);
and U14180 (N_14180,N_10340,N_11881);
and U14181 (N_14181,N_10838,N_8893);
nand U14182 (N_14182,N_10068,N_8679);
or U14183 (N_14183,N_9644,N_8852);
and U14184 (N_14184,N_8715,N_8416);
or U14185 (N_14185,N_10008,N_10444);
or U14186 (N_14186,N_8032,N_11870);
nand U14187 (N_14187,N_8016,N_10623);
nand U14188 (N_14188,N_9309,N_8634);
nand U14189 (N_14189,N_11550,N_9344);
or U14190 (N_14190,N_11547,N_10441);
nor U14191 (N_14191,N_9678,N_11749);
and U14192 (N_14192,N_11966,N_8381);
nor U14193 (N_14193,N_10383,N_11036);
nor U14194 (N_14194,N_9137,N_10931);
xor U14195 (N_14195,N_9581,N_9567);
and U14196 (N_14196,N_9624,N_9018);
nand U14197 (N_14197,N_11936,N_8697);
nand U14198 (N_14198,N_10251,N_8041);
or U14199 (N_14199,N_9445,N_9526);
and U14200 (N_14200,N_11424,N_11105);
and U14201 (N_14201,N_10482,N_11207);
and U14202 (N_14202,N_10034,N_8779);
or U14203 (N_14203,N_9225,N_8989);
nand U14204 (N_14204,N_10775,N_10421);
nand U14205 (N_14205,N_8364,N_9579);
and U14206 (N_14206,N_10163,N_9402);
nand U14207 (N_14207,N_8963,N_10951);
nor U14208 (N_14208,N_9244,N_9646);
nor U14209 (N_14209,N_11782,N_10238);
xor U14210 (N_14210,N_11110,N_11942);
nor U14211 (N_14211,N_9316,N_8041);
and U14212 (N_14212,N_9528,N_8163);
nand U14213 (N_14213,N_8891,N_8133);
and U14214 (N_14214,N_9404,N_11224);
or U14215 (N_14215,N_9366,N_10996);
nand U14216 (N_14216,N_11934,N_8346);
and U14217 (N_14217,N_10403,N_10497);
nand U14218 (N_14218,N_10227,N_10299);
and U14219 (N_14219,N_11037,N_11659);
nand U14220 (N_14220,N_9225,N_9621);
xnor U14221 (N_14221,N_10115,N_8149);
nand U14222 (N_14222,N_9250,N_10504);
nand U14223 (N_14223,N_9462,N_9623);
or U14224 (N_14224,N_10161,N_10775);
or U14225 (N_14225,N_10696,N_11031);
and U14226 (N_14226,N_10441,N_8974);
or U14227 (N_14227,N_11576,N_11312);
nor U14228 (N_14228,N_11884,N_8423);
and U14229 (N_14229,N_9330,N_9443);
nand U14230 (N_14230,N_10377,N_8150);
or U14231 (N_14231,N_9064,N_9818);
nor U14232 (N_14232,N_11554,N_10184);
nor U14233 (N_14233,N_11322,N_9223);
nand U14234 (N_14234,N_10110,N_11475);
or U14235 (N_14235,N_8100,N_8307);
nand U14236 (N_14236,N_10133,N_10437);
and U14237 (N_14237,N_11474,N_10978);
and U14238 (N_14238,N_8381,N_10108);
xnor U14239 (N_14239,N_8543,N_8817);
or U14240 (N_14240,N_9028,N_8234);
and U14241 (N_14241,N_11213,N_9918);
xnor U14242 (N_14242,N_9527,N_8022);
or U14243 (N_14243,N_10874,N_8887);
nand U14244 (N_14244,N_11710,N_8116);
or U14245 (N_14245,N_9441,N_11556);
nand U14246 (N_14246,N_10224,N_11077);
nand U14247 (N_14247,N_10312,N_10924);
nand U14248 (N_14248,N_10614,N_8345);
xor U14249 (N_14249,N_10909,N_8535);
nor U14250 (N_14250,N_10682,N_10218);
nand U14251 (N_14251,N_10062,N_10521);
or U14252 (N_14252,N_10149,N_8846);
nand U14253 (N_14253,N_9822,N_8345);
nor U14254 (N_14254,N_8009,N_10102);
or U14255 (N_14255,N_8499,N_11527);
nand U14256 (N_14256,N_11186,N_8053);
nand U14257 (N_14257,N_10509,N_10824);
and U14258 (N_14258,N_9194,N_11451);
nand U14259 (N_14259,N_11146,N_11004);
and U14260 (N_14260,N_11432,N_8500);
nand U14261 (N_14261,N_8809,N_9078);
nor U14262 (N_14262,N_8875,N_9261);
nand U14263 (N_14263,N_8607,N_10781);
or U14264 (N_14264,N_8412,N_9719);
nand U14265 (N_14265,N_10530,N_11113);
or U14266 (N_14266,N_10651,N_10338);
nor U14267 (N_14267,N_11021,N_11335);
nor U14268 (N_14268,N_9893,N_10905);
or U14269 (N_14269,N_8396,N_9919);
xor U14270 (N_14270,N_8002,N_11594);
and U14271 (N_14271,N_9996,N_11920);
and U14272 (N_14272,N_9248,N_8864);
xor U14273 (N_14273,N_11369,N_9954);
and U14274 (N_14274,N_9565,N_9104);
and U14275 (N_14275,N_11062,N_11071);
nand U14276 (N_14276,N_11845,N_9870);
nor U14277 (N_14277,N_9586,N_11119);
nand U14278 (N_14278,N_9582,N_9211);
nor U14279 (N_14279,N_10663,N_9416);
or U14280 (N_14280,N_10780,N_11667);
nor U14281 (N_14281,N_10901,N_11465);
nor U14282 (N_14282,N_11028,N_10644);
or U14283 (N_14283,N_11326,N_9433);
or U14284 (N_14284,N_11199,N_8660);
xor U14285 (N_14285,N_11869,N_10086);
and U14286 (N_14286,N_9350,N_10661);
nor U14287 (N_14287,N_9219,N_11974);
nor U14288 (N_14288,N_8832,N_11165);
nand U14289 (N_14289,N_11171,N_8080);
xor U14290 (N_14290,N_9669,N_9596);
nor U14291 (N_14291,N_10465,N_8787);
nand U14292 (N_14292,N_8847,N_8566);
and U14293 (N_14293,N_10966,N_11484);
nand U14294 (N_14294,N_11457,N_9181);
nand U14295 (N_14295,N_9211,N_11517);
nor U14296 (N_14296,N_11577,N_11463);
nand U14297 (N_14297,N_10800,N_10367);
and U14298 (N_14298,N_9949,N_10034);
or U14299 (N_14299,N_9225,N_11319);
or U14300 (N_14300,N_8475,N_10867);
nor U14301 (N_14301,N_8498,N_11700);
and U14302 (N_14302,N_9023,N_8067);
and U14303 (N_14303,N_9993,N_11260);
nand U14304 (N_14304,N_11277,N_8928);
nor U14305 (N_14305,N_8645,N_10111);
nand U14306 (N_14306,N_9590,N_9917);
nor U14307 (N_14307,N_10774,N_9248);
nand U14308 (N_14308,N_10288,N_11239);
nor U14309 (N_14309,N_9689,N_8267);
and U14310 (N_14310,N_10370,N_9573);
and U14311 (N_14311,N_10179,N_9401);
and U14312 (N_14312,N_10371,N_9528);
nand U14313 (N_14313,N_9639,N_10257);
nand U14314 (N_14314,N_9017,N_9311);
and U14315 (N_14315,N_9825,N_10565);
xor U14316 (N_14316,N_11675,N_11141);
nand U14317 (N_14317,N_9491,N_8843);
or U14318 (N_14318,N_9674,N_10435);
nand U14319 (N_14319,N_10289,N_9150);
or U14320 (N_14320,N_10427,N_10803);
and U14321 (N_14321,N_8918,N_10356);
nor U14322 (N_14322,N_8655,N_9810);
nor U14323 (N_14323,N_9079,N_10976);
or U14324 (N_14324,N_10128,N_8028);
or U14325 (N_14325,N_9837,N_9057);
nor U14326 (N_14326,N_9813,N_8602);
nor U14327 (N_14327,N_10099,N_11662);
nor U14328 (N_14328,N_8865,N_8792);
nor U14329 (N_14329,N_11723,N_11032);
and U14330 (N_14330,N_10570,N_10170);
and U14331 (N_14331,N_11891,N_8770);
or U14332 (N_14332,N_10908,N_11475);
nor U14333 (N_14333,N_9382,N_9095);
or U14334 (N_14334,N_10159,N_11197);
and U14335 (N_14335,N_9765,N_10647);
or U14336 (N_14336,N_11141,N_9404);
nor U14337 (N_14337,N_8578,N_11380);
nand U14338 (N_14338,N_11897,N_8505);
nor U14339 (N_14339,N_8684,N_11906);
nand U14340 (N_14340,N_10856,N_8215);
nor U14341 (N_14341,N_11773,N_10415);
or U14342 (N_14342,N_10852,N_9566);
nor U14343 (N_14343,N_8100,N_11461);
and U14344 (N_14344,N_11819,N_10463);
nand U14345 (N_14345,N_10464,N_9657);
or U14346 (N_14346,N_11888,N_10320);
nor U14347 (N_14347,N_10331,N_9943);
nor U14348 (N_14348,N_10693,N_10175);
nand U14349 (N_14349,N_10671,N_8994);
nor U14350 (N_14350,N_11838,N_8977);
and U14351 (N_14351,N_11976,N_11683);
nand U14352 (N_14352,N_11919,N_11376);
nand U14353 (N_14353,N_8619,N_8446);
nor U14354 (N_14354,N_8949,N_11366);
xnor U14355 (N_14355,N_8407,N_8223);
nand U14356 (N_14356,N_10706,N_10926);
and U14357 (N_14357,N_11748,N_11362);
nor U14358 (N_14358,N_9224,N_8578);
or U14359 (N_14359,N_8549,N_11967);
and U14360 (N_14360,N_10127,N_10418);
nor U14361 (N_14361,N_10023,N_11553);
and U14362 (N_14362,N_9281,N_9208);
nand U14363 (N_14363,N_10199,N_10872);
and U14364 (N_14364,N_8402,N_11133);
nand U14365 (N_14365,N_8481,N_10665);
or U14366 (N_14366,N_8327,N_11813);
nor U14367 (N_14367,N_10092,N_10656);
nand U14368 (N_14368,N_10393,N_8877);
nand U14369 (N_14369,N_9032,N_10076);
xnor U14370 (N_14370,N_11035,N_11689);
nor U14371 (N_14371,N_11555,N_8026);
nor U14372 (N_14372,N_11333,N_10348);
nand U14373 (N_14373,N_11210,N_9888);
or U14374 (N_14374,N_10555,N_10193);
nand U14375 (N_14375,N_10591,N_9013);
and U14376 (N_14376,N_9801,N_9562);
or U14377 (N_14377,N_8015,N_9807);
and U14378 (N_14378,N_8234,N_9735);
nor U14379 (N_14379,N_11352,N_10738);
and U14380 (N_14380,N_9520,N_9772);
xor U14381 (N_14381,N_10366,N_11718);
or U14382 (N_14382,N_10721,N_10986);
and U14383 (N_14383,N_8324,N_9736);
nor U14384 (N_14384,N_10583,N_11303);
and U14385 (N_14385,N_10967,N_8110);
nor U14386 (N_14386,N_9456,N_10259);
and U14387 (N_14387,N_9085,N_11624);
or U14388 (N_14388,N_11886,N_8388);
and U14389 (N_14389,N_9111,N_8739);
nor U14390 (N_14390,N_9949,N_8258);
nor U14391 (N_14391,N_10046,N_9198);
nand U14392 (N_14392,N_8021,N_11131);
nand U14393 (N_14393,N_10402,N_8287);
or U14394 (N_14394,N_10781,N_9197);
nor U14395 (N_14395,N_11002,N_11866);
nor U14396 (N_14396,N_8307,N_9318);
nand U14397 (N_14397,N_9225,N_10451);
or U14398 (N_14398,N_11803,N_10229);
or U14399 (N_14399,N_11424,N_10420);
nand U14400 (N_14400,N_9818,N_9169);
or U14401 (N_14401,N_10998,N_10526);
nor U14402 (N_14402,N_8196,N_11006);
nor U14403 (N_14403,N_10411,N_10263);
nor U14404 (N_14404,N_10194,N_8636);
or U14405 (N_14405,N_8407,N_10010);
or U14406 (N_14406,N_11549,N_9190);
nand U14407 (N_14407,N_8601,N_8282);
nand U14408 (N_14408,N_10210,N_11143);
and U14409 (N_14409,N_10080,N_11920);
nand U14410 (N_14410,N_8848,N_9851);
and U14411 (N_14411,N_8395,N_8975);
nand U14412 (N_14412,N_8214,N_9773);
and U14413 (N_14413,N_9617,N_8284);
and U14414 (N_14414,N_10873,N_11956);
and U14415 (N_14415,N_10191,N_9107);
or U14416 (N_14416,N_10779,N_10758);
or U14417 (N_14417,N_10881,N_10759);
or U14418 (N_14418,N_10716,N_11470);
xnor U14419 (N_14419,N_10629,N_9234);
nor U14420 (N_14420,N_11875,N_11829);
nand U14421 (N_14421,N_10629,N_11660);
nor U14422 (N_14422,N_10570,N_8222);
nor U14423 (N_14423,N_10320,N_11891);
xnor U14424 (N_14424,N_10643,N_11304);
xnor U14425 (N_14425,N_10437,N_10447);
xor U14426 (N_14426,N_8963,N_10699);
nor U14427 (N_14427,N_9739,N_11060);
nand U14428 (N_14428,N_9535,N_9468);
or U14429 (N_14429,N_8725,N_8311);
or U14430 (N_14430,N_8881,N_11868);
nand U14431 (N_14431,N_8380,N_8408);
nand U14432 (N_14432,N_11245,N_11837);
nor U14433 (N_14433,N_11685,N_8709);
and U14434 (N_14434,N_11543,N_10010);
and U14435 (N_14435,N_9118,N_9946);
nor U14436 (N_14436,N_11244,N_8943);
and U14437 (N_14437,N_10560,N_9706);
nand U14438 (N_14438,N_11221,N_11943);
nor U14439 (N_14439,N_8390,N_10107);
nor U14440 (N_14440,N_9210,N_8011);
nor U14441 (N_14441,N_10188,N_8228);
nand U14442 (N_14442,N_9984,N_9619);
or U14443 (N_14443,N_11196,N_9121);
and U14444 (N_14444,N_9051,N_9591);
or U14445 (N_14445,N_8683,N_8661);
nand U14446 (N_14446,N_11389,N_11135);
nor U14447 (N_14447,N_10696,N_10370);
and U14448 (N_14448,N_11280,N_9663);
nor U14449 (N_14449,N_11197,N_10262);
or U14450 (N_14450,N_9531,N_9148);
and U14451 (N_14451,N_10643,N_10114);
and U14452 (N_14452,N_8405,N_11663);
nand U14453 (N_14453,N_9005,N_9244);
nand U14454 (N_14454,N_11320,N_10875);
nand U14455 (N_14455,N_11825,N_10428);
and U14456 (N_14456,N_11796,N_9968);
and U14457 (N_14457,N_10243,N_11128);
xnor U14458 (N_14458,N_11435,N_10640);
and U14459 (N_14459,N_11554,N_9841);
nor U14460 (N_14460,N_10041,N_10554);
nand U14461 (N_14461,N_9189,N_10380);
nor U14462 (N_14462,N_10915,N_8612);
nor U14463 (N_14463,N_8733,N_11489);
or U14464 (N_14464,N_10541,N_9743);
nor U14465 (N_14465,N_8254,N_10929);
nand U14466 (N_14466,N_8324,N_8438);
nand U14467 (N_14467,N_8045,N_11387);
and U14468 (N_14468,N_10021,N_9261);
nand U14469 (N_14469,N_9201,N_8791);
nor U14470 (N_14470,N_9957,N_8606);
and U14471 (N_14471,N_9482,N_8728);
or U14472 (N_14472,N_10258,N_10603);
and U14473 (N_14473,N_11163,N_10673);
and U14474 (N_14474,N_9305,N_8902);
nor U14475 (N_14475,N_10249,N_9221);
nand U14476 (N_14476,N_9122,N_9054);
nand U14477 (N_14477,N_10544,N_9789);
or U14478 (N_14478,N_10448,N_10249);
or U14479 (N_14479,N_11046,N_10568);
xnor U14480 (N_14480,N_10504,N_11927);
xor U14481 (N_14481,N_8491,N_8615);
nor U14482 (N_14482,N_11625,N_10870);
or U14483 (N_14483,N_11267,N_10698);
nand U14484 (N_14484,N_9991,N_9993);
nand U14485 (N_14485,N_11269,N_10132);
nor U14486 (N_14486,N_8063,N_9853);
or U14487 (N_14487,N_10609,N_10531);
nor U14488 (N_14488,N_9181,N_8075);
nor U14489 (N_14489,N_11138,N_10490);
nor U14490 (N_14490,N_8006,N_11994);
or U14491 (N_14491,N_8958,N_8657);
nand U14492 (N_14492,N_8010,N_10938);
nand U14493 (N_14493,N_9554,N_10916);
or U14494 (N_14494,N_9260,N_10295);
and U14495 (N_14495,N_9971,N_11631);
or U14496 (N_14496,N_10761,N_11475);
nand U14497 (N_14497,N_9980,N_11264);
and U14498 (N_14498,N_11524,N_9290);
xnor U14499 (N_14499,N_11930,N_11954);
or U14500 (N_14500,N_9153,N_8316);
nor U14501 (N_14501,N_9879,N_8512);
or U14502 (N_14502,N_10303,N_8304);
nor U14503 (N_14503,N_8816,N_11943);
nand U14504 (N_14504,N_10578,N_9910);
or U14505 (N_14505,N_11836,N_10945);
or U14506 (N_14506,N_8023,N_10610);
nand U14507 (N_14507,N_10339,N_10301);
nand U14508 (N_14508,N_10461,N_11193);
nand U14509 (N_14509,N_8210,N_10480);
or U14510 (N_14510,N_11149,N_11549);
nand U14511 (N_14511,N_9614,N_10008);
nor U14512 (N_14512,N_11101,N_9200);
or U14513 (N_14513,N_9003,N_9220);
nand U14514 (N_14514,N_8523,N_9504);
nor U14515 (N_14515,N_11576,N_9451);
and U14516 (N_14516,N_11862,N_10139);
or U14517 (N_14517,N_8111,N_11634);
nor U14518 (N_14518,N_8975,N_10073);
nor U14519 (N_14519,N_11450,N_10908);
or U14520 (N_14520,N_11618,N_10629);
nor U14521 (N_14521,N_8609,N_9504);
and U14522 (N_14522,N_8360,N_10681);
nor U14523 (N_14523,N_9986,N_11236);
xor U14524 (N_14524,N_9616,N_8957);
nand U14525 (N_14525,N_11254,N_11705);
or U14526 (N_14526,N_11825,N_11791);
and U14527 (N_14527,N_9915,N_9990);
nor U14528 (N_14528,N_10013,N_10365);
xnor U14529 (N_14529,N_10849,N_11350);
nor U14530 (N_14530,N_10718,N_8610);
or U14531 (N_14531,N_8210,N_9594);
and U14532 (N_14532,N_10960,N_11679);
nand U14533 (N_14533,N_8630,N_11518);
or U14534 (N_14534,N_9708,N_11116);
nand U14535 (N_14535,N_11299,N_9286);
and U14536 (N_14536,N_11843,N_9621);
and U14537 (N_14537,N_8236,N_8881);
xnor U14538 (N_14538,N_8352,N_10201);
nand U14539 (N_14539,N_8423,N_8982);
xnor U14540 (N_14540,N_10292,N_11330);
or U14541 (N_14541,N_11764,N_10940);
nand U14542 (N_14542,N_9858,N_11331);
and U14543 (N_14543,N_10584,N_9723);
or U14544 (N_14544,N_9637,N_9289);
nor U14545 (N_14545,N_8081,N_11357);
or U14546 (N_14546,N_11494,N_11373);
or U14547 (N_14547,N_9597,N_9039);
nand U14548 (N_14548,N_10863,N_10268);
nor U14549 (N_14549,N_9356,N_9635);
and U14550 (N_14550,N_10147,N_9644);
or U14551 (N_14551,N_9699,N_11744);
nor U14552 (N_14552,N_9311,N_9830);
nor U14553 (N_14553,N_10500,N_10027);
nor U14554 (N_14554,N_11948,N_8242);
xnor U14555 (N_14555,N_9982,N_9626);
nor U14556 (N_14556,N_9686,N_8184);
or U14557 (N_14557,N_10736,N_8457);
and U14558 (N_14558,N_8545,N_8299);
and U14559 (N_14559,N_9471,N_8049);
nand U14560 (N_14560,N_8503,N_9668);
or U14561 (N_14561,N_11970,N_8467);
nand U14562 (N_14562,N_9780,N_10389);
nor U14563 (N_14563,N_11912,N_8367);
nor U14564 (N_14564,N_9632,N_8726);
nor U14565 (N_14565,N_8424,N_8609);
nand U14566 (N_14566,N_9334,N_11988);
xor U14567 (N_14567,N_8519,N_9655);
and U14568 (N_14568,N_9918,N_9493);
nor U14569 (N_14569,N_8031,N_10908);
and U14570 (N_14570,N_10866,N_8400);
nand U14571 (N_14571,N_11832,N_10826);
nor U14572 (N_14572,N_10941,N_10747);
nand U14573 (N_14573,N_9581,N_9990);
or U14574 (N_14574,N_9221,N_10585);
nand U14575 (N_14575,N_10048,N_10981);
xor U14576 (N_14576,N_9745,N_8760);
nand U14577 (N_14577,N_10477,N_11426);
or U14578 (N_14578,N_11797,N_11580);
or U14579 (N_14579,N_10339,N_10251);
nand U14580 (N_14580,N_9225,N_10976);
or U14581 (N_14581,N_9552,N_10456);
or U14582 (N_14582,N_8108,N_11504);
nand U14583 (N_14583,N_8156,N_9460);
nor U14584 (N_14584,N_9351,N_8663);
and U14585 (N_14585,N_8236,N_11920);
and U14586 (N_14586,N_8815,N_9736);
xor U14587 (N_14587,N_11064,N_10536);
and U14588 (N_14588,N_11703,N_11833);
and U14589 (N_14589,N_11740,N_10480);
or U14590 (N_14590,N_9967,N_10019);
nor U14591 (N_14591,N_9630,N_9389);
and U14592 (N_14592,N_8591,N_11285);
nand U14593 (N_14593,N_8827,N_9322);
nor U14594 (N_14594,N_8883,N_10482);
nand U14595 (N_14595,N_10071,N_9730);
xor U14596 (N_14596,N_9056,N_8406);
or U14597 (N_14597,N_9437,N_11386);
nor U14598 (N_14598,N_9541,N_9183);
nor U14599 (N_14599,N_9423,N_10761);
xnor U14600 (N_14600,N_9611,N_9617);
nor U14601 (N_14601,N_11502,N_10575);
nor U14602 (N_14602,N_11059,N_10985);
or U14603 (N_14603,N_10673,N_9894);
and U14604 (N_14604,N_11823,N_9070);
nor U14605 (N_14605,N_10475,N_9076);
xnor U14606 (N_14606,N_11754,N_8862);
nor U14607 (N_14607,N_9653,N_11949);
nand U14608 (N_14608,N_8036,N_8471);
and U14609 (N_14609,N_9705,N_8547);
or U14610 (N_14610,N_9267,N_10888);
xor U14611 (N_14611,N_10515,N_10653);
and U14612 (N_14612,N_10101,N_8457);
nand U14613 (N_14613,N_8961,N_8334);
nor U14614 (N_14614,N_10524,N_11382);
nor U14615 (N_14615,N_8691,N_8248);
xnor U14616 (N_14616,N_8353,N_9936);
or U14617 (N_14617,N_11975,N_9536);
nand U14618 (N_14618,N_10735,N_11864);
and U14619 (N_14619,N_9223,N_10443);
nor U14620 (N_14620,N_8861,N_8962);
nor U14621 (N_14621,N_11748,N_8408);
nand U14622 (N_14622,N_11266,N_10390);
nand U14623 (N_14623,N_8640,N_8993);
or U14624 (N_14624,N_11625,N_9506);
and U14625 (N_14625,N_11236,N_11660);
or U14626 (N_14626,N_11804,N_10096);
and U14627 (N_14627,N_11906,N_11031);
or U14628 (N_14628,N_9555,N_8142);
xnor U14629 (N_14629,N_11500,N_9404);
nor U14630 (N_14630,N_9303,N_8285);
nor U14631 (N_14631,N_10695,N_10339);
and U14632 (N_14632,N_11250,N_11061);
nand U14633 (N_14633,N_11128,N_11631);
nor U14634 (N_14634,N_8804,N_8312);
nand U14635 (N_14635,N_10633,N_8329);
xnor U14636 (N_14636,N_10462,N_11580);
nor U14637 (N_14637,N_9294,N_9464);
nor U14638 (N_14638,N_10884,N_8857);
and U14639 (N_14639,N_8555,N_9613);
nand U14640 (N_14640,N_9104,N_11347);
or U14641 (N_14641,N_11536,N_11613);
and U14642 (N_14642,N_8905,N_8412);
and U14643 (N_14643,N_8038,N_9612);
or U14644 (N_14644,N_11394,N_9429);
xor U14645 (N_14645,N_8926,N_10646);
nor U14646 (N_14646,N_9215,N_10599);
nor U14647 (N_14647,N_10770,N_8080);
xor U14648 (N_14648,N_8449,N_8633);
nor U14649 (N_14649,N_9144,N_9310);
xnor U14650 (N_14650,N_8280,N_11678);
and U14651 (N_14651,N_9023,N_8658);
xor U14652 (N_14652,N_8311,N_8604);
and U14653 (N_14653,N_8619,N_9787);
and U14654 (N_14654,N_10620,N_11673);
or U14655 (N_14655,N_11543,N_10342);
and U14656 (N_14656,N_11106,N_9354);
and U14657 (N_14657,N_9634,N_10663);
xor U14658 (N_14658,N_8441,N_11540);
or U14659 (N_14659,N_10965,N_8059);
and U14660 (N_14660,N_8119,N_11624);
and U14661 (N_14661,N_9471,N_8926);
nand U14662 (N_14662,N_9432,N_11757);
nor U14663 (N_14663,N_10867,N_9834);
or U14664 (N_14664,N_10879,N_10656);
nor U14665 (N_14665,N_11918,N_9603);
or U14666 (N_14666,N_8646,N_8022);
nor U14667 (N_14667,N_11064,N_8431);
and U14668 (N_14668,N_11028,N_9235);
nand U14669 (N_14669,N_11574,N_10919);
or U14670 (N_14670,N_8121,N_10613);
xor U14671 (N_14671,N_9220,N_11512);
nor U14672 (N_14672,N_8600,N_10418);
or U14673 (N_14673,N_9030,N_8097);
nor U14674 (N_14674,N_9453,N_9236);
and U14675 (N_14675,N_9210,N_11785);
or U14676 (N_14676,N_9992,N_10980);
nand U14677 (N_14677,N_10944,N_8993);
or U14678 (N_14678,N_8891,N_9727);
xnor U14679 (N_14679,N_9282,N_8766);
and U14680 (N_14680,N_8180,N_9266);
and U14681 (N_14681,N_11937,N_10909);
and U14682 (N_14682,N_10722,N_8682);
nor U14683 (N_14683,N_8021,N_8447);
nor U14684 (N_14684,N_8004,N_8479);
or U14685 (N_14685,N_11673,N_11649);
nand U14686 (N_14686,N_9541,N_10938);
nor U14687 (N_14687,N_9310,N_11502);
and U14688 (N_14688,N_10661,N_11967);
or U14689 (N_14689,N_11653,N_8850);
and U14690 (N_14690,N_10090,N_8795);
or U14691 (N_14691,N_11066,N_9125);
nor U14692 (N_14692,N_11459,N_8434);
or U14693 (N_14693,N_10362,N_8976);
and U14694 (N_14694,N_9274,N_11423);
and U14695 (N_14695,N_8740,N_9024);
and U14696 (N_14696,N_9500,N_10871);
and U14697 (N_14697,N_10545,N_11490);
nor U14698 (N_14698,N_8235,N_10677);
nand U14699 (N_14699,N_11382,N_11256);
or U14700 (N_14700,N_10905,N_8785);
nor U14701 (N_14701,N_10704,N_8880);
and U14702 (N_14702,N_10992,N_9598);
nor U14703 (N_14703,N_10199,N_9283);
or U14704 (N_14704,N_8965,N_10225);
xnor U14705 (N_14705,N_11284,N_9148);
and U14706 (N_14706,N_10525,N_11127);
xor U14707 (N_14707,N_11931,N_10191);
nand U14708 (N_14708,N_8478,N_10324);
nor U14709 (N_14709,N_10660,N_9185);
nor U14710 (N_14710,N_11547,N_11446);
xor U14711 (N_14711,N_8488,N_10463);
and U14712 (N_14712,N_10337,N_11612);
and U14713 (N_14713,N_10611,N_10955);
and U14714 (N_14714,N_8307,N_11159);
or U14715 (N_14715,N_10164,N_11109);
or U14716 (N_14716,N_8291,N_10214);
nor U14717 (N_14717,N_11083,N_8113);
and U14718 (N_14718,N_10128,N_8880);
nor U14719 (N_14719,N_9962,N_8652);
nor U14720 (N_14720,N_9698,N_8689);
or U14721 (N_14721,N_10910,N_8577);
or U14722 (N_14722,N_11389,N_10879);
and U14723 (N_14723,N_11139,N_9265);
and U14724 (N_14724,N_8874,N_10123);
or U14725 (N_14725,N_9297,N_10383);
nand U14726 (N_14726,N_10617,N_9552);
nor U14727 (N_14727,N_11657,N_11170);
or U14728 (N_14728,N_11258,N_8799);
nand U14729 (N_14729,N_9799,N_8751);
nand U14730 (N_14730,N_9587,N_10529);
nor U14731 (N_14731,N_10713,N_10160);
nor U14732 (N_14732,N_10756,N_11390);
xor U14733 (N_14733,N_10408,N_8943);
and U14734 (N_14734,N_10258,N_8895);
xor U14735 (N_14735,N_9103,N_11259);
and U14736 (N_14736,N_11952,N_11440);
nand U14737 (N_14737,N_9733,N_11665);
nand U14738 (N_14738,N_11775,N_9605);
and U14739 (N_14739,N_10061,N_9258);
or U14740 (N_14740,N_8993,N_9068);
or U14741 (N_14741,N_8548,N_11634);
or U14742 (N_14742,N_10717,N_8224);
and U14743 (N_14743,N_9693,N_8664);
xnor U14744 (N_14744,N_11984,N_9526);
xnor U14745 (N_14745,N_8720,N_11445);
nor U14746 (N_14746,N_9179,N_9793);
nand U14747 (N_14747,N_11454,N_9784);
nand U14748 (N_14748,N_8516,N_11997);
or U14749 (N_14749,N_10438,N_8289);
nor U14750 (N_14750,N_9017,N_8110);
and U14751 (N_14751,N_8996,N_11844);
nand U14752 (N_14752,N_8959,N_10126);
and U14753 (N_14753,N_11565,N_11836);
and U14754 (N_14754,N_10679,N_10994);
nor U14755 (N_14755,N_9391,N_9225);
or U14756 (N_14756,N_11696,N_11080);
xnor U14757 (N_14757,N_9174,N_8091);
and U14758 (N_14758,N_10655,N_8065);
or U14759 (N_14759,N_8234,N_9234);
or U14760 (N_14760,N_11041,N_10434);
nor U14761 (N_14761,N_9841,N_10279);
nand U14762 (N_14762,N_11190,N_8564);
and U14763 (N_14763,N_11854,N_8421);
nand U14764 (N_14764,N_9947,N_11630);
nand U14765 (N_14765,N_9347,N_10170);
and U14766 (N_14766,N_9316,N_9638);
or U14767 (N_14767,N_8037,N_8204);
nor U14768 (N_14768,N_10322,N_9374);
or U14769 (N_14769,N_8563,N_9762);
and U14770 (N_14770,N_11433,N_9204);
nand U14771 (N_14771,N_8285,N_11717);
nor U14772 (N_14772,N_11558,N_11230);
nor U14773 (N_14773,N_10415,N_10807);
nor U14774 (N_14774,N_9574,N_10443);
nor U14775 (N_14775,N_11603,N_11834);
or U14776 (N_14776,N_9261,N_8635);
nand U14777 (N_14777,N_9621,N_10410);
or U14778 (N_14778,N_8973,N_9086);
xnor U14779 (N_14779,N_9313,N_8723);
xnor U14780 (N_14780,N_8272,N_10001);
xnor U14781 (N_14781,N_11369,N_9670);
or U14782 (N_14782,N_8321,N_9425);
nand U14783 (N_14783,N_8833,N_11691);
or U14784 (N_14784,N_8109,N_11123);
or U14785 (N_14785,N_11121,N_8333);
nor U14786 (N_14786,N_10519,N_10514);
and U14787 (N_14787,N_9936,N_9150);
xor U14788 (N_14788,N_8713,N_10323);
nor U14789 (N_14789,N_11411,N_8976);
or U14790 (N_14790,N_8022,N_8822);
or U14791 (N_14791,N_11076,N_11044);
nand U14792 (N_14792,N_8567,N_11831);
or U14793 (N_14793,N_8854,N_8282);
xor U14794 (N_14794,N_9844,N_9228);
or U14795 (N_14795,N_9835,N_11093);
or U14796 (N_14796,N_9855,N_9132);
and U14797 (N_14797,N_8608,N_9395);
or U14798 (N_14798,N_8857,N_10208);
nand U14799 (N_14799,N_10510,N_9383);
and U14800 (N_14800,N_9307,N_10578);
nor U14801 (N_14801,N_8222,N_8139);
nor U14802 (N_14802,N_9256,N_11617);
and U14803 (N_14803,N_8863,N_11955);
xnor U14804 (N_14804,N_10987,N_10887);
and U14805 (N_14805,N_8965,N_11550);
nand U14806 (N_14806,N_11768,N_10539);
and U14807 (N_14807,N_9986,N_11462);
nor U14808 (N_14808,N_10800,N_10935);
and U14809 (N_14809,N_9888,N_8507);
or U14810 (N_14810,N_10166,N_10022);
nand U14811 (N_14811,N_10219,N_8496);
nor U14812 (N_14812,N_10507,N_9321);
and U14813 (N_14813,N_8632,N_10531);
xnor U14814 (N_14814,N_10967,N_10571);
nand U14815 (N_14815,N_9321,N_10660);
or U14816 (N_14816,N_8506,N_8141);
nand U14817 (N_14817,N_9861,N_8638);
nor U14818 (N_14818,N_9789,N_10493);
nor U14819 (N_14819,N_8445,N_10811);
or U14820 (N_14820,N_11957,N_10508);
and U14821 (N_14821,N_11555,N_11928);
and U14822 (N_14822,N_11926,N_11422);
nand U14823 (N_14823,N_8695,N_10738);
and U14824 (N_14824,N_11501,N_8626);
nor U14825 (N_14825,N_9564,N_11648);
or U14826 (N_14826,N_10946,N_8614);
nand U14827 (N_14827,N_9338,N_10147);
or U14828 (N_14828,N_11719,N_9780);
nand U14829 (N_14829,N_10506,N_8300);
and U14830 (N_14830,N_10428,N_8387);
nand U14831 (N_14831,N_9519,N_9954);
or U14832 (N_14832,N_9315,N_9997);
or U14833 (N_14833,N_10835,N_11738);
and U14834 (N_14834,N_11599,N_10314);
and U14835 (N_14835,N_10250,N_11868);
or U14836 (N_14836,N_11244,N_10828);
or U14837 (N_14837,N_11602,N_8635);
nor U14838 (N_14838,N_10861,N_11747);
or U14839 (N_14839,N_8561,N_11730);
or U14840 (N_14840,N_11193,N_10413);
nand U14841 (N_14841,N_9222,N_8029);
nor U14842 (N_14842,N_10722,N_8613);
nor U14843 (N_14843,N_8861,N_8944);
or U14844 (N_14844,N_9361,N_11484);
nor U14845 (N_14845,N_10094,N_8498);
and U14846 (N_14846,N_10897,N_11254);
and U14847 (N_14847,N_9417,N_11733);
and U14848 (N_14848,N_10355,N_8305);
or U14849 (N_14849,N_9751,N_10704);
or U14850 (N_14850,N_9628,N_9073);
and U14851 (N_14851,N_11604,N_8919);
or U14852 (N_14852,N_10017,N_10864);
or U14853 (N_14853,N_11275,N_10804);
nor U14854 (N_14854,N_8068,N_8719);
nor U14855 (N_14855,N_11415,N_10036);
nand U14856 (N_14856,N_11894,N_8627);
nand U14857 (N_14857,N_10638,N_11582);
nand U14858 (N_14858,N_10044,N_11238);
and U14859 (N_14859,N_10303,N_11596);
or U14860 (N_14860,N_8980,N_10040);
xnor U14861 (N_14861,N_10319,N_10501);
nand U14862 (N_14862,N_8370,N_8872);
nand U14863 (N_14863,N_10430,N_8945);
xor U14864 (N_14864,N_8249,N_9956);
and U14865 (N_14865,N_11358,N_8209);
and U14866 (N_14866,N_8611,N_8891);
nor U14867 (N_14867,N_9653,N_8798);
and U14868 (N_14868,N_9883,N_8784);
nor U14869 (N_14869,N_9903,N_11159);
or U14870 (N_14870,N_10500,N_8668);
nor U14871 (N_14871,N_11772,N_10787);
xnor U14872 (N_14872,N_11640,N_11775);
nor U14873 (N_14873,N_8609,N_9148);
xor U14874 (N_14874,N_11850,N_9407);
and U14875 (N_14875,N_10098,N_11226);
nor U14876 (N_14876,N_10020,N_10595);
nand U14877 (N_14877,N_11357,N_8478);
nor U14878 (N_14878,N_10297,N_9894);
or U14879 (N_14879,N_10044,N_8561);
and U14880 (N_14880,N_9719,N_10491);
xor U14881 (N_14881,N_10667,N_10577);
or U14882 (N_14882,N_10291,N_9820);
nand U14883 (N_14883,N_10621,N_11277);
or U14884 (N_14884,N_10804,N_9777);
or U14885 (N_14885,N_8777,N_9376);
nor U14886 (N_14886,N_10750,N_10352);
or U14887 (N_14887,N_9959,N_11534);
nor U14888 (N_14888,N_9404,N_10151);
nand U14889 (N_14889,N_11852,N_9674);
nand U14890 (N_14890,N_11597,N_8873);
and U14891 (N_14891,N_8376,N_8063);
nor U14892 (N_14892,N_11539,N_9570);
xnor U14893 (N_14893,N_9659,N_8763);
nand U14894 (N_14894,N_9286,N_8448);
or U14895 (N_14895,N_9963,N_8829);
nand U14896 (N_14896,N_10404,N_11238);
and U14897 (N_14897,N_8494,N_10488);
nand U14898 (N_14898,N_11125,N_8947);
or U14899 (N_14899,N_9518,N_9016);
nor U14900 (N_14900,N_8717,N_9298);
xor U14901 (N_14901,N_11991,N_10787);
nor U14902 (N_14902,N_10751,N_8681);
and U14903 (N_14903,N_10707,N_8297);
or U14904 (N_14904,N_9482,N_9377);
or U14905 (N_14905,N_11288,N_11559);
nor U14906 (N_14906,N_11846,N_9922);
nor U14907 (N_14907,N_8355,N_10239);
xor U14908 (N_14908,N_8649,N_10714);
or U14909 (N_14909,N_10585,N_9844);
and U14910 (N_14910,N_9176,N_8741);
and U14911 (N_14911,N_8260,N_8747);
nand U14912 (N_14912,N_10011,N_8714);
xnor U14913 (N_14913,N_9987,N_10697);
nand U14914 (N_14914,N_8519,N_10732);
nor U14915 (N_14915,N_8378,N_10616);
and U14916 (N_14916,N_11394,N_9405);
nand U14917 (N_14917,N_11979,N_10939);
nor U14918 (N_14918,N_11220,N_10687);
and U14919 (N_14919,N_9187,N_10285);
nor U14920 (N_14920,N_10402,N_8717);
nor U14921 (N_14921,N_9687,N_8155);
and U14922 (N_14922,N_8380,N_10165);
nand U14923 (N_14923,N_11557,N_11770);
and U14924 (N_14924,N_11954,N_11289);
or U14925 (N_14925,N_11593,N_9030);
nor U14926 (N_14926,N_10535,N_9163);
nor U14927 (N_14927,N_9849,N_8280);
or U14928 (N_14928,N_9778,N_10652);
or U14929 (N_14929,N_8896,N_9480);
and U14930 (N_14930,N_9776,N_9307);
nand U14931 (N_14931,N_8559,N_9375);
and U14932 (N_14932,N_10229,N_9486);
nand U14933 (N_14933,N_11575,N_9942);
nor U14934 (N_14934,N_8597,N_11759);
nor U14935 (N_14935,N_9062,N_8953);
nor U14936 (N_14936,N_9558,N_11890);
nor U14937 (N_14937,N_8560,N_8029);
xnor U14938 (N_14938,N_11842,N_9376);
nand U14939 (N_14939,N_8436,N_11078);
nor U14940 (N_14940,N_9552,N_8450);
or U14941 (N_14941,N_8751,N_11710);
nor U14942 (N_14942,N_10817,N_10266);
nand U14943 (N_14943,N_8520,N_9499);
nand U14944 (N_14944,N_8586,N_9649);
and U14945 (N_14945,N_10639,N_11785);
nor U14946 (N_14946,N_11458,N_8583);
nor U14947 (N_14947,N_11626,N_8139);
or U14948 (N_14948,N_10523,N_9823);
or U14949 (N_14949,N_11929,N_8290);
nor U14950 (N_14950,N_8519,N_10821);
or U14951 (N_14951,N_8774,N_11251);
nand U14952 (N_14952,N_9926,N_10522);
nor U14953 (N_14953,N_9944,N_10847);
nor U14954 (N_14954,N_9172,N_10198);
nand U14955 (N_14955,N_11771,N_9655);
nor U14956 (N_14956,N_10424,N_9985);
and U14957 (N_14957,N_8160,N_8081);
nand U14958 (N_14958,N_8148,N_10515);
and U14959 (N_14959,N_10440,N_11577);
or U14960 (N_14960,N_11875,N_9760);
xor U14961 (N_14961,N_10385,N_8631);
nand U14962 (N_14962,N_8515,N_9697);
or U14963 (N_14963,N_11314,N_9724);
and U14964 (N_14964,N_10892,N_10005);
nor U14965 (N_14965,N_11929,N_8911);
nor U14966 (N_14966,N_8612,N_11487);
nor U14967 (N_14967,N_11849,N_8017);
xnor U14968 (N_14968,N_9544,N_9002);
and U14969 (N_14969,N_9427,N_9661);
xor U14970 (N_14970,N_9625,N_8550);
and U14971 (N_14971,N_9335,N_11788);
and U14972 (N_14972,N_10709,N_10082);
nand U14973 (N_14973,N_11587,N_9802);
nand U14974 (N_14974,N_8547,N_8049);
nor U14975 (N_14975,N_11413,N_10836);
xor U14976 (N_14976,N_9352,N_8579);
and U14977 (N_14977,N_9528,N_10464);
nor U14978 (N_14978,N_9979,N_9386);
xnor U14979 (N_14979,N_9020,N_8072);
xnor U14980 (N_14980,N_8506,N_11959);
and U14981 (N_14981,N_10230,N_11431);
or U14982 (N_14982,N_11396,N_10802);
and U14983 (N_14983,N_9233,N_8372);
nor U14984 (N_14984,N_9724,N_9250);
nor U14985 (N_14985,N_9979,N_8581);
xnor U14986 (N_14986,N_10564,N_8841);
nand U14987 (N_14987,N_10371,N_9142);
nor U14988 (N_14988,N_8006,N_9371);
xnor U14989 (N_14989,N_11556,N_11006);
xor U14990 (N_14990,N_8200,N_8207);
and U14991 (N_14991,N_10401,N_10056);
or U14992 (N_14992,N_10959,N_10636);
and U14993 (N_14993,N_9147,N_9862);
nor U14994 (N_14994,N_11901,N_8020);
nor U14995 (N_14995,N_8746,N_9085);
or U14996 (N_14996,N_9638,N_10444);
or U14997 (N_14997,N_9507,N_10441);
and U14998 (N_14998,N_9398,N_8841);
nor U14999 (N_14999,N_9959,N_9056);
and U15000 (N_15000,N_8555,N_8678);
or U15001 (N_15001,N_10338,N_11971);
nor U15002 (N_15002,N_11138,N_8034);
xor U15003 (N_15003,N_11705,N_10994);
and U15004 (N_15004,N_10329,N_9371);
nand U15005 (N_15005,N_10792,N_8804);
or U15006 (N_15006,N_9096,N_11449);
or U15007 (N_15007,N_11216,N_10440);
nor U15008 (N_15008,N_8962,N_11487);
nor U15009 (N_15009,N_8853,N_10436);
or U15010 (N_15010,N_8404,N_11156);
nor U15011 (N_15011,N_11947,N_8159);
nand U15012 (N_15012,N_11726,N_10835);
or U15013 (N_15013,N_8399,N_10230);
nand U15014 (N_15014,N_11458,N_8516);
or U15015 (N_15015,N_11039,N_10744);
and U15016 (N_15016,N_9309,N_10839);
nand U15017 (N_15017,N_11767,N_8757);
nor U15018 (N_15018,N_8095,N_10883);
nand U15019 (N_15019,N_9693,N_10858);
nand U15020 (N_15020,N_11473,N_9407);
nor U15021 (N_15021,N_11438,N_8064);
and U15022 (N_15022,N_11623,N_11977);
or U15023 (N_15023,N_10146,N_11897);
or U15024 (N_15024,N_8978,N_11866);
nor U15025 (N_15025,N_10394,N_8748);
or U15026 (N_15026,N_8598,N_10061);
or U15027 (N_15027,N_8863,N_11124);
xor U15028 (N_15028,N_9560,N_8181);
nor U15029 (N_15029,N_9526,N_8751);
xnor U15030 (N_15030,N_10757,N_9459);
xnor U15031 (N_15031,N_11355,N_11226);
or U15032 (N_15032,N_11304,N_11585);
or U15033 (N_15033,N_11474,N_10226);
and U15034 (N_15034,N_10637,N_9853);
and U15035 (N_15035,N_10103,N_10876);
nor U15036 (N_15036,N_9700,N_9409);
or U15037 (N_15037,N_9593,N_10488);
nor U15038 (N_15038,N_8128,N_11572);
or U15039 (N_15039,N_10391,N_11570);
nor U15040 (N_15040,N_10924,N_10176);
nor U15041 (N_15041,N_9874,N_10659);
nand U15042 (N_15042,N_10306,N_11067);
or U15043 (N_15043,N_9298,N_9384);
nand U15044 (N_15044,N_10370,N_8133);
nand U15045 (N_15045,N_9815,N_9065);
or U15046 (N_15046,N_11597,N_8632);
nand U15047 (N_15047,N_10072,N_9045);
and U15048 (N_15048,N_10622,N_9208);
or U15049 (N_15049,N_8698,N_8240);
or U15050 (N_15050,N_8967,N_9121);
nand U15051 (N_15051,N_10878,N_10164);
or U15052 (N_15052,N_11562,N_11298);
or U15053 (N_15053,N_9078,N_9316);
nand U15054 (N_15054,N_11501,N_10006);
nand U15055 (N_15055,N_9918,N_9504);
nand U15056 (N_15056,N_11509,N_11459);
nor U15057 (N_15057,N_9114,N_8163);
or U15058 (N_15058,N_10676,N_11234);
or U15059 (N_15059,N_10298,N_10970);
nand U15060 (N_15060,N_9038,N_9799);
or U15061 (N_15061,N_11207,N_8515);
or U15062 (N_15062,N_9434,N_8270);
xnor U15063 (N_15063,N_9666,N_9882);
or U15064 (N_15064,N_9308,N_8409);
nor U15065 (N_15065,N_10980,N_8081);
or U15066 (N_15066,N_9488,N_9671);
or U15067 (N_15067,N_10776,N_11991);
xnor U15068 (N_15068,N_8267,N_8701);
and U15069 (N_15069,N_10290,N_9422);
nand U15070 (N_15070,N_11966,N_11391);
nand U15071 (N_15071,N_8664,N_11222);
xor U15072 (N_15072,N_8201,N_8215);
nor U15073 (N_15073,N_9759,N_9826);
or U15074 (N_15074,N_10846,N_8068);
or U15075 (N_15075,N_8857,N_10817);
nor U15076 (N_15076,N_10766,N_8889);
or U15077 (N_15077,N_8452,N_10439);
or U15078 (N_15078,N_9010,N_10375);
nand U15079 (N_15079,N_11089,N_9225);
nor U15080 (N_15080,N_8134,N_8836);
xor U15081 (N_15081,N_10602,N_8331);
nor U15082 (N_15082,N_10041,N_11258);
nand U15083 (N_15083,N_9125,N_8763);
nand U15084 (N_15084,N_11476,N_8471);
nor U15085 (N_15085,N_10437,N_9578);
or U15086 (N_15086,N_10556,N_10946);
nand U15087 (N_15087,N_8568,N_9560);
and U15088 (N_15088,N_9099,N_11643);
and U15089 (N_15089,N_10105,N_9589);
and U15090 (N_15090,N_9402,N_9161);
nand U15091 (N_15091,N_9532,N_10084);
or U15092 (N_15092,N_8648,N_8171);
and U15093 (N_15093,N_8852,N_9799);
nor U15094 (N_15094,N_8620,N_10725);
or U15095 (N_15095,N_9769,N_9821);
nand U15096 (N_15096,N_11155,N_10404);
nand U15097 (N_15097,N_9965,N_8507);
nand U15098 (N_15098,N_11028,N_11870);
nor U15099 (N_15099,N_10813,N_11248);
and U15100 (N_15100,N_11447,N_10161);
xor U15101 (N_15101,N_11237,N_11102);
and U15102 (N_15102,N_11403,N_8203);
or U15103 (N_15103,N_9235,N_9817);
nand U15104 (N_15104,N_10668,N_10117);
nand U15105 (N_15105,N_10093,N_10523);
nand U15106 (N_15106,N_10020,N_11226);
nand U15107 (N_15107,N_11938,N_11943);
or U15108 (N_15108,N_11781,N_11737);
or U15109 (N_15109,N_8045,N_10545);
xor U15110 (N_15110,N_10819,N_9828);
and U15111 (N_15111,N_9112,N_11302);
nor U15112 (N_15112,N_9059,N_9223);
nand U15113 (N_15113,N_11912,N_8047);
nor U15114 (N_15114,N_9038,N_10022);
and U15115 (N_15115,N_11119,N_10028);
nor U15116 (N_15116,N_11609,N_10985);
nand U15117 (N_15117,N_8434,N_11073);
nor U15118 (N_15118,N_11799,N_11380);
nor U15119 (N_15119,N_11931,N_8544);
and U15120 (N_15120,N_10400,N_10017);
or U15121 (N_15121,N_9816,N_10132);
nand U15122 (N_15122,N_8922,N_9903);
nor U15123 (N_15123,N_8540,N_9829);
xnor U15124 (N_15124,N_10313,N_8570);
xor U15125 (N_15125,N_10234,N_9516);
xnor U15126 (N_15126,N_8847,N_10691);
nand U15127 (N_15127,N_11840,N_10339);
xor U15128 (N_15128,N_11700,N_8395);
and U15129 (N_15129,N_8854,N_9633);
and U15130 (N_15130,N_11104,N_10188);
xor U15131 (N_15131,N_8460,N_10659);
nand U15132 (N_15132,N_9204,N_10902);
nand U15133 (N_15133,N_8948,N_9737);
and U15134 (N_15134,N_9414,N_10164);
nand U15135 (N_15135,N_11567,N_11124);
or U15136 (N_15136,N_8834,N_8492);
nor U15137 (N_15137,N_9857,N_8671);
and U15138 (N_15138,N_9929,N_10990);
nand U15139 (N_15139,N_11359,N_11319);
nor U15140 (N_15140,N_11432,N_10671);
and U15141 (N_15141,N_11953,N_10501);
and U15142 (N_15142,N_10647,N_8133);
nand U15143 (N_15143,N_8691,N_9162);
and U15144 (N_15144,N_10850,N_11563);
or U15145 (N_15145,N_9477,N_9385);
or U15146 (N_15146,N_8407,N_10599);
xnor U15147 (N_15147,N_10081,N_10489);
nand U15148 (N_15148,N_10579,N_11118);
nor U15149 (N_15149,N_9959,N_10094);
nor U15150 (N_15150,N_9102,N_8445);
and U15151 (N_15151,N_11995,N_10202);
xor U15152 (N_15152,N_11391,N_11557);
nand U15153 (N_15153,N_9364,N_9295);
and U15154 (N_15154,N_8541,N_8781);
nand U15155 (N_15155,N_9786,N_8490);
xnor U15156 (N_15156,N_9051,N_11817);
nor U15157 (N_15157,N_10572,N_11747);
or U15158 (N_15158,N_9212,N_10813);
and U15159 (N_15159,N_10782,N_9416);
or U15160 (N_15160,N_11733,N_8239);
nor U15161 (N_15161,N_9473,N_10517);
nand U15162 (N_15162,N_11921,N_8335);
nor U15163 (N_15163,N_8610,N_10443);
nand U15164 (N_15164,N_10232,N_9450);
nand U15165 (N_15165,N_11035,N_10765);
nand U15166 (N_15166,N_8445,N_9208);
nor U15167 (N_15167,N_11862,N_11212);
xnor U15168 (N_15168,N_9719,N_9032);
and U15169 (N_15169,N_9964,N_9204);
or U15170 (N_15170,N_8638,N_8143);
nand U15171 (N_15171,N_11520,N_11561);
xnor U15172 (N_15172,N_10655,N_8207);
or U15173 (N_15173,N_10141,N_8345);
and U15174 (N_15174,N_9851,N_8536);
nand U15175 (N_15175,N_11722,N_9773);
or U15176 (N_15176,N_11562,N_10498);
or U15177 (N_15177,N_8719,N_10077);
nor U15178 (N_15178,N_8617,N_8870);
nand U15179 (N_15179,N_11456,N_8681);
nor U15180 (N_15180,N_11742,N_10807);
nor U15181 (N_15181,N_8190,N_10000);
nor U15182 (N_15182,N_10204,N_10208);
xor U15183 (N_15183,N_11365,N_11992);
xor U15184 (N_15184,N_10600,N_11326);
nand U15185 (N_15185,N_10178,N_11409);
and U15186 (N_15186,N_9241,N_10290);
nand U15187 (N_15187,N_10648,N_9643);
nor U15188 (N_15188,N_11709,N_8543);
and U15189 (N_15189,N_8840,N_10913);
nand U15190 (N_15190,N_9798,N_9907);
nor U15191 (N_15191,N_9081,N_10201);
nor U15192 (N_15192,N_8603,N_8014);
or U15193 (N_15193,N_8030,N_9990);
or U15194 (N_15194,N_11077,N_10607);
nand U15195 (N_15195,N_9331,N_11973);
and U15196 (N_15196,N_8624,N_9403);
and U15197 (N_15197,N_9609,N_8113);
nor U15198 (N_15198,N_10807,N_10079);
nor U15199 (N_15199,N_11203,N_10076);
nor U15200 (N_15200,N_8700,N_9955);
or U15201 (N_15201,N_9763,N_11976);
xor U15202 (N_15202,N_11026,N_10367);
nor U15203 (N_15203,N_10362,N_9694);
or U15204 (N_15204,N_9545,N_8622);
nand U15205 (N_15205,N_11817,N_8180);
nand U15206 (N_15206,N_10528,N_8752);
or U15207 (N_15207,N_9288,N_11205);
or U15208 (N_15208,N_9727,N_9744);
nor U15209 (N_15209,N_10297,N_11463);
nand U15210 (N_15210,N_9099,N_9675);
and U15211 (N_15211,N_9970,N_10797);
xor U15212 (N_15212,N_8431,N_9756);
nand U15213 (N_15213,N_9593,N_9014);
nor U15214 (N_15214,N_10920,N_11110);
or U15215 (N_15215,N_8931,N_9730);
nand U15216 (N_15216,N_9097,N_10722);
nand U15217 (N_15217,N_9601,N_10698);
nand U15218 (N_15218,N_11580,N_9959);
or U15219 (N_15219,N_11035,N_10044);
nor U15220 (N_15220,N_8232,N_10227);
nand U15221 (N_15221,N_9160,N_8482);
or U15222 (N_15222,N_8253,N_9796);
xor U15223 (N_15223,N_9050,N_11013);
nand U15224 (N_15224,N_8144,N_8836);
xor U15225 (N_15225,N_8392,N_10092);
and U15226 (N_15226,N_10175,N_8352);
nand U15227 (N_15227,N_9513,N_9985);
and U15228 (N_15228,N_11254,N_8184);
nor U15229 (N_15229,N_11117,N_10739);
nor U15230 (N_15230,N_8238,N_9810);
nor U15231 (N_15231,N_10320,N_11412);
nor U15232 (N_15232,N_11620,N_8578);
nand U15233 (N_15233,N_10766,N_11586);
and U15234 (N_15234,N_9372,N_8566);
nand U15235 (N_15235,N_10587,N_8390);
or U15236 (N_15236,N_10004,N_9593);
nor U15237 (N_15237,N_11668,N_8896);
or U15238 (N_15238,N_10828,N_10871);
or U15239 (N_15239,N_11381,N_11356);
nor U15240 (N_15240,N_10919,N_9350);
or U15241 (N_15241,N_10916,N_10172);
nand U15242 (N_15242,N_9514,N_10141);
or U15243 (N_15243,N_8236,N_8930);
and U15244 (N_15244,N_11450,N_11255);
and U15245 (N_15245,N_10890,N_8914);
xor U15246 (N_15246,N_8969,N_11072);
nor U15247 (N_15247,N_9374,N_8930);
xnor U15248 (N_15248,N_11619,N_11798);
nor U15249 (N_15249,N_11272,N_9093);
nor U15250 (N_15250,N_9831,N_9197);
or U15251 (N_15251,N_11285,N_11108);
nor U15252 (N_15252,N_9844,N_11871);
and U15253 (N_15253,N_9240,N_11245);
or U15254 (N_15254,N_9593,N_9967);
and U15255 (N_15255,N_8680,N_9280);
xor U15256 (N_15256,N_11952,N_11116);
xnor U15257 (N_15257,N_11551,N_9013);
and U15258 (N_15258,N_10299,N_9956);
xor U15259 (N_15259,N_11752,N_10690);
xnor U15260 (N_15260,N_9602,N_8102);
and U15261 (N_15261,N_10108,N_11111);
nand U15262 (N_15262,N_10295,N_11082);
xor U15263 (N_15263,N_9784,N_10785);
nand U15264 (N_15264,N_9298,N_11392);
nor U15265 (N_15265,N_11048,N_9263);
nor U15266 (N_15266,N_9914,N_8384);
xnor U15267 (N_15267,N_11530,N_10247);
nor U15268 (N_15268,N_9183,N_11306);
or U15269 (N_15269,N_8940,N_11180);
and U15270 (N_15270,N_10213,N_9766);
nand U15271 (N_15271,N_10955,N_9198);
nand U15272 (N_15272,N_11125,N_8544);
and U15273 (N_15273,N_9563,N_10457);
nor U15274 (N_15274,N_11052,N_10220);
or U15275 (N_15275,N_10568,N_9494);
and U15276 (N_15276,N_10280,N_8565);
nor U15277 (N_15277,N_8117,N_8214);
nand U15278 (N_15278,N_10135,N_11110);
nor U15279 (N_15279,N_10122,N_8750);
and U15280 (N_15280,N_9518,N_8557);
nor U15281 (N_15281,N_8831,N_11346);
or U15282 (N_15282,N_10280,N_10554);
or U15283 (N_15283,N_10620,N_8105);
and U15284 (N_15284,N_10935,N_11454);
or U15285 (N_15285,N_9198,N_11564);
xor U15286 (N_15286,N_11932,N_9673);
or U15287 (N_15287,N_10068,N_11730);
xnor U15288 (N_15288,N_9053,N_8726);
nor U15289 (N_15289,N_11997,N_9461);
nand U15290 (N_15290,N_9794,N_9316);
nor U15291 (N_15291,N_11887,N_8712);
or U15292 (N_15292,N_11671,N_11642);
xnor U15293 (N_15293,N_8674,N_8778);
nor U15294 (N_15294,N_8699,N_9778);
nand U15295 (N_15295,N_8966,N_11650);
or U15296 (N_15296,N_8340,N_9108);
or U15297 (N_15297,N_8479,N_9949);
nand U15298 (N_15298,N_9091,N_10113);
and U15299 (N_15299,N_9525,N_8573);
or U15300 (N_15300,N_9032,N_11818);
nand U15301 (N_15301,N_9603,N_8755);
and U15302 (N_15302,N_9809,N_10517);
and U15303 (N_15303,N_9367,N_9221);
nor U15304 (N_15304,N_10900,N_9352);
nor U15305 (N_15305,N_11411,N_9514);
and U15306 (N_15306,N_10111,N_11912);
or U15307 (N_15307,N_10763,N_8884);
and U15308 (N_15308,N_10808,N_11983);
nor U15309 (N_15309,N_9044,N_10248);
nand U15310 (N_15310,N_9614,N_10223);
nor U15311 (N_15311,N_11822,N_11467);
and U15312 (N_15312,N_10252,N_9620);
nor U15313 (N_15313,N_9819,N_11094);
nor U15314 (N_15314,N_10637,N_8873);
and U15315 (N_15315,N_9678,N_11539);
nand U15316 (N_15316,N_10177,N_11597);
nor U15317 (N_15317,N_9688,N_9090);
nor U15318 (N_15318,N_10326,N_10794);
nand U15319 (N_15319,N_8787,N_8877);
nor U15320 (N_15320,N_9330,N_10277);
nor U15321 (N_15321,N_11599,N_10462);
and U15322 (N_15322,N_10351,N_8813);
nand U15323 (N_15323,N_10385,N_11322);
or U15324 (N_15324,N_11631,N_9133);
xor U15325 (N_15325,N_11714,N_10612);
and U15326 (N_15326,N_8687,N_9021);
or U15327 (N_15327,N_10348,N_8728);
nor U15328 (N_15328,N_8081,N_10947);
nor U15329 (N_15329,N_10948,N_11274);
xor U15330 (N_15330,N_11532,N_11703);
nand U15331 (N_15331,N_8729,N_10620);
nand U15332 (N_15332,N_9629,N_11436);
nor U15333 (N_15333,N_11110,N_11002);
nand U15334 (N_15334,N_10796,N_9356);
xor U15335 (N_15335,N_9222,N_9132);
or U15336 (N_15336,N_10008,N_8065);
or U15337 (N_15337,N_8646,N_11638);
xnor U15338 (N_15338,N_8808,N_9263);
and U15339 (N_15339,N_10618,N_10110);
or U15340 (N_15340,N_10817,N_9436);
or U15341 (N_15341,N_10325,N_8578);
or U15342 (N_15342,N_10237,N_10779);
xor U15343 (N_15343,N_11948,N_9860);
and U15344 (N_15344,N_10286,N_8405);
nor U15345 (N_15345,N_10438,N_10155);
nor U15346 (N_15346,N_8400,N_11375);
and U15347 (N_15347,N_9318,N_9250);
and U15348 (N_15348,N_10398,N_11562);
and U15349 (N_15349,N_10718,N_8956);
or U15350 (N_15350,N_8423,N_8585);
nand U15351 (N_15351,N_8344,N_10216);
nor U15352 (N_15352,N_9944,N_9519);
nor U15353 (N_15353,N_9273,N_10394);
nor U15354 (N_15354,N_11267,N_10069);
xor U15355 (N_15355,N_8069,N_8810);
nor U15356 (N_15356,N_9205,N_8247);
or U15357 (N_15357,N_10309,N_8393);
or U15358 (N_15358,N_8803,N_8092);
nand U15359 (N_15359,N_9054,N_11747);
and U15360 (N_15360,N_10218,N_9308);
nor U15361 (N_15361,N_8871,N_10261);
or U15362 (N_15362,N_11927,N_11994);
or U15363 (N_15363,N_9048,N_9619);
or U15364 (N_15364,N_10014,N_10208);
and U15365 (N_15365,N_8767,N_11955);
and U15366 (N_15366,N_9003,N_11033);
nor U15367 (N_15367,N_8188,N_11977);
nand U15368 (N_15368,N_8954,N_9666);
nor U15369 (N_15369,N_9765,N_10879);
or U15370 (N_15370,N_10794,N_9442);
nand U15371 (N_15371,N_9141,N_11200);
nand U15372 (N_15372,N_9413,N_8654);
nor U15373 (N_15373,N_9957,N_10075);
nor U15374 (N_15374,N_8992,N_9848);
or U15375 (N_15375,N_10983,N_10522);
or U15376 (N_15376,N_10064,N_8659);
nor U15377 (N_15377,N_8409,N_10308);
nor U15378 (N_15378,N_8462,N_8842);
or U15379 (N_15379,N_11519,N_10821);
and U15380 (N_15380,N_8780,N_11914);
xnor U15381 (N_15381,N_10619,N_11227);
and U15382 (N_15382,N_8796,N_8382);
and U15383 (N_15383,N_10571,N_10867);
nand U15384 (N_15384,N_9452,N_9793);
nor U15385 (N_15385,N_8226,N_9206);
and U15386 (N_15386,N_8016,N_10209);
xor U15387 (N_15387,N_9679,N_10345);
xnor U15388 (N_15388,N_10212,N_8089);
xor U15389 (N_15389,N_8701,N_10435);
and U15390 (N_15390,N_8158,N_9949);
nand U15391 (N_15391,N_11651,N_10671);
or U15392 (N_15392,N_9702,N_9254);
xnor U15393 (N_15393,N_8239,N_10570);
nand U15394 (N_15394,N_8728,N_9455);
nand U15395 (N_15395,N_9978,N_9273);
nor U15396 (N_15396,N_8821,N_8308);
or U15397 (N_15397,N_9774,N_9249);
nor U15398 (N_15398,N_9193,N_10710);
xor U15399 (N_15399,N_11669,N_10029);
xor U15400 (N_15400,N_8824,N_11933);
nor U15401 (N_15401,N_10754,N_10749);
or U15402 (N_15402,N_11883,N_11554);
nand U15403 (N_15403,N_9756,N_11500);
and U15404 (N_15404,N_10886,N_8890);
nand U15405 (N_15405,N_8853,N_9833);
and U15406 (N_15406,N_11313,N_11494);
and U15407 (N_15407,N_9504,N_8496);
nand U15408 (N_15408,N_9251,N_8653);
or U15409 (N_15409,N_8076,N_11512);
nand U15410 (N_15410,N_9793,N_10518);
nand U15411 (N_15411,N_10186,N_10618);
nor U15412 (N_15412,N_8302,N_10683);
and U15413 (N_15413,N_9821,N_8701);
nand U15414 (N_15414,N_8458,N_9296);
or U15415 (N_15415,N_8285,N_10746);
nand U15416 (N_15416,N_8513,N_8511);
nand U15417 (N_15417,N_9442,N_9290);
or U15418 (N_15418,N_8215,N_9435);
nand U15419 (N_15419,N_9593,N_11617);
or U15420 (N_15420,N_11422,N_11262);
xnor U15421 (N_15421,N_8455,N_10303);
or U15422 (N_15422,N_11300,N_11898);
and U15423 (N_15423,N_11395,N_9018);
nand U15424 (N_15424,N_9294,N_9926);
nand U15425 (N_15425,N_11080,N_11012);
and U15426 (N_15426,N_9528,N_9044);
nor U15427 (N_15427,N_8688,N_8836);
and U15428 (N_15428,N_10511,N_10823);
nand U15429 (N_15429,N_9427,N_10955);
xor U15430 (N_15430,N_10216,N_8971);
nand U15431 (N_15431,N_10229,N_9117);
or U15432 (N_15432,N_9177,N_10695);
nor U15433 (N_15433,N_9292,N_9868);
xnor U15434 (N_15434,N_9040,N_10791);
or U15435 (N_15435,N_10352,N_11774);
nand U15436 (N_15436,N_11929,N_8298);
and U15437 (N_15437,N_8548,N_11697);
and U15438 (N_15438,N_11251,N_11802);
nor U15439 (N_15439,N_10337,N_9844);
or U15440 (N_15440,N_8883,N_11552);
and U15441 (N_15441,N_10452,N_8773);
nand U15442 (N_15442,N_11322,N_8111);
nand U15443 (N_15443,N_10057,N_10534);
and U15444 (N_15444,N_10677,N_10397);
nor U15445 (N_15445,N_9391,N_10585);
nor U15446 (N_15446,N_11458,N_9928);
or U15447 (N_15447,N_9671,N_11607);
nor U15448 (N_15448,N_8307,N_8396);
or U15449 (N_15449,N_9703,N_11803);
and U15450 (N_15450,N_9421,N_10360);
xnor U15451 (N_15451,N_10545,N_10942);
xor U15452 (N_15452,N_11770,N_9655);
nand U15453 (N_15453,N_10245,N_10354);
or U15454 (N_15454,N_11214,N_8722);
xnor U15455 (N_15455,N_10099,N_10518);
nor U15456 (N_15456,N_8121,N_9051);
or U15457 (N_15457,N_10512,N_10491);
nand U15458 (N_15458,N_9621,N_11719);
nand U15459 (N_15459,N_11755,N_10110);
and U15460 (N_15460,N_8263,N_9202);
nand U15461 (N_15461,N_8756,N_11789);
or U15462 (N_15462,N_9771,N_8384);
or U15463 (N_15463,N_8297,N_10569);
and U15464 (N_15464,N_9790,N_10084);
nand U15465 (N_15465,N_11969,N_8263);
nand U15466 (N_15466,N_10416,N_11120);
or U15467 (N_15467,N_11568,N_8363);
nor U15468 (N_15468,N_10109,N_8277);
and U15469 (N_15469,N_8183,N_9184);
or U15470 (N_15470,N_9341,N_10704);
and U15471 (N_15471,N_10423,N_10868);
nor U15472 (N_15472,N_8379,N_11224);
and U15473 (N_15473,N_9868,N_10377);
nand U15474 (N_15474,N_10413,N_9808);
nor U15475 (N_15475,N_11550,N_8632);
and U15476 (N_15476,N_8733,N_11896);
or U15477 (N_15477,N_11759,N_11918);
or U15478 (N_15478,N_11368,N_10016);
nor U15479 (N_15479,N_10941,N_9302);
nand U15480 (N_15480,N_11355,N_8321);
and U15481 (N_15481,N_8980,N_9103);
and U15482 (N_15482,N_8525,N_10194);
nor U15483 (N_15483,N_11672,N_11182);
or U15484 (N_15484,N_8121,N_9385);
nand U15485 (N_15485,N_8312,N_8435);
nor U15486 (N_15486,N_8628,N_9261);
and U15487 (N_15487,N_11294,N_11445);
nand U15488 (N_15488,N_8626,N_11692);
xor U15489 (N_15489,N_9320,N_8331);
xor U15490 (N_15490,N_8933,N_10074);
nor U15491 (N_15491,N_11615,N_8164);
or U15492 (N_15492,N_9205,N_11702);
nor U15493 (N_15493,N_9042,N_8311);
or U15494 (N_15494,N_9740,N_10511);
nand U15495 (N_15495,N_8363,N_9253);
and U15496 (N_15496,N_11262,N_8239);
nor U15497 (N_15497,N_8909,N_11275);
nand U15498 (N_15498,N_8231,N_11271);
or U15499 (N_15499,N_10166,N_8634);
nand U15500 (N_15500,N_8769,N_8955);
nand U15501 (N_15501,N_8506,N_10180);
and U15502 (N_15502,N_9442,N_11426);
or U15503 (N_15503,N_8561,N_8660);
and U15504 (N_15504,N_9129,N_10476);
nor U15505 (N_15505,N_8929,N_10853);
nor U15506 (N_15506,N_11397,N_10997);
nand U15507 (N_15507,N_11060,N_9176);
and U15508 (N_15508,N_10871,N_10013);
xnor U15509 (N_15509,N_10016,N_11456);
and U15510 (N_15510,N_11736,N_8822);
and U15511 (N_15511,N_10771,N_8649);
xnor U15512 (N_15512,N_10129,N_11353);
nor U15513 (N_15513,N_11088,N_9762);
nor U15514 (N_15514,N_8113,N_9537);
nand U15515 (N_15515,N_9235,N_11834);
nor U15516 (N_15516,N_10417,N_10456);
nand U15517 (N_15517,N_9770,N_9877);
nor U15518 (N_15518,N_10475,N_9040);
or U15519 (N_15519,N_10924,N_8452);
and U15520 (N_15520,N_9851,N_11126);
nor U15521 (N_15521,N_9306,N_10292);
nor U15522 (N_15522,N_11758,N_9180);
nor U15523 (N_15523,N_11259,N_11175);
nand U15524 (N_15524,N_10026,N_10510);
or U15525 (N_15525,N_8290,N_8004);
and U15526 (N_15526,N_9140,N_11305);
and U15527 (N_15527,N_11273,N_8797);
and U15528 (N_15528,N_11385,N_9937);
and U15529 (N_15529,N_10623,N_11350);
and U15530 (N_15530,N_9482,N_11037);
nor U15531 (N_15531,N_10374,N_10615);
and U15532 (N_15532,N_9653,N_9530);
nand U15533 (N_15533,N_11051,N_10855);
and U15534 (N_15534,N_8584,N_8468);
xor U15535 (N_15535,N_8302,N_11936);
xor U15536 (N_15536,N_8818,N_9814);
nor U15537 (N_15537,N_10763,N_10432);
nand U15538 (N_15538,N_9430,N_11660);
nor U15539 (N_15539,N_11069,N_8713);
nand U15540 (N_15540,N_8561,N_10915);
nand U15541 (N_15541,N_11646,N_10763);
and U15542 (N_15542,N_8762,N_8456);
and U15543 (N_15543,N_9341,N_9455);
and U15544 (N_15544,N_8288,N_11010);
and U15545 (N_15545,N_11772,N_8728);
and U15546 (N_15546,N_10602,N_11208);
xor U15547 (N_15547,N_8257,N_10156);
nand U15548 (N_15548,N_11868,N_11606);
and U15549 (N_15549,N_10376,N_9872);
and U15550 (N_15550,N_11452,N_9971);
nor U15551 (N_15551,N_8966,N_10506);
and U15552 (N_15552,N_10098,N_8960);
nand U15553 (N_15553,N_11216,N_11357);
nand U15554 (N_15554,N_11617,N_9948);
or U15555 (N_15555,N_8278,N_11312);
or U15556 (N_15556,N_11937,N_9488);
nor U15557 (N_15557,N_11869,N_10849);
nand U15558 (N_15558,N_9815,N_9916);
or U15559 (N_15559,N_8043,N_9946);
nand U15560 (N_15560,N_8447,N_9685);
nor U15561 (N_15561,N_10673,N_8038);
xnor U15562 (N_15562,N_9334,N_8866);
and U15563 (N_15563,N_10967,N_11918);
nand U15564 (N_15564,N_11263,N_11417);
nor U15565 (N_15565,N_11409,N_8470);
nor U15566 (N_15566,N_11940,N_10385);
xnor U15567 (N_15567,N_8435,N_9933);
and U15568 (N_15568,N_10000,N_10233);
xor U15569 (N_15569,N_10512,N_9836);
nand U15570 (N_15570,N_10337,N_11308);
or U15571 (N_15571,N_9378,N_10836);
nand U15572 (N_15572,N_10801,N_10047);
nand U15573 (N_15573,N_9586,N_8987);
nor U15574 (N_15574,N_9789,N_11014);
nor U15575 (N_15575,N_9771,N_11454);
and U15576 (N_15576,N_9374,N_9439);
nor U15577 (N_15577,N_11612,N_9087);
or U15578 (N_15578,N_11814,N_11000);
nor U15579 (N_15579,N_9511,N_8897);
nor U15580 (N_15580,N_8674,N_10296);
or U15581 (N_15581,N_10924,N_9413);
or U15582 (N_15582,N_11885,N_11909);
nor U15583 (N_15583,N_8820,N_10365);
or U15584 (N_15584,N_9609,N_11773);
and U15585 (N_15585,N_8176,N_10731);
xnor U15586 (N_15586,N_9593,N_11832);
and U15587 (N_15587,N_10213,N_9112);
nor U15588 (N_15588,N_9185,N_10577);
xnor U15589 (N_15589,N_8555,N_9824);
or U15590 (N_15590,N_10015,N_11816);
nor U15591 (N_15591,N_9298,N_8986);
and U15592 (N_15592,N_11471,N_11942);
nor U15593 (N_15593,N_8597,N_10385);
or U15594 (N_15594,N_10329,N_9243);
nor U15595 (N_15595,N_8988,N_10181);
and U15596 (N_15596,N_11844,N_9169);
or U15597 (N_15597,N_9821,N_10990);
or U15598 (N_15598,N_11097,N_9610);
and U15599 (N_15599,N_11478,N_9977);
xnor U15600 (N_15600,N_9879,N_11239);
xor U15601 (N_15601,N_8140,N_8742);
and U15602 (N_15602,N_11249,N_8241);
xor U15603 (N_15603,N_9320,N_11956);
nor U15604 (N_15604,N_9532,N_10070);
nand U15605 (N_15605,N_10132,N_8626);
or U15606 (N_15606,N_10028,N_8955);
and U15607 (N_15607,N_10358,N_9105);
xor U15608 (N_15608,N_8395,N_11583);
nor U15609 (N_15609,N_11707,N_10962);
nand U15610 (N_15610,N_8098,N_10620);
nor U15611 (N_15611,N_9100,N_8589);
nand U15612 (N_15612,N_9171,N_8978);
or U15613 (N_15613,N_11592,N_9381);
nand U15614 (N_15614,N_10196,N_11966);
nor U15615 (N_15615,N_10963,N_9684);
nor U15616 (N_15616,N_10509,N_11461);
nor U15617 (N_15617,N_9694,N_9621);
nor U15618 (N_15618,N_11389,N_8844);
or U15619 (N_15619,N_9253,N_11481);
and U15620 (N_15620,N_10455,N_10595);
nand U15621 (N_15621,N_9778,N_11717);
nor U15622 (N_15622,N_9297,N_8982);
or U15623 (N_15623,N_8310,N_11103);
nor U15624 (N_15624,N_9090,N_8868);
or U15625 (N_15625,N_10433,N_8514);
xnor U15626 (N_15626,N_8724,N_10282);
xnor U15627 (N_15627,N_10164,N_11262);
xor U15628 (N_15628,N_9773,N_9665);
nor U15629 (N_15629,N_9234,N_11919);
nor U15630 (N_15630,N_9845,N_10796);
nand U15631 (N_15631,N_8159,N_11005);
nand U15632 (N_15632,N_8172,N_8163);
nor U15633 (N_15633,N_8504,N_9217);
nor U15634 (N_15634,N_11473,N_8810);
or U15635 (N_15635,N_11113,N_9577);
nor U15636 (N_15636,N_10837,N_11315);
and U15637 (N_15637,N_8618,N_11351);
nor U15638 (N_15638,N_8279,N_8782);
xnor U15639 (N_15639,N_9040,N_8218);
nand U15640 (N_15640,N_9475,N_11396);
nor U15641 (N_15641,N_10049,N_9596);
or U15642 (N_15642,N_11577,N_8540);
or U15643 (N_15643,N_10219,N_8779);
or U15644 (N_15644,N_11132,N_9509);
nand U15645 (N_15645,N_11994,N_8363);
or U15646 (N_15646,N_11804,N_8423);
or U15647 (N_15647,N_9539,N_9162);
or U15648 (N_15648,N_9895,N_9586);
and U15649 (N_15649,N_10779,N_8662);
nand U15650 (N_15650,N_10802,N_9818);
and U15651 (N_15651,N_11452,N_8075);
and U15652 (N_15652,N_8625,N_9431);
xnor U15653 (N_15653,N_10533,N_10451);
or U15654 (N_15654,N_10607,N_11344);
nand U15655 (N_15655,N_10161,N_9607);
and U15656 (N_15656,N_11305,N_11872);
nor U15657 (N_15657,N_10341,N_11246);
and U15658 (N_15658,N_8689,N_9390);
nand U15659 (N_15659,N_9776,N_9226);
xnor U15660 (N_15660,N_9081,N_10741);
nor U15661 (N_15661,N_11256,N_8897);
and U15662 (N_15662,N_11697,N_9702);
or U15663 (N_15663,N_10187,N_9056);
or U15664 (N_15664,N_11224,N_11510);
nor U15665 (N_15665,N_10773,N_9316);
and U15666 (N_15666,N_9450,N_11524);
nand U15667 (N_15667,N_10090,N_8683);
nor U15668 (N_15668,N_8592,N_8966);
or U15669 (N_15669,N_10233,N_9788);
or U15670 (N_15670,N_9806,N_8307);
and U15671 (N_15671,N_9720,N_8726);
xnor U15672 (N_15672,N_8252,N_9707);
nand U15673 (N_15673,N_8647,N_8289);
nor U15674 (N_15674,N_10312,N_9052);
and U15675 (N_15675,N_10053,N_11474);
nor U15676 (N_15676,N_11753,N_11471);
xnor U15677 (N_15677,N_11982,N_9935);
nand U15678 (N_15678,N_11303,N_11576);
and U15679 (N_15679,N_9717,N_11378);
and U15680 (N_15680,N_10249,N_9024);
nand U15681 (N_15681,N_8574,N_9201);
nand U15682 (N_15682,N_11079,N_9836);
and U15683 (N_15683,N_11562,N_11079);
or U15684 (N_15684,N_8742,N_8229);
nor U15685 (N_15685,N_11446,N_11663);
or U15686 (N_15686,N_10784,N_10120);
and U15687 (N_15687,N_9277,N_11533);
and U15688 (N_15688,N_8198,N_11567);
and U15689 (N_15689,N_10137,N_11719);
and U15690 (N_15690,N_10495,N_10671);
nor U15691 (N_15691,N_10763,N_8717);
or U15692 (N_15692,N_9610,N_11803);
and U15693 (N_15693,N_11329,N_9672);
and U15694 (N_15694,N_8514,N_9896);
nand U15695 (N_15695,N_11162,N_9418);
xnor U15696 (N_15696,N_9043,N_11703);
xnor U15697 (N_15697,N_9341,N_10147);
nor U15698 (N_15698,N_10008,N_10229);
xor U15699 (N_15699,N_9476,N_10556);
and U15700 (N_15700,N_11061,N_8165);
nor U15701 (N_15701,N_11109,N_10768);
xor U15702 (N_15702,N_10262,N_8954);
and U15703 (N_15703,N_8154,N_10094);
nor U15704 (N_15704,N_8405,N_10865);
nor U15705 (N_15705,N_10442,N_9007);
nand U15706 (N_15706,N_8623,N_11061);
nand U15707 (N_15707,N_9160,N_8715);
or U15708 (N_15708,N_10489,N_9307);
nor U15709 (N_15709,N_11437,N_8346);
xor U15710 (N_15710,N_11160,N_11613);
and U15711 (N_15711,N_10764,N_11778);
nor U15712 (N_15712,N_9044,N_11170);
or U15713 (N_15713,N_11505,N_9652);
nor U15714 (N_15714,N_10135,N_10292);
and U15715 (N_15715,N_11663,N_8736);
nand U15716 (N_15716,N_10004,N_8612);
nor U15717 (N_15717,N_9953,N_9571);
nor U15718 (N_15718,N_10190,N_8153);
and U15719 (N_15719,N_10226,N_8676);
and U15720 (N_15720,N_10946,N_10985);
or U15721 (N_15721,N_8103,N_9559);
nor U15722 (N_15722,N_11376,N_11408);
nand U15723 (N_15723,N_8585,N_8184);
nand U15724 (N_15724,N_11636,N_9615);
or U15725 (N_15725,N_8548,N_8252);
and U15726 (N_15726,N_10468,N_8140);
nor U15727 (N_15727,N_9524,N_10456);
nand U15728 (N_15728,N_11946,N_10424);
or U15729 (N_15729,N_11725,N_9503);
nand U15730 (N_15730,N_8920,N_10507);
or U15731 (N_15731,N_8372,N_11226);
or U15732 (N_15732,N_10991,N_9548);
xnor U15733 (N_15733,N_9736,N_9281);
nand U15734 (N_15734,N_10000,N_11488);
or U15735 (N_15735,N_10588,N_10939);
nand U15736 (N_15736,N_11418,N_10417);
or U15737 (N_15737,N_9426,N_8224);
xor U15738 (N_15738,N_8829,N_9494);
nand U15739 (N_15739,N_11599,N_9079);
xor U15740 (N_15740,N_9269,N_11671);
xor U15741 (N_15741,N_9146,N_9448);
nand U15742 (N_15742,N_11389,N_9145);
nor U15743 (N_15743,N_10645,N_9705);
nand U15744 (N_15744,N_11243,N_10779);
nor U15745 (N_15745,N_11098,N_9394);
and U15746 (N_15746,N_8845,N_10318);
nand U15747 (N_15747,N_8876,N_11437);
nand U15748 (N_15748,N_10135,N_9086);
nand U15749 (N_15749,N_10272,N_10162);
xnor U15750 (N_15750,N_11715,N_11060);
and U15751 (N_15751,N_10713,N_11532);
nor U15752 (N_15752,N_8485,N_8829);
and U15753 (N_15753,N_11732,N_11418);
nand U15754 (N_15754,N_11726,N_11858);
and U15755 (N_15755,N_9332,N_11354);
nand U15756 (N_15756,N_9246,N_9181);
nand U15757 (N_15757,N_8089,N_8781);
xnor U15758 (N_15758,N_9318,N_9452);
or U15759 (N_15759,N_9881,N_10467);
nor U15760 (N_15760,N_10613,N_11829);
nand U15761 (N_15761,N_11653,N_9055);
and U15762 (N_15762,N_11308,N_9952);
or U15763 (N_15763,N_9504,N_11037);
and U15764 (N_15764,N_10662,N_8806);
and U15765 (N_15765,N_11043,N_9191);
nand U15766 (N_15766,N_8218,N_11795);
nor U15767 (N_15767,N_8588,N_11058);
or U15768 (N_15768,N_10295,N_10471);
or U15769 (N_15769,N_9797,N_10898);
nor U15770 (N_15770,N_11098,N_8466);
or U15771 (N_15771,N_10154,N_9804);
and U15772 (N_15772,N_8782,N_10165);
nor U15773 (N_15773,N_8321,N_11433);
and U15774 (N_15774,N_8278,N_11299);
xor U15775 (N_15775,N_11502,N_10117);
nand U15776 (N_15776,N_8570,N_8652);
or U15777 (N_15777,N_8153,N_9692);
nand U15778 (N_15778,N_10216,N_10918);
xnor U15779 (N_15779,N_11331,N_11657);
nand U15780 (N_15780,N_10570,N_10096);
nor U15781 (N_15781,N_9098,N_11989);
nand U15782 (N_15782,N_11803,N_10573);
xnor U15783 (N_15783,N_10075,N_8996);
and U15784 (N_15784,N_10569,N_8263);
and U15785 (N_15785,N_10837,N_11029);
nor U15786 (N_15786,N_9034,N_10460);
nand U15787 (N_15787,N_10505,N_8382);
nand U15788 (N_15788,N_10936,N_10355);
nor U15789 (N_15789,N_9874,N_11542);
nor U15790 (N_15790,N_10613,N_9282);
nand U15791 (N_15791,N_11187,N_9270);
and U15792 (N_15792,N_11200,N_11620);
and U15793 (N_15793,N_11139,N_8098);
nor U15794 (N_15794,N_10758,N_9579);
xor U15795 (N_15795,N_9110,N_10412);
nand U15796 (N_15796,N_10991,N_9078);
nor U15797 (N_15797,N_9961,N_8063);
and U15798 (N_15798,N_8600,N_8512);
nand U15799 (N_15799,N_10818,N_9108);
nand U15800 (N_15800,N_10700,N_11917);
nor U15801 (N_15801,N_8617,N_11922);
xnor U15802 (N_15802,N_10010,N_10251);
nand U15803 (N_15803,N_11465,N_11877);
and U15804 (N_15804,N_8924,N_11380);
xor U15805 (N_15805,N_9240,N_10826);
and U15806 (N_15806,N_11976,N_11620);
xor U15807 (N_15807,N_8731,N_10025);
or U15808 (N_15808,N_9549,N_11801);
nor U15809 (N_15809,N_8992,N_11477);
nand U15810 (N_15810,N_8991,N_9695);
nor U15811 (N_15811,N_10629,N_8588);
and U15812 (N_15812,N_11756,N_9531);
or U15813 (N_15813,N_10342,N_8335);
and U15814 (N_15814,N_8677,N_11384);
and U15815 (N_15815,N_8385,N_9495);
and U15816 (N_15816,N_8631,N_9374);
and U15817 (N_15817,N_9951,N_8297);
or U15818 (N_15818,N_10418,N_9143);
nor U15819 (N_15819,N_11404,N_10998);
nor U15820 (N_15820,N_10652,N_8496);
nand U15821 (N_15821,N_11774,N_10116);
and U15822 (N_15822,N_8886,N_9124);
or U15823 (N_15823,N_9722,N_9569);
nand U15824 (N_15824,N_10685,N_11941);
nor U15825 (N_15825,N_10638,N_10192);
or U15826 (N_15826,N_9034,N_10154);
nor U15827 (N_15827,N_11692,N_11516);
nor U15828 (N_15828,N_11295,N_10384);
and U15829 (N_15829,N_11162,N_9677);
nand U15830 (N_15830,N_8589,N_9041);
and U15831 (N_15831,N_9379,N_8224);
and U15832 (N_15832,N_8327,N_9878);
and U15833 (N_15833,N_9301,N_8684);
nand U15834 (N_15834,N_8550,N_11565);
or U15835 (N_15835,N_9814,N_10992);
nor U15836 (N_15836,N_10631,N_10252);
and U15837 (N_15837,N_8659,N_8301);
and U15838 (N_15838,N_8687,N_9068);
or U15839 (N_15839,N_8603,N_10928);
and U15840 (N_15840,N_8554,N_9656);
nand U15841 (N_15841,N_11896,N_8664);
or U15842 (N_15842,N_11890,N_11223);
xnor U15843 (N_15843,N_10726,N_11188);
or U15844 (N_15844,N_10183,N_11116);
or U15845 (N_15845,N_8440,N_11211);
nand U15846 (N_15846,N_8319,N_11438);
or U15847 (N_15847,N_10010,N_11637);
nand U15848 (N_15848,N_8487,N_8761);
or U15849 (N_15849,N_8963,N_11509);
nand U15850 (N_15850,N_8045,N_8489);
nand U15851 (N_15851,N_11824,N_8722);
nor U15852 (N_15852,N_9965,N_9223);
and U15853 (N_15853,N_11900,N_11628);
or U15854 (N_15854,N_11213,N_8875);
nand U15855 (N_15855,N_8516,N_11302);
and U15856 (N_15856,N_8258,N_10257);
nand U15857 (N_15857,N_11610,N_11894);
and U15858 (N_15858,N_8846,N_11793);
and U15859 (N_15859,N_8457,N_10903);
and U15860 (N_15860,N_11372,N_10433);
nor U15861 (N_15861,N_11463,N_8272);
nor U15862 (N_15862,N_8340,N_10638);
and U15863 (N_15863,N_9260,N_11646);
and U15864 (N_15864,N_9056,N_11465);
and U15865 (N_15865,N_10039,N_8375);
and U15866 (N_15866,N_8612,N_11318);
nand U15867 (N_15867,N_9611,N_9630);
and U15868 (N_15868,N_8871,N_10952);
and U15869 (N_15869,N_10607,N_11459);
nor U15870 (N_15870,N_9874,N_9367);
and U15871 (N_15871,N_11904,N_11049);
nor U15872 (N_15872,N_9060,N_8115);
nor U15873 (N_15873,N_11763,N_11349);
nor U15874 (N_15874,N_10332,N_8966);
nor U15875 (N_15875,N_11182,N_11458);
nand U15876 (N_15876,N_10514,N_9803);
and U15877 (N_15877,N_8530,N_9202);
nor U15878 (N_15878,N_9923,N_10074);
nor U15879 (N_15879,N_9869,N_11883);
and U15880 (N_15880,N_8500,N_9960);
nor U15881 (N_15881,N_9978,N_9265);
or U15882 (N_15882,N_10039,N_10356);
nand U15883 (N_15883,N_11899,N_8719);
xor U15884 (N_15884,N_9046,N_8390);
and U15885 (N_15885,N_11359,N_10247);
or U15886 (N_15886,N_10809,N_11733);
xnor U15887 (N_15887,N_10439,N_11089);
or U15888 (N_15888,N_10477,N_8453);
and U15889 (N_15889,N_8476,N_11758);
and U15890 (N_15890,N_8188,N_11955);
or U15891 (N_15891,N_11608,N_11092);
xor U15892 (N_15892,N_11842,N_8299);
nand U15893 (N_15893,N_10133,N_9860);
xnor U15894 (N_15894,N_9779,N_8619);
and U15895 (N_15895,N_9426,N_8854);
and U15896 (N_15896,N_8756,N_8465);
and U15897 (N_15897,N_10763,N_9460);
xor U15898 (N_15898,N_11553,N_11613);
and U15899 (N_15899,N_10203,N_9812);
nand U15900 (N_15900,N_8882,N_8172);
nand U15901 (N_15901,N_10613,N_11852);
and U15902 (N_15902,N_10119,N_8619);
or U15903 (N_15903,N_9413,N_9779);
nand U15904 (N_15904,N_11020,N_8392);
and U15905 (N_15905,N_9007,N_11121);
and U15906 (N_15906,N_11320,N_10815);
nand U15907 (N_15907,N_10859,N_10344);
and U15908 (N_15908,N_10101,N_11122);
nand U15909 (N_15909,N_8466,N_8588);
or U15910 (N_15910,N_8864,N_11274);
or U15911 (N_15911,N_11383,N_8332);
nor U15912 (N_15912,N_10442,N_10989);
and U15913 (N_15913,N_10053,N_10070);
nand U15914 (N_15914,N_11265,N_10803);
nor U15915 (N_15915,N_11504,N_11404);
nor U15916 (N_15916,N_10685,N_8065);
nand U15917 (N_15917,N_11312,N_9418);
nor U15918 (N_15918,N_11535,N_10124);
or U15919 (N_15919,N_8756,N_11305);
nor U15920 (N_15920,N_8505,N_11847);
or U15921 (N_15921,N_10294,N_8414);
nand U15922 (N_15922,N_9043,N_11743);
and U15923 (N_15923,N_8294,N_8974);
nor U15924 (N_15924,N_9158,N_8407);
and U15925 (N_15925,N_8763,N_8040);
nand U15926 (N_15926,N_11457,N_11580);
and U15927 (N_15927,N_9693,N_11426);
xnor U15928 (N_15928,N_10908,N_8246);
nor U15929 (N_15929,N_8939,N_9963);
nand U15930 (N_15930,N_10230,N_11616);
xnor U15931 (N_15931,N_10976,N_8310);
nand U15932 (N_15932,N_10271,N_8088);
nand U15933 (N_15933,N_9579,N_9556);
or U15934 (N_15934,N_8084,N_11732);
nor U15935 (N_15935,N_11813,N_8292);
nor U15936 (N_15936,N_8924,N_8733);
nand U15937 (N_15937,N_8996,N_10988);
and U15938 (N_15938,N_9390,N_9685);
nand U15939 (N_15939,N_9838,N_8126);
or U15940 (N_15940,N_9604,N_9497);
or U15941 (N_15941,N_11487,N_11801);
xnor U15942 (N_15942,N_9196,N_11510);
and U15943 (N_15943,N_10344,N_9990);
and U15944 (N_15944,N_9521,N_9538);
nand U15945 (N_15945,N_9280,N_9870);
nor U15946 (N_15946,N_10336,N_8667);
and U15947 (N_15947,N_10252,N_11943);
nand U15948 (N_15948,N_10161,N_8317);
nor U15949 (N_15949,N_8176,N_8341);
or U15950 (N_15950,N_8261,N_9046);
nand U15951 (N_15951,N_10874,N_8581);
or U15952 (N_15952,N_11876,N_9283);
nor U15953 (N_15953,N_8720,N_11928);
nor U15954 (N_15954,N_11466,N_9649);
or U15955 (N_15955,N_11045,N_9884);
nor U15956 (N_15956,N_9835,N_9144);
nor U15957 (N_15957,N_10509,N_8437);
or U15958 (N_15958,N_11934,N_8381);
xnor U15959 (N_15959,N_9367,N_9565);
xor U15960 (N_15960,N_9978,N_9739);
nor U15961 (N_15961,N_10264,N_9415);
and U15962 (N_15962,N_9971,N_11751);
and U15963 (N_15963,N_10907,N_10026);
nor U15964 (N_15964,N_11775,N_10086);
or U15965 (N_15965,N_10524,N_10569);
nor U15966 (N_15966,N_9136,N_9170);
and U15967 (N_15967,N_8270,N_11276);
and U15968 (N_15968,N_11557,N_10837);
or U15969 (N_15969,N_10488,N_8587);
or U15970 (N_15970,N_10370,N_9641);
nor U15971 (N_15971,N_11870,N_9615);
nand U15972 (N_15972,N_11932,N_8204);
xnor U15973 (N_15973,N_9852,N_11298);
nor U15974 (N_15974,N_10677,N_9246);
xnor U15975 (N_15975,N_10707,N_9250);
and U15976 (N_15976,N_8406,N_11639);
and U15977 (N_15977,N_10332,N_8995);
and U15978 (N_15978,N_11764,N_8336);
nand U15979 (N_15979,N_11030,N_10237);
or U15980 (N_15980,N_8701,N_11982);
or U15981 (N_15981,N_8786,N_10520);
nor U15982 (N_15982,N_10960,N_9974);
nand U15983 (N_15983,N_9174,N_9108);
nor U15984 (N_15984,N_9825,N_10442);
and U15985 (N_15985,N_10620,N_8229);
or U15986 (N_15986,N_8540,N_9085);
or U15987 (N_15987,N_8440,N_9883);
and U15988 (N_15988,N_11581,N_10573);
nand U15989 (N_15989,N_11363,N_9420);
or U15990 (N_15990,N_9582,N_8073);
nand U15991 (N_15991,N_10269,N_10306);
nor U15992 (N_15992,N_10165,N_10587);
and U15993 (N_15993,N_8913,N_8115);
or U15994 (N_15994,N_11417,N_11078);
nand U15995 (N_15995,N_8318,N_11286);
and U15996 (N_15996,N_9254,N_10303);
or U15997 (N_15997,N_11511,N_11244);
and U15998 (N_15998,N_9711,N_9409);
and U15999 (N_15999,N_10081,N_8871);
nor U16000 (N_16000,N_12213,N_15165);
nand U16001 (N_16001,N_12640,N_15519);
and U16002 (N_16002,N_13814,N_14920);
or U16003 (N_16003,N_13446,N_13014);
nor U16004 (N_16004,N_14610,N_14144);
and U16005 (N_16005,N_15623,N_13623);
nand U16006 (N_16006,N_13862,N_12052);
nand U16007 (N_16007,N_12317,N_14199);
nor U16008 (N_16008,N_15375,N_13418);
or U16009 (N_16009,N_13806,N_15803);
nand U16010 (N_16010,N_15755,N_12014);
and U16011 (N_16011,N_14376,N_12827);
nor U16012 (N_16012,N_14935,N_14222);
nand U16013 (N_16013,N_13502,N_12542);
and U16014 (N_16014,N_14903,N_12965);
and U16015 (N_16015,N_12584,N_13302);
or U16016 (N_16016,N_12600,N_14491);
and U16017 (N_16017,N_13507,N_12651);
and U16018 (N_16018,N_14927,N_12670);
nand U16019 (N_16019,N_12249,N_14671);
and U16020 (N_16020,N_12383,N_13849);
nand U16021 (N_16021,N_15643,N_13669);
and U16022 (N_16022,N_13140,N_15204);
nor U16023 (N_16023,N_15368,N_12268);
and U16024 (N_16024,N_13064,N_15957);
xnor U16025 (N_16025,N_12215,N_14215);
or U16026 (N_16026,N_13406,N_13206);
nand U16027 (N_16027,N_14220,N_15489);
or U16028 (N_16028,N_15638,N_13096);
nand U16029 (N_16029,N_12593,N_13033);
nor U16030 (N_16030,N_14519,N_15828);
and U16031 (N_16031,N_13467,N_13540);
and U16032 (N_16032,N_13311,N_13444);
and U16033 (N_16033,N_14119,N_12531);
or U16034 (N_16034,N_12981,N_15230);
and U16035 (N_16035,N_12064,N_15433);
xnor U16036 (N_16036,N_14345,N_14625);
nand U16037 (N_16037,N_14623,N_15684);
nor U16038 (N_16038,N_14476,N_14153);
nor U16039 (N_16039,N_13553,N_12001);
nor U16040 (N_16040,N_13437,N_14657);
or U16041 (N_16041,N_12252,N_13589);
xnor U16042 (N_16042,N_13821,N_14471);
nor U16043 (N_16043,N_12655,N_15327);
xnor U16044 (N_16044,N_14238,N_13092);
or U16045 (N_16045,N_12716,N_14255);
xor U16046 (N_16046,N_12950,N_12100);
nor U16047 (N_16047,N_14979,N_12028);
nor U16048 (N_16048,N_13296,N_12217);
nand U16049 (N_16049,N_15309,N_12909);
and U16050 (N_16050,N_15482,N_15942);
xnor U16051 (N_16051,N_14869,N_13027);
or U16052 (N_16052,N_12534,N_13115);
nor U16053 (N_16053,N_12994,N_13369);
nor U16054 (N_16054,N_13591,N_15915);
nor U16055 (N_16055,N_14373,N_14197);
or U16056 (N_16056,N_13327,N_15123);
nor U16057 (N_16057,N_13166,N_12646);
and U16058 (N_16058,N_13390,N_15979);
or U16059 (N_16059,N_15164,N_14660);
nor U16060 (N_16060,N_13240,N_13537);
nor U16061 (N_16061,N_12857,N_13161);
xnor U16062 (N_16062,N_12068,N_12492);
and U16063 (N_16063,N_13928,N_12725);
and U16064 (N_16064,N_15462,N_14021);
or U16065 (N_16065,N_15751,N_12979);
xnor U16066 (N_16066,N_14123,N_12825);
nor U16067 (N_16067,N_13035,N_14630);
nand U16068 (N_16068,N_12080,N_13813);
or U16069 (N_16069,N_14567,N_15619);
nor U16070 (N_16070,N_13457,N_15146);
or U16071 (N_16071,N_14730,N_15762);
nor U16072 (N_16072,N_14246,N_14067);
or U16073 (N_16073,N_15155,N_12387);
nand U16074 (N_16074,N_12490,N_14666);
and U16075 (N_16075,N_13668,N_15088);
or U16076 (N_16076,N_15074,N_12206);
and U16077 (N_16077,N_12937,N_15894);
or U16078 (N_16078,N_13337,N_14125);
nand U16079 (N_16079,N_12609,N_12495);
and U16080 (N_16080,N_12897,N_12508);
nand U16081 (N_16081,N_14158,N_12737);
or U16082 (N_16082,N_14540,N_14839);
and U16083 (N_16083,N_12910,N_14670);
xnor U16084 (N_16084,N_12294,N_12266);
nand U16085 (N_16085,N_15882,N_14472);
nor U16086 (N_16086,N_15516,N_12930);
and U16087 (N_16087,N_15350,N_15596);
nand U16088 (N_16088,N_13153,N_15170);
or U16089 (N_16089,N_13009,N_12493);
nand U16090 (N_16090,N_13313,N_14664);
nand U16091 (N_16091,N_13995,N_12873);
nor U16092 (N_16092,N_15817,N_15635);
nand U16093 (N_16093,N_12742,N_14554);
or U16094 (N_16094,N_15238,N_14769);
nand U16095 (N_16095,N_14804,N_15911);
or U16096 (N_16096,N_14480,N_12037);
and U16097 (N_16097,N_13550,N_14892);
and U16098 (N_16098,N_15562,N_12688);
and U16099 (N_16099,N_14915,N_14088);
nand U16100 (N_16100,N_13579,N_14542);
and U16101 (N_16101,N_15026,N_15244);
or U16102 (N_16102,N_12704,N_12118);
or U16103 (N_16103,N_13950,N_15852);
or U16104 (N_16104,N_14284,N_12024);
and U16105 (N_16105,N_13341,N_14016);
and U16106 (N_16106,N_15655,N_15842);
and U16107 (N_16107,N_14868,N_13793);
nor U16108 (N_16108,N_13721,N_12861);
xor U16109 (N_16109,N_13134,N_15767);
and U16110 (N_16110,N_13643,N_13970);
or U16111 (N_16111,N_15268,N_14260);
nand U16112 (N_16112,N_13097,N_14663);
nor U16113 (N_16113,N_12958,N_15058);
nand U16114 (N_16114,N_14518,N_15838);
and U16115 (N_16115,N_13656,N_15272);
nand U16116 (N_16116,N_12447,N_12788);
nor U16117 (N_16117,N_15428,N_13866);
and U16118 (N_16118,N_15484,N_12479);
nand U16119 (N_16119,N_15880,N_13275);
and U16120 (N_16120,N_12871,N_15395);
nand U16121 (N_16121,N_12812,N_12814);
and U16122 (N_16122,N_15711,N_14589);
nand U16123 (N_16123,N_13262,N_13081);
or U16124 (N_16124,N_13394,N_13864);
nor U16125 (N_16125,N_15132,N_15879);
and U16126 (N_16126,N_12803,N_14668);
and U16127 (N_16127,N_13521,N_15399);
xor U16128 (N_16128,N_12468,N_15210);
and U16129 (N_16129,N_12603,N_15658);
xor U16130 (N_16130,N_14866,N_12648);
nor U16131 (N_16131,N_12560,N_13519);
and U16132 (N_16132,N_14507,N_13675);
or U16133 (N_16133,N_15137,N_13831);
or U16134 (N_16134,N_14971,N_14406);
xor U16135 (N_16135,N_15426,N_15015);
and U16136 (N_16136,N_12955,N_13011);
xor U16137 (N_16137,N_12503,N_12340);
or U16138 (N_16138,N_14891,N_15025);
and U16139 (N_16139,N_14973,N_15190);
and U16140 (N_16140,N_13044,N_12039);
nand U16141 (N_16141,N_15172,N_13853);
and U16142 (N_16142,N_12343,N_13982);
and U16143 (N_16143,N_14161,N_15427);
nor U16144 (N_16144,N_12304,N_15504);
or U16145 (N_16145,N_15715,N_15053);
nor U16146 (N_16146,N_12279,N_14386);
nand U16147 (N_16147,N_13084,N_12019);
xor U16148 (N_16148,N_15682,N_13737);
or U16149 (N_16149,N_15291,N_12359);
and U16150 (N_16150,N_12283,N_13780);
nor U16151 (N_16151,N_12058,N_12150);
nand U16152 (N_16152,N_15582,N_14078);
or U16153 (N_16153,N_14555,N_12949);
xor U16154 (N_16154,N_15602,N_15898);
nor U16155 (N_16155,N_13316,N_13389);
or U16156 (N_16156,N_14430,N_14940);
or U16157 (N_16157,N_12777,N_13487);
or U16158 (N_16158,N_12325,N_15523);
nand U16159 (N_16159,N_14688,N_13056);
nand U16160 (N_16160,N_13817,N_15495);
xnor U16161 (N_16161,N_14323,N_15685);
nor U16162 (N_16162,N_15361,N_13095);
nor U16163 (N_16163,N_15922,N_12020);
nand U16164 (N_16164,N_12625,N_12254);
nor U16165 (N_16165,N_13354,N_14445);
nor U16166 (N_16166,N_13459,N_12008);
and U16167 (N_16167,N_13734,N_13387);
xnor U16168 (N_16168,N_12945,N_12824);
xor U16169 (N_16169,N_15534,N_15198);
and U16170 (N_16170,N_14290,N_13070);
nand U16171 (N_16171,N_15833,N_12792);
nand U16172 (N_16172,N_15413,N_12121);
and U16173 (N_16173,N_15084,N_13255);
and U16174 (N_16174,N_12339,N_12029);
xnor U16175 (N_16175,N_15745,N_13810);
nor U16176 (N_16176,N_12209,N_14121);
nand U16177 (N_16177,N_15932,N_14586);
and U16178 (N_16178,N_13673,N_12377);
or U16179 (N_16179,N_13979,N_15722);
nand U16180 (N_16180,N_14652,N_14746);
or U16181 (N_16181,N_14527,N_15440);
or U16182 (N_16182,N_13401,N_13561);
nor U16183 (N_16183,N_12663,N_15093);
nor U16184 (N_16184,N_14191,N_12280);
nor U16185 (N_16185,N_14342,N_12816);
nand U16186 (N_16186,N_15527,N_12373);
nand U16187 (N_16187,N_12232,N_15650);
or U16188 (N_16188,N_15985,N_15970);
and U16189 (N_16189,N_12302,N_15532);
nor U16190 (N_16190,N_14607,N_15799);
and U16191 (N_16191,N_12726,N_13426);
nor U16192 (N_16192,N_12316,N_14938);
and U16193 (N_16193,N_14013,N_13788);
xnor U16194 (N_16194,N_14431,N_12502);
nor U16195 (N_16195,N_15329,N_14307);
nor U16196 (N_16196,N_13990,N_15631);
nand U16197 (N_16197,N_15748,N_15664);
or U16198 (N_16198,N_12174,N_14020);
and U16199 (N_16199,N_13125,N_13048);
and U16200 (N_16200,N_15987,N_15537);
and U16201 (N_16201,N_14043,N_13482);
and U16202 (N_16202,N_13740,N_12970);
xor U16203 (N_16203,N_15013,N_12832);
nor U16204 (N_16204,N_15760,N_15934);
or U16205 (N_16205,N_13073,N_13230);
nand U16206 (N_16206,N_12661,N_14250);
nand U16207 (N_16207,N_15859,N_12540);
and U16208 (N_16208,N_13367,N_13716);
nand U16209 (N_16209,N_13888,N_14218);
xor U16210 (N_16210,N_13832,N_15316);
nand U16211 (N_16211,N_14985,N_13495);
and U16212 (N_16212,N_13914,N_13368);
xnor U16213 (N_16213,N_13119,N_12443);
and U16214 (N_16214,N_13712,N_12840);
and U16215 (N_16215,N_14117,N_12672);
nor U16216 (N_16216,N_15207,N_13065);
and U16217 (N_16217,N_12025,N_13785);
nand U16218 (N_16218,N_14488,N_14443);
or U16219 (N_16219,N_13775,N_13568);
nor U16220 (N_16220,N_14885,N_12846);
nand U16221 (N_16221,N_15921,N_12126);
and U16222 (N_16222,N_15955,N_12854);
or U16223 (N_16223,N_12426,N_13315);
and U16224 (N_16224,N_15118,N_14105);
nor U16225 (N_16225,N_13042,N_12628);
nor U16226 (N_16226,N_15119,N_12896);
and U16227 (N_16227,N_13657,N_14756);
and U16228 (N_16228,N_13098,N_12251);
or U16229 (N_16229,N_14860,N_15385);
and U16230 (N_16230,N_15502,N_12235);
nand U16231 (N_16231,N_12826,N_15304);
and U16232 (N_16232,N_13967,N_12394);
and U16233 (N_16233,N_12624,N_14673);
xnor U16234 (N_16234,N_13309,N_15345);
nand U16235 (N_16235,N_15468,N_15873);
nand U16236 (N_16236,N_12000,N_13542);
nor U16237 (N_16237,N_15910,N_15477);
or U16238 (N_16238,N_13857,N_15470);
or U16239 (N_16239,N_15402,N_13878);
nor U16240 (N_16240,N_13225,N_12587);
or U16241 (N_16241,N_12759,N_14981);
and U16242 (N_16242,N_12267,N_14948);
and U16243 (N_16243,N_14887,N_14919);
nand U16244 (N_16244,N_13620,N_13923);
nor U16245 (N_16245,N_12244,N_14411);
and U16246 (N_16246,N_12644,N_12130);
nor U16247 (N_16247,N_15714,N_13346);
nand U16248 (N_16248,N_13450,N_12033);
and U16249 (N_16249,N_15798,N_12925);
and U16250 (N_16250,N_13644,N_15743);
nand U16251 (N_16251,N_14438,N_14539);
nor U16252 (N_16252,N_13304,N_14720);
and U16253 (N_16253,N_14205,N_14764);
or U16254 (N_16254,N_14790,N_14683);
and U16255 (N_16255,N_14520,N_12233);
and U16256 (N_16256,N_15016,N_15450);
or U16257 (N_16257,N_12013,N_12987);
nand U16258 (N_16258,N_14134,N_14487);
xnor U16259 (N_16259,N_14045,N_15615);
or U16260 (N_16260,N_12207,N_13451);
and U16261 (N_16261,N_12372,N_14845);
or U16262 (N_16262,N_14352,N_12833);
nor U16263 (N_16263,N_12689,N_14553);
and U16264 (N_16264,N_13475,N_12484);
xnor U16265 (N_16265,N_13985,N_12711);
nor U16266 (N_16266,N_14559,N_15763);
or U16267 (N_16267,N_12049,N_15456);
xor U16268 (N_16268,N_15771,N_13611);
or U16269 (N_16269,N_12533,N_14881);
nand U16270 (N_16270,N_14613,N_15135);
nand U16271 (N_16271,N_12708,N_12415);
or U16272 (N_16272,N_12481,N_13366);
nor U16273 (N_16273,N_14747,N_14094);
nor U16274 (N_16274,N_13267,N_13896);
or U16275 (N_16275,N_15768,N_14861);
and U16276 (N_16276,N_12388,N_14030);
nand U16277 (N_16277,N_13358,N_15436);
nand U16278 (N_16278,N_15073,N_14497);
nand U16279 (N_16279,N_12868,N_12613);
xnor U16280 (N_16280,N_14057,N_12056);
nor U16281 (N_16281,N_15222,N_14532);
or U16282 (N_16282,N_12307,N_13922);
nand U16283 (N_16283,N_12616,N_12082);
xor U16284 (N_16284,N_12798,N_12715);
and U16285 (N_16285,N_14783,N_13241);
and U16286 (N_16286,N_14970,N_13508);
nand U16287 (N_16287,N_13235,N_15454);
nand U16288 (N_16288,N_15759,N_15824);
or U16289 (N_16289,N_14461,N_14003);
and U16290 (N_16290,N_15072,N_14318);
nand U16291 (N_16291,N_12248,N_12734);
nor U16292 (N_16292,N_14063,N_13308);
nor U16293 (N_16293,N_12924,N_12632);
nand U16294 (N_16294,N_15366,N_13800);
xnor U16295 (N_16295,N_13086,N_14015);
nand U16296 (N_16296,N_15218,N_14401);
nor U16297 (N_16297,N_14339,N_13666);
or U16298 (N_16298,N_13584,N_14047);
and U16299 (N_16299,N_13172,N_15183);
and U16300 (N_16300,N_13162,N_13528);
and U16301 (N_16301,N_13184,N_14362);
and U16302 (N_16302,N_12599,N_12173);
or U16303 (N_16303,N_13176,N_12653);
nor U16304 (N_16304,N_15707,N_15314);
nand U16305 (N_16305,N_13477,N_12457);
nor U16306 (N_16306,N_13069,N_14953);
nand U16307 (N_16307,N_13074,N_14841);
nand U16308 (N_16308,N_13695,N_15278);
xor U16309 (N_16309,N_15524,N_13112);
and U16310 (N_16310,N_12167,N_14229);
and U16311 (N_16311,N_15895,N_15827);
xor U16312 (N_16312,N_15837,N_13471);
nor U16313 (N_16313,N_14065,N_12112);
or U16314 (N_16314,N_14468,N_15288);
nand U16315 (N_16315,N_15540,N_13952);
xnor U16316 (N_16316,N_12169,N_14457);
nand U16317 (N_16317,N_14615,N_14701);
nor U16318 (N_16318,N_12386,N_13362);
and U16319 (N_16319,N_13855,N_12131);
or U16320 (N_16320,N_12630,N_15121);
xor U16321 (N_16321,N_15592,N_12581);
nand U16322 (N_16322,N_12471,N_12664);
nor U16323 (N_16323,N_14090,N_13469);
and U16324 (N_16324,N_14363,N_12212);
nor U16325 (N_16325,N_13732,N_15575);
and U16326 (N_16326,N_15744,N_14622);
nor U16327 (N_16327,N_13156,N_14834);
nand U16328 (N_16328,N_13493,N_15560);
and U16329 (N_16329,N_12706,N_12894);
and U16330 (N_16330,N_13433,N_15251);
nand U16331 (N_16331,N_13283,N_12852);
and U16332 (N_16332,N_13747,N_13147);
nand U16333 (N_16333,N_13333,N_15716);
or U16334 (N_16334,N_12439,N_13852);
or U16335 (N_16335,N_15579,N_12515);
nor U16336 (N_16336,N_15099,N_15122);
or U16337 (N_16337,N_12809,N_12695);
nor U16338 (N_16338,N_12477,N_13399);
xor U16339 (N_16339,N_15812,N_12768);
nor U16340 (N_16340,N_14122,N_15514);
nor U16341 (N_16341,N_14482,N_13295);
or U16342 (N_16342,N_14904,N_15293);
and U16343 (N_16343,N_14112,N_12189);
or U16344 (N_16344,N_12018,N_14330);
xnor U16345 (N_16345,N_14071,N_13105);
nor U16346 (N_16346,N_12686,N_13870);
nor U16347 (N_16347,N_13355,N_14710);
nor U16348 (N_16348,N_13205,N_12047);
and U16349 (N_16349,N_15253,N_12272);
nand U16350 (N_16350,N_14163,N_13751);
and U16351 (N_16351,N_13563,N_14794);
and U16352 (N_16352,N_14313,N_14998);
nand U16353 (N_16353,N_15811,N_15881);
nand U16354 (N_16354,N_12195,N_13894);
nor U16355 (N_16355,N_12867,N_12142);
or U16356 (N_16356,N_13610,N_13543);
nor U16357 (N_16357,N_13946,N_15506);
and U16358 (N_16358,N_14762,N_12269);
nor U16359 (N_16359,N_12276,N_13876);
and U16360 (N_16360,N_15012,N_14890);
and U16361 (N_16361,N_14140,N_12005);
and U16362 (N_16362,N_14875,N_12512);
or U16363 (N_16363,N_15313,N_13758);
nand U16364 (N_16364,N_14923,N_15545);
nand U16365 (N_16365,N_15324,N_14317);
nand U16366 (N_16366,N_14606,N_14751);
and U16367 (N_16367,N_12766,N_13204);
nand U16368 (N_16368,N_14976,N_14242);
and U16369 (N_16369,N_15149,N_15629);
or U16370 (N_16370,N_15216,N_15416);
and U16371 (N_16371,N_15045,N_15286);
xor U16372 (N_16372,N_15177,N_14656);
or U16373 (N_16373,N_14262,N_15212);
nand U16374 (N_16374,N_14634,N_13614);
nand U16375 (N_16375,N_12094,N_14789);
xnor U16376 (N_16376,N_13167,N_14035);
nand U16377 (N_16377,N_15723,N_12680);
and U16378 (N_16378,N_13208,N_14618);
and U16379 (N_16379,N_13660,N_12764);
and U16380 (N_16380,N_12323,N_12348);
or U16381 (N_16381,N_15694,N_15719);
or U16382 (N_16382,N_14395,N_12658);
nand U16383 (N_16383,N_15501,N_13847);
xor U16384 (N_16384,N_12619,N_14434);
nand U16385 (N_16385,N_15642,N_13639);
and U16386 (N_16386,N_12717,N_13199);
nor U16387 (N_16387,N_12836,N_12134);
or U16388 (N_16388,N_12181,N_14966);
or U16389 (N_16389,N_14770,N_15322);
or U16390 (N_16390,N_12057,N_13298);
nor U16391 (N_16391,N_12983,N_14547);
nor U16392 (N_16392,N_15163,N_14824);
xnor U16393 (N_16393,N_14611,N_13300);
nor U16394 (N_16394,N_12163,N_13158);
nand U16395 (N_16395,N_13343,N_13812);
nor U16396 (N_16396,N_12137,N_15732);
and U16397 (N_16397,N_14076,N_13571);
and U16398 (N_16398,N_14235,N_13574);
and U16399 (N_16399,N_13642,N_15011);
and U16400 (N_16400,N_15425,N_12501);
or U16401 (N_16401,N_15756,N_13375);
nor U16402 (N_16402,N_13748,N_14712);
and U16403 (N_16403,N_13776,N_14941);
nor U16404 (N_16404,N_13247,N_14695);
nor U16405 (N_16405,N_14299,N_13207);
xor U16406 (N_16406,N_12907,N_13129);
nand U16407 (N_16407,N_14475,N_15994);
and U16408 (N_16408,N_14148,N_13628);
nand U16409 (N_16409,N_14316,N_13828);
nor U16410 (N_16410,N_13622,N_13049);
nand U16411 (N_16411,N_14552,N_12575);
nand U16412 (N_16412,N_15917,N_12841);
or U16413 (N_16413,N_12469,N_14734);
xor U16414 (N_16414,N_15953,N_14055);
nand U16415 (N_16415,N_14172,N_13565);
and U16416 (N_16416,N_15776,N_15958);
nor U16417 (N_16417,N_15387,N_14802);
nand U16418 (N_16418,N_14835,N_14268);
xnor U16419 (N_16419,N_14538,N_13490);
or U16420 (N_16420,N_13834,N_12434);
nand U16421 (N_16421,N_12499,N_12723);
or U16422 (N_16422,N_14223,N_13792);
and U16423 (N_16423,N_12456,N_14964);
nor U16424 (N_16424,N_15371,N_12417);
or U16425 (N_16425,N_13711,N_15036);
xor U16426 (N_16426,N_15459,N_15059);
nor U16427 (N_16427,N_15362,N_14576);
nor U16428 (N_16428,N_14369,N_15054);
and U16429 (N_16429,N_14375,N_14658);
nand U16430 (N_16430,N_14798,N_14501);
nand U16431 (N_16431,N_13517,N_15182);
or U16432 (N_16432,N_14558,N_12102);
nand U16433 (N_16433,N_13652,N_15938);
nor U16434 (N_16434,N_14533,N_15503);
xor U16435 (N_16435,N_12576,N_12548);
nor U16436 (N_16436,N_13567,N_12539);
or U16437 (N_16437,N_14895,N_12627);
nor U16438 (N_16438,N_13374,N_14907);
xnor U16439 (N_16439,N_14654,N_14455);
and U16440 (N_16440,N_14721,N_13050);
nor U16441 (N_16441,N_14777,N_12859);
or U16442 (N_16442,N_14597,N_13741);
xor U16443 (N_16443,N_13835,N_15185);
or U16444 (N_16444,N_12884,N_13953);
and U16445 (N_16445,N_12771,N_14208);
nor U16446 (N_16446,N_12569,N_14537);
or U16447 (N_16447,N_13601,N_15249);
nor U16448 (N_16448,N_13029,N_14510);
or U16449 (N_16449,N_12675,N_14529);
xnor U16450 (N_16450,N_15047,N_14944);
nor U16451 (N_16451,N_15050,N_12199);
nand U16452 (N_16452,N_15761,N_13186);
and U16453 (N_16453,N_14871,N_15197);
or U16454 (N_16454,N_13724,N_14489);
nand U16455 (N_16455,N_13645,N_12193);
and U16456 (N_16456,N_13276,N_15167);
nand U16457 (N_16457,N_15874,N_13873);
or U16458 (N_16458,N_12003,N_13015);
nor U16459 (N_16459,N_15193,N_12180);
or U16460 (N_16460,N_13417,N_14761);
nor U16461 (N_16461,N_15092,N_12525);
and U16462 (N_16462,N_14239,N_12291);
nand U16463 (N_16463,N_14681,N_14031);
nor U16464 (N_16464,N_12308,N_15107);
or U16465 (N_16465,N_15273,N_12785);
nor U16466 (N_16466,N_12293,N_13197);
xor U16467 (N_16467,N_15261,N_13903);
and U16468 (N_16468,N_12720,N_12522);
xor U16469 (N_16469,N_14398,N_15300);
nand U16470 (N_16470,N_14522,N_13576);
nor U16471 (N_16471,N_15990,N_12571);
nor U16472 (N_16472,N_13700,N_14864);
nand U16473 (N_16473,N_12911,N_14916);
nor U16474 (N_16474,N_13759,N_14484);
xnor U16475 (N_16475,N_13702,N_13955);
and U16476 (N_16476,N_14167,N_14034);
and U16477 (N_16477,N_12971,N_13845);
nand U16478 (N_16478,N_12772,N_12615);
and U16479 (N_16479,N_13089,N_13706);
or U16480 (N_16480,N_14120,N_13753);
xor U16481 (N_16481,N_15781,N_14820);
nand U16482 (N_16482,N_14856,N_12152);
and U16483 (N_16483,N_12787,N_15774);
xnor U16484 (N_16484,N_14580,N_12350);
or U16485 (N_16485,N_15378,N_12574);
or U16486 (N_16486,N_15680,N_13384);
xor U16487 (N_16487,N_12756,N_14414);
xnor U16488 (N_16488,N_13257,N_14292);
or U16489 (N_16489,N_15094,N_14174);
nor U16490 (N_16490,N_14946,N_15862);
and U16491 (N_16491,N_13285,N_14462);
nand U16492 (N_16492,N_13504,N_13397);
nor U16493 (N_16493,N_14346,N_14050);
or U16494 (N_16494,N_12744,N_12530);
nand U16495 (N_16495,N_14686,N_12881);
and U16496 (N_16496,N_14758,N_13575);
or U16497 (N_16497,N_13965,N_14089);
nor U16498 (N_16498,N_13104,N_12486);
xnor U16499 (N_16499,N_13604,N_12988);
nand U16500 (N_16500,N_15577,N_13400);
or U16501 (N_16501,N_15384,N_15208);
nor U16502 (N_16502,N_12682,N_12284);
or U16503 (N_16503,N_15255,N_13020);
nor U16504 (N_16504,N_12327,N_13807);
nor U16505 (N_16505,N_13558,N_13939);
nand U16506 (N_16506,N_12972,N_15389);
nor U16507 (N_16507,N_12968,N_12470);
nand U16508 (N_16508,N_15279,N_12423);
nand U16509 (N_16509,N_14809,N_13008);
xnor U16510 (N_16510,N_14236,N_13697);
xnor U16511 (N_16511,N_14165,N_14156);
or U16512 (N_16512,N_14499,N_15202);
nand U16513 (N_16513,N_13920,N_14295);
nor U16514 (N_16514,N_12805,N_15297);
nand U16515 (N_16515,N_14347,N_14225);
nand U16516 (N_16516,N_15347,N_14176);
nand U16517 (N_16517,N_15931,N_14743);
or U16518 (N_16518,N_13808,N_13088);
and U16519 (N_16519,N_13155,N_13228);
or U16520 (N_16520,N_14727,N_12538);
or U16521 (N_16521,N_14584,N_14275);
nand U16522 (N_16522,N_15554,N_15893);
nand U16523 (N_16523,N_15174,N_13037);
xor U16524 (N_16524,N_13330,N_12099);
or U16525 (N_16525,N_15754,N_14674);
or U16526 (N_16526,N_14526,N_14179);
xnor U16527 (N_16527,N_13299,N_14744);
nand U16528 (N_16528,N_12136,N_13826);
nor U16529 (N_16529,N_15486,N_12853);
or U16530 (N_16530,N_15949,N_15405);
or U16531 (N_16531,N_13829,N_15865);
or U16532 (N_16532,N_14209,N_12657);
and U16533 (N_16533,N_15057,N_15900);
or U16534 (N_16534,N_13071,N_14616);
and U16535 (N_16535,N_14415,N_15237);
xnor U16536 (N_16536,N_13391,N_14378);
and U16537 (N_16537,N_12239,N_13465);
nor U16538 (N_16538,N_15705,N_12356);
and U16539 (N_16539,N_12745,N_12401);
and U16540 (N_16540,N_13599,N_12464);
nand U16541 (N_16541,N_13183,N_13841);
nand U16542 (N_16542,N_14083,N_15129);
nand U16543 (N_16543,N_14367,N_12306);
nor U16544 (N_16544,N_13510,N_15688);
nor U16545 (N_16545,N_12138,N_14886);
nor U16546 (N_16546,N_15678,N_13927);
and U16547 (N_16547,N_12202,N_14138);
or U16548 (N_16548,N_13522,N_13177);
nor U16549 (N_16549,N_13342,N_12281);
nor U16550 (N_16550,N_12601,N_12273);
or U16551 (N_16551,N_14277,N_14354);
and U16552 (N_16552,N_12200,N_15959);
and U16553 (N_16553,N_14109,N_15843);
or U16554 (N_16554,N_14326,N_14577);
nand U16555 (N_16555,N_15930,N_12042);
or U16556 (N_16556,N_14393,N_15937);
nand U16557 (N_16557,N_14311,N_12436);
nor U16558 (N_16558,N_15956,N_12659);
or U16559 (N_16559,N_14548,N_13421);
and U16560 (N_16560,N_12879,N_13272);
and U16561 (N_16561,N_12608,N_15262);
nor U16562 (N_16562,N_15332,N_14635);
and U16563 (N_16563,N_12957,N_12724);
or U16564 (N_16564,N_13270,N_13485);
and U16565 (N_16565,N_14914,N_13704);
or U16566 (N_16566,N_12831,N_12880);
or U16567 (N_16567,N_13709,N_14857);
and U16568 (N_16568,N_12544,N_15909);
or U16569 (N_16569,N_13944,N_15860);
or U16570 (N_16570,N_15617,N_12980);
xor U16571 (N_16571,N_12595,N_15718);
xnor U16572 (N_16572,N_14838,N_15819);
nor U16573 (N_16573,N_12558,N_13555);
and U16574 (N_16574,N_13743,N_15147);
and U16575 (N_16575,N_15338,N_13670);
nand U16576 (N_16576,N_15055,N_12159);
or U16577 (N_16577,N_13356,N_13395);
and U16578 (N_16578,N_14717,N_15071);
nor U16579 (N_16579,N_13572,N_13902);
or U16580 (N_16580,N_12518,N_13223);
nor U16581 (N_16581,N_14100,N_15976);
and U16582 (N_16582,N_15896,N_15872);
xnor U16583 (N_16583,N_15281,N_12917);
and U16584 (N_16584,N_13244,N_12074);
and U16585 (N_16585,N_14160,N_13231);
and U16586 (N_16586,N_13160,N_15815);
xor U16587 (N_16587,N_15087,N_13925);
nor U16588 (N_16588,N_14578,N_12326);
nand U16589 (N_16589,N_12184,N_12799);
nand U16590 (N_16590,N_12905,N_15280);
and U16591 (N_16591,N_15919,N_15795);
nor U16592 (N_16592,N_13677,N_12355);
nand U16593 (N_16593,N_12384,N_14359);
nor U16594 (N_16594,N_13441,N_13000);
and U16595 (N_16595,N_12259,N_15328);
xnor U16596 (N_16596,N_12367,N_15525);
nand U16597 (N_16597,N_13679,N_12874);
and U16598 (N_16598,N_12270,N_12578);
nand U16599 (N_16599,N_14142,N_13004);
nor U16600 (N_16600,N_14322,N_13220);
nand U16601 (N_16601,N_15644,N_12151);
nor U16602 (N_16602,N_13765,N_12176);
and U16603 (N_16603,N_12298,N_14943);
xor U16604 (N_16604,N_12400,N_12730);
and U16605 (N_16605,N_15188,N_15801);
nor U16606 (N_16606,N_15116,N_14560);
xor U16607 (N_16607,N_12098,N_13691);
or U16608 (N_16608,N_13784,N_12618);
or U16609 (N_16609,N_12506,N_13600);
nor U16610 (N_16610,N_15376,N_15697);
xnor U16611 (N_16611,N_14787,N_12374);
xnor U16612 (N_16612,N_14563,N_13149);
nand U16613 (N_16613,N_14990,N_15947);
and U16614 (N_16614,N_15720,N_14801);
nand U16615 (N_16615,N_13822,N_12095);
nand U16616 (N_16616,N_15821,N_15248);
and U16617 (N_16617,N_12105,N_13719);
or U16618 (N_16618,N_13655,N_13797);
nor U16619 (N_16619,N_14425,N_15452);
or U16620 (N_16620,N_12566,N_15613);
and U16621 (N_16621,N_12260,N_12106);
and U16622 (N_16622,N_15493,N_13322);
xnor U16623 (N_16623,N_15713,N_15943);
or U16624 (N_16624,N_15306,N_12687);
xnor U16625 (N_16625,N_12246,N_13379);
nor U16626 (N_16626,N_13919,N_12243);
and U16627 (N_16627,N_13975,N_13376);
and U16628 (N_16628,N_15924,N_14131);
or U16629 (N_16629,N_12241,N_13334);
and U16630 (N_16630,N_13328,N_12902);
or U16631 (N_16631,N_14285,N_13138);
and U16632 (N_16632,N_14807,N_13884);
or U16633 (N_16633,N_14441,N_13991);
or U16634 (N_16634,N_14949,N_12592);
or U16635 (N_16635,N_15675,N_14894);
and U16636 (N_16636,N_13573,N_13659);
nor U16637 (N_16637,N_12662,N_12822);
nor U16638 (N_16638,N_13182,N_12203);
and U16639 (N_16639,N_15557,N_12310);
or U16640 (N_16640,N_15144,N_15153);
nor U16641 (N_16641,N_15136,N_12709);
nand U16642 (N_16642,N_14006,N_12190);
nor U16643 (N_16643,N_13752,N_12110);
or U16644 (N_16644,N_13325,N_13492);
or U16645 (N_16645,N_12315,N_14389);
and U16646 (N_16646,N_15853,N_14227);
or U16647 (N_16647,N_14240,N_15323);
nor U16648 (N_16648,N_15727,N_12256);
or U16649 (N_16649,N_14152,N_12414);
or U16650 (N_16650,N_13116,N_12346);
or U16651 (N_16651,N_12514,N_13305);
xnor U16652 (N_16652,N_13214,N_14588);
nand U16653 (N_16653,N_15844,N_14741);
nand U16654 (N_16654,N_14004,N_12432);
or U16655 (N_16655,N_14099,N_14655);
or U16656 (N_16656,N_15739,N_15660);
or U16657 (N_16657,N_14207,N_15049);
and U16658 (N_16658,N_13022,N_12153);
and U16659 (N_16659,N_13338,N_14827);
nor U16660 (N_16660,N_15246,N_13764);
and U16661 (N_16661,N_13908,N_15757);
nand U16662 (N_16662,N_14780,N_13034);
nor U16663 (N_16663,N_13468,N_15848);
nor U16664 (N_16664,N_13916,N_12851);
nor U16665 (N_16665,N_13032,N_14687);
nand U16666 (N_16666,N_15221,N_13547);
nor U16667 (N_16667,N_12551,N_12990);
and U16668 (N_16668,N_14258,N_14699);
and U16669 (N_16669,N_13148,N_15390);
xnor U16670 (N_16670,N_14079,N_12487);
and U16671 (N_16671,N_15335,N_13431);
nor U16672 (N_16672,N_14102,N_12966);
or U16673 (N_16673,N_15892,N_13624);
or U16674 (N_16674,N_12650,N_13667);
nand U16675 (N_16675,N_13803,N_12678);
and U16676 (N_16676,N_15151,N_15806);
xnor U16677 (N_16677,N_13968,N_12228);
xor U16678 (N_16678,N_14582,N_15349);
xnor U16679 (N_16679,N_14596,N_13195);
and U16680 (N_16680,N_14778,N_13236);
nand U16681 (N_16681,N_15551,N_15858);
and U16682 (N_16682,N_15992,N_13637);
nand U16683 (N_16683,N_14848,N_12758);
or U16684 (N_16684,N_14974,N_12763);
nand U16685 (N_16685,N_15126,N_15584);
or U16686 (N_16686,N_14568,N_14512);
or U16687 (N_16687,N_13647,N_14093);
nand U16688 (N_16688,N_13259,N_13382);
and U16689 (N_16689,N_12453,N_15006);
and U16690 (N_16690,N_13860,N_12375);
nor U16691 (N_16691,N_15555,N_14763);
and U16692 (N_16692,N_14486,N_13549);
nor U16693 (N_16693,N_13641,N_12148);
xor U16694 (N_16694,N_14939,N_14594);
or U16695 (N_16695,N_15111,N_12883);
and U16696 (N_16696,N_13609,N_14779);
and U16697 (N_16697,N_12864,N_13595);
nor U16698 (N_16698,N_12075,N_14182);
and U16699 (N_16699,N_13006,N_14994);
nand U16700 (N_16700,N_15232,N_15341);
nor U16701 (N_16701,N_15564,N_14930);
xor U16702 (N_16702,N_14310,N_14950);
nand U16703 (N_16703,N_15864,N_15175);
nand U16704 (N_16704,N_13363,N_12511);
nand U16705 (N_16705,N_12774,N_14186);
and U16706 (N_16706,N_15861,N_14169);
nand U16707 (N_16707,N_15673,N_15483);
nand U16708 (N_16708,N_14280,N_13181);
nand U16709 (N_16709,N_14194,N_15003);
nor U16710 (N_16710,N_15778,N_15832);
nor U16711 (N_16711,N_13560,N_15269);
nand U16712 (N_16712,N_14832,N_13940);
and U16713 (N_16713,N_14682,N_15689);
or U16714 (N_16714,N_14184,N_15033);
nor U16715 (N_16715,N_14056,N_14054);
nor U16716 (N_16716,N_12030,N_12942);
and U16717 (N_16717,N_14496,N_14115);
nor U16718 (N_16718,N_12264,N_14958);
nor U16719 (N_16719,N_15725,N_14924);
and U16720 (N_16720,N_13613,N_15765);
nand U16721 (N_16721,N_14972,N_12046);
nor U16722 (N_16722,N_14929,N_15666);
and U16723 (N_16723,N_12416,N_13907);
nor U16724 (N_16724,N_13414,N_15481);
or U16725 (N_16725,N_12904,N_12975);
nand U16726 (N_16726,N_15823,N_13271);
nor U16727 (N_16727,N_12685,N_14517);
nor U16728 (N_16728,N_14977,N_14980);
or U16729 (N_16729,N_13344,N_15196);
or U16730 (N_16730,N_14637,N_14357);
and U16731 (N_16731,N_14201,N_12223);
or U16732 (N_16732,N_13128,N_15863);
nand U16733 (N_16733,N_14139,N_13978);
or U16734 (N_16734,N_13481,N_13615);
or U16735 (N_16735,N_15260,N_13838);
nand U16736 (N_16736,N_14458,N_14995);
and U16737 (N_16737,N_13851,N_13754);
nor U16738 (N_16738,N_12081,N_15636);
nand U16739 (N_16739,N_15576,N_12710);
nor U16740 (N_16740,N_12089,N_14206);
and U16741 (N_16741,N_13472,N_13093);
or U16742 (N_16742,N_15406,N_12257);
and U16743 (N_16743,N_15736,N_13891);
and U16744 (N_16744,N_15158,N_12914);
or U16745 (N_16745,N_14245,N_13061);
or U16746 (N_16746,N_12536,N_14988);
nand U16747 (N_16747,N_13900,N_14101);
xnor U16748 (N_16748,N_13062,N_15508);
xor U16749 (N_16749,N_15690,N_14525);
and U16750 (N_16750,N_13635,N_12078);
or U16751 (N_16751,N_15339,N_12626);
and U16752 (N_16752,N_14111,N_12069);
or U16753 (N_16753,N_14309,N_12336);
nand U16754 (N_16754,N_12036,N_12253);
or U16755 (N_16755,N_12337,N_14060);
nor U16756 (N_16756,N_13405,N_15140);
xor U16757 (N_16757,N_14439,N_14621);
nand U16758 (N_16758,N_12997,N_14450);
or U16759 (N_16759,N_15787,N_13879);
or U16760 (N_16760,N_15531,N_13885);
nand U16761 (N_16761,N_13514,N_15672);
and U16762 (N_16762,N_12998,N_13288);
and U16763 (N_16763,N_13324,N_15046);
nor U16764 (N_16764,N_13320,N_12568);
nor U16765 (N_16765,N_12964,N_13730);
or U16766 (N_16766,N_14321,N_14523);
xor U16767 (N_16767,N_13131,N_15465);
xor U16768 (N_16768,N_13312,N_12398);
nand U16769 (N_16769,N_13524,N_15078);
nor U16770 (N_16770,N_15373,N_14011);
nand U16771 (N_16771,N_12397,N_14978);
nand U16772 (N_16772,N_14272,N_14987);
and U16773 (N_16773,N_15106,N_15621);
nor U16774 (N_16774,N_12231,N_14693);
and U16775 (N_16775,N_14253,N_12140);
nor U16776 (N_16776,N_13013,N_14865);
nor U16777 (N_16777,N_15777,N_13250);
and U16778 (N_16778,N_12807,N_15840);
and U16779 (N_16779,N_13554,N_14951);
nand U16780 (N_16780,N_12219,N_15042);
or U16781 (N_16781,N_14639,N_14937);
xor U16782 (N_16782,N_15512,N_13263);
nand U16783 (N_16783,N_14166,N_15822);
xor U16784 (N_16784,N_12504,N_13219);
nand U16785 (N_16785,N_14446,N_13703);
and U16786 (N_16786,N_14786,N_13654);
and U16787 (N_16787,N_15645,N_13031);
or U16788 (N_16788,N_15319,N_15258);
nand U16789 (N_16789,N_14859,N_13180);
xnor U16790 (N_16790,N_14025,N_15159);
nor U16791 (N_16791,N_15845,N_15496);
nor U16792 (N_16792,N_13996,N_14561);
and U16793 (N_16793,N_13947,N_15234);
nand U16794 (N_16794,N_14470,N_14800);
or U16795 (N_16795,N_12370,N_13662);
nor U16796 (N_16796,N_13323,N_15810);
nor U16797 (N_16797,N_14703,N_12396);
nand U16798 (N_16798,N_12262,N_15307);
nor U16799 (N_16799,N_14294,N_12292);
and U16800 (N_16800,N_12927,N_15458);
or U16801 (N_16801,N_15746,N_15355);
nor U16802 (N_16802,N_13597,N_15034);
nor U16803 (N_16803,N_15614,N_15948);
nor U16804 (N_16804,N_13253,N_13217);
or U16805 (N_16805,N_12585,N_14107);
or U16806 (N_16806,N_15975,N_15847);
nor U16807 (N_16807,N_13453,N_13824);
nor U16808 (N_16808,N_12072,N_13473);
nor U16809 (N_16809,N_14405,N_12543);
and U16810 (N_16810,N_13969,N_12288);
nand U16811 (N_16811,N_13559,N_15001);
nand U16812 (N_16812,N_14151,N_15826);
nor U16813 (N_16813,N_13889,N_15905);
and U16814 (N_16814,N_15926,N_12813);
nand U16815 (N_16815,N_12478,N_14417);
nor U16816 (N_16816,N_14797,N_14234);
or U16817 (N_16817,N_12698,N_12580);
and U16818 (N_16818,N_14659,N_13261);
or U16819 (N_16819,N_15331,N_14391);
nor U16820 (N_16820,N_13566,N_13513);
or U16821 (N_16821,N_12931,N_13237);
nor U16822 (N_16822,N_12035,N_15648);
and U16823 (N_16823,N_14360,N_14750);
nand U16824 (N_16824,N_15543,N_13681);
and U16825 (N_16825,N_15572,N_14181);
nor U16826 (N_16826,N_12351,N_12338);
xnor U16827 (N_16827,N_15788,N_13790);
or U16828 (N_16828,N_14231,N_14402);
and U16829 (N_16829,N_14469,N_13209);
nor U16830 (N_16830,N_12043,N_14684);
nand U16831 (N_16831,N_13766,N_13386);
and U16832 (N_16832,N_14147,N_15687);
nand U16833 (N_16833,N_12225,N_13142);
or U16834 (N_16834,N_12527,N_12050);
nor U16835 (N_16835,N_13003,N_12860);
nand U16836 (N_16836,N_14975,N_14620);
nor U16837 (N_16837,N_15899,N_12915);
and U16838 (N_16838,N_13778,N_12007);
nand U16839 (N_16839,N_12783,N_13762);
nor U16840 (N_16840,N_15231,N_13266);
xor U16841 (N_16841,N_12299,N_14766);
nand U16842 (N_16842,N_12586,N_12594);
or U16843 (N_16843,N_14084,N_12305);
and U16844 (N_16844,N_13525,N_14226);
or U16845 (N_16845,N_15633,N_12642);
or U16846 (N_16846,N_13114,N_14626);
or U16847 (N_16847,N_15391,N_15139);
and U16848 (N_16848,N_13424,N_15305);
nor U16849 (N_16849,N_13122,N_15079);
nor U16850 (N_16850,N_12940,N_12087);
nand U16851 (N_16851,N_12621,N_12165);
nand U16852 (N_16852,N_14614,N_12119);
nor U16853 (N_16853,N_15728,N_15891);
or U16854 (N_16854,N_13570,N_14708);
nand U16855 (N_16855,N_14211,N_14314);
nand U16856 (N_16856,N_14212,N_13749);
nor U16857 (N_16857,N_14989,N_15961);
or U16858 (N_16858,N_14513,N_12275);
nor U16859 (N_16859,N_14024,N_14095);
nor U16860 (N_16860,N_15603,N_13699);
or U16861 (N_16861,N_12395,N_13768);
or U16862 (N_16862,N_13592,N_12969);
nor U16863 (N_16863,N_14947,N_15276);
and U16864 (N_16864,N_15752,N_15243);
nand U16865 (N_16865,N_14889,N_15369);
nor U16866 (N_16866,N_15354,N_15372);
or U16867 (N_16867,N_12839,N_13625);
nand U16868 (N_16868,N_13159,N_15474);
xor U16869 (N_16869,N_13992,N_13552);
nand U16870 (N_16870,N_15789,N_15651);
nor U16871 (N_16871,N_12572,N_14265);
and U16872 (N_16872,N_12967,N_12229);
nand U16873 (N_16873,N_14017,N_15802);
nor U16874 (N_16874,N_15161,N_15095);
nor U16875 (N_16875,N_15626,N_15008);
nor U16876 (N_16876,N_15939,N_15377);
or U16877 (N_16877,N_12038,N_12999);
and U16878 (N_16878,N_12820,N_14279);
and U16879 (N_16879,N_12510,N_15952);
nand U16880 (N_16880,N_14286,N_13480);
xnor U16881 (N_16881,N_14738,N_12977);
nand U16882 (N_16882,N_14905,N_15710);
nor U16883 (N_16883,N_15076,N_13819);
nor U16884 (N_16884,N_13151,N_12696);
xor U16885 (N_16885,N_15461,N_13520);
nor U16886 (N_16886,N_12297,N_13193);
nand U16887 (N_16887,N_15404,N_12371);
xor U16888 (N_16888,N_13360,N_15984);
nand U16889 (N_16889,N_15967,N_13117);
or U16890 (N_16890,N_14130,N_13023);
xor U16891 (N_16891,N_13370,N_14609);
and U16892 (N_16892,N_12438,N_14704);
or U16893 (N_16893,N_12129,N_14504);
nand U16894 (N_16894,N_14189,N_15692);
and U16895 (N_16895,N_14759,N_14202);
nor U16896 (N_16896,N_15233,N_13763);
xnor U16897 (N_16897,N_13229,N_14350);
or U16898 (N_16898,N_12472,N_12437);
nor U16899 (N_16899,N_13314,N_13989);
and U16900 (N_16900,N_14773,N_12196);
nor U16901 (N_16901,N_12321,N_12090);
nand U16902 (N_16902,N_13658,N_15721);
xnor U16903 (N_16903,N_13456,N_15769);
nor U16904 (N_16904,N_15211,N_13883);
nand U16905 (N_16905,N_15571,N_13959);
nor U16906 (N_16906,N_14514,N_13458);
or U16907 (N_16907,N_13856,N_14287);
and U16908 (N_16908,N_14157,N_13745);
nor U16909 (N_16909,N_12077,N_14073);
nor U16910 (N_16910,N_15770,N_15683);
and U16911 (N_16911,N_13491,N_14435);
xor U16912 (N_16912,N_15263,N_15418);
and U16913 (N_16913,N_14822,N_12023);
nand U16914 (N_16914,N_14961,N_14534);
nand U16915 (N_16915,N_13791,N_12561);
or U16916 (N_16916,N_14288,N_12886);
nor U16917 (N_16917,N_15392,N_13804);
or U16918 (N_16918,N_15374,N_13895);
xnor U16919 (N_16919,N_13738,N_12221);
and U16920 (N_16920,N_14388,N_14906);
nor U16921 (N_16921,N_14075,N_13077);
nand U16922 (N_16922,N_15605,N_15589);
or U16923 (N_16923,N_12690,N_13041);
or U16924 (N_16924,N_14381,N_15235);
nand U16925 (N_16925,N_13971,N_13935);
nand U16926 (N_16926,N_12409,N_14249);
and U16927 (N_16927,N_12598,N_15993);
and U16928 (N_16928,N_14546,N_14291);
nor U16929 (N_16929,N_12700,N_13735);
nor U16930 (N_16930,N_12076,N_12422);
nor U16931 (N_16931,N_15004,N_12494);
or U16932 (N_16932,N_13012,N_14500);
and U16933 (N_16933,N_13787,N_15060);
or U16934 (N_16934,N_14690,N_13260);
and U16935 (N_16935,N_15447,N_12428);
or U16936 (N_16936,N_13958,N_14813);
nor U16937 (N_16937,N_13218,N_15649);
or U16938 (N_16938,N_15659,N_13755);
nor U16939 (N_16939,N_15301,N_13173);
or U16940 (N_16940,N_13340,N_15654);
and U16941 (N_16941,N_14198,N_12435);
nor U16942 (N_16942,N_15299,N_15620);
or U16943 (N_16943,N_13430,N_12762);
or U16944 (N_16944,N_15733,N_13633);
and U16945 (N_16945,N_12145,N_12012);
nor U16946 (N_16946,N_12995,N_12402);
and U16947 (N_16947,N_15067,N_14053);
and U16948 (N_16948,N_12888,N_14641);
and U16949 (N_16949,N_13501,N_13603);
or U16950 (N_16950,N_15275,N_12086);
or U16951 (N_16951,N_15292,N_15382);
nand U16952 (N_16952,N_13523,N_15676);
or U16953 (N_16953,N_13974,N_13121);
or U16954 (N_16954,N_15138,N_14549);
nand U16955 (N_16955,N_14082,N_15887);
nand U16956 (N_16956,N_12748,N_13999);
and U16957 (N_16957,N_13779,N_14806);
nor U16958 (N_16958,N_12286,N_12017);
nor U16959 (N_16959,N_15424,N_15423);
or U16960 (N_16960,N_14705,N_14038);
nor U16961 (N_16961,N_15412,N_14066);
or U16962 (N_16962,N_15110,N_14028);
nand U16963 (N_16963,N_12899,N_15500);
and U16964 (N_16964,N_12780,N_15400);
and U16965 (N_16965,N_15679,N_13051);
nand U16966 (N_16966,N_13111,N_12564);
or U16967 (N_16967,N_14404,N_13854);
and U16968 (N_16968,N_13447,N_13987);
nor U16969 (N_16969,N_12022,N_13474);
or U16970 (N_16970,N_12817,N_13187);
nand U16971 (N_16971,N_15708,N_15181);
nand U16972 (N_16972,N_14453,N_12669);
and U16973 (N_16973,N_13731,N_15228);
nor U16974 (N_16974,N_14793,N_12679);
and U16975 (N_16975,N_12216,N_13054);
xnor U16976 (N_16976,N_14349,N_12107);
or U16977 (N_16977,N_14524,N_14436);
nand U16978 (N_16978,N_14593,N_13868);
and U16979 (N_16979,N_14049,N_13157);
nor U16980 (N_16980,N_12111,N_15134);
nand U16981 (N_16981,N_15187,N_15108);
and U16982 (N_16982,N_15435,N_15031);
or U16983 (N_16983,N_12198,N_13385);
or U16984 (N_16984,N_15010,N_14213);
nand U16985 (N_16985,N_15978,N_14858);
nor U16986 (N_16986,N_12289,N_13396);
nor U16987 (N_16987,N_12559,N_12194);
and U16988 (N_16988,N_13918,N_12429);
nor U16989 (N_16989,N_15020,N_12683);
or U16990 (N_16990,N_14863,N_15996);
nand U16991 (N_16991,N_15310,N_15505);
nand U16992 (N_16992,N_12932,N_14190);
and U16993 (N_16993,N_12922,N_15935);
or U16994 (N_16994,N_14237,N_13039);
and U16995 (N_16995,N_14259,N_15914);
and U16996 (N_16996,N_15698,N_13143);
and U16997 (N_16997,N_14707,N_12164);
and U16998 (N_16998,N_15102,N_14324);
nor U16999 (N_16999,N_14816,N_12973);
nand U17000 (N_17000,N_13551,N_15681);
and U17001 (N_17001,N_14926,N_15820);
or U17002 (N_17002,N_12300,N_15065);
or U17003 (N_17003,N_12334,N_15903);
nor U17004 (N_17004,N_14805,N_14372);
xor U17005 (N_17005,N_15925,N_15816);
nand U17006 (N_17006,N_12441,N_12458);
and U17007 (N_17007,N_13213,N_13983);
nand U17008 (N_17008,N_13720,N_15206);
nand U17009 (N_17009,N_14302,N_13326);
nand U17010 (N_17010,N_14642,N_14168);
nor U17011 (N_17011,N_13781,N_12197);
and U17012 (N_17012,N_12125,N_14289);
or U17013 (N_17013,N_15308,N_12926);
or U17014 (N_17014,N_12363,N_13877);
or U17015 (N_17015,N_13943,N_12555);
nand U17016 (N_17016,N_14348,N_15561);
nor U17017 (N_17017,N_13688,N_14046);
nor U17018 (N_17018,N_15849,N_12287);
xnor U17019 (N_17019,N_14217,N_14830);
or U17020 (N_17020,N_15342,N_14241);
xnor U17021 (N_17021,N_15825,N_13349);
and U17022 (N_17022,N_13931,N_14516);
and U17023 (N_17023,N_12133,N_12002);
and U17024 (N_17024,N_15526,N_15888);
nor U17025 (N_17025,N_12448,N_12250);
xor U17026 (N_17026,N_14451,N_13694);
and U17027 (N_17027,N_13818,N_14377);
nor U17028 (N_17028,N_12330,N_15125);
nand U17029 (N_17029,N_14833,N_14150);
nand U17030 (N_17030,N_14014,N_12893);
nand U17031 (N_17031,N_14001,N_15453);
or U17032 (N_17032,N_15539,N_12366);
xor U17033 (N_17033,N_15213,N_15180);
and U17034 (N_17034,N_14467,N_15009);
nor U17035 (N_17035,N_15062,N_13972);
nand U17036 (N_17036,N_14772,N_13535);
nor U17037 (N_17037,N_14962,N_15618);
nor U17038 (N_17038,N_12113,N_14672);
nor U17039 (N_17039,N_12093,N_14776);
nand U17040 (N_17040,N_15209,N_14037);
nor U17041 (N_17041,N_12143,N_13245);
nor U17042 (N_17042,N_13040,N_15550);
or U17043 (N_17043,N_15030,N_12793);
nand U17044 (N_17044,N_13976,N_13692);
nor U17045 (N_17045,N_14087,N_13248);
and U17046 (N_17046,N_12420,N_14269);
and U17047 (N_17047,N_13678,N_13258);
nor U17048 (N_17048,N_15241,N_13707);
nor U17049 (N_17049,N_12166,N_15380);
and U17050 (N_17050,N_14880,N_14494);
nor U17051 (N_17051,N_14917,N_15085);
nor U17052 (N_17052,N_13306,N_13500);
nand U17053 (N_17053,N_14498,N_15989);
nor U17054 (N_17054,N_14154,N_14146);
nor U17055 (N_17055,N_12892,N_15652);
and U17056 (N_17056,N_14301,N_15186);
nor U17057 (N_17057,N_14210,N_13052);
or U17058 (N_17058,N_14808,N_15346);
and U17059 (N_17059,N_13419,N_15334);
nand U17060 (N_17060,N_14042,N_12204);
or U17061 (N_17061,N_12838,N_15473);
nor U17062 (N_17062,N_14051,N_13185);
nand U17063 (N_17063,N_12645,N_13708);
nor U17064 (N_17064,N_14645,N_15738);
nor U17065 (N_17065,N_14132,N_14679);
xor U17066 (N_17066,N_14203,N_14464);
nand U17067 (N_17067,N_14649,N_14788);
nand U17068 (N_17068,N_12620,N_13961);
nor U17069 (N_17069,N_15583,N_15267);
nand U17070 (N_17070,N_12791,N_14719);
and U17071 (N_17071,N_15693,N_12691);
nand U17072 (N_17072,N_15367,N_13443);
nand U17073 (N_17073,N_14545,N_13106);
nor U17074 (N_17074,N_15568,N_15974);
nor U17075 (N_17075,N_14706,N_15148);
nor U17076 (N_17076,N_12636,N_13145);
nor U17077 (N_17077,N_14515,N_14583);
nor U17078 (N_17078,N_14792,N_14678);
xnor U17079 (N_17079,N_14379,N_15105);
xnor U17080 (N_17080,N_14338,N_15630);
nand U17081 (N_17081,N_14922,N_13893);
and U17082 (N_17082,N_12956,N_15429);
nand U17083 (N_17083,N_13123,N_15381);
or U17084 (N_17084,N_15451,N_13212);
or U17085 (N_17085,N_13532,N_15612);
xnor U17086 (N_17086,N_12410,N_14170);
and U17087 (N_17087,N_14752,N_14303);
xnor U17088 (N_17088,N_15665,N_12175);
and U17089 (N_17089,N_13211,N_12916);
or U17090 (N_17090,N_15510,N_15191);
or U17091 (N_17091,N_12011,N_15358);
or U17092 (N_17092,N_13665,N_12324);
and U17093 (N_17093,N_13332,N_13651);
or U17094 (N_17094,N_15284,N_14270);
and U17095 (N_17095,N_12722,N_13210);
and U17096 (N_17096,N_14811,N_12461);
nor U17097 (N_17097,N_15445,N_15007);
nand U17098 (N_17098,N_13463,N_15981);
nor U17099 (N_17099,N_13284,N_12455);
or U17100 (N_17100,N_14448,N_13683);
xor U17101 (N_17101,N_14331,N_14251);
and U17102 (N_17102,N_12031,N_14999);
nand U17103 (N_17103,N_12928,N_14601);
or U17104 (N_17104,N_15290,N_15002);
or U17105 (N_17105,N_13455,N_13242);
and U17106 (N_17106,N_14573,N_12168);
and U17107 (N_17107,N_15444,N_14336);
or U17108 (N_17108,N_13407,N_12639);
nor U17109 (N_17109,N_14149,N_12092);
or U17110 (N_17110,N_12403,N_12693);
or U17111 (N_17111,N_15661,N_12044);
or U17112 (N_17112,N_14327,N_15923);
nor U17113 (N_17113,N_15321,N_12733);
nand U17114 (N_17114,N_13310,N_13005);
or U17115 (N_17115,N_13682,N_12392);
xor U17116 (N_17116,N_13957,N_13977);
nor U17117 (N_17117,N_14399,N_12234);
nand U17118 (N_17118,N_12913,N_15086);
xor U17119 (N_17119,N_15791,N_13301);
nor U17120 (N_17120,N_13075,N_13689);
nor U17121 (N_17121,N_14909,N_14960);
or U17122 (N_17122,N_13949,N_13282);
and U17123 (N_17123,N_13274,N_12135);
nand U17124 (N_17124,N_13091,N_15463);
and U17125 (N_17125,N_12699,N_13674);
or U17126 (N_17126,N_13722,N_12120);
and U17127 (N_17127,N_13789,N_14413);
and U17128 (N_17128,N_15022,N_14749);
and U17129 (N_17129,N_14364,N_13698);
and U17130 (N_17130,N_15070,N_14188);
nor U17131 (N_17131,N_12144,N_12034);
nand U17132 (N_17132,N_13353,N_15250);
and U17133 (N_17133,N_12547,N_14479);
or U17134 (N_17134,N_12643,N_12320);
and U17135 (N_17135,N_14722,N_12285);
nor U17136 (N_17136,N_14709,N_15794);
and U17137 (N_17137,N_15498,N_14901);
nand U17138 (N_17138,N_12473,N_14007);
and U17139 (N_17139,N_12802,N_13842);
or U17140 (N_17140,N_15113,N_12829);
nor U17141 (N_17141,N_14332,N_12753);
or U17142 (N_17142,N_12681,N_15908);
or U17143 (N_17143,N_15131,N_15479);
or U17144 (N_17144,N_14456,N_12263);
xnor U17145 (N_17145,N_13505,N_14628);
nand U17146 (N_17146,N_14012,N_12060);
or U17147 (N_17147,N_13043,N_12808);
nor U17148 (N_17148,N_12918,N_12155);
nand U17149 (N_17149,N_13118,N_15604);
xor U17150 (N_17150,N_13596,N_12781);
nand U17151 (N_17151,N_15779,N_12071);
xnor U17152 (N_17152,N_15729,N_14221);
nand U17153 (N_17153,N_12450,N_14685);
nand U17154 (N_17154,N_15634,N_15028);
and U17155 (N_17155,N_14661,N_14380);
or U17156 (N_17156,N_12440,N_14298);
or U17157 (N_17157,N_15487,N_13053);
and U17158 (N_17158,N_13002,N_13580);
nor U17159 (N_17159,N_12391,N_13191);
nor U17160 (N_17160,N_15225,N_12790);
or U17161 (N_17161,N_15709,N_15061);
nor U17162 (N_17162,N_14403,N_12622);
nand U17163 (N_17163,N_15668,N_15855);
and U17164 (N_17164,N_12357,N_13036);
nor U17165 (N_17165,N_13196,N_15393);
nand U17166 (N_17166,N_13239,N_15726);
nand U17167 (N_17167,N_12674,N_12065);
nor U17168 (N_17168,N_14585,N_12545);
and U17169 (N_17169,N_13773,N_12887);
xnor U17170 (N_17170,N_12309,N_12201);
and U17171 (N_17171,N_14765,N_14416);
and U17172 (N_17172,N_13174,N_12694);
nor U17173 (N_17173,N_13126,N_13503);
and U17174 (N_17174,N_15359,N_13317);
nor U17175 (N_17175,N_15035,N_12713);
xnor U17176 (N_17176,N_12614,N_12240);
nor U17177 (N_17177,N_15409,N_14022);
xor U17178 (N_17178,N_15983,N_12590);
nand U17179 (N_17179,N_12891,N_14647);
or U17180 (N_17180,N_13729,N_14600);
and U17181 (N_17181,N_14252,N_12290);
nand U17182 (N_17182,N_13127,N_13164);
and U17183 (N_17183,N_12948,N_12147);
or U17184 (N_17184,N_15245,N_15607);
nand U17185 (N_17185,N_13690,N_15609);
or U17186 (N_17186,N_12605,N_13087);
and U17187 (N_17187,N_13823,N_13411);
or U17188 (N_17188,N_15877,N_14410);
nor U17189 (N_17189,N_12465,N_15677);
or U17190 (N_17190,N_12654,N_14116);
or U17191 (N_17191,N_14141,N_15702);
and U17192 (N_17192,N_12850,N_13799);
and U17193 (N_17193,N_14228,N_12692);
and U17194 (N_17194,N_14928,N_13388);
nor U17195 (N_17195,N_15220,N_15420);
nand U17196 (N_17196,N_13007,N_15730);
and U17197 (N_17197,N_14256,N_14735);
xnor U17198 (N_17198,N_14185,N_12656);
and U17199 (N_17199,N_12773,N_14757);
and U17200 (N_17200,N_14113,N_15089);
xor U17201 (N_17201,N_13010,N_13224);
and U17202 (N_17202,N_15364,N_12961);
nand U17203 (N_17203,N_14428,N_12908);
or U17204 (N_17204,N_12179,N_12382);
nand U17205 (N_17205,N_13536,N_12236);
xor U17206 (N_17206,N_13820,N_15530);
or U17207 (N_17207,N_15850,N_14575);
or U17208 (N_17208,N_15039,N_12516);
nor U17209 (N_17209,N_14781,N_12789);
nor U17210 (N_17210,N_12532,N_14264);
and U17211 (N_17211,N_15457,N_12349);
or U17212 (N_17212,N_14925,N_13412);
or U17213 (N_17213,N_14447,N_12376);
and U17214 (N_17214,N_15480,N_13339);
nand U17215 (N_17215,N_12103,N_14400);
and U17216 (N_17216,N_14814,N_13398);
or U17217 (N_17217,N_12182,N_14091);
and U17218 (N_17218,N_13984,N_12466);
or U17219 (N_17219,N_12649,N_14910);
or U17220 (N_17220,N_13771,N_14092);
nor U17221 (N_17221,N_14691,N_13078);
and U17222 (N_17222,N_12360,N_12985);
nand U17223 (N_17223,N_12379,N_13428);
nand U17224 (N_17224,N_15224,N_14572);
or U17225 (N_17225,N_12635,N_15383);
and U17226 (N_17226,N_13435,N_13028);
or U17227 (N_17227,N_13954,N_13124);
nor U17228 (N_17228,N_15363,N_12045);
nor U17229 (N_17229,N_14714,N_12083);
or U17230 (N_17230,N_12797,N_12061);
xor U17231 (N_17231,N_14328,N_12364);
and U17232 (N_17232,N_15357,N_13693);
and U17233 (N_17233,N_15805,N_14676);
nor U17234 (N_17234,N_13351,N_12452);
xor U17235 (N_17235,N_15109,N_12404);
xnor U17236 (N_17236,N_13530,N_14032);
and U17237 (N_17237,N_13287,N_12208);
or U17238 (N_17238,N_12427,N_13684);
xor U17239 (N_17239,N_13882,N_13190);
and U17240 (N_17240,N_13294,N_12128);
or U17241 (N_17241,N_12941,N_14044);
nor U17242 (N_17242,N_14912,N_12920);
or U17243 (N_17243,N_13531,N_13066);
nand U17244 (N_17244,N_15973,N_14466);
or U17245 (N_17245,N_13278,N_15000);
or U17246 (N_17246,N_14855,N_14897);
xnor U17247 (N_17247,N_13811,N_12063);
nor U17248 (N_17248,N_13068,N_14183);
xor U17249 (N_17249,N_12353,N_12124);
and U17250 (N_17250,N_13998,N_15622);
nor U17251 (N_17251,N_14293,N_14965);
and U17252 (N_17252,N_13055,N_12546);
or U17253 (N_17253,N_12953,N_13422);
nand U17254 (N_17254,N_13728,N_12978);
nor U17255 (N_17255,N_15854,N_14591);
nor U17256 (N_17256,N_14677,N_14969);
xnor U17257 (N_17257,N_13345,N_15878);
and U17258 (N_17258,N_15403,N_15906);
xor U17259 (N_17259,N_15256,N_15704);
nor U17260 (N_17260,N_12460,N_15201);
nand U17261 (N_17261,N_13234,N_15696);
nand U17262 (N_17262,N_15189,N_12411);
and U17263 (N_17263,N_15410,N_15488);
or U17264 (N_17264,N_14059,N_14085);
or U17265 (N_17265,N_14442,N_15977);
or U17266 (N_17266,N_13090,N_15950);
nor U17267 (N_17267,N_13956,N_13025);
and U17268 (N_17268,N_14263,N_15553);
and U17269 (N_17269,N_12301,N_15786);
nand U17270 (N_17270,N_13538,N_14702);
xor U17271 (N_17271,N_12021,N_12890);
nor U17272 (N_17272,N_15052,N_15901);
and U17273 (N_17273,N_12389,N_14602);
nor U17274 (N_17274,N_14592,N_14711);
nor U17275 (N_17275,N_14440,N_15920);
nor U17276 (N_17276,N_14232,N_13629);
or U17277 (N_17277,N_13941,N_15706);
nand U17278 (N_17278,N_14337,N_12053);
or U17279 (N_17279,N_15315,N_12755);
or U17280 (N_17280,N_12519,N_14791);
or U17281 (N_17281,N_12265,N_15178);
and U17282 (N_17282,N_15548,N_14986);
nand U17283 (N_17283,N_15439,N_15100);
xnor U17284 (N_17284,N_13676,N_14506);
xnor U17285 (N_17285,N_15538,N_15448);
and U17286 (N_17286,N_15169,N_14837);
or U17287 (N_17287,N_13898,N_15184);
nand U17288 (N_17288,N_12210,N_15916);
and U17289 (N_17289,N_14956,N_15699);
or U17290 (N_17290,N_12329,N_15336);
and U17291 (N_17291,N_15162,N_15963);
and U17292 (N_17292,N_12318,N_14483);
xnor U17293 (N_17293,N_15063,N_15266);
xnor U17294 (N_17294,N_13080,N_14775);
and U17295 (N_17295,N_12729,N_13132);
nand U17296 (N_17296,N_14812,N_14768);
xor U17297 (N_17297,N_15897,N_13964);
nand U17298 (N_17298,N_12055,N_14118);
nor U17299 (N_17299,N_13466,N_15951);
or U17300 (N_17300,N_12740,N_14878);
xor U17301 (N_17301,N_15379,N_13133);
or U17302 (N_17302,N_14810,N_13746);
nor U17303 (N_17303,N_15394,N_14392);
or U17304 (N_17304,N_14200,N_12754);
nor U17305 (N_17305,N_15813,N_13650);
nand U17306 (N_17306,N_13767,N_14849);
nor U17307 (N_17307,N_13427,N_15972);
nor U17308 (N_17308,N_13843,N_15533);
xor U17309 (N_17309,N_15646,N_15731);
or U17310 (N_17310,N_15173,N_15091);
nand U17311 (N_17311,N_14124,N_13705);
nand U17312 (N_17312,N_15703,N_15928);
or U17313 (N_17313,N_12919,N_15205);
nor U17314 (N_17314,N_13141,N_13297);
and U17315 (N_17315,N_14819,N_14390);
or U17316 (N_17316,N_12006,N_13926);
nand U17317 (N_17317,N_12721,N_15521);
and U17318 (N_17318,N_13470,N_13019);
nand U17319 (N_17319,N_12738,N_13815);
xnor U17320 (N_17320,N_13222,N_13319);
and U17321 (N_17321,N_15590,N_13067);
nor U17322 (N_17322,N_13606,N_14566);
nor U17323 (N_17323,N_12623,N_13404);
or U17324 (N_17324,N_12059,N_13352);
nor U17325 (N_17325,N_12010,N_12935);
nor U17326 (N_17326,N_14843,N_13671);
nand U17327 (N_17327,N_14282,N_13782);
and U17328 (N_17328,N_12475,N_15104);
xor U17329 (N_17329,N_14842,N_12187);
nand U17330 (N_17330,N_15289,N_13130);
or U17331 (N_17331,N_13973,N_12459);
or U17332 (N_17332,N_14921,N_12728);
nor U17333 (N_17333,N_12211,N_12277);
nor U17334 (N_17334,N_13801,N_12009);
nor U17335 (N_17335,N_14541,N_12296);
xor U17336 (N_17336,N_14433,N_14178);
and U17337 (N_17337,N_13863,N_12834);
or U17338 (N_17338,N_14640,N_15239);
and U17339 (N_17339,N_13335,N_14196);
nand U17340 (N_17340,N_13046,N_14984);
or U17341 (N_17341,N_14384,N_14068);
nand U17342 (N_17342,N_13680,N_13442);
nor U17343 (N_17343,N_13640,N_14224);
xnor U17344 (N_17344,N_15333,N_12517);
or U17345 (N_17345,N_13188,N_15686);
nand U17346 (N_17346,N_13756,N_15396);
and U17347 (N_17347,N_14412,N_13264);
and U17348 (N_17348,N_13904,N_12736);
nand U17349 (N_17349,N_15270,N_13774);
nor U17350 (N_17350,N_15971,N_15330);
or U17351 (N_17351,N_15397,N_13410);
nand U17352 (N_17352,N_15254,N_13392);
nand U17353 (N_17353,N_13439,N_12746);
nor U17354 (N_17354,N_13809,N_14650);
nand U17355 (N_17355,N_12876,N_12923);
or U17356 (N_17356,N_14370,N_12513);
or U17357 (N_17357,N_14536,N_13476);
or U17358 (N_17358,N_13496,N_13945);
or U17359 (N_17359,N_13265,N_14052);
nand U17360 (N_17360,N_13739,N_12474);
xor U17361 (N_17361,N_13120,N_13924);
or U17362 (N_17362,N_14254,N_15841);
and U17363 (N_17363,N_12227,N_13585);
xnor U17364 (N_17364,N_12146,N_15541);
xnor U17365 (N_17365,N_13303,N_14266);
nand U17366 (N_17366,N_15753,N_15467);
xnor U17367 (N_17367,N_13146,N_13170);
or U17368 (N_17368,N_12313,N_14799);
or U17369 (N_17369,N_15356,N_13577);
nand U17370 (N_17370,N_12117,N_12842);
and U17371 (N_17371,N_13913,N_14385);
and U17372 (N_17372,N_13291,N_13802);
or U17373 (N_17373,N_14608,N_13938);
nand U17374 (N_17374,N_14248,N_15120);
or U17375 (N_17375,N_13872,N_15785);
nand U17376 (N_17376,N_13638,N_14341);
or U17377 (N_17377,N_13590,N_14605);
and U17378 (N_17378,N_12091,N_14418);
nor U17379 (N_17379,N_15830,N_15215);
nand U17380 (N_17380,N_12186,N_13415);
and U17381 (N_17381,N_12529,N_15818);
or U17382 (N_17382,N_12795,N_14356);
nand U17383 (N_17383,N_14104,N_14918);
and U17384 (N_17384,N_15370,N_14180);
or U17385 (N_17385,N_13233,N_12819);
nand U17386 (N_17386,N_15295,N_13578);
or U17387 (N_17387,N_13348,N_15758);
or U17388 (N_17388,N_13686,N_13409);
nand U17389 (N_17389,N_12344,N_14437);
nor U17390 (N_17390,N_12462,N_14774);
xor U17391 (N_17391,N_14847,N_15656);
or U17392 (N_17392,N_15980,N_15351);
nor U17393 (N_17393,N_14908,N_13714);
or U17394 (N_17394,N_15712,N_13533);
nand U17395 (N_17395,N_14581,N_13227);
nand U17396 (N_17396,N_12258,N_13281);
nor U17397 (N_17397,N_13626,N_15552);
nand U17398 (N_17398,N_13359,N_14852);
and U17399 (N_17399,N_15936,N_14665);
or U17400 (N_17400,N_12984,N_15271);
xor U17401 (N_17401,N_12929,N_12488);
or U17402 (N_17402,N_13839,N_13402);
nand U17403 (N_17403,N_15096,N_15069);
nand U17404 (N_17404,N_12784,N_13361);
nor U17405 (N_17405,N_15982,N_12747);
or U17406 (N_17406,N_14569,N_14728);
or U17407 (N_17407,N_14304,N_14604);
nor U17408 (N_17408,N_13200,N_12073);
nor U17409 (N_17409,N_14407,N_13994);
nor U17410 (N_17410,N_12413,N_12895);
or U17411 (N_17411,N_12431,N_13201);
and U17412 (N_17412,N_12255,N_13541);
nor U17413 (N_17413,N_14477,N_14216);
nand U17414 (N_17414,N_14579,N_14329);
nand U17415 (N_17415,N_15041,N_12116);
and U17416 (N_17416,N_13672,N_15559);
xor U17417 (N_17417,N_12385,N_12843);
or U17418 (N_17418,N_13840,N_15637);
nand U17419 (N_17419,N_12665,N_13892);
and U17420 (N_17420,N_14846,N_13742);
nand U17421 (N_17421,N_13569,N_15986);
and U17422 (N_17422,N_15075,N_15141);
nor U17423 (N_17423,N_13664,N_15653);
nor U17424 (N_17424,N_13047,N_13331);
nand U17425 (N_17425,N_14041,N_13932);
or U17426 (N_17426,N_14551,N_15742);
nand U17427 (N_17427,N_14358,N_15283);
and U17428 (N_17428,N_14353,N_12390);
nor U17429 (N_17429,N_12104,N_12991);
nand U17430 (N_17430,N_14502,N_15434);
nand U17431 (N_17431,N_13544,N_12811);
nor U17432 (N_17432,N_13171,N_15628);
or U17433 (N_17433,N_12214,N_13960);
and U17434 (N_17434,N_15968,N_15422);
and U17435 (N_17435,N_14713,N_12237);
and U17436 (N_17436,N_12703,N_14409);
nand U17437 (N_17437,N_13464,N_15018);
nor U17438 (N_17438,N_14243,N_12900);
nand U17439 (N_17439,N_14675,N_13602);
xor U17440 (N_17440,N_15581,N_14557);
nor U17441 (N_17441,N_15056,N_14097);
nor U17442 (N_17442,N_12084,N_15965);
nor U17443 (N_17443,N_12962,N_14599);
or U17444 (N_17444,N_13850,N_13017);
xnor U17445 (N_17445,N_14933,N_15098);
nor U17446 (N_17446,N_14742,N_15365);
nor U17447 (N_17447,N_15192,N_12399);
nand U17448 (N_17448,N_15437,N_15219);
nand U17449 (N_17449,N_13837,N_15154);
or U17450 (N_17450,N_12454,N_15773);
xnor U17451 (N_17451,N_15419,N_12523);
and U17452 (N_17452,N_14565,N_14698);
and U17453 (N_17453,N_13277,N_14027);
or U17454 (N_17454,N_14831,N_14932);
nand U17455 (N_17455,N_13290,N_15871);
or U17456 (N_17456,N_15171,N_12631);
or U17457 (N_17457,N_12629,N_12606);
nor U17458 (N_17458,N_15766,N_12274);
xnor U17459 (N_17459,N_12673,N_15226);
nor U17460 (N_17460,N_13962,N_12192);
and U17461 (N_17461,N_15492,N_15081);
nor U17462 (N_17462,N_12127,N_13076);
nor U17463 (N_17463,N_12500,N_14700);
nand U17464 (N_17464,N_12425,N_12342);
and U17465 (N_17465,N_15695,N_15775);
or U17466 (N_17466,N_15542,N_14803);
or U17467 (N_17467,N_12870,N_13381);
and U17468 (N_17468,N_12048,N_14374);
and U17469 (N_17469,N_15836,N_13226);
nand U17470 (N_17470,N_14556,N_12446);
or U17471 (N_17471,N_13216,N_12185);
xnor U17472 (N_17472,N_14383,N_12041);
and U17473 (N_17473,N_14725,N_15242);
nand U17474 (N_17474,N_15469,N_15969);
or U17475 (N_17475,N_13581,N_14305);
nand U17476 (N_17476,N_14945,N_12677);
or U17477 (N_17477,N_14667,N_13867);
and U17478 (N_17478,N_12739,N_12660);
nand U17479 (N_17479,N_13192,N_14963);
xnor U17480 (N_17480,N_15857,N_12845);
and U17481 (N_17481,N_15449,N_12951);
or U17482 (N_17482,N_12974,N_14175);
nand U17483 (N_17483,N_14511,N_15851);
or U17484 (N_17484,N_13082,N_13687);
or U17485 (N_17485,N_13268,N_15797);
xnor U17486 (N_17486,N_14876,N_14785);
nand U17487 (N_17487,N_12123,N_13833);
and U17488 (N_17488,N_15700,N_12875);
nor U17489 (N_17489,N_14884,N_15343);
or U17490 (N_17490,N_14074,N_13434);
nand U17491 (N_17491,N_13378,N_14603);
or U17492 (N_17492,N_15344,N_12633);
nor U17493 (N_17493,N_12172,N_13511);
and U17494 (N_17494,N_12963,N_12638);
and U17495 (N_17495,N_15114,N_15780);
or U17496 (N_17496,N_14072,N_13663);
nor U17497 (N_17497,N_13110,N_14936);
and U17498 (N_17498,N_13058,N_12583);
xor U17499 (N_17499,N_12830,N_13783);
nand U17500 (N_17500,N_15565,N_12430);
and U17501 (N_17501,N_13060,N_14137);
nor U17502 (N_17502,N_15431,N_12936);
nand U17503 (N_17503,N_15464,N_12062);
and U17504 (N_17504,N_15455,N_13937);
and U17505 (N_17505,N_15294,N_14952);
nand U17506 (N_17506,N_14096,N_13488);
nor U17507 (N_17507,N_14274,N_15217);
nor U17508 (N_17508,N_15037,N_12835);
and U17509 (N_17509,N_15179,N_12993);
nand U17510 (N_17510,N_12541,N_12761);
and U17511 (N_17511,N_15038,N_12602);
nand U17512 (N_17512,N_12731,N_14795);
or U17513 (N_17513,N_12610,N_13715);
nor U17514 (N_17514,N_14888,N_15048);
xor U17515 (N_17515,N_12796,N_13038);
or U17516 (N_17516,N_15415,N_15160);
nand U17517 (N_17517,N_13632,N_13423);
or U17518 (N_17518,N_13906,N_12332);
and U17519 (N_17519,N_15156,N_14753);
nand U17520 (N_17520,N_15032,N_14233);
nand U17521 (N_17521,N_15734,N_13631);
nor U17522 (N_17522,N_12497,N_12444);
xor U17523 (N_17523,N_14361,N_13993);
and U17524 (N_17524,N_14817,N_13744);
or U17525 (N_17525,N_12191,N_14694);
and U17526 (N_17526,N_15517,N_12858);
nor U17527 (N_17527,N_14954,N_15476);
nor U17528 (N_17528,N_15593,N_13246);
xnor U17529 (N_17529,N_12996,N_14697);
and U17530 (N_17530,N_14828,N_13107);
nand U17531 (N_17531,N_13621,N_15475);
and U17532 (N_17532,N_15312,N_13848);
and U17533 (N_17533,N_15944,N_15883);
or U17534 (N_17534,N_12849,N_15115);
nand U17535 (N_17535,N_12550,N_14033);
and U17536 (N_17536,N_12421,N_13289);
nand U17537 (N_17537,N_13725,N_12004);
nand U17538 (N_17538,N_14997,N_14177);
or U17539 (N_17539,N_12158,N_12177);
xor U17540 (N_17540,N_13936,N_15625);
and U17541 (N_17541,N_14570,N_14968);
and U17542 (N_17542,N_13630,N_13461);
nand U17543 (N_17543,N_12369,N_15890);
or U17544 (N_17544,N_14931,N_13045);
nor U17545 (N_17545,N_14574,N_15200);
nand U17546 (N_17546,N_15991,N_12684);
or U17547 (N_17547,N_14192,N_13269);
nand U17548 (N_17548,N_15124,N_12067);
nor U17549 (N_17549,N_12565,N_14505);
nor U17550 (N_17550,N_13805,N_15662);
nor U17551 (N_17551,N_12898,N_15005);
nand U17552 (N_17552,N_12804,N_13880);
xor U17553 (N_17553,N_14879,N_15411);
and U17554 (N_17554,N_15407,N_15616);
or U17555 (N_17555,N_12946,N_13794);
and U17556 (N_17556,N_12701,N_14595);
nor U17557 (N_17557,N_13350,N_13772);
or U17558 (N_17558,N_15257,N_14955);
nor U17559 (N_17559,N_12507,N_14531);
or U17560 (N_17560,N_12938,N_14543);
nor U17561 (N_17561,N_14992,N_13252);
or U17562 (N_17562,N_15090,N_15485);
nand U17563 (N_17563,N_14114,N_12282);
nand U17564 (N_17564,N_14732,N_14745);
nand U17565 (N_17565,N_12161,N_13438);
or U17566 (N_17566,N_13607,N_14911);
and U17567 (N_17567,N_12607,N_13347);
and U17568 (N_17568,N_14064,N_15964);
or U17569 (N_17569,N_15834,N_14723);
xor U17570 (N_17570,N_12070,N_13425);
or U17571 (N_17571,N_14315,N_14902);
xnor U17572 (N_17572,N_15674,N_15152);
or U17573 (N_17573,N_14394,N_12591);
nand U17574 (N_17574,N_15884,N_12765);
and U17575 (N_17575,N_12096,N_13942);
and U17576 (N_17576,N_12866,N_13256);
or U17577 (N_17577,N_15627,N_14853);
and U17578 (N_17578,N_12449,N_15867);
nor U17579 (N_17579,N_13588,N_15466);
xnor U17580 (N_17580,N_15563,N_12528);
and U17581 (N_17581,N_12877,N_14133);
nand U17582 (N_17582,N_12823,N_15408);
or U17583 (N_17583,N_12760,N_13016);
nand U17584 (N_17584,N_12345,N_15478);
or U17585 (N_17585,N_15214,N_15520);
and U17586 (N_17586,N_13869,N_12960);
or U17587 (N_17587,N_14562,N_14423);
nor U17588 (N_17588,N_12224,N_15021);
nand U17589 (N_17589,N_12312,N_12242);
nand U17590 (N_17590,N_12220,N_15325);
nand U17591 (N_17591,N_12906,N_13545);
nand U17592 (N_17592,N_12570,N_14261);
xor U17593 (N_17593,N_14726,N_15302);
or U17594 (N_17594,N_15608,N_12362);
nor U17595 (N_17595,N_14366,N_15017);
nor U17596 (N_17596,N_14627,N_15277);
and U17597 (N_17597,N_13825,N_13024);
nand U17598 (N_17598,N_14844,N_12815);
nand U17599 (N_17599,N_13713,N_13717);
or U17600 (N_17600,N_15259,N_12496);
nand U17601 (N_17601,N_13169,N_15029);
nor U17602 (N_17602,N_12743,N_13912);
nor U17603 (N_17603,N_12612,N_14271);
nand U17604 (N_17604,N_14840,N_13915);
nand U17605 (N_17605,N_14821,N_12903);
nand U17606 (N_17606,N_15966,N_14729);
nand U17607 (N_17607,N_15869,N_15611);
and U17608 (N_17608,N_12480,N_15998);
and U17609 (N_17609,N_12944,N_12652);
nand U17610 (N_17610,N_12442,N_14760);
nand U17611 (N_17611,N_13634,N_13102);
or U17612 (N_17612,N_12844,N_15929);
nand U17613 (N_17613,N_13440,N_12054);
or U17614 (N_17614,N_14873,N_15051);
nand U17615 (N_17615,N_15023,N_12992);
or U17616 (N_17616,N_14110,N_13383);
xnor U17617 (N_17617,N_13557,N_14883);
and U17618 (N_17618,N_12750,N_14365);
and U17619 (N_17619,N_13454,N_14633);
nor U17620 (N_17620,N_14340,N_14862);
and U17621 (N_17621,N_12365,N_14422);
or U17622 (N_17622,N_14689,N_14619);
or U17623 (N_17623,N_13109,N_14587);
xor U17624 (N_17624,N_14481,N_13858);
or U17625 (N_17625,N_15764,N_15509);
nor U17626 (N_17626,N_12959,N_12445);
nor U17627 (N_17627,N_14771,N_14173);
xor U17628 (N_17628,N_14036,N_13449);
or U17629 (N_17629,N_12617,N_14334);
or U17630 (N_17630,N_13135,N_13136);
or U17631 (N_17631,N_14737,N_14193);
and U17632 (N_17632,N_15988,N_13198);
nor U17633 (N_17633,N_13512,N_15814);
and U17634 (N_17634,N_15578,N_14653);
nand U17635 (N_17635,N_13899,N_15027);
and U17636 (N_17636,N_12154,N_15588);
nor U17637 (N_17637,N_12451,N_14230);
nand U17638 (N_17638,N_12149,N_13329);
or U17639 (N_17639,N_14967,N_13909);
nand U17640 (N_17640,N_13254,N_15839);
nand U17641 (N_17641,N_14325,N_13661);
xnor U17642 (N_17642,N_12408,N_12579);
nor U17643 (N_17643,N_14432,N_14731);
nor U17644 (N_17644,N_13336,N_14993);
nand U17645 (N_17645,N_15927,N_13462);
nor U17646 (N_17646,N_12556,N_12878);
or U17647 (N_17647,N_14739,N_12573);
xnor U17648 (N_17648,N_13215,N_13079);
and U17649 (N_17649,N_12139,N_15885);
nor U17650 (N_17650,N_13905,N_12132);
nand U17651 (N_17651,N_14278,N_15913);
nor U17652 (N_17652,N_15528,N_13509);
nand U17653 (N_17653,N_14195,N_15229);
nor U17654 (N_17654,N_13546,N_14454);
xor U17655 (N_17655,N_13516,N_13727);
xor U17656 (N_17656,N_12026,N_15421);
nand U17657 (N_17657,N_14636,N_15077);
and U17658 (N_17658,N_15518,N_13063);
and U17659 (N_17659,N_15632,N_14267);
nand U17660 (N_17660,N_14544,N_12549);
or U17661 (N_17661,N_13059,N_13865);
or U17662 (N_17662,N_14836,N_12331);
or U17663 (N_17663,N_12712,N_14159);
or U17664 (N_17664,N_14474,N_13859);
nand U17665 (N_17665,N_14874,N_14896);
nor U17666 (N_17666,N_15194,N_14829);
nand U17667 (N_17667,N_15960,N_15735);
or U17668 (N_17668,N_14276,N_13483);
nor U17669 (N_17669,N_14550,N_13515);
or U17670 (N_17670,N_15040,N_12741);
nor U17671 (N_17671,N_14108,N_12727);
nor U17672 (N_17672,N_15491,N_15522);
and U17673 (N_17673,N_12040,N_13769);
or U17674 (N_17674,N_14508,N_13619);
and U17675 (N_17675,N_12702,N_12770);
nor U17676 (N_17676,N_14490,N_13612);
and U17677 (N_17677,N_14081,N_12535);
nor U17678 (N_17678,N_13890,N_15995);
nand U17679 (N_17679,N_14103,N_15195);
nor U17680 (N_17680,N_13139,N_12596);
xor U17681 (N_17681,N_15808,N_15398);
xnor U17682 (N_17682,N_15663,N_13413);
nor U17683 (N_17683,N_12295,N_15782);
nand U17684 (N_17684,N_13179,N_12563);
and U17685 (N_17685,N_14669,N_14135);
or U17686 (N_17686,N_14421,N_12767);
or U17687 (N_17687,N_14308,N_14643);
and U17688 (N_17688,N_15591,N_15907);
nand U17689 (N_17689,N_15529,N_12122);
nor U17690 (N_17690,N_13726,N_13653);
nand U17691 (N_17691,N_15796,N_12476);
nand U17692 (N_17692,N_12222,N_12954);
and U17693 (N_17693,N_14715,N_14368);
or U17694 (N_17694,N_13021,N_14452);
or U17695 (N_17695,N_15902,N_13593);
xnor U17696 (N_17696,N_14273,N_14145);
or U17697 (N_17697,N_15999,N_13478);
nand U17698 (N_17698,N_12407,N_12577);
and U17699 (N_17699,N_13875,N_15282);
nand U17700 (N_17700,N_14624,N_12085);
nor U17701 (N_17701,N_14171,N_12828);
or U17702 (N_17702,N_14058,N_12412);
or U17703 (N_17703,N_15800,N_13526);
or U17704 (N_17704,N_14913,N_12732);
and U17705 (N_17705,N_14754,N_15954);
or U17706 (N_17706,N_15176,N_15082);
or U17707 (N_17707,N_13168,N_13618);
or U17708 (N_17708,N_15868,N_14629);
nand U17709 (N_17709,N_14244,N_13587);
nor U17710 (N_17710,N_13948,N_15945);
xnor U17711 (N_17711,N_15117,N_13279);
or U17712 (N_17712,N_12718,N_15080);
nand U17713 (N_17713,N_15997,N_14077);
and U17714 (N_17714,N_15594,N_12667);
nand U17715 (N_17715,N_12032,N_15352);
nor U17716 (N_17716,N_12933,N_12303);
nand U17717 (N_17717,N_15130,N_15793);
nand U17718 (N_17718,N_14283,N_12109);
and U17719 (N_17719,N_15624,N_14449);
or U17720 (N_17720,N_13886,N_12557);
and U17721 (N_17721,N_15442,N_15784);
or U17722 (N_17722,N_14571,N_12491);
and U17723 (N_17723,N_12157,N_12378);
nand U17724 (N_17724,N_12863,N_13598);
or U17725 (N_17725,N_12597,N_14748);
or U17726 (N_17726,N_14128,N_14062);
nand U17727 (N_17727,N_15783,N_15097);
and U17728 (N_17728,N_14982,N_14900);
nand U17729 (N_17729,N_14281,N_15142);
xor U17730 (N_17730,N_13175,N_15717);
and U17731 (N_17731,N_12889,N_14319);
nor U17732 (N_17732,N_15443,N_15112);
and U17733 (N_17733,N_14459,N_13710);
nand U17734 (N_17734,N_12989,N_12424);
and U17735 (N_17735,N_14023,N_13293);
and U17736 (N_17736,N_14826,N_13026);
and U17737 (N_17737,N_12634,N_12982);
nor U17738 (N_17738,N_15303,N_13836);
or U17739 (N_17739,N_12160,N_15918);
nand U17740 (N_17740,N_12463,N_14371);
and U17741 (N_17741,N_14503,N_15640);
nor U17742 (N_17742,N_12368,N_15790);
or U17743 (N_17743,N_12637,N_14850);
or U17744 (N_17744,N_14420,N_15285);
or U17745 (N_17745,N_13420,N_12786);
and U17746 (N_17746,N_15133,N_13760);
and U17747 (N_17747,N_12885,N_14335);
nor U17748 (N_17748,N_12751,N_13897);
and U17749 (N_17749,N_12354,N_15145);
nor U17750 (N_17750,N_14870,N_13980);
nand U17751 (N_17751,N_15143,N_12489);
nand U17752 (N_17752,N_12976,N_15150);
nand U17753 (N_17753,N_14427,N_13636);
or U17754 (N_17754,N_14598,N_13202);
nand U17755 (N_17755,N_13377,N_12554);
or U17756 (N_17756,N_12156,N_15318);
nor U17757 (N_17757,N_12016,N_15264);
or U17758 (N_17758,N_14485,N_12666);
or U17759 (N_17759,N_15360,N_13357);
or U17760 (N_17760,N_12901,N_12358);
and U17761 (N_17761,N_15401,N_13616);
nor U17762 (N_17762,N_14069,N_12115);
xnor U17763 (N_17763,N_13094,N_12162);
nand U17764 (N_17764,N_12952,N_12800);
nand U17765 (N_17765,N_13534,N_14002);
and U17766 (N_17766,N_14312,N_15019);
nand U17767 (N_17767,N_12776,N_15691);
and U17768 (N_17768,N_14136,N_14818);
nor U17769 (N_17769,N_12226,N_12205);
and U17770 (N_17770,N_14473,N_13144);
and U17771 (N_17771,N_15043,N_12641);
xor U17772 (N_17772,N_12218,N_15962);
and U17773 (N_17773,N_15598,N_15870);
nor U17774 (N_17774,N_14029,N_15597);
or U17775 (N_17775,N_14899,N_13617);
or U17776 (N_17776,N_13911,N_12524);
nor U17777 (N_17777,N_14530,N_13373);
nand U17778 (N_17778,N_12697,N_15064);
nand U17779 (N_17779,N_14396,N_15430);
xor U17780 (N_17780,N_13489,N_14959);
and U17781 (N_17781,N_14724,N_13249);
and U17782 (N_17782,N_12381,N_12097);
nor U17783 (N_17783,N_14898,N_13594);
xor U17784 (N_17784,N_14796,N_15570);
nand U17785 (N_17785,N_12188,N_12757);
xor U17786 (N_17786,N_12183,N_12526);
nor U17787 (N_17787,N_13981,N_14696);
nor U17788 (N_17788,N_14851,N_12088);
or U17789 (N_17789,N_12779,N_15667);
or U17790 (N_17790,N_15601,N_12582);
or U17791 (N_17791,N_12520,N_15639);
or U17792 (N_17792,N_15513,N_13318);
and U17793 (N_17793,N_14646,N_15585);
nand U17794 (N_17794,N_12245,N_12562);
nor U17795 (N_17795,N_15252,N_13416);
and U17796 (N_17796,N_13113,N_15227);
or U17797 (N_17797,N_14214,N_12066);
nor U17798 (N_17798,N_14039,N_13583);
or U17799 (N_17799,N_13137,N_12855);
and U17800 (N_17800,N_13874,N_12311);
and U17801 (N_17801,N_12509,N_13988);
nor U17802 (N_17802,N_12707,N_14631);
and U17803 (N_17803,N_12668,N_12406);
xnor U17804 (N_17804,N_13445,N_15298);
nand U17805 (N_17805,N_13786,N_15472);
nand U17806 (N_17806,N_12278,N_12986);
nor U17807 (N_17807,N_14333,N_13494);
nor U17808 (N_17808,N_12393,N_14648);
nand U17809 (N_17809,N_13723,N_15912);
xor U17810 (N_17810,N_15587,N_14300);
nand U17811 (N_17811,N_12015,N_13649);
or U17812 (N_17812,N_14040,N_14784);
nand U17813 (N_17813,N_12769,N_13527);
xnor U17814 (N_17814,N_14957,N_14872);
or U17815 (N_17815,N_14740,N_14509);
nor U17816 (N_17816,N_14408,N_14893);
nand U17817 (N_17817,N_12947,N_14996);
nand U17818 (N_17818,N_15311,N_12352);
and U17819 (N_17819,N_15101,N_13646);
or U17820 (N_17820,N_15414,N_14521);
and U17821 (N_17821,N_14983,N_15586);
nand U17822 (N_17822,N_15296,N_14219);
nand U17823 (N_17823,N_13154,N_15432);
or U17824 (N_17824,N_13795,N_12079);
and U17825 (N_17825,N_13910,N_14823);
nand U17826 (N_17826,N_15024,N_12856);
or U17827 (N_17827,N_12775,N_14247);
nor U17828 (N_17828,N_14005,N_13030);
or U17829 (N_17829,N_14492,N_14782);
and U17830 (N_17830,N_14465,N_15438);
or U17831 (N_17831,N_13605,N_14934);
nand U17832 (N_17832,N_15460,N_13498);
nand U17833 (N_17833,N_12749,N_14127);
nand U17834 (N_17834,N_12347,N_13648);
or U17835 (N_17835,N_14815,N_12114);
nand U17836 (N_17836,N_14867,N_13057);
xor U17837 (N_17837,N_13364,N_15471);
nand U17838 (N_17838,N_13194,N_12552);
nor U17839 (N_17839,N_14009,N_12782);
and U17840 (N_17840,N_13861,N_13232);
xnor U17841 (N_17841,N_15386,N_15641);
and U17842 (N_17842,N_15606,N_14320);
or U17843 (N_17843,N_15580,N_15670);
nand U17844 (N_17844,N_14991,N_15595);
or U17845 (N_17845,N_13562,N_13997);
and U17846 (N_17846,N_13203,N_14460);
or U17847 (N_17847,N_12333,N_13777);
nand U17848 (N_17848,N_14098,N_12433);
nor U17849 (N_17849,N_12862,N_13685);
or U17850 (N_17850,N_15068,N_15886);
and U17851 (N_17851,N_13103,N_14106);
nand U17852 (N_17852,N_14008,N_14493);
nand U17853 (N_17853,N_13917,N_15547);
nor U17854 (N_17854,N_14429,N_15536);
xor U17855 (N_17855,N_15265,N_14162);
nor U17856 (N_17856,N_13371,N_15317);
or U17857 (N_17857,N_12778,N_13582);
and U17858 (N_17858,N_13830,N_15274);
nand U17859 (N_17859,N_13001,N_14877);
nand U17860 (N_17860,N_12419,N_14463);
or U17861 (N_17861,N_13529,N_13933);
and U17862 (N_17862,N_15876,N_15724);
xor U17863 (N_17863,N_12806,N_15544);
or U17864 (N_17864,N_14343,N_15740);
nand U17865 (N_17865,N_13460,N_13816);
nor U17866 (N_17866,N_15866,N_14444);
xnor U17867 (N_17867,N_12328,N_13286);
nand U17868 (N_17868,N_12912,N_12939);
and U17869 (N_17869,N_15941,N_12847);
and U17870 (N_17870,N_12869,N_14632);
nand U17871 (N_17871,N_13871,N_14692);
nor U17872 (N_17872,N_13251,N_15511);
xor U17873 (N_17873,N_12821,N_14854);
nand U17874 (N_17874,N_14296,N_13099);
or U17875 (N_17875,N_15066,N_15804);
nand U17876 (N_17876,N_15566,N_13452);
nand U17877 (N_17877,N_12230,N_15166);
nor U17878 (N_17878,N_13548,N_12498);
nor U17879 (N_17879,N_15747,N_15574);
nor U17880 (N_17880,N_15904,N_14718);
xnor U17881 (N_17881,N_12170,N_14767);
nor U17882 (N_17882,N_14351,N_12714);
and U17883 (N_17883,N_12108,N_14736);
or U17884 (N_17884,N_14086,N_15320);
nor U17885 (N_17885,N_13273,N_12537);
nand U17886 (N_17886,N_13951,N_13929);
nor U17887 (N_17887,N_12921,N_12521);
xnor U17888 (N_17888,N_13429,N_14387);
and U17889 (N_17889,N_14080,N_12943);
nand U17890 (N_17890,N_13307,N_13189);
nand U17891 (N_17891,N_12810,N_13827);
and U17892 (N_17892,N_15940,N_15671);
nand U17893 (N_17893,N_13770,N_14397);
nand U17894 (N_17894,N_13627,N_12467);
nor U17895 (N_17895,N_15236,N_14026);
or U17896 (N_17896,N_15044,N_14617);
nand U17897 (N_17897,N_15792,N_15946);
and U17898 (N_17898,N_13101,N_13798);
and U17899 (N_17899,N_15168,N_14419);
or U17900 (N_17900,N_12051,N_13750);
or U17901 (N_17901,N_15497,N_14070);
and U17902 (N_17902,N_15809,N_12671);
and U17903 (N_17903,N_15240,N_12335);
or U17904 (N_17904,N_13556,N_13479);
nor U17905 (N_17905,N_13921,N_13506);
nor U17906 (N_17906,N_12934,N_13497);
or U17907 (N_17907,N_12482,N_15610);
nand U17908 (N_17908,N_14564,N_14535);
nand U17909 (N_17909,N_14048,N_15558);
nor U17910 (N_17910,N_12719,N_15573);
or U17911 (N_17911,N_12848,N_14755);
and U17912 (N_17912,N_14257,N_12882);
nand U17913 (N_17913,N_12872,N_14126);
nand U17914 (N_17914,N_14662,N_15875);
and U17915 (N_17915,N_14155,N_14297);
nand U17916 (N_17916,N_13518,N_14716);
nor U17917 (N_17917,N_13165,N_13966);
and U17918 (N_17918,N_12178,N_12611);
and U17919 (N_17919,N_15600,N_15569);
or U17920 (N_17920,N_12676,N_12405);
and U17921 (N_17921,N_14882,N_13280);
xor U17922 (N_17922,N_13432,N_15340);
and U17923 (N_17923,N_12553,N_15417);
and U17924 (N_17924,N_15157,N_13408);
nor U17925 (N_17925,N_15494,N_12505);
nand U17926 (N_17926,N_15657,N_13986);
nor U17927 (N_17927,N_15287,N_15490);
nor U17928 (N_17928,N_12589,N_13403);
nor U17929 (N_17929,N_15103,N_13736);
and U17930 (N_17930,N_13901,N_15337);
or U17931 (N_17931,N_14644,N_13718);
xnor U17932 (N_17932,N_14355,N_14143);
xnor U17933 (N_17933,N_13564,N_14164);
nand U17934 (N_17934,N_13178,N_15441);
nor U17935 (N_17935,N_13152,N_13887);
nor U17936 (N_17936,N_15889,N_12735);
and U17937 (N_17937,N_13243,N_13393);
nor U17938 (N_17938,N_12647,N_15388);
or U17939 (N_17939,N_15750,N_14204);
nand U17940 (N_17940,N_14680,N_15199);
or U17941 (N_17941,N_15856,N_12361);
or U17942 (N_17942,N_15546,N_14825);
and U17943 (N_17943,N_14424,N_12794);
or U17944 (N_17944,N_14000,N_13761);
and U17945 (N_17945,N_13930,N_13238);
xnor U17946 (N_17946,N_12567,N_15203);
nor U17947 (N_17947,N_12705,N_14019);
xnor U17948 (N_17948,N_15535,N_12418);
and U17949 (N_17949,N_15599,N_13733);
or U17950 (N_17950,N_12247,N_13085);
nand U17951 (N_17951,N_15127,N_13844);
and U17952 (N_17952,N_12588,N_15549);
and U17953 (N_17953,N_12171,N_14187);
nand U17954 (N_17954,N_12314,N_15499);
nor U17955 (N_17955,N_12604,N_14733);
nor U17956 (N_17956,N_12752,N_12485);
and U17957 (N_17957,N_13150,N_12341);
nor U17958 (N_17958,N_13586,N_12238);
and U17959 (N_17959,N_14018,N_15831);
nor U17960 (N_17960,N_12271,N_13701);
nand U17961 (N_17961,N_13448,N_12483);
and U17962 (N_17962,N_13486,N_14344);
and U17963 (N_17963,N_13796,N_15669);
and U17964 (N_17964,N_15353,N_13436);
and U17965 (N_17965,N_13380,N_15701);
nor U17966 (N_17966,N_15223,N_15014);
nand U17967 (N_17967,N_12865,N_15446);
and U17968 (N_17968,N_15348,N_13108);
xor U17969 (N_17969,N_15507,N_15741);
nor U17970 (N_17970,N_13757,N_13365);
and U17971 (N_17971,N_14061,N_13100);
xnor U17972 (N_17972,N_13539,N_15846);
and U17973 (N_17973,N_12801,N_12322);
nor U17974 (N_17974,N_14528,N_15647);
nor U17975 (N_17975,N_15247,N_14129);
nor U17976 (N_17976,N_15829,N_14478);
and U17977 (N_17977,N_14010,N_13372);
nand U17978 (N_17978,N_13499,N_14612);
nand U17979 (N_17979,N_12261,N_12319);
nor U17980 (N_17980,N_14942,N_13083);
nor U17981 (N_17981,N_14495,N_13292);
nand U17982 (N_17982,N_15737,N_14651);
and U17983 (N_17983,N_12141,N_15933);
nand U17984 (N_17984,N_15749,N_13846);
nor U17985 (N_17985,N_15835,N_12818);
and U17986 (N_17986,N_14590,N_13163);
and U17987 (N_17987,N_15083,N_15128);
xor U17988 (N_17988,N_13321,N_14306);
xor U17989 (N_17989,N_13608,N_15326);
xnor U17990 (N_17990,N_13484,N_12837);
nor U17991 (N_17991,N_13963,N_13221);
nor U17992 (N_17992,N_14426,N_13018);
nor U17993 (N_17993,N_12380,N_15567);
nor U17994 (N_17994,N_13072,N_15556);
and U17995 (N_17995,N_12101,N_15515);
nand U17996 (N_17996,N_13934,N_12027);
and U17997 (N_17997,N_14382,N_15772);
nor U17998 (N_17998,N_13696,N_14638);
and U17999 (N_17999,N_13881,N_15807);
and U18000 (N_18000,N_12799,N_12688);
xor U18001 (N_18001,N_12266,N_12684);
or U18002 (N_18002,N_12552,N_15981);
or U18003 (N_18003,N_15009,N_14821);
or U18004 (N_18004,N_15146,N_15876);
nor U18005 (N_18005,N_13157,N_12939);
and U18006 (N_18006,N_14364,N_12970);
nand U18007 (N_18007,N_15920,N_13847);
or U18008 (N_18008,N_13569,N_14697);
nor U18009 (N_18009,N_13941,N_12640);
nor U18010 (N_18010,N_13146,N_12088);
or U18011 (N_18011,N_14069,N_12718);
and U18012 (N_18012,N_15865,N_14805);
and U18013 (N_18013,N_15197,N_15501);
nor U18014 (N_18014,N_15676,N_14522);
nand U18015 (N_18015,N_14417,N_14182);
and U18016 (N_18016,N_13005,N_13122);
or U18017 (N_18017,N_12512,N_12605);
xnor U18018 (N_18018,N_13564,N_13457);
nor U18019 (N_18019,N_12012,N_14809);
xnor U18020 (N_18020,N_15760,N_15317);
and U18021 (N_18021,N_13651,N_15780);
or U18022 (N_18022,N_13962,N_14650);
nand U18023 (N_18023,N_15838,N_15785);
or U18024 (N_18024,N_15246,N_13793);
or U18025 (N_18025,N_14851,N_15268);
xor U18026 (N_18026,N_13325,N_15903);
nor U18027 (N_18027,N_15571,N_15787);
or U18028 (N_18028,N_14108,N_15031);
or U18029 (N_18029,N_15408,N_15448);
nor U18030 (N_18030,N_12211,N_14635);
nand U18031 (N_18031,N_12535,N_14896);
nand U18032 (N_18032,N_14336,N_12165);
xor U18033 (N_18033,N_12835,N_14285);
and U18034 (N_18034,N_13436,N_14096);
nor U18035 (N_18035,N_14020,N_12679);
and U18036 (N_18036,N_13305,N_15885);
nand U18037 (N_18037,N_14699,N_13123);
and U18038 (N_18038,N_14895,N_15772);
nand U18039 (N_18039,N_12313,N_15029);
nand U18040 (N_18040,N_15246,N_15578);
nor U18041 (N_18041,N_15870,N_12853);
nor U18042 (N_18042,N_12583,N_12399);
nor U18043 (N_18043,N_12088,N_15335);
nor U18044 (N_18044,N_13057,N_15095);
nand U18045 (N_18045,N_12037,N_12251);
nand U18046 (N_18046,N_15696,N_13968);
and U18047 (N_18047,N_13054,N_13825);
and U18048 (N_18048,N_13741,N_13184);
xor U18049 (N_18049,N_14317,N_12137);
or U18050 (N_18050,N_14162,N_12634);
or U18051 (N_18051,N_13787,N_15372);
nand U18052 (N_18052,N_12859,N_15097);
xor U18053 (N_18053,N_12205,N_15889);
nand U18054 (N_18054,N_15373,N_13255);
nor U18055 (N_18055,N_15990,N_12082);
nand U18056 (N_18056,N_13211,N_12569);
nor U18057 (N_18057,N_12522,N_14876);
nand U18058 (N_18058,N_13413,N_13233);
nand U18059 (N_18059,N_13942,N_15593);
and U18060 (N_18060,N_12497,N_12403);
and U18061 (N_18061,N_13780,N_14794);
or U18062 (N_18062,N_14590,N_13808);
nand U18063 (N_18063,N_13597,N_13967);
and U18064 (N_18064,N_12224,N_14344);
nand U18065 (N_18065,N_15203,N_12933);
nor U18066 (N_18066,N_14752,N_13585);
and U18067 (N_18067,N_15077,N_15340);
or U18068 (N_18068,N_14856,N_14498);
nor U18069 (N_18069,N_12769,N_12169);
nand U18070 (N_18070,N_12371,N_15021);
and U18071 (N_18071,N_14886,N_13818);
nand U18072 (N_18072,N_12361,N_13804);
and U18073 (N_18073,N_13193,N_13752);
xor U18074 (N_18074,N_13163,N_13273);
and U18075 (N_18075,N_12308,N_14319);
and U18076 (N_18076,N_13758,N_13639);
and U18077 (N_18077,N_12708,N_14390);
or U18078 (N_18078,N_12230,N_13020);
or U18079 (N_18079,N_14824,N_15184);
nand U18080 (N_18080,N_15080,N_14678);
xnor U18081 (N_18081,N_13877,N_12236);
and U18082 (N_18082,N_12000,N_12379);
nand U18083 (N_18083,N_12058,N_13927);
nor U18084 (N_18084,N_13799,N_14530);
or U18085 (N_18085,N_13807,N_14546);
nand U18086 (N_18086,N_13289,N_13833);
nand U18087 (N_18087,N_15392,N_12671);
nor U18088 (N_18088,N_12628,N_12753);
xor U18089 (N_18089,N_15869,N_12674);
and U18090 (N_18090,N_15249,N_15865);
xnor U18091 (N_18091,N_15992,N_12042);
and U18092 (N_18092,N_13021,N_12627);
xor U18093 (N_18093,N_15039,N_12167);
and U18094 (N_18094,N_13431,N_12597);
and U18095 (N_18095,N_13890,N_13168);
nand U18096 (N_18096,N_13037,N_14894);
nor U18097 (N_18097,N_15048,N_12793);
xor U18098 (N_18098,N_15250,N_12467);
nor U18099 (N_18099,N_14667,N_12295);
nand U18100 (N_18100,N_12499,N_14063);
and U18101 (N_18101,N_14466,N_14789);
or U18102 (N_18102,N_15170,N_14212);
and U18103 (N_18103,N_12953,N_14349);
nand U18104 (N_18104,N_14777,N_12152);
nor U18105 (N_18105,N_13296,N_14754);
nand U18106 (N_18106,N_14180,N_13248);
nor U18107 (N_18107,N_12850,N_14162);
xnor U18108 (N_18108,N_14031,N_12024);
nor U18109 (N_18109,N_15294,N_12884);
nand U18110 (N_18110,N_13178,N_12812);
or U18111 (N_18111,N_13100,N_12170);
and U18112 (N_18112,N_15533,N_12202);
and U18113 (N_18113,N_15657,N_14112);
xnor U18114 (N_18114,N_14052,N_13642);
or U18115 (N_18115,N_14260,N_14569);
nor U18116 (N_18116,N_12606,N_12361);
xnor U18117 (N_18117,N_12120,N_15774);
and U18118 (N_18118,N_15716,N_14378);
nor U18119 (N_18119,N_13777,N_13468);
nor U18120 (N_18120,N_13429,N_12387);
or U18121 (N_18121,N_14576,N_15350);
nor U18122 (N_18122,N_14742,N_15120);
nand U18123 (N_18123,N_14095,N_13140);
nor U18124 (N_18124,N_13190,N_14681);
and U18125 (N_18125,N_15480,N_15857);
nor U18126 (N_18126,N_15729,N_15091);
or U18127 (N_18127,N_15131,N_13190);
nor U18128 (N_18128,N_13877,N_15377);
nor U18129 (N_18129,N_13476,N_13014);
nand U18130 (N_18130,N_12278,N_14438);
or U18131 (N_18131,N_12758,N_14896);
and U18132 (N_18132,N_14876,N_12924);
or U18133 (N_18133,N_14238,N_13263);
nor U18134 (N_18134,N_12868,N_12174);
and U18135 (N_18135,N_14743,N_14384);
xnor U18136 (N_18136,N_12867,N_13366);
and U18137 (N_18137,N_12780,N_15618);
xnor U18138 (N_18138,N_15612,N_13064);
nand U18139 (N_18139,N_13369,N_13329);
nand U18140 (N_18140,N_15524,N_15937);
and U18141 (N_18141,N_13491,N_14879);
nor U18142 (N_18142,N_15517,N_13120);
nand U18143 (N_18143,N_13610,N_15651);
xor U18144 (N_18144,N_13059,N_14341);
and U18145 (N_18145,N_15175,N_15228);
xor U18146 (N_18146,N_15189,N_14260);
or U18147 (N_18147,N_12471,N_13631);
and U18148 (N_18148,N_15121,N_13254);
nor U18149 (N_18149,N_12241,N_12254);
nand U18150 (N_18150,N_14898,N_14750);
nand U18151 (N_18151,N_13933,N_12778);
xor U18152 (N_18152,N_14921,N_12554);
nor U18153 (N_18153,N_15624,N_14999);
or U18154 (N_18154,N_13017,N_15316);
nand U18155 (N_18155,N_13714,N_13670);
and U18156 (N_18156,N_15148,N_15764);
and U18157 (N_18157,N_15648,N_14051);
and U18158 (N_18158,N_14630,N_13500);
and U18159 (N_18159,N_13433,N_12857);
or U18160 (N_18160,N_12808,N_12804);
nor U18161 (N_18161,N_15198,N_12888);
xor U18162 (N_18162,N_14024,N_15054);
xor U18163 (N_18163,N_12429,N_15652);
nor U18164 (N_18164,N_13014,N_12514);
nor U18165 (N_18165,N_15062,N_14971);
or U18166 (N_18166,N_15354,N_14719);
xor U18167 (N_18167,N_13031,N_14209);
xnor U18168 (N_18168,N_13349,N_13021);
or U18169 (N_18169,N_14252,N_13397);
xnor U18170 (N_18170,N_13632,N_13294);
nor U18171 (N_18171,N_15169,N_12475);
and U18172 (N_18172,N_13503,N_12477);
xor U18173 (N_18173,N_14954,N_12189);
nand U18174 (N_18174,N_14966,N_14017);
and U18175 (N_18175,N_13294,N_12478);
nand U18176 (N_18176,N_12930,N_15586);
xnor U18177 (N_18177,N_12074,N_15397);
nor U18178 (N_18178,N_14145,N_12681);
nor U18179 (N_18179,N_15241,N_15562);
nand U18180 (N_18180,N_12772,N_14450);
nor U18181 (N_18181,N_15913,N_13850);
or U18182 (N_18182,N_13304,N_12054);
and U18183 (N_18183,N_12194,N_12434);
nor U18184 (N_18184,N_15660,N_15404);
nor U18185 (N_18185,N_14152,N_14881);
nor U18186 (N_18186,N_14193,N_12164);
and U18187 (N_18187,N_12837,N_14426);
or U18188 (N_18188,N_15251,N_13825);
nor U18189 (N_18189,N_13930,N_12411);
xnor U18190 (N_18190,N_12769,N_14473);
xor U18191 (N_18191,N_14938,N_12450);
and U18192 (N_18192,N_13747,N_15310);
or U18193 (N_18193,N_13894,N_12253);
xor U18194 (N_18194,N_12867,N_13738);
nand U18195 (N_18195,N_14653,N_12918);
and U18196 (N_18196,N_14407,N_12433);
and U18197 (N_18197,N_12670,N_14835);
or U18198 (N_18198,N_13720,N_13403);
nand U18199 (N_18199,N_12097,N_15977);
xnor U18200 (N_18200,N_15248,N_12871);
nand U18201 (N_18201,N_12186,N_14666);
nor U18202 (N_18202,N_13484,N_12755);
nand U18203 (N_18203,N_14702,N_13225);
or U18204 (N_18204,N_13373,N_12638);
nand U18205 (N_18205,N_13977,N_13620);
nor U18206 (N_18206,N_12026,N_13781);
and U18207 (N_18207,N_12432,N_12634);
nor U18208 (N_18208,N_14401,N_15344);
nand U18209 (N_18209,N_15887,N_14324);
nor U18210 (N_18210,N_15044,N_14727);
and U18211 (N_18211,N_13756,N_14018);
and U18212 (N_18212,N_12786,N_13106);
xor U18213 (N_18213,N_12694,N_12258);
nor U18214 (N_18214,N_14188,N_12975);
nor U18215 (N_18215,N_15279,N_12779);
nor U18216 (N_18216,N_12945,N_15965);
nand U18217 (N_18217,N_12497,N_13652);
nor U18218 (N_18218,N_15264,N_12454);
nor U18219 (N_18219,N_13155,N_14213);
or U18220 (N_18220,N_15326,N_14086);
nand U18221 (N_18221,N_13412,N_13226);
and U18222 (N_18222,N_12264,N_13010);
and U18223 (N_18223,N_13187,N_14702);
or U18224 (N_18224,N_14965,N_13297);
nand U18225 (N_18225,N_14572,N_13997);
nor U18226 (N_18226,N_15366,N_14621);
and U18227 (N_18227,N_15288,N_12397);
xor U18228 (N_18228,N_13581,N_12212);
and U18229 (N_18229,N_12690,N_14385);
nor U18230 (N_18230,N_15080,N_13561);
xor U18231 (N_18231,N_15878,N_14158);
nor U18232 (N_18232,N_14590,N_13953);
and U18233 (N_18233,N_15372,N_12819);
nand U18234 (N_18234,N_12042,N_12669);
nand U18235 (N_18235,N_13150,N_12147);
and U18236 (N_18236,N_12459,N_15663);
or U18237 (N_18237,N_15522,N_13624);
nand U18238 (N_18238,N_12623,N_12869);
or U18239 (N_18239,N_15215,N_12551);
and U18240 (N_18240,N_13533,N_14956);
nor U18241 (N_18241,N_15059,N_13006);
nor U18242 (N_18242,N_13214,N_14430);
xnor U18243 (N_18243,N_14161,N_14380);
and U18244 (N_18244,N_12351,N_13143);
nor U18245 (N_18245,N_13120,N_15415);
xor U18246 (N_18246,N_14955,N_12375);
and U18247 (N_18247,N_13537,N_15437);
or U18248 (N_18248,N_15514,N_15822);
and U18249 (N_18249,N_14148,N_12121);
nand U18250 (N_18250,N_14645,N_13967);
and U18251 (N_18251,N_12685,N_12074);
xnor U18252 (N_18252,N_14904,N_13224);
xnor U18253 (N_18253,N_12326,N_15351);
nand U18254 (N_18254,N_14204,N_12409);
and U18255 (N_18255,N_12919,N_13098);
and U18256 (N_18256,N_15558,N_13334);
or U18257 (N_18257,N_14274,N_13244);
and U18258 (N_18258,N_15864,N_14175);
nor U18259 (N_18259,N_12812,N_12671);
and U18260 (N_18260,N_14816,N_12779);
nand U18261 (N_18261,N_15910,N_12622);
or U18262 (N_18262,N_15864,N_12072);
and U18263 (N_18263,N_13275,N_13789);
or U18264 (N_18264,N_12054,N_13655);
and U18265 (N_18265,N_13657,N_13082);
xnor U18266 (N_18266,N_15365,N_15271);
nand U18267 (N_18267,N_15256,N_12240);
and U18268 (N_18268,N_13316,N_12922);
nor U18269 (N_18269,N_15602,N_12205);
nand U18270 (N_18270,N_15260,N_14335);
and U18271 (N_18271,N_14707,N_13066);
or U18272 (N_18272,N_15075,N_12645);
nor U18273 (N_18273,N_12268,N_12347);
and U18274 (N_18274,N_13771,N_15673);
nand U18275 (N_18275,N_12568,N_13174);
nand U18276 (N_18276,N_15851,N_12224);
and U18277 (N_18277,N_13787,N_13607);
or U18278 (N_18278,N_12703,N_14852);
nor U18279 (N_18279,N_13128,N_13006);
nor U18280 (N_18280,N_15124,N_15027);
or U18281 (N_18281,N_14496,N_13898);
and U18282 (N_18282,N_14830,N_14786);
or U18283 (N_18283,N_12562,N_13931);
and U18284 (N_18284,N_13778,N_15060);
nor U18285 (N_18285,N_15741,N_13095);
or U18286 (N_18286,N_14403,N_12516);
nor U18287 (N_18287,N_12118,N_12397);
xnor U18288 (N_18288,N_12050,N_15850);
or U18289 (N_18289,N_14754,N_15859);
nor U18290 (N_18290,N_13926,N_15040);
nor U18291 (N_18291,N_13841,N_12102);
nand U18292 (N_18292,N_14724,N_13560);
xor U18293 (N_18293,N_12953,N_12987);
nand U18294 (N_18294,N_13389,N_15237);
nor U18295 (N_18295,N_14041,N_12937);
nor U18296 (N_18296,N_13396,N_15219);
and U18297 (N_18297,N_12742,N_12537);
nor U18298 (N_18298,N_13187,N_12339);
xor U18299 (N_18299,N_12747,N_15307);
nand U18300 (N_18300,N_15597,N_14108);
xor U18301 (N_18301,N_12991,N_13811);
or U18302 (N_18302,N_12195,N_13202);
nor U18303 (N_18303,N_13583,N_13301);
nand U18304 (N_18304,N_15802,N_13496);
and U18305 (N_18305,N_15186,N_13633);
and U18306 (N_18306,N_13800,N_15261);
and U18307 (N_18307,N_13954,N_13631);
or U18308 (N_18308,N_13127,N_15224);
nand U18309 (N_18309,N_12365,N_14518);
and U18310 (N_18310,N_12652,N_13627);
nor U18311 (N_18311,N_14073,N_14207);
and U18312 (N_18312,N_13273,N_14895);
nand U18313 (N_18313,N_14856,N_14216);
and U18314 (N_18314,N_14521,N_15520);
nand U18315 (N_18315,N_12712,N_12265);
nand U18316 (N_18316,N_12110,N_13168);
or U18317 (N_18317,N_13218,N_12531);
xnor U18318 (N_18318,N_13437,N_13463);
or U18319 (N_18319,N_15578,N_13430);
nor U18320 (N_18320,N_12628,N_13995);
nand U18321 (N_18321,N_12003,N_13832);
and U18322 (N_18322,N_13569,N_12450);
and U18323 (N_18323,N_15677,N_14744);
nand U18324 (N_18324,N_15932,N_13391);
nand U18325 (N_18325,N_12334,N_13706);
and U18326 (N_18326,N_12333,N_12481);
nor U18327 (N_18327,N_13183,N_12517);
and U18328 (N_18328,N_14705,N_15081);
or U18329 (N_18329,N_14742,N_13249);
nor U18330 (N_18330,N_15910,N_14406);
and U18331 (N_18331,N_12233,N_13895);
nor U18332 (N_18332,N_13871,N_14199);
nor U18333 (N_18333,N_15073,N_12753);
or U18334 (N_18334,N_12529,N_14088);
xnor U18335 (N_18335,N_13207,N_12838);
nor U18336 (N_18336,N_12949,N_14799);
nand U18337 (N_18337,N_13871,N_12614);
or U18338 (N_18338,N_12300,N_14348);
or U18339 (N_18339,N_12142,N_14688);
nor U18340 (N_18340,N_15390,N_14605);
nor U18341 (N_18341,N_13609,N_12837);
and U18342 (N_18342,N_15703,N_14997);
and U18343 (N_18343,N_12908,N_15035);
and U18344 (N_18344,N_15439,N_13931);
or U18345 (N_18345,N_12257,N_15258);
xor U18346 (N_18346,N_15189,N_15467);
nor U18347 (N_18347,N_13193,N_15806);
or U18348 (N_18348,N_13124,N_13714);
nand U18349 (N_18349,N_12483,N_12369);
nor U18350 (N_18350,N_15069,N_14420);
and U18351 (N_18351,N_13594,N_12929);
and U18352 (N_18352,N_13339,N_13016);
and U18353 (N_18353,N_12063,N_12598);
and U18354 (N_18354,N_15567,N_15973);
nand U18355 (N_18355,N_13268,N_12578);
nor U18356 (N_18356,N_14191,N_13944);
nand U18357 (N_18357,N_14972,N_12482);
and U18358 (N_18358,N_15854,N_14897);
xnor U18359 (N_18359,N_15005,N_14900);
xor U18360 (N_18360,N_14443,N_14968);
nor U18361 (N_18361,N_13669,N_14600);
and U18362 (N_18362,N_15044,N_12311);
nand U18363 (N_18363,N_13836,N_15128);
and U18364 (N_18364,N_13495,N_12572);
and U18365 (N_18365,N_14622,N_12124);
or U18366 (N_18366,N_12467,N_14674);
and U18367 (N_18367,N_12423,N_13117);
or U18368 (N_18368,N_13413,N_15891);
or U18369 (N_18369,N_15713,N_12878);
nor U18370 (N_18370,N_15917,N_14137);
or U18371 (N_18371,N_14737,N_13268);
nand U18372 (N_18372,N_12613,N_12327);
nand U18373 (N_18373,N_15240,N_13106);
nor U18374 (N_18374,N_13533,N_13885);
and U18375 (N_18375,N_12514,N_14277);
and U18376 (N_18376,N_13954,N_15719);
and U18377 (N_18377,N_12178,N_12282);
nor U18378 (N_18378,N_15258,N_12962);
and U18379 (N_18379,N_13878,N_14868);
nand U18380 (N_18380,N_12400,N_14445);
or U18381 (N_18381,N_14388,N_14491);
and U18382 (N_18382,N_13081,N_12527);
and U18383 (N_18383,N_14739,N_12764);
and U18384 (N_18384,N_14702,N_14296);
nand U18385 (N_18385,N_14917,N_12424);
or U18386 (N_18386,N_14020,N_12055);
xor U18387 (N_18387,N_12646,N_14045);
nor U18388 (N_18388,N_12710,N_13672);
xor U18389 (N_18389,N_12133,N_14886);
nor U18390 (N_18390,N_13403,N_14794);
or U18391 (N_18391,N_14261,N_12662);
nor U18392 (N_18392,N_14537,N_12699);
or U18393 (N_18393,N_14392,N_13541);
or U18394 (N_18394,N_12548,N_15703);
nor U18395 (N_18395,N_15838,N_13044);
and U18396 (N_18396,N_12442,N_12341);
nor U18397 (N_18397,N_14296,N_13639);
xor U18398 (N_18398,N_15629,N_12487);
and U18399 (N_18399,N_15085,N_15570);
nor U18400 (N_18400,N_15829,N_15090);
nand U18401 (N_18401,N_15313,N_14938);
or U18402 (N_18402,N_12322,N_13849);
nand U18403 (N_18403,N_15538,N_12927);
or U18404 (N_18404,N_13037,N_15971);
nor U18405 (N_18405,N_14373,N_12457);
nand U18406 (N_18406,N_13957,N_15198);
nand U18407 (N_18407,N_14623,N_14894);
or U18408 (N_18408,N_14789,N_14048);
or U18409 (N_18409,N_14806,N_13847);
and U18410 (N_18410,N_14852,N_13701);
and U18411 (N_18411,N_12527,N_15554);
nor U18412 (N_18412,N_13874,N_14489);
or U18413 (N_18413,N_12257,N_15936);
nor U18414 (N_18414,N_15036,N_15238);
and U18415 (N_18415,N_13539,N_13916);
nor U18416 (N_18416,N_12742,N_12555);
or U18417 (N_18417,N_15343,N_15145);
and U18418 (N_18418,N_15651,N_15096);
and U18419 (N_18419,N_12811,N_14113);
xnor U18420 (N_18420,N_15605,N_15238);
nand U18421 (N_18421,N_15376,N_14559);
nor U18422 (N_18422,N_12229,N_13470);
or U18423 (N_18423,N_13765,N_14907);
nor U18424 (N_18424,N_12873,N_15669);
nand U18425 (N_18425,N_15444,N_14814);
nor U18426 (N_18426,N_12039,N_14234);
and U18427 (N_18427,N_15127,N_13574);
or U18428 (N_18428,N_13778,N_15380);
or U18429 (N_18429,N_12194,N_14209);
nor U18430 (N_18430,N_14926,N_13053);
nand U18431 (N_18431,N_12579,N_13629);
and U18432 (N_18432,N_12494,N_15967);
nor U18433 (N_18433,N_12152,N_13774);
nor U18434 (N_18434,N_13093,N_13514);
nor U18435 (N_18435,N_14638,N_12241);
nand U18436 (N_18436,N_14697,N_12274);
or U18437 (N_18437,N_14889,N_12701);
or U18438 (N_18438,N_13962,N_13671);
and U18439 (N_18439,N_12873,N_13704);
or U18440 (N_18440,N_13595,N_13441);
or U18441 (N_18441,N_15122,N_13847);
nor U18442 (N_18442,N_12809,N_12995);
nor U18443 (N_18443,N_12194,N_13663);
and U18444 (N_18444,N_15412,N_12239);
or U18445 (N_18445,N_15107,N_15833);
nand U18446 (N_18446,N_15819,N_14233);
nor U18447 (N_18447,N_14264,N_14828);
or U18448 (N_18448,N_15929,N_14694);
nand U18449 (N_18449,N_12496,N_12467);
nand U18450 (N_18450,N_14354,N_12550);
nor U18451 (N_18451,N_13248,N_14593);
nand U18452 (N_18452,N_14602,N_15649);
or U18453 (N_18453,N_12069,N_12847);
nand U18454 (N_18454,N_13358,N_15934);
and U18455 (N_18455,N_13703,N_14051);
and U18456 (N_18456,N_12502,N_13631);
and U18457 (N_18457,N_15641,N_13965);
xor U18458 (N_18458,N_13863,N_14187);
nor U18459 (N_18459,N_12573,N_13652);
nor U18460 (N_18460,N_15341,N_15995);
or U18461 (N_18461,N_12967,N_12575);
or U18462 (N_18462,N_13922,N_12852);
or U18463 (N_18463,N_14020,N_12128);
and U18464 (N_18464,N_12941,N_14937);
nor U18465 (N_18465,N_12998,N_13443);
and U18466 (N_18466,N_13624,N_15438);
nor U18467 (N_18467,N_13008,N_12774);
or U18468 (N_18468,N_13146,N_14030);
nor U18469 (N_18469,N_15660,N_15024);
nor U18470 (N_18470,N_12699,N_12328);
or U18471 (N_18471,N_12030,N_12627);
and U18472 (N_18472,N_15824,N_12649);
nor U18473 (N_18473,N_13265,N_15203);
nor U18474 (N_18474,N_14531,N_12350);
nor U18475 (N_18475,N_12512,N_14628);
nand U18476 (N_18476,N_15440,N_12497);
nor U18477 (N_18477,N_15665,N_12599);
and U18478 (N_18478,N_12872,N_14300);
or U18479 (N_18479,N_13622,N_14423);
or U18480 (N_18480,N_14717,N_15968);
and U18481 (N_18481,N_15425,N_15312);
or U18482 (N_18482,N_15279,N_13077);
and U18483 (N_18483,N_14933,N_13982);
nand U18484 (N_18484,N_13672,N_13847);
or U18485 (N_18485,N_12457,N_14489);
xnor U18486 (N_18486,N_14630,N_15348);
nor U18487 (N_18487,N_12743,N_14170);
and U18488 (N_18488,N_15225,N_12769);
nor U18489 (N_18489,N_12232,N_15728);
or U18490 (N_18490,N_15960,N_15629);
nor U18491 (N_18491,N_12950,N_15313);
nand U18492 (N_18492,N_13185,N_13579);
nor U18493 (N_18493,N_13923,N_14334);
and U18494 (N_18494,N_15455,N_14559);
nor U18495 (N_18495,N_15902,N_14743);
and U18496 (N_18496,N_13200,N_13592);
and U18497 (N_18497,N_12735,N_13041);
nand U18498 (N_18498,N_12986,N_12654);
or U18499 (N_18499,N_15410,N_12859);
nor U18500 (N_18500,N_13234,N_13575);
nand U18501 (N_18501,N_14977,N_12036);
nand U18502 (N_18502,N_14931,N_14065);
or U18503 (N_18503,N_12247,N_13597);
nand U18504 (N_18504,N_14967,N_14713);
or U18505 (N_18505,N_12877,N_14254);
nor U18506 (N_18506,N_13566,N_14178);
or U18507 (N_18507,N_14530,N_13894);
nand U18508 (N_18508,N_15875,N_14774);
xnor U18509 (N_18509,N_15495,N_14671);
nand U18510 (N_18510,N_14879,N_12145);
and U18511 (N_18511,N_12123,N_14985);
nand U18512 (N_18512,N_13239,N_13575);
or U18513 (N_18513,N_15800,N_14780);
xor U18514 (N_18514,N_13896,N_13245);
xnor U18515 (N_18515,N_12624,N_15963);
and U18516 (N_18516,N_14876,N_12592);
or U18517 (N_18517,N_12596,N_14235);
or U18518 (N_18518,N_15901,N_15313);
nor U18519 (N_18519,N_12886,N_13480);
and U18520 (N_18520,N_13100,N_15850);
and U18521 (N_18521,N_14068,N_14846);
or U18522 (N_18522,N_15351,N_13690);
and U18523 (N_18523,N_13941,N_13699);
and U18524 (N_18524,N_13399,N_15513);
nor U18525 (N_18525,N_14167,N_12511);
and U18526 (N_18526,N_14779,N_14731);
nand U18527 (N_18527,N_14220,N_12386);
nor U18528 (N_18528,N_13847,N_15861);
and U18529 (N_18529,N_12964,N_14809);
and U18530 (N_18530,N_15899,N_12699);
nand U18531 (N_18531,N_15335,N_15538);
nor U18532 (N_18532,N_13518,N_14953);
nand U18533 (N_18533,N_12111,N_14057);
or U18534 (N_18534,N_14278,N_14698);
and U18535 (N_18535,N_12769,N_14130);
and U18536 (N_18536,N_12179,N_13359);
nor U18537 (N_18537,N_15955,N_13017);
nor U18538 (N_18538,N_15424,N_12321);
nand U18539 (N_18539,N_14467,N_12449);
nand U18540 (N_18540,N_13280,N_13128);
and U18541 (N_18541,N_14522,N_13788);
nand U18542 (N_18542,N_15694,N_13782);
or U18543 (N_18543,N_15284,N_14547);
nand U18544 (N_18544,N_14937,N_14071);
nand U18545 (N_18545,N_13557,N_12496);
or U18546 (N_18546,N_15212,N_12150);
nand U18547 (N_18547,N_13089,N_12165);
nor U18548 (N_18548,N_15346,N_15302);
nand U18549 (N_18549,N_15247,N_15380);
xor U18550 (N_18550,N_13985,N_12323);
xnor U18551 (N_18551,N_14718,N_15388);
and U18552 (N_18552,N_12096,N_15941);
nand U18553 (N_18553,N_12832,N_12733);
or U18554 (N_18554,N_13364,N_14160);
xor U18555 (N_18555,N_15992,N_12918);
or U18556 (N_18556,N_15832,N_15140);
nor U18557 (N_18557,N_14407,N_14913);
nor U18558 (N_18558,N_12516,N_14719);
or U18559 (N_18559,N_12968,N_15853);
nand U18560 (N_18560,N_13053,N_15375);
nand U18561 (N_18561,N_14678,N_15928);
nand U18562 (N_18562,N_13455,N_15612);
and U18563 (N_18563,N_12689,N_14994);
nor U18564 (N_18564,N_14876,N_12234);
nor U18565 (N_18565,N_14444,N_15602);
nor U18566 (N_18566,N_15565,N_14790);
xor U18567 (N_18567,N_13853,N_12871);
nand U18568 (N_18568,N_14682,N_13968);
or U18569 (N_18569,N_14255,N_14577);
nand U18570 (N_18570,N_15445,N_15022);
and U18571 (N_18571,N_14495,N_12503);
and U18572 (N_18572,N_14773,N_14997);
or U18573 (N_18573,N_14500,N_12976);
and U18574 (N_18574,N_13386,N_15323);
nand U18575 (N_18575,N_15349,N_12232);
nand U18576 (N_18576,N_15061,N_15641);
nand U18577 (N_18577,N_14403,N_13263);
nand U18578 (N_18578,N_12485,N_13604);
nand U18579 (N_18579,N_12679,N_14763);
and U18580 (N_18580,N_12483,N_15424);
xnor U18581 (N_18581,N_12297,N_15927);
nor U18582 (N_18582,N_15835,N_15140);
nand U18583 (N_18583,N_13749,N_13461);
and U18584 (N_18584,N_12443,N_14593);
and U18585 (N_18585,N_12853,N_13355);
nor U18586 (N_18586,N_15132,N_12037);
or U18587 (N_18587,N_15549,N_12156);
nand U18588 (N_18588,N_13061,N_12986);
nor U18589 (N_18589,N_15353,N_15766);
nor U18590 (N_18590,N_13831,N_12606);
and U18591 (N_18591,N_14890,N_15558);
nand U18592 (N_18592,N_13155,N_13085);
nand U18593 (N_18593,N_14685,N_13273);
nor U18594 (N_18594,N_13361,N_15267);
nor U18595 (N_18595,N_15670,N_13161);
xor U18596 (N_18596,N_12932,N_15110);
or U18597 (N_18597,N_12507,N_14959);
and U18598 (N_18598,N_15074,N_13884);
or U18599 (N_18599,N_12032,N_13008);
nand U18600 (N_18600,N_14897,N_15530);
xnor U18601 (N_18601,N_15801,N_15162);
and U18602 (N_18602,N_13816,N_12693);
nor U18603 (N_18603,N_14997,N_14971);
nand U18604 (N_18604,N_15736,N_12711);
nor U18605 (N_18605,N_15354,N_12897);
nand U18606 (N_18606,N_14984,N_14600);
nand U18607 (N_18607,N_12951,N_12897);
or U18608 (N_18608,N_13057,N_13033);
nand U18609 (N_18609,N_13696,N_14278);
nand U18610 (N_18610,N_15508,N_15297);
or U18611 (N_18611,N_13975,N_15654);
nand U18612 (N_18612,N_12359,N_15010);
and U18613 (N_18613,N_14567,N_12365);
nand U18614 (N_18614,N_15851,N_13860);
and U18615 (N_18615,N_12804,N_15553);
and U18616 (N_18616,N_13004,N_12221);
and U18617 (N_18617,N_15651,N_13067);
nor U18618 (N_18618,N_14181,N_12630);
and U18619 (N_18619,N_13888,N_13192);
nand U18620 (N_18620,N_14625,N_15862);
and U18621 (N_18621,N_13476,N_15146);
and U18622 (N_18622,N_14344,N_15642);
nor U18623 (N_18623,N_13984,N_12343);
nand U18624 (N_18624,N_13390,N_15637);
xor U18625 (N_18625,N_15749,N_12230);
nor U18626 (N_18626,N_14665,N_13956);
nand U18627 (N_18627,N_15874,N_14404);
or U18628 (N_18628,N_13387,N_12885);
or U18629 (N_18629,N_12872,N_12452);
nor U18630 (N_18630,N_15572,N_14624);
or U18631 (N_18631,N_14585,N_12969);
or U18632 (N_18632,N_15949,N_13291);
and U18633 (N_18633,N_13108,N_12479);
and U18634 (N_18634,N_12922,N_13034);
or U18635 (N_18635,N_12934,N_14621);
nor U18636 (N_18636,N_12009,N_15036);
xnor U18637 (N_18637,N_15857,N_13277);
nand U18638 (N_18638,N_15040,N_15699);
nand U18639 (N_18639,N_13365,N_12313);
or U18640 (N_18640,N_15742,N_12259);
xnor U18641 (N_18641,N_15749,N_13438);
xor U18642 (N_18642,N_12154,N_12511);
and U18643 (N_18643,N_14748,N_12297);
nand U18644 (N_18644,N_13692,N_14314);
or U18645 (N_18645,N_15576,N_15614);
nand U18646 (N_18646,N_15174,N_15619);
and U18647 (N_18647,N_12771,N_15484);
xor U18648 (N_18648,N_15676,N_13931);
and U18649 (N_18649,N_14797,N_15497);
nor U18650 (N_18650,N_12919,N_15081);
xor U18651 (N_18651,N_13973,N_13310);
nor U18652 (N_18652,N_15911,N_14236);
or U18653 (N_18653,N_15804,N_13474);
nor U18654 (N_18654,N_12953,N_12056);
or U18655 (N_18655,N_12771,N_13068);
nor U18656 (N_18656,N_14716,N_13083);
xor U18657 (N_18657,N_12214,N_13567);
nand U18658 (N_18658,N_15132,N_12673);
or U18659 (N_18659,N_13803,N_13572);
or U18660 (N_18660,N_15171,N_15569);
and U18661 (N_18661,N_15544,N_15781);
nor U18662 (N_18662,N_13046,N_12339);
or U18663 (N_18663,N_14732,N_14533);
nor U18664 (N_18664,N_13457,N_14053);
nand U18665 (N_18665,N_15411,N_12813);
and U18666 (N_18666,N_14744,N_15117);
xnor U18667 (N_18667,N_15364,N_13099);
and U18668 (N_18668,N_14724,N_14466);
xor U18669 (N_18669,N_13607,N_12208);
xor U18670 (N_18670,N_15586,N_13967);
xnor U18671 (N_18671,N_13664,N_15478);
nand U18672 (N_18672,N_15874,N_13017);
nand U18673 (N_18673,N_12963,N_13730);
or U18674 (N_18674,N_12945,N_12001);
nor U18675 (N_18675,N_14597,N_15503);
nand U18676 (N_18676,N_15780,N_13990);
nor U18677 (N_18677,N_14157,N_14633);
or U18678 (N_18678,N_14338,N_15578);
xnor U18679 (N_18679,N_15215,N_15881);
nand U18680 (N_18680,N_12169,N_14032);
and U18681 (N_18681,N_12864,N_13308);
and U18682 (N_18682,N_12332,N_15262);
nand U18683 (N_18683,N_13524,N_15687);
or U18684 (N_18684,N_14938,N_14905);
nand U18685 (N_18685,N_14095,N_14854);
and U18686 (N_18686,N_12190,N_13603);
nand U18687 (N_18687,N_13018,N_12069);
and U18688 (N_18688,N_12409,N_13961);
nand U18689 (N_18689,N_13713,N_14228);
nor U18690 (N_18690,N_14288,N_12229);
nor U18691 (N_18691,N_14669,N_15895);
or U18692 (N_18692,N_15003,N_15927);
nand U18693 (N_18693,N_12280,N_12083);
nor U18694 (N_18694,N_15378,N_14525);
nand U18695 (N_18695,N_12122,N_15628);
and U18696 (N_18696,N_12064,N_14089);
or U18697 (N_18697,N_13515,N_12279);
or U18698 (N_18698,N_13459,N_13210);
xor U18699 (N_18699,N_13893,N_14197);
nor U18700 (N_18700,N_13327,N_14107);
nor U18701 (N_18701,N_15419,N_15514);
and U18702 (N_18702,N_13806,N_12970);
or U18703 (N_18703,N_14108,N_15177);
xnor U18704 (N_18704,N_15731,N_15982);
nand U18705 (N_18705,N_13708,N_12941);
nor U18706 (N_18706,N_12760,N_15924);
xnor U18707 (N_18707,N_15475,N_15441);
nand U18708 (N_18708,N_14339,N_14732);
or U18709 (N_18709,N_14278,N_13123);
nor U18710 (N_18710,N_14953,N_15008);
nand U18711 (N_18711,N_14329,N_14548);
and U18712 (N_18712,N_15196,N_12406);
nor U18713 (N_18713,N_15983,N_14332);
or U18714 (N_18714,N_15126,N_15513);
nand U18715 (N_18715,N_12077,N_12674);
or U18716 (N_18716,N_13998,N_14165);
xnor U18717 (N_18717,N_12868,N_13469);
nor U18718 (N_18718,N_12397,N_12955);
xnor U18719 (N_18719,N_15585,N_15743);
nand U18720 (N_18720,N_15954,N_13373);
nor U18721 (N_18721,N_13598,N_12601);
and U18722 (N_18722,N_12640,N_15731);
xnor U18723 (N_18723,N_13729,N_12316);
xor U18724 (N_18724,N_14107,N_13369);
or U18725 (N_18725,N_12536,N_12230);
nand U18726 (N_18726,N_13329,N_12729);
or U18727 (N_18727,N_14260,N_13960);
xor U18728 (N_18728,N_15822,N_13746);
and U18729 (N_18729,N_13291,N_13731);
nand U18730 (N_18730,N_14636,N_13290);
nand U18731 (N_18731,N_14531,N_12579);
and U18732 (N_18732,N_13409,N_14970);
and U18733 (N_18733,N_14384,N_12482);
nor U18734 (N_18734,N_13343,N_15186);
or U18735 (N_18735,N_15581,N_13005);
or U18736 (N_18736,N_15434,N_15531);
or U18737 (N_18737,N_15119,N_14132);
nor U18738 (N_18738,N_12315,N_14365);
nand U18739 (N_18739,N_14003,N_14191);
nand U18740 (N_18740,N_12869,N_13362);
or U18741 (N_18741,N_12026,N_12552);
or U18742 (N_18742,N_12363,N_14033);
nor U18743 (N_18743,N_12397,N_12020);
or U18744 (N_18744,N_14832,N_13717);
or U18745 (N_18745,N_12031,N_13849);
or U18746 (N_18746,N_13729,N_12645);
nor U18747 (N_18747,N_15677,N_13216);
or U18748 (N_18748,N_15814,N_13558);
nand U18749 (N_18749,N_12453,N_12741);
or U18750 (N_18750,N_12017,N_14282);
and U18751 (N_18751,N_12714,N_13204);
nand U18752 (N_18752,N_14529,N_15352);
and U18753 (N_18753,N_15292,N_12163);
and U18754 (N_18754,N_12613,N_12045);
or U18755 (N_18755,N_12601,N_13979);
or U18756 (N_18756,N_15812,N_12725);
and U18757 (N_18757,N_14938,N_13497);
xor U18758 (N_18758,N_15610,N_15410);
nand U18759 (N_18759,N_13337,N_12041);
nand U18760 (N_18760,N_12585,N_13633);
and U18761 (N_18761,N_14664,N_15779);
nand U18762 (N_18762,N_15250,N_12665);
and U18763 (N_18763,N_14366,N_12163);
or U18764 (N_18764,N_15899,N_15724);
nand U18765 (N_18765,N_13947,N_14234);
nor U18766 (N_18766,N_14114,N_12441);
nand U18767 (N_18767,N_12006,N_12933);
nand U18768 (N_18768,N_15260,N_13775);
and U18769 (N_18769,N_14756,N_14187);
xor U18770 (N_18770,N_14685,N_15431);
nand U18771 (N_18771,N_14731,N_15500);
xor U18772 (N_18772,N_12107,N_13453);
or U18773 (N_18773,N_14082,N_12447);
and U18774 (N_18774,N_15910,N_12553);
or U18775 (N_18775,N_15795,N_15497);
nand U18776 (N_18776,N_13478,N_14361);
and U18777 (N_18777,N_12497,N_13146);
xor U18778 (N_18778,N_12376,N_13602);
nand U18779 (N_18779,N_13797,N_15701);
and U18780 (N_18780,N_14903,N_14572);
nor U18781 (N_18781,N_12865,N_12342);
nand U18782 (N_18782,N_13201,N_15781);
xor U18783 (N_18783,N_14543,N_15112);
and U18784 (N_18784,N_15034,N_12228);
xor U18785 (N_18785,N_14662,N_13030);
and U18786 (N_18786,N_13828,N_12741);
xnor U18787 (N_18787,N_12606,N_15760);
nand U18788 (N_18788,N_13664,N_14080);
xnor U18789 (N_18789,N_14834,N_12043);
or U18790 (N_18790,N_12801,N_13345);
nor U18791 (N_18791,N_15952,N_13183);
nand U18792 (N_18792,N_14381,N_12060);
nand U18793 (N_18793,N_13688,N_13754);
nor U18794 (N_18794,N_14927,N_12495);
and U18795 (N_18795,N_15833,N_15542);
and U18796 (N_18796,N_12910,N_12199);
xnor U18797 (N_18797,N_14349,N_12210);
nor U18798 (N_18798,N_14346,N_13915);
and U18799 (N_18799,N_12418,N_13511);
xnor U18800 (N_18800,N_12648,N_14730);
and U18801 (N_18801,N_15212,N_15642);
xor U18802 (N_18802,N_14017,N_14334);
xnor U18803 (N_18803,N_12984,N_12199);
nor U18804 (N_18804,N_13033,N_15608);
and U18805 (N_18805,N_15051,N_13767);
nand U18806 (N_18806,N_12814,N_15789);
nand U18807 (N_18807,N_13533,N_13419);
or U18808 (N_18808,N_15031,N_15134);
nand U18809 (N_18809,N_15814,N_13553);
and U18810 (N_18810,N_13516,N_14333);
nor U18811 (N_18811,N_14049,N_12467);
xor U18812 (N_18812,N_13393,N_14978);
nand U18813 (N_18813,N_12703,N_15560);
or U18814 (N_18814,N_13961,N_14590);
nand U18815 (N_18815,N_15428,N_15400);
nand U18816 (N_18816,N_15712,N_12043);
and U18817 (N_18817,N_13762,N_15177);
xnor U18818 (N_18818,N_12875,N_12313);
nor U18819 (N_18819,N_12697,N_12776);
and U18820 (N_18820,N_13278,N_14553);
nor U18821 (N_18821,N_13830,N_13826);
and U18822 (N_18822,N_15519,N_14207);
and U18823 (N_18823,N_13898,N_12306);
or U18824 (N_18824,N_14107,N_15366);
and U18825 (N_18825,N_14295,N_14771);
nor U18826 (N_18826,N_13736,N_13836);
nand U18827 (N_18827,N_15042,N_13496);
and U18828 (N_18828,N_12384,N_15935);
nand U18829 (N_18829,N_14577,N_15726);
nor U18830 (N_18830,N_15500,N_15572);
and U18831 (N_18831,N_15609,N_14914);
or U18832 (N_18832,N_15154,N_14933);
nor U18833 (N_18833,N_14721,N_15330);
nor U18834 (N_18834,N_14305,N_12802);
nor U18835 (N_18835,N_12171,N_14059);
and U18836 (N_18836,N_12800,N_13327);
or U18837 (N_18837,N_13210,N_13453);
or U18838 (N_18838,N_14382,N_12038);
or U18839 (N_18839,N_12255,N_15466);
nand U18840 (N_18840,N_14802,N_15561);
nand U18841 (N_18841,N_13577,N_15389);
or U18842 (N_18842,N_14204,N_15283);
or U18843 (N_18843,N_15092,N_13481);
and U18844 (N_18844,N_12818,N_15727);
and U18845 (N_18845,N_13834,N_15481);
or U18846 (N_18846,N_15879,N_15643);
or U18847 (N_18847,N_12309,N_14077);
nand U18848 (N_18848,N_14793,N_14859);
or U18849 (N_18849,N_13870,N_15286);
or U18850 (N_18850,N_12469,N_14151);
and U18851 (N_18851,N_13224,N_13030);
nand U18852 (N_18852,N_13782,N_15376);
and U18853 (N_18853,N_12555,N_14507);
nor U18854 (N_18854,N_15975,N_12328);
xnor U18855 (N_18855,N_15161,N_15353);
and U18856 (N_18856,N_15134,N_12993);
nor U18857 (N_18857,N_15336,N_12610);
and U18858 (N_18858,N_14271,N_13644);
and U18859 (N_18859,N_15624,N_14895);
xor U18860 (N_18860,N_14276,N_15774);
nand U18861 (N_18861,N_15575,N_14130);
nand U18862 (N_18862,N_15121,N_14355);
nor U18863 (N_18863,N_13491,N_13038);
or U18864 (N_18864,N_14349,N_14439);
nor U18865 (N_18865,N_15370,N_13031);
or U18866 (N_18866,N_13119,N_13169);
nand U18867 (N_18867,N_14829,N_13410);
nand U18868 (N_18868,N_13151,N_14180);
nor U18869 (N_18869,N_12248,N_12238);
or U18870 (N_18870,N_15194,N_15809);
and U18871 (N_18871,N_15475,N_13142);
nand U18872 (N_18872,N_15074,N_13988);
and U18873 (N_18873,N_15905,N_12583);
nor U18874 (N_18874,N_13487,N_13498);
nand U18875 (N_18875,N_12090,N_15327);
and U18876 (N_18876,N_13113,N_12977);
and U18877 (N_18877,N_12618,N_13840);
or U18878 (N_18878,N_12402,N_14368);
nand U18879 (N_18879,N_14612,N_12613);
nand U18880 (N_18880,N_12715,N_15259);
nand U18881 (N_18881,N_14759,N_14974);
nand U18882 (N_18882,N_12956,N_15822);
nor U18883 (N_18883,N_14956,N_15828);
and U18884 (N_18884,N_15772,N_14811);
or U18885 (N_18885,N_14034,N_12191);
and U18886 (N_18886,N_15829,N_14906);
nand U18887 (N_18887,N_12416,N_12966);
or U18888 (N_18888,N_12120,N_15072);
and U18889 (N_18889,N_13825,N_13226);
nand U18890 (N_18890,N_12461,N_14046);
nor U18891 (N_18891,N_15819,N_15135);
and U18892 (N_18892,N_12183,N_12331);
xor U18893 (N_18893,N_12239,N_12568);
xnor U18894 (N_18894,N_15782,N_14125);
or U18895 (N_18895,N_15331,N_13239);
or U18896 (N_18896,N_13864,N_15162);
nor U18897 (N_18897,N_15455,N_15195);
nand U18898 (N_18898,N_15804,N_13241);
nor U18899 (N_18899,N_12025,N_14638);
nor U18900 (N_18900,N_15416,N_15953);
and U18901 (N_18901,N_12923,N_13163);
nor U18902 (N_18902,N_14267,N_15144);
nand U18903 (N_18903,N_14364,N_14968);
nand U18904 (N_18904,N_14373,N_14642);
or U18905 (N_18905,N_15022,N_15914);
nand U18906 (N_18906,N_15236,N_12898);
or U18907 (N_18907,N_14064,N_14096);
and U18908 (N_18908,N_12608,N_12061);
nand U18909 (N_18909,N_14607,N_14891);
nand U18910 (N_18910,N_13441,N_15619);
nor U18911 (N_18911,N_12566,N_15596);
nor U18912 (N_18912,N_15038,N_12148);
nand U18913 (N_18913,N_12786,N_14806);
nand U18914 (N_18914,N_12685,N_12765);
nand U18915 (N_18915,N_13925,N_14017);
nor U18916 (N_18916,N_15624,N_12578);
nor U18917 (N_18917,N_15214,N_14097);
xor U18918 (N_18918,N_14019,N_13726);
and U18919 (N_18919,N_15470,N_15090);
and U18920 (N_18920,N_13807,N_14833);
xor U18921 (N_18921,N_14941,N_12934);
nor U18922 (N_18922,N_12228,N_12521);
nor U18923 (N_18923,N_14981,N_13803);
nand U18924 (N_18924,N_13622,N_14845);
or U18925 (N_18925,N_14814,N_15456);
or U18926 (N_18926,N_13951,N_15142);
and U18927 (N_18927,N_12284,N_15796);
nand U18928 (N_18928,N_12183,N_13128);
nor U18929 (N_18929,N_12233,N_15767);
nor U18930 (N_18930,N_15498,N_12319);
nor U18931 (N_18931,N_12668,N_15936);
and U18932 (N_18932,N_14452,N_13193);
or U18933 (N_18933,N_15460,N_15883);
nor U18934 (N_18934,N_13800,N_15595);
xor U18935 (N_18935,N_12754,N_12300);
or U18936 (N_18936,N_14534,N_15256);
xor U18937 (N_18937,N_15400,N_13599);
and U18938 (N_18938,N_14193,N_15761);
nor U18939 (N_18939,N_15363,N_13534);
nand U18940 (N_18940,N_15943,N_15139);
or U18941 (N_18941,N_13383,N_12358);
nor U18942 (N_18942,N_14929,N_15450);
xor U18943 (N_18943,N_15294,N_15028);
or U18944 (N_18944,N_15741,N_14174);
nand U18945 (N_18945,N_14473,N_13119);
xor U18946 (N_18946,N_15385,N_14714);
and U18947 (N_18947,N_14583,N_13457);
nand U18948 (N_18948,N_15829,N_15029);
and U18949 (N_18949,N_14211,N_15835);
and U18950 (N_18950,N_13002,N_12766);
and U18951 (N_18951,N_13302,N_13033);
nand U18952 (N_18952,N_12290,N_13417);
nor U18953 (N_18953,N_12426,N_15668);
and U18954 (N_18954,N_12474,N_15460);
nand U18955 (N_18955,N_12803,N_14370);
nor U18956 (N_18956,N_12432,N_15656);
nand U18957 (N_18957,N_13639,N_13830);
nor U18958 (N_18958,N_14177,N_13833);
or U18959 (N_18959,N_14770,N_12332);
nand U18960 (N_18960,N_15125,N_14464);
nor U18961 (N_18961,N_15542,N_15453);
and U18962 (N_18962,N_15590,N_12558);
nor U18963 (N_18963,N_15847,N_13164);
nand U18964 (N_18964,N_12826,N_13920);
and U18965 (N_18965,N_13796,N_14739);
and U18966 (N_18966,N_13297,N_15807);
or U18967 (N_18967,N_14007,N_15040);
nor U18968 (N_18968,N_13981,N_12803);
and U18969 (N_18969,N_14761,N_15962);
or U18970 (N_18970,N_12986,N_12089);
and U18971 (N_18971,N_14984,N_12184);
xnor U18972 (N_18972,N_13227,N_14995);
and U18973 (N_18973,N_15384,N_14819);
xnor U18974 (N_18974,N_13197,N_14833);
and U18975 (N_18975,N_14965,N_13921);
and U18976 (N_18976,N_14184,N_15816);
or U18977 (N_18977,N_15962,N_13400);
nor U18978 (N_18978,N_14790,N_12259);
and U18979 (N_18979,N_12644,N_14339);
nand U18980 (N_18980,N_14411,N_12989);
or U18981 (N_18981,N_14711,N_14509);
and U18982 (N_18982,N_15729,N_14171);
and U18983 (N_18983,N_12742,N_15940);
and U18984 (N_18984,N_12367,N_12200);
and U18985 (N_18985,N_13059,N_13790);
and U18986 (N_18986,N_15837,N_13355);
nand U18987 (N_18987,N_14680,N_14290);
nand U18988 (N_18988,N_12641,N_12161);
nor U18989 (N_18989,N_13427,N_12893);
nand U18990 (N_18990,N_13072,N_13090);
nand U18991 (N_18991,N_13535,N_12739);
nand U18992 (N_18992,N_15129,N_13669);
and U18993 (N_18993,N_13254,N_14846);
or U18994 (N_18994,N_14395,N_15268);
and U18995 (N_18995,N_14784,N_13395);
nand U18996 (N_18996,N_14315,N_12537);
nand U18997 (N_18997,N_13563,N_14611);
nor U18998 (N_18998,N_14505,N_14929);
or U18999 (N_18999,N_14942,N_13404);
and U19000 (N_19000,N_13791,N_14258);
nand U19001 (N_19001,N_12109,N_13839);
xnor U19002 (N_19002,N_12941,N_13509);
nand U19003 (N_19003,N_15616,N_15672);
and U19004 (N_19004,N_15539,N_15410);
nor U19005 (N_19005,N_12500,N_12059);
nand U19006 (N_19006,N_12576,N_15068);
nor U19007 (N_19007,N_15980,N_14496);
nor U19008 (N_19008,N_14519,N_15512);
xor U19009 (N_19009,N_15367,N_14033);
nor U19010 (N_19010,N_14424,N_14752);
nor U19011 (N_19011,N_15038,N_13807);
xnor U19012 (N_19012,N_13861,N_14946);
nor U19013 (N_19013,N_15303,N_14049);
xor U19014 (N_19014,N_12758,N_12355);
xor U19015 (N_19015,N_12820,N_14326);
nand U19016 (N_19016,N_12324,N_13497);
xor U19017 (N_19017,N_13597,N_13748);
nand U19018 (N_19018,N_14391,N_12875);
or U19019 (N_19019,N_14980,N_12319);
or U19020 (N_19020,N_12730,N_12773);
nor U19021 (N_19021,N_13926,N_14133);
nand U19022 (N_19022,N_15858,N_12771);
or U19023 (N_19023,N_15835,N_15862);
xor U19024 (N_19024,N_14196,N_15361);
and U19025 (N_19025,N_14802,N_12940);
or U19026 (N_19026,N_12075,N_14862);
nand U19027 (N_19027,N_12884,N_15000);
nand U19028 (N_19028,N_14356,N_13573);
and U19029 (N_19029,N_14244,N_12751);
nand U19030 (N_19030,N_15782,N_12374);
and U19031 (N_19031,N_14279,N_14153);
nand U19032 (N_19032,N_15036,N_15567);
nor U19033 (N_19033,N_15686,N_14388);
nand U19034 (N_19034,N_14043,N_14385);
or U19035 (N_19035,N_13817,N_13243);
nand U19036 (N_19036,N_12306,N_15726);
nand U19037 (N_19037,N_15545,N_13902);
nor U19038 (N_19038,N_15560,N_13908);
nor U19039 (N_19039,N_12515,N_14016);
nand U19040 (N_19040,N_14994,N_12036);
and U19041 (N_19041,N_12334,N_12115);
or U19042 (N_19042,N_15541,N_15148);
or U19043 (N_19043,N_13728,N_12637);
or U19044 (N_19044,N_13867,N_14022);
and U19045 (N_19045,N_12884,N_15595);
xnor U19046 (N_19046,N_13305,N_12871);
and U19047 (N_19047,N_13509,N_15901);
or U19048 (N_19048,N_13210,N_12307);
or U19049 (N_19049,N_13228,N_13815);
and U19050 (N_19050,N_12715,N_15937);
nand U19051 (N_19051,N_15622,N_12563);
nor U19052 (N_19052,N_13815,N_12268);
nor U19053 (N_19053,N_14599,N_14309);
nor U19054 (N_19054,N_12565,N_12833);
xor U19055 (N_19055,N_15018,N_15291);
xnor U19056 (N_19056,N_15945,N_14298);
nor U19057 (N_19057,N_13363,N_12627);
and U19058 (N_19058,N_13075,N_13855);
and U19059 (N_19059,N_14771,N_13328);
xor U19060 (N_19060,N_13571,N_15306);
and U19061 (N_19061,N_14809,N_13729);
xnor U19062 (N_19062,N_15728,N_15409);
and U19063 (N_19063,N_12242,N_14449);
or U19064 (N_19064,N_14214,N_13744);
or U19065 (N_19065,N_14972,N_12678);
or U19066 (N_19066,N_14659,N_14689);
nor U19067 (N_19067,N_15854,N_12997);
and U19068 (N_19068,N_15481,N_13149);
nand U19069 (N_19069,N_13558,N_15227);
and U19070 (N_19070,N_14850,N_14128);
and U19071 (N_19071,N_13661,N_15291);
nand U19072 (N_19072,N_14615,N_12416);
nor U19073 (N_19073,N_12884,N_13304);
or U19074 (N_19074,N_12633,N_15563);
nor U19075 (N_19075,N_14328,N_14071);
nand U19076 (N_19076,N_13894,N_13411);
or U19077 (N_19077,N_15527,N_12018);
or U19078 (N_19078,N_15513,N_13978);
nor U19079 (N_19079,N_14561,N_12529);
nor U19080 (N_19080,N_12846,N_13671);
or U19081 (N_19081,N_12698,N_15357);
nand U19082 (N_19082,N_12549,N_12543);
or U19083 (N_19083,N_14330,N_13325);
nand U19084 (N_19084,N_13139,N_13644);
or U19085 (N_19085,N_14797,N_13497);
and U19086 (N_19086,N_12282,N_12928);
or U19087 (N_19087,N_12209,N_14377);
and U19088 (N_19088,N_13187,N_15862);
nor U19089 (N_19089,N_15969,N_13444);
nor U19090 (N_19090,N_13270,N_15153);
nand U19091 (N_19091,N_14591,N_12183);
and U19092 (N_19092,N_15954,N_15398);
nand U19093 (N_19093,N_14438,N_15218);
or U19094 (N_19094,N_15463,N_12532);
nand U19095 (N_19095,N_12052,N_14901);
nand U19096 (N_19096,N_14440,N_13144);
or U19097 (N_19097,N_15519,N_12511);
nor U19098 (N_19098,N_15627,N_14975);
and U19099 (N_19099,N_13499,N_14474);
nor U19100 (N_19100,N_15405,N_13544);
nand U19101 (N_19101,N_14693,N_13614);
and U19102 (N_19102,N_12960,N_14116);
xor U19103 (N_19103,N_13993,N_13398);
nand U19104 (N_19104,N_15668,N_14356);
or U19105 (N_19105,N_14884,N_13289);
or U19106 (N_19106,N_15200,N_15383);
nor U19107 (N_19107,N_14058,N_15753);
and U19108 (N_19108,N_12212,N_12068);
or U19109 (N_19109,N_15031,N_13810);
and U19110 (N_19110,N_14804,N_15627);
xor U19111 (N_19111,N_14755,N_15944);
nand U19112 (N_19112,N_15995,N_12483);
or U19113 (N_19113,N_14269,N_13911);
nand U19114 (N_19114,N_12071,N_13434);
or U19115 (N_19115,N_14947,N_15631);
or U19116 (N_19116,N_12679,N_12397);
or U19117 (N_19117,N_13908,N_13869);
nor U19118 (N_19118,N_14212,N_14473);
and U19119 (N_19119,N_15401,N_12634);
nor U19120 (N_19120,N_15834,N_14172);
nor U19121 (N_19121,N_13109,N_15100);
nand U19122 (N_19122,N_13029,N_15393);
or U19123 (N_19123,N_13145,N_14668);
and U19124 (N_19124,N_15599,N_13218);
nand U19125 (N_19125,N_14708,N_14212);
nor U19126 (N_19126,N_13659,N_14811);
or U19127 (N_19127,N_15161,N_15943);
or U19128 (N_19128,N_15012,N_14554);
or U19129 (N_19129,N_15506,N_12788);
xnor U19130 (N_19130,N_12811,N_15669);
nand U19131 (N_19131,N_12856,N_12117);
nor U19132 (N_19132,N_15948,N_14448);
nand U19133 (N_19133,N_15491,N_15703);
nand U19134 (N_19134,N_15789,N_12232);
nand U19135 (N_19135,N_13861,N_13773);
and U19136 (N_19136,N_13380,N_15634);
nor U19137 (N_19137,N_13523,N_15531);
or U19138 (N_19138,N_12696,N_12380);
nand U19139 (N_19139,N_13640,N_14372);
and U19140 (N_19140,N_12950,N_13552);
xnor U19141 (N_19141,N_12606,N_14632);
or U19142 (N_19142,N_13811,N_13061);
nand U19143 (N_19143,N_13395,N_13896);
nand U19144 (N_19144,N_15452,N_12874);
nor U19145 (N_19145,N_12947,N_12156);
nand U19146 (N_19146,N_15686,N_14124);
and U19147 (N_19147,N_12670,N_15818);
nor U19148 (N_19148,N_15889,N_12144);
or U19149 (N_19149,N_13028,N_14205);
nand U19150 (N_19150,N_13941,N_13562);
and U19151 (N_19151,N_13290,N_15155);
xor U19152 (N_19152,N_14163,N_12564);
and U19153 (N_19153,N_12853,N_15253);
and U19154 (N_19154,N_14446,N_15518);
or U19155 (N_19155,N_15864,N_13269);
xnor U19156 (N_19156,N_12616,N_15348);
xor U19157 (N_19157,N_12135,N_13115);
nor U19158 (N_19158,N_13562,N_14591);
nand U19159 (N_19159,N_12993,N_15911);
nand U19160 (N_19160,N_12883,N_12985);
nor U19161 (N_19161,N_14755,N_13675);
or U19162 (N_19162,N_14911,N_12142);
and U19163 (N_19163,N_14917,N_13719);
or U19164 (N_19164,N_15051,N_15749);
and U19165 (N_19165,N_12181,N_15853);
nand U19166 (N_19166,N_12394,N_15919);
nand U19167 (N_19167,N_12372,N_15820);
nor U19168 (N_19168,N_14621,N_15341);
nor U19169 (N_19169,N_12989,N_13874);
nand U19170 (N_19170,N_15440,N_14746);
nor U19171 (N_19171,N_12158,N_15735);
nor U19172 (N_19172,N_14738,N_15297);
nand U19173 (N_19173,N_13080,N_12389);
nor U19174 (N_19174,N_13245,N_13465);
nor U19175 (N_19175,N_15627,N_13140);
or U19176 (N_19176,N_12493,N_15683);
xor U19177 (N_19177,N_12699,N_15613);
nor U19178 (N_19178,N_12245,N_12527);
xnor U19179 (N_19179,N_12499,N_14006);
or U19180 (N_19180,N_15511,N_12604);
and U19181 (N_19181,N_14916,N_13882);
or U19182 (N_19182,N_13807,N_12418);
and U19183 (N_19183,N_12523,N_12111);
nor U19184 (N_19184,N_12010,N_13282);
and U19185 (N_19185,N_15400,N_13911);
nor U19186 (N_19186,N_12517,N_13347);
xor U19187 (N_19187,N_12147,N_14157);
nor U19188 (N_19188,N_14555,N_14334);
nand U19189 (N_19189,N_14069,N_15131);
nand U19190 (N_19190,N_14804,N_12350);
or U19191 (N_19191,N_13354,N_14890);
nor U19192 (N_19192,N_13701,N_12694);
nand U19193 (N_19193,N_14662,N_13998);
nor U19194 (N_19194,N_14272,N_13623);
or U19195 (N_19195,N_13101,N_14813);
or U19196 (N_19196,N_15335,N_12538);
nand U19197 (N_19197,N_14316,N_14023);
or U19198 (N_19198,N_13222,N_13010);
xor U19199 (N_19199,N_13717,N_14608);
nor U19200 (N_19200,N_12150,N_15535);
and U19201 (N_19201,N_13681,N_12865);
nor U19202 (N_19202,N_15309,N_14648);
xnor U19203 (N_19203,N_13125,N_14622);
nand U19204 (N_19204,N_15455,N_15345);
and U19205 (N_19205,N_14883,N_14598);
or U19206 (N_19206,N_14755,N_13860);
nand U19207 (N_19207,N_12690,N_12399);
nor U19208 (N_19208,N_14560,N_13400);
nor U19209 (N_19209,N_13156,N_14940);
nand U19210 (N_19210,N_12269,N_12172);
nor U19211 (N_19211,N_12297,N_12226);
nor U19212 (N_19212,N_12197,N_15302);
and U19213 (N_19213,N_12126,N_12165);
nor U19214 (N_19214,N_14054,N_12542);
nor U19215 (N_19215,N_14413,N_15859);
or U19216 (N_19216,N_14697,N_15140);
and U19217 (N_19217,N_12030,N_15998);
xor U19218 (N_19218,N_13842,N_14605);
and U19219 (N_19219,N_13427,N_14786);
nor U19220 (N_19220,N_14507,N_14970);
and U19221 (N_19221,N_14148,N_15134);
xor U19222 (N_19222,N_12541,N_12495);
nand U19223 (N_19223,N_15157,N_12286);
nand U19224 (N_19224,N_12606,N_13944);
nor U19225 (N_19225,N_14650,N_15172);
or U19226 (N_19226,N_13844,N_13808);
or U19227 (N_19227,N_13358,N_15087);
xor U19228 (N_19228,N_15720,N_15753);
xor U19229 (N_19229,N_13397,N_13415);
nor U19230 (N_19230,N_15230,N_14650);
nor U19231 (N_19231,N_15161,N_15246);
nand U19232 (N_19232,N_15768,N_13833);
and U19233 (N_19233,N_12810,N_14266);
or U19234 (N_19234,N_15582,N_15306);
nor U19235 (N_19235,N_13564,N_13881);
or U19236 (N_19236,N_15816,N_14484);
nor U19237 (N_19237,N_15443,N_15493);
nor U19238 (N_19238,N_13652,N_15691);
and U19239 (N_19239,N_15993,N_12602);
or U19240 (N_19240,N_14577,N_12041);
nand U19241 (N_19241,N_15942,N_12477);
or U19242 (N_19242,N_12683,N_14879);
and U19243 (N_19243,N_13981,N_12171);
and U19244 (N_19244,N_12387,N_13265);
nand U19245 (N_19245,N_13802,N_13707);
nor U19246 (N_19246,N_15555,N_13631);
and U19247 (N_19247,N_15599,N_13571);
and U19248 (N_19248,N_15084,N_13609);
and U19249 (N_19249,N_14418,N_13747);
nor U19250 (N_19250,N_15548,N_13524);
or U19251 (N_19251,N_14809,N_13644);
and U19252 (N_19252,N_13881,N_12079);
nand U19253 (N_19253,N_14302,N_15379);
or U19254 (N_19254,N_15790,N_14040);
nand U19255 (N_19255,N_12706,N_13686);
or U19256 (N_19256,N_15380,N_15728);
nand U19257 (N_19257,N_12116,N_15960);
nor U19258 (N_19258,N_13488,N_12495);
nor U19259 (N_19259,N_14315,N_14782);
or U19260 (N_19260,N_12451,N_12426);
nand U19261 (N_19261,N_15116,N_13784);
nor U19262 (N_19262,N_15101,N_15035);
xor U19263 (N_19263,N_14631,N_13194);
xor U19264 (N_19264,N_13198,N_14310);
nor U19265 (N_19265,N_15985,N_12449);
or U19266 (N_19266,N_12773,N_14729);
or U19267 (N_19267,N_14007,N_15279);
and U19268 (N_19268,N_13800,N_13791);
nand U19269 (N_19269,N_14750,N_14031);
nand U19270 (N_19270,N_15058,N_12523);
and U19271 (N_19271,N_15776,N_13254);
xnor U19272 (N_19272,N_15599,N_14536);
or U19273 (N_19273,N_14530,N_12228);
nand U19274 (N_19274,N_12226,N_15066);
nand U19275 (N_19275,N_13260,N_13558);
and U19276 (N_19276,N_15116,N_15343);
xor U19277 (N_19277,N_12108,N_15764);
nor U19278 (N_19278,N_12372,N_13593);
nand U19279 (N_19279,N_13690,N_12114);
nor U19280 (N_19280,N_12403,N_12271);
nand U19281 (N_19281,N_14192,N_12689);
nand U19282 (N_19282,N_14116,N_13899);
nor U19283 (N_19283,N_12065,N_14293);
xor U19284 (N_19284,N_14733,N_12830);
xor U19285 (N_19285,N_14804,N_13635);
and U19286 (N_19286,N_15223,N_13935);
xnor U19287 (N_19287,N_15183,N_14599);
and U19288 (N_19288,N_12021,N_14512);
and U19289 (N_19289,N_14916,N_15881);
nand U19290 (N_19290,N_12410,N_12424);
and U19291 (N_19291,N_13694,N_13151);
and U19292 (N_19292,N_13130,N_15518);
nand U19293 (N_19293,N_15420,N_15209);
or U19294 (N_19294,N_12350,N_15446);
nor U19295 (N_19295,N_13562,N_12213);
and U19296 (N_19296,N_12629,N_12144);
or U19297 (N_19297,N_12359,N_12055);
nor U19298 (N_19298,N_13124,N_13258);
or U19299 (N_19299,N_15988,N_14194);
nor U19300 (N_19300,N_12767,N_12819);
and U19301 (N_19301,N_13038,N_13159);
nor U19302 (N_19302,N_13979,N_15112);
nand U19303 (N_19303,N_15489,N_13326);
nor U19304 (N_19304,N_12941,N_14895);
or U19305 (N_19305,N_15073,N_15263);
or U19306 (N_19306,N_14790,N_15911);
and U19307 (N_19307,N_14900,N_15536);
and U19308 (N_19308,N_15211,N_14429);
nor U19309 (N_19309,N_13990,N_14627);
nor U19310 (N_19310,N_13322,N_15369);
or U19311 (N_19311,N_13183,N_12755);
or U19312 (N_19312,N_15950,N_13664);
or U19313 (N_19313,N_13925,N_15852);
nand U19314 (N_19314,N_14339,N_15045);
or U19315 (N_19315,N_13483,N_15931);
nor U19316 (N_19316,N_14817,N_15432);
and U19317 (N_19317,N_13183,N_12318);
or U19318 (N_19318,N_12795,N_13235);
nor U19319 (N_19319,N_13199,N_14295);
or U19320 (N_19320,N_13215,N_13429);
or U19321 (N_19321,N_15775,N_15317);
or U19322 (N_19322,N_15386,N_12677);
or U19323 (N_19323,N_13763,N_14189);
or U19324 (N_19324,N_12537,N_12070);
and U19325 (N_19325,N_12323,N_14731);
or U19326 (N_19326,N_15877,N_13833);
nand U19327 (N_19327,N_14231,N_12829);
nor U19328 (N_19328,N_12108,N_15536);
and U19329 (N_19329,N_15015,N_12942);
and U19330 (N_19330,N_15491,N_13684);
and U19331 (N_19331,N_15273,N_13094);
nand U19332 (N_19332,N_13709,N_12509);
and U19333 (N_19333,N_15744,N_12608);
nor U19334 (N_19334,N_13341,N_14648);
and U19335 (N_19335,N_14009,N_13485);
xor U19336 (N_19336,N_15590,N_15093);
xor U19337 (N_19337,N_13399,N_12841);
nor U19338 (N_19338,N_13303,N_12632);
nand U19339 (N_19339,N_12370,N_12348);
and U19340 (N_19340,N_13981,N_12149);
xor U19341 (N_19341,N_15878,N_14412);
nor U19342 (N_19342,N_13109,N_12336);
xnor U19343 (N_19343,N_15217,N_15863);
nor U19344 (N_19344,N_12611,N_12892);
nand U19345 (N_19345,N_14885,N_15088);
or U19346 (N_19346,N_13064,N_15155);
or U19347 (N_19347,N_14052,N_14525);
and U19348 (N_19348,N_14562,N_14419);
or U19349 (N_19349,N_12950,N_13549);
xnor U19350 (N_19350,N_14171,N_12394);
and U19351 (N_19351,N_12041,N_12255);
and U19352 (N_19352,N_14537,N_13830);
and U19353 (N_19353,N_15930,N_13995);
nand U19354 (N_19354,N_15880,N_14124);
nor U19355 (N_19355,N_14029,N_15669);
xor U19356 (N_19356,N_14276,N_13477);
nand U19357 (N_19357,N_13676,N_14947);
or U19358 (N_19358,N_14721,N_14361);
and U19359 (N_19359,N_12752,N_12036);
nand U19360 (N_19360,N_14426,N_12647);
and U19361 (N_19361,N_15836,N_13424);
and U19362 (N_19362,N_13483,N_14605);
or U19363 (N_19363,N_13327,N_13556);
and U19364 (N_19364,N_13978,N_12172);
and U19365 (N_19365,N_14246,N_14113);
nand U19366 (N_19366,N_13880,N_14882);
nand U19367 (N_19367,N_13207,N_12772);
nor U19368 (N_19368,N_14755,N_12956);
nand U19369 (N_19369,N_15016,N_13956);
and U19370 (N_19370,N_13768,N_13968);
nand U19371 (N_19371,N_15683,N_15294);
nor U19372 (N_19372,N_12149,N_14247);
and U19373 (N_19373,N_13223,N_12258);
xor U19374 (N_19374,N_12524,N_12886);
nor U19375 (N_19375,N_15412,N_14962);
or U19376 (N_19376,N_14553,N_14321);
nand U19377 (N_19377,N_14627,N_15636);
nand U19378 (N_19378,N_12911,N_14609);
nor U19379 (N_19379,N_12554,N_12925);
nor U19380 (N_19380,N_15906,N_12359);
nor U19381 (N_19381,N_12479,N_12558);
nand U19382 (N_19382,N_13037,N_13822);
nor U19383 (N_19383,N_12357,N_15252);
nor U19384 (N_19384,N_13084,N_14704);
and U19385 (N_19385,N_13118,N_15217);
xnor U19386 (N_19386,N_15486,N_13894);
nand U19387 (N_19387,N_15580,N_12103);
nor U19388 (N_19388,N_15735,N_12252);
or U19389 (N_19389,N_13766,N_15692);
nand U19390 (N_19390,N_15287,N_15800);
nand U19391 (N_19391,N_15397,N_15844);
nand U19392 (N_19392,N_12434,N_13385);
nor U19393 (N_19393,N_15255,N_12681);
xnor U19394 (N_19394,N_12349,N_13323);
nor U19395 (N_19395,N_15146,N_15137);
nand U19396 (N_19396,N_14125,N_12776);
and U19397 (N_19397,N_13731,N_12413);
nor U19398 (N_19398,N_12058,N_12782);
or U19399 (N_19399,N_12036,N_13023);
xor U19400 (N_19400,N_14218,N_12691);
or U19401 (N_19401,N_14280,N_13486);
or U19402 (N_19402,N_13024,N_14258);
and U19403 (N_19403,N_12308,N_12173);
nor U19404 (N_19404,N_14287,N_14811);
and U19405 (N_19405,N_13610,N_15896);
and U19406 (N_19406,N_13983,N_14509);
and U19407 (N_19407,N_13299,N_12607);
nand U19408 (N_19408,N_15126,N_12432);
nor U19409 (N_19409,N_15023,N_15080);
nor U19410 (N_19410,N_12892,N_13628);
xor U19411 (N_19411,N_13065,N_14769);
and U19412 (N_19412,N_12891,N_12426);
or U19413 (N_19413,N_13192,N_15749);
or U19414 (N_19414,N_15872,N_12195);
nand U19415 (N_19415,N_15354,N_12344);
nand U19416 (N_19416,N_15276,N_12794);
and U19417 (N_19417,N_15809,N_14025);
nand U19418 (N_19418,N_13091,N_15627);
nand U19419 (N_19419,N_12413,N_15523);
nand U19420 (N_19420,N_12021,N_12305);
nor U19421 (N_19421,N_14631,N_12437);
nor U19422 (N_19422,N_15217,N_14009);
nand U19423 (N_19423,N_12992,N_12908);
nor U19424 (N_19424,N_13571,N_12354);
and U19425 (N_19425,N_12340,N_12539);
and U19426 (N_19426,N_13500,N_14404);
xor U19427 (N_19427,N_14719,N_12275);
nor U19428 (N_19428,N_12814,N_12216);
nor U19429 (N_19429,N_14282,N_13478);
and U19430 (N_19430,N_14847,N_13898);
nor U19431 (N_19431,N_14843,N_14799);
or U19432 (N_19432,N_12220,N_14263);
nand U19433 (N_19433,N_14382,N_15586);
nand U19434 (N_19434,N_15927,N_14202);
or U19435 (N_19435,N_12246,N_15597);
nand U19436 (N_19436,N_15507,N_13036);
or U19437 (N_19437,N_15259,N_14016);
or U19438 (N_19438,N_14538,N_14110);
nor U19439 (N_19439,N_13039,N_14487);
nor U19440 (N_19440,N_14291,N_13339);
and U19441 (N_19441,N_13328,N_15365);
nand U19442 (N_19442,N_13225,N_12341);
nand U19443 (N_19443,N_14321,N_13562);
and U19444 (N_19444,N_14077,N_13425);
nand U19445 (N_19445,N_13254,N_15832);
and U19446 (N_19446,N_12640,N_13468);
nor U19447 (N_19447,N_14892,N_12910);
or U19448 (N_19448,N_13481,N_15767);
xor U19449 (N_19449,N_15003,N_14067);
and U19450 (N_19450,N_12715,N_13313);
nand U19451 (N_19451,N_15603,N_14939);
nor U19452 (N_19452,N_15587,N_14765);
nand U19453 (N_19453,N_12777,N_14943);
and U19454 (N_19454,N_15757,N_15175);
nor U19455 (N_19455,N_14173,N_15405);
and U19456 (N_19456,N_14618,N_14400);
or U19457 (N_19457,N_12340,N_13543);
or U19458 (N_19458,N_14537,N_15438);
xor U19459 (N_19459,N_14542,N_12451);
xnor U19460 (N_19460,N_14899,N_14527);
nand U19461 (N_19461,N_15649,N_14040);
and U19462 (N_19462,N_12020,N_13144);
nor U19463 (N_19463,N_13310,N_12057);
or U19464 (N_19464,N_12418,N_12356);
nor U19465 (N_19465,N_15953,N_14493);
or U19466 (N_19466,N_13651,N_13553);
and U19467 (N_19467,N_12061,N_12172);
nand U19468 (N_19468,N_14426,N_14705);
nand U19469 (N_19469,N_12549,N_12873);
nand U19470 (N_19470,N_14708,N_13277);
nor U19471 (N_19471,N_14998,N_13022);
or U19472 (N_19472,N_15875,N_13394);
and U19473 (N_19473,N_14222,N_14937);
nand U19474 (N_19474,N_15849,N_12552);
xnor U19475 (N_19475,N_12847,N_13369);
or U19476 (N_19476,N_14253,N_13104);
nor U19477 (N_19477,N_14379,N_13003);
nand U19478 (N_19478,N_14119,N_15651);
or U19479 (N_19479,N_13608,N_12120);
and U19480 (N_19480,N_13583,N_15222);
xor U19481 (N_19481,N_14742,N_12959);
or U19482 (N_19482,N_12948,N_13619);
xor U19483 (N_19483,N_12463,N_13578);
and U19484 (N_19484,N_15810,N_14331);
or U19485 (N_19485,N_13449,N_12617);
and U19486 (N_19486,N_15456,N_15189);
nand U19487 (N_19487,N_12691,N_14174);
nand U19488 (N_19488,N_15981,N_14693);
nand U19489 (N_19489,N_12651,N_12504);
or U19490 (N_19490,N_14447,N_14926);
nand U19491 (N_19491,N_12822,N_13548);
and U19492 (N_19492,N_14559,N_14322);
nand U19493 (N_19493,N_12918,N_15859);
nand U19494 (N_19494,N_14218,N_12222);
nor U19495 (N_19495,N_14543,N_14029);
xnor U19496 (N_19496,N_15087,N_12070);
and U19497 (N_19497,N_13751,N_13899);
or U19498 (N_19498,N_13980,N_12773);
nor U19499 (N_19499,N_15674,N_15992);
or U19500 (N_19500,N_14349,N_12206);
nand U19501 (N_19501,N_14958,N_12265);
nand U19502 (N_19502,N_14412,N_14726);
or U19503 (N_19503,N_15884,N_13507);
nor U19504 (N_19504,N_13962,N_13164);
nand U19505 (N_19505,N_12412,N_15988);
xnor U19506 (N_19506,N_15636,N_12943);
and U19507 (N_19507,N_13866,N_14098);
nand U19508 (N_19508,N_14988,N_13488);
xnor U19509 (N_19509,N_15470,N_15466);
and U19510 (N_19510,N_13481,N_15163);
nand U19511 (N_19511,N_14438,N_12034);
and U19512 (N_19512,N_15222,N_14003);
or U19513 (N_19513,N_13738,N_12499);
and U19514 (N_19514,N_13202,N_13318);
and U19515 (N_19515,N_12917,N_13097);
and U19516 (N_19516,N_15435,N_12269);
nand U19517 (N_19517,N_15406,N_15528);
or U19518 (N_19518,N_14223,N_13460);
nand U19519 (N_19519,N_15930,N_12926);
or U19520 (N_19520,N_12280,N_13055);
nand U19521 (N_19521,N_12985,N_13949);
xnor U19522 (N_19522,N_14065,N_14852);
nand U19523 (N_19523,N_15123,N_12677);
or U19524 (N_19524,N_13988,N_15558);
nor U19525 (N_19525,N_15887,N_14568);
nand U19526 (N_19526,N_13336,N_14817);
nor U19527 (N_19527,N_14974,N_14869);
nand U19528 (N_19528,N_13517,N_12683);
or U19529 (N_19529,N_12064,N_12848);
nor U19530 (N_19530,N_12121,N_12923);
or U19531 (N_19531,N_13645,N_13797);
or U19532 (N_19532,N_12654,N_14196);
nand U19533 (N_19533,N_12351,N_12484);
nor U19534 (N_19534,N_12829,N_14348);
and U19535 (N_19535,N_12250,N_15626);
and U19536 (N_19536,N_13103,N_15571);
nor U19537 (N_19537,N_15766,N_15408);
xor U19538 (N_19538,N_13713,N_14200);
or U19539 (N_19539,N_12454,N_12144);
nor U19540 (N_19540,N_14449,N_12083);
nor U19541 (N_19541,N_13100,N_13401);
nand U19542 (N_19542,N_12225,N_13246);
and U19543 (N_19543,N_15662,N_15021);
and U19544 (N_19544,N_15067,N_13431);
nand U19545 (N_19545,N_13267,N_15889);
and U19546 (N_19546,N_14379,N_13583);
or U19547 (N_19547,N_14763,N_13866);
nor U19548 (N_19548,N_15846,N_13620);
nand U19549 (N_19549,N_13664,N_13474);
nand U19550 (N_19550,N_15791,N_13175);
xnor U19551 (N_19551,N_14993,N_14080);
xor U19552 (N_19552,N_15513,N_13579);
or U19553 (N_19553,N_14075,N_15069);
nand U19554 (N_19554,N_14047,N_13914);
nor U19555 (N_19555,N_14474,N_12964);
and U19556 (N_19556,N_13336,N_14062);
or U19557 (N_19557,N_12860,N_13736);
and U19558 (N_19558,N_12394,N_13546);
or U19559 (N_19559,N_12073,N_15989);
or U19560 (N_19560,N_13599,N_14780);
xnor U19561 (N_19561,N_15828,N_13240);
and U19562 (N_19562,N_12583,N_15758);
nand U19563 (N_19563,N_15433,N_14228);
or U19564 (N_19564,N_14643,N_12217);
nor U19565 (N_19565,N_15427,N_12332);
nor U19566 (N_19566,N_15384,N_12363);
nand U19567 (N_19567,N_14262,N_12169);
nand U19568 (N_19568,N_13542,N_12096);
nor U19569 (N_19569,N_15649,N_14168);
or U19570 (N_19570,N_13973,N_12343);
or U19571 (N_19571,N_13868,N_12739);
nor U19572 (N_19572,N_14126,N_12678);
xnor U19573 (N_19573,N_13992,N_14319);
nand U19574 (N_19574,N_15702,N_15608);
nand U19575 (N_19575,N_15706,N_13951);
or U19576 (N_19576,N_12212,N_12469);
or U19577 (N_19577,N_14584,N_15080);
and U19578 (N_19578,N_15817,N_15573);
or U19579 (N_19579,N_14146,N_13283);
nor U19580 (N_19580,N_15055,N_12310);
or U19581 (N_19581,N_13418,N_12786);
nand U19582 (N_19582,N_12504,N_13501);
nand U19583 (N_19583,N_14396,N_13199);
nor U19584 (N_19584,N_14359,N_12576);
or U19585 (N_19585,N_14499,N_14530);
or U19586 (N_19586,N_15554,N_14720);
or U19587 (N_19587,N_14073,N_13790);
nand U19588 (N_19588,N_12778,N_12342);
or U19589 (N_19589,N_13606,N_12465);
and U19590 (N_19590,N_12470,N_12378);
nor U19591 (N_19591,N_12116,N_12480);
nor U19592 (N_19592,N_12083,N_14427);
nor U19593 (N_19593,N_13983,N_15099);
nand U19594 (N_19594,N_12701,N_15261);
or U19595 (N_19595,N_15638,N_15245);
nand U19596 (N_19596,N_13596,N_12586);
and U19597 (N_19597,N_12777,N_13580);
and U19598 (N_19598,N_15784,N_12746);
or U19599 (N_19599,N_12311,N_12897);
nand U19600 (N_19600,N_12630,N_14827);
nor U19601 (N_19601,N_14263,N_15210);
nand U19602 (N_19602,N_12362,N_15468);
nor U19603 (N_19603,N_15557,N_15664);
and U19604 (N_19604,N_14115,N_13040);
and U19605 (N_19605,N_12705,N_14776);
and U19606 (N_19606,N_13979,N_14688);
xnor U19607 (N_19607,N_15512,N_13573);
nor U19608 (N_19608,N_12861,N_14163);
nor U19609 (N_19609,N_13529,N_12737);
or U19610 (N_19610,N_14069,N_12362);
nor U19611 (N_19611,N_15778,N_14770);
nor U19612 (N_19612,N_14900,N_13804);
or U19613 (N_19613,N_13430,N_13418);
nor U19614 (N_19614,N_12614,N_14390);
nand U19615 (N_19615,N_13203,N_15766);
xor U19616 (N_19616,N_14608,N_13147);
xor U19617 (N_19617,N_15546,N_15958);
nor U19618 (N_19618,N_15768,N_13861);
nand U19619 (N_19619,N_13251,N_13838);
and U19620 (N_19620,N_13426,N_12923);
or U19621 (N_19621,N_14196,N_14132);
nor U19622 (N_19622,N_12967,N_14382);
xnor U19623 (N_19623,N_15948,N_12608);
nor U19624 (N_19624,N_13420,N_12235);
nor U19625 (N_19625,N_14390,N_12970);
xnor U19626 (N_19626,N_14594,N_13073);
xnor U19627 (N_19627,N_13890,N_13327);
or U19628 (N_19628,N_13319,N_14706);
nor U19629 (N_19629,N_15867,N_14304);
nor U19630 (N_19630,N_12161,N_15013);
nand U19631 (N_19631,N_13339,N_13104);
xnor U19632 (N_19632,N_15256,N_14906);
and U19633 (N_19633,N_14577,N_13806);
and U19634 (N_19634,N_14976,N_13135);
and U19635 (N_19635,N_13720,N_12057);
and U19636 (N_19636,N_15359,N_13545);
and U19637 (N_19637,N_13267,N_15366);
and U19638 (N_19638,N_12514,N_14874);
nor U19639 (N_19639,N_15737,N_13213);
and U19640 (N_19640,N_14634,N_12969);
and U19641 (N_19641,N_15738,N_14354);
and U19642 (N_19642,N_14340,N_15580);
and U19643 (N_19643,N_15487,N_15111);
and U19644 (N_19644,N_13144,N_12468);
and U19645 (N_19645,N_14703,N_14570);
and U19646 (N_19646,N_15810,N_14505);
and U19647 (N_19647,N_12209,N_14250);
nand U19648 (N_19648,N_13070,N_13347);
nand U19649 (N_19649,N_14768,N_15190);
nand U19650 (N_19650,N_12381,N_14455);
and U19651 (N_19651,N_14298,N_15478);
xnor U19652 (N_19652,N_13642,N_14492);
or U19653 (N_19653,N_12092,N_12590);
and U19654 (N_19654,N_15110,N_15182);
and U19655 (N_19655,N_12996,N_13489);
or U19656 (N_19656,N_15132,N_14541);
and U19657 (N_19657,N_13026,N_15700);
and U19658 (N_19658,N_15663,N_15503);
and U19659 (N_19659,N_12584,N_13607);
and U19660 (N_19660,N_15841,N_12252);
and U19661 (N_19661,N_15234,N_14320);
or U19662 (N_19662,N_13408,N_13674);
nor U19663 (N_19663,N_15099,N_14984);
and U19664 (N_19664,N_12191,N_15977);
xnor U19665 (N_19665,N_12344,N_15820);
nor U19666 (N_19666,N_12853,N_15242);
or U19667 (N_19667,N_14179,N_15638);
nor U19668 (N_19668,N_13680,N_13205);
and U19669 (N_19669,N_15360,N_15877);
nand U19670 (N_19670,N_13945,N_12486);
and U19671 (N_19671,N_12994,N_14323);
nand U19672 (N_19672,N_14681,N_14318);
or U19673 (N_19673,N_12555,N_13147);
and U19674 (N_19674,N_13352,N_15793);
and U19675 (N_19675,N_15257,N_12593);
nand U19676 (N_19676,N_15033,N_14192);
and U19677 (N_19677,N_12785,N_12055);
and U19678 (N_19678,N_12899,N_13103);
and U19679 (N_19679,N_13347,N_12730);
xor U19680 (N_19680,N_14248,N_14724);
nor U19681 (N_19681,N_12144,N_13025);
nor U19682 (N_19682,N_12428,N_12015);
nor U19683 (N_19683,N_13672,N_12691);
and U19684 (N_19684,N_15694,N_12756);
nor U19685 (N_19685,N_14266,N_15040);
nor U19686 (N_19686,N_15645,N_12482);
and U19687 (N_19687,N_13738,N_14288);
nor U19688 (N_19688,N_12048,N_12055);
xor U19689 (N_19689,N_12199,N_15272);
or U19690 (N_19690,N_14460,N_13690);
or U19691 (N_19691,N_13518,N_14751);
nor U19692 (N_19692,N_13674,N_14869);
or U19693 (N_19693,N_14463,N_14589);
nand U19694 (N_19694,N_12676,N_12686);
and U19695 (N_19695,N_14326,N_12584);
and U19696 (N_19696,N_12249,N_15520);
nand U19697 (N_19697,N_13350,N_15914);
nand U19698 (N_19698,N_15715,N_15150);
and U19699 (N_19699,N_14207,N_13399);
nor U19700 (N_19700,N_13730,N_15304);
nor U19701 (N_19701,N_12741,N_14337);
or U19702 (N_19702,N_15816,N_12889);
nor U19703 (N_19703,N_12480,N_13061);
nor U19704 (N_19704,N_12886,N_13543);
or U19705 (N_19705,N_13532,N_13282);
xnor U19706 (N_19706,N_13846,N_14602);
xor U19707 (N_19707,N_12868,N_14695);
nor U19708 (N_19708,N_14065,N_12480);
or U19709 (N_19709,N_12177,N_13395);
nor U19710 (N_19710,N_12203,N_14885);
and U19711 (N_19711,N_13405,N_14510);
or U19712 (N_19712,N_12884,N_13295);
nor U19713 (N_19713,N_13218,N_15011);
nand U19714 (N_19714,N_15856,N_14878);
nor U19715 (N_19715,N_13278,N_15160);
and U19716 (N_19716,N_13173,N_12273);
or U19717 (N_19717,N_12886,N_15776);
or U19718 (N_19718,N_15078,N_13761);
xnor U19719 (N_19719,N_12058,N_13210);
nor U19720 (N_19720,N_15204,N_13714);
nor U19721 (N_19721,N_12418,N_14046);
and U19722 (N_19722,N_14570,N_14224);
and U19723 (N_19723,N_14768,N_14175);
or U19724 (N_19724,N_13197,N_14725);
and U19725 (N_19725,N_15115,N_15215);
nand U19726 (N_19726,N_13127,N_12705);
or U19727 (N_19727,N_14389,N_12037);
and U19728 (N_19728,N_12581,N_15638);
nand U19729 (N_19729,N_13269,N_13667);
xor U19730 (N_19730,N_14048,N_13215);
xor U19731 (N_19731,N_14606,N_15165);
nor U19732 (N_19732,N_13137,N_15034);
or U19733 (N_19733,N_15159,N_15426);
nor U19734 (N_19734,N_14155,N_14158);
and U19735 (N_19735,N_14953,N_13706);
or U19736 (N_19736,N_14261,N_14494);
and U19737 (N_19737,N_13037,N_15557);
and U19738 (N_19738,N_15793,N_12360);
nand U19739 (N_19739,N_15611,N_15125);
and U19740 (N_19740,N_13649,N_13190);
and U19741 (N_19741,N_12474,N_12307);
nor U19742 (N_19742,N_14856,N_15422);
xor U19743 (N_19743,N_15612,N_15305);
and U19744 (N_19744,N_14215,N_14509);
or U19745 (N_19745,N_13720,N_13207);
and U19746 (N_19746,N_14020,N_15085);
or U19747 (N_19747,N_15846,N_15446);
nor U19748 (N_19748,N_14909,N_13151);
and U19749 (N_19749,N_13718,N_12253);
or U19750 (N_19750,N_14343,N_12937);
or U19751 (N_19751,N_12831,N_14335);
nand U19752 (N_19752,N_13345,N_13034);
or U19753 (N_19753,N_12499,N_13595);
nor U19754 (N_19754,N_15602,N_12662);
nor U19755 (N_19755,N_13428,N_14215);
nand U19756 (N_19756,N_14171,N_12111);
nor U19757 (N_19757,N_15903,N_15108);
nor U19758 (N_19758,N_12455,N_14005);
xnor U19759 (N_19759,N_15959,N_15120);
xnor U19760 (N_19760,N_15053,N_14947);
nand U19761 (N_19761,N_12897,N_13652);
or U19762 (N_19762,N_13263,N_12811);
and U19763 (N_19763,N_15856,N_12921);
xor U19764 (N_19764,N_13842,N_13210);
nand U19765 (N_19765,N_12391,N_12445);
nor U19766 (N_19766,N_12833,N_14112);
and U19767 (N_19767,N_13586,N_13562);
and U19768 (N_19768,N_12359,N_13034);
or U19769 (N_19769,N_14663,N_12744);
and U19770 (N_19770,N_15422,N_14773);
and U19771 (N_19771,N_12784,N_14535);
or U19772 (N_19772,N_14036,N_14629);
and U19773 (N_19773,N_13754,N_13180);
or U19774 (N_19774,N_14530,N_12891);
or U19775 (N_19775,N_12537,N_15760);
nand U19776 (N_19776,N_14678,N_14054);
nand U19777 (N_19777,N_12924,N_15092);
and U19778 (N_19778,N_13822,N_13998);
or U19779 (N_19779,N_14184,N_15709);
and U19780 (N_19780,N_15654,N_12292);
and U19781 (N_19781,N_15422,N_15033);
and U19782 (N_19782,N_14260,N_14733);
nor U19783 (N_19783,N_13367,N_13639);
and U19784 (N_19784,N_15976,N_12364);
nor U19785 (N_19785,N_12453,N_13796);
nand U19786 (N_19786,N_15195,N_14169);
nor U19787 (N_19787,N_13611,N_15880);
nor U19788 (N_19788,N_13563,N_14716);
nand U19789 (N_19789,N_15022,N_13279);
nand U19790 (N_19790,N_13569,N_13201);
nand U19791 (N_19791,N_12876,N_15957);
nor U19792 (N_19792,N_12798,N_13107);
and U19793 (N_19793,N_15017,N_14776);
xnor U19794 (N_19794,N_15265,N_15711);
or U19795 (N_19795,N_15780,N_12529);
and U19796 (N_19796,N_12679,N_13887);
nor U19797 (N_19797,N_12307,N_14161);
xor U19798 (N_19798,N_13007,N_13800);
and U19799 (N_19799,N_15464,N_14067);
or U19800 (N_19800,N_14690,N_12994);
nand U19801 (N_19801,N_12485,N_12908);
or U19802 (N_19802,N_12129,N_13625);
nand U19803 (N_19803,N_12495,N_12277);
or U19804 (N_19804,N_15482,N_12338);
nor U19805 (N_19805,N_15247,N_13928);
or U19806 (N_19806,N_13635,N_13103);
and U19807 (N_19807,N_12764,N_12749);
or U19808 (N_19808,N_14312,N_14119);
or U19809 (N_19809,N_15961,N_13484);
nor U19810 (N_19810,N_12091,N_13159);
nor U19811 (N_19811,N_13417,N_12288);
and U19812 (N_19812,N_14036,N_15939);
nand U19813 (N_19813,N_13355,N_13096);
and U19814 (N_19814,N_12069,N_14294);
or U19815 (N_19815,N_12696,N_13946);
nor U19816 (N_19816,N_12858,N_13737);
nor U19817 (N_19817,N_15854,N_14090);
and U19818 (N_19818,N_13677,N_12535);
or U19819 (N_19819,N_14290,N_15180);
nand U19820 (N_19820,N_13909,N_13211);
nand U19821 (N_19821,N_12914,N_13520);
or U19822 (N_19822,N_15403,N_14090);
nor U19823 (N_19823,N_13195,N_14240);
and U19824 (N_19824,N_14710,N_12352);
nor U19825 (N_19825,N_13312,N_15969);
nand U19826 (N_19826,N_15346,N_15852);
and U19827 (N_19827,N_15551,N_13168);
nor U19828 (N_19828,N_14589,N_12298);
nand U19829 (N_19829,N_12478,N_15841);
nor U19830 (N_19830,N_14138,N_14522);
nand U19831 (N_19831,N_14162,N_13667);
nand U19832 (N_19832,N_13825,N_14739);
nor U19833 (N_19833,N_14784,N_13772);
nor U19834 (N_19834,N_13209,N_12691);
and U19835 (N_19835,N_13884,N_14004);
nand U19836 (N_19836,N_13307,N_15209);
and U19837 (N_19837,N_15356,N_13728);
and U19838 (N_19838,N_15507,N_15368);
nor U19839 (N_19839,N_12140,N_14679);
or U19840 (N_19840,N_12266,N_12769);
nand U19841 (N_19841,N_13761,N_15156);
or U19842 (N_19842,N_14916,N_14918);
nor U19843 (N_19843,N_13028,N_13646);
or U19844 (N_19844,N_14131,N_14013);
nor U19845 (N_19845,N_15399,N_12813);
and U19846 (N_19846,N_14398,N_14006);
nand U19847 (N_19847,N_14720,N_12330);
nor U19848 (N_19848,N_13735,N_12366);
nor U19849 (N_19849,N_12283,N_14522);
nor U19850 (N_19850,N_12022,N_13867);
xor U19851 (N_19851,N_12503,N_14930);
xnor U19852 (N_19852,N_13627,N_12448);
nand U19853 (N_19853,N_15646,N_15289);
nor U19854 (N_19854,N_12967,N_13977);
or U19855 (N_19855,N_14795,N_13901);
nand U19856 (N_19856,N_12273,N_15826);
nor U19857 (N_19857,N_12237,N_14969);
nor U19858 (N_19858,N_14648,N_15579);
nand U19859 (N_19859,N_14964,N_15353);
and U19860 (N_19860,N_15212,N_14095);
nor U19861 (N_19861,N_14371,N_15160);
and U19862 (N_19862,N_12634,N_15143);
nand U19863 (N_19863,N_14235,N_13083);
or U19864 (N_19864,N_14702,N_14938);
and U19865 (N_19865,N_14025,N_13138);
and U19866 (N_19866,N_12315,N_12630);
nor U19867 (N_19867,N_14642,N_13283);
nand U19868 (N_19868,N_13180,N_12170);
nand U19869 (N_19869,N_15245,N_12889);
and U19870 (N_19870,N_12588,N_12192);
nand U19871 (N_19871,N_12356,N_15889);
nor U19872 (N_19872,N_13144,N_12832);
and U19873 (N_19873,N_13284,N_12556);
nand U19874 (N_19874,N_13524,N_14706);
xor U19875 (N_19875,N_14926,N_12744);
nor U19876 (N_19876,N_15138,N_14447);
nor U19877 (N_19877,N_13909,N_12516);
nor U19878 (N_19878,N_15003,N_12131);
or U19879 (N_19879,N_13736,N_15198);
nand U19880 (N_19880,N_13675,N_13215);
or U19881 (N_19881,N_12517,N_12732);
and U19882 (N_19882,N_13071,N_13564);
and U19883 (N_19883,N_13550,N_13553);
and U19884 (N_19884,N_13933,N_13176);
nor U19885 (N_19885,N_12351,N_13608);
and U19886 (N_19886,N_14919,N_13222);
and U19887 (N_19887,N_14219,N_15041);
nor U19888 (N_19888,N_15750,N_14218);
or U19889 (N_19889,N_12949,N_15286);
nor U19890 (N_19890,N_13731,N_15767);
or U19891 (N_19891,N_15202,N_13537);
nor U19892 (N_19892,N_13302,N_15322);
nand U19893 (N_19893,N_12430,N_12199);
nor U19894 (N_19894,N_12801,N_12552);
nor U19895 (N_19895,N_14297,N_15814);
or U19896 (N_19896,N_13944,N_13846);
nor U19897 (N_19897,N_15333,N_15597);
xor U19898 (N_19898,N_15541,N_12226);
nand U19899 (N_19899,N_15090,N_15035);
nor U19900 (N_19900,N_12119,N_13889);
and U19901 (N_19901,N_13557,N_15010);
or U19902 (N_19902,N_12232,N_15311);
xor U19903 (N_19903,N_13154,N_14616);
and U19904 (N_19904,N_14699,N_15405);
nand U19905 (N_19905,N_12936,N_14322);
or U19906 (N_19906,N_15167,N_13355);
or U19907 (N_19907,N_14466,N_13433);
nand U19908 (N_19908,N_13944,N_15015);
or U19909 (N_19909,N_12979,N_13462);
and U19910 (N_19910,N_15888,N_12652);
nor U19911 (N_19911,N_14069,N_13741);
and U19912 (N_19912,N_12458,N_14984);
and U19913 (N_19913,N_15168,N_15283);
nand U19914 (N_19914,N_15172,N_13110);
nand U19915 (N_19915,N_13005,N_14251);
nand U19916 (N_19916,N_12853,N_13598);
or U19917 (N_19917,N_15926,N_15639);
and U19918 (N_19918,N_14755,N_12928);
xnor U19919 (N_19919,N_12121,N_13276);
nand U19920 (N_19920,N_15802,N_13307);
nand U19921 (N_19921,N_15308,N_14641);
nand U19922 (N_19922,N_13318,N_14082);
nor U19923 (N_19923,N_13783,N_13433);
nand U19924 (N_19924,N_14509,N_12408);
nor U19925 (N_19925,N_14947,N_13897);
nand U19926 (N_19926,N_13943,N_13805);
nor U19927 (N_19927,N_12961,N_13947);
nand U19928 (N_19928,N_15744,N_12564);
nand U19929 (N_19929,N_14086,N_13307);
and U19930 (N_19930,N_14776,N_14305);
nor U19931 (N_19931,N_12970,N_13086);
nand U19932 (N_19932,N_13922,N_14058);
or U19933 (N_19933,N_13318,N_12365);
xnor U19934 (N_19934,N_14691,N_14247);
or U19935 (N_19935,N_14610,N_15143);
and U19936 (N_19936,N_12840,N_13931);
xnor U19937 (N_19937,N_14867,N_12074);
or U19938 (N_19938,N_12292,N_14161);
or U19939 (N_19939,N_14618,N_12288);
and U19940 (N_19940,N_15586,N_14894);
and U19941 (N_19941,N_15392,N_15262);
nand U19942 (N_19942,N_14300,N_14603);
nor U19943 (N_19943,N_14272,N_12323);
or U19944 (N_19944,N_14353,N_13103);
nor U19945 (N_19945,N_14171,N_13947);
or U19946 (N_19946,N_12714,N_12970);
and U19947 (N_19947,N_12005,N_12074);
or U19948 (N_19948,N_13477,N_13445);
nor U19949 (N_19949,N_15545,N_13985);
and U19950 (N_19950,N_15642,N_14923);
and U19951 (N_19951,N_13822,N_13139);
nand U19952 (N_19952,N_14499,N_12282);
or U19953 (N_19953,N_14985,N_14544);
nand U19954 (N_19954,N_12764,N_14732);
or U19955 (N_19955,N_14538,N_15480);
nor U19956 (N_19956,N_14766,N_12991);
nor U19957 (N_19957,N_15292,N_12344);
nand U19958 (N_19958,N_15520,N_14212);
and U19959 (N_19959,N_15926,N_13296);
nor U19960 (N_19960,N_12700,N_13329);
or U19961 (N_19961,N_12685,N_12853);
and U19962 (N_19962,N_15121,N_12975);
and U19963 (N_19963,N_12506,N_15409);
or U19964 (N_19964,N_13489,N_15703);
nand U19965 (N_19965,N_12898,N_12305);
and U19966 (N_19966,N_13291,N_13460);
and U19967 (N_19967,N_12570,N_14825);
and U19968 (N_19968,N_15498,N_13382);
and U19969 (N_19969,N_14910,N_13906);
and U19970 (N_19970,N_12705,N_13174);
xor U19971 (N_19971,N_15960,N_13360);
nor U19972 (N_19972,N_13479,N_15449);
and U19973 (N_19973,N_14901,N_13334);
nand U19974 (N_19974,N_13596,N_13756);
or U19975 (N_19975,N_14371,N_13629);
and U19976 (N_19976,N_13111,N_15597);
and U19977 (N_19977,N_15018,N_14833);
nand U19978 (N_19978,N_13776,N_12617);
or U19979 (N_19979,N_14852,N_15822);
nor U19980 (N_19980,N_13019,N_12597);
xnor U19981 (N_19981,N_12687,N_14440);
xor U19982 (N_19982,N_14053,N_15934);
nor U19983 (N_19983,N_13884,N_14232);
nor U19984 (N_19984,N_13216,N_15714);
xor U19985 (N_19985,N_12113,N_13503);
and U19986 (N_19986,N_13886,N_15573);
or U19987 (N_19987,N_14190,N_15731);
nor U19988 (N_19988,N_14867,N_12193);
and U19989 (N_19989,N_13050,N_15518);
xor U19990 (N_19990,N_14804,N_12783);
or U19991 (N_19991,N_14009,N_13966);
nor U19992 (N_19992,N_12706,N_13333);
nand U19993 (N_19993,N_15514,N_14817);
nand U19994 (N_19994,N_15551,N_14480);
and U19995 (N_19995,N_15257,N_13771);
nand U19996 (N_19996,N_12562,N_13856);
and U19997 (N_19997,N_12556,N_13418);
and U19998 (N_19998,N_15457,N_12095);
nand U19999 (N_19999,N_14313,N_12770);
or UO_0 (O_0,N_19334,N_19485);
nor UO_1 (O_1,N_19758,N_16481);
or UO_2 (O_2,N_18633,N_16932);
nand UO_3 (O_3,N_18483,N_16482);
or UO_4 (O_4,N_18968,N_19886);
and UO_5 (O_5,N_17999,N_18618);
and UO_6 (O_6,N_17371,N_18791);
nor UO_7 (O_7,N_17148,N_19703);
or UO_8 (O_8,N_17520,N_17865);
and UO_9 (O_9,N_19123,N_19373);
or UO_10 (O_10,N_17717,N_16365);
or UO_11 (O_11,N_19005,N_17483);
or UO_12 (O_12,N_16814,N_18585);
and UO_13 (O_13,N_17008,N_17210);
nand UO_14 (O_14,N_19844,N_17073);
or UO_15 (O_15,N_16632,N_18136);
and UO_16 (O_16,N_19283,N_17860);
or UO_17 (O_17,N_19942,N_19785);
and UO_18 (O_18,N_17002,N_19291);
nand UO_19 (O_19,N_17643,N_19549);
nor UO_20 (O_20,N_17415,N_16379);
and UO_21 (O_21,N_18463,N_17453);
xor UO_22 (O_22,N_16108,N_16529);
nor UO_23 (O_23,N_17428,N_16967);
or UO_24 (O_24,N_19576,N_16975);
nand UO_25 (O_25,N_18389,N_17747);
and UO_26 (O_26,N_16807,N_19352);
nand UO_27 (O_27,N_19524,N_18787);
nand UO_28 (O_28,N_16968,N_17866);
or UO_29 (O_29,N_19574,N_19353);
nor UO_30 (O_30,N_17726,N_17753);
xor UO_31 (O_31,N_16327,N_19708);
nor UO_32 (O_32,N_16019,N_16935);
or UO_33 (O_33,N_18356,N_17142);
or UO_34 (O_34,N_16897,N_16462);
or UO_35 (O_35,N_18632,N_17886);
nor UO_36 (O_36,N_17572,N_18885);
and UO_37 (O_37,N_16562,N_19384);
nand UO_38 (O_38,N_19985,N_16691);
nand UO_39 (O_39,N_18249,N_16472);
nand UO_40 (O_40,N_19997,N_16816);
nand UO_41 (O_41,N_17405,N_18847);
nor UO_42 (O_42,N_16701,N_17198);
or UO_43 (O_43,N_16372,N_18478);
nand UO_44 (O_44,N_16704,N_18371);
and UO_45 (O_45,N_19022,N_17580);
and UO_46 (O_46,N_18010,N_19316);
or UO_47 (O_47,N_17131,N_18309);
nand UO_48 (O_48,N_16493,N_18383);
nand UO_49 (O_49,N_16722,N_16026);
nand UO_50 (O_50,N_18454,N_19233);
or UO_51 (O_51,N_19422,N_19602);
nand UO_52 (O_52,N_18416,N_16188);
nand UO_53 (O_53,N_18964,N_17793);
nand UO_54 (O_54,N_18451,N_18536);
or UO_55 (O_55,N_16063,N_17461);
and UO_56 (O_56,N_18688,N_19300);
xnor UO_57 (O_57,N_19766,N_18734);
nor UO_58 (O_58,N_18019,N_17554);
nand UO_59 (O_59,N_19404,N_16485);
nor UO_60 (O_60,N_19925,N_18750);
and UO_61 (O_61,N_16764,N_17792);
nand UO_62 (O_62,N_16219,N_17834);
and UO_63 (O_63,N_19967,N_19717);
and UO_64 (O_64,N_18548,N_17235);
xnor UO_65 (O_65,N_17806,N_17034);
nand UO_66 (O_66,N_18907,N_16155);
xor UO_67 (O_67,N_17993,N_17233);
and UO_68 (O_68,N_16329,N_17840);
or UO_69 (O_69,N_18859,N_19526);
and UO_70 (O_70,N_17634,N_19666);
or UO_71 (O_71,N_19116,N_16099);
and UO_72 (O_72,N_17317,N_19722);
or UO_73 (O_73,N_19782,N_19581);
nor UO_74 (O_74,N_16004,N_16668);
nand UO_75 (O_75,N_16328,N_16688);
nand UO_76 (O_76,N_16696,N_18944);
and UO_77 (O_77,N_17045,N_18628);
and UO_78 (O_78,N_18367,N_18197);
nand UO_79 (O_79,N_16030,N_18870);
nor UO_80 (O_80,N_18426,N_19519);
nand UO_81 (O_81,N_16166,N_16777);
and UO_82 (O_82,N_19220,N_17535);
and UO_83 (O_83,N_17375,N_16159);
nand UO_84 (O_84,N_19684,N_19775);
nor UO_85 (O_85,N_16123,N_19090);
and UO_86 (O_86,N_18857,N_16721);
or UO_87 (O_87,N_16341,N_18247);
and UO_88 (O_88,N_17963,N_18834);
and UO_89 (O_89,N_18557,N_16474);
and UO_90 (O_90,N_18140,N_18578);
or UO_91 (O_91,N_16259,N_18098);
or UO_92 (O_92,N_16793,N_17651);
nand UO_93 (O_93,N_16920,N_16959);
and UO_94 (O_94,N_17009,N_18363);
xnor UO_95 (O_95,N_16009,N_18241);
nor UO_96 (O_96,N_16150,N_17475);
nor UO_97 (O_97,N_17638,N_19618);
nand UO_98 (O_98,N_16742,N_17410);
nor UO_99 (O_99,N_18313,N_19660);
and UO_100 (O_100,N_16496,N_16825);
nand UO_101 (O_101,N_17144,N_19041);
nand UO_102 (O_102,N_16037,N_16244);
nand UO_103 (O_103,N_17991,N_16455);
or UO_104 (O_104,N_16132,N_18992);
or UO_105 (O_105,N_16989,N_16450);
nor UO_106 (O_106,N_19608,N_18147);
xnor UO_107 (O_107,N_17463,N_18473);
nand UO_108 (O_108,N_16772,N_18533);
or UO_109 (O_109,N_17730,N_18038);
nand UO_110 (O_110,N_16076,N_19266);
nand UO_111 (O_111,N_18550,N_16656);
nand UO_112 (O_112,N_19583,N_17671);
and UO_113 (O_113,N_17703,N_19294);
nor UO_114 (O_114,N_18767,N_16014);
or UO_115 (O_115,N_18500,N_16670);
xor UO_116 (O_116,N_16468,N_17675);
nand UO_117 (O_117,N_19950,N_16012);
and UO_118 (O_118,N_17681,N_16234);
nor UO_119 (O_119,N_19657,N_16380);
or UO_120 (O_120,N_16494,N_17464);
and UO_121 (O_121,N_16867,N_18599);
nand UO_122 (O_122,N_17560,N_18259);
nand UO_123 (O_123,N_19752,N_19446);
and UO_124 (O_124,N_17723,N_17394);
or UO_125 (O_125,N_18017,N_16408);
nand UO_126 (O_126,N_19386,N_17725);
nand UO_127 (O_127,N_17534,N_16045);
nor UO_128 (O_128,N_19186,N_19955);
or UO_129 (O_129,N_17745,N_18030);
nor UO_130 (O_130,N_17610,N_19535);
or UO_131 (O_131,N_16331,N_19982);
nor UO_132 (O_132,N_19258,N_16981);
nor UO_133 (O_133,N_16788,N_17019);
and UO_134 (O_134,N_16401,N_18830);
or UO_135 (O_135,N_19147,N_18231);
nor UO_136 (O_136,N_18607,N_16690);
and UO_137 (O_137,N_19757,N_18602);
nand UO_138 (O_138,N_19239,N_16755);
or UO_139 (O_139,N_16241,N_17485);
or UO_140 (O_140,N_19410,N_19028);
nand UO_141 (O_141,N_16820,N_19655);
and UO_142 (O_142,N_17001,N_17076);
nand UO_143 (O_143,N_18687,N_17332);
and UO_144 (O_144,N_17835,N_16808);
nor UO_145 (O_145,N_17875,N_18155);
nand UO_146 (O_146,N_17874,N_17425);
nand UO_147 (O_147,N_19099,N_19144);
nand UO_148 (O_148,N_19207,N_17686);
nand UO_149 (O_149,N_17622,N_18950);
xor UO_150 (O_150,N_19833,N_17462);
xor UO_151 (O_151,N_19457,N_16924);
nand UO_152 (O_152,N_19452,N_17598);
nor UO_153 (O_153,N_17734,N_17669);
nor UO_154 (O_154,N_18138,N_16432);
nor UO_155 (O_155,N_19633,N_18515);
nand UO_156 (O_156,N_16758,N_19781);
and UO_157 (O_157,N_17207,N_19448);
or UO_158 (O_158,N_17872,N_16899);
nand UO_159 (O_159,N_18216,N_18142);
xnor UO_160 (O_160,N_18581,N_19183);
xor UO_161 (O_161,N_18221,N_16386);
or UO_162 (O_162,N_16054,N_19718);
or UO_163 (O_163,N_17075,N_19619);
or UO_164 (O_164,N_17058,N_18446);
and UO_165 (O_165,N_16734,N_17798);
and UO_166 (O_166,N_16437,N_19821);
or UO_167 (O_167,N_17459,N_19237);
nor UO_168 (O_168,N_16747,N_17214);
nor UO_169 (O_169,N_18975,N_19023);
nand UO_170 (O_170,N_18388,N_19394);
xor UO_171 (O_171,N_17500,N_19841);
xnor UO_172 (O_172,N_19382,N_17361);
nand UO_173 (O_173,N_17642,N_19548);
nor UO_174 (O_174,N_16141,N_18493);
nand UO_175 (O_175,N_18883,N_16532);
and UO_176 (O_176,N_18002,N_17647);
nand UO_177 (O_177,N_19351,N_17111);
and UO_178 (O_178,N_17347,N_17659);
or UO_179 (O_179,N_18580,N_17273);
and UO_180 (O_180,N_17672,N_18215);
xnor UO_181 (O_181,N_18627,N_17608);
xnor UO_182 (O_182,N_17417,N_16446);
nand UO_183 (O_183,N_18596,N_17934);
or UO_184 (O_184,N_16441,N_18670);
nand UO_185 (O_185,N_16991,N_19857);
nor UO_186 (O_186,N_16160,N_18936);
xnor UO_187 (O_187,N_18480,N_18253);
and UO_188 (O_188,N_18319,N_19056);
and UO_189 (O_189,N_17773,N_16303);
nand UO_190 (O_190,N_18368,N_17697);
and UO_191 (O_191,N_19432,N_19991);
nand UO_192 (O_192,N_17440,N_17618);
or UO_193 (O_193,N_18920,N_19530);
nand UO_194 (O_194,N_18576,N_19811);
or UO_195 (O_195,N_16459,N_17640);
nand UO_196 (O_196,N_16640,N_18005);
xnor UO_197 (O_197,N_18986,N_19177);
nand UO_198 (O_198,N_16785,N_17949);
xnor UO_199 (O_199,N_18212,N_16598);
or UO_200 (O_200,N_16499,N_17794);
xnor UO_201 (O_201,N_18887,N_18981);
nand UO_202 (O_202,N_17849,N_19280);
nand UO_203 (O_203,N_18046,N_17031);
or UO_204 (O_204,N_18760,N_19122);
nor UO_205 (O_205,N_19687,N_16034);
and UO_206 (O_206,N_17983,N_16585);
and UO_207 (O_207,N_19355,N_18937);
nand UO_208 (O_208,N_16646,N_16636);
xor UO_209 (O_209,N_17816,N_19934);
and UO_210 (O_210,N_19585,N_18331);
and UO_211 (O_211,N_19038,N_16369);
nor UO_212 (O_212,N_17612,N_18504);
xor UO_213 (O_213,N_18900,N_18292);
and UO_214 (O_214,N_16339,N_17842);
and UO_215 (O_215,N_18822,N_17550);
xnor UO_216 (O_216,N_18648,N_16489);
or UO_217 (O_217,N_16537,N_16752);
nand UO_218 (O_218,N_17000,N_18198);
xor UO_219 (O_219,N_19492,N_17270);
nand UO_220 (O_220,N_16792,N_19986);
or UO_221 (O_221,N_17218,N_19630);
or UO_222 (O_222,N_19094,N_16892);
nand UO_223 (O_223,N_18288,N_19265);
nand UO_224 (O_224,N_19286,N_19045);
and UO_225 (O_225,N_19388,N_16837);
or UO_226 (O_226,N_17575,N_17503);
or UO_227 (O_227,N_19802,N_19317);
or UO_228 (O_228,N_19299,N_17829);
and UO_229 (O_229,N_18358,N_17323);
and UO_230 (O_230,N_17900,N_18722);
nor UO_231 (O_231,N_18803,N_18814);
nor UO_232 (O_232,N_17106,N_18893);
or UO_233 (O_233,N_17225,N_17257);
and UO_234 (O_234,N_19001,N_17917);
or UO_235 (O_235,N_17470,N_17698);
or UO_236 (O_236,N_18004,N_16354);
nand UO_237 (O_237,N_17613,N_16046);
nand UO_238 (O_238,N_16194,N_19928);
or UO_239 (O_239,N_16878,N_19674);
or UO_240 (O_240,N_17139,N_16209);
nand UO_241 (O_241,N_19016,N_17518);
or UO_242 (O_242,N_17399,N_19146);
and UO_243 (O_243,N_18284,N_17899);
and UO_244 (O_244,N_18530,N_19486);
nand UO_245 (O_245,N_16253,N_19212);
or UO_246 (O_246,N_17298,N_19557);
and UO_247 (O_247,N_18220,N_17067);
nor UO_248 (O_248,N_16749,N_19990);
and UO_249 (O_249,N_18167,N_18894);
nor UO_250 (O_250,N_19285,N_16488);
nand UO_251 (O_251,N_17928,N_16727);
or UO_252 (O_252,N_17379,N_19203);
xnor UO_253 (O_253,N_17552,N_19228);
nand UO_254 (O_254,N_19085,N_16366);
nand UO_255 (O_255,N_17607,N_18733);
and UO_256 (O_256,N_17517,N_16604);
or UO_257 (O_257,N_19101,N_19849);
nand UO_258 (O_258,N_18774,N_17190);
xnor UO_259 (O_259,N_18380,N_19463);
or UO_260 (O_260,N_18637,N_18616);
xnor UO_261 (O_261,N_17958,N_19272);
nand UO_262 (O_262,N_17123,N_16301);
or UO_263 (O_263,N_19027,N_17576);
nor UO_264 (O_264,N_17915,N_16821);
xnor UO_265 (O_265,N_19540,N_16884);
nand UO_266 (O_266,N_17937,N_16249);
nor UO_267 (O_267,N_16660,N_18877);
or UO_268 (O_268,N_16900,N_18890);
nand UO_269 (O_269,N_17290,N_18012);
nor UO_270 (O_270,N_18556,N_17978);
and UO_271 (O_271,N_19973,N_17163);
nand UO_272 (O_272,N_19431,N_16635);
or UO_273 (O_273,N_19277,N_19555);
nor UO_274 (O_274,N_17484,N_16578);
and UO_275 (O_275,N_16676,N_16436);
xnor UO_276 (O_276,N_17781,N_18832);
or UO_277 (O_277,N_16838,N_17695);
and UO_278 (O_278,N_18617,N_16733);
nand UO_279 (O_279,N_19826,N_19761);
nor UO_280 (O_280,N_18267,N_16666);
nand UO_281 (O_281,N_17595,N_16665);
and UO_282 (O_282,N_19140,N_18559);
nand UO_283 (O_283,N_19975,N_18678);
nor UO_284 (O_284,N_19765,N_17340);
nand UO_285 (O_285,N_19776,N_17907);
or UO_286 (O_286,N_18586,N_16414);
nor UO_287 (O_287,N_18328,N_17922);
or UO_288 (O_288,N_17049,N_19161);
or UO_289 (O_289,N_18621,N_16855);
nor UO_290 (O_290,N_18732,N_19582);
and UO_291 (O_291,N_19364,N_18940);
and UO_292 (O_292,N_18558,N_18049);
or UO_293 (O_293,N_16579,N_16297);
and UO_294 (O_294,N_18965,N_19251);
nor UO_295 (O_295,N_19029,N_17504);
xor UO_296 (O_296,N_16138,N_18307);
nor UO_297 (O_297,N_18202,N_18507);
and UO_298 (O_298,N_18043,N_17449);
and UO_299 (O_299,N_18720,N_16395);
or UO_300 (O_300,N_19868,N_19972);
or UO_301 (O_301,N_18845,N_16960);
nor UO_302 (O_302,N_17351,N_17573);
xnor UO_303 (O_303,N_16066,N_18978);
xor UO_304 (O_304,N_18600,N_17339);
nor UO_305 (O_305,N_16038,N_17217);
xor UO_306 (O_306,N_16010,N_18495);
nor UO_307 (O_307,N_16064,N_19960);
xnor UO_308 (O_308,N_18036,N_19411);
nor UO_309 (O_309,N_17166,N_16248);
nand UO_310 (O_310,N_17699,N_17436);
nand UO_311 (O_311,N_18946,N_18692);
nand UO_312 (O_312,N_19504,N_17714);
nor UO_313 (O_313,N_17308,N_19813);
xnor UO_314 (O_314,N_17341,N_19238);
and UO_315 (O_315,N_18948,N_16471);
or UO_316 (O_316,N_17358,N_18315);
or UO_317 (O_317,N_17895,N_17855);
or UO_318 (O_318,N_17941,N_19676);
or UO_319 (O_319,N_18869,N_19862);
and UO_320 (O_320,N_16885,N_19979);
nand UO_321 (O_321,N_18290,N_18126);
nor UO_322 (O_322,N_18994,N_16905);
and UO_323 (O_323,N_18177,N_19401);
nor UO_324 (O_324,N_16970,N_19141);
nor UO_325 (O_325,N_19406,N_17412);
or UO_326 (O_326,N_16547,N_16115);
or UO_327 (O_327,N_16754,N_19458);
nand UO_328 (O_328,N_17487,N_19806);
nor UO_329 (O_329,N_16461,N_18743);
nor UO_330 (O_330,N_18606,N_16332);
nand UO_331 (O_331,N_18825,N_18551);
nor UO_332 (O_332,N_16086,N_16065);
nand UO_333 (O_333,N_17376,N_17022);
xnor UO_334 (O_334,N_18574,N_18158);
and UO_335 (O_335,N_16263,N_17950);
and UO_336 (O_336,N_17283,N_16528);
nor UO_337 (O_337,N_16658,N_16337);
or UO_338 (O_338,N_16768,N_16036);
and UO_339 (O_339,N_16286,N_18006);
xnor UO_340 (O_340,N_16470,N_18310);
or UO_341 (O_341,N_19390,N_18476);
and UO_342 (O_342,N_18271,N_16412);
nand UO_343 (O_343,N_17989,N_17023);
and UO_344 (O_344,N_19187,N_18148);
xnor UO_345 (O_345,N_18087,N_16161);
or UO_346 (O_346,N_19075,N_16685);
and UO_347 (O_347,N_18625,N_18377);
or UO_348 (O_348,N_19043,N_17530);
and UO_349 (O_349,N_16611,N_16879);
xor UO_350 (O_350,N_19319,N_18453);
or UO_351 (O_351,N_17348,N_17059);
nor UO_352 (O_352,N_19741,N_19692);
and UO_353 (O_353,N_19196,N_16023);
nand UO_354 (O_354,N_16302,N_19901);
nor UO_355 (O_355,N_18171,N_18945);
nand UO_356 (O_356,N_18154,N_19668);
xnor UO_357 (O_357,N_16677,N_19387);
and UO_358 (O_358,N_17812,N_17246);
and UO_359 (O_359,N_16292,N_16724);
or UO_360 (O_360,N_18084,N_16678);
and UO_361 (O_361,N_16373,N_19935);
nand UO_362 (O_362,N_16125,N_19250);
nand UO_363 (O_363,N_17896,N_17267);
or UO_364 (O_364,N_17418,N_17799);
nand UO_365 (O_365,N_19261,N_19026);
and UO_366 (O_366,N_16922,N_16048);
and UO_367 (O_367,N_16422,N_18429);
nand UO_368 (O_368,N_16260,N_18631);
nand UO_369 (O_369,N_18462,N_17118);
xor UO_370 (O_370,N_16951,N_17419);
xnor UO_371 (O_371,N_19520,N_16312);
nand UO_372 (O_372,N_16214,N_19638);
and UO_373 (O_373,N_17541,N_16504);
nand UO_374 (O_374,N_18788,N_16164);
nor UO_375 (O_375,N_19624,N_16024);
nand UO_376 (O_376,N_18194,N_17241);
nand UO_377 (O_377,N_17946,N_16864);
or UO_378 (O_378,N_17815,N_18470);
nand UO_379 (O_379,N_16091,N_17141);
and UO_380 (O_380,N_19740,N_18387);
xnor UO_381 (O_381,N_18686,N_16008);
and UO_382 (O_382,N_16671,N_19424);
and UO_383 (O_383,N_19751,N_18527);
nand UO_384 (O_384,N_16149,N_18145);
nand UO_385 (O_385,N_16299,N_19483);
or UO_386 (O_386,N_17708,N_17495);
nand UO_387 (O_387,N_17972,N_16028);
nor UO_388 (O_388,N_19575,N_16972);
and UO_389 (O_389,N_19529,N_19333);
nand UO_390 (O_390,N_16805,N_17515);
and UO_391 (O_391,N_16124,N_18868);
nand UO_392 (O_392,N_16720,N_18698);
or UO_393 (O_393,N_19738,N_17005);
xnor UO_394 (O_394,N_16073,N_19628);
nand UO_395 (O_395,N_17837,N_18534);
or UO_396 (O_396,N_19107,N_19544);
and UO_397 (O_397,N_19667,N_18996);
nor UO_398 (O_398,N_17104,N_16845);
nand UO_399 (O_399,N_17489,N_17955);
or UO_400 (O_400,N_19778,N_19393);
or UO_401 (O_401,N_17635,N_17862);
xor UO_402 (O_402,N_18901,N_17382);
and UO_403 (O_403,N_19421,N_16424);
and UO_404 (O_404,N_17344,N_16243);
or UO_405 (O_405,N_18958,N_18370);
or UO_406 (O_406,N_18614,N_19126);
or UO_407 (O_407,N_18105,N_18011);
and UO_408 (O_408,N_19774,N_19683);
or UO_409 (O_409,N_18914,N_18236);
or UO_410 (O_410,N_18897,N_17599);
nand UO_411 (O_411,N_18187,N_16511);
or UO_412 (O_412,N_19399,N_19307);
and UO_413 (O_413,N_17318,N_17491);
nor UO_414 (O_414,N_18206,N_19400);
or UO_415 (O_415,N_18967,N_17882);
and UO_416 (O_416,N_19691,N_18680);
nand UO_417 (O_417,N_16031,N_16645);
xor UO_418 (O_418,N_18816,N_19527);
and UO_419 (O_419,N_17555,N_18653);
xnor UO_420 (O_420,N_18683,N_19108);
and UO_421 (O_421,N_19603,N_16693);
xor UO_422 (O_422,N_17822,N_16664);
xor UO_423 (O_423,N_17513,N_18780);
xor UO_424 (O_424,N_16990,N_16220);
nand UO_425 (O_425,N_16916,N_16827);
nor UO_426 (O_426,N_19652,N_17346);
and UO_427 (O_427,N_18779,N_18176);
or UO_428 (O_428,N_17960,N_17856);
nand UO_429 (O_429,N_16120,N_19343);
nor UO_430 (O_430,N_19621,N_18754);
or UO_431 (O_431,N_18844,N_19310);
nor UO_432 (O_432,N_18665,N_18498);
or UO_433 (O_433,N_18961,N_18114);
or UO_434 (O_434,N_18445,N_18015);
and UO_435 (O_435,N_19647,N_18406);
nand UO_436 (O_436,N_17039,N_18287);
and UO_437 (O_437,N_17254,N_17673);
nand UO_438 (O_438,N_19842,N_17615);
or UO_439 (O_439,N_17546,N_17401);
xnor UO_440 (O_440,N_19805,N_18184);
or UO_441 (O_441,N_19533,N_17061);
and UO_442 (O_442,N_16451,N_16876);
and UO_443 (O_443,N_16997,N_16180);
nor UO_444 (O_444,N_16443,N_18752);
nor UO_445 (O_445,N_16226,N_18721);
and UO_446 (O_446,N_18379,N_19787);
nand UO_447 (O_447,N_19747,N_17755);
nand UO_448 (O_448,N_19501,N_16254);
and UO_449 (O_449,N_17693,N_16240);
nand UO_450 (O_450,N_16137,N_17446);
and UO_451 (O_451,N_16183,N_19302);
or UO_452 (O_452,N_16929,N_18728);
nor UO_453 (O_453,N_16163,N_19512);
or UO_454 (O_454,N_17762,N_18349);
or UO_455 (O_455,N_16439,N_19951);
or UO_456 (O_456,N_18188,N_17701);
and UO_457 (O_457,N_17288,N_18783);
nand UO_458 (O_458,N_17300,N_16338);
nand UO_459 (O_459,N_16784,N_19423);
nand UO_460 (O_460,N_19433,N_19742);
xnor UO_461 (O_461,N_18839,N_19102);
and UO_462 (O_462,N_17468,N_18793);
nand UO_463 (O_463,N_17398,N_17441);
and UO_464 (O_464,N_17420,N_18689);
nor UO_465 (O_465,N_18702,N_19321);
and UO_466 (O_466,N_16309,N_19830);
or UO_467 (O_467,N_17265,N_16594);
or UO_468 (O_468,N_16333,N_17656);
nand UO_469 (O_469,N_19052,N_16396);
xor UO_470 (O_470,N_19002,N_17334);
or UO_471 (O_471,N_16564,N_18466);
or UO_472 (O_472,N_19464,N_19030);
or UO_473 (O_473,N_18402,N_16089);
nand UO_474 (O_474,N_18073,N_17437);
nand UO_475 (O_475,N_17724,N_17179);
nand UO_476 (O_476,N_16973,N_16130);
and UO_477 (O_477,N_18805,N_16002);
nor UO_478 (O_478,N_19796,N_17797);
nand UO_479 (O_479,N_16427,N_18299);
and UO_480 (O_480,N_19389,N_18304);
nor UO_481 (O_481,N_16616,N_19591);
nor UO_482 (O_482,N_16072,N_18726);
and UO_483 (O_483,N_18737,N_19430);
and UO_484 (O_484,N_18647,N_17191);
and UO_485 (O_485,N_18041,N_18419);
nor UO_486 (O_486,N_18260,N_16445);
or UO_487 (O_487,N_19593,N_17378);
or UO_488 (O_488,N_19920,N_16113);
or UO_489 (O_489,N_17078,N_18861);
and UO_490 (O_490,N_17954,N_19672);
nor UO_491 (O_491,N_16107,N_17748);
xnor UO_492 (O_492,N_19565,N_16533);
or UO_493 (O_493,N_16110,N_19764);
or UO_494 (O_494,N_17426,N_18238);
nor UO_495 (O_495,N_17825,N_17846);
or UO_496 (O_496,N_19340,N_17442);
nor UO_497 (O_497,N_18740,N_18146);
nand UO_498 (O_498,N_17884,N_16035);
and UO_499 (O_499,N_16565,N_18372);
and UO_500 (O_500,N_18492,N_18519);
nor UO_501 (O_501,N_16887,N_18410);
nand UO_502 (O_502,N_16428,N_18452);
nor UO_503 (O_503,N_18508,N_19112);
nand UO_504 (O_504,N_16315,N_18723);
or UO_505 (O_505,N_17289,N_19074);
nor UO_506 (O_506,N_16500,N_19876);
or UO_507 (O_507,N_18640,N_17976);
nor UO_508 (O_508,N_17390,N_19707);
nor UO_509 (O_509,N_17013,N_18159);
nand UO_510 (O_510,N_16633,N_19613);
or UO_511 (O_511,N_17266,N_16810);
and UO_512 (O_512,N_17984,N_18050);
nand UO_513 (O_513,N_19275,N_16698);
nand UO_514 (O_514,N_19428,N_18682);
nand UO_515 (O_515,N_18119,N_19048);
or UO_516 (O_516,N_18938,N_17906);
and UO_517 (O_517,N_17056,N_18025);
nand UO_518 (O_518,N_17088,N_18369);
and UO_519 (O_519,N_17628,N_16914);
and UO_520 (O_520,N_18817,N_18677);
nand UO_521 (O_521,N_18560,N_16591);
and UO_522 (O_522,N_19768,N_16711);
nand UO_523 (O_523,N_19962,N_16712);
nand UO_524 (O_524,N_19215,N_18000);
xnor UO_525 (O_525,N_17313,N_16353);
and UO_526 (O_526,N_19996,N_16262);
and UO_527 (O_527,N_19154,N_16618);
or UO_528 (O_528,N_16517,N_17095);
and UO_529 (O_529,N_16824,N_16223);
nor UO_530 (O_530,N_19255,N_17383);
and UO_531 (O_531,N_16551,N_17359);
and UO_532 (O_532,N_18809,N_18930);
or UO_533 (O_533,N_19208,N_16773);
nand UO_534 (O_534,N_17066,N_17567);
nor UO_535 (O_535,N_16675,N_17565);
nand UO_536 (O_536,N_18818,N_16582);
and UO_537 (O_537,N_16478,N_16473);
nand UO_538 (O_538,N_16918,N_18465);
nand UO_539 (O_539,N_16403,N_18264);
nor UO_540 (O_540,N_17055,N_17929);
and UO_541 (O_541,N_19298,N_16908);
or UO_542 (O_542,N_16596,N_19599);
xor UO_543 (O_543,N_19607,N_19297);
xnor UO_544 (O_544,N_19829,N_16804);
nand UO_545 (O_545,N_17305,N_16800);
nor UO_546 (O_546,N_17090,N_19569);
xor UO_547 (O_547,N_18746,N_18421);
nor UO_548 (O_548,N_18769,N_16836);
and UO_549 (O_549,N_18293,N_18033);
xnor UO_550 (O_550,N_16409,N_18355);
nand UO_551 (O_551,N_17588,N_16285);
and UO_552 (O_552,N_19392,N_18302);
nand UO_553 (O_553,N_18348,N_16456);
xor UO_554 (O_554,N_18441,N_17234);
nor UO_555 (O_555,N_17721,N_16607);
or UO_556 (O_556,N_16893,N_17700);
nor UO_557 (O_557,N_19727,N_16273);
nor UO_558 (O_558,N_17038,N_19558);
or UO_559 (O_559,N_19326,N_17942);
nand UO_560 (O_560,N_16119,N_18806);
nand UO_561 (O_561,N_19577,N_16206);
xnor UO_562 (O_562,N_18163,N_16326);
nand UO_563 (O_563,N_17918,N_18375);
nand UO_564 (O_564,N_19594,N_16980);
or UO_565 (O_565,N_17735,N_17519);
or UO_566 (O_566,N_18317,N_17706);
nor UO_567 (O_567,N_19929,N_19176);
nand UO_568 (O_568,N_16574,N_16165);
or UO_569 (O_569,N_18991,N_19910);
or UO_570 (O_570,N_18748,N_17889);
nand UO_571 (O_571,N_16889,N_19139);
xnor UO_572 (O_572,N_16425,N_17583);
and UO_573 (O_573,N_18998,N_17804);
xor UO_574 (O_574,N_16118,N_17593);
xor UO_575 (O_575,N_17665,N_18982);
nand UO_576 (O_576,N_16770,N_16718);
xor UO_577 (O_577,N_16860,N_18956);
and UO_578 (O_578,N_17505,N_17510);
nand UO_579 (O_579,N_19938,N_19164);
xnor UO_580 (O_580,N_17467,N_17050);
nand UO_581 (O_581,N_18669,N_16553);
nor UO_582 (O_582,N_18753,N_16946);
and UO_583 (O_583,N_18713,N_17556);
or UO_584 (O_584,N_18778,N_18285);
nand UO_585 (O_585,N_16707,N_18189);
nand UO_586 (O_586,N_17867,N_17287);
and UO_587 (O_587,N_17947,N_17481);
or UO_588 (O_588,N_18850,N_17240);
xor UO_589 (O_589,N_19339,N_19970);
nor UO_590 (O_590,N_16881,N_19663);
and UO_591 (O_591,N_16029,N_19695);
xor UO_592 (O_592,N_18820,N_16622);
or UO_593 (O_593,N_19851,N_18070);
or UO_594 (O_594,N_16146,N_16581);
nor UO_595 (O_595,N_18579,N_18988);
or UO_596 (O_596,N_17232,N_16082);
and UO_597 (O_597,N_19677,N_19542);
and UO_598 (O_598,N_18409,N_18161);
xnor UO_599 (O_599,N_16978,N_19360);
nor UO_600 (O_600,N_17367,N_16798);
or UO_601 (O_601,N_19358,N_16211);
and UO_602 (O_602,N_16167,N_16308);
nand UO_603 (O_603,N_17156,N_18186);
nand UO_604 (O_604,N_19436,N_19348);
or UO_605 (O_605,N_16094,N_17536);
xnor UO_606 (O_606,N_17291,N_16895);
and UO_607 (O_607,N_18794,N_19748);
or UO_608 (O_608,N_19831,N_19616);
and UO_609 (O_609,N_16192,N_16919);
nand UO_610 (O_610,N_16126,N_19644);
nor UO_611 (O_611,N_17424,N_17032);
nor UO_612 (O_612,N_16886,N_17278);
nand UO_613 (O_613,N_16558,N_16322);
xor UO_614 (O_614,N_16575,N_19994);
nand UO_615 (O_615,N_16087,N_19804);
xnor UO_616 (O_616,N_18575,N_17474);
nand UO_617 (O_617,N_16859,N_19332);
xnor UO_618 (O_618,N_17429,N_19060);
or UO_619 (O_619,N_18183,N_17641);
nor UO_620 (O_620,N_18984,N_18539);
and UO_621 (O_621,N_19590,N_16961);
nor UO_622 (O_622,N_19337,N_16971);
nand UO_623 (O_623,N_19745,N_18570);
nand UO_624 (O_624,N_18164,N_17967);
or UO_625 (O_625,N_19615,N_17243);
nand UO_626 (O_626,N_16287,N_18107);
and UO_627 (O_627,N_16440,N_19083);
and UO_628 (O_628,N_18076,N_16399);
and UO_629 (O_629,N_16682,N_18843);
or UO_630 (O_630,N_18125,N_16270);
nor UO_631 (O_631,N_18035,N_19562);
xnor UO_632 (O_632,N_17497,N_17727);
or UO_633 (O_633,N_18028,N_17260);
and UO_634 (O_634,N_17786,N_16101);
nor UO_635 (O_635,N_18411,N_18336);
or UO_636 (O_636,N_18269,N_18925);
and UO_637 (O_637,N_16829,N_16977);
nor UO_638 (O_638,N_18096,N_16697);
and UO_639 (O_639,N_19162,N_16280);
and UO_640 (O_640,N_17596,N_19252);
nand UO_641 (O_641,N_19359,N_19361);
xnor UO_642 (O_642,N_18959,N_18540);
nand UO_643 (O_643,N_18395,N_17819);
or UO_644 (O_644,N_17948,N_17997);
nand UO_645 (O_645,N_19915,N_17769);
xor UO_646 (O_646,N_17448,N_19345);
and UO_647 (O_647,N_17115,N_16710);
nor UO_648 (O_648,N_18749,N_18622);
and UO_649 (O_649,N_17070,N_18807);
or UO_650 (O_650,N_18386,N_19809);
nand UO_651 (O_651,N_17403,N_16526);
and UO_652 (O_652,N_16984,N_19437);
nor UO_653 (O_653,N_18044,N_16955);
xnor UO_654 (O_654,N_16552,N_19926);
xor UO_655 (O_655,N_18828,N_19690);
or UO_656 (O_656,N_16694,N_19671);
xnor UO_657 (O_657,N_19794,N_18512);
and UO_658 (O_658,N_16833,N_16986);
xnor UO_659 (O_659,N_18630,N_17188);
or UO_660 (O_660,N_18650,N_19331);
and UO_661 (O_661,N_17625,N_17350);
nand UO_662 (O_662,N_18178,N_18432);
nand UO_663 (O_663,N_18535,N_16839);
or UO_664 (O_664,N_18516,N_16314);
nor UO_665 (O_665,N_19713,N_17590);
nor UO_666 (O_666,N_17127,N_18134);
nor UO_667 (O_667,N_18305,N_18248);
and UO_668 (O_668,N_19509,N_19367);
or UO_669 (O_669,N_18866,N_18056);
or UO_670 (O_670,N_18080,N_19133);
and UO_671 (O_671,N_19965,N_17956);
and UO_672 (O_672,N_17823,N_19788);
xnor UO_673 (O_673,N_18157,N_18542);
nor UO_674 (O_674,N_18761,N_19864);
nand UO_675 (O_675,N_16716,N_17150);
xnor UO_676 (O_676,N_19473,N_19014);
nand UO_677 (O_677,N_19008,N_18916);
nand UO_678 (O_678,N_16296,N_19219);
xor UO_679 (O_679,N_19916,N_18773);
nand UO_680 (O_680,N_19610,N_19209);
nand UO_681 (O_681,N_16342,N_17814);
and UO_682 (O_682,N_16597,N_18117);
or UO_683 (O_683,N_18577,N_19719);
nand UO_684 (O_684,N_19648,N_16725);
nand UO_685 (O_685,N_16657,N_17633);
or UO_686 (O_686,N_18731,N_16874);
nand UO_687 (O_687,N_19349,N_19443);
nand UO_688 (O_688,N_18442,N_19070);
and UO_689 (O_689,N_18053,N_16469);
or UO_690 (O_690,N_18656,N_19983);
nor UO_691 (O_691,N_19882,N_18052);
nor UO_692 (O_692,N_19853,N_18108);
or UO_693 (O_693,N_16735,N_18872);
nor UO_694 (O_694,N_16531,N_19296);
nand UO_695 (O_695,N_16143,N_18792);
and UO_696 (O_696,N_16964,N_17421);
or UO_697 (O_697,N_19403,N_18211);
nor UO_698 (O_698,N_17015,N_17173);
nor UO_699 (O_699,N_16757,N_17925);
nand UO_700 (O_700,N_19453,N_16079);
nand UO_701 (O_701,N_19379,N_19034);
or UO_702 (O_702,N_19637,N_18324);
or UO_703 (O_703,N_16982,N_19245);
or UO_704 (O_704,N_19790,N_17024);
nor UO_705 (O_705,N_17052,N_16095);
nand UO_706 (O_706,N_19664,N_19871);
or UO_707 (O_707,N_17432,N_18635);
nand UO_708 (O_708,N_19313,N_17649);
xnor UO_709 (O_709,N_19860,N_16032);
nor UO_710 (O_710,N_18497,N_18645);
and UO_711 (O_711,N_16402,N_17372);
nor UO_712 (O_712,N_17782,N_16147);
nor UO_713 (O_713,N_16255,N_17103);
nor UO_714 (O_714,N_19263,N_17355);
nor UO_715 (O_715,N_19614,N_17201);
nand UO_716 (O_716,N_18919,N_18711);
nand UO_717 (O_717,N_18785,N_18437);
and UO_718 (O_718,N_18971,N_16317);
and UO_719 (O_719,N_18876,N_17482);
and UO_720 (O_720,N_18662,N_19009);
or UO_721 (O_721,N_16911,N_18744);
xnor UO_722 (O_722,N_19750,N_17422);
or UO_723 (O_723,N_17713,N_18927);
or UO_724 (O_724,N_17902,N_17858);
or UO_725 (O_725,N_19494,N_19700);
nand UO_726 (O_726,N_16174,N_19696);
nor UO_727 (O_727,N_17286,N_18889);
nand UO_728 (O_728,N_16162,N_17362);
or UO_729 (O_729,N_16550,N_19560);
or UO_730 (O_730,N_17345,N_18297);
or UO_731 (O_731,N_18460,N_17116);
or UO_732 (O_732,N_19900,N_18330);
nor UO_733 (O_733,N_18139,N_17733);
xor UO_734 (O_734,N_19198,N_17731);
nor UO_735 (O_735,N_17302,N_16522);
or UO_736 (O_736,N_17676,N_19335);
nor UO_737 (O_737,N_16857,N_17087);
and UO_738 (O_738,N_16787,N_17368);
and UO_739 (O_739,N_18258,N_17992);
and UO_740 (O_740,N_16179,N_16205);
nand UO_741 (O_741,N_19278,N_19779);
nor UO_742 (O_742,N_16475,N_17927);
nor UO_743 (O_743,N_17888,N_19170);
nor UO_744 (O_744,N_18291,N_16883);
or UO_745 (O_745,N_17561,N_19870);
nor UO_746 (O_746,N_19184,N_17741);
nor UO_747 (O_747,N_18768,N_16846);
nand UO_748 (O_748,N_19863,N_18149);
or UO_749 (O_749,N_18265,N_16005);
or UO_750 (O_750,N_18162,N_18970);
xor UO_751 (O_751,N_18321,N_18709);
nor UO_752 (O_752,N_17502,N_17395);
nor UO_753 (O_753,N_18423,N_16514);
nand UO_754 (O_754,N_16071,N_16988);
nor UO_755 (O_755,N_16872,N_18244);
or UO_756 (O_756,N_19429,N_16683);
and UO_757 (O_757,N_16719,N_16614);
nand UO_758 (O_758,N_16068,N_17423);
and UO_759 (O_759,N_18058,N_19685);
nand UO_760 (O_760,N_17998,N_19229);
and UO_761 (O_761,N_17328,N_18929);
nand UO_762 (O_762,N_19730,N_19964);
or UO_763 (O_763,N_17250,N_18407);
and UO_764 (O_764,N_19218,N_16605);
nor UO_765 (O_765,N_18273,N_17450);
and UO_766 (O_766,N_18831,N_16080);
and UO_767 (O_767,N_18747,N_16902);
and UO_768 (O_768,N_17839,N_16181);
nor UO_769 (O_769,N_18086,N_19721);
and UO_770 (O_770,N_19175,N_19329);
and UO_771 (O_771,N_19488,N_16663);
nand UO_772 (O_772,N_18346,N_19847);
nor UO_773 (O_773,N_16778,N_19514);
and UO_774 (O_774,N_18770,N_16561);
xor UO_775 (O_775,N_19037,N_16823);
xnor UO_776 (O_776,N_19015,N_17479);
or UO_777 (O_777,N_17683,N_19445);
and UO_778 (O_778,N_18062,N_17663);
nor UO_779 (O_779,N_19046,N_17791);
xnor UO_780 (O_780,N_18931,N_16996);
nand UO_781 (O_781,N_17959,N_19984);
xor UO_782 (O_782,N_17891,N_16942);
nand UO_783 (O_783,N_17262,N_19204);
and UO_784 (O_784,N_19089,N_16486);
nor UO_785 (O_785,N_18067,N_18715);
nor UO_786 (O_786,N_18181,N_19087);
and UO_787 (O_787,N_16490,N_16416);
and UO_788 (O_788,N_18908,N_19927);
nor UO_789 (O_789,N_17543,N_16318);
and UO_790 (O_790,N_18132,N_18111);
and UO_791 (O_791,N_16349,N_19323);
and UO_792 (O_792,N_18079,N_16520);
nand UO_793 (O_793,N_17692,N_19236);
or UO_794 (O_794,N_19573,N_18124);
and UO_795 (O_795,N_18763,N_18308);
nor UO_796 (O_796,N_16257,N_18093);
nor UO_797 (O_797,N_17662,N_17828);
nand UO_798 (O_798,N_16256,N_16915);
nor UO_799 (O_799,N_18626,N_19288);
nand UO_800 (O_800,N_18739,N_16173);
or UO_801 (O_801,N_17194,N_19744);
xor UO_802 (O_802,N_18401,N_16813);
and UO_803 (O_803,N_16311,N_17028);
xnor UO_804 (O_804,N_19705,N_16802);
nor UO_805 (O_805,N_17310,N_16952);
xnor UO_806 (O_806,N_16122,N_18312);
and UO_807 (O_807,N_18193,N_17728);
xnor UO_808 (O_808,N_17939,N_17961);
nor UO_809 (O_809,N_17808,N_18520);
and UO_810 (O_810,N_18568,N_19312);
and UO_811 (O_811,N_19822,N_18810);
and UO_812 (O_812,N_16075,N_16554);
or UO_813 (O_813,N_17285,N_19773);
and UO_814 (O_814,N_19579,N_17936);
and UO_815 (O_815,N_18165,N_18027);
nand UO_816 (O_816,N_17719,N_19073);
or UO_817 (O_817,N_19369,N_17873);
nand UO_818 (O_818,N_19797,N_19571);
nor UO_819 (O_819,N_16284,N_18673);
nand UO_820 (O_820,N_18795,N_19385);
and UO_821 (O_821,N_17740,N_18422);
and UO_822 (O_822,N_18420,N_16620);
nand UO_823 (O_823,N_19441,N_19919);
nor UO_824 (O_824,N_18802,N_17311);
nand UO_825 (O_825,N_16251,N_17851);
or UO_826 (O_826,N_19631,N_19240);
and UO_827 (O_827,N_17710,N_19160);
nand UO_828 (O_828,N_17545,N_16927);
nor UO_829 (O_829,N_16258,N_18471);
nand UO_830 (O_830,N_17658,N_19409);
and UO_831 (O_831,N_16433,N_19466);
nand UO_832 (O_832,N_18620,N_19273);
and UO_833 (O_833,N_16750,N_17757);
and UO_834 (O_834,N_19444,N_19772);
and UO_835 (O_835,N_19305,N_19756);
and UO_836 (O_836,N_18553,N_19958);
and UO_837 (O_837,N_18322,N_18852);
or UO_838 (O_838,N_19961,N_18325);
and UO_839 (O_839,N_16221,N_16363);
nand UO_840 (O_840,N_19899,N_18864);
xor UO_841 (O_841,N_19493,N_16634);
nand UO_842 (O_842,N_17433,N_16629);
and UO_843 (O_843,N_18924,N_16189);
or UO_844 (O_844,N_19905,N_17296);
xnor UO_845 (O_845,N_19729,N_16630);
nor UO_846 (O_846,N_16882,N_17743);
and UO_847 (O_847,N_17732,N_16659);
nand UO_848 (O_848,N_16306,N_17680);
nor UO_849 (O_849,N_18156,N_19835);
nand UO_850 (O_850,N_16264,N_17870);
nor UO_851 (O_851,N_16852,N_19992);
nor UO_852 (O_852,N_16420,N_16350);
or UO_853 (O_853,N_16129,N_19706);
nand UO_854 (O_854,N_17594,N_16623);
nand UO_855 (O_855,N_19867,N_16556);
nand UO_856 (O_856,N_19010,N_17511);
nand UO_857 (O_857,N_19714,N_18085);
nor UO_858 (O_858,N_19525,N_17393);
and UO_859 (O_859,N_19376,N_18359);
and UO_860 (O_860,N_19268,N_19803);
and UO_861 (O_861,N_16818,N_18333);
or UO_862 (O_862,N_17551,N_16831);
and UO_863 (O_863,N_18091,N_18450);
xnor UO_864 (O_864,N_16364,N_19148);
and UO_865 (O_865,N_16523,N_19226);
nor UO_866 (O_866,N_16834,N_17411);
nor UO_867 (O_867,N_19179,N_16340);
and UO_868 (O_868,N_19018,N_17830);
nand UO_869 (O_869,N_17553,N_18222);
nor UO_870 (O_870,N_17151,N_18243);
and UO_871 (O_871,N_16567,N_16418);
and UO_872 (O_872,N_17330,N_19024);
or UO_873 (O_873,N_19368,N_19039);
and UO_874 (O_874,N_17205,N_19489);
and UO_875 (O_875,N_17604,N_19665);
nor UO_876 (O_876,N_17363,N_19762);
nor UO_877 (O_877,N_19138,N_18081);
nor UO_878 (O_878,N_18547,N_19063);
nor UO_879 (O_879,N_16413,N_16172);
or UO_880 (O_880,N_16235,N_18213);
or UO_881 (O_881,N_16465,N_19328);
or UO_882 (O_882,N_18784,N_17097);
or UO_883 (O_883,N_17994,N_16177);
nor UO_884 (O_884,N_16215,N_16608);
and UO_885 (O_885,N_16653,N_16692);
or UO_886 (O_886,N_17624,N_16444);
nor UO_887 (O_887,N_18804,N_19528);
xnor UO_888 (O_888,N_17563,N_18169);
nand UO_889 (O_889,N_18252,N_18997);
nor UO_890 (O_890,N_19572,N_17540);
nor UO_891 (O_891,N_18913,N_17297);
nor UO_892 (O_892,N_17987,N_18664);
nor UO_893 (O_893,N_19320,N_16783);
or UO_894 (O_894,N_19879,N_18838);
and UO_895 (O_895,N_19482,N_17838);
or UO_896 (O_896,N_19999,N_16661);
nor UO_897 (O_897,N_17370,N_16457);
and UO_898 (O_898,N_16245,N_18858);
and UO_899 (O_899,N_19080,N_16109);
or UO_900 (O_900,N_19396,N_18400);
nand UO_901 (O_901,N_17183,N_18065);
nor UO_902 (O_902,N_16238,N_17161);
or UO_903 (O_903,N_16157,N_19889);
or UO_904 (O_904,N_17574,N_16515);
and UO_905 (O_905,N_18428,N_17269);
or UO_906 (O_906,N_19817,N_18880);
and UO_907 (O_907,N_17229,N_19079);
or UO_908 (O_908,N_18268,N_18584);
xor UO_909 (O_909,N_18112,N_16385);
or UO_910 (O_910,N_18522,N_19391);
xor UO_911 (O_911,N_18708,N_16599);
and UO_912 (O_912,N_17181,N_17811);
nor UO_913 (O_913,N_17455,N_18911);
or UO_914 (O_914,N_16812,N_17775);
nand UO_915 (O_915,N_18408,N_16684);
nand UO_916 (O_916,N_16389,N_17795);
and UO_917 (O_917,N_17711,N_16057);
xnor UO_918 (O_918,N_18431,N_16641);
and UO_919 (O_919,N_16070,N_19407);
nor UO_920 (O_920,N_18538,N_18615);
nand UO_921 (O_921,N_18168,N_17040);
nand UO_922 (O_922,N_16512,N_19894);
nand UO_923 (O_923,N_19020,N_18077);
nor UO_924 (O_924,N_19807,N_18976);
nor UO_925 (O_925,N_18314,N_16464);
nand UO_926 (O_926,N_18738,N_18227);
and UO_927 (O_927,N_18484,N_19017);
and UO_928 (O_928,N_18357,N_17919);
nand UO_929 (O_929,N_17661,N_17524);
or UO_930 (O_930,N_17208,N_16625);
xor UO_931 (O_931,N_16466,N_19315);
nand UO_932 (O_932,N_18133,N_16357);
or UO_933 (O_933,N_16376,N_18955);
nand UO_934 (O_934,N_18381,N_18031);
or UO_935 (O_935,N_18593,N_19137);
nor UO_936 (O_936,N_16356,N_19082);
and UO_937 (O_937,N_18846,N_16903);
or UO_938 (O_938,N_17859,N_17020);
and UO_939 (O_939,N_17903,N_19210);
and UO_940 (O_940,N_16483,N_18364);
and UO_941 (O_941,N_17887,N_18777);
and UO_942 (O_942,N_18083,N_17558);
and UO_943 (O_943,N_18525,N_16210);
and UO_944 (O_944,N_18283,N_16383);
nand UO_945 (O_945,N_19734,N_17165);
nor UO_946 (O_946,N_17155,N_19130);
or UO_947 (O_947,N_18066,N_18217);
or UO_948 (O_948,N_19067,N_18396);
nor UO_949 (O_949,N_18467,N_19732);
nand UO_950 (O_950,N_18878,N_18826);
and UO_951 (O_951,N_19325,N_16822);
nand UO_952 (O_952,N_18261,N_18341);
nor UO_953 (O_953,N_17657,N_17177);
xnor UO_954 (O_954,N_18234,N_19643);
and UO_955 (O_955,N_17071,N_18871);
nand UO_956 (O_956,N_17790,N_18660);
xor UO_957 (O_957,N_17785,N_17427);
or UO_958 (O_958,N_19963,N_18382);
or UO_959 (O_959,N_16199,N_19426);
nor UO_960 (O_960,N_19923,N_19397);
nand UO_961 (O_961,N_16153,N_18137);
nor UO_962 (O_962,N_16305,N_19640);
and UO_963 (O_963,N_18469,N_18690);
nor UO_964 (O_964,N_19784,N_18782);
or UO_965 (O_965,N_18932,N_17255);
nand UO_966 (O_966,N_16826,N_18378);
or UO_967 (O_967,N_16304,N_18173);
nand UO_968 (O_968,N_18564,N_16862);
xnor UO_969 (O_969,N_18433,N_19260);
and UO_970 (O_970,N_16954,N_16207);
nand UO_971 (O_971,N_18781,N_17319);
nor UO_972 (O_972,N_17365,N_16025);
nand UO_973 (O_973,N_19214,N_17430);
nor UO_974 (O_974,N_17802,N_17224);
or UO_975 (O_975,N_16053,N_18741);
xnor UO_976 (O_976,N_17158,N_18072);
nor UO_977 (O_977,N_18127,N_17157);
xnor UO_978 (O_978,N_17490,N_16400);
or UO_979 (O_979,N_16202,N_18756);
and UO_980 (O_980,N_18905,N_19971);
and UO_981 (O_981,N_17974,N_19632);
nand UO_982 (O_982,N_16600,N_18710);
or UO_983 (O_983,N_16586,N_18591);
and UO_984 (O_984,N_19119,N_17471);
nand UO_985 (O_985,N_16131,N_18604);
and UO_986 (O_986,N_17060,N_19521);
nor UO_987 (O_987,N_19221,N_19953);
and UO_988 (O_988,N_17271,N_16589);
nand UO_989 (O_989,N_16169,N_16835);
nand UO_990 (O_990,N_18326,N_18301);
xor UO_991 (O_991,N_16728,N_19943);
nor UO_992 (O_992,N_19789,N_18815);
nand UO_993 (O_993,N_19134,N_18279);
and UO_994 (O_994,N_19042,N_18029);
and UO_995 (O_995,N_19936,N_16487);
nor UO_996 (O_996,N_18440,N_16921);
or UO_997 (O_997,N_16930,N_18638);
xnor UO_998 (O_998,N_18235,N_19456);
nand UO_999 (O_999,N_18701,N_17003);
xor UO_1000 (O_1000,N_18122,N_18655);
and UO_1001 (O_1001,N_19654,N_18563);
or UO_1002 (O_1002,N_16726,N_17128);
nand UO_1003 (O_1003,N_17488,N_18047);
or UO_1004 (O_1004,N_18218,N_19051);
xnor UO_1005 (O_1005,N_16858,N_16231);
nor UO_1006 (O_1006,N_19948,N_19206);
and UO_1007 (O_1007,N_16442,N_18311);
nand UO_1008 (O_1008,N_16330,N_16948);
and UO_1009 (O_1009,N_16291,N_17877);
and UO_1010 (O_1010,N_17977,N_19344);
or UO_1011 (O_1011,N_16139,N_16193);
nor UO_1012 (O_1012,N_16809,N_19701);
nor UO_1013 (O_1013,N_17321,N_18589);
and UO_1014 (O_1014,N_19510,N_16060);
nand UO_1015 (O_1015,N_17538,N_16431);
nand UO_1016 (O_1016,N_18207,N_18745);
or UO_1017 (O_1017,N_18957,N_17206);
and UO_1018 (O_1018,N_17631,N_16237);
and UO_1019 (O_1019,N_19088,N_19192);
nand UO_1020 (O_1020,N_16406,N_18074);
nor UO_1021 (O_1021,N_19469,N_17639);
and UO_1022 (O_1022,N_16507,N_17579);
xnor UO_1023 (O_1023,N_18835,N_16452);
or UO_1024 (O_1024,N_18842,N_19739);
nor UO_1025 (O_1025,N_18256,N_17244);
xnor UO_1026 (O_1026,N_19875,N_19907);
xnor UO_1027 (O_1027,N_16875,N_18059);
nand UO_1028 (O_1028,N_16377,N_16580);
nor UO_1029 (O_1029,N_17029,N_18435);
nor UO_1030 (O_1030,N_17492,N_16121);
xor UO_1031 (O_1031,N_17619,N_16410);
and UO_1032 (O_1032,N_17146,N_17626);
nor UO_1033 (O_1033,N_17037,N_18917);
and UO_1034 (O_1034,N_17136,N_16944);
and UO_1035 (O_1035,N_17164,N_16178);
nand UO_1036 (O_1036,N_16910,N_17926);
and UO_1037 (O_1037,N_18404,N_19125);
xor UO_1038 (O_1038,N_19306,N_17027);
nor UO_1039 (O_1039,N_17222,N_19704);
nor UO_1040 (O_1040,N_17456,N_19760);
or UO_1041 (O_1041,N_16979,N_19551);
and UO_1042 (O_1042,N_16117,N_18128);
and UO_1043 (O_1043,N_18712,N_18130);
nor UO_1044 (O_1044,N_17154,N_18415);
or UO_1045 (O_1045,N_16197,N_18798);
and UO_1046 (O_1046,N_17284,N_16039);
or UO_1047 (O_1047,N_19012,N_16624);
xor UO_1048 (O_1048,N_16843,N_17636);
nand UO_1049 (O_1049,N_18131,N_19230);
nor UO_1050 (O_1050,N_18623,N_18209);
and UO_1051 (O_1051,N_19434,N_17688);
nor UO_1052 (O_1052,N_19071,N_18718);
nor UO_1053 (O_1053,N_19969,N_18129);
nor UO_1054 (O_1054,N_17568,N_18611);
nor UO_1055 (O_1055,N_19188,N_19662);
and UO_1056 (O_1056,N_16227,N_17729);
nor UO_1057 (O_1057,N_18634,N_16144);
nor UO_1058 (O_1058,N_19697,N_16538);
xor UO_1059 (O_1059,N_18007,N_16931);
and UO_1060 (O_1060,N_18765,N_16495);
or UO_1061 (O_1061,N_17476,N_18764);
nand UO_1062 (O_1062,N_17343,N_17542);
or UO_1063 (O_1063,N_18345,N_16974);
or UO_1064 (O_1064,N_17152,N_18477);
nor UO_1065 (O_1065,N_19314,N_17107);
and UO_1066 (O_1066,N_18390,N_17203);
nand UO_1067 (O_1067,N_16116,N_19620);
or UO_1068 (O_1068,N_19698,N_17801);
and UO_1069 (O_1069,N_19646,N_17951);
nor UO_1070 (O_1070,N_18337,N_16869);
nor UO_1071 (O_1071,N_16969,N_17253);
or UO_1072 (O_1072,N_18910,N_17564);
nor UO_1073 (O_1073,N_18487,N_16775);
nand UO_1074 (O_1074,N_19786,N_16938);
nor UO_1075 (O_1075,N_16152,N_17186);
nand UO_1076 (O_1076,N_18413,N_18639);
nor UO_1077 (O_1077,N_16477,N_18595);
or UO_1078 (O_1078,N_19290,N_19124);
and UO_1079 (O_1079,N_19712,N_17650);
nor UO_1080 (O_1080,N_18999,N_17200);
or UO_1081 (O_1081,N_19904,N_16388);
or UO_1082 (O_1082,N_16746,N_19189);
nand UO_1083 (O_1083,N_19580,N_17170);
or UO_1084 (O_1084,N_18863,N_17507);
nor UO_1085 (O_1085,N_17276,N_16744);
or UO_1086 (O_1086,N_19869,N_17242);
xnor UO_1087 (O_1087,N_19065,N_17396);
nand UO_1088 (O_1088,N_17644,N_18281);
nand UO_1089 (O_1089,N_19304,N_17600);
nand UO_1090 (O_1090,N_19374,N_16799);
and UO_1091 (O_1091,N_19898,N_16347);
or UO_1092 (O_1092,N_16017,N_19468);
and UO_1093 (O_1093,N_18952,N_19269);
or UO_1094 (O_1094,N_16527,N_16786);
and UO_1095 (O_1095,N_17016,N_16913);
and UO_1096 (O_1096,N_18569,N_18566);
nor UO_1097 (O_1097,N_16513,N_18609);
nand UO_1098 (O_1098,N_18772,N_17508);
nor UO_1099 (O_1099,N_19249,N_16447);
or UO_1100 (O_1100,N_16925,N_17980);
nand UO_1101 (O_1101,N_18141,N_18329);
nand UO_1102 (O_1102,N_16516,N_19816);
or UO_1103 (O_1103,N_16319,N_17864);
xnor UO_1104 (O_1104,N_17668,N_17666);
or UO_1105 (O_1105,N_19924,N_16870);
nor UO_1106 (O_1106,N_17048,N_16266);
nor UO_1107 (O_1107,N_17609,N_18675);
or UO_1108 (O_1108,N_18856,N_18691);
nand UO_1109 (O_1109,N_19543,N_18942);
xnor UO_1110 (O_1110,N_17749,N_16134);
and UO_1111 (O_1111,N_17988,N_16606);
nor UO_1112 (O_1112,N_18502,N_16576);
or UO_1113 (O_1113,N_18613,N_17329);
and UO_1114 (O_1114,N_19861,N_17854);
and UO_1115 (O_1115,N_18366,N_19639);
and UO_1116 (O_1116,N_17962,N_17041);
nor UO_1117 (O_1117,N_17349,N_16359);
or UO_1118 (O_1118,N_18821,N_16705);
and UO_1119 (O_1119,N_18642,N_18102);
and UO_1120 (O_1120,N_17720,N_19155);
nor UO_1121 (O_1121,N_17130,N_19596);
nor UO_1122 (O_1122,N_17645,N_16647);
or UO_1123 (O_1123,N_17354,N_19295);
nand UO_1124 (O_1124,N_18813,N_19586);
or UO_1125 (O_1125,N_16013,N_16230);
nand UO_1126 (O_1126,N_18659,N_16639);
and UO_1127 (O_1127,N_17970,N_17965);
nand UO_1128 (O_1128,N_18347,N_18990);
nand UO_1129 (O_1129,N_18021,N_17281);
or UO_1130 (O_1130,N_19064,N_19069);
nor UO_1131 (O_1131,N_16229,N_18819);
or UO_1132 (O_1132,N_18094,N_16939);
nand UO_1133 (O_1133,N_17818,N_16703);
nor UO_1134 (O_1134,N_19425,N_19450);
and UO_1135 (O_1135,N_17702,N_16615);
and UO_1136 (O_1136,N_16168,N_18262);
and UO_1137 (O_1137,N_17121,N_18506);
nand UO_1138 (O_1138,N_18837,N_17316);
nor UO_1139 (O_1139,N_18771,N_18903);
or UO_1140 (O_1140,N_16142,N_17026);
xor UO_1141 (O_1141,N_19832,N_19885);
or UO_1142 (O_1142,N_18318,N_19800);
xnor UO_1143 (O_1143,N_19174,N_19438);
nand UO_1144 (O_1144,N_18588,N_18481);
or UO_1145 (O_1145,N_16853,N_19225);
or UO_1146 (O_1146,N_18152,N_17897);
and UO_1147 (O_1147,N_17592,N_16127);
or UO_1148 (O_1148,N_17384,N_19777);
nor UO_1149 (O_1149,N_16956,N_18684);
nor UO_1150 (O_1150,N_16498,N_16612);
nor UO_1151 (O_1151,N_19922,N_17844);
and UO_1152 (O_1152,N_18543,N_19995);
or UO_1153 (O_1153,N_17231,N_16112);
or UO_1154 (O_1154,N_19006,N_16861);
nand UO_1155 (O_1155,N_19246,N_18537);
xor UO_1156 (O_1156,N_19159,N_17292);
nand UO_1157 (O_1157,N_19180,N_16509);
nand UO_1158 (O_1158,N_16375,N_16819);
nand UO_1159 (O_1159,N_18054,N_18926);
and UO_1160 (O_1160,N_16832,N_19848);
nor UO_1161 (O_1161,N_19244,N_18759);
or UO_1162 (O_1162,N_16868,N_19799);
nand UO_1163 (O_1163,N_17460,N_16392);
or UO_1164 (O_1164,N_19749,N_16617);
and UO_1165 (O_1165,N_19217,N_19053);
or UO_1166 (O_1166,N_19380,N_19460);
nand UO_1167 (O_1167,N_18016,N_19629);
nand UO_1168 (O_1168,N_16213,N_16055);
nor UO_1169 (O_1169,N_18104,N_16051);
nand UO_1170 (O_1170,N_19050,N_16796);
and UO_1171 (O_1171,N_19592,N_17763);
nor UO_1172 (O_1172,N_19276,N_16736);
nor UO_1173 (O_1173,N_17277,N_16275);
and UO_1174 (O_1174,N_17577,N_17653);
and UO_1175 (O_1175,N_18674,N_19442);
or UO_1176 (O_1176,N_18034,N_19181);
nand UO_1177 (O_1177,N_18572,N_17135);
nand UO_1178 (O_1178,N_16541,N_17584);
nor UO_1179 (O_1179,N_19780,N_18972);
and UO_1180 (O_1180,N_17685,N_17879);
xnor UO_1181 (O_1181,N_17445,N_17820);
and UO_1182 (O_1182,N_16828,N_16058);
xnor UO_1183 (O_1183,N_18912,N_18199);
nor UO_1184 (O_1184,N_19930,N_19827);
and UO_1185 (O_1185,N_19836,N_19845);
or UO_1186 (O_1186,N_17030,N_19538);
nand UO_1187 (O_1187,N_19194,N_19142);
or UO_1188 (O_1188,N_19531,N_17678);
nand UO_1189 (O_1189,N_17548,N_18443);
nand UO_1190 (O_1190,N_18775,N_18867);
nand UO_1191 (O_1191,N_18208,N_18518);
or UO_1192 (O_1192,N_17185,N_16686);
and UO_1193 (O_1193,N_18896,N_16626);
or UO_1194 (O_1194,N_17413,N_18109);
xor UO_1195 (O_1195,N_18592,N_19702);
and UO_1196 (O_1196,N_17199,N_18987);
xor UO_1197 (O_1197,N_18546,N_18242);
or UO_1198 (O_1198,N_16570,N_19954);
nor UO_1199 (O_1199,N_18294,N_16610);
or UO_1200 (O_1200,N_17247,N_18118);
nand UO_1201 (O_1201,N_18223,N_19854);
nand UO_1202 (O_1202,N_18503,N_18192);
or UO_1203 (O_1203,N_16078,N_16549);
nor UO_1204 (O_1204,N_18757,N_18549);
nand UO_1205 (O_1205,N_19680,N_16265);
and UO_1206 (O_1206,N_17010,N_16367);
nand UO_1207 (O_1207,N_19378,N_19262);
nand UO_1208 (O_1208,N_19476,N_19937);
nand UO_1209 (O_1209,N_18344,N_18340);
nor UO_1210 (O_1210,N_17122,N_17477);
nor UO_1211 (O_1211,N_17025,N_17175);
nor UO_1212 (O_1212,N_19222,N_19891);
nor UO_1213 (O_1213,N_17051,N_19381);
or UO_1214 (O_1214,N_19478,N_18884);
or UO_1215 (O_1215,N_17783,N_17913);
or UO_1216 (O_1216,N_19104,N_17098);
and UO_1217 (O_1217,N_18933,N_17516);
nand UO_1218 (O_1218,N_16345,N_19921);
and UO_1219 (O_1219,N_18009,N_18796);
nor UO_1220 (O_1220,N_18565,N_16987);
and UO_1221 (O_1221,N_18590,N_19645);
nor UO_1222 (O_1222,N_18729,N_16560);
nor UO_1223 (O_1223,N_17754,N_16780);
and UO_1224 (O_1224,N_16863,N_19949);
and UO_1225 (O_1225,N_18384,N_17143);
xor UO_1226 (O_1226,N_16776,N_19518);
or UO_1227 (O_1227,N_16609,N_17973);
nand UO_1228 (O_1228,N_16088,N_17279);
nand UO_1229 (O_1229,N_17228,N_19759);
xnor UO_1230 (O_1230,N_19173,N_17458);
nor UO_1231 (O_1231,N_16042,N_17630);
nor UO_1232 (O_1232,N_16102,N_17248);
nand UO_1233 (O_1233,N_17539,N_18949);
nand UO_1234 (O_1234,N_16277,N_19408);
or UO_1235 (O_1235,N_18824,N_16548);
and UO_1236 (O_1236,N_16355,N_19873);
nor UO_1237 (O_1237,N_17438,N_17469);
nor UO_1238 (O_1238,N_18841,N_16662);
nor UO_1239 (O_1239,N_17881,N_19318);
xor UO_1240 (O_1240,N_16936,N_17571);
nand UO_1241 (O_1241,N_16949,N_16407);
nand UO_1242 (O_1242,N_16923,N_17787);
xor UO_1243 (O_1243,N_18985,N_18255);
nand UO_1244 (O_1244,N_16759,N_17133);
and UO_1245 (O_1245,N_16114,N_17898);
or UO_1246 (O_1246,N_18339,N_19545);
nand UO_1247 (O_1247,N_18941,N_19823);
nor UO_1248 (O_1248,N_18928,N_16985);
nand UO_1249 (O_1249,N_19271,N_17768);
or UO_1250 (O_1250,N_16901,N_18174);
nor UO_1251 (O_1251,N_19681,N_16510);
xnor UO_1252 (O_1252,N_16602,N_19195);
and UO_1253 (O_1253,N_16467,N_17100);
nand UO_1254 (O_1254,N_16953,N_17404);
or UO_1255 (O_1255,N_17408,N_16346);
and UO_1256 (O_1256,N_19019,N_18166);
or UO_1257 (O_1257,N_18418,N_17360);
nor UO_1258 (O_1258,N_19715,N_19098);
nand UO_1259 (O_1259,N_17342,N_18048);
and UO_1260 (O_1260,N_18587,N_17826);
and UO_1261 (O_1261,N_17079,N_17522);
nor UO_1262 (O_1262,N_17314,N_18092);
and UO_1263 (O_1263,N_17744,N_17682);
nand UO_1264 (O_1264,N_18397,N_16293);
nor UO_1265 (O_1265,N_17077,N_19767);
nor UO_1266 (O_1266,N_19642,N_16085);
nand UO_1267 (O_1267,N_18694,N_18891);
nand UO_1268 (O_1268,N_17213,N_19726);
nor UO_1269 (O_1269,N_18693,N_16393);
nand UO_1270 (O_1270,N_18099,N_17125);
nand UO_1271 (O_1271,N_18376,N_16271);
nand UO_1272 (O_1272,N_16730,N_16438);
or UO_1273 (O_1273,N_18121,N_16426);
nand UO_1274 (O_1274,N_17282,N_18352);
nor UO_1275 (O_1275,N_19941,N_17591);
nand UO_1276 (O_1276,N_19118,N_17333);
nand UO_1277 (O_1277,N_16204,N_16158);
xnor UO_1278 (O_1278,N_17261,N_19686);
or UO_1279 (O_1279,N_19897,N_18879);
nor UO_1280 (O_1280,N_16052,N_17004);
or UO_1281 (O_1281,N_19737,N_17256);
nor UO_1282 (O_1282,N_18524,N_19451);
nand UO_1283 (O_1283,N_19231,N_17623);
nor UO_1284 (O_1284,N_18008,N_17894);
or UO_1285 (O_1285,N_19414,N_16148);
xor UO_1286 (O_1286,N_19190,N_19011);
nor UO_1287 (O_1287,N_17765,N_19202);
nor UO_1288 (O_1288,N_18026,N_19455);
and UO_1289 (O_1289,N_16098,N_17957);
nor UO_1290 (O_1290,N_19462,N_16298);
xnor UO_1291 (O_1291,N_19945,N_16502);
nand UO_1292 (O_1292,N_19793,N_18528);
or UO_1293 (O_1293,N_16595,N_18666);
nor UO_1294 (O_1294,N_17388,N_16795);
nor UO_1295 (O_1295,N_18545,N_17578);
nand UO_1296 (O_1296,N_17084,N_19649);
and UO_1297 (O_1297,N_17559,N_17209);
and UO_1298 (O_1298,N_19241,N_17400);
or UO_1299 (O_1299,N_18373,N_18474);
nand UO_1300 (O_1300,N_18225,N_16047);
or UO_1301 (O_1301,N_19931,N_19057);
xnor UO_1302 (O_1302,N_17171,N_18724);
nor UO_1303 (O_1303,N_19993,N_16555);
nand UO_1304 (O_1304,N_16195,N_19193);
or UO_1305 (O_1305,N_19753,N_18457);
nor UO_1306 (O_1306,N_16503,N_19912);
nor UO_1307 (O_1307,N_18039,N_16866);
nand UO_1308 (O_1308,N_18619,N_19626);
or UO_1309 (O_1309,N_17402,N_19211);
xor UO_1310 (O_1310,N_18598,N_19086);
nor UO_1311 (O_1311,N_19940,N_16933);
or UO_1312 (O_1312,N_18182,N_17011);
nand UO_1313 (O_1313,N_19883,N_18361);
nor UO_1314 (O_1314,N_16535,N_16563);
and UO_1315 (O_1315,N_17529,N_17299);
and UO_1316 (O_1316,N_17923,N_19887);
nand UO_1317 (O_1317,N_19634,N_16247);
or UO_1318 (O_1318,N_19711,N_19588);
and UO_1319 (O_1319,N_19550,N_17465);
nor UO_1320 (O_1320,N_16761,N_19007);
and UO_1321 (O_1321,N_18491,N_16524);
nand UO_1322 (O_1322,N_17852,N_16590);
nor UO_1323 (O_1323,N_17969,N_16679);
nor UO_1324 (O_1324,N_17021,N_16840);
nand UO_1325 (O_1325,N_19487,N_18089);
nand UO_1326 (O_1326,N_18385,N_17674);
nor UO_1327 (O_1327,N_18270,N_17064);
nor UO_1328 (O_1328,N_17444,N_19716);
and UO_1329 (O_1329,N_16449,N_19597);
nand UO_1330 (O_1330,N_17863,N_17220);
nor UO_1331 (O_1331,N_19892,N_16268);
xor UO_1332 (O_1332,N_19679,N_19025);
nor UO_1333 (O_1333,N_18365,N_16140);
or UO_1334 (O_1334,N_18343,N_16673);
nand UO_1335 (O_1335,N_17821,N_19669);
nand UO_1336 (O_1336,N_17275,N_18399);
or UO_1337 (O_1337,N_16603,N_18479);
nor UO_1338 (O_1338,N_18730,N_16766);
nor UO_1339 (O_1339,N_19859,N_18851);
nand UO_1340 (O_1340,N_16272,N_19746);
and UO_1341 (O_1341,N_16966,N_16890);
and UO_1342 (O_1342,N_18263,N_17172);
xnor UO_1343 (O_1343,N_16203,N_18456);
nand UO_1344 (O_1344,N_18286,N_19136);
or UO_1345 (O_1345,N_16358,N_17606);
xor UO_1346 (O_1346,N_16022,N_16756);
or UO_1347 (O_1347,N_19243,N_16233);
or UO_1348 (O_1348,N_19622,N_16519);
nand UO_1349 (O_1349,N_19589,N_18953);
or UO_1350 (O_1350,N_18023,N_19508);
or UO_1351 (O_1351,N_19881,N_17245);
or UO_1352 (O_1352,N_19709,N_16848);
and UO_1353 (O_1353,N_18398,N_16760);
or UO_1354 (O_1354,N_16983,N_18071);
and UO_1355 (O_1355,N_19417,N_19365);
nor UO_1356 (O_1356,N_18969,N_19371);
and UO_1357 (O_1357,N_18219,N_16239);
and UO_1358 (O_1358,N_19395,N_16880);
and UO_1359 (O_1359,N_16917,N_18742);
and UO_1360 (O_1360,N_19281,N_19484);
nand UO_1361 (O_1361,N_17921,N_17327);
nand UO_1362 (O_1362,N_18191,N_17124);
xnor UO_1363 (O_1363,N_19470,N_16648);
or UO_1364 (O_1364,N_16062,N_17086);
or UO_1365 (O_1365,N_16871,N_16667);
and UO_1366 (O_1366,N_18719,N_16763);
xnor UO_1367 (O_1367,N_18811,N_18298);
nand UO_1368 (O_1368,N_19828,N_16849);
nand UO_1369 (O_1369,N_18663,N_16043);
nor UO_1370 (O_1370,N_17263,N_17533);
nand UO_1371 (O_1371,N_18020,N_19856);
or UO_1372 (O_1372,N_16557,N_19977);
and UO_1373 (O_1373,N_16015,N_19890);
or UO_1374 (O_1374,N_18103,N_17767);
nand UO_1375 (O_1375,N_18562,N_19223);
nor UO_1376 (O_1376,N_16781,N_17570);
or UO_1377 (O_1377,N_18391,N_18040);
xor UO_1378 (O_1378,N_17528,N_17069);
or UO_1379 (O_1379,N_18644,N_19604);
nor UO_1380 (O_1380,N_18943,N_18254);
or UO_1381 (O_1381,N_17451,N_19635);
and UO_1382 (O_1382,N_19658,N_18490);
xnor UO_1383 (O_1383,N_16136,N_16743);
or UO_1384 (O_1384,N_16530,N_17853);
and UO_1385 (O_1385,N_17377,N_17788);
and UO_1386 (O_1386,N_18882,N_16842);
or UO_1387 (O_1387,N_19459,N_17226);
xnor UO_1388 (O_1388,N_19840,N_18608);
nor UO_1389 (O_1389,N_17655,N_18195);
and UO_1390 (O_1390,N_18541,N_16212);
nand UO_1391 (O_1391,N_18438,N_16713);
nor UO_1392 (O_1392,N_19235,N_19552);
xor UO_1393 (O_1393,N_18051,N_17195);
or UO_1394 (O_1394,N_19502,N_17679);
and UO_1395 (O_1395,N_17374,N_18320);
nand UO_1396 (O_1396,N_17857,N_19474);
nand UO_1397 (O_1397,N_16856,N_18963);
and UO_1398 (O_1398,N_19952,N_18170);
nor UO_1399 (O_1399,N_18667,N_19947);
nand UO_1400 (O_1400,N_19427,N_16740);
or UO_1401 (O_1401,N_16294,N_18865);
and UO_1402 (O_1402,N_19149,N_17498);
or UO_1403 (O_1403,N_16714,N_18706);
or UO_1404 (O_1404,N_19914,N_17392);
nor UO_1405 (O_1405,N_16011,N_19171);
nor UO_1406 (O_1406,N_18973,N_17187);
nor UO_1407 (O_1407,N_16463,N_18979);
xnor UO_1408 (O_1408,N_17068,N_18523);
nand UO_1409 (O_1409,N_19988,N_18276);
and UO_1410 (O_1410,N_18529,N_17509);
or UO_1411 (O_1411,N_18205,N_17715);
and UO_1412 (O_1412,N_19109,N_16628);
xor UO_1413 (O_1413,N_16435,N_19998);
or UO_1414 (O_1414,N_16344,N_17696);
or UO_1415 (O_1415,N_18658,N_16361);
or UO_1416 (O_1416,N_16894,N_18240);
and UO_1417 (O_1417,N_16044,N_16729);
nor UO_1418 (O_1418,N_17912,N_16405);
xor UO_1419 (O_1419,N_19850,N_17101);
or UO_1420 (O_1420,N_16279,N_19957);
or UO_1421 (O_1421,N_17531,N_17557);
or UO_1422 (O_1422,N_17807,N_18323);
nor UO_1423 (O_1423,N_18707,N_16321);
or UO_1424 (O_1424,N_19743,N_19731);
xor UO_1425 (O_1425,N_17739,N_18977);
nand UO_1426 (O_1426,N_17132,N_17083);
and UO_1427 (O_1427,N_17848,N_16631);
or UO_1428 (O_1428,N_16791,N_19523);
and UO_1429 (O_1429,N_17996,N_19496);
or UO_1430 (O_1430,N_17501,N_17120);
and UO_1431 (O_1431,N_19077,N_17953);
and UO_1432 (O_1432,N_17366,N_18980);
and UO_1433 (O_1433,N_17871,N_17985);
and UO_1434 (O_1434,N_17589,N_19058);
nand UO_1435 (O_1435,N_18624,N_18327);
or UO_1436 (O_1436,N_19274,N_18393);
nand UO_1437 (O_1437,N_17357,N_17751);
xnor UO_1438 (O_1438,N_19843,N_18351);
or UO_1439 (O_1439,N_16384,N_17544);
and UO_1440 (O_1440,N_17182,N_18934);
and UO_1441 (O_1441,N_19322,N_18951);
nand UO_1442 (O_1442,N_18179,N_19878);
nand UO_1443 (O_1443,N_18499,N_18510);
and UO_1444 (O_1444,N_19197,N_16360);
nor UO_1445 (O_1445,N_17966,N_17547);
or UO_1446 (O_1446,N_17119,N_16191);
xor UO_1447 (O_1447,N_17979,N_19033);
nor UO_1448 (O_1448,N_19346,N_16397);
or UO_1449 (O_1449,N_17916,N_18316);
or UO_1450 (O_1450,N_19903,N_16965);
or UO_1451 (O_1451,N_19720,N_19818);
nand UO_1452 (O_1452,N_19791,N_16274);
nand UO_1453 (O_1453,N_16689,N_16281);
and UO_1454 (O_1454,N_19815,N_17196);
xnor UO_1455 (O_1455,N_19292,N_19513);
nor UO_1456 (O_1456,N_17774,N_19625);
or UO_1457 (O_1457,N_19242,N_16877);
nand UO_1458 (O_1458,N_19132,N_19182);
or UO_1459 (O_1459,N_19061,N_17833);
or UO_1460 (O_1460,N_17920,N_18245);
and UO_1461 (O_1461,N_17585,N_16289);
or UO_1462 (O_1462,N_16056,N_18735);
or UO_1463 (O_1463,N_17617,N_16854);
or UO_1464 (O_1464,N_17306,N_17705);
nand UO_1465 (O_1465,N_19227,N_18013);
and UO_1466 (O_1466,N_18116,N_18335);
and UO_1467 (O_1467,N_18573,N_18374);
or UO_1468 (O_1468,N_19185,N_16536);
nor UO_1469 (O_1469,N_16587,N_19688);
xnor UO_1470 (O_1470,N_16999,N_16077);
xor UO_1471 (O_1471,N_17667,N_19515);
and UO_1472 (O_1472,N_17053,N_17072);
nor UO_1473 (O_1473,N_16937,N_18853);
nand UO_1474 (O_1474,N_17760,N_16198);
nor UO_1475 (O_1475,N_19987,N_16106);
nand UO_1476 (O_1476,N_17036,N_18571);
and UO_1477 (O_1477,N_19354,N_18362);
and UO_1478 (O_1478,N_16290,N_17472);
nor UO_1479 (O_1479,N_16896,N_17761);
or UO_1480 (O_1480,N_17237,N_19595);
or UO_1481 (O_1481,N_18700,N_16111);
and UO_1482 (O_1482,N_19129,N_16074);
nand UO_1483 (O_1483,N_18494,N_16888);
nand UO_1484 (O_1484,N_16588,N_17352);
nand UO_1485 (O_1485,N_17880,N_17845);
nor UO_1486 (O_1486,N_19653,N_19311);
and UO_1487 (O_1487,N_16545,N_16269);
nand UO_1488 (O_1488,N_19172,N_16906);
or UO_1489 (O_1489,N_18995,N_17496);
or UO_1490 (O_1490,N_17223,N_17304);
and UO_1491 (O_1491,N_16006,N_19454);
xnor UO_1492 (O_1492,N_16324,N_19440);
nor UO_1493 (O_1493,N_19736,N_16651);
nand UO_1494 (O_1494,N_18651,N_19157);
or UO_1495 (O_1495,N_16368,N_18175);
or UO_1496 (O_1496,N_16769,N_18278);
and UO_1497 (O_1497,N_19059,N_16544);
and UO_1498 (O_1498,N_19968,N_18605);
nor UO_1499 (O_1499,N_17784,N_17335);
nand UO_1500 (O_1500,N_17457,N_19866);
nor UO_1501 (O_1501,N_19812,N_17109);
nand UO_1502 (O_1502,N_16539,N_19783);
xor UO_1503 (O_1503,N_19495,N_17160);
nand UO_1504 (O_1504,N_19611,N_18888);
and UO_1505 (O_1505,N_19547,N_16170);
nand UO_1506 (O_1506,N_17080,N_17611);
or UO_1507 (O_1507,N_17876,N_19402);
nor UO_1508 (O_1508,N_19201,N_17074);
nand UO_1509 (O_1509,N_19932,N_16378);
nor UO_1510 (O_1510,N_16950,N_17326);
or UO_1511 (O_1511,N_18717,N_17147);
nand UO_1512 (O_1512,N_18045,N_19308);
nand UO_1513 (O_1513,N_18716,N_18203);
and UO_1514 (O_1514,N_18544,N_16176);
nand UO_1515 (O_1515,N_17473,N_19570);
and UO_1516 (O_1516,N_17047,N_16963);
or UO_1517 (O_1517,N_18923,N_19612);
nand UO_1518 (O_1518,N_17722,N_16815);
or UO_1519 (O_1519,N_19532,N_16479);
nor UO_1520 (O_1520,N_18909,N_17841);
and UO_1521 (O_1521,N_17054,N_19301);
and UO_1522 (O_1522,N_19956,N_17406);
nand UO_1523 (O_1523,N_16518,N_17046);
xor UO_1524 (O_1524,N_19511,N_17901);
and UO_1525 (O_1525,N_17042,N_19336);
nand UO_1526 (O_1526,N_17478,N_16501);
and UO_1527 (O_1527,N_16128,N_18610);
or UO_1528 (O_1528,N_18153,N_16841);
xnor UO_1529 (O_1529,N_17112,N_19383);
nor UO_1530 (O_1530,N_18003,N_17527);
or UO_1531 (O_1531,N_16336,N_17063);
and UO_1532 (O_1532,N_19724,N_19362);
nand UO_1533 (O_1533,N_19341,N_19366);
xor UO_1534 (O_1534,N_16343,N_19858);
and UO_1535 (O_1535,N_18190,N_18303);
nor UO_1536 (O_1536,N_16782,N_18989);
nand UO_1537 (O_1537,N_18427,N_18629);
and UO_1538 (O_1538,N_18699,N_16391);
xor UO_1539 (O_1539,N_16084,N_18246);
or UO_1540 (O_1540,N_19420,N_16261);
nand UO_1541 (O_1541,N_19072,N_18436);
and UO_1542 (O_1542,N_19449,N_19670);
and UO_1543 (O_1543,N_19200,N_19100);
or UO_1544 (O_1544,N_19327,N_17736);
nor UO_1545 (O_1545,N_19888,N_19651);
and UO_1546 (O_1546,N_17861,N_17776);
nand UO_1547 (O_1547,N_18334,N_16316);
or UO_1548 (O_1548,N_17995,N_19047);
nand UO_1549 (O_1549,N_16423,N_18144);
nor UO_1550 (O_1550,N_16674,N_17249);
nand UO_1551 (O_1551,N_16928,N_16069);
xor UO_1552 (O_1552,N_18280,N_18983);
or UO_1553 (O_1553,N_18854,N_18226);
nor UO_1554 (O_1554,N_16700,N_17944);
nand UO_1555 (O_1555,N_18394,N_19264);
xor UO_1556 (O_1556,N_18661,N_16186);
or UO_1557 (O_1557,N_18758,N_16751);
nor UO_1558 (O_1558,N_17221,N_18786);
xnor UO_1559 (O_1559,N_16649,N_19959);
and UO_1560 (O_1560,N_17094,N_17506);
nor UO_1561 (O_1561,N_17114,N_17990);
nor UO_1562 (O_1562,N_17831,N_16092);
and UO_1563 (O_1563,N_16374,N_18860);
or UO_1564 (O_1564,N_16709,N_17012);
nor UO_1565 (O_1565,N_17813,N_17746);
or UO_1566 (O_1566,N_16601,N_19563);
nand UO_1567 (O_1567,N_18921,N_19289);
nand UO_1568 (O_1568,N_17523,N_17236);
or UO_1569 (O_1569,N_17796,N_18966);
or UO_1570 (O_1570,N_19479,N_19917);
nor UO_1571 (O_1571,N_18840,N_19537);
nor UO_1572 (O_1572,N_17690,N_18160);
nor UO_1573 (O_1573,N_17336,N_19825);
and UO_1574 (O_1574,N_18652,N_19499);
nand UO_1575 (O_1575,N_16584,N_16672);
nand UO_1576 (O_1576,N_17707,N_19834);
nor UO_1577 (O_1577,N_18430,N_17409);
or UO_1578 (O_1578,N_17035,N_19413);
nor UO_1579 (O_1579,N_19893,N_19095);
or UO_1580 (O_1580,N_17892,N_19093);
nand UO_1581 (O_1581,N_17134,N_18037);
nand UO_1582 (O_1582,N_18915,N_17911);
xnor UO_1583 (O_1583,N_18275,N_19199);
nand UO_1584 (O_1584,N_19733,N_16154);
and UO_1585 (O_1585,N_17353,N_17836);
nand UO_1586 (O_1586,N_16506,N_17605);
or UO_1587 (O_1587,N_18095,N_18272);
and UO_1588 (O_1588,N_18078,N_19810);
nor UO_1589 (O_1589,N_16654,N_19902);
nand UO_1590 (O_1590,N_17931,N_19152);
nand UO_1591 (O_1591,N_16806,N_16850);
nor UO_1592 (O_1592,N_17621,N_19659);
and UO_1593 (O_1593,N_17227,N_17252);
nand UO_1594 (O_1594,N_18239,N_19694);
or UO_1595 (O_1595,N_17439,N_19497);
or UO_1596 (O_1596,N_16430,N_16453);
or UO_1597 (O_1597,N_17932,N_17909);
or UO_1598 (O_1598,N_16067,N_16638);
nor UO_1599 (O_1599,N_18060,N_19896);
and UO_1600 (O_1600,N_17454,N_18918);
nor UO_1601 (O_1601,N_19553,N_19003);
nor UO_1602 (O_1602,N_19839,N_18899);
or UO_1603 (O_1603,N_16803,N_17691);
nand UO_1604 (O_1604,N_19578,N_16267);
nand UO_1605 (O_1605,N_18736,N_17110);
or UO_1606 (O_1606,N_16105,N_19769);
xnor UO_1607 (O_1607,N_16000,N_16295);
or UO_1608 (O_1608,N_19682,N_18230);
or UO_1609 (O_1609,N_17162,N_17168);
nand UO_1610 (O_1610,N_18057,N_16190);
xor UO_1611 (O_1611,N_19000,N_18827);
nor UO_1612 (O_1612,N_16525,N_18123);
and UO_1613 (O_1613,N_19556,N_19415);
or UO_1614 (O_1614,N_19416,N_16018);
nand UO_1615 (O_1615,N_17759,N_19078);
xnor UO_1616 (O_1616,N_17364,N_16334);
and UO_1617 (O_1617,N_19234,N_17397);
and UO_1618 (O_1618,N_17648,N_16090);
nand UO_1619 (O_1619,N_17566,N_16947);
nand UO_1620 (O_1620,N_16637,N_19324);
nor UO_1621 (O_1621,N_18697,N_19350);
nor UO_1622 (O_1622,N_16571,N_16232);
nand UO_1623 (O_1623,N_18922,N_16797);
or UO_1624 (O_1624,N_17219,N_18180);
nor UO_1625 (O_1625,N_17637,N_17295);
xor UO_1626 (O_1626,N_18892,N_17738);
or UO_1627 (O_1627,N_17789,N_17914);
nand UO_1628 (O_1628,N_18018,N_18014);
xnor UO_1629 (O_1629,N_18799,N_17189);
xor UO_1630 (O_1630,N_19855,N_19946);
nand UO_1631 (O_1631,N_18886,N_18672);
or UO_1632 (O_1632,N_18567,N_16739);
and UO_1633 (O_1633,N_19405,N_17202);
nor UO_1634 (O_1634,N_17369,N_19105);
nand UO_1635 (O_1635,N_17910,N_17443);
and UO_1636 (O_1636,N_17174,N_18101);
and UO_1637 (O_1637,N_19377,N_19167);
xnor UO_1638 (O_1638,N_18960,N_17712);
or UO_1639 (O_1639,N_19153,N_17268);
and UO_1640 (O_1640,N_17085,N_16208);
or UO_1641 (O_1641,N_18597,N_17803);
nor UO_1642 (O_1642,N_19755,N_19471);
or UO_1643 (O_1643,N_17597,N_16282);
xnor UO_1644 (O_1644,N_19117,N_17239);
nand UO_1645 (O_1645,N_16941,N_16097);
xor UO_1646 (O_1646,N_17687,N_19933);
nor UO_1647 (O_1647,N_19412,N_18204);
nor UO_1648 (O_1648,N_18228,N_18705);
or UO_1649 (O_1649,N_17113,N_17452);
and UO_1650 (O_1650,N_17832,N_17301);
nor UO_1651 (O_1651,N_19491,N_19507);
or UO_1652 (O_1652,N_19498,N_19795);
nor UO_1653 (O_1653,N_18485,N_17407);
or UO_1654 (O_1654,N_16790,N_19689);
nand UO_1655 (O_1655,N_19673,N_18755);
nor UO_1656 (O_1656,N_16288,N_19248);
xnor UO_1657 (O_1657,N_18075,N_19837);
nand UO_1658 (O_1658,N_19044,N_19880);
and UO_1659 (O_1659,N_16001,N_16476);
nand UO_1660 (O_1660,N_19505,N_18704);
nor UO_1661 (O_1661,N_16681,N_19372);
xnor UO_1662 (O_1662,N_17885,N_19976);
and UO_1663 (O_1663,N_16175,N_17169);
nand UO_1664 (O_1664,N_16016,N_19490);
nand UO_1665 (O_1665,N_19232,N_19605);
nor UO_1666 (O_1666,N_16909,N_18954);
nor UO_1667 (O_1667,N_18300,N_19609);
nor UO_1668 (O_1668,N_16007,N_19522);
or UO_1669 (O_1669,N_19168,N_19111);
or UO_1670 (O_1670,N_19656,N_18468);
xor UO_1671 (O_1671,N_17843,N_19820);
nor UO_1672 (O_1672,N_17167,N_17908);
nand UO_1673 (O_1673,N_19978,N_18766);
xor UO_1674 (O_1674,N_18482,N_18115);
nand UO_1675 (O_1675,N_19375,N_17805);
or UO_1676 (O_1676,N_19623,N_17627);
and UO_1677 (O_1677,N_16801,N_16998);
and UO_1678 (O_1678,N_16020,N_17197);
and UO_1679 (O_1679,N_17737,N_18855);
or UO_1680 (O_1680,N_17670,N_17391);
nor UO_1681 (O_1681,N_18594,N_19981);
or UO_1682 (O_1682,N_19293,N_17620);
or UO_1683 (O_1683,N_19480,N_18405);
xnor UO_1684 (O_1684,N_16323,N_19091);
nand UO_1685 (O_1685,N_19906,N_16104);
and UO_1686 (O_1686,N_16394,N_18902);
nor UO_1687 (O_1687,N_18353,N_16748);
and UO_1688 (O_1688,N_19342,N_16216);
or UO_1689 (O_1689,N_18679,N_18521);
or UO_1690 (O_1690,N_17312,N_17824);
nand UO_1691 (O_1691,N_19598,N_19114);
nor UO_1692 (O_1692,N_17176,N_16508);
nor UO_1693 (O_1693,N_18350,N_16559);
nor UO_1694 (O_1694,N_18448,N_19877);
nor UO_1695 (O_1695,N_16222,N_19106);
nor UO_1696 (O_1696,N_19516,N_19120);
nor UO_1697 (O_1697,N_18488,N_18727);
xor UO_1698 (O_1698,N_17251,N_17215);
or UO_1699 (O_1699,N_18063,N_16093);
and UO_1700 (O_1700,N_17512,N_18612);
nor UO_1701 (O_1701,N_18801,N_17758);
nor UO_1702 (O_1702,N_17096,N_19216);
nor UO_1703 (O_1703,N_16491,N_19763);
nand UO_1704 (O_1704,N_17582,N_18064);
and UO_1705 (O_1705,N_18354,N_18751);
and UO_1706 (O_1706,N_19546,N_18561);
nand UO_1707 (O_1707,N_16699,N_17800);
and UO_1708 (O_1708,N_17303,N_16387);
nand UO_1709 (O_1709,N_17062,N_17521);
or UO_1710 (O_1710,N_17192,N_16370);
xor UO_1711 (O_1711,N_16040,N_17943);
or UO_1712 (O_1712,N_18583,N_17716);
or UO_1713 (O_1713,N_18449,N_17586);
and UO_1714 (O_1714,N_16779,N_19213);
nor UO_1715 (O_1715,N_18042,N_18338);
or UO_1716 (O_1716,N_19636,N_16912);
nor UO_1717 (O_1717,N_17153,N_16351);
nand UO_1718 (O_1718,N_18459,N_16577);
or UO_1719 (O_1719,N_19895,N_16429);
xor UO_1720 (O_1720,N_18266,N_16033);
or UO_1721 (O_1721,N_16851,N_18110);
and UO_1722 (O_1722,N_18848,N_17149);
nand UO_1723 (O_1723,N_17827,N_19270);
nor UO_1724 (O_1724,N_16593,N_17986);
or UO_1725 (O_1725,N_19330,N_19092);
or UO_1726 (O_1726,N_17381,N_16958);
xor UO_1727 (O_1727,N_18862,N_18505);
xor UO_1728 (O_1728,N_19178,N_16313);
xor UO_1729 (O_1729,N_17525,N_19257);
and UO_1730 (O_1730,N_16619,N_17883);
or UO_1731 (O_1731,N_16540,N_19127);
and UO_1732 (O_1732,N_16767,N_16217);
nor UO_1733 (O_1733,N_16421,N_18695);
or UO_1734 (O_1734,N_18881,N_19559);
and UO_1735 (O_1735,N_18150,N_16650);
xnor UO_1736 (O_1736,N_18526,N_18898);
or UO_1737 (O_1737,N_18531,N_17414);
and UO_1738 (O_1738,N_16583,N_17091);
nor UO_1739 (O_1739,N_19465,N_19678);
nor UO_1740 (O_1740,N_18135,N_16732);
nor UO_1741 (O_1741,N_17809,N_18461);
nor UO_1742 (O_1742,N_17043,N_16492);
and UO_1743 (O_1743,N_16940,N_16096);
or UO_1744 (O_1744,N_19481,N_19554);
and UO_1745 (O_1745,N_17018,N_16484);
nor UO_1746 (O_1746,N_18603,N_16184);
nor UO_1747 (O_1747,N_18295,N_19872);
nor UO_1748 (O_1748,N_16242,N_16059);
and UO_1749 (O_1749,N_19254,N_16145);
or UO_1750 (O_1750,N_16572,N_16460);
nand UO_1751 (O_1751,N_16655,N_17756);
nand UO_1752 (O_1752,N_19004,N_16049);
or UO_1753 (O_1753,N_16371,N_16228);
nand UO_1754 (O_1754,N_16543,N_19728);
xnor UO_1755 (O_1755,N_19641,N_17581);
or UO_1756 (O_1756,N_19467,N_17017);
or UO_1757 (O_1757,N_18646,N_16715);
and UO_1758 (O_1758,N_18464,N_17238);
nand UO_1759 (O_1759,N_17764,N_19035);
or UO_1760 (O_1760,N_18489,N_18475);
and UO_1761 (O_1761,N_16236,N_16171);
nand UO_1762 (O_1762,N_16811,N_18657);
nor UO_1763 (O_1763,N_17373,N_18201);
xnor UO_1764 (O_1764,N_18643,N_16613);
nor UO_1765 (O_1765,N_19735,N_17935);
and UO_1766 (O_1766,N_17632,N_19770);
and UO_1767 (O_1767,N_18993,N_17385);
xnor UO_1768 (O_1768,N_17212,N_17230);
and UO_1769 (O_1769,N_18904,N_16382);
and UO_1770 (O_1770,N_19584,N_18224);
nand UO_1771 (O_1771,N_19600,N_18455);
nor UO_1772 (O_1772,N_16081,N_19568);
or UO_1773 (O_1773,N_16325,N_19156);
and UO_1774 (O_1774,N_19435,N_18641);
nor UO_1775 (O_1775,N_17968,N_19165);
or UO_1776 (O_1776,N_18514,N_16390);
nor UO_1777 (O_1777,N_16454,N_17259);
nand UO_1778 (O_1778,N_18061,N_18090);
or UO_1779 (O_1779,N_19980,N_16404);
xnor UO_1780 (O_1780,N_19911,N_19398);
nor UO_1781 (O_1781,N_19121,N_16904);
and UO_1782 (O_1782,N_18636,N_19439);
or UO_1783 (O_1783,N_18797,N_17945);
nand UO_1784 (O_1784,N_19874,N_19036);
xnor UO_1785 (O_1785,N_19031,N_16224);
xor UO_1786 (O_1786,N_16061,N_18342);
xnor UO_1787 (O_1787,N_16962,N_16246);
and UO_1788 (O_1788,N_17514,N_19566);
or UO_1789 (O_1789,N_17386,N_19534);
nor UO_1790 (O_1790,N_16250,N_18676);
nor UO_1791 (O_1791,N_17603,N_19163);
or UO_1792 (O_1792,N_18296,N_17486);
nor UO_1793 (O_1793,N_16276,N_17850);
nor UO_1794 (O_1794,N_19814,N_18229);
nand UO_1795 (O_1795,N_16381,N_17324);
and UO_1796 (O_1796,N_19055,N_17933);
nor UO_1797 (O_1797,N_17315,N_16771);
xnor UO_1798 (O_1798,N_16865,N_17138);
nand UO_1799 (O_1799,N_18100,N_19798);
xor UO_1800 (O_1800,N_18582,N_16300);
or UO_1801 (O_1801,N_18414,N_17689);
nand UO_1802 (O_1802,N_19021,N_17416);
nor UO_1803 (O_1803,N_17878,N_19974);
and UO_1804 (O_1804,N_17140,N_17952);
nor UO_1805 (O_1805,N_16185,N_18113);
or UO_1806 (O_1806,N_16844,N_19675);
and UO_1807 (O_1807,N_17081,N_19049);
or UO_1808 (O_1808,N_17587,N_18873);
nor UO_1809 (O_1809,N_16573,N_16201);
nand UO_1810 (O_1810,N_17601,N_19503);
and UO_1811 (O_1811,N_17868,N_18001);
nand UO_1812 (O_1812,N_18250,N_16050);
and UO_1813 (O_1813,N_19068,N_18601);
xor UO_1814 (O_1814,N_16335,N_17435);
and UO_1815 (O_1815,N_17193,N_16627);
nand UO_1816 (O_1816,N_16156,N_16310);
xor UO_1817 (O_1817,N_19128,N_19303);
or UO_1818 (O_1818,N_18439,N_17890);
and UO_1819 (O_1819,N_17006,N_19224);
nand UO_1820 (O_1820,N_19096,N_17549);
nand UO_1821 (O_1821,N_18055,N_16745);
or UO_1822 (O_1822,N_16706,N_17654);
and UO_1823 (O_1823,N_18257,N_18509);
and UO_1824 (O_1824,N_17810,N_17159);
or UO_1825 (O_1825,N_19801,N_17562);
or UO_1826 (O_1826,N_19517,N_17964);
and UO_1827 (O_1827,N_17272,N_17778);
nor UO_1828 (O_1828,N_16417,N_17337);
or UO_1829 (O_1829,N_16891,N_17099);
nand UO_1830 (O_1830,N_17108,N_19084);
nor UO_1831 (O_1831,N_17431,N_19725);
and UO_1832 (O_1832,N_17258,N_18200);
nand UO_1833 (O_1833,N_19913,N_18447);
and UO_1834 (O_1834,N_17092,N_17904);
and UO_1835 (O_1835,N_17537,N_17646);
xnor UO_1836 (O_1836,N_19475,N_16200);
and UO_1837 (O_1837,N_16497,N_18425);
nor UO_1838 (O_1838,N_19103,N_16994);
or UO_1839 (O_1839,N_19166,N_17322);
xnor UO_1840 (O_1840,N_16992,N_18412);
nor UO_1841 (O_1841,N_19909,N_16103);
nand UO_1842 (O_1842,N_17704,N_19650);
and UO_1843 (O_1843,N_17660,N_16458);
and UO_1844 (O_1844,N_19309,N_16027);
or UO_1845 (O_1845,N_17338,N_16411);
nor UO_1846 (O_1846,N_19135,N_19506);
nand UO_1847 (O_1847,N_17331,N_17817);
and UO_1848 (O_1848,N_19536,N_17684);
nand UO_1849 (O_1849,N_17930,N_18776);
nand UO_1850 (O_1850,N_16644,N_19824);
or UO_1851 (O_1851,N_18444,N_19472);
nand UO_1852 (O_1852,N_17893,N_18808);
xnor UO_1853 (O_1853,N_19852,N_19040);
nand UO_1854 (O_1854,N_19939,N_16737);
nand UO_1855 (O_1855,N_19710,N_18210);
nand UO_1856 (O_1856,N_16307,N_16723);
and UO_1857 (O_1857,N_19253,N_17434);
nor UO_1858 (O_1858,N_18472,N_19097);
nand UO_1859 (O_1859,N_16762,N_16480);
and UO_1860 (O_1860,N_18517,N_16182);
nand UO_1861 (O_1861,N_17105,N_16592);
xnor UO_1862 (O_1862,N_18282,N_19661);
and UO_1863 (O_1863,N_18143,N_17602);
nand UO_1864 (O_1864,N_18289,N_18496);
and UO_1865 (O_1865,N_17938,N_16320);
nand UO_1866 (O_1866,N_17184,N_19282);
nand UO_1867 (O_1867,N_16278,N_16542);
or UO_1868 (O_1868,N_17057,N_19418);
xnor UO_1869 (O_1869,N_17216,N_19347);
and UO_1870 (O_1870,N_19627,N_17677);
nand UO_1871 (O_1871,N_17777,N_16021);
or UO_1872 (O_1872,N_18974,N_17211);
nor UO_1873 (O_1873,N_19205,N_19115);
nand UO_1874 (O_1874,N_18947,N_16687);
and UO_1875 (O_1875,N_18424,N_17280);
nand UO_1876 (O_1876,N_18836,N_18555);
nand UO_1877 (O_1877,N_19500,N_17014);
nor UO_1878 (O_1878,N_17082,N_19150);
nand UO_1879 (O_1879,N_17102,N_16642);
nand UO_1880 (O_1880,N_19601,N_16434);
or UO_1881 (O_1881,N_18106,N_16717);
xnor UO_1882 (O_1882,N_19145,N_18511);
nand UO_1883 (O_1883,N_19279,N_16419);
or UO_1884 (O_1884,N_17770,N_19143);
or UO_1885 (O_1885,N_19561,N_17694);
or UO_1886 (O_1886,N_18668,N_17664);
nor UO_1887 (O_1887,N_17652,N_17126);
nand UO_1888 (O_1888,N_19606,N_17466);
nand UO_1889 (O_1889,N_17629,N_18022);
and UO_1890 (O_1890,N_17771,N_18790);
nor UO_1891 (O_1891,N_16041,N_16847);
nand UO_1892 (O_1892,N_16943,N_17309);
and UO_1893 (O_1893,N_19461,N_17750);
and UO_1894 (O_1894,N_17526,N_18082);
or UO_1895 (O_1895,N_16695,N_16133);
nand UO_1896 (O_1896,N_19808,N_19771);
xor UO_1897 (O_1897,N_18671,N_19754);
or UO_1898 (O_1898,N_18274,N_18392);
nand UO_1899 (O_1899,N_16830,N_16218);
nand UO_1900 (O_1900,N_16448,N_19564);
and UO_1901 (O_1901,N_18552,N_19256);
nand UO_1902 (O_1902,N_17780,N_18024);
nand UO_1903 (O_1903,N_16738,N_19110);
and UO_1904 (O_1904,N_18232,N_19013);
and UO_1905 (O_1905,N_19447,N_16534);
xnor UO_1906 (O_1906,N_18332,N_19032);
nor UO_1907 (O_1907,N_17293,N_16566);
or UO_1908 (O_1908,N_18151,N_17766);
or UO_1909 (O_1909,N_19723,N_19918);
xor UO_1910 (O_1910,N_19169,N_17294);
nand UO_1911 (O_1911,N_19370,N_17499);
or UO_1912 (O_1912,N_19081,N_18486);
nor UO_1913 (O_1913,N_17779,N_18532);
xnor UO_1914 (O_1914,N_18458,N_19356);
or UO_1915 (O_1915,N_16252,N_17137);
nor UO_1916 (O_1916,N_17356,N_17924);
nand UO_1917 (O_1917,N_19191,N_19846);
nand UO_1918 (O_1918,N_19076,N_17532);
or UO_1919 (O_1919,N_18895,N_18277);
nor UO_1920 (O_1920,N_17264,N_19062);
and UO_1921 (O_1921,N_18833,N_17614);
or UO_1922 (O_1922,N_18233,N_16521);
nor UO_1923 (O_1923,N_16789,N_17129);
nor UO_1924 (O_1924,N_18654,N_19357);
or UO_1925 (O_1925,N_17982,N_18306);
xnor UO_1926 (O_1926,N_19908,N_18513);
nor UO_1927 (O_1927,N_16196,N_16753);
nor UO_1928 (O_1928,N_16505,N_18874);
xnor UO_1929 (O_1929,N_17380,N_17742);
or UO_1930 (O_1930,N_19066,N_19884);
nand UO_1931 (O_1931,N_17869,N_16621);
or UO_1932 (O_1932,N_17033,N_16926);
nor UO_1933 (O_1933,N_16003,N_16765);
and UO_1934 (O_1934,N_19693,N_16398);
nand UO_1935 (O_1935,N_16993,N_17847);
xor UO_1936 (O_1936,N_18417,N_19819);
and UO_1937 (O_1937,N_17325,N_16669);
or UO_1938 (O_1938,N_16187,N_19539);
or UO_1939 (O_1939,N_19287,N_18823);
nand UO_1940 (O_1940,N_18185,N_17274);
and UO_1941 (O_1941,N_18800,N_19617);
and UO_1942 (O_1942,N_16151,N_19158);
nor UO_1943 (O_1943,N_18032,N_17180);
nand UO_1944 (O_1944,N_16995,N_19587);
and UO_1945 (O_1945,N_17447,N_16348);
or UO_1946 (O_1946,N_17718,N_19338);
and UO_1947 (O_1947,N_18906,N_18251);
nor UO_1948 (O_1948,N_18935,N_16702);
nor UO_1949 (O_1949,N_18703,N_19699);
or UO_1950 (O_1950,N_19838,N_19113);
and UO_1951 (O_1951,N_16945,N_18939);
and UO_1952 (O_1952,N_17389,N_18849);
and UO_1953 (O_1953,N_19477,N_17981);
nand UO_1954 (O_1954,N_16907,N_19131);
nor UO_1955 (O_1955,N_17204,N_16283);
or UO_1956 (O_1956,N_17616,N_17089);
nand UO_1957 (O_1957,N_16680,N_17320);
and UO_1958 (O_1958,N_16652,N_18120);
nor UO_1959 (O_1959,N_16352,N_19419);
nor UO_1960 (O_1960,N_19966,N_18725);
nand UO_1961 (O_1961,N_17752,N_19567);
nand UO_1962 (O_1962,N_16731,N_16362);
nor UO_1963 (O_1963,N_16083,N_16568);
and UO_1964 (O_1964,N_16225,N_16898);
nand UO_1965 (O_1965,N_19989,N_17971);
nand UO_1966 (O_1966,N_16957,N_18962);
and UO_1967 (O_1967,N_16569,N_16100);
nor UO_1968 (O_1968,N_18714,N_19247);
or UO_1969 (O_1969,N_18360,N_18696);
nand UO_1970 (O_1970,N_19792,N_17044);
or UO_1971 (O_1971,N_17065,N_16415);
or UO_1972 (O_1972,N_18172,N_17117);
nand UO_1973 (O_1973,N_18829,N_17480);
nor UO_1974 (O_1974,N_19944,N_19865);
or UO_1975 (O_1975,N_18501,N_19284);
nand UO_1976 (O_1976,N_16873,N_17307);
or UO_1977 (O_1977,N_18649,N_16976);
xor UO_1978 (O_1978,N_18237,N_16934);
nand UO_1979 (O_1979,N_18403,N_16135);
and UO_1980 (O_1980,N_19151,N_19267);
xor UO_1981 (O_1981,N_17178,N_18068);
nor UO_1982 (O_1982,N_17093,N_16794);
nand UO_1983 (O_1983,N_17709,N_16708);
and UO_1984 (O_1984,N_18069,N_18685);
xnor UO_1985 (O_1985,N_16643,N_18812);
and UO_1986 (O_1986,N_17975,N_17494);
or UO_1987 (O_1987,N_19259,N_18088);
nor UO_1988 (O_1988,N_18097,N_17007);
nand UO_1989 (O_1989,N_17387,N_16774);
and UO_1990 (O_1990,N_18214,N_19541);
and UO_1991 (O_1991,N_17940,N_18196);
nor UO_1992 (O_1992,N_18762,N_17772);
nor UO_1993 (O_1993,N_18434,N_18789);
and UO_1994 (O_1994,N_18681,N_16817);
and UO_1995 (O_1995,N_17569,N_17493);
nand UO_1996 (O_1996,N_16546,N_17145);
and UO_1997 (O_1997,N_19363,N_16741);
and UO_1998 (O_1998,N_18554,N_17905);
or UO_1999 (O_1999,N_18875,N_19054);
nor UO_2000 (O_2000,N_19973,N_17437);
and UO_2001 (O_2001,N_17758,N_19851);
or UO_2002 (O_2002,N_18566,N_19304);
nor UO_2003 (O_2003,N_18766,N_19537);
and UO_2004 (O_2004,N_18119,N_17749);
and UO_2005 (O_2005,N_16803,N_18615);
and UO_2006 (O_2006,N_19090,N_18426);
nand UO_2007 (O_2007,N_18313,N_16521);
or UO_2008 (O_2008,N_18964,N_19893);
and UO_2009 (O_2009,N_17667,N_17184);
and UO_2010 (O_2010,N_18789,N_17832);
xor UO_2011 (O_2011,N_18727,N_18521);
or UO_2012 (O_2012,N_19759,N_17815);
nor UO_2013 (O_2013,N_17189,N_19861);
nor UO_2014 (O_2014,N_19885,N_16157);
nand UO_2015 (O_2015,N_16036,N_17263);
and UO_2016 (O_2016,N_17747,N_18708);
nand UO_2017 (O_2017,N_19757,N_16518);
or UO_2018 (O_2018,N_18252,N_19263);
nand UO_2019 (O_2019,N_17973,N_19502);
nand UO_2020 (O_2020,N_18025,N_18342);
nand UO_2021 (O_2021,N_18967,N_16435);
or UO_2022 (O_2022,N_16528,N_18417);
or UO_2023 (O_2023,N_19967,N_17698);
or UO_2024 (O_2024,N_17914,N_16726);
nand UO_2025 (O_2025,N_17704,N_19732);
nand UO_2026 (O_2026,N_16837,N_18994);
and UO_2027 (O_2027,N_16709,N_19620);
or UO_2028 (O_2028,N_18600,N_19377);
or UO_2029 (O_2029,N_18405,N_17402);
nor UO_2030 (O_2030,N_17276,N_16703);
nor UO_2031 (O_2031,N_16529,N_17978);
and UO_2032 (O_2032,N_16702,N_18829);
nor UO_2033 (O_2033,N_19235,N_18606);
nor UO_2034 (O_2034,N_17269,N_16464);
or UO_2035 (O_2035,N_18375,N_18275);
or UO_2036 (O_2036,N_19981,N_19596);
nand UO_2037 (O_2037,N_17757,N_16435);
and UO_2038 (O_2038,N_16690,N_19870);
xnor UO_2039 (O_2039,N_17874,N_16188);
nor UO_2040 (O_2040,N_19823,N_16417);
or UO_2041 (O_2041,N_16502,N_16573);
nor UO_2042 (O_2042,N_19961,N_16064);
nand UO_2043 (O_2043,N_18653,N_17457);
nand UO_2044 (O_2044,N_17744,N_16463);
xor UO_2045 (O_2045,N_19394,N_16094);
or UO_2046 (O_2046,N_18508,N_19997);
nor UO_2047 (O_2047,N_19967,N_16099);
and UO_2048 (O_2048,N_17755,N_17228);
or UO_2049 (O_2049,N_17042,N_17386);
or UO_2050 (O_2050,N_17623,N_17273);
nor UO_2051 (O_2051,N_18809,N_16622);
nor UO_2052 (O_2052,N_17508,N_18848);
or UO_2053 (O_2053,N_17175,N_19224);
nand UO_2054 (O_2054,N_18512,N_16112);
nand UO_2055 (O_2055,N_19973,N_16059);
nor UO_2056 (O_2056,N_19703,N_17349);
and UO_2057 (O_2057,N_19155,N_19111);
nand UO_2058 (O_2058,N_17329,N_17827);
or UO_2059 (O_2059,N_16220,N_18273);
or UO_2060 (O_2060,N_18179,N_17893);
nand UO_2061 (O_2061,N_19275,N_16262);
nand UO_2062 (O_2062,N_17559,N_17696);
nand UO_2063 (O_2063,N_16243,N_17568);
and UO_2064 (O_2064,N_17115,N_16621);
nor UO_2065 (O_2065,N_16716,N_18643);
and UO_2066 (O_2066,N_16605,N_19660);
xor UO_2067 (O_2067,N_17902,N_16295);
nand UO_2068 (O_2068,N_19519,N_18064);
nand UO_2069 (O_2069,N_18088,N_17563);
and UO_2070 (O_2070,N_18949,N_19329);
nand UO_2071 (O_2071,N_18367,N_18864);
nand UO_2072 (O_2072,N_19581,N_17587);
and UO_2073 (O_2073,N_16209,N_17599);
or UO_2074 (O_2074,N_16983,N_17340);
nor UO_2075 (O_2075,N_17365,N_17909);
and UO_2076 (O_2076,N_18306,N_19508);
and UO_2077 (O_2077,N_17097,N_18319);
or UO_2078 (O_2078,N_18776,N_19238);
nor UO_2079 (O_2079,N_18724,N_16755);
nor UO_2080 (O_2080,N_19554,N_17156);
xnor UO_2081 (O_2081,N_17343,N_17824);
or UO_2082 (O_2082,N_17505,N_19072);
and UO_2083 (O_2083,N_17758,N_16341);
nor UO_2084 (O_2084,N_16030,N_17902);
and UO_2085 (O_2085,N_19640,N_19733);
nor UO_2086 (O_2086,N_16738,N_19987);
xnor UO_2087 (O_2087,N_19829,N_18188);
and UO_2088 (O_2088,N_16116,N_19563);
or UO_2089 (O_2089,N_17238,N_19561);
and UO_2090 (O_2090,N_16438,N_17555);
nand UO_2091 (O_2091,N_18547,N_18918);
nand UO_2092 (O_2092,N_19511,N_17767);
nor UO_2093 (O_2093,N_16764,N_16296);
or UO_2094 (O_2094,N_16955,N_16184);
xor UO_2095 (O_2095,N_19635,N_17528);
and UO_2096 (O_2096,N_17945,N_19182);
nor UO_2097 (O_2097,N_16594,N_16364);
nand UO_2098 (O_2098,N_16154,N_16291);
xnor UO_2099 (O_2099,N_16254,N_17988);
nand UO_2100 (O_2100,N_17531,N_18686);
and UO_2101 (O_2101,N_17456,N_17555);
or UO_2102 (O_2102,N_17031,N_19867);
or UO_2103 (O_2103,N_19708,N_19790);
and UO_2104 (O_2104,N_17070,N_18162);
nand UO_2105 (O_2105,N_17772,N_17832);
or UO_2106 (O_2106,N_19363,N_19100);
nor UO_2107 (O_2107,N_18386,N_17725);
xnor UO_2108 (O_2108,N_17236,N_19174);
nand UO_2109 (O_2109,N_17489,N_18783);
nand UO_2110 (O_2110,N_16143,N_19182);
and UO_2111 (O_2111,N_18050,N_17478);
and UO_2112 (O_2112,N_16963,N_19804);
xnor UO_2113 (O_2113,N_17323,N_18560);
nand UO_2114 (O_2114,N_19269,N_19521);
or UO_2115 (O_2115,N_18763,N_19842);
and UO_2116 (O_2116,N_17516,N_17240);
nand UO_2117 (O_2117,N_18589,N_17170);
nor UO_2118 (O_2118,N_18986,N_18344);
or UO_2119 (O_2119,N_16857,N_16461);
or UO_2120 (O_2120,N_18518,N_16279);
or UO_2121 (O_2121,N_18955,N_16877);
xnor UO_2122 (O_2122,N_17115,N_19331);
and UO_2123 (O_2123,N_19716,N_17151);
nand UO_2124 (O_2124,N_18890,N_17490);
nor UO_2125 (O_2125,N_19780,N_19751);
and UO_2126 (O_2126,N_17112,N_18530);
nand UO_2127 (O_2127,N_18205,N_19809);
nor UO_2128 (O_2128,N_16895,N_17235);
nor UO_2129 (O_2129,N_19080,N_17473);
nand UO_2130 (O_2130,N_18068,N_19049);
nor UO_2131 (O_2131,N_16448,N_17945);
nor UO_2132 (O_2132,N_16313,N_16286);
nor UO_2133 (O_2133,N_16729,N_17461);
and UO_2134 (O_2134,N_16851,N_18379);
and UO_2135 (O_2135,N_16201,N_17547);
nor UO_2136 (O_2136,N_16197,N_17769);
and UO_2137 (O_2137,N_19882,N_18720);
xnor UO_2138 (O_2138,N_16574,N_17854);
nand UO_2139 (O_2139,N_18984,N_18299);
xnor UO_2140 (O_2140,N_19854,N_19559);
nor UO_2141 (O_2141,N_16029,N_19494);
or UO_2142 (O_2142,N_19621,N_19313);
and UO_2143 (O_2143,N_18150,N_19354);
and UO_2144 (O_2144,N_16253,N_19743);
nand UO_2145 (O_2145,N_18072,N_18052);
or UO_2146 (O_2146,N_17965,N_16941);
and UO_2147 (O_2147,N_19318,N_17066);
xnor UO_2148 (O_2148,N_18581,N_19416);
nor UO_2149 (O_2149,N_16691,N_16721);
or UO_2150 (O_2150,N_16272,N_19153);
or UO_2151 (O_2151,N_16318,N_19133);
and UO_2152 (O_2152,N_18077,N_19448);
xor UO_2153 (O_2153,N_16464,N_16752);
or UO_2154 (O_2154,N_16049,N_16668);
or UO_2155 (O_2155,N_17713,N_19743);
and UO_2156 (O_2156,N_17489,N_17784);
nor UO_2157 (O_2157,N_18069,N_16259);
or UO_2158 (O_2158,N_18106,N_16512);
xnor UO_2159 (O_2159,N_16096,N_18975);
xor UO_2160 (O_2160,N_19582,N_16597);
nor UO_2161 (O_2161,N_17360,N_17722);
or UO_2162 (O_2162,N_17350,N_19049);
and UO_2163 (O_2163,N_19056,N_19601);
and UO_2164 (O_2164,N_18216,N_18155);
xnor UO_2165 (O_2165,N_17092,N_17592);
or UO_2166 (O_2166,N_16297,N_18726);
nand UO_2167 (O_2167,N_16496,N_18115);
nand UO_2168 (O_2168,N_19520,N_18064);
nor UO_2169 (O_2169,N_17355,N_17011);
and UO_2170 (O_2170,N_18963,N_17353);
nor UO_2171 (O_2171,N_16070,N_16051);
nand UO_2172 (O_2172,N_17651,N_19971);
xnor UO_2173 (O_2173,N_19500,N_16895);
or UO_2174 (O_2174,N_19519,N_19382);
or UO_2175 (O_2175,N_17690,N_18497);
xor UO_2176 (O_2176,N_17621,N_19603);
nand UO_2177 (O_2177,N_18634,N_17086);
xor UO_2178 (O_2178,N_17815,N_19510);
nor UO_2179 (O_2179,N_16697,N_17252);
or UO_2180 (O_2180,N_18016,N_16980);
nor UO_2181 (O_2181,N_19267,N_18047);
nand UO_2182 (O_2182,N_16188,N_16428);
and UO_2183 (O_2183,N_18737,N_18865);
nor UO_2184 (O_2184,N_18172,N_16183);
or UO_2185 (O_2185,N_19022,N_19344);
or UO_2186 (O_2186,N_18374,N_19053);
and UO_2187 (O_2187,N_16356,N_17962);
or UO_2188 (O_2188,N_16529,N_18393);
nand UO_2189 (O_2189,N_18516,N_16762);
nor UO_2190 (O_2190,N_16936,N_16476);
or UO_2191 (O_2191,N_17945,N_16091);
and UO_2192 (O_2192,N_17810,N_16183);
nand UO_2193 (O_2193,N_17483,N_19314);
or UO_2194 (O_2194,N_16741,N_18313);
nand UO_2195 (O_2195,N_16532,N_18285);
nand UO_2196 (O_2196,N_16954,N_18182);
or UO_2197 (O_2197,N_18731,N_19203);
nor UO_2198 (O_2198,N_17104,N_17192);
nor UO_2199 (O_2199,N_17171,N_16164);
nor UO_2200 (O_2200,N_16105,N_19097);
nor UO_2201 (O_2201,N_16261,N_18083);
nand UO_2202 (O_2202,N_16569,N_16963);
nor UO_2203 (O_2203,N_16687,N_18957);
nor UO_2204 (O_2204,N_17874,N_16331);
or UO_2205 (O_2205,N_17083,N_16858);
nor UO_2206 (O_2206,N_17190,N_18210);
nand UO_2207 (O_2207,N_19698,N_18810);
nand UO_2208 (O_2208,N_19340,N_18982);
or UO_2209 (O_2209,N_17946,N_16823);
nand UO_2210 (O_2210,N_17580,N_16058);
and UO_2211 (O_2211,N_16658,N_19831);
nand UO_2212 (O_2212,N_17964,N_17857);
or UO_2213 (O_2213,N_18151,N_16595);
nor UO_2214 (O_2214,N_17645,N_17928);
or UO_2215 (O_2215,N_18463,N_16003);
or UO_2216 (O_2216,N_18443,N_18145);
or UO_2217 (O_2217,N_17056,N_16837);
and UO_2218 (O_2218,N_18392,N_19286);
nand UO_2219 (O_2219,N_17256,N_16964);
and UO_2220 (O_2220,N_17788,N_17961);
nand UO_2221 (O_2221,N_17542,N_17914);
nor UO_2222 (O_2222,N_18484,N_16420);
nand UO_2223 (O_2223,N_18759,N_18113);
and UO_2224 (O_2224,N_18428,N_17247);
nand UO_2225 (O_2225,N_16281,N_16892);
nand UO_2226 (O_2226,N_17885,N_17833);
or UO_2227 (O_2227,N_19738,N_18496);
or UO_2228 (O_2228,N_16364,N_17532);
nor UO_2229 (O_2229,N_18141,N_17533);
or UO_2230 (O_2230,N_18634,N_18061);
and UO_2231 (O_2231,N_16847,N_19447);
or UO_2232 (O_2232,N_18710,N_18358);
and UO_2233 (O_2233,N_18797,N_18505);
nand UO_2234 (O_2234,N_19458,N_19982);
or UO_2235 (O_2235,N_18274,N_18680);
nand UO_2236 (O_2236,N_16188,N_19766);
and UO_2237 (O_2237,N_18242,N_16427);
or UO_2238 (O_2238,N_18179,N_19867);
nor UO_2239 (O_2239,N_18413,N_16251);
or UO_2240 (O_2240,N_19750,N_17837);
nor UO_2241 (O_2241,N_16775,N_17534);
nand UO_2242 (O_2242,N_16692,N_17871);
or UO_2243 (O_2243,N_18997,N_17902);
or UO_2244 (O_2244,N_16404,N_18800);
nor UO_2245 (O_2245,N_17398,N_17267);
or UO_2246 (O_2246,N_19779,N_16119);
nand UO_2247 (O_2247,N_17139,N_17546);
nand UO_2248 (O_2248,N_16892,N_19590);
nand UO_2249 (O_2249,N_17821,N_19482);
nor UO_2250 (O_2250,N_19564,N_16283);
nand UO_2251 (O_2251,N_17515,N_17069);
nand UO_2252 (O_2252,N_18908,N_19939);
nand UO_2253 (O_2253,N_16264,N_16469);
nor UO_2254 (O_2254,N_19072,N_18604);
nor UO_2255 (O_2255,N_18373,N_19134);
nor UO_2256 (O_2256,N_19724,N_16265);
nand UO_2257 (O_2257,N_18403,N_19090);
or UO_2258 (O_2258,N_19173,N_17897);
xor UO_2259 (O_2259,N_19397,N_16487);
or UO_2260 (O_2260,N_17634,N_17914);
nor UO_2261 (O_2261,N_16144,N_17939);
xnor UO_2262 (O_2262,N_18819,N_19060);
nand UO_2263 (O_2263,N_18745,N_18248);
and UO_2264 (O_2264,N_18364,N_16720);
nor UO_2265 (O_2265,N_16049,N_18740);
and UO_2266 (O_2266,N_17993,N_18668);
or UO_2267 (O_2267,N_19753,N_16379);
nand UO_2268 (O_2268,N_16742,N_19307);
xnor UO_2269 (O_2269,N_16838,N_19750);
or UO_2270 (O_2270,N_19695,N_18722);
nor UO_2271 (O_2271,N_19792,N_18622);
xnor UO_2272 (O_2272,N_19120,N_17678);
nand UO_2273 (O_2273,N_17855,N_17142);
and UO_2274 (O_2274,N_18762,N_19159);
or UO_2275 (O_2275,N_17825,N_16240);
and UO_2276 (O_2276,N_19143,N_19394);
xnor UO_2277 (O_2277,N_16518,N_17993);
nand UO_2278 (O_2278,N_17497,N_19607);
nor UO_2279 (O_2279,N_17310,N_16543);
and UO_2280 (O_2280,N_19554,N_16931);
nor UO_2281 (O_2281,N_19345,N_16503);
nand UO_2282 (O_2282,N_17012,N_16558);
or UO_2283 (O_2283,N_19040,N_19083);
nor UO_2284 (O_2284,N_18436,N_19124);
nand UO_2285 (O_2285,N_17130,N_16058);
nand UO_2286 (O_2286,N_18789,N_18594);
and UO_2287 (O_2287,N_18011,N_18344);
nor UO_2288 (O_2288,N_16020,N_18844);
nor UO_2289 (O_2289,N_19759,N_17681);
nand UO_2290 (O_2290,N_18581,N_18431);
nand UO_2291 (O_2291,N_19957,N_19097);
xnor UO_2292 (O_2292,N_17939,N_16322);
nor UO_2293 (O_2293,N_19169,N_18162);
and UO_2294 (O_2294,N_16234,N_19332);
nand UO_2295 (O_2295,N_16664,N_19305);
nor UO_2296 (O_2296,N_17966,N_16569);
and UO_2297 (O_2297,N_19473,N_16376);
nand UO_2298 (O_2298,N_19160,N_16713);
xnor UO_2299 (O_2299,N_19836,N_17625);
or UO_2300 (O_2300,N_16166,N_18470);
nor UO_2301 (O_2301,N_16634,N_19328);
nand UO_2302 (O_2302,N_18813,N_16580);
or UO_2303 (O_2303,N_17103,N_17925);
and UO_2304 (O_2304,N_19396,N_19732);
nor UO_2305 (O_2305,N_18891,N_18935);
nand UO_2306 (O_2306,N_16534,N_17856);
nor UO_2307 (O_2307,N_18721,N_17245);
nand UO_2308 (O_2308,N_17000,N_16004);
nor UO_2309 (O_2309,N_16894,N_17519);
and UO_2310 (O_2310,N_18556,N_16221);
and UO_2311 (O_2311,N_17323,N_16549);
or UO_2312 (O_2312,N_17809,N_16827);
and UO_2313 (O_2313,N_19039,N_17354);
or UO_2314 (O_2314,N_16491,N_16553);
nand UO_2315 (O_2315,N_19972,N_17630);
and UO_2316 (O_2316,N_17537,N_18387);
nand UO_2317 (O_2317,N_19718,N_18746);
nor UO_2318 (O_2318,N_17550,N_16211);
nand UO_2319 (O_2319,N_18080,N_18011);
and UO_2320 (O_2320,N_19259,N_19288);
and UO_2321 (O_2321,N_16879,N_18032);
nor UO_2322 (O_2322,N_16367,N_17317);
nor UO_2323 (O_2323,N_16132,N_19709);
nand UO_2324 (O_2324,N_16211,N_16942);
nor UO_2325 (O_2325,N_18539,N_17498);
or UO_2326 (O_2326,N_18603,N_18048);
or UO_2327 (O_2327,N_18110,N_19508);
and UO_2328 (O_2328,N_18592,N_19322);
nor UO_2329 (O_2329,N_19714,N_17044);
or UO_2330 (O_2330,N_17044,N_19059);
and UO_2331 (O_2331,N_18401,N_19112);
or UO_2332 (O_2332,N_16771,N_19966);
or UO_2333 (O_2333,N_16896,N_18101);
and UO_2334 (O_2334,N_18014,N_18275);
or UO_2335 (O_2335,N_18126,N_17674);
nand UO_2336 (O_2336,N_16789,N_19176);
or UO_2337 (O_2337,N_17838,N_16107);
nand UO_2338 (O_2338,N_19780,N_16783);
nor UO_2339 (O_2339,N_17753,N_16549);
nand UO_2340 (O_2340,N_17312,N_18554);
or UO_2341 (O_2341,N_16562,N_19204);
or UO_2342 (O_2342,N_16474,N_19565);
nand UO_2343 (O_2343,N_19438,N_17738);
nand UO_2344 (O_2344,N_18442,N_16385);
and UO_2345 (O_2345,N_17169,N_16514);
or UO_2346 (O_2346,N_16534,N_16076);
nor UO_2347 (O_2347,N_16730,N_17460);
nor UO_2348 (O_2348,N_19153,N_18233);
or UO_2349 (O_2349,N_19443,N_19328);
or UO_2350 (O_2350,N_18324,N_18389);
or UO_2351 (O_2351,N_16763,N_16846);
and UO_2352 (O_2352,N_16132,N_17227);
nor UO_2353 (O_2353,N_16704,N_18524);
nand UO_2354 (O_2354,N_17887,N_19768);
or UO_2355 (O_2355,N_19355,N_17371);
nor UO_2356 (O_2356,N_16338,N_17051);
and UO_2357 (O_2357,N_19454,N_17245);
and UO_2358 (O_2358,N_19649,N_17541);
nor UO_2359 (O_2359,N_17197,N_16496);
nand UO_2360 (O_2360,N_19884,N_19589);
nand UO_2361 (O_2361,N_17875,N_18618);
and UO_2362 (O_2362,N_16277,N_18010);
or UO_2363 (O_2363,N_17998,N_19524);
nand UO_2364 (O_2364,N_18515,N_17943);
nand UO_2365 (O_2365,N_16740,N_17775);
nor UO_2366 (O_2366,N_18682,N_16056);
or UO_2367 (O_2367,N_19835,N_19518);
xor UO_2368 (O_2368,N_18570,N_19537);
nor UO_2369 (O_2369,N_17965,N_19211);
nor UO_2370 (O_2370,N_17866,N_17307);
and UO_2371 (O_2371,N_16249,N_18653);
nand UO_2372 (O_2372,N_19634,N_17547);
nand UO_2373 (O_2373,N_17107,N_17713);
nand UO_2374 (O_2374,N_18231,N_18145);
xnor UO_2375 (O_2375,N_19611,N_18320);
or UO_2376 (O_2376,N_16765,N_19733);
or UO_2377 (O_2377,N_18942,N_19816);
and UO_2378 (O_2378,N_18491,N_16831);
or UO_2379 (O_2379,N_16820,N_16103);
nand UO_2380 (O_2380,N_16757,N_19818);
or UO_2381 (O_2381,N_19104,N_19793);
nor UO_2382 (O_2382,N_19013,N_19145);
and UO_2383 (O_2383,N_16438,N_18848);
nand UO_2384 (O_2384,N_16340,N_16748);
or UO_2385 (O_2385,N_18444,N_17246);
and UO_2386 (O_2386,N_18118,N_18574);
and UO_2387 (O_2387,N_18812,N_16973);
nand UO_2388 (O_2388,N_17599,N_16942);
xnor UO_2389 (O_2389,N_19833,N_19157);
and UO_2390 (O_2390,N_19956,N_16637);
nand UO_2391 (O_2391,N_17511,N_19963);
or UO_2392 (O_2392,N_17185,N_16627);
and UO_2393 (O_2393,N_16062,N_17187);
or UO_2394 (O_2394,N_16288,N_16891);
nor UO_2395 (O_2395,N_19475,N_17313);
and UO_2396 (O_2396,N_18145,N_17782);
nor UO_2397 (O_2397,N_17706,N_17378);
xor UO_2398 (O_2398,N_17445,N_17831);
and UO_2399 (O_2399,N_18979,N_17484);
nor UO_2400 (O_2400,N_17491,N_17188);
and UO_2401 (O_2401,N_16054,N_17654);
nand UO_2402 (O_2402,N_19045,N_17115);
nand UO_2403 (O_2403,N_16152,N_17970);
nor UO_2404 (O_2404,N_18453,N_18586);
nand UO_2405 (O_2405,N_16268,N_16058);
nand UO_2406 (O_2406,N_17068,N_17738);
nand UO_2407 (O_2407,N_16198,N_18724);
nor UO_2408 (O_2408,N_18080,N_18092);
and UO_2409 (O_2409,N_16662,N_19202);
nor UO_2410 (O_2410,N_17769,N_19444);
or UO_2411 (O_2411,N_16172,N_19167);
or UO_2412 (O_2412,N_18691,N_17195);
and UO_2413 (O_2413,N_16647,N_17518);
nand UO_2414 (O_2414,N_16069,N_17360);
nand UO_2415 (O_2415,N_18962,N_19999);
and UO_2416 (O_2416,N_16991,N_16017);
xor UO_2417 (O_2417,N_16421,N_19554);
or UO_2418 (O_2418,N_18568,N_17188);
and UO_2419 (O_2419,N_19361,N_19135);
and UO_2420 (O_2420,N_19415,N_19098);
or UO_2421 (O_2421,N_19553,N_19181);
or UO_2422 (O_2422,N_18958,N_16766);
nand UO_2423 (O_2423,N_18092,N_17293);
nand UO_2424 (O_2424,N_19227,N_17350);
xor UO_2425 (O_2425,N_17755,N_19392);
nor UO_2426 (O_2426,N_18495,N_18849);
nor UO_2427 (O_2427,N_16213,N_17335);
nand UO_2428 (O_2428,N_17084,N_16979);
nand UO_2429 (O_2429,N_17956,N_17083);
xor UO_2430 (O_2430,N_16746,N_19628);
xor UO_2431 (O_2431,N_16438,N_17747);
xnor UO_2432 (O_2432,N_18078,N_19269);
or UO_2433 (O_2433,N_17575,N_16349);
nand UO_2434 (O_2434,N_18814,N_19388);
nor UO_2435 (O_2435,N_19300,N_18028);
or UO_2436 (O_2436,N_17065,N_19566);
nor UO_2437 (O_2437,N_16136,N_16215);
or UO_2438 (O_2438,N_17903,N_16318);
nand UO_2439 (O_2439,N_17434,N_17150);
nor UO_2440 (O_2440,N_19511,N_18746);
or UO_2441 (O_2441,N_19877,N_18900);
nand UO_2442 (O_2442,N_17602,N_18135);
and UO_2443 (O_2443,N_17956,N_18341);
nand UO_2444 (O_2444,N_17079,N_18679);
nand UO_2445 (O_2445,N_19045,N_18119);
nor UO_2446 (O_2446,N_19606,N_18855);
or UO_2447 (O_2447,N_16864,N_16752);
and UO_2448 (O_2448,N_18069,N_19629);
nor UO_2449 (O_2449,N_17388,N_16042);
xnor UO_2450 (O_2450,N_17336,N_18258);
or UO_2451 (O_2451,N_17917,N_16931);
or UO_2452 (O_2452,N_19886,N_16949);
and UO_2453 (O_2453,N_18376,N_17245);
and UO_2454 (O_2454,N_17016,N_16345);
nor UO_2455 (O_2455,N_19940,N_19119);
xor UO_2456 (O_2456,N_17370,N_19912);
xor UO_2457 (O_2457,N_16160,N_18735);
nand UO_2458 (O_2458,N_17919,N_17952);
or UO_2459 (O_2459,N_18931,N_17943);
nand UO_2460 (O_2460,N_19352,N_16323);
nor UO_2461 (O_2461,N_16303,N_16829);
and UO_2462 (O_2462,N_16297,N_19651);
or UO_2463 (O_2463,N_16887,N_16991);
nand UO_2464 (O_2464,N_16489,N_18663);
nand UO_2465 (O_2465,N_18583,N_18704);
nand UO_2466 (O_2466,N_19258,N_18418);
nand UO_2467 (O_2467,N_19897,N_16389);
or UO_2468 (O_2468,N_19050,N_19932);
or UO_2469 (O_2469,N_17634,N_16897);
and UO_2470 (O_2470,N_19444,N_19084);
nand UO_2471 (O_2471,N_18475,N_17122);
and UO_2472 (O_2472,N_17319,N_18315);
and UO_2473 (O_2473,N_17948,N_18852);
and UO_2474 (O_2474,N_18298,N_16304);
and UO_2475 (O_2475,N_17491,N_17619);
and UO_2476 (O_2476,N_19592,N_17428);
nand UO_2477 (O_2477,N_16509,N_16820);
and UO_2478 (O_2478,N_18898,N_19744);
nor UO_2479 (O_2479,N_16888,N_18019);
nand UO_2480 (O_2480,N_19367,N_17986);
xor UO_2481 (O_2481,N_18258,N_17665);
nor UO_2482 (O_2482,N_19514,N_16963);
and UO_2483 (O_2483,N_17980,N_17369);
nand UO_2484 (O_2484,N_19374,N_17178);
nand UO_2485 (O_2485,N_19049,N_16914);
nand UO_2486 (O_2486,N_19778,N_19089);
nand UO_2487 (O_2487,N_16813,N_17957);
xnor UO_2488 (O_2488,N_18306,N_19015);
nand UO_2489 (O_2489,N_16245,N_18507);
xnor UO_2490 (O_2490,N_16224,N_17399);
nor UO_2491 (O_2491,N_16315,N_18323);
or UO_2492 (O_2492,N_18599,N_16874);
or UO_2493 (O_2493,N_16663,N_19375);
and UO_2494 (O_2494,N_17201,N_16014);
nand UO_2495 (O_2495,N_17541,N_19731);
nand UO_2496 (O_2496,N_19293,N_18958);
nand UO_2497 (O_2497,N_19819,N_19161);
or UO_2498 (O_2498,N_18795,N_19655);
or UO_2499 (O_2499,N_18382,N_17499);
endmodule