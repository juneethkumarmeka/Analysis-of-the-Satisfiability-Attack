module basic_2500_25000_3000_4_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18835,N_18836,N_18837,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18864,N_18866,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18983,N_18984,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19230,N_19231,N_19232,N_19233,N_19234,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19315,N_19316,N_19317,N_19318,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19425,N_19426,N_19427,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19517,N_19518,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19697,N_19698,N_19699,N_19700,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19847,N_19848,N_19849,N_19850,N_19851,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19873,N_19874,N_19875,N_19876,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20012,N_20013,N_20014,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20346,N_20347,N_20348,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20654,N_20655,N_20656,N_20657,N_20658,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20693,N_20694,N_20695,N_20696,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20871,N_20872,N_20873,N_20874,N_20875,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21102,N_21103,N_21104,N_21105,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21306,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21463,N_21464,N_21465,N_21466,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21654,N_21655,N_21657,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22020,N_22021,N_22022,N_22023,N_22024,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22117,N_22118,N_22119,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22269,N_22270,N_22271,N_22272,N_22274,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22283,N_22284,N_22285,N_22286,N_22287,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22646,N_22647,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22683,N_22684,N_22685,N_22686,N_22687,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22809,N_22810,N_22811,N_22812,N_22813,N_22815,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23140,N_23141,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23352,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23374,N_23375,N_23376,N_23377,N_23378,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23387,N_23388,N_23389,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23427,N_23428,N_23429,N_23430,N_23431,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23530,N_23531,N_23533,N_23534,N_23536,N_23537,N_23538,N_23539,N_23541,N_23542,N_23543,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23564,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23698,N_23699,N_23700,N_23701,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23733,N_23734,N_23735,N_23736,N_23737,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23805,N_23806,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23976,N_23977,N_23978,N_23979,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23991,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24573,N_24574,N_24575,N_24576,N_24577,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24725,N_24726,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24753,N_24754,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24781,N_24782,N_24783,N_24784,N_24785,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24844,N_24845,N_24846,N_24847,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24943,N_24944,N_24945,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_1158,In_2121);
or U1 (N_1,In_504,In_1574);
and U2 (N_2,In_1436,In_1081);
nor U3 (N_3,In_1383,In_100);
and U4 (N_4,In_2239,In_1189);
xnor U5 (N_5,In_2120,In_2045);
nor U6 (N_6,In_275,In_159);
nor U7 (N_7,In_655,In_976);
nor U8 (N_8,In_2448,In_2280);
or U9 (N_9,In_459,In_1555);
nor U10 (N_10,In_1918,In_1530);
and U11 (N_11,In_1341,In_2252);
nor U12 (N_12,In_720,In_709);
xnor U13 (N_13,In_227,In_1859);
nor U14 (N_14,In_70,In_2283);
and U15 (N_15,In_253,In_1039);
nor U16 (N_16,In_1803,In_405);
or U17 (N_17,In_527,In_466);
and U18 (N_18,In_1786,In_2140);
nor U19 (N_19,In_2472,In_2309);
xor U20 (N_20,In_982,In_2231);
nand U21 (N_21,In_1031,In_1708);
or U22 (N_22,In_1849,In_2135);
or U23 (N_23,In_2311,In_330);
nor U24 (N_24,In_254,In_1736);
xnor U25 (N_25,In_1930,In_553);
nand U26 (N_26,In_1575,In_931);
and U27 (N_27,In_994,In_162);
or U28 (N_28,In_194,In_2131);
nand U29 (N_29,In_1005,In_185);
and U30 (N_30,In_317,In_1288);
and U31 (N_31,In_1257,In_2144);
and U32 (N_32,In_2425,In_963);
or U33 (N_33,In_1871,In_1538);
nor U34 (N_34,In_1417,In_2401);
and U35 (N_35,In_1946,In_643);
and U36 (N_36,In_2107,In_1298);
and U37 (N_37,In_690,In_1489);
or U38 (N_38,In_1048,In_838);
nand U39 (N_39,In_1848,In_349);
and U40 (N_40,In_2111,In_993);
nand U41 (N_41,In_1093,In_2319);
or U42 (N_42,In_2117,In_2352);
nand U43 (N_43,In_981,In_948);
nor U44 (N_44,In_1690,In_540);
or U45 (N_45,In_1651,In_1255);
xnor U46 (N_46,In_1442,In_1509);
and U47 (N_47,In_112,In_1380);
and U48 (N_48,In_2156,In_1642);
nor U49 (N_49,In_18,In_1078);
xor U50 (N_50,In_2400,In_2226);
or U51 (N_51,In_915,In_2330);
xor U52 (N_52,In_1394,In_2478);
nor U53 (N_53,In_140,In_1129);
or U54 (N_54,In_1890,In_150);
xor U55 (N_55,In_2076,In_1443);
nor U56 (N_56,In_1504,In_1390);
nand U57 (N_57,In_262,In_546);
xnor U58 (N_58,In_2381,In_344);
xnor U59 (N_59,In_2146,In_1604);
or U60 (N_60,In_2353,In_1987);
and U61 (N_61,In_1344,In_1090);
and U62 (N_62,In_312,In_1416);
nand U63 (N_63,In_377,In_955);
xor U64 (N_64,In_280,In_737);
xor U65 (N_65,In_2051,In_1198);
xnor U66 (N_66,In_2260,In_1688);
or U67 (N_67,In_1258,In_927);
and U68 (N_68,In_2211,In_106);
and U69 (N_69,In_2181,In_1364);
xor U70 (N_70,In_2449,In_2093);
nand U71 (N_71,In_2245,In_2494);
and U72 (N_72,In_1401,In_2023);
nand U73 (N_73,In_2265,In_249);
nor U74 (N_74,In_1307,In_157);
or U75 (N_75,In_1217,In_677);
or U76 (N_76,In_1084,In_14);
and U77 (N_77,In_85,In_1350);
and U78 (N_78,In_1044,In_214);
and U79 (N_79,In_2468,In_769);
or U80 (N_80,In_2394,In_347);
nand U81 (N_81,In_1784,In_61);
nor U82 (N_82,In_1154,In_1799);
xor U83 (N_83,In_841,In_1694);
or U84 (N_84,In_1679,In_4);
nand U85 (N_85,In_1334,In_324);
nor U86 (N_86,In_933,In_2099);
or U87 (N_87,In_901,In_2476);
and U88 (N_88,In_863,In_730);
nand U89 (N_89,In_1333,In_1527);
xnor U90 (N_90,In_1473,In_1850);
nor U91 (N_91,In_1451,In_1980);
nand U92 (N_92,In_1098,In_1389);
nor U93 (N_93,In_1900,In_232);
or U94 (N_94,In_2403,In_1347);
nor U95 (N_95,In_2000,In_726);
or U96 (N_96,In_289,In_1950);
nand U97 (N_97,In_1243,In_1211);
nor U98 (N_98,In_1181,In_154);
and U99 (N_99,In_44,In_938);
or U100 (N_100,In_1487,In_1052);
or U101 (N_101,In_1928,In_114);
xnor U102 (N_102,In_998,In_247);
and U103 (N_103,In_1471,In_2248);
or U104 (N_104,In_631,In_609);
and U105 (N_105,In_566,In_772);
nor U106 (N_106,In_1224,In_761);
and U107 (N_107,In_305,In_1810);
nor U108 (N_108,In_1660,In_2004);
and U109 (N_109,In_2047,In_868);
nor U110 (N_110,In_2233,In_241);
and U111 (N_111,In_1674,In_1858);
xnor U112 (N_112,In_2190,In_1220);
nand U113 (N_113,In_618,In_1362);
nand U114 (N_114,In_779,In_2488);
nor U115 (N_115,In_1329,In_717);
nor U116 (N_116,In_1226,In_1529);
and U117 (N_117,In_684,In_1103);
nor U118 (N_118,In_1826,In_1237);
and U119 (N_119,In_1601,In_1054);
nor U120 (N_120,In_1261,In_2081);
or U121 (N_121,In_34,In_2413);
and U122 (N_122,In_23,In_616);
xor U123 (N_123,In_745,In_1836);
nor U124 (N_124,In_485,In_1203);
nand U125 (N_125,In_2464,In_2218);
nand U126 (N_126,In_1139,In_2206);
or U127 (N_127,In_2049,In_1000);
and U128 (N_128,In_2274,In_445);
and U129 (N_129,In_207,In_339);
nor U130 (N_130,In_2219,In_768);
nand U131 (N_131,In_1917,In_143);
xnor U132 (N_132,In_607,In_854);
and U133 (N_133,In_1315,In_399);
nand U134 (N_134,In_222,In_288);
xnor U135 (N_135,In_2297,In_2487);
or U136 (N_136,In_65,In_1038);
nor U137 (N_137,In_2227,In_1359);
nor U138 (N_138,In_1309,In_1614);
xnor U139 (N_139,In_1147,In_2042);
and U140 (N_140,In_669,In_52);
nand U141 (N_141,In_1134,In_448);
nand U142 (N_142,In_56,In_2064);
xor U143 (N_143,In_754,In_1883);
xnor U144 (N_144,In_398,In_903);
and U145 (N_145,In_887,In_116);
nand U146 (N_146,In_2171,In_2044);
xnor U147 (N_147,In_1144,In_2402);
and U148 (N_148,In_1585,In_1322);
and U149 (N_149,In_469,In_1889);
nand U150 (N_150,In_1131,In_2175);
nand U151 (N_151,In_1841,In_316);
or U152 (N_152,In_800,In_1760);
nand U153 (N_153,In_2216,In_1812);
or U154 (N_154,In_96,In_1995);
xor U155 (N_155,In_453,In_235);
or U156 (N_156,In_464,In_115);
or U157 (N_157,In_2436,In_205);
and U158 (N_158,In_1214,In_1662);
nand U159 (N_159,In_728,In_889);
xnor U160 (N_160,In_1827,In_1375);
nor U161 (N_161,In_251,In_230);
or U162 (N_162,In_359,In_2496);
nor U163 (N_163,In_217,In_2054);
nor U164 (N_164,In_1639,In_1895);
nand U165 (N_165,In_1744,In_763);
or U166 (N_166,In_1748,In_2056);
or U167 (N_167,In_1764,In_844);
and U168 (N_168,In_952,In_2225);
nand U169 (N_169,In_1933,In_865);
nor U170 (N_170,In_1299,In_1548);
nor U171 (N_171,In_1046,In_1986);
or U172 (N_172,In_835,In_975);
nor U173 (N_173,In_1612,In_2183);
nor U174 (N_174,In_877,In_1379);
nor U175 (N_175,In_2253,In_2290);
or U176 (N_176,In_849,In_681);
nor U177 (N_177,In_379,In_1776);
nor U178 (N_178,In_389,In_2258);
or U179 (N_179,In_1017,In_2482);
xor U180 (N_180,In_965,In_1308);
nor U181 (N_181,In_1397,In_2307);
or U182 (N_182,In_110,In_2017);
nor U183 (N_183,In_287,In_492);
or U184 (N_184,In_1998,In_1608);
xor U185 (N_185,In_1778,In_170);
nor U186 (N_186,In_807,In_652);
xor U187 (N_187,In_1204,In_1292);
nor U188 (N_188,In_1482,In_519);
nor U189 (N_189,In_1837,In_1981);
nor U190 (N_190,In_1587,In_2424);
nor U191 (N_191,In_1043,In_2124);
and U192 (N_192,In_2396,In_1636);
nand U193 (N_193,In_163,In_93);
and U194 (N_194,In_1969,In_1781);
nand U195 (N_195,In_462,In_699);
or U196 (N_196,In_1263,In_174);
xnor U197 (N_197,In_480,In_2459);
xnor U198 (N_198,In_1285,In_1524);
or U199 (N_199,In_1453,In_2208);
nor U200 (N_200,In_2244,In_787);
or U201 (N_201,In_129,In_87);
and U202 (N_202,In_2439,In_1241);
or U203 (N_203,In_82,In_1627);
xor U204 (N_204,In_511,In_2278);
or U205 (N_205,In_897,In_1558);
nand U206 (N_206,In_2230,In_2318);
nor U207 (N_207,In_1256,In_525);
nand U208 (N_208,In_431,In_563);
xor U209 (N_209,In_1404,In_2103);
nor U210 (N_210,In_550,In_400);
xnor U211 (N_211,In_733,In_1954);
xor U212 (N_212,In_1644,In_294);
nand U213 (N_213,In_1065,In_1172);
or U214 (N_214,In_2059,In_1846);
or U215 (N_215,In_2463,In_1123);
nand U216 (N_216,In_1430,In_211);
nor U217 (N_217,In_1042,In_181);
or U218 (N_218,In_848,In_2006);
and U219 (N_219,In_1311,In_722);
and U220 (N_220,In_2087,In_2256);
nand U221 (N_221,In_2043,In_1097);
nand U222 (N_222,In_223,In_1068);
and U223 (N_223,In_1881,In_802);
nand U224 (N_224,In_1268,In_215);
xnor U225 (N_225,In_1686,In_506);
or U226 (N_226,In_995,In_266);
nand U227 (N_227,In_10,In_291);
or U228 (N_228,In_246,In_49);
nor U229 (N_229,In_752,In_689);
xor U230 (N_230,In_1654,In_2391);
xnor U231 (N_231,In_2327,In_2074);
and U232 (N_232,In_862,In_2378);
nand U233 (N_233,In_1165,In_583);
and U234 (N_234,In_1483,In_1768);
or U235 (N_235,In_128,In_300);
or U236 (N_236,In_1598,In_691);
xor U237 (N_237,In_1310,In_1354);
xor U238 (N_238,In_688,In_1272);
nor U239 (N_239,In_515,In_1032);
and U240 (N_240,In_1798,In_322);
nor U241 (N_241,In_176,In_813);
xor U242 (N_242,In_1029,In_554);
xor U243 (N_243,In_2423,In_1630);
and U244 (N_244,In_792,In_956);
or U245 (N_245,In_198,In_1689);
or U246 (N_246,In_259,In_1516);
and U247 (N_247,In_1728,In_1004);
nand U248 (N_248,In_449,In_1792);
nand U249 (N_249,In_496,In_188);
and U250 (N_250,In_1168,In_1425);
nand U251 (N_251,In_1982,In_1136);
nand U252 (N_252,In_33,In_1008);
xnor U253 (N_253,In_2287,In_636);
or U254 (N_254,In_2469,In_1515);
or U255 (N_255,In_869,In_447);
or U256 (N_256,In_307,In_135);
nand U257 (N_257,In_2426,In_909);
and U258 (N_258,In_94,In_2441);
xnor U259 (N_259,In_723,In_329);
xor U260 (N_260,In_1944,In_641);
xnor U261 (N_261,In_966,In_2055);
and U262 (N_262,In_1368,In_2161);
and U263 (N_263,In_560,In_2089);
nor U264 (N_264,In_2421,In_1905);
or U265 (N_265,In_2203,In_523);
nor U266 (N_266,In_53,In_1523);
or U267 (N_267,In_1794,In_2243);
xor U268 (N_268,In_1113,In_2357);
nor U269 (N_269,In_1891,In_1590);
and U270 (N_270,In_1929,In_634);
nand U271 (N_271,In_1703,In_2215);
and U272 (N_272,In_375,In_1740);
and U273 (N_273,In_1325,In_2384);
or U274 (N_274,In_1869,In_811);
or U275 (N_275,In_1,In_873);
and U276 (N_276,In_1185,In_1970);
xor U277 (N_277,In_1621,In_2165);
or U278 (N_278,In_713,In_73);
xnor U279 (N_279,In_893,In_576);
nand U280 (N_280,In_1875,In_1996);
and U281 (N_281,In_160,In_764);
nor U282 (N_282,In_2471,In_1749);
and U283 (N_283,In_444,In_1484);
or U284 (N_284,In_1437,In_2300);
nand U285 (N_285,In_961,In_46);
nand U286 (N_286,In_1475,In_1340);
nor U287 (N_287,In_72,In_192);
nor U288 (N_288,In_505,In_1872);
nor U289 (N_289,In_169,In_2027);
nand U290 (N_290,In_1420,In_881);
nand U291 (N_291,In_1106,In_700);
nand U292 (N_292,In_929,In_2363);
and U293 (N_293,In_1470,In_810);
and U294 (N_294,In_1695,In_286);
or U295 (N_295,In_120,In_1301);
nor U296 (N_296,In_979,In_2450);
and U297 (N_297,In_794,In_1545);
and U298 (N_298,In_99,In_1221);
xnor U299 (N_299,In_899,In_1559);
xor U300 (N_300,In_833,In_1312);
and U301 (N_301,In_142,In_1976);
and U302 (N_302,In_2143,In_1888);
xor U303 (N_303,In_2149,In_179);
or U304 (N_304,In_821,In_2429);
nand U305 (N_305,In_1336,In_1646);
xnor U306 (N_306,In_870,In_1045);
nand U307 (N_307,In_177,In_2343);
or U308 (N_308,In_1452,In_1159);
nor U309 (N_309,In_337,In_775);
nor U310 (N_310,In_1148,In_1153);
nand U311 (N_311,In_2362,In_663);
and U312 (N_312,In_1829,In_1035);
nand U313 (N_313,In_1990,In_1407);
nor U314 (N_314,In_415,In_1622);
nand U315 (N_315,In_2458,In_601);
nor U316 (N_316,In_107,In_478);
xnor U317 (N_317,In_650,In_595);
nand U318 (N_318,In_2210,In_315);
nand U319 (N_319,In_562,In_67);
and U320 (N_320,In_762,In_1015);
nor U321 (N_321,In_2164,In_1454);
xnor U322 (N_322,In_1745,In_2035);
nand U323 (N_323,In_1324,In_985);
nor U324 (N_324,In_209,In_408);
and U325 (N_325,In_1219,In_2142);
and U326 (N_326,In_486,In_1632);
xor U327 (N_327,In_2177,In_2479);
xnor U328 (N_328,In_2451,In_356);
xor U329 (N_329,In_2393,In_1266);
xor U330 (N_330,In_2337,In_543);
nand U331 (N_331,In_1076,In_1066);
xor U332 (N_332,In_101,In_1462);
or U333 (N_333,In_1025,In_1171);
and U334 (N_334,In_2323,In_1493);
or U335 (N_335,In_1719,In_2010);
xor U336 (N_336,In_2063,In_1867);
or U337 (N_337,In_1002,In_2024);
or U338 (N_338,In_670,In_2483);
nand U339 (N_339,In_1957,In_1857);
and U340 (N_340,In_2242,In_2303);
xor U341 (N_341,In_1478,In_2302);
nand U342 (N_342,In_1704,In_1244);
and U343 (N_343,In_959,In_1835);
nor U344 (N_344,In_591,In_2002);
or U345 (N_345,In_673,In_1318);
nand U346 (N_346,In_465,In_1876);
xor U347 (N_347,In_570,In_236);
or U348 (N_348,In_1761,In_210);
and U349 (N_349,In_796,In_1873);
nand U350 (N_350,In_653,In_1655);
nor U351 (N_351,In_123,In_1157);
nor U352 (N_352,In_2335,In_1556);
or U353 (N_353,In_50,In_2048);
or U354 (N_354,In_858,In_1819);
and U355 (N_355,In_1095,In_21);
xnor U356 (N_356,In_1591,In_1186);
and U357 (N_357,In_747,In_1967);
or U358 (N_358,In_1958,In_64);
and U359 (N_359,In_1787,In_654);
nand U360 (N_360,In_1723,In_417);
xor U361 (N_361,In_2058,In_1520);
and U362 (N_362,In_2345,In_362);
nand U363 (N_363,In_788,In_2014);
xnor U364 (N_364,In_917,In_86);
and U365 (N_365,In_750,In_2229);
xor U366 (N_366,In_2015,In_1135);
and U367 (N_367,In_1691,In_1376);
or U368 (N_368,In_2374,In_1817);
or U369 (N_369,In_2277,In_1856);
nor U370 (N_370,In_436,In_716);
and U371 (N_371,In_1641,In_144);
nand U372 (N_372,In_1729,In_103);
nand U373 (N_373,In_1128,In_2418);
nand U374 (N_374,In_1485,In_491);
or U375 (N_375,In_182,In_1822);
xor U376 (N_376,In_350,In_311);
and U377 (N_377,In_1193,In_1248);
and U378 (N_378,In_495,In_659);
nand U379 (N_379,In_1806,In_1433);
and U380 (N_380,In_1699,In_1977);
nand U381 (N_381,In_1964,In_1012);
xnor U382 (N_382,In_675,In_191);
nand U383 (N_383,In_850,In_2321);
nand U384 (N_384,In_735,In_647);
nand U385 (N_385,In_2016,In_1353);
or U386 (N_386,In_950,In_1206);
and U387 (N_387,In_1143,In_1349);
and U388 (N_388,In_1109,In_1233);
or U389 (N_389,In_1542,In_1789);
nor U390 (N_390,In_1326,In_1381);
nor U391 (N_391,In_878,In_1510);
nor U392 (N_392,In_1357,In_776);
or U393 (N_393,In_805,In_1146);
nor U394 (N_394,In_1907,In_949);
or U395 (N_395,In_1438,In_392);
and U396 (N_396,In_252,In_2470);
xor U397 (N_397,In_148,In_1293);
and U398 (N_398,In_1971,In_795);
or U399 (N_399,In_575,In_573);
and U400 (N_400,In_1501,In_474);
nor U401 (N_401,In_628,In_195);
xor U402 (N_402,In_1600,In_969);
nor U403 (N_403,In_204,In_2320);
xnor U404 (N_404,In_1595,In_271);
nor U405 (N_405,In_1251,In_299);
xnor U406 (N_406,In_490,In_1282);
nor U407 (N_407,In_2032,In_834);
and U408 (N_408,In_1274,In_388);
xnor U409 (N_409,In_2430,In_1974);
and U410 (N_410,In_2134,In_2091);
nand U411 (N_411,In_2288,In_1490);
or U412 (N_412,In_782,In_1586);
nand U413 (N_413,In_193,In_2174);
and U414 (N_414,In_1580,In_2326);
xnor U415 (N_415,In_1772,In_1560);
xnor U416 (N_416,In_310,In_2271);
and U417 (N_417,In_2263,In_2259);
or U418 (N_418,In_2261,In_1276);
xnor U419 (N_419,In_1180,In_2457);
nand U420 (N_420,In_1972,In_1184);
nor U421 (N_421,In_1155,In_798);
nor U422 (N_422,In_202,In_2067);
nand U423 (N_423,In_944,In_2433);
xor U424 (N_424,In_226,In_1124);
and U425 (N_425,In_1864,In_1993);
nand U426 (N_426,In_2061,In_612);
nand U427 (N_427,In_1528,In_1434);
or U428 (N_428,In_1339,In_2011);
nand U429 (N_429,In_2036,In_1137);
or U430 (N_430,In_1200,In_1303);
and U431 (N_431,In_672,In_567);
or U432 (N_432,In_2419,In_1975);
nor U433 (N_433,In_2185,In_1071);
xnor U434 (N_434,In_146,In_1242);
nand U435 (N_435,In_2028,In_1427);
or U436 (N_436,In_451,In_538);
nor U437 (N_437,In_853,In_2235);
nor U438 (N_438,In_1581,In_824);
xnor U439 (N_439,In_664,In_2347);
xor U440 (N_440,In_1297,In_1960);
or U441 (N_441,In_1223,In_2132);
xnor U442 (N_442,In_1435,In_978);
nand U443 (N_443,In_2493,In_648);
or U444 (N_444,In_791,In_81);
and U445 (N_445,In_1472,In_561);
and U446 (N_446,In_1887,In_1345);
and U447 (N_447,In_2399,In_421);
nand U448 (N_448,In_2198,In_345);
nand U449 (N_449,In_623,In_471);
nor U450 (N_450,In_704,In_393);
nand U451 (N_451,In_1110,In_827);
nand U452 (N_452,In_1733,In_1459);
and U453 (N_453,In_1141,In_1839);
nand U454 (N_454,In_2057,In_1814);
xnor U455 (N_455,In_2029,In_727);
nand U456 (N_456,In_113,In_31);
and U457 (N_457,In_1605,In_1774);
xnor U458 (N_458,In_1874,In_1860);
and U459 (N_459,In_602,In_1395);
nand U460 (N_460,In_912,In_2207);
nor U461 (N_461,In_79,In_166);
xor U462 (N_462,In_1447,In_517);
nand U463 (N_463,In_264,In_422);
nand U464 (N_464,In_1229,In_1003);
nor U465 (N_465,In_1685,In_977);
nor U466 (N_466,In_1105,In_1557);
nor U467 (N_467,In_2193,In_1369);
nand U468 (N_468,In_2166,In_1021);
xor U469 (N_469,In_1423,In_1321);
or U470 (N_470,In_1800,In_529);
xor U471 (N_471,In_1680,In_57);
xnor U472 (N_472,In_1592,In_964);
xor U473 (N_473,In_2349,In_1702);
xor U474 (N_474,In_971,In_828);
or U475 (N_475,In_342,In_1892);
nor U476 (N_476,In_1119,In_890);
nand U477 (N_477,In_147,In_907);
or U478 (N_478,In_401,In_2053);
and U479 (N_479,In_581,In_1488);
nor U480 (N_480,In_816,In_742);
or U481 (N_481,In_1080,In_1613);
or U482 (N_482,In_1968,In_233);
xor U483 (N_483,In_1941,In_1541);
and U484 (N_484,In_172,In_2112);
xor U485 (N_485,In_967,In_1295);
or U486 (N_486,In_698,In_1913);
nand U487 (N_487,In_1955,In_467);
nor U488 (N_488,In_2334,In_1101);
and U489 (N_489,In_2370,In_1777);
nor U490 (N_490,In_161,In_1116);
nor U491 (N_491,In_1626,In_1652);
or U492 (N_492,In_1666,In_657);
xnor U493 (N_493,In_2269,In_1610);
and U494 (N_494,In_411,In_1020);
and U495 (N_495,In_1973,In_725);
nor U496 (N_496,In_2444,In_168);
or U497 (N_497,In_229,In_2150);
nand U498 (N_498,In_171,In_666);
nand U499 (N_499,In_1196,In_942);
xor U500 (N_500,In_248,In_1028);
and U501 (N_501,In_1648,In_1419);
or U502 (N_502,In_333,In_2405);
and U503 (N_503,In_1717,In_1897);
or U504 (N_504,In_645,In_2408);
or U505 (N_505,In_441,In_845);
nand U506 (N_506,In_1951,In_277);
or U507 (N_507,In_76,In_124);
nand U508 (N_508,In_744,In_856);
nand U509 (N_509,In_2246,In_1640);
or U510 (N_510,In_1578,In_1809);
nor U511 (N_511,In_1681,In_403);
nor U512 (N_512,In_766,In_658);
nand U513 (N_513,In_443,In_1413);
and U514 (N_514,In_1683,In_313);
and U515 (N_515,In_1534,In_139);
nand U516 (N_516,In_2018,In_224);
nor U517 (N_517,In_423,In_397);
xnor U518 (N_518,In_1331,In_2160);
xor U519 (N_519,In_1619,In_2404);
nand U520 (N_520,In_1834,In_285);
or U521 (N_521,In_1563,In_1985);
xnor U522 (N_522,In_559,In_1161);
xor U523 (N_523,In_751,In_2033);
or U524 (N_524,In_270,In_428);
and U525 (N_525,In_1479,In_173);
or U526 (N_526,In_1716,In_1752);
nand U527 (N_527,In_2434,In_303);
nor U528 (N_528,In_1920,In_829);
nand U529 (N_529,In_904,In_1718);
and U530 (N_530,In_2358,In_2308);
nand U531 (N_531,In_1676,In_1351);
and U532 (N_532,In_2392,In_2420);
and U533 (N_533,In_1593,In_2209);
xor U534 (N_534,In_674,In_1631);
or U535 (N_535,In_2455,In_2191);
nand U536 (N_536,In_1227,In_1396);
and U537 (N_537,In_1802,In_136);
nand U538 (N_538,In_360,In_1073);
and U539 (N_539,In_2456,In_1894);
and U540 (N_540,In_1818,In_30);
xor U541 (N_541,In_2499,In_1300);
nor U542 (N_542,In_804,In_578);
or U543 (N_543,In_258,In_420);
nor U544 (N_544,In_1306,In_557);
or U545 (N_545,In_1576,In_749);
nor U546 (N_546,In_820,In_697);
or U547 (N_547,In_635,In_1500);
and U548 (N_548,In_551,In_925);
nand U549 (N_549,In_2069,In_22);
or U550 (N_550,In_340,In_785);
nor U551 (N_551,In_472,In_973);
nand U552 (N_552,In_1664,In_1816);
or U553 (N_553,In_58,In_1305);
xnor U554 (N_554,In_2477,In_1378);
nand U555 (N_555,In_1464,In_613);
nand U556 (N_556,In_2254,In_2212);
and U557 (N_557,In_1770,In_1507);
nor U558 (N_558,In_2324,In_88);
or U559 (N_559,In_1290,In_2008);
nand U560 (N_560,In_1743,In_2025);
nand U561 (N_561,In_1304,In_1899);
or U562 (N_562,In_2003,In_319);
and U563 (N_563,In_284,In_59);
nor U564 (N_564,In_918,In_983);
nand U565 (N_565,In_2092,In_1606);
nand U566 (N_566,In_19,In_2090);
and U567 (N_567,In_1014,In_1201);
nor U568 (N_568,In_2312,In_535);
or U569 (N_569,In_1893,In_2298);
nor U570 (N_570,In_274,In_908);
xnor U571 (N_571,In_1497,In_2179);
nand U572 (N_572,In_1700,In_1034);
xnor U573 (N_573,In_1584,In_260);
nor U574 (N_574,In_2096,In_1953);
or U575 (N_575,In_2336,In_1176);
nand U576 (N_576,In_7,In_2372);
xnor U577 (N_577,In_2240,In_2104);
and U578 (N_578,In_1863,In_66);
xnor U579 (N_579,In_2250,In_1440);
and U580 (N_580,In_1030,In_2196);
xor U581 (N_581,In_1205,In_138);
nor U582 (N_582,In_710,In_1589);
nand U583 (N_583,In_926,In_639);
and U584 (N_584,In_2406,In_2490);
nor U585 (N_585,In_651,In_598);
xnor U586 (N_586,In_1934,In_861);
nor U587 (N_587,In_1579,In_895);
or U588 (N_588,In_1079,In_1988);
nor U589 (N_589,In_2158,In_2346);
and U590 (N_590,In_1855,In_493);
xor U591 (N_591,In_1117,In_846);
nor U592 (N_592,In_649,In_1550);
or U593 (N_593,In_26,In_45);
nor U594 (N_594,In_999,In_2109);
nor U595 (N_595,In_793,In_361);
nand U596 (N_596,In_427,In_2079);
nor U597 (N_597,In_1943,In_433);
xor U598 (N_598,In_1554,In_531);
or U599 (N_599,In_1426,In_1705);
and U600 (N_600,In_282,In_801);
or U601 (N_601,In_781,In_592);
xnor U602 (N_602,In_1094,In_2340);
xor U603 (N_603,In_1912,In_624);
nor U604 (N_604,In_2446,In_1118);
or U605 (N_605,In_1677,In_468);
or U606 (N_606,In_263,In_2106);
and U607 (N_607,In_92,In_152);
xor U608 (N_608,In_131,In_1444);
and U609 (N_609,In_2178,In_2162);
or U610 (N_610,In_1253,In_257);
xor U611 (N_611,In_2492,In_518);
and U612 (N_612,In_218,In_323);
nor U613 (N_613,In_1635,In_178);
xor U614 (N_614,In_2202,In_1492);
nand U615 (N_615,In_1387,In_2338);
and U616 (N_616,In_1361,In_1757);
nor U617 (N_617,In_706,In_1788);
and U618 (N_618,In_1474,In_682);
xor U619 (N_619,In_2368,In_565);
or U620 (N_620,In_2145,In_2122);
or U621 (N_621,In_1187,In_109);
or U622 (N_622,In_424,In_2125);
nand U623 (N_623,In_1517,In_11);
and U624 (N_624,In_589,In_2118);
xnor U625 (N_625,In_332,In_711);
and U626 (N_626,In_1026,In_499);
nor U627 (N_627,In_1284,In_290);
or U628 (N_628,In_552,In_1278);
or U629 (N_629,In_2197,In_2169);
and U630 (N_630,In_216,In_2331);
and U631 (N_631,In_1178,In_2447);
nand U632 (N_632,In_376,In_455);
or U633 (N_633,In_2031,In_857);
and U634 (N_634,In_919,In_326);
or U635 (N_635,In_442,In_1793);
or U636 (N_636,In_1352,In_1795);
and U637 (N_637,In_2491,In_1273);
or U638 (N_638,In_2344,In_1130);
nor U639 (N_639,In_1328,In_2);
nand U640 (N_640,In_1840,In_1179);
or U641 (N_641,In_71,In_888);
nand U642 (N_642,In_1568,In_225);
or U643 (N_643,In_1138,In_364);
nand U644 (N_644,In_2097,In_8);
and U645 (N_645,In_189,In_279);
or U646 (N_646,In_1932,In_1216);
and U647 (N_647,In_456,In_619);
and U648 (N_648,In_871,In_1763);
nor U649 (N_649,In_549,In_611);
or U650 (N_650,In_1830,In_1089);
and U651 (N_651,In_1682,In_2021);
and U652 (N_652,In_1410,In_1072);
nor U653 (N_653,In_341,In_1916);
xor U654 (N_654,In_2382,In_1661);
or U655 (N_655,In_2282,In_708);
xnor U656 (N_656,In_2050,In_593);
or U657 (N_657,In_1085,In_692);
and U658 (N_658,In_1024,In_2005);
and U659 (N_659,In_1773,In_814);
and U660 (N_660,In_1825,In_1561);
nand U661 (N_661,In_1663,In_366);
nor U662 (N_662,In_1540,In_1270);
xor U663 (N_663,In_1152,In_2084);
nand U664 (N_664,In_920,In_2388);
or U665 (N_665,In_2101,In_1195);
and U666 (N_666,In_1486,In_2237);
and U667 (N_667,In_15,In_2199);
or U668 (N_668,In_1163,In_1966);
xnor U669 (N_669,In_928,In_1617);
xnor U670 (N_670,In_2443,In_386);
or U671 (N_671,In_1649,In_268);
xnor U672 (N_672,In_1225,In_201);
xor U673 (N_673,In_1519,In_1922);
or U674 (N_674,In_2128,In_859);
nor U675 (N_675,In_2116,In_736);
nand U676 (N_676,In_537,In_1463);
or U677 (N_677,In_1174,In_686);
and U678 (N_678,In_1316,In_2385);
and U679 (N_679,In_1370,In_1552);
nor U680 (N_680,In_2264,In_1096);
and U681 (N_681,In_127,In_1449);
and U682 (N_682,In_1607,In_1623);
and U683 (N_683,In_2275,In_1235);
and U684 (N_684,In_991,In_1936);
nor U685 (N_685,In_1518,In_213);
xnor U686 (N_686,In_1197,In_2022);
and U687 (N_687,In_585,In_2442);
or U688 (N_688,In_1832,In_2377);
xnor U689 (N_689,In_1687,In_383);
nand U690 (N_690,In_1750,In_2306);
nand U691 (N_691,In_396,In_228);
and U692 (N_692,In_75,In_42);
xnor U693 (N_693,In_1865,In_2313);
nor U694 (N_694,In_1983,In_1570);
or U695 (N_695,In_1150,In_1126);
nand U696 (N_696,In_348,In_2126);
nand U697 (N_697,In_1040,In_2461);
nand U698 (N_698,In_1252,In_867);
nand U699 (N_699,In_1758,In_134);
and U700 (N_700,In_1269,In_1823);
xor U701 (N_701,In_1908,In_1693);
xnor U702 (N_702,In_740,In_1919);
nor U703 (N_703,In_604,In_1461);
and U704 (N_704,In_302,In_1314);
xor U705 (N_705,In_539,In_1707);
or U706 (N_706,In_378,In_461);
nor U707 (N_707,In_1939,In_1037);
nor U708 (N_708,In_632,In_1780);
xor U709 (N_709,In_1108,In_855);
or U710 (N_710,In_1537,In_864);
and U711 (N_711,In_167,In_434);
xnor U712 (N_712,In_958,In_121);
nand U713 (N_713,In_656,In_1533);
xnor U714 (N_714,In_2266,In_267);
or U715 (N_715,In_2348,In_1208);
nor U716 (N_716,In_2078,In_2155);
and U717 (N_717,In_1467,In_2296);
xor U718 (N_718,In_2220,In_524);
nor U719 (N_719,In_1102,In_1731);
nand U720 (N_720,In_874,In_1246);
xor U721 (N_721,In_1979,In_826);
and U722 (N_722,In_2082,In_482);
nor U723 (N_723,In_118,In_2108);
nand U724 (N_724,In_2034,In_1019);
and U725 (N_725,In_1280,In_2141);
nor U726 (N_726,In_295,In_1289);
nand U727 (N_727,In_1553,In_2083);
and U728 (N_728,In_614,In_2234);
and U729 (N_729,In_1843,In_1259);
or U730 (N_730,In_402,In_701);
or U731 (N_731,In_2276,In_1247);
xor U732 (N_732,In_2437,In_1572);
nand U733 (N_733,In_2428,In_1514);
nand U734 (N_734,In_1111,In_665);
or U735 (N_735,In_1460,In_945);
or U736 (N_736,In_1373,In_440);
nor U737 (N_737,In_2012,In_1701);
xor U738 (N_738,In_812,In_2257);
nand U739 (N_739,In_2085,In_885);
or U740 (N_740,In_1525,In_584);
nor U741 (N_741,In_622,In_54);
nand U742 (N_742,In_2273,In_789);
and U743 (N_743,In_272,In_1759);
or U744 (N_744,In_1665,In_429);
and U745 (N_745,In_715,In_62);
and U746 (N_746,In_2342,In_1360);
or U747 (N_747,In_2262,In_1064);
nor U748 (N_748,In_1597,In_321);
or U749 (N_749,In_2038,In_1755);
or U750 (N_750,In_685,In_1050);
or U751 (N_751,In_1320,In_2285);
nand U752 (N_752,In_1386,In_1061);
or U753 (N_753,In_1532,In_1901);
and U754 (N_754,In_1730,In_406);
or U755 (N_755,In_866,In_921);
and U756 (N_756,In_521,In_817);
xnor U757 (N_757,In_1711,In_501);
and U758 (N_758,In_186,In_2293);
or U759 (N_759,In_68,In_1742);
or U760 (N_760,In_1726,In_916);
xnor U761 (N_761,In_1927,In_1053);
or U762 (N_762,In_368,In_1721);
and U763 (N_763,In_1151,In_2194);
nor U764 (N_764,In_2380,In_996);
xor U765 (N_765,In_640,In_1965);
nor U766 (N_766,In_2188,In_1720);
nand U767 (N_767,In_77,In_569);
nand U768 (N_768,In_2114,In_1009);
nor U769 (N_769,In_6,In_1455);
nand U770 (N_770,In_1657,In_1115);
and U771 (N_771,In_2214,In_780);
nand U772 (N_772,In_1880,In_1959);
xor U773 (N_773,In_2100,In_1997);
nor U774 (N_774,In_1886,In_293);
nor U775 (N_775,In_2497,In_1747);
and U776 (N_776,In_1565,In_1480);
or U777 (N_777,In_2473,In_1678);
nand U778 (N_778,In_1767,In_1450);
nor U779 (N_779,In_1384,In_1808);
xor U780 (N_780,In_1599,In_1051);
xor U781 (N_781,In_1698,In_719);
nand U782 (N_782,In_633,In_1820);
and U783 (N_783,In_2291,In_297);
and U784 (N_784,In_1275,In_133);
nor U785 (N_785,In_548,In_2445);
or U786 (N_786,In_1402,In_48);
xor U787 (N_787,In_2322,In_308);
or U788 (N_788,In_1801,In_439);
nor U789 (N_789,In_2030,In_1712);
xnor U790 (N_790,In_1088,In_425);
and U791 (N_791,In_1813,In_1942);
xnor U792 (N_792,In_1060,In_1104);
and U793 (N_793,In_38,In_69);
nand U794 (N_794,In_2453,In_2105);
or U795 (N_795,In_513,In_63);
nor U796 (N_796,In_759,In_1495);
or U797 (N_797,In_837,In_497);
xnor U798 (N_798,In_1618,In_1338);
nor U799 (N_799,In_1033,In_1746);
xnor U800 (N_800,In_974,In_2238);
or U801 (N_801,In_1637,In_1232);
xor U802 (N_802,In_476,In_843);
and U803 (N_803,In_1409,In_627);
nand U804 (N_804,In_5,In_2241);
nand U805 (N_805,In_487,In_1505);
nor U806 (N_806,In_1611,In_1160);
xor U807 (N_807,In_603,In_1625);
and U808 (N_808,In_2037,In_1805);
or U809 (N_809,In_104,In_283);
nor U810 (N_810,In_1083,In_579);
nor U811 (N_811,In_1771,In_158);
and U812 (N_812,In_1457,In_1769);
and U813 (N_813,In_947,In_1175);
nand U814 (N_814,In_2375,In_2485);
nor U815 (N_815,In_2041,In_1335);
xnor U816 (N_816,In_1086,In_1866);
nand U817 (N_817,In_1170,In_564);
and U818 (N_818,In_2325,In_183);
or U819 (N_819,In_40,In_1112);
xor U820 (N_820,In_80,In_1218);
and U821 (N_821,In_1082,In_1188);
and U822 (N_822,In_125,In_790);
nor U823 (N_823,In_338,In_1710);
or U824 (N_824,In_292,In_234);
and U825 (N_825,In_2376,In_1725);
or U826 (N_826,In_898,In_599);
or U827 (N_827,In_1481,In_2170);
xnor U828 (N_828,In_1062,In_1190);
nor U829 (N_829,In_678,In_494);
or U830 (N_830,In_1670,In_1935);
and U831 (N_831,In_2184,In_1429);
nor U832 (N_832,In_78,In_32);
and U833 (N_833,In_799,In_2452);
nand U834 (N_834,In_1363,In_1992);
xor U835 (N_835,In_318,In_438);
nor U836 (N_836,In_1671,In_2026);
nor U837 (N_837,In_102,In_597);
or U838 (N_838,In_84,In_774);
xnor U839 (N_839,In_1628,In_724);
xnor U840 (N_840,In_2071,In_2232);
xor U841 (N_841,In_1807,In_1001);
and U842 (N_842,In_477,In_1715);
xnor U843 (N_843,In_164,In_36);
and U844 (N_844,In_1183,In_2039);
nand U845 (N_845,In_1709,In_2486);
xor U846 (N_846,In_2127,In_1194);
and U847 (N_847,In_2075,In_90);
nand U848 (N_848,In_1569,In_2440);
and U849 (N_849,In_1797,In_1739);
nor U850 (N_850,In_896,In_2466);
or U851 (N_851,In_668,In_1191);
xnor U852 (N_852,In_2065,In_2431);
nand U853 (N_853,In_528,In_739);
nor U854 (N_854,In_346,In_1779);
nor U855 (N_855,In_1367,In_2186);
nor U856 (N_856,In_394,In_2379);
or U857 (N_857,In_43,In_556);
or U858 (N_858,In_1222,In_1469);
xor U859 (N_859,In_1456,In_1100);
and U860 (N_860,In_2139,In_1697);
xor U861 (N_861,In_369,In_363);
nand U862 (N_862,In_1653,In_243);
xnor U863 (N_863,In_530,In_296);
nor U864 (N_864,In_1099,In_91);
xnor U865 (N_865,In_968,In_1114);
xnor U866 (N_866,In_765,In_237);
nand U867 (N_867,In_309,In_1087);
nand U868 (N_868,In_1911,In_534);
xnor U869 (N_869,In_2310,In_240);
nand U870 (N_870,In_2438,In_60);
xor U871 (N_871,In_1041,In_367);
and U872 (N_872,In_507,In_55);
or U873 (N_873,In_1945,In_1371);
or U874 (N_874,In_479,In_1667);
xor U875 (N_875,In_1164,In_414);
and U876 (N_876,In_1016,In_2355);
nand U877 (N_877,In_2329,In_1783);
and U878 (N_878,In_197,In_930);
xnor U879 (N_879,In_2136,In_1878);
and U880 (N_880,In_1342,In_2173);
nand U881 (N_881,In_2072,In_404);
xnor U882 (N_882,In_1879,In_741);
and U883 (N_883,In_880,In_1782);
xor U884 (N_884,In_12,In_910);
or U885 (N_885,In_1543,In_1313);
or U886 (N_886,In_734,In_1790);
and U887 (N_887,In_1399,In_2270);
xor U888 (N_888,In_1156,In_2339);
nor U889 (N_889,In_2317,In_2094);
or U890 (N_890,In_1948,In_1140);
nand U891 (N_891,In_2119,In_1431);
xor U892 (N_892,In_51,In_1392);
or U893 (N_893,In_1526,In_2247);
and U894 (N_894,In_2066,In_2295);
and U895 (N_895,In_1714,In_541);
nor U896 (N_896,In_255,In_29);
and U897 (N_897,In_1279,In_1120);
and U898 (N_898,In_1938,In_1735);
or U899 (N_899,In_932,In_391);
or U900 (N_900,In_1262,In_488);
nor U901 (N_901,In_1650,In_1925);
xor U902 (N_902,In_2110,In_2286);
or U903 (N_903,In_514,In_988);
nor U904 (N_904,In_902,In_703);
xor U905 (N_905,In_924,In_165);
nor U906 (N_906,In_809,In_145);
xnor U907 (N_907,In_1398,In_2407);
nor U908 (N_908,In_2304,In_395);
nor U909 (N_909,In_1281,In_1348);
xnor U910 (N_910,In_1766,In_1441);
and U911 (N_911,In_1465,In_757);
xnor U912 (N_912,In_1238,In_696);
xor U913 (N_913,In_662,In_2060);
xnor U914 (N_914,In_1006,In_1978);
or U915 (N_915,In_387,In_2223);
xnor U916 (N_916,In_1287,In_629);
or U917 (N_917,In_1209,In_637);
nand U918 (N_918,In_732,In_1994);
or U919 (N_919,In_1991,In_276);
xor U920 (N_920,In_784,In_2159);
nor U921 (N_921,In_1291,In_2138);
nand U922 (N_922,In_939,In_2480);
xor U923 (N_923,In_526,In_1791);
and U924 (N_924,In_2095,In_508);
xnor U925 (N_925,In_783,In_555);
or U926 (N_926,In_2020,In_646);
or U927 (N_927,In_1506,In_2432);
nand U928 (N_928,In_2268,In_797);
nor U929 (N_929,In_1374,In_1924);
nand U930 (N_930,In_1499,In_1265);
xnor U931 (N_931,In_1811,In_1672);
and U932 (N_932,In_2395,In_1634);
and U933 (N_933,In_2294,In_2369);
and U934 (N_934,In_460,In_1508);
and U935 (N_935,In_2484,In_1323);
or U936 (N_936,In_1713,In_1458);
xor U937 (N_937,In_1999,In_2390);
or U938 (N_938,In_2373,In_1166);
nand U939 (N_939,In_1624,In_306);
or U940 (N_940,In_199,In_1077);
xnor U941 (N_941,In_382,In_2387);
and U942 (N_942,In_437,In_1121);
nor U943 (N_943,In_1940,In_2204);
xnor U944 (N_944,In_906,In_2279);
or U945 (N_945,In_1915,In_1902);
and U946 (N_946,In_2176,In_1330);
nand U947 (N_947,In_2200,In_304);
or U948 (N_948,In_760,In_137);
nand U949 (N_949,In_2086,In_1842);
xnor U950 (N_950,In_384,In_1754);
nand U951 (N_951,In_1127,In_1596);
nand U952 (N_952,In_660,In_1055);
or U953 (N_953,In_2153,In_1264);
and U954 (N_954,In_2070,In_770);
or U955 (N_955,In_2180,In_327);
or U956 (N_956,In_1271,In_1914);
and U957 (N_957,In_694,In_105);
nor U958 (N_958,In_1013,In_936);
nor U959 (N_959,In_2130,In_615);
and U960 (N_960,In_2427,In_851);
xnor U961 (N_961,In_588,In_1844);
xnor U962 (N_962,In_2213,In_301);
or U963 (N_963,In_314,In_335);
or U964 (N_964,In_590,In_1962);
nand U965 (N_965,In_1414,In_923);
nand U966 (N_966,In_231,In_1851);
nand U967 (N_967,In_1877,In_2462);
nor U968 (N_968,In_1522,In_244);
nor U969 (N_969,In_2046,In_2366);
nand U970 (N_970,In_1796,In_17);
and U971 (N_971,In_758,In_2217);
nand U972 (N_972,In_1296,In_1403);
and U973 (N_973,In_1468,In_1910);
xor U974 (N_974,In_1904,In_1854);
xor U975 (N_975,In_1337,In_1358);
or U976 (N_976,In_151,In_2172);
and U977 (N_977,In_1210,In_2351);
and U978 (N_978,In_238,In_1067);
nor U979 (N_979,In_884,In_1566);
nor U980 (N_980,In_940,In_620);
or U981 (N_981,In_1762,In_281);
nand U982 (N_982,In_2009,In_1833);
or U983 (N_983,In_126,In_2416);
xor U984 (N_984,In_385,In_1609);
and U985 (N_985,In_1885,In_1388);
and U986 (N_986,In_343,In_1861);
nor U987 (N_987,In_221,In_1847);
xor U988 (N_988,In_2148,In_1056);
and U989 (N_989,In_1544,In_577);
nor U990 (N_990,In_1250,In_2163);
nor U991 (N_991,In_2062,In_457);
xnor U992 (N_992,In_1477,In_960);
xor U993 (N_993,In_1133,In_1207);
xor U994 (N_994,In_876,In_712);
nand U995 (N_995,In_1984,In_2467);
nor U996 (N_996,In_1853,In_1643);
or U997 (N_997,In_1405,In_1446);
nand U998 (N_998,In_2474,In_671);
and U999 (N_999,In_1961,In_432);
nor U1000 (N_1000,In_1332,In_1785);
nand U1001 (N_1001,In_1884,In_606);
xnor U1002 (N_1002,In_1421,In_98);
nand U1003 (N_1003,In_1845,In_2102);
and U1004 (N_1004,In_1852,In_1023);
nor U1005 (N_1005,In_1732,In_1937);
xor U1006 (N_1006,In_1063,In_473);
or U1007 (N_1007,In_587,In_605);
and U1008 (N_1008,In_27,In_358);
xnor U1009 (N_1009,In_2221,In_803);
or U1010 (N_1010,In_512,In_594);
or U1011 (N_1011,In_2187,In_117);
xnor U1012 (N_1012,In_3,In_1132);
nand U1013 (N_1013,In_502,In_2272);
nand U1014 (N_1014,In_1059,In_1503);
or U1015 (N_1015,In_1070,In_2397);
nand U1016 (N_1016,In_1267,In_1418);
nor U1017 (N_1017,In_219,In_2341);
and U1018 (N_1018,In_2314,In_498);
nor U1019 (N_1019,In_1751,In_353);
xnor U1020 (N_1020,In_509,In_1149);
or U1021 (N_1021,In_693,In_2411);
xor U1022 (N_1022,In_1828,In_2489);
nand U1023 (N_1023,In_984,In_155);
xnor U1024 (N_1024,In_334,In_822);
or U1025 (N_1025,In_815,In_269);
and U1026 (N_1026,In_1007,In_2098);
nand U1027 (N_1027,In_1949,In_1393);
nor U1028 (N_1028,In_187,In_1466);
nor U1029 (N_1029,In_1602,In_1432);
and U1030 (N_1030,In_1022,In_558);
and U1031 (N_1031,In_2195,In_2077);
and U1032 (N_1032,In_1400,In_2201);
or U1033 (N_1033,In_2359,In_2435);
nand U1034 (N_1034,In_913,In_1213);
and U1035 (N_1035,In_220,In_1675);
and U1036 (N_1036,In_2073,In_419);
xnor U1037 (N_1037,In_1724,In_644);
and U1038 (N_1038,In_987,In_1753);
and U1039 (N_1039,In_1365,In_1722);
or U1040 (N_1040,In_1535,In_2409);
nor U1041 (N_1041,In_755,In_568);
nor U1042 (N_1042,In_542,In_1018);
xor U1043 (N_1043,In_2398,In_2133);
nand U1044 (N_1044,In_1327,In_250);
and U1045 (N_1045,In_1476,In_2365);
xor U1046 (N_1046,In_1239,In_1122);
xor U1047 (N_1047,In_830,In_980);
nand U1048 (N_1048,In_2386,In_695);
xnor U1049 (N_1049,In_2333,In_2013);
nand U1050 (N_1050,In_1531,In_1428);
nor U1051 (N_1051,In_2052,In_1821);
and U1052 (N_1052,In_2465,In_2154);
xnor U1053 (N_1053,In_1074,In_1511);
xor U1054 (N_1054,In_922,In_1734);
or U1055 (N_1055,In_47,In_522);
or U1056 (N_1056,In_894,In_1727);
nand U1057 (N_1057,In_879,In_997);
xor U1058 (N_1058,In_954,In_1075);
or U1059 (N_1059,In_336,In_676);
xor U1060 (N_1060,In_1539,In_1202);
xnor U1061 (N_1061,In_1756,In_532);
xnor U1062 (N_1062,In_16,In_1696);
and U1063 (N_1063,In_1228,In_905);
xor U1064 (N_1064,In_2222,In_2167);
or U1065 (N_1065,In_545,In_1921);
nand U1066 (N_1066,In_1947,In_184);
nand U1067 (N_1067,In_1571,In_132);
and U1068 (N_1068,In_986,In_1870);
nor U1069 (N_1069,In_108,In_331);
nand U1070 (N_1070,In_2354,In_806);
nor U1071 (N_1071,In_705,In_351);
nand U1072 (N_1072,In_610,In_1377);
or U1073 (N_1073,In_261,In_1952);
xnor U1074 (N_1074,In_2389,In_1831);
xor U1075 (N_1075,In_1125,In_1346);
nand U1076 (N_1076,In_2289,In_621);
xnor U1077 (N_1077,In_1562,In_582);
or U1078 (N_1078,In_718,In_1277);
or U1079 (N_1079,In_156,In_1107);
or U1080 (N_1080,In_2417,In_24);
nor U1081 (N_1081,In_1177,In_2151);
nand U1082 (N_1082,In_454,In_600);
and U1083 (N_1083,In_808,In_2137);
nand U1084 (N_1084,In_2182,In_972);
nand U1085 (N_1085,In_1356,In_1838);
nor U1086 (N_1086,In_687,In_2356);
xor U1087 (N_1087,In_1372,In_452);
and U1088 (N_1088,In_1658,In_1573);
and U1089 (N_1089,In_771,In_510);
and U1090 (N_1090,In_1931,In_1260);
nand U1091 (N_1091,In_2364,In_95);
or U1092 (N_1092,In_1234,In_839);
and U1093 (N_1093,In_818,In_840);
nor U1094 (N_1094,In_1765,In_970);
xor U1095 (N_1095,In_83,In_357);
and U1096 (N_1096,In_74,In_416);
and U1097 (N_1097,In_1903,In_1512);
xor U1098 (N_1098,In_2332,In_638);
nor U1099 (N_1099,In_380,In_1659);
and U1100 (N_1100,In_122,In_1286);
or U1101 (N_1101,In_503,In_1036);
nor U1102 (N_1102,In_130,In_1249);
nor U1103 (N_1103,In_1192,In_2007);
nand U1104 (N_1104,In_1896,In_731);
xnor U1105 (N_1105,In_245,In_667);
or U1106 (N_1106,In_410,In_891);
xnor U1107 (N_1107,In_2205,In_500);
xor U1108 (N_1108,In_753,In_1513);
and U1109 (N_1109,In_1898,In_679);
or U1110 (N_1110,In_2460,In_1882);
and U1111 (N_1111,In_608,In_1366);
and U1112 (N_1112,In_2152,In_571);
nand U1113 (N_1113,In_900,In_1498);
and U1114 (N_1114,In_1092,In_1343);
or U1115 (N_1115,In_2305,In_175);
nor U1116 (N_1116,In_989,In_852);
and U1117 (N_1117,In_28,In_767);
nand U1118 (N_1118,In_990,In_435);
xor U1119 (N_1119,In_256,In_1167);
nor U1120 (N_1120,In_911,In_1382);
nor U1121 (N_1121,In_239,In_2189);
nand U1122 (N_1122,In_2316,In_934);
and U1123 (N_1123,In_1620,In_371);
and U1124 (N_1124,In_1245,In_1741);
xor U1125 (N_1125,In_1142,In_738);
and U1126 (N_1126,In_149,In_1804);
and U1127 (N_1127,In_1212,In_1319);
nand U1128 (N_1128,In_847,In_208);
or U1129 (N_1129,In_1594,In_1706);
nor U1130 (N_1130,In_580,In_957);
nand U1131 (N_1131,In_475,In_2410);
or U1132 (N_1132,In_489,In_1254);
xnor U1133 (N_1133,In_381,In_1496);
nand U1134 (N_1134,In_1956,In_265);
xor U1135 (N_1135,In_426,In_2255);
nor U1136 (N_1136,In_483,In_2328);
or U1137 (N_1137,In_547,In_372);
or U1138 (N_1138,In_1673,In_196);
or U1139 (N_1139,In_1011,In_680);
and U1140 (N_1140,In_1385,In_2123);
nand U1141 (N_1141,In_1549,In_273);
nor U1142 (N_1142,In_1638,In_875);
nand U1143 (N_1143,In_2236,In_1162);
nand U1144 (N_1144,In_407,In_2481);
nor U1145 (N_1145,In_2249,In_9);
nor U1146 (N_1146,In_819,In_1408);
nand U1147 (N_1147,In_203,In_1057);
xor U1148 (N_1148,In_1547,In_937);
and U1149 (N_1149,In_1411,In_2157);
nand U1150 (N_1150,In_773,In_872);
nand U1151 (N_1151,In_626,In_212);
and U1152 (N_1152,In_2475,In_1775);
or U1153 (N_1153,In_832,In_180);
xnor U1154 (N_1154,In_1603,In_1169);
xnor U1155 (N_1155,In_458,In_2315);
nand U1156 (N_1156,In_373,In_1502);
or U1157 (N_1157,In_355,In_1424);
nand U1158 (N_1158,In_119,In_1422);
or U1159 (N_1159,In_206,In_1551);
nor U1160 (N_1160,In_1656,In_446);
xor U1161 (N_1161,In_352,In_1491);
xor U1162 (N_1162,In_2299,In_2068);
and U1163 (N_1163,In_390,In_642);
nand U1164 (N_1164,In_2422,In_586);
and U1165 (N_1165,In_141,In_536);
xnor U1166 (N_1166,In_1738,In_1027);
and U1167 (N_1167,In_883,In_836);
and U1168 (N_1168,In_412,In_430);
xor U1169 (N_1169,In_1963,In_484);
nor U1170 (N_1170,In_1215,In_37);
and U1171 (N_1171,In_2454,In_2115);
nand U1172 (N_1172,In_882,In_190);
or U1173 (N_1173,In_1047,In_1824);
and U1174 (N_1174,In_2147,In_1145);
or U1175 (N_1175,In_1240,In_1294);
nand U1176 (N_1176,In_1049,In_574);
and U1177 (N_1177,In_1415,In_1633);
nand U1178 (N_1178,In_860,In_1564);
nor U1179 (N_1179,In_470,In_946);
xor U1180 (N_1180,In_13,In_625);
and U1181 (N_1181,In_630,In_365);
xnor U1182 (N_1182,In_298,In_481);
xor U1183 (N_1183,In_1494,In_743);
nor U1184 (N_1184,In_707,In_1536);
nand U1185 (N_1185,In_2284,In_572);
nor U1186 (N_1186,In_992,In_596);
and U1187 (N_1187,In_1317,In_111);
xor U1188 (N_1188,In_1989,In_943);
nand U1189 (N_1189,In_953,In_1616);
and U1190 (N_1190,In_1448,In_2292);
nor U1191 (N_1191,In_721,In_463);
xor U1192 (N_1192,In_2019,In_320);
and U1193 (N_1193,In_2367,In_533);
xor U1194 (N_1194,In_20,In_1406);
nor U1195 (N_1195,In_2251,In_842);
nand U1196 (N_1196,In_2113,In_413);
nor U1197 (N_1197,In_951,In_892);
nor U1198 (N_1198,In_778,In_2267);
or U1199 (N_1199,In_516,In_1684);
and U1200 (N_1200,In_1391,In_1645);
nor U1201 (N_1201,In_2228,In_1577);
and U1202 (N_1202,In_1668,In_2371);
xor U1203 (N_1203,In_1199,In_2495);
xnor U1204 (N_1204,In_2080,In_2224);
nand U1205 (N_1205,In_825,In_661);
xor U1206 (N_1206,In_1647,In_374);
nand U1207 (N_1207,In_1815,In_1283);
nand U1208 (N_1208,In_1182,In_1692);
nand U1209 (N_1209,In_39,In_278);
nand U1210 (N_1210,In_1567,In_325);
or U1211 (N_1211,In_1412,In_1439);
and U1212 (N_1212,In_25,In_328);
or U1213 (N_1213,In_2168,In_2301);
nand U1214 (N_1214,In_1230,In_2001);
nand U1215 (N_1215,In_200,In_1058);
xnor U1216 (N_1216,In_2281,In_941);
or U1217 (N_1217,In_409,In_748);
nand U1218 (N_1218,In_2360,In_786);
nor U1219 (N_1219,In_2040,In_1862);
or U1220 (N_1220,In_1355,In_2415);
nor U1221 (N_1221,In_746,In_97);
nand U1222 (N_1222,In_1669,In_370);
xnor U1223 (N_1223,In_823,In_1582);
nand U1224 (N_1224,In_1926,In_418);
xnor U1225 (N_1225,In_1546,In_2350);
nand U1226 (N_1226,In_89,In_2414);
nand U1227 (N_1227,In_520,In_702);
and U1228 (N_1228,In_831,In_2498);
nor U1229 (N_1229,In_2412,In_962);
nor U1230 (N_1230,In_1302,In_1909);
nand U1231 (N_1231,In_914,In_1583);
or U1232 (N_1232,In_41,In_617);
xnor U1233 (N_1233,In_1231,In_1521);
and U1234 (N_1234,In_2129,In_2088);
or U1235 (N_1235,In_1091,In_729);
and U1236 (N_1236,In_714,In_683);
xnor U1237 (N_1237,In_2192,In_935);
or U1238 (N_1238,In_777,In_242);
nor U1239 (N_1239,In_2361,In_35);
and U1240 (N_1240,In_1069,In_1868);
nand U1241 (N_1241,In_886,In_1906);
and U1242 (N_1242,In_1737,In_1445);
nand U1243 (N_1243,In_1173,In_153);
xor U1244 (N_1244,In_1010,In_354);
xnor U1245 (N_1245,In_0,In_450);
or U1246 (N_1246,In_544,In_756);
or U1247 (N_1247,In_2383,In_1629);
or U1248 (N_1248,In_1588,In_1923);
nand U1249 (N_1249,In_1236,In_1615);
nor U1250 (N_1250,In_1809,In_1556);
and U1251 (N_1251,In_283,In_2286);
nor U1252 (N_1252,In_691,In_2185);
xnor U1253 (N_1253,In_1375,In_2262);
nor U1254 (N_1254,In_540,In_1508);
xnor U1255 (N_1255,In_1613,In_1762);
xor U1256 (N_1256,In_34,In_416);
and U1257 (N_1257,In_1328,In_1059);
and U1258 (N_1258,In_207,In_144);
and U1259 (N_1259,In_836,In_2250);
xor U1260 (N_1260,In_1409,In_1174);
nand U1261 (N_1261,In_1962,In_1551);
nor U1262 (N_1262,In_935,In_1840);
nor U1263 (N_1263,In_664,In_2265);
and U1264 (N_1264,In_973,In_1263);
or U1265 (N_1265,In_175,In_1607);
xnor U1266 (N_1266,In_1009,In_1959);
nor U1267 (N_1267,In_2296,In_1209);
or U1268 (N_1268,In_1938,In_370);
nor U1269 (N_1269,In_2455,In_1977);
and U1270 (N_1270,In_902,In_2108);
xnor U1271 (N_1271,In_331,In_1842);
nand U1272 (N_1272,In_2210,In_1557);
nor U1273 (N_1273,In_1076,In_1356);
nand U1274 (N_1274,In_1936,In_278);
nor U1275 (N_1275,In_2451,In_1287);
xor U1276 (N_1276,In_1945,In_1085);
nand U1277 (N_1277,In_1070,In_2114);
and U1278 (N_1278,In_257,In_896);
and U1279 (N_1279,In_2128,In_1771);
nand U1280 (N_1280,In_137,In_1755);
or U1281 (N_1281,In_1493,In_2159);
xor U1282 (N_1282,In_2233,In_110);
nand U1283 (N_1283,In_39,In_1849);
nor U1284 (N_1284,In_911,In_1790);
or U1285 (N_1285,In_763,In_2029);
nand U1286 (N_1286,In_761,In_746);
and U1287 (N_1287,In_243,In_1936);
xor U1288 (N_1288,In_1199,In_1442);
nand U1289 (N_1289,In_1030,In_1762);
nand U1290 (N_1290,In_2446,In_1348);
xor U1291 (N_1291,In_1535,In_992);
nor U1292 (N_1292,In_420,In_1970);
xor U1293 (N_1293,In_1344,In_365);
or U1294 (N_1294,In_1854,In_1974);
or U1295 (N_1295,In_2020,In_253);
or U1296 (N_1296,In_359,In_1467);
xnor U1297 (N_1297,In_1448,In_713);
or U1298 (N_1298,In_680,In_400);
and U1299 (N_1299,In_534,In_264);
nor U1300 (N_1300,In_461,In_413);
nor U1301 (N_1301,In_1477,In_580);
xor U1302 (N_1302,In_889,In_409);
nor U1303 (N_1303,In_1385,In_1173);
nor U1304 (N_1304,In_1352,In_1613);
nand U1305 (N_1305,In_158,In_476);
xnor U1306 (N_1306,In_2221,In_2212);
nand U1307 (N_1307,In_2360,In_107);
xnor U1308 (N_1308,In_888,In_1983);
and U1309 (N_1309,In_330,In_2466);
xnor U1310 (N_1310,In_1204,In_914);
xnor U1311 (N_1311,In_1899,In_915);
nor U1312 (N_1312,In_773,In_1349);
nor U1313 (N_1313,In_1292,In_1694);
or U1314 (N_1314,In_1737,In_1033);
and U1315 (N_1315,In_109,In_1997);
nor U1316 (N_1316,In_1481,In_1883);
nor U1317 (N_1317,In_1620,In_650);
and U1318 (N_1318,In_1856,In_2339);
xnor U1319 (N_1319,In_2021,In_72);
xor U1320 (N_1320,In_2401,In_1069);
xnor U1321 (N_1321,In_644,In_2016);
and U1322 (N_1322,In_1349,In_2374);
and U1323 (N_1323,In_2457,In_58);
nand U1324 (N_1324,In_2294,In_1888);
and U1325 (N_1325,In_1154,In_1016);
and U1326 (N_1326,In_1744,In_717);
or U1327 (N_1327,In_706,In_357);
and U1328 (N_1328,In_741,In_1555);
and U1329 (N_1329,In_688,In_1376);
and U1330 (N_1330,In_1881,In_92);
or U1331 (N_1331,In_885,In_1290);
or U1332 (N_1332,In_862,In_742);
nor U1333 (N_1333,In_693,In_2460);
nand U1334 (N_1334,In_320,In_652);
xor U1335 (N_1335,In_770,In_390);
nor U1336 (N_1336,In_1497,In_1855);
and U1337 (N_1337,In_1838,In_573);
nand U1338 (N_1338,In_1638,In_278);
xnor U1339 (N_1339,In_2023,In_695);
and U1340 (N_1340,In_1338,In_92);
or U1341 (N_1341,In_2462,In_2405);
xnor U1342 (N_1342,In_1174,In_580);
nor U1343 (N_1343,In_38,In_2147);
xnor U1344 (N_1344,In_723,In_686);
and U1345 (N_1345,In_410,In_88);
nor U1346 (N_1346,In_1447,In_1971);
nand U1347 (N_1347,In_1957,In_481);
and U1348 (N_1348,In_1133,In_456);
nand U1349 (N_1349,In_1299,In_1775);
nand U1350 (N_1350,In_361,In_1445);
xnor U1351 (N_1351,In_1941,In_256);
nor U1352 (N_1352,In_671,In_1698);
nor U1353 (N_1353,In_397,In_1362);
and U1354 (N_1354,In_2245,In_1801);
and U1355 (N_1355,In_1366,In_2075);
or U1356 (N_1356,In_577,In_1010);
and U1357 (N_1357,In_1975,In_1061);
xor U1358 (N_1358,In_2162,In_1529);
nor U1359 (N_1359,In_1594,In_1561);
or U1360 (N_1360,In_1718,In_1469);
and U1361 (N_1361,In_1073,In_2079);
xor U1362 (N_1362,In_1547,In_2073);
and U1363 (N_1363,In_2232,In_256);
xnor U1364 (N_1364,In_139,In_269);
nor U1365 (N_1365,In_37,In_1206);
and U1366 (N_1366,In_2326,In_1236);
nor U1367 (N_1367,In_1175,In_1573);
xor U1368 (N_1368,In_487,In_1726);
and U1369 (N_1369,In_2406,In_1757);
nor U1370 (N_1370,In_458,In_2224);
xor U1371 (N_1371,In_206,In_202);
xnor U1372 (N_1372,In_1075,In_254);
and U1373 (N_1373,In_2442,In_592);
nand U1374 (N_1374,In_1618,In_1769);
nand U1375 (N_1375,In_1040,In_52);
and U1376 (N_1376,In_1812,In_930);
nand U1377 (N_1377,In_2478,In_602);
nand U1378 (N_1378,In_1720,In_137);
nor U1379 (N_1379,In_2142,In_2088);
xor U1380 (N_1380,In_650,In_1302);
or U1381 (N_1381,In_1375,In_1243);
and U1382 (N_1382,In_1684,In_1468);
nand U1383 (N_1383,In_2117,In_469);
and U1384 (N_1384,In_2147,In_1926);
and U1385 (N_1385,In_1816,In_307);
or U1386 (N_1386,In_676,In_1940);
or U1387 (N_1387,In_2338,In_1540);
or U1388 (N_1388,In_1971,In_1856);
xnor U1389 (N_1389,In_959,In_1852);
nor U1390 (N_1390,In_1044,In_2258);
and U1391 (N_1391,In_1968,In_149);
nand U1392 (N_1392,In_1404,In_1356);
nand U1393 (N_1393,In_1357,In_1665);
nand U1394 (N_1394,In_2493,In_471);
and U1395 (N_1395,In_1183,In_141);
nor U1396 (N_1396,In_894,In_1967);
and U1397 (N_1397,In_484,In_1925);
and U1398 (N_1398,In_1121,In_578);
and U1399 (N_1399,In_2373,In_1665);
nor U1400 (N_1400,In_44,In_1465);
nand U1401 (N_1401,In_1534,In_1361);
or U1402 (N_1402,In_332,In_456);
and U1403 (N_1403,In_994,In_1118);
and U1404 (N_1404,In_2490,In_1829);
nor U1405 (N_1405,In_957,In_1651);
xnor U1406 (N_1406,In_2208,In_855);
nor U1407 (N_1407,In_1059,In_1090);
nand U1408 (N_1408,In_1349,In_2464);
xnor U1409 (N_1409,In_260,In_2361);
and U1410 (N_1410,In_677,In_1523);
nand U1411 (N_1411,In_76,In_2323);
nor U1412 (N_1412,In_1345,In_999);
nor U1413 (N_1413,In_1582,In_741);
nor U1414 (N_1414,In_996,In_437);
and U1415 (N_1415,In_2392,In_2065);
nor U1416 (N_1416,In_2090,In_1186);
nor U1417 (N_1417,In_1024,In_456);
nand U1418 (N_1418,In_2262,In_1892);
xor U1419 (N_1419,In_266,In_1903);
and U1420 (N_1420,In_590,In_2294);
nor U1421 (N_1421,In_1749,In_1139);
or U1422 (N_1422,In_1589,In_520);
or U1423 (N_1423,In_879,In_465);
and U1424 (N_1424,In_798,In_1474);
xor U1425 (N_1425,In_1381,In_1524);
nand U1426 (N_1426,In_2125,In_1223);
xnor U1427 (N_1427,In_2347,In_1891);
and U1428 (N_1428,In_2008,In_1649);
nand U1429 (N_1429,In_168,In_562);
and U1430 (N_1430,In_765,In_1433);
or U1431 (N_1431,In_1741,In_2083);
and U1432 (N_1432,In_1239,In_459);
nand U1433 (N_1433,In_2016,In_1784);
and U1434 (N_1434,In_508,In_621);
xor U1435 (N_1435,In_908,In_1926);
nor U1436 (N_1436,In_1635,In_1802);
and U1437 (N_1437,In_2467,In_1867);
nor U1438 (N_1438,In_2118,In_1128);
or U1439 (N_1439,In_1125,In_33);
nand U1440 (N_1440,In_870,In_908);
nor U1441 (N_1441,In_1096,In_1206);
xor U1442 (N_1442,In_776,In_1535);
or U1443 (N_1443,In_1031,In_2160);
xor U1444 (N_1444,In_2250,In_136);
and U1445 (N_1445,In_972,In_724);
or U1446 (N_1446,In_950,In_1493);
nand U1447 (N_1447,In_2088,In_1342);
and U1448 (N_1448,In_1968,In_1555);
nand U1449 (N_1449,In_2478,In_232);
nand U1450 (N_1450,In_883,In_1461);
and U1451 (N_1451,In_2345,In_1314);
or U1452 (N_1452,In_1854,In_488);
xor U1453 (N_1453,In_1588,In_969);
xnor U1454 (N_1454,In_1196,In_133);
or U1455 (N_1455,In_174,In_1844);
and U1456 (N_1456,In_2082,In_2032);
and U1457 (N_1457,In_1302,In_424);
xnor U1458 (N_1458,In_793,In_2109);
xnor U1459 (N_1459,In_1343,In_2230);
or U1460 (N_1460,In_1677,In_1081);
nand U1461 (N_1461,In_1943,In_291);
xnor U1462 (N_1462,In_268,In_1436);
and U1463 (N_1463,In_381,In_244);
or U1464 (N_1464,In_1968,In_1104);
nor U1465 (N_1465,In_296,In_821);
and U1466 (N_1466,In_2423,In_1119);
nand U1467 (N_1467,In_1871,In_1233);
xor U1468 (N_1468,In_341,In_999);
nor U1469 (N_1469,In_1846,In_484);
xnor U1470 (N_1470,In_1791,In_379);
or U1471 (N_1471,In_1570,In_1851);
or U1472 (N_1472,In_2068,In_1881);
nor U1473 (N_1473,In_2466,In_2316);
and U1474 (N_1474,In_672,In_459);
and U1475 (N_1475,In_2032,In_1977);
or U1476 (N_1476,In_1137,In_830);
nor U1477 (N_1477,In_2361,In_1929);
or U1478 (N_1478,In_760,In_2391);
or U1479 (N_1479,In_1476,In_1281);
or U1480 (N_1480,In_1548,In_1077);
nand U1481 (N_1481,In_1523,In_1128);
or U1482 (N_1482,In_1317,In_1210);
or U1483 (N_1483,In_1622,In_1330);
and U1484 (N_1484,In_2048,In_583);
xor U1485 (N_1485,In_1821,In_2384);
or U1486 (N_1486,In_470,In_467);
xor U1487 (N_1487,In_636,In_2030);
or U1488 (N_1488,In_2492,In_400);
and U1489 (N_1489,In_2454,In_1501);
and U1490 (N_1490,In_67,In_1665);
xor U1491 (N_1491,In_1734,In_1408);
nand U1492 (N_1492,In_1578,In_26);
nor U1493 (N_1493,In_2493,In_2451);
nand U1494 (N_1494,In_814,In_1872);
and U1495 (N_1495,In_1678,In_1751);
or U1496 (N_1496,In_2489,In_1842);
or U1497 (N_1497,In_934,In_82);
nand U1498 (N_1498,In_1470,In_911);
nor U1499 (N_1499,In_172,In_445);
and U1500 (N_1500,In_2039,In_1530);
nand U1501 (N_1501,In_1576,In_205);
xnor U1502 (N_1502,In_1362,In_2060);
nor U1503 (N_1503,In_269,In_2258);
and U1504 (N_1504,In_864,In_1963);
or U1505 (N_1505,In_1110,In_2149);
nor U1506 (N_1506,In_1234,In_304);
or U1507 (N_1507,In_1847,In_2412);
xnor U1508 (N_1508,In_2230,In_445);
nand U1509 (N_1509,In_730,In_2131);
or U1510 (N_1510,In_2397,In_2487);
nor U1511 (N_1511,In_988,In_1149);
and U1512 (N_1512,In_490,In_430);
xnor U1513 (N_1513,In_1952,In_2213);
or U1514 (N_1514,In_290,In_535);
or U1515 (N_1515,In_442,In_876);
nor U1516 (N_1516,In_616,In_2109);
nor U1517 (N_1517,In_87,In_785);
nor U1518 (N_1518,In_990,In_767);
xnor U1519 (N_1519,In_286,In_1804);
or U1520 (N_1520,In_2290,In_797);
and U1521 (N_1521,In_2059,In_1338);
nor U1522 (N_1522,In_948,In_821);
xor U1523 (N_1523,In_606,In_1135);
xnor U1524 (N_1524,In_2410,In_1290);
xnor U1525 (N_1525,In_139,In_2092);
and U1526 (N_1526,In_2323,In_2271);
xor U1527 (N_1527,In_1901,In_1249);
nand U1528 (N_1528,In_1845,In_804);
or U1529 (N_1529,In_2173,In_1333);
and U1530 (N_1530,In_477,In_1041);
nand U1531 (N_1531,In_2229,In_718);
or U1532 (N_1532,In_1654,In_1868);
and U1533 (N_1533,In_1487,In_2328);
nand U1534 (N_1534,In_1139,In_2487);
or U1535 (N_1535,In_992,In_851);
and U1536 (N_1536,In_927,In_1632);
nor U1537 (N_1537,In_748,In_2177);
nor U1538 (N_1538,In_2412,In_535);
xor U1539 (N_1539,In_1172,In_942);
nor U1540 (N_1540,In_1432,In_769);
and U1541 (N_1541,In_1874,In_1273);
or U1542 (N_1542,In_1507,In_406);
and U1543 (N_1543,In_736,In_470);
nand U1544 (N_1544,In_660,In_206);
xor U1545 (N_1545,In_953,In_1330);
or U1546 (N_1546,In_663,In_1891);
and U1547 (N_1547,In_1870,In_1397);
nand U1548 (N_1548,In_178,In_15);
xnor U1549 (N_1549,In_1623,In_1713);
and U1550 (N_1550,In_472,In_1449);
and U1551 (N_1551,In_1131,In_168);
nor U1552 (N_1552,In_1618,In_2427);
and U1553 (N_1553,In_1721,In_1226);
xor U1554 (N_1554,In_1143,In_794);
or U1555 (N_1555,In_2006,In_1428);
xor U1556 (N_1556,In_1917,In_1271);
xnor U1557 (N_1557,In_1297,In_2124);
xnor U1558 (N_1558,In_1976,In_2337);
or U1559 (N_1559,In_1194,In_2085);
or U1560 (N_1560,In_172,In_1091);
nand U1561 (N_1561,In_1845,In_1357);
nand U1562 (N_1562,In_1778,In_727);
xor U1563 (N_1563,In_430,In_1342);
nor U1564 (N_1564,In_271,In_2412);
and U1565 (N_1565,In_1963,In_1707);
or U1566 (N_1566,In_878,In_661);
nand U1567 (N_1567,In_191,In_708);
or U1568 (N_1568,In_479,In_515);
or U1569 (N_1569,In_9,In_152);
or U1570 (N_1570,In_1809,In_1712);
xnor U1571 (N_1571,In_2306,In_1394);
and U1572 (N_1572,In_532,In_298);
xor U1573 (N_1573,In_634,In_309);
nand U1574 (N_1574,In_2254,In_1803);
or U1575 (N_1575,In_107,In_1893);
xnor U1576 (N_1576,In_1189,In_1607);
xnor U1577 (N_1577,In_2333,In_2117);
nand U1578 (N_1578,In_559,In_2168);
and U1579 (N_1579,In_244,In_610);
or U1580 (N_1580,In_2130,In_2228);
and U1581 (N_1581,In_143,In_517);
xnor U1582 (N_1582,In_1320,In_1226);
xor U1583 (N_1583,In_1030,In_1790);
xor U1584 (N_1584,In_774,In_1799);
or U1585 (N_1585,In_1010,In_1146);
and U1586 (N_1586,In_1090,In_1705);
and U1587 (N_1587,In_479,In_796);
nor U1588 (N_1588,In_2247,In_1272);
and U1589 (N_1589,In_2481,In_2418);
or U1590 (N_1590,In_1361,In_519);
and U1591 (N_1591,In_1087,In_687);
or U1592 (N_1592,In_743,In_1491);
nor U1593 (N_1593,In_278,In_2335);
or U1594 (N_1594,In_727,In_2369);
or U1595 (N_1595,In_718,In_2318);
or U1596 (N_1596,In_968,In_245);
xor U1597 (N_1597,In_461,In_2484);
nor U1598 (N_1598,In_1026,In_1674);
and U1599 (N_1599,In_107,In_424);
nor U1600 (N_1600,In_1920,In_2446);
or U1601 (N_1601,In_1871,In_334);
xor U1602 (N_1602,In_762,In_246);
or U1603 (N_1603,In_1685,In_853);
nand U1604 (N_1604,In_1654,In_1556);
nand U1605 (N_1605,In_1857,In_954);
nand U1606 (N_1606,In_1700,In_2114);
xnor U1607 (N_1607,In_1510,In_111);
nor U1608 (N_1608,In_417,In_2074);
nor U1609 (N_1609,In_2456,In_2126);
nand U1610 (N_1610,In_1662,In_462);
xor U1611 (N_1611,In_762,In_1884);
and U1612 (N_1612,In_363,In_2446);
xnor U1613 (N_1613,In_1802,In_2238);
nand U1614 (N_1614,In_408,In_1169);
and U1615 (N_1615,In_264,In_1094);
xnor U1616 (N_1616,In_3,In_2201);
nor U1617 (N_1617,In_629,In_883);
or U1618 (N_1618,In_2041,In_527);
nor U1619 (N_1619,In_593,In_1358);
xnor U1620 (N_1620,In_1117,In_852);
nor U1621 (N_1621,In_897,In_583);
nand U1622 (N_1622,In_1506,In_826);
or U1623 (N_1623,In_2379,In_351);
xor U1624 (N_1624,In_2038,In_337);
and U1625 (N_1625,In_1575,In_2086);
nand U1626 (N_1626,In_1971,In_2029);
nor U1627 (N_1627,In_488,In_2263);
nand U1628 (N_1628,In_64,In_920);
xnor U1629 (N_1629,In_572,In_2263);
nor U1630 (N_1630,In_2439,In_49);
nand U1631 (N_1631,In_799,In_1919);
xnor U1632 (N_1632,In_17,In_1869);
and U1633 (N_1633,In_1862,In_1588);
and U1634 (N_1634,In_2408,In_1812);
or U1635 (N_1635,In_2390,In_1427);
nand U1636 (N_1636,In_2362,In_571);
xor U1637 (N_1637,In_95,In_2230);
or U1638 (N_1638,In_2272,In_611);
or U1639 (N_1639,In_1242,In_2169);
xor U1640 (N_1640,In_774,In_2);
nor U1641 (N_1641,In_871,In_490);
nor U1642 (N_1642,In_2478,In_1900);
xor U1643 (N_1643,In_2358,In_2064);
xnor U1644 (N_1644,In_702,In_522);
nor U1645 (N_1645,In_1172,In_1275);
nor U1646 (N_1646,In_532,In_673);
or U1647 (N_1647,In_554,In_1237);
xor U1648 (N_1648,In_305,In_2441);
or U1649 (N_1649,In_803,In_318);
nor U1650 (N_1650,In_1424,In_775);
nand U1651 (N_1651,In_2136,In_2274);
or U1652 (N_1652,In_595,In_236);
xnor U1653 (N_1653,In_1218,In_2016);
nand U1654 (N_1654,In_1377,In_1506);
or U1655 (N_1655,In_879,In_2321);
or U1656 (N_1656,In_1753,In_302);
nand U1657 (N_1657,In_1129,In_962);
nor U1658 (N_1658,In_247,In_972);
nand U1659 (N_1659,In_1946,In_2247);
or U1660 (N_1660,In_338,In_1870);
nor U1661 (N_1661,In_2151,In_1492);
nand U1662 (N_1662,In_602,In_2293);
xnor U1663 (N_1663,In_2491,In_1330);
nand U1664 (N_1664,In_212,In_350);
nand U1665 (N_1665,In_155,In_1606);
or U1666 (N_1666,In_1497,In_2301);
nand U1667 (N_1667,In_575,In_837);
and U1668 (N_1668,In_2142,In_1703);
xnor U1669 (N_1669,In_726,In_2157);
xnor U1670 (N_1670,In_579,In_833);
xnor U1671 (N_1671,In_994,In_481);
or U1672 (N_1672,In_1725,In_1733);
nor U1673 (N_1673,In_910,In_77);
or U1674 (N_1674,In_1420,In_1146);
or U1675 (N_1675,In_410,In_1089);
nand U1676 (N_1676,In_124,In_259);
nor U1677 (N_1677,In_1014,In_834);
nor U1678 (N_1678,In_1779,In_1855);
nand U1679 (N_1679,In_1675,In_2320);
or U1680 (N_1680,In_552,In_2219);
nor U1681 (N_1681,In_666,In_49);
nand U1682 (N_1682,In_998,In_2472);
nor U1683 (N_1683,In_826,In_2276);
and U1684 (N_1684,In_1573,In_1799);
and U1685 (N_1685,In_667,In_1631);
nor U1686 (N_1686,In_1168,In_1464);
or U1687 (N_1687,In_36,In_2293);
nor U1688 (N_1688,In_1978,In_2425);
and U1689 (N_1689,In_2224,In_1892);
or U1690 (N_1690,In_342,In_1584);
or U1691 (N_1691,In_1406,In_906);
nor U1692 (N_1692,In_353,In_1236);
and U1693 (N_1693,In_1822,In_1600);
nand U1694 (N_1694,In_1607,In_1706);
nand U1695 (N_1695,In_133,In_1360);
nand U1696 (N_1696,In_1349,In_1325);
nand U1697 (N_1697,In_1125,In_719);
nand U1698 (N_1698,In_441,In_609);
and U1699 (N_1699,In_1894,In_937);
nor U1700 (N_1700,In_2022,In_1296);
nand U1701 (N_1701,In_1602,In_2477);
xnor U1702 (N_1702,In_908,In_1172);
nor U1703 (N_1703,In_891,In_713);
xnor U1704 (N_1704,In_1233,In_282);
and U1705 (N_1705,In_967,In_347);
nand U1706 (N_1706,In_1435,In_1411);
nor U1707 (N_1707,In_1672,In_854);
or U1708 (N_1708,In_506,In_1922);
or U1709 (N_1709,In_1638,In_2024);
xnor U1710 (N_1710,In_2481,In_735);
and U1711 (N_1711,In_1506,In_1022);
and U1712 (N_1712,In_596,In_2086);
xnor U1713 (N_1713,In_1758,In_2273);
nand U1714 (N_1714,In_1839,In_1511);
nand U1715 (N_1715,In_1103,In_556);
and U1716 (N_1716,In_122,In_1094);
xor U1717 (N_1717,In_234,In_1298);
xnor U1718 (N_1718,In_2477,In_2307);
xnor U1719 (N_1719,In_1070,In_60);
nand U1720 (N_1720,In_2218,In_578);
nand U1721 (N_1721,In_295,In_550);
nor U1722 (N_1722,In_756,In_899);
nand U1723 (N_1723,In_1322,In_132);
xor U1724 (N_1724,In_2426,In_1932);
or U1725 (N_1725,In_1554,In_753);
and U1726 (N_1726,In_7,In_904);
xnor U1727 (N_1727,In_963,In_1401);
and U1728 (N_1728,In_2112,In_2476);
xnor U1729 (N_1729,In_2227,In_1035);
and U1730 (N_1730,In_1113,In_2003);
xor U1731 (N_1731,In_962,In_1118);
and U1732 (N_1732,In_600,In_1233);
nand U1733 (N_1733,In_998,In_2346);
xnor U1734 (N_1734,In_1185,In_2175);
and U1735 (N_1735,In_2145,In_2024);
nor U1736 (N_1736,In_1191,In_539);
nor U1737 (N_1737,In_355,In_148);
nand U1738 (N_1738,In_2158,In_2188);
nor U1739 (N_1739,In_1005,In_201);
nor U1740 (N_1740,In_2418,In_161);
nand U1741 (N_1741,In_1333,In_140);
nor U1742 (N_1742,In_812,In_1454);
and U1743 (N_1743,In_526,In_2325);
nor U1744 (N_1744,In_2043,In_2454);
or U1745 (N_1745,In_219,In_1321);
and U1746 (N_1746,In_217,In_865);
or U1747 (N_1747,In_1572,In_65);
xor U1748 (N_1748,In_1756,In_548);
and U1749 (N_1749,In_2221,In_2279);
xnor U1750 (N_1750,In_1454,In_1844);
and U1751 (N_1751,In_1330,In_1126);
nor U1752 (N_1752,In_50,In_1507);
nand U1753 (N_1753,In_558,In_1379);
nand U1754 (N_1754,In_29,In_245);
or U1755 (N_1755,In_2081,In_2414);
nand U1756 (N_1756,In_1604,In_1317);
or U1757 (N_1757,In_1005,In_152);
nand U1758 (N_1758,In_600,In_1503);
nor U1759 (N_1759,In_2374,In_2177);
nor U1760 (N_1760,In_157,In_1534);
nand U1761 (N_1761,In_1699,In_1404);
xor U1762 (N_1762,In_95,In_280);
and U1763 (N_1763,In_1955,In_2130);
nand U1764 (N_1764,In_1074,In_1858);
nand U1765 (N_1765,In_454,In_699);
or U1766 (N_1766,In_1414,In_1926);
nor U1767 (N_1767,In_1879,In_169);
or U1768 (N_1768,In_393,In_2100);
xor U1769 (N_1769,In_2164,In_553);
nor U1770 (N_1770,In_34,In_2192);
xor U1771 (N_1771,In_1460,In_303);
and U1772 (N_1772,In_277,In_122);
nand U1773 (N_1773,In_388,In_543);
xnor U1774 (N_1774,In_851,In_243);
or U1775 (N_1775,In_1541,In_574);
xnor U1776 (N_1776,In_1863,In_2134);
xor U1777 (N_1777,In_286,In_924);
and U1778 (N_1778,In_1477,In_2397);
nor U1779 (N_1779,In_437,In_2324);
nand U1780 (N_1780,In_1317,In_161);
and U1781 (N_1781,In_1106,In_263);
nand U1782 (N_1782,In_1003,In_1521);
nand U1783 (N_1783,In_1890,In_1523);
nand U1784 (N_1784,In_764,In_188);
nand U1785 (N_1785,In_1234,In_666);
nand U1786 (N_1786,In_1175,In_2437);
xor U1787 (N_1787,In_2159,In_239);
nor U1788 (N_1788,In_2412,In_1998);
nand U1789 (N_1789,In_533,In_786);
nand U1790 (N_1790,In_900,In_188);
nand U1791 (N_1791,In_490,In_1407);
xnor U1792 (N_1792,In_293,In_1795);
or U1793 (N_1793,In_2339,In_1870);
xor U1794 (N_1794,In_75,In_1602);
or U1795 (N_1795,In_2436,In_1866);
and U1796 (N_1796,In_290,In_1628);
nand U1797 (N_1797,In_345,In_1977);
nor U1798 (N_1798,In_1814,In_867);
or U1799 (N_1799,In_80,In_1851);
nor U1800 (N_1800,In_1483,In_451);
and U1801 (N_1801,In_1120,In_34);
or U1802 (N_1802,In_90,In_2);
xnor U1803 (N_1803,In_949,In_669);
and U1804 (N_1804,In_1338,In_1048);
or U1805 (N_1805,In_45,In_1809);
nand U1806 (N_1806,In_2135,In_474);
xnor U1807 (N_1807,In_1695,In_1608);
nand U1808 (N_1808,In_2137,In_1255);
nor U1809 (N_1809,In_1567,In_1654);
and U1810 (N_1810,In_1170,In_419);
and U1811 (N_1811,In_1296,In_1064);
nor U1812 (N_1812,In_1205,In_494);
nor U1813 (N_1813,In_1194,In_667);
and U1814 (N_1814,In_1806,In_1931);
nand U1815 (N_1815,In_2178,In_1413);
xor U1816 (N_1816,In_535,In_32);
and U1817 (N_1817,In_1187,In_747);
or U1818 (N_1818,In_1031,In_285);
and U1819 (N_1819,In_1932,In_863);
nand U1820 (N_1820,In_398,In_588);
and U1821 (N_1821,In_47,In_1741);
xor U1822 (N_1822,In_2481,In_1692);
nand U1823 (N_1823,In_1872,In_907);
nand U1824 (N_1824,In_1579,In_1654);
nand U1825 (N_1825,In_917,In_1835);
nor U1826 (N_1826,In_1885,In_82);
nor U1827 (N_1827,In_1751,In_393);
or U1828 (N_1828,In_1080,In_2428);
xnor U1829 (N_1829,In_1994,In_892);
and U1830 (N_1830,In_1716,In_1503);
and U1831 (N_1831,In_367,In_747);
and U1832 (N_1832,In_1240,In_669);
nand U1833 (N_1833,In_2333,In_444);
xnor U1834 (N_1834,In_270,In_954);
and U1835 (N_1835,In_1534,In_2099);
or U1836 (N_1836,In_1617,In_915);
nor U1837 (N_1837,In_1840,In_1197);
xor U1838 (N_1838,In_1901,In_238);
or U1839 (N_1839,In_1994,In_1275);
nand U1840 (N_1840,In_153,In_2231);
and U1841 (N_1841,In_653,In_1023);
or U1842 (N_1842,In_2163,In_746);
nor U1843 (N_1843,In_2054,In_2455);
or U1844 (N_1844,In_2326,In_984);
and U1845 (N_1845,In_579,In_1742);
and U1846 (N_1846,In_843,In_561);
nand U1847 (N_1847,In_288,In_582);
nor U1848 (N_1848,In_284,In_1794);
xor U1849 (N_1849,In_867,In_2150);
nor U1850 (N_1850,In_938,In_1704);
nor U1851 (N_1851,In_79,In_375);
or U1852 (N_1852,In_695,In_1185);
nand U1853 (N_1853,In_893,In_2051);
nand U1854 (N_1854,In_704,In_254);
nor U1855 (N_1855,In_2378,In_303);
or U1856 (N_1856,In_732,In_2220);
or U1857 (N_1857,In_535,In_1147);
or U1858 (N_1858,In_213,In_461);
or U1859 (N_1859,In_2250,In_678);
and U1860 (N_1860,In_1466,In_281);
and U1861 (N_1861,In_2350,In_1519);
or U1862 (N_1862,In_1969,In_2333);
nor U1863 (N_1863,In_439,In_81);
nor U1864 (N_1864,In_2178,In_2211);
nand U1865 (N_1865,In_350,In_1458);
and U1866 (N_1866,In_393,In_11);
nor U1867 (N_1867,In_1934,In_1506);
nand U1868 (N_1868,In_1354,In_1421);
xor U1869 (N_1869,In_1401,In_2161);
and U1870 (N_1870,In_1212,In_138);
or U1871 (N_1871,In_2226,In_37);
and U1872 (N_1872,In_764,In_1241);
xnor U1873 (N_1873,In_1698,In_2068);
xnor U1874 (N_1874,In_2006,In_516);
xor U1875 (N_1875,In_1692,In_2073);
or U1876 (N_1876,In_1724,In_1986);
or U1877 (N_1877,In_1049,In_1570);
and U1878 (N_1878,In_530,In_1736);
and U1879 (N_1879,In_911,In_1296);
xor U1880 (N_1880,In_2279,In_1499);
nor U1881 (N_1881,In_2303,In_2152);
or U1882 (N_1882,In_2377,In_1236);
and U1883 (N_1883,In_2237,In_746);
or U1884 (N_1884,In_2259,In_1524);
xnor U1885 (N_1885,In_1328,In_1801);
nor U1886 (N_1886,In_125,In_1198);
or U1887 (N_1887,In_805,In_917);
or U1888 (N_1888,In_2216,In_2234);
nor U1889 (N_1889,In_1019,In_1259);
nand U1890 (N_1890,In_1162,In_386);
nor U1891 (N_1891,In_2027,In_495);
and U1892 (N_1892,In_1791,In_1111);
nand U1893 (N_1893,In_1721,In_603);
xnor U1894 (N_1894,In_311,In_2118);
nor U1895 (N_1895,In_345,In_414);
xor U1896 (N_1896,In_898,In_1033);
or U1897 (N_1897,In_808,In_802);
or U1898 (N_1898,In_535,In_2416);
or U1899 (N_1899,In_1759,In_1030);
xor U1900 (N_1900,In_2233,In_2201);
and U1901 (N_1901,In_2375,In_2081);
nand U1902 (N_1902,In_1912,In_1819);
xor U1903 (N_1903,In_1112,In_622);
and U1904 (N_1904,In_1450,In_1103);
nor U1905 (N_1905,In_2041,In_1385);
nor U1906 (N_1906,In_232,In_1750);
nand U1907 (N_1907,In_325,In_2021);
and U1908 (N_1908,In_521,In_1089);
xnor U1909 (N_1909,In_1541,In_1059);
nand U1910 (N_1910,In_1563,In_2031);
nand U1911 (N_1911,In_826,In_1004);
xor U1912 (N_1912,In_1082,In_938);
nand U1913 (N_1913,In_208,In_1381);
or U1914 (N_1914,In_109,In_165);
nand U1915 (N_1915,In_950,In_248);
or U1916 (N_1916,In_1000,In_231);
nand U1917 (N_1917,In_288,In_1073);
nor U1918 (N_1918,In_1581,In_42);
nand U1919 (N_1919,In_2113,In_32);
nor U1920 (N_1920,In_562,In_1095);
and U1921 (N_1921,In_924,In_1260);
nand U1922 (N_1922,In_489,In_1214);
nand U1923 (N_1923,In_222,In_37);
or U1924 (N_1924,In_439,In_1210);
or U1925 (N_1925,In_1603,In_1397);
nand U1926 (N_1926,In_133,In_2136);
or U1927 (N_1927,In_2254,In_499);
xnor U1928 (N_1928,In_2056,In_367);
xnor U1929 (N_1929,In_1512,In_2096);
nor U1930 (N_1930,In_1844,In_2386);
or U1931 (N_1931,In_1572,In_1001);
or U1932 (N_1932,In_407,In_1641);
nor U1933 (N_1933,In_2016,In_1075);
xnor U1934 (N_1934,In_669,In_1326);
or U1935 (N_1935,In_2076,In_673);
nand U1936 (N_1936,In_834,In_593);
nand U1937 (N_1937,In_140,In_15);
xor U1938 (N_1938,In_1175,In_230);
or U1939 (N_1939,In_2412,In_331);
and U1940 (N_1940,In_2430,In_888);
and U1941 (N_1941,In_630,In_1546);
nand U1942 (N_1942,In_722,In_889);
nor U1943 (N_1943,In_1707,In_2118);
nor U1944 (N_1944,In_1754,In_438);
nor U1945 (N_1945,In_2325,In_511);
and U1946 (N_1946,In_1062,In_988);
nand U1947 (N_1947,In_2276,In_59);
xor U1948 (N_1948,In_1162,In_1031);
and U1949 (N_1949,In_817,In_1651);
xor U1950 (N_1950,In_1316,In_2432);
and U1951 (N_1951,In_2235,In_1537);
nand U1952 (N_1952,In_174,In_275);
and U1953 (N_1953,In_2211,In_1744);
or U1954 (N_1954,In_2314,In_729);
nor U1955 (N_1955,In_1978,In_1679);
nor U1956 (N_1956,In_1069,In_719);
nand U1957 (N_1957,In_2166,In_716);
and U1958 (N_1958,In_1748,In_1593);
xnor U1959 (N_1959,In_2158,In_493);
or U1960 (N_1960,In_682,In_2490);
and U1961 (N_1961,In_1438,In_2053);
xor U1962 (N_1962,In_2435,In_316);
nand U1963 (N_1963,In_2016,In_2180);
nor U1964 (N_1964,In_182,In_1176);
nor U1965 (N_1965,In_1,In_1967);
nand U1966 (N_1966,In_227,In_594);
or U1967 (N_1967,In_12,In_853);
or U1968 (N_1968,In_1890,In_1642);
xnor U1969 (N_1969,In_684,In_611);
and U1970 (N_1970,In_442,In_1942);
and U1971 (N_1971,In_691,In_326);
nor U1972 (N_1972,In_1090,In_1154);
or U1973 (N_1973,In_77,In_1614);
and U1974 (N_1974,In_2463,In_970);
xnor U1975 (N_1975,In_1215,In_199);
nor U1976 (N_1976,In_1383,In_74);
nor U1977 (N_1977,In_1494,In_1353);
and U1978 (N_1978,In_905,In_1035);
nor U1979 (N_1979,In_1087,In_793);
nor U1980 (N_1980,In_1735,In_1996);
and U1981 (N_1981,In_1336,In_239);
nor U1982 (N_1982,In_669,In_153);
xor U1983 (N_1983,In_1488,In_848);
or U1984 (N_1984,In_1429,In_84);
or U1985 (N_1985,In_796,In_537);
or U1986 (N_1986,In_457,In_1317);
nand U1987 (N_1987,In_1834,In_659);
nor U1988 (N_1988,In_1360,In_2318);
and U1989 (N_1989,In_1982,In_1701);
xnor U1990 (N_1990,In_1601,In_1379);
nor U1991 (N_1991,In_603,In_154);
and U1992 (N_1992,In_1848,In_2044);
and U1993 (N_1993,In_1919,In_1391);
nand U1994 (N_1994,In_1061,In_493);
or U1995 (N_1995,In_846,In_1763);
nor U1996 (N_1996,In_885,In_1363);
or U1997 (N_1997,In_591,In_2029);
and U1998 (N_1998,In_2346,In_9);
and U1999 (N_1999,In_2213,In_613);
and U2000 (N_2000,In_755,In_1093);
xor U2001 (N_2001,In_1759,In_239);
nor U2002 (N_2002,In_205,In_2047);
xnor U2003 (N_2003,In_445,In_1926);
or U2004 (N_2004,In_2461,In_1296);
nand U2005 (N_2005,In_226,In_701);
nor U2006 (N_2006,In_141,In_2472);
xnor U2007 (N_2007,In_2145,In_1977);
nand U2008 (N_2008,In_235,In_1564);
nand U2009 (N_2009,In_342,In_56);
and U2010 (N_2010,In_611,In_1028);
and U2011 (N_2011,In_238,In_659);
and U2012 (N_2012,In_67,In_1249);
xnor U2013 (N_2013,In_2252,In_1179);
xor U2014 (N_2014,In_21,In_2018);
nor U2015 (N_2015,In_2104,In_1682);
nor U2016 (N_2016,In_361,In_734);
and U2017 (N_2017,In_800,In_1723);
nand U2018 (N_2018,In_2491,In_408);
or U2019 (N_2019,In_120,In_268);
xor U2020 (N_2020,In_766,In_1032);
xnor U2021 (N_2021,In_482,In_1728);
nor U2022 (N_2022,In_316,In_1476);
nor U2023 (N_2023,In_1736,In_1855);
or U2024 (N_2024,In_1735,In_1409);
nand U2025 (N_2025,In_2284,In_428);
or U2026 (N_2026,In_215,In_1312);
and U2027 (N_2027,In_922,In_878);
nand U2028 (N_2028,In_1690,In_172);
xor U2029 (N_2029,In_2116,In_617);
nor U2030 (N_2030,In_391,In_2392);
nor U2031 (N_2031,In_446,In_2045);
and U2032 (N_2032,In_1393,In_1938);
or U2033 (N_2033,In_1860,In_727);
and U2034 (N_2034,In_196,In_68);
or U2035 (N_2035,In_480,In_2416);
nand U2036 (N_2036,In_2489,In_1343);
or U2037 (N_2037,In_754,In_1000);
xor U2038 (N_2038,In_1631,In_1848);
nor U2039 (N_2039,In_2226,In_1257);
nor U2040 (N_2040,In_2468,In_2353);
nand U2041 (N_2041,In_740,In_361);
nand U2042 (N_2042,In_1541,In_347);
nor U2043 (N_2043,In_729,In_13);
nand U2044 (N_2044,In_345,In_740);
xnor U2045 (N_2045,In_1076,In_48);
nand U2046 (N_2046,In_1926,In_1507);
nand U2047 (N_2047,In_1045,In_12);
nor U2048 (N_2048,In_985,In_1671);
and U2049 (N_2049,In_95,In_1926);
or U2050 (N_2050,In_2472,In_255);
nor U2051 (N_2051,In_633,In_1817);
nand U2052 (N_2052,In_821,In_1146);
nand U2053 (N_2053,In_133,In_507);
and U2054 (N_2054,In_1326,In_2216);
xnor U2055 (N_2055,In_2468,In_1136);
xor U2056 (N_2056,In_427,In_1935);
nand U2057 (N_2057,In_1234,In_1338);
or U2058 (N_2058,In_261,In_1835);
nand U2059 (N_2059,In_245,In_2123);
nand U2060 (N_2060,In_1698,In_2455);
nor U2061 (N_2061,In_944,In_462);
xnor U2062 (N_2062,In_1709,In_467);
xor U2063 (N_2063,In_2358,In_2377);
and U2064 (N_2064,In_1682,In_735);
and U2065 (N_2065,In_2281,In_446);
or U2066 (N_2066,In_1654,In_1264);
nor U2067 (N_2067,In_243,In_901);
nand U2068 (N_2068,In_1187,In_2269);
and U2069 (N_2069,In_297,In_1750);
xor U2070 (N_2070,In_2361,In_1664);
xnor U2071 (N_2071,In_1796,In_2194);
or U2072 (N_2072,In_1570,In_2439);
and U2073 (N_2073,In_1141,In_1092);
nor U2074 (N_2074,In_331,In_1407);
xnor U2075 (N_2075,In_1888,In_1775);
xnor U2076 (N_2076,In_541,In_2405);
xnor U2077 (N_2077,In_1434,In_849);
xnor U2078 (N_2078,In_434,In_544);
or U2079 (N_2079,In_2128,In_1031);
nor U2080 (N_2080,In_696,In_505);
nor U2081 (N_2081,In_700,In_566);
nand U2082 (N_2082,In_338,In_1740);
and U2083 (N_2083,In_628,In_1137);
nor U2084 (N_2084,In_239,In_442);
nand U2085 (N_2085,In_1255,In_1838);
nor U2086 (N_2086,In_2396,In_2384);
nor U2087 (N_2087,In_3,In_1258);
and U2088 (N_2088,In_1313,In_37);
or U2089 (N_2089,In_630,In_1973);
and U2090 (N_2090,In_1108,In_2319);
xnor U2091 (N_2091,In_385,In_1011);
nand U2092 (N_2092,In_2120,In_29);
and U2093 (N_2093,In_55,In_487);
nor U2094 (N_2094,In_2203,In_1586);
nand U2095 (N_2095,In_2012,In_1332);
nor U2096 (N_2096,In_1861,In_2039);
or U2097 (N_2097,In_37,In_677);
or U2098 (N_2098,In_1945,In_1292);
and U2099 (N_2099,In_233,In_2305);
nor U2100 (N_2100,In_2411,In_2218);
nand U2101 (N_2101,In_629,In_2280);
and U2102 (N_2102,In_1700,In_1287);
nand U2103 (N_2103,In_2142,In_1991);
and U2104 (N_2104,In_2360,In_491);
nor U2105 (N_2105,In_20,In_300);
xnor U2106 (N_2106,In_1518,In_126);
and U2107 (N_2107,In_204,In_220);
and U2108 (N_2108,In_2489,In_1030);
nand U2109 (N_2109,In_914,In_1068);
and U2110 (N_2110,In_707,In_385);
or U2111 (N_2111,In_924,In_1913);
and U2112 (N_2112,In_1870,In_2029);
nor U2113 (N_2113,In_1386,In_1392);
xnor U2114 (N_2114,In_991,In_1355);
and U2115 (N_2115,In_781,In_404);
and U2116 (N_2116,In_875,In_1392);
and U2117 (N_2117,In_16,In_2111);
and U2118 (N_2118,In_1976,In_512);
or U2119 (N_2119,In_2086,In_121);
xnor U2120 (N_2120,In_497,In_2331);
xnor U2121 (N_2121,In_2464,In_1869);
and U2122 (N_2122,In_2161,In_1472);
nand U2123 (N_2123,In_2255,In_310);
or U2124 (N_2124,In_2395,In_1993);
or U2125 (N_2125,In_629,In_278);
and U2126 (N_2126,In_956,In_319);
nand U2127 (N_2127,In_617,In_1058);
xnor U2128 (N_2128,In_554,In_626);
or U2129 (N_2129,In_498,In_1887);
nand U2130 (N_2130,In_1265,In_2105);
and U2131 (N_2131,In_1363,In_866);
nand U2132 (N_2132,In_886,In_1163);
xnor U2133 (N_2133,In_700,In_466);
xnor U2134 (N_2134,In_1024,In_1199);
xnor U2135 (N_2135,In_893,In_1717);
nor U2136 (N_2136,In_869,In_1411);
nor U2137 (N_2137,In_246,In_1845);
and U2138 (N_2138,In_901,In_2376);
and U2139 (N_2139,In_2177,In_1790);
and U2140 (N_2140,In_1216,In_2436);
xnor U2141 (N_2141,In_2471,In_2169);
xnor U2142 (N_2142,In_2210,In_298);
or U2143 (N_2143,In_144,In_597);
and U2144 (N_2144,In_1163,In_1847);
xnor U2145 (N_2145,In_2341,In_1309);
xor U2146 (N_2146,In_1623,In_985);
and U2147 (N_2147,In_1498,In_1723);
xnor U2148 (N_2148,In_2376,In_1406);
or U2149 (N_2149,In_303,In_1458);
nand U2150 (N_2150,In_1771,In_1531);
xor U2151 (N_2151,In_1346,In_2243);
or U2152 (N_2152,In_502,In_2483);
nor U2153 (N_2153,In_1883,In_1572);
or U2154 (N_2154,In_212,In_1842);
or U2155 (N_2155,In_748,In_349);
and U2156 (N_2156,In_931,In_1805);
nand U2157 (N_2157,In_675,In_1875);
and U2158 (N_2158,In_849,In_693);
or U2159 (N_2159,In_2391,In_641);
or U2160 (N_2160,In_1755,In_1329);
and U2161 (N_2161,In_2483,In_1355);
nand U2162 (N_2162,In_1071,In_692);
nand U2163 (N_2163,In_1912,In_1391);
nor U2164 (N_2164,In_337,In_2);
or U2165 (N_2165,In_2000,In_74);
and U2166 (N_2166,In_1812,In_1901);
xnor U2167 (N_2167,In_2325,In_670);
nand U2168 (N_2168,In_1534,In_1684);
xor U2169 (N_2169,In_1185,In_2468);
and U2170 (N_2170,In_668,In_66);
nand U2171 (N_2171,In_1129,In_1831);
or U2172 (N_2172,In_2158,In_262);
nor U2173 (N_2173,In_643,In_58);
nor U2174 (N_2174,In_693,In_15);
nand U2175 (N_2175,In_498,In_2023);
xor U2176 (N_2176,In_686,In_2025);
nor U2177 (N_2177,In_1023,In_2235);
nand U2178 (N_2178,In_1915,In_1061);
nand U2179 (N_2179,In_430,In_1271);
nand U2180 (N_2180,In_2420,In_2139);
or U2181 (N_2181,In_2330,In_2205);
and U2182 (N_2182,In_30,In_2400);
or U2183 (N_2183,In_1395,In_863);
nand U2184 (N_2184,In_662,In_1800);
and U2185 (N_2185,In_1664,In_1316);
and U2186 (N_2186,In_2479,In_270);
nand U2187 (N_2187,In_2471,In_1795);
or U2188 (N_2188,In_1806,In_52);
nand U2189 (N_2189,In_2383,In_611);
xnor U2190 (N_2190,In_1950,In_330);
nor U2191 (N_2191,In_722,In_1034);
nand U2192 (N_2192,In_705,In_1362);
or U2193 (N_2193,In_1993,In_2283);
nand U2194 (N_2194,In_1659,In_247);
and U2195 (N_2195,In_1208,In_2498);
nand U2196 (N_2196,In_1594,In_1082);
and U2197 (N_2197,In_1035,In_1096);
nor U2198 (N_2198,In_2249,In_185);
and U2199 (N_2199,In_1573,In_2419);
and U2200 (N_2200,In_2254,In_2289);
xor U2201 (N_2201,In_331,In_469);
xnor U2202 (N_2202,In_323,In_1129);
or U2203 (N_2203,In_210,In_1740);
nor U2204 (N_2204,In_831,In_1787);
and U2205 (N_2205,In_1342,In_1829);
xnor U2206 (N_2206,In_2339,In_1852);
or U2207 (N_2207,In_2059,In_2335);
nor U2208 (N_2208,In_2147,In_861);
nand U2209 (N_2209,In_858,In_2319);
or U2210 (N_2210,In_1692,In_2250);
xnor U2211 (N_2211,In_2199,In_1913);
and U2212 (N_2212,In_851,In_421);
nand U2213 (N_2213,In_570,In_1763);
nor U2214 (N_2214,In_1981,In_1819);
nor U2215 (N_2215,In_1713,In_1540);
nand U2216 (N_2216,In_861,In_1044);
nor U2217 (N_2217,In_357,In_1231);
xnor U2218 (N_2218,In_1274,In_788);
or U2219 (N_2219,In_2279,In_1046);
or U2220 (N_2220,In_1089,In_1463);
nand U2221 (N_2221,In_1615,In_949);
nor U2222 (N_2222,In_1042,In_183);
nor U2223 (N_2223,In_850,In_992);
nand U2224 (N_2224,In_871,In_1874);
nor U2225 (N_2225,In_297,In_1616);
nor U2226 (N_2226,In_221,In_1981);
nor U2227 (N_2227,In_1864,In_791);
xor U2228 (N_2228,In_1045,In_1532);
nor U2229 (N_2229,In_1309,In_1888);
xor U2230 (N_2230,In_1294,In_328);
nand U2231 (N_2231,In_8,In_855);
and U2232 (N_2232,In_826,In_1745);
nor U2233 (N_2233,In_184,In_110);
nor U2234 (N_2234,In_2,In_1909);
nor U2235 (N_2235,In_2306,In_2345);
and U2236 (N_2236,In_19,In_895);
and U2237 (N_2237,In_2410,In_476);
nor U2238 (N_2238,In_1851,In_1219);
or U2239 (N_2239,In_1784,In_171);
or U2240 (N_2240,In_1603,In_543);
and U2241 (N_2241,In_1837,In_1950);
and U2242 (N_2242,In_751,In_141);
xor U2243 (N_2243,In_2000,In_960);
or U2244 (N_2244,In_1599,In_1552);
xor U2245 (N_2245,In_1416,In_1604);
or U2246 (N_2246,In_1611,In_897);
xnor U2247 (N_2247,In_138,In_1674);
xor U2248 (N_2248,In_1779,In_0);
and U2249 (N_2249,In_6,In_1165);
xor U2250 (N_2250,In_641,In_303);
xor U2251 (N_2251,In_649,In_1462);
and U2252 (N_2252,In_1496,In_1610);
nand U2253 (N_2253,In_587,In_2121);
xnor U2254 (N_2254,In_2007,In_567);
nor U2255 (N_2255,In_312,In_140);
and U2256 (N_2256,In_1529,In_2122);
xnor U2257 (N_2257,In_805,In_1669);
nor U2258 (N_2258,In_1427,In_755);
or U2259 (N_2259,In_533,In_1708);
or U2260 (N_2260,In_613,In_2409);
nor U2261 (N_2261,In_1913,In_2173);
nand U2262 (N_2262,In_2189,In_676);
and U2263 (N_2263,In_534,In_1170);
nand U2264 (N_2264,In_757,In_846);
nand U2265 (N_2265,In_1490,In_409);
xor U2266 (N_2266,In_2158,In_89);
and U2267 (N_2267,In_1490,In_2253);
nand U2268 (N_2268,In_530,In_470);
nand U2269 (N_2269,In_1401,In_830);
nand U2270 (N_2270,In_1648,In_1420);
nor U2271 (N_2271,In_672,In_768);
nand U2272 (N_2272,In_1182,In_2251);
xnor U2273 (N_2273,In_1066,In_716);
or U2274 (N_2274,In_825,In_65);
xnor U2275 (N_2275,In_218,In_988);
xnor U2276 (N_2276,In_1622,In_557);
or U2277 (N_2277,In_2150,In_2027);
nor U2278 (N_2278,In_1108,In_195);
nand U2279 (N_2279,In_967,In_1906);
nand U2280 (N_2280,In_2001,In_2489);
and U2281 (N_2281,In_1990,In_254);
nor U2282 (N_2282,In_997,In_573);
xor U2283 (N_2283,In_153,In_2447);
nand U2284 (N_2284,In_2006,In_2344);
or U2285 (N_2285,In_2203,In_2177);
and U2286 (N_2286,In_2335,In_2292);
xor U2287 (N_2287,In_695,In_561);
nand U2288 (N_2288,In_415,In_1209);
nor U2289 (N_2289,In_607,In_697);
nor U2290 (N_2290,In_1497,In_631);
or U2291 (N_2291,In_1668,In_1594);
nand U2292 (N_2292,In_817,In_2107);
nor U2293 (N_2293,In_1560,In_705);
or U2294 (N_2294,In_1220,In_1047);
nand U2295 (N_2295,In_138,In_1636);
and U2296 (N_2296,In_1477,In_1694);
nor U2297 (N_2297,In_34,In_1267);
xor U2298 (N_2298,In_19,In_946);
nor U2299 (N_2299,In_1275,In_1361);
and U2300 (N_2300,In_406,In_332);
nand U2301 (N_2301,In_828,In_1377);
or U2302 (N_2302,In_1734,In_246);
or U2303 (N_2303,In_1947,In_1345);
xor U2304 (N_2304,In_1159,In_1580);
and U2305 (N_2305,In_572,In_76);
nand U2306 (N_2306,In_530,In_2130);
and U2307 (N_2307,In_2467,In_726);
xnor U2308 (N_2308,In_1495,In_1729);
and U2309 (N_2309,In_2099,In_265);
nand U2310 (N_2310,In_722,In_1049);
xnor U2311 (N_2311,In_2260,In_1242);
or U2312 (N_2312,In_280,In_529);
xor U2313 (N_2313,In_2296,In_2387);
and U2314 (N_2314,In_454,In_260);
nand U2315 (N_2315,In_1758,In_1601);
xor U2316 (N_2316,In_1991,In_2455);
or U2317 (N_2317,In_372,In_1943);
or U2318 (N_2318,In_1089,In_2347);
nor U2319 (N_2319,In_2360,In_1762);
and U2320 (N_2320,In_144,In_1796);
xnor U2321 (N_2321,In_190,In_2427);
or U2322 (N_2322,In_1270,In_1142);
and U2323 (N_2323,In_2195,In_1560);
or U2324 (N_2324,In_220,In_2396);
xor U2325 (N_2325,In_517,In_899);
nor U2326 (N_2326,In_131,In_536);
and U2327 (N_2327,In_2067,In_1224);
and U2328 (N_2328,In_443,In_2116);
or U2329 (N_2329,In_780,In_1178);
or U2330 (N_2330,In_2025,In_2136);
nand U2331 (N_2331,In_829,In_76);
and U2332 (N_2332,In_1859,In_197);
nor U2333 (N_2333,In_1044,In_1022);
nor U2334 (N_2334,In_2037,In_482);
nor U2335 (N_2335,In_2091,In_2346);
xnor U2336 (N_2336,In_525,In_773);
xnor U2337 (N_2337,In_2030,In_655);
nand U2338 (N_2338,In_1995,In_1205);
xnor U2339 (N_2339,In_10,In_136);
or U2340 (N_2340,In_1732,In_1742);
nor U2341 (N_2341,In_2139,In_2413);
xor U2342 (N_2342,In_1443,In_2430);
nor U2343 (N_2343,In_68,In_486);
nor U2344 (N_2344,In_1975,In_44);
xor U2345 (N_2345,In_50,In_2455);
xor U2346 (N_2346,In_403,In_1435);
nand U2347 (N_2347,In_27,In_2065);
and U2348 (N_2348,In_183,In_629);
or U2349 (N_2349,In_787,In_747);
nor U2350 (N_2350,In_534,In_2356);
nand U2351 (N_2351,In_484,In_2132);
xor U2352 (N_2352,In_1534,In_1212);
xor U2353 (N_2353,In_2322,In_1290);
and U2354 (N_2354,In_1025,In_1787);
nor U2355 (N_2355,In_462,In_1196);
and U2356 (N_2356,In_18,In_122);
and U2357 (N_2357,In_35,In_261);
nand U2358 (N_2358,In_1152,In_2402);
or U2359 (N_2359,In_5,In_1616);
or U2360 (N_2360,In_1969,In_253);
and U2361 (N_2361,In_1756,In_1168);
or U2362 (N_2362,In_1424,In_1792);
and U2363 (N_2363,In_2243,In_1442);
nand U2364 (N_2364,In_2353,In_1928);
nand U2365 (N_2365,In_2100,In_1718);
nand U2366 (N_2366,In_1492,In_606);
nand U2367 (N_2367,In_2010,In_1893);
xnor U2368 (N_2368,In_2048,In_1599);
nand U2369 (N_2369,In_426,In_721);
nand U2370 (N_2370,In_1836,In_1608);
or U2371 (N_2371,In_1606,In_114);
and U2372 (N_2372,In_2334,In_2439);
xor U2373 (N_2373,In_2334,In_248);
nor U2374 (N_2374,In_2198,In_1540);
and U2375 (N_2375,In_2290,In_850);
or U2376 (N_2376,In_250,In_1791);
nor U2377 (N_2377,In_1112,In_472);
and U2378 (N_2378,In_1282,In_1444);
nor U2379 (N_2379,In_942,In_2096);
or U2380 (N_2380,In_200,In_206);
xnor U2381 (N_2381,In_2340,In_1819);
xor U2382 (N_2382,In_1838,In_18);
nor U2383 (N_2383,In_1520,In_1047);
xor U2384 (N_2384,In_2434,In_1223);
and U2385 (N_2385,In_1784,In_453);
or U2386 (N_2386,In_2139,In_1309);
nand U2387 (N_2387,In_2130,In_187);
and U2388 (N_2388,In_1467,In_1387);
or U2389 (N_2389,In_757,In_1405);
nand U2390 (N_2390,In_163,In_933);
nand U2391 (N_2391,In_667,In_800);
or U2392 (N_2392,In_2107,In_992);
and U2393 (N_2393,In_1788,In_1211);
nand U2394 (N_2394,In_2311,In_1247);
nand U2395 (N_2395,In_1450,In_725);
or U2396 (N_2396,In_1391,In_1938);
or U2397 (N_2397,In_1754,In_1627);
nor U2398 (N_2398,In_1406,In_1577);
nor U2399 (N_2399,In_1699,In_287);
or U2400 (N_2400,In_203,In_1177);
or U2401 (N_2401,In_1138,In_1817);
nor U2402 (N_2402,In_2055,In_263);
nand U2403 (N_2403,In_752,In_1489);
or U2404 (N_2404,In_928,In_1752);
and U2405 (N_2405,In_2302,In_1298);
and U2406 (N_2406,In_2106,In_127);
nor U2407 (N_2407,In_1226,In_1929);
xnor U2408 (N_2408,In_486,In_1762);
nor U2409 (N_2409,In_697,In_483);
xnor U2410 (N_2410,In_1450,In_672);
nand U2411 (N_2411,In_2340,In_1218);
xor U2412 (N_2412,In_1290,In_745);
or U2413 (N_2413,In_563,In_1156);
or U2414 (N_2414,In_992,In_2178);
nor U2415 (N_2415,In_2010,In_2313);
xnor U2416 (N_2416,In_32,In_1270);
nor U2417 (N_2417,In_1165,In_1527);
nor U2418 (N_2418,In_1663,In_173);
and U2419 (N_2419,In_1355,In_1528);
or U2420 (N_2420,In_181,In_1604);
and U2421 (N_2421,In_2302,In_224);
xnor U2422 (N_2422,In_1224,In_424);
nand U2423 (N_2423,In_114,In_2186);
xor U2424 (N_2424,In_1710,In_2333);
and U2425 (N_2425,In_24,In_1477);
or U2426 (N_2426,In_2053,In_2169);
nor U2427 (N_2427,In_929,In_1761);
nor U2428 (N_2428,In_1001,In_1767);
or U2429 (N_2429,In_2031,In_632);
nand U2430 (N_2430,In_56,In_1975);
nor U2431 (N_2431,In_2377,In_2164);
nor U2432 (N_2432,In_2469,In_1356);
or U2433 (N_2433,In_270,In_885);
nand U2434 (N_2434,In_2091,In_777);
nor U2435 (N_2435,In_997,In_1786);
xor U2436 (N_2436,In_2338,In_1170);
nand U2437 (N_2437,In_441,In_1607);
and U2438 (N_2438,In_1767,In_2247);
nand U2439 (N_2439,In_1381,In_1943);
xor U2440 (N_2440,In_1699,In_129);
nor U2441 (N_2441,In_1072,In_2094);
nor U2442 (N_2442,In_1277,In_119);
or U2443 (N_2443,In_1849,In_72);
or U2444 (N_2444,In_344,In_667);
xor U2445 (N_2445,In_1621,In_1749);
or U2446 (N_2446,In_952,In_1628);
nor U2447 (N_2447,In_2303,In_1314);
and U2448 (N_2448,In_1294,In_2221);
nand U2449 (N_2449,In_838,In_9);
nor U2450 (N_2450,In_2356,In_477);
nor U2451 (N_2451,In_401,In_6);
xnor U2452 (N_2452,In_996,In_1787);
nand U2453 (N_2453,In_2469,In_2427);
nand U2454 (N_2454,In_277,In_67);
nand U2455 (N_2455,In_2153,In_2076);
nor U2456 (N_2456,In_1019,In_744);
nand U2457 (N_2457,In_938,In_1032);
or U2458 (N_2458,In_2384,In_467);
nor U2459 (N_2459,In_668,In_1277);
xnor U2460 (N_2460,In_1941,In_1152);
nand U2461 (N_2461,In_416,In_2358);
xor U2462 (N_2462,In_2115,In_2049);
xnor U2463 (N_2463,In_2118,In_561);
xnor U2464 (N_2464,In_1463,In_894);
nand U2465 (N_2465,In_1464,In_168);
nand U2466 (N_2466,In_980,In_1680);
or U2467 (N_2467,In_904,In_2024);
nand U2468 (N_2468,In_1892,In_1063);
nor U2469 (N_2469,In_1186,In_1471);
and U2470 (N_2470,In_557,In_2018);
and U2471 (N_2471,In_1517,In_2262);
or U2472 (N_2472,In_823,In_1700);
nor U2473 (N_2473,In_864,In_55);
nand U2474 (N_2474,In_1942,In_2146);
xor U2475 (N_2475,In_1117,In_632);
xor U2476 (N_2476,In_2129,In_1000);
nor U2477 (N_2477,In_2311,In_620);
or U2478 (N_2478,In_2275,In_645);
nor U2479 (N_2479,In_569,In_510);
nor U2480 (N_2480,In_1241,In_1563);
or U2481 (N_2481,In_2380,In_2223);
nor U2482 (N_2482,In_1706,In_1061);
and U2483 (N_2483,In_2366,In_506);
or U2484 (N_2484,In_1159,In_464);
and U2485 (N_2485,In_85,In_1962);
xor U2486 (N_2486,In_1145,In_1605);
or U2487 (N_2487,In_506,In_1231);
nand U2488 (N_2488,In_1115,In_2497);
xnor U2489 (N_2489,In_2041,In_891);
and U2490 (N_2490,In_454,In_653);
nand U2491 (N_2491,In_1306,In_2289);
xor U2492 (N_2492,In_1284,In_1774);
xor U2493 (N_2493,In_1122,In_2343);
xor U2494 (N_2494,In_1449,In_549);
nor U2495 (N_2495,In_577,In_2452);
nor U2496 (N_2496,In_851,In_89);
nand U2497 (N_2497,In_1813,In_1396);
xor U2498 (N_2498,In_293,In_2436);
xnor U2499 (N_2499,In_987,In_145);
xor U2500 (N_2500,In_628,In_957);
xnor U2501 (N_2501,In_2240,In_1751);
or U2502 (N_2502,In_991,In_2373);
xor U2503 (N_2503,In_1361,In_591);
nand U2504 (N_2504,In_363,In_9);
nand U2505 (N_2505,In_2297,In_2366);
and U2506 (N_2506,In_1752,In_622);
nand U2507 (N_2507,In_2082,In_751);
xor U2508 (N_2508,In_1377,In_2031);
nand U2509 (N_2509,In_537,In_431);
or U2510 (N_2510,In_1564,In_517);
nor U2511 (N_2511,In_1493,In_1329);
nor U2512 (N_2512,In_1989,In_537);
nand U2513 (N_2513,In_1219,In_2064);
nand U2514 (N_2514,In_642,In_263);
or U2515 (N_2515,In_384,In_2015);
nand U2516 (N_2516,In_985,In_1667);
or U2517 (N_2517,In_710,In_884);
nand U2518 (N_2518,In_1267,In_230);
nand U2519 (N_2519,In_2323,In_1944);
or U2520 (N_2520,In_1183,In_1670);
and U2521 (N_2521,In_1274,In_2091);
and U2522 (N_2522,In_2388,In_1893);
or U2523 (N_2523,In_2082,In_2351);
or U2524 (N_2524,In_1284,In_547);
nand U2525 (N_2525,In_11,In_1204);
or U2526 (N_2526,In_1939,In_1769);
nand U2527 (N_2527,In_779,In_759);
nand U2528 (N_2528,In_859,In_982);
xor U2529 (N_2529,In_2365,In_1928);
or U2530 (N_2530,In_2387,In_165);
xnor U2531 (N_2531,In_204,In_1547);
nor U2532 (N_2532,In_187,In_2175);
and U2533 (N_2533,In_1058,In_1585);
xor U2534 (N_2534,In_544,In_1609);
xor U2535 (N_2535,In_2257,In_634);
and U2536 (N_2536,In_115,In_1656);
xor U2537 (N_2537,In_1051,In_1610);
and U2538 (N_2538,In_229,In_1737);
xnor U2539 (N_2539,In_1777,In_1079);
nand U2540 (N_2540,In_1729,In_1316);
nor U2541 (N_2541,In_1856,In_2242);
nor U2542 (N_2542,In_611,In_1475);
and U2543 (N_2543,In_2308,In_983);
xnor U2544 (N_2544,In_1088,In_1386);
or U2545 (N_2545,In_511,In_1339);
nor U2546 (N_2546,In_80,In_1951);
nand U2547 (N_2547,In_784,In_1917);
or U2548 (N_2548,In_2308,In_365);
nor U2549 (N_2549,In_742,In_1434);
nor U2550 (N_2550,In_36,In_248);
nand U2551 (N_2551,In_908,In_2065);
or U2552 (N_2552,In_1961,In_1634);
or U2553 (N_2553,In_379,In_1032);
and U2554 (N_2554,In_784,In_2350);
nor U2555 (N_2555,In_848,In_262);
or U2556 (N_2556,In_995,In_632);
and U2557 (N_2557,In_1081,In_385);
and U2558 (N_2558,In_1662,In_1390);
xor U2559 (N_2559,In_1880,In_1649);
xnor U2560 (N_2560,In_283,In_1384);
xnor U2561 (N_2561,In_541,In_1828);
nand U2562 (N_2562,In_88,In_1796);
nor U2563 (N_2563,In_1633,In_2297);
xor U2564 (N_2564,In_1513,In_808);
nor U2565 (N_2565,In_2120,In_1208);
xor U2566 (N_2566,In_2010,In_1174);
xnor U2567 (N_2567,In_2229,In_187);
nand U2568 (N_2568,In_410,In_306);
and U2569 (N_2569,In_503,In_1470);
xnor U2570 (N_2570,In_646,In_556);
and U2571 (N_2571,In_2394,In_2209);
and U2572 (N_2572,In_1390,In_1714);
or U2573 (N_2573,In_1190,In_618);
nor U2574 (N_2574,In_2190,In_332);
nor U2575 (N_2575,In_1304,In_1928);
nand U2576 (N_2576,In_1397,In_1634);
xnor U2577 (N_2577,In_515,In_20);
or U2578 (N_2578,In_1418,In_2416);
nand U2579 (N_2579,In_899,In_2461);
nand U2580 (N_2580,In_1285,In_2061);
and U2581 (N_2581,In_1022,In_93);
or U2582 (N_2582,In_1165,In_769);
nor U2583 (N_2583,In_712,In_1702);
and U2584 (N_2584,In_1630,In_2129);
nand U2585 (N_2585,In_1535,In_1269);
or U2586 (N_2586,In_1811,In_714);
nor U2587 (N_2587,In_2315,In_2121);
and U2588 (N_2588,In_1719,In_1078);
nor U2589 (N_2589,In_1057,In_993);
nand U2590 (N_2590,In_1296,In_1662);
nor U2591 (N_2591,In_618,In_2413);
xnor U2592 (N_2592,In_1459,In_1158);
xor U2593 (N_2593,In_2072,In_1354);
or U2594 (N_2594,In_1007,In_332);
and U2595 (N_2595,In_2025,In_1915);
nor U2596 (N_2596,In_1704,In_2301);
and U2597 (N_2597,In_1964,In_974);
and U2598 (N_2598,In_1974,In_1673);
and U2599 (N_2599,In_1223,In_1101);
xnor U2600 (N_2600,In_1905,In_72);
xnor U2601 (N_2601,In_1070,In_726);
nand U2602 (N_2602,In_404,In_1915);
nor U2603 (N_2603,In_232,In_445);
nor U2604 (N_2604,In_1298,In_2442);
nand U2605 (N_2605,In_1904,In_384);
nand U2606 (N_2606,In_2117,In_1814);
and U2607 (N_2607,In_1916,In_1870);
or U2608 (N_2608,In_295,In_856);
xor U2609 (N_2609,In_2440,In_2223);
nor U2610 (N_2610,In_2369,In_290);
and U2611 (N_2611,In_2295,In_1983);
nand U2612 (N_2612,In_518,In_1811);
or U2613 (N_2613,In_62,In_1298);
xnor U2614 (N_2614,In_341,In_697);
or U2615 (N_2615,In_1984,In_2040);
xor U2616 (N_2616,In_2178,In_2290);
nor U2617 (N_2617,In_148,In_901);
xor U2618 (N_2618,In_1700,In_35);
nand U2619 (N_2619,In_2043,In_919);
nor U2620 (N_2620,In_1240,In_1473);
nand U2621 (N_2621,In_2391,In_1111);
xor U2622 (N_2622,In_769,In_2138);
and U2623 (N_2623,In_1706,In_618);
nand U2624 (N_2624,In_2127,In_983);
or U2625 (N_2625,In_2216,In_2448);
xor U2626 (N_2626,In_1704,In_2052);
xnor U2627 (N_2627,In_2096,In_897);
xor U2628 (N_2628,In_753,In_804);
and U2629 (N_2629,In_1159,In_2095);
nand U2630 (N_2630,In_2334,In_763);
or U2631 (N_2631,In_181,In_12);
and U2632 (N_2632,In_524,In_1034);
nand U2633 (N_2633,In_1235,In_1209);
or U2634 (N_2634,In_1384,In_107);
and U2635 (N_2635,In_1643,In_1632);
nor U2636 (N_2636,In_499,In_679);
or U2637 (N_2637,In_1715,In_1004);
nand U2638 (N_2638,In_792,In_2401);
nor U2639 (N_2639,In_1629,In_1086);
or U2640 (N_2640,In_2305,In_1684);
nor U2641 (N_2641,In_945,In_1505);
nand U2642 (N_2642,In_97,In_435);
nand U2643 (N_2643,In_229,In_1270);
and U2644 (N_2644,In_1019,In_862);
and U2645 (N_2645,In_695,In_1140);
or U2646 (N_2646,In_296,In_685);
xor U2647 (N_2647,In_1676,In_286);
nand U2648 (N_2648,In_534,In_1714);
and U2649 (N_2649,In_1068,In_1536);
nor U2650 (N_2650,In_1477,In_306);
xor U2651 (N_2651,In_1018,In_242);
nor U2652 (N_2652,In_1116,In_208);
nand U2653 (N_2653,In_2499,In_2149);
nor U2654 (N_2654,In_611,In_1809);
xnor U2655 (N_2655,In_425,In_923);
xnor U2656 (N_2656,In_926,In_1833);
nor U2657 (N_2657,In_837,In_536);
or U2658 (N_2658,In_2103,In_1620);
nor U2659 (N_2659,In_1522,In_1785);
xnor U2660 (N_2660,In_1111,In_1525);
xor U2661 (N_2661,In_652,In_1714);
nor U2662 (N_2662,In_1756,In_354);
nand U2663 (N_2663,In_351,In_442);
nand U2664 (N_2664,In_137,In_1365);
nor U2665 (N_2665,In_2209,In_553);
xor U2666 (N_2666,In_76,In_1266);
and U2667 (N_2667,In_1969,In_1440);
or U2668 (N_2668,In_2375,In_1006);
nand U2669 (N_2669,In_1387,In_382);
and U2670 (N_2670,In_2149,In_1463);
nand U2671 (N_2671,In_2416,In_1067);
nand U2672 (N_2672,In_1158,In_108);
and U2673 (N_2673,In_61,In_182);
nor U2674 (N_2674,In_380,In_1562);
and U2675 (N_2675,In_1196,In_89);
nor U2676 (N_2676,In_1490,In_2045);
xor U2677 (N_2677,In_83,In_1268);
nand U2678 (N_2678,In_627,In_668);
nand U2679 (N_2679,In_865,In_1329);
nor U2680 (N_2680,In_1211,In_822);
xnor U2681 (N_2681,In_1868,In_2033);
or U2682 (N_2682,In_535,In_2026);
and U2683 (N_2683,In_354,In_1102);
nand U2684 (N_2684,In_2197,In_487);
xor U2685 (N_2685,In_1270,In_868);
xor U2686 (N_2686,In_1313,In_429);
nand U2687 (N_2687,In_1196,In_1704);
nor U2688 (N_2688,In_777,In_381);
or U2689 (N_2689,In_754,In_2144);
or U2690 (N_2690,In_2322,In_1691);
xnor U2691 (N_2691,In_520,In_1638);
or U2692 (N_2692,In_1641,In_1538);
nor U2693 (N_2693,In_2172,In_150);
xor U2694 (N_2694,In_1898,In_1735);
xnor U2695 (N_2695,In_190,In_612);
nand U2696 (N_2696,In_1869,In_1613);
nor U2697 (N_2697,In_178,In_262);
nor U2698 (N_2698,In_656,In_2333);
nand U2699 (N_2699,In_2398,In_2029);
nand U2700 (N_2700,In_141,In_1914);
or U2701 (N_2701,In_146,In_556);
and U2702 (N_2702,In_1973,In_2157);
nor U2703 (N_2703,In_2051,In_851);
xnor U2704 (N_2704,In_1268,In_221);
or U2705 (N_2705,In_355,In_2425);
nand U2706 (N_2706,In_1262,In_2229);
nor U2707 (N_2707,In_1776,In_1985);
or U2708 (N_2708,In_782,In_2153);
nand U2709 (N_2709,In_1618,In_49);
nand U2710 (N_2710,In_1210,In_2192);
or U2711 (N_2711,In_264,In_1067);
xor U2712 (N_2712,In_1591,In_2452);
nand U2713 (N_2713,In_1853,In_70);
xor U2714 (N_2714,In_54,In_606);
nand U2715 (N_2715,In_2116,In_781);
or U2716 (N_2716,In_580,In_946);
xor U2717 (N_2717,In_1647,In_2014);
and U2718 (N_2718,In_529,In_473);
nor U2719 (N_2719,In_1735,In_870);
and U2720 (N_2720,In_274,In_354);
or U2721 (N_2721,In_741,In_650);
nand U2722 (N_2722,In_125,In_1727);
nor U2723 (N_2723,In_633,In_2437);
nand U2724 (N_2724,In_762,In_2037);
nor U2725 (N_2725,In_2228,In_253);
or U2726 (N_2726,In_650,In_631);
and U2727 (N_2727,In_1476,In_12);
xor U2728 (N_2728,In_1532,In_333);
xnor U2729 (N_2729,In_1074,In_1884);
nand U2730 (N_2730,In_623,In_1592);
xnor U2731 (N_2731,In_990,In_2152);
nor U2732 (N_2732,In_694,In_156);
and U2733 (N_2733,In_1618,In_117);
and U2734 (N_2734,In_1419,In_1042);
xor U2735 (N_2735,In_1240,In_701);
nor U2736 (N_2736,In_2174,In_1162);
nand U2737 (N_2737,In_1958,In_1819);
and U2738 (N_2738,In_905,In_1448);
nand U2739 (N_2739,In_1387,In_1436);
and U2740 (N_2740,In_599,In_93);
nand U2741 (N_2741,In_904,In_2333);
nand U2742 (N_2742,In_1168,In_1823);
and U2743 (N_2743,In_2471,In_124);
nor U2744 (N_2744,In_1736,In_802);
nor U2745 (N_2745,In_1624,In_1634);
nor U2746 (N_2746,In_368,In_2139);
nand U2747 (N_2747,In_132,In_1875);
or U2748 (N_2748,In_1510,In_1000);
or U2749 (N_2749,In_184,In_1878);
xnor U2750 (N_2750,In_2352,In_299);
nand U2751 (N_2751,In_649,In_316);
nor U2752 (N_2752,In_171,In_2013);
xor U2753 (N_2753,In_2388,In_1813);
or U2754 (N_2754,In_428,In_2243);
nor U2755 (N_2755,In_1434,In_1592);
or U2756 (N_2756,In_1638,In_2317);
nor U2757 (N_2757,In_804,In_1520);
xor U2758 (N_2758,In_2207,In_783);
and U2759 (N_2759,In_1522,In_2339);
or U2760 (N_2760,In_779,In_1391);
nor U2761 (N_2761,In_1229,In_505);
nand U2762 (N_2762,In_1803,In_1392);
xor U2763 (N_2763,In_2010,In_1568);
and U2764 (N_2764,In_371,In_560);
and U2765 (N_2765,In_1833,In_530);
xor U2766 (N_2766,In_1704,In_66);
or U2767 (N_2767,In_185,In_2096);
xnor U2768 (N_2768,In_1669,In_1644);
xnor U2769 (N_2769,In_1165,In_2298);
xnor U2770 (N_2770,In_2391,In_529);
nand U2771 (N_2771,In_2488,In_1773);
or U2772 (N_2772,In_386,In_2461);
nand U2773 (N_2773,In_396,In_960);
nand U2774 (N_2774,In_2416,In_755);
or U2775 (N_2775,In_884,In_673);
nand U2776 (N_2776,In_1539,In_260);
nand U2777 (N_2777,In_5,In_167);
or U2778 (N_2778,In_2056,In_648);
or U2779 (N_2779,In_751,In_1232);
or U2780 (N_2780,In_2000,In_2451);
and U2781 (N_2781,In_916,In_1552);
nand U2782 (N_2782,In_777,In_1646);
or U2783 (N_2783,In_615,In_1689);
xnor U2784 (N_2784,In_2162,In_671);
or U2785 (N_2785,In_978,In_2410);
or U2786 (N_2786,In_482,In_1417);
nand U2787 (N_2787,In_200,In_816);
or U2788 (N_2788,In_1735,In_931);
xnor U2789 (N_2789,In_628,In_253);
or U2790 (N_2790,In_1184,In_1095);
and U2791 (N_2791,In_2092,In_1392);
or U2792 (N_2792,In_1290,In_1332);
or U2793 (N_2793,In_1969,In_2334);
and U2794 (N_2794,In_2353,In_593);
xnor U2795 (N_2795,In_1972,In_192);
xor U2796 (N_2796,In_1733,In_980);
nor U2797 (N_2797,In_533,In_1469);
xnor U2798 (N_2798,In_1479,In_836);
nand U2799 (N_2799,In_1881,In_361);
nor U2800 (N_2800,In_1134,In_1736);
and U2801 (N_2801,In_1165,In_1215);
or U2802 (N_2802,In_23,In_777);
xor U2803 (N_2803,In_1618,In_582);
xnor U2804 (N_2804,In_1991,In_2361);
nand U2805 (N_2805,In_276,In_653);
nor U2806 (N_2806,In_1404,In_668);
or U2807 (N_2807,In_2092,In_1820);
xor U2808 (N_2808,In_794,In_159);
nand U2809 (N_2809,In_1072,In_2299);
nor U2810 (N_2810,In_1511,In_355);
nand U2811 (N_2811,In_1011,In_167);
nor U2812 (N_2812,In_1624,In_539);
nand U2813 (N_2813,In_678,In_1275);
or U2814 (N_2814,In_2125,In_658);
nor U2815 (N_2815,In_838,In_1301);
and U2816 (N_2816,In_242,In_973);
nor U2817 (N_2817,In_1698,In_1584);
nor U2818 (N_2818,In_603,In_1922);
xnor U2819 (N_2819,In_2439,In_2200);
nor U2820 (N_2820,In_1131,In_1355);
or U2821 (N_2821,In_705,In_596);
and U2822 (N_2822,In_1237,In_602);
xor U2823 (N_2823,In_1172,In_1404);
nor U2824 (N_2824,In_982,In_5);
xor U2825 (N_2825,In_536,In_730);
nor U2826 (N_2826,In_433,In_1618);
nand U2827 (N_2827,In_1290,In_1033);
and U2828 (N_2828,In_1256,In_2220);
nor U2829 (N_2829,In_2269,In_1824);
nand U2830 (N_2830,In_2416,In_795);
or U2831 (N_2831,In_888,In_1585);
nand U2832 (N_2832,In_639,In_1314);
or U2833 (N_2833,In_118,In_350);
nor U2834 (N_2834,In_797,In_537);
xor U2835 (N_2835,In_575,In_179);
or U2836 (N_2836,In_1688,In_168);
xnor U2837 (N_2837,In_231,In_125);
xnor U2838 (N_2838,In_68,In_640);
or U2839 (N_2839,In_106,In_423);
or U2840 (N_2840,In_1003,In_1958);
and U2841 (N_2841,In_2081,In_1918);
or U2842 (N_2842,In_973,In_2018);
and U2843 (N_2843,In_626,In_1904);
xor U2844 (N_2844,In_2145,In_2222);
nand U2845 (N_2845,In_2495,In_555);
nand U2846 (N_2846,In_739,In_2106);
and U2847 (N_2847,In_944,In_2417);
or U2848 (N_2848,In_2374,In_736);
nand U2849 (N_2849,In_1051,In_2039);
nand U2850 (N_2850,In_135,In_261);
and U2851 (N_2851,In_386,In_1900);
nand U2852 (N_2852,In_1491,In_671);
xnor U2853 (N_2853,In_1543,In_25);
and U2854 (N_2854,In_392,In_1139);
nor U2855 (N_2855,In_666,In_1489);
xor U2856 (N_2856,In_1140,In_2278);
and U2857 (N_2857,In_1543,In_718);
nor U2858 (N_2858,In_1741,In_423);
nor U2859 (N_2859,In_308,In_2136);
nor U2860 (N_2860,In_584,In_1260);
nand U2861 (N_2861,In_1256,In_502);
or U2862 (N_2862,In_1874,In_351);
xnor U2863 (N_2863,In_1520,In_2284);
or U2864 (N_2864,In_2137,In_1119);
and U2865 (N_2865,In_971,In_1630);
nand U2866 (N_2866,In_2165,In_1347);
nand U2867 (N_2867,In_1595,In_2283);
nor U2868 (N_2868,In_1275,In_1281);
nor U2869 (N_2869,In_1037,In_1968);
and U2870 (N_2870,In_190,In_1598);
nand U2871 (N_2871,In_638,In_1146);
nor U2872 (N_2872,In_671,In_1711);
nor U2873 (N_2873,In_2209,In_1515);
or U2874 (N_2874,In_417,In_2159);
or U2875 (N_2875,In_479,In_933);
nor U2876 (N_2876,In_1998,In_1054);
or U2877 (N_2877,In_160,In_1270);
nor U2878 (N_2878,In_94,In_616);
xor U2879 (N_2879,In_864,In_1917);
xnor U2880 (N_2880,In_782,In_1463);
xnor U2881 (N_2881,In_168,In_1567);
or U2882 (N_2882,In_1807,In_1820);
nand U2883 (N_2883,In_1120,In_98);
nand U2884 (N_2884,In_1681,In_2043);
nor U2885 (N_2885,In_1794,In_116);
xor U2886 (N_2886,In_1074,In_559);
nor U2887 (N_2887,In_624,In_1337);
nor U2888 (N_2888,In_1126,In_1440);
nand U2889 (N_2889,In_399,In_1548);
nor U2890 (N_2890,In_2219,In_1084);
xor U2891 (N_2891,In_2018,In_1143);
xnor U2892 (N_2892,In_486,In_1644);
and U2893 (N_2893,In_320,In_450);
or U2894 (N_2894,In_601,In_1766);
and U2895 (N_2895,In_2046,In_1261);
nand U2896 (N_2896,In_197,In_1207);
xnor U2897 (N_2897,In_1266,In_1462);
and U2898 (N_2898,In_226,In_723);
or U2899 (N_2899,In_712,In_1582);
nand U2900 (N_2900,In_880,In_1846);
xnor U2901 (N_2901,In_1487,In_394);
nand U2902 (N_2902,In_1034,In_614);
nor U2903 (N_2903,In_2315,In_827);
or U2904 (N_2904,In_60,In_1685);
and U2905 (N_2905,In_1553,In_231);
and U2906 (N_2906,In_993,In_740);
nor U2907 (N_2907,In_925,In_1093);
xnor U2908 (N_2908,In_1801,In_2018);
nand U2909 (N_2909,In_576,In_2250);
and U2910 (N_2910,In_1672,In_2491);
xor U2911 (N_2911,In_647,In_576);
nor U2912 (N_2912,In_2437,In_2151);
or U2913 (N_2913,In_916,In_774);
or U2914 (N_2914,In_2198,In_886);
and U2915 (N_2915,In_17,In_236);
nand U2916 (N_2916,In_1644,In_1942);
nor U2917 (N_2917,In_1321,In_783);
or U2918 (N_2918,In_263,In_1200);
xnor U2919 (N_2919,In_2406,In_160);
or U2920 (N_2920,In_1364,In_1935);
or U2921 (N_2921,In_1471,In_1769);
nor U2922 (N_2922,In_959,In_2441);
and U2923 (N_2923,In_723,In_2205);
xnor U2924 (N_2924,In_1011,In_1849);
nor U2925 (N_2925,In_2482,In_756);
and U2926 (N_2926,In_494,In_140);
or U2927 (N_2927,In_537,In_1684);
nand U2928 (N_2928,In_1093,In_1124);
nor U2929 (N_2929,In_2300,In_605);
nand U2930 (N_2930,In_2207,In_1424);
and U2931 (N_2931,In_1693,In_1645);
and U2932 (N_2932,In_75,In_1720);
nor U2933 (N_2933,In_2213,In_105);
nor U2934 (N_2934,In_555,In_63);
nand U2935 (N_2935,In_1033,In_909);
xor U2936 (N_2936,In_1793,In_113);
xor U2937 (N_2937,In_2070,In_605);
or U2938 (N_2938,In_287,In_922);
and U2939 (N_2939,In_1237,In_1876);
nor U2940 (N_2940,In_613,In_1046);
xor U2941 (N_2941,In_502,In_1574);
xnor U2942 (N_2942,In_2176,In_451);
nor U2943 (N_2943,In_1854,In_1107);
xnor U2944 (N_2944,In_970,In_1111);
and U2945 (N_2945,In_704,In_609);
and U2946 (N_2946,In_2082,In_2135);
or U2947 (N_2947,In_266,In_2472);
xnor U2948 (N_2948,In_1750,In_1652);
and U2949 (N_2949,In_289,In_506);
and U2950 (N_2950,In_534,In_199);
or U2951 (N_2951,In_1524,In_514);
nor U2952 (N_2952,In_1358,In_1841);
nor U2953 (N_2953,In_1477,In_326);
or U2954 (N_2954,In_224,In_933);
nor U2955 (N_2955,In_559,In_254);
and U2956 (N_2956,In_838,In_1625);
xnor U2957 (N_2957,In_272,In_2347);
or U2958 (N_2958,In_437,In_1022);
xor U2959 (N_2959,In_2326,In_1220);
nand U2960 (N_2960,In_2224,In_130);
nor U2961 (N_2961,In_514,In_1958);
or U2962 (N_2962,In_1901,In_1540);
nand U2963 (N_2963,In_1882,In_410);
xor U2964 (N_2964,In_13,In_833);
xnor U2965 (N_2965,In_1309,In_1873);
nand U2966 (N_2966,In_1226,In_1262);
xnor U2967 (N_2967,In_443,In_1790);
nor U2968 (N_2968,In_1796,In_2106);
and U2969 (N_2969,In_2368,In_629);
or U2970 (N_2970,In_1725,In_1874);
nand U2971 (N_2971,In_135,In_182);
xnor U2972 (N_2972,In_254,In_1360);
xnor U2973 (N_2973,In_1683,In_1024);
and U2974 (N_2974,In_186,In_672);
or U2975 (N_2975,In_869,In_1671);
nor U2976 (N_2976,In_1443,In_262);
nand U2977 (N_2977,In_2256,In_627);
nand U2978 (N_2978,In_2374,In_2259);
or U2979 (N_2979,In_2187,In_1604);
xnor U2980 (N_2980,In_2444,In_238);
nor U2981 (N_2981,In_1764,In_1282);
xnor U2982 (N_2982,In_1667,In_2146);
xnor U2983 (N_2983,In_1636,In_2012);
and U2984 (N_2984,In_1900,In_1140);
xor U2985 (N_2985,In_935,In_2332);
nor U2986 (N_2986,In_708,In_795);
nor U2987 (N_2987,In_376,In_1529);
xnor U2988 (N_2988,In_1784,In_2219);
or U2989 (N_2989,In_147,In_1412);
or U2990 (N_2990,In_510,In_2466);
or U2991 (N_2991,In_1581,In_2158);
and U2992 (N_2992,In_1568,In_2047);
xor U2993 (N_2993,In_353,In_1828);
or U2994 (N_2994,In_874,In_1138);
nor U2995 (N_2995,In_2123,In_2160);
nor U2996 (N_2996,In_1830,In_1173);
or U2997 (N_2997,In_377,In_1362);
and U2998 (N_2998,In_1258,In_79);
nor U2999 (N_2999,In_828,In_294);
nor U3000 (N_3000,In_1117,In_936);
nor U3001 (N_3001,In_188,In_2302);
nand U3002 (N_3002,In_1579,In_1331);
nand U3003 (N_3003,In_1563,In_2150);
nor U3004 (N_3004,In_781,In_917);
and U3005 (N_3005,In_430,In_2083);
or U3006 (N_3006,In_739,In_456);
xor U3007 (N_3007,In_2276,In_889);
nor U3008 (N_3008,In_2337,In_2168);
nor U3009 (N_3009,In_2346,In_2224);
nor U3010 (N_3010,In_930,In_413);
and U3011 (N_3011,In_867,In_721);
nand U3012 (N_3012,In_852,In_1247);
and U3013 (N_3013,In_1238,In_265);
or U3014 (N_3014,In_184,In_486);
and U3015 (N_3015,In_136,In_484);
nor U3016 (N_3016,In_1703,In_723);
or U3017 (N_3017,In_1800,In_1745);
and U3018 (N_3018,In_1470,In_1103);
or U3019 (N_3019,In_176,In_1755);
nand U3020 (N_3020,In_1519,In_93);
and U3021 (N_3021,In_1640,In_960);
or U3022 (N_3022,In_2082,In_392);
or U3023 (N_3023,In_2167,In_914);
and U3024 (N_3024,In_301,In_1581);
or U3025 (N_3025,In_1311,In_1256);
and U3026 (N_3026,In_1800,In_160);
or U3027 (N_3027,In_521,In_514);
nor U3028 (N_3028,In_1880,In_1170);
nor U3029 (N_3029,In_1494,In_1374);
xnor U3030 (N_3030,In_2350,In_1826);
xor U3031 (N_3031,In_1690,In_189);
xnor U3032 (N_3032,In_299,In_68);
xnor U3033 (N_3033,In_2339,In_1488);
nand U3034 (N_3034,In_1593,In_2052);
xnor U3035 (N_3035,In_1965,In_151);
and U3036 (N_3036,In_1478,In_1010);
nor U3037 (N_3037,In_625,In_2312);
or U3038 (N_3038,In_856,In_1884);
nor U3039 (N_3039,In_512,In_2204);
and U3040 (N_3040,In_788,In_349);
and U3041 (N_3041,In_332,In_1395);
or U3042 (N_3042,In_2231,In_60);
xor U3043 (N_3043,In_1036,In_1354);
xnor U3044 (N_3044,In_502,In_1477);
and U3045 (N_3045,In_2349,In_1756);
nand U3046 (N_3046,In_1235,In_72);
nand U3047 (N_3047,In_1966,In_2181);
xor U3048 (N_3048,In_1984,In_933);
xnor U3049 (N_3049,In_1627,In_1913);
xnor U3050 (N_3050,In_1480,In_1818);
nand U3051 (N_3051,In_833,In_1115);
and U3052 (N_3052,In_559,In_1108);
and U3053 (N_3053,In_908,In_958);
nor U3054 (N_3054,In_560,In_2111);
and U3055 (N_3055,In_2083,In_530);
nand U3056 (N_3056,In_2028,In_1154);
nor U3057 (N_3057,In_138,In_1707);
xor U3058 (N_3058,In_1325,In_2053);
or U3059 (N_3059,In_362,In_676);
xor U3060 (N_3060,In_1394,In_1077);
xnor U3061 (N_3061,In_1004,In_273);
nand U3062 (N_3062,In_583,In_965);
and U3063 (N_3063,In_342,In_1830);
xnor U3064 (N_3064,In_50,In_2163);
xnor U3065 (N_3065,In_234,In_2274);
xnor U3066 (N_3066,In_241,In_1263);
xnor U3067 (N_3067,In_1650,In_2056);
or U3068 (N_3068,In_2090,In_2202);
or U3069 (N_3069,In_2449,In_425);
nand U3070 (N_3070,In_131,In_2347);
nor U3071 (N_3071,In_341,In_1817);
nand U3072 (N_3072,In_1963,In_196);
nand U3073 (N_3073,In_227,In_1338);
and U3074 (N_3074,In_1659,In_1165);
or U3075 (N_3075,In_248,In_226);
nand U3076 (N_3076,In_2027,In_660);
xor U3077 (N_3077,In_2399,In_2104);
and U3078 (N_3078,In_1378,In_1629);
xor U3079 (N_3079,In_4,In_666);
or U3080 (N_3080,In_463,In_1123);
xor U3081 (N_3081,In_2065,In_109);
or U3082 (N_3082,In_1176,In_689);
or U3083 (N_3083,In_1335,In_335);
or U3084 (N_3084,In_2237,In_2494);
and U3085 (N_3085,In_1795,In_1452);
nand U3086 (N_3086,In_1803,In_525);
xor U3087 (N_3087,In_555,In_2496);
nand U3088 (N_3088,In_2049,In_259);
nor U3089 (N_3089,In_1911,In_2476);
and U3090 (N_3090,In_586,In_339);
nor U3091 (N_3091,In_2262,In_1963);
nor U3092 (N_3092,In_96,In_753);
xnor U3093 (N_3093,In_2410,In_1672);
nor U3094 (N_3094,In_1389,In_1392);
xor U3095 (N_3095,In_1185,In_1039);
and U3096 (N_3096,In_2009,In_1490);
and U3097 (N_3097,In_1112,In_1621);
xor U3098 (N_3098,In_1148,In_971);
nor U3099 (N_3099,In_2033,In_1522);
and U3100 (N_3100,In_1902,In_1841);
nor U3101 (N_3101,In_1776,In_1280);
nor U3102 (N_3102,In_2202,In_1410);
and U3103 (N_3103,In_1661,In_1155);
or U3104 (N_3104,In_655,In_2038);
nand U3105 (N_3105,In_2362,In_152);
nor U3106 (N_3106,In_1390,In_2071);
nor U3107 (N_3107,In_2044,In_2053);
or U3108 (N_3108,In_980,In_2447);
nor U3109 (N_3109,In_356,In_783);
and U3110 (N_3110,In_103,In_1684);
or U3111 (N_3111,In_2361,In_1527);
nand U3112 (N_3112,In_859,In_1813);
and U3113 (N_3113,In_2499,In_87);
nand U3114 (N_3114,In_607,In_1102);
xnor U3115 (N_3115,In_423,In_2145);
nor U3116 (N_3116,In_1407,In_2013);
or U3117 (N_3117,In_1666,In_1199);
nand U3118 (N_3118,In_271,In_215);
nor U3119 (N_3119,In_2218,In_1221);
and U3120 (N_3120,In_1287,In_109);
nand U3121 (N_3121,In_1113,In_1055);
xor U3122 (N_3122,In_2406,In_545);
xnor U3123 (N_3123,In_1235,In_982);
nor U3124 (N_3124,In_2310,In_2122);
and U3125 (N_3125,In_1810,In_1145);
and U3126 (N_3126,In_792,In_141);
nor U3127 (N_3127,In_1338,In_624);
nand U3128 (N_3128,In_2345,In_1416);
and U3129 (N_3129,In_622,In_2474);
and U3130 (N_3130,In_1169,In_1100);
nand U3131 (N_3131,In_1728,In_272);
and U3132 (N_3132,In_648,In_1891);
nand U3133 (N_3133,In_775,In_864);
xor U3134 (N_3134,In_259,In_889);
nor U3135 (N_3135,In_407,In_1456);
nor U3136 (N_3136,In_896,In_1412);
nand U3137 (N_3137,In_1619,In_1883);
nor U3138 (N_3138,In_1431,In_1467);
xnor U3139 (N_3139,In_992,In_224);
xnor U3140 (N_3140,In_889,In_1811);
nand U3141 (N_3141,In_1699,In_1133);
nor U3142 (N_3142,In_628,In_755);
xnor U3143 (N_3143,In_1171,In_1884);
nand U3144 (N_3144,In_77,In_1772);
and U3145 (N_3145,In_1752,In_263);
nand U3146 (N_3146,In_1221,In_1058);
xor U3147 (N_3147,In_1644,In_1187);
nand U3148 (N_3148,In_1243,In_2401);
nor U3149 (N_3149,In_528,In_1131);
nand U3150 (N_3150,In_2158,In_1189);
and U3151 (N_3151,In_2217,In_132);
nand U3152 (N_3152,In_1318,In_535);
or U3153 (N_3153,In_2399,In_2217);
nor U3154 (N_3154,In_1449,In_2377);
nor U3155 (N_3155,In_197,In_931);
or U3156 (N_3156,In_617,In_155);
and U3157 (N_3157,In_907,In_1993);
nand U3158 (N_3158,In_1003,In_168);
xor U3159 (N_3159,In_191,In_1026);
and U3160 (N_3160,In_1876,In_1796);
nand U3161 (N_3161,In_630,In_1046);
xor U3162 (N_3162,In_1541,In_444);
nor U3163 (N_3163,In_264,In_140);
nor U3164 (N_3164,In_2217,In_2229);
nor U3165 (N_3165,In_272,In_1867);
and U3166 (N_3166,In_1175,In_1185);
xnor U3167 (N_3167,In_2482,In_810);
or U3168 (N_3168,In_1158,In_710);
nand U3169 (N_3169,In_1707,In_1771);
xor U3170 (N_3170,In_173,In_2389);
xor U3171 (N_3171,In_768,In_866);
and U3172 (N_3172,In_1404,In_916);
nor U3173 (N_3173,In_2028,In_1672);
or U3174 (N_3174,In_563,In_1781);
xor U3175 (N_3175,In_238,In_311);
and U3176 (N_3176,In_211,In_154);
nand U3177 (N_3177,In_1544,In_1825);
xnor U3178 (N_3178,In_2043,In_1140);
nand U3179 (N_3179,In_1192,In_738);
nand U3180 (N_3180,In_1636,In_939);
and U3181 (N_3181,In_1966,In_1916);
or U3182 (N_3182,In_1187,In_490);
nand U3183 (N_3183,In_613,In_953);
nor U3184 (N_3184,In_516,In_2183);
nor U3185 (N_3185,In_2047,In_1108);
or U3186 (N_3186,In_1191,In_251);
and U3187 (N_3187,In_2342,In_610);
nand U3188 (N_3188,In_992,In_810);
nand U3189 (N_3189,In_935,In_2433);
nand U3190 (N_3190,In_1511,In_1703);
and U3191 (N_3191,In_1639,In_1619);
nor U3192 (N_3192,In_2390,In_1341);
nor U3193 (N_3193,In_1950,In_1285);
or U3194 (N_3194,In_857,In_2290);
and U3195 (N_3195,In_542,In_66);
xor U3196 (N_3196,In_1421,In_493);
or U3197 (N_3197,In_2399,In_1999);
and U3198 (N_3198,In_548,In_676);
nor U3199 (N_3199,In_203,In_659);
nand U3200 (N_3200,In_630,In_964);
xnor U3201 (N_3201,In_2089,In_1736);
and U3202 (N_3202,In_1905,In_1553);
xor U3203 (N_3203,In_1293,In_1475);
xor U3204 (N_3204,In_2429,In_114);
and U3205 (N_3205,In_1679,In_691);
or U3206 (N_3206,In_2186,In_2137);
nor U3207 (N_3207,In_2104,In_2042);
xnor U3208 (N_3208,In_1231,In_2441);
and U3209 (N_3209,In_1287,In_1172);
nor U3210 (N_3210,In_332,In_1455);
and U3211 (N_3211,In_692,In_1824);
or U3212 (N_3212,In_2205,In_145);
and U3213 (N_3213,In_663,In_1954);
or U3214 (N_3214,In_702,In_344);
and U3215 (N_3215,In_841,In_1874);
or U3216 (N_3216,In_70,In_462);
nand U3217 (N_3217,In_41,In_1394);
nand U3218 (N_3218,In_916,In_1689);
or U3219 (N_3219,In_516,In_506);
nand U3220 (N_3220,In_298,In_1729);
nor U3221 (N_3221,In_2019,In_635);
or U3222 (N_3222,In_435,In_393);
and U3223 (N_3223,In_634,In_2275);
nand U3224 (N_3224,In_1691,In_1466);
nor U3225 (N_3225,In_247,In_595);
xor U3226 (N_3226,In_1039,In_2322);
nor U3227 (N_3227,In_1975,In_2111);
nor U3228 (N_3228,In_530,In_2441);
nor U3229 (N_3229,In_1868,In_1147);
nand U3230 (N_3230,In_803,In_457);
or U3231 (N_3231,In_1374,In_1114);
nor U3232 (N_3232,In_1621,In_2013);
or U3233 (N_3233,In_1464,In_1140);
xor U3234 (N_3234,In_1493,In_1229);
nor U3235 (N_3235,In_1482,In_1159);
or U3236 (N_3236,In_1574,In_2271);
or U3237 (N_3237,In_591,In_1131);
xor U3238 (N_3238,In_1768,In_2238);
nor U3239 (N_3239,In_2365,In_634);
or U3240 (N_3240,In_644,In_1124);
or U3241 (N_3241,In_2450,In_823);
and U3242 (N_3242,In_1391,In_2268);
and U3243 (N_3243,In_263,In_1536);
and U3244 (N_3244,In_1844,In_187);
nand U3245 (N_3245,In_2324,In_1010);
nand U3246 (N_3246,In_969,In_487);
and U3247 (N_3247,In_770,In_785);
nand U3248 (N_3248,In_1311,In_1933);
nand U3249 (N_3249,In_942,In_982);
nor U3250 (N_3250,In_1281,In_248);
or U3251 (N_3251,In_269,In_868);
xnor U3252 (N_3252,In_1431,In_1411);
nand U3253 (N_3253,In_2037,In_194);
xnor U3254 (N_3254,In_22,In_84);
or U3255 (N_3255,In_1195,In_92);
or U3256 (N_3256,In_2075,In_1260);
or U3257 (N_3257,In_1158,In_1593);
nor U3258 (N_3258,In_1511,In_1870);
nor U3259 (N_3259,In_1596,In_2180);
nor U3260 (N_3260,In_1669,In_838);
or U3261 (N_3261,In_1041,In_710);
nand U3262 (N_3262,In_2480,In_2245);
and U3263 (N_3263,In_210,In_2241);
nand U3264 (N_3264,In_1834,In_1754);
or U3265 (N_3265,In_2132,In_1207);
nor U3266 (N_3266,In_463,In_938);
nand U3267 (N_3267,In_2247,In_1582);
xnor U3268 (N_3268,In_449,In_113);
and U3269 (N_3269,In_567,In_828);
or U3270 (N_3270,In_224,In_2437);
nor U3271 (N_3271,In_820,In_1911);
xor U3272 (N_3272,In_2458,In_1446);
xor U3273 (N_3273,In_2009,In_658);
and U3274 (N_3274,In_1490,In_687);
nand U3275 (N_3275,In_2121,In_1328);
or U3276 (N_3276,In_1722,In_2193);
nand U3277 (N_3277,In_2350,In_2419);
and U3278 (N_3278,In_830,In_2002);
or U3279 (N_3279,In_284,In_1346);
nand U3280 (N_3280,In_1380,In_1402);
nor U3281 (N_3281,In_1558,In_1489);
nand U3282 (N_3282,In_161,In_1235);
xnor U3283 (N_3283,In_2487,In_1125);
nand U3284 (N_3284,In_699,In_915);
and U3285 (N_3285,In_1980,In_937);
xnor U3286 (N_3286,In_266,In_996);
or U3287 (N_3287,In_2011,In_2223);
or U3288 (N_3288,In_717,In_2304);
and U3289 (N_3289,In_2033,In_1357);
or U3290 (N_3290,In_641,In_1474);
nor U3291 (N_3291,In_751,In_586);
or U3292 (N_3292,In_2158,In_831);
xor U3293 (N_3293,In_1723,In_1832);
nor U3294 (N_3294,In_1824,In_2300);
or U3295 (N_3295,In_2461,In_1790);
nand U3296 (N_3296,In_2104,In_1338);
and U3297 (N_3297,In_1728,In_230);
and U3298 (N_3298,In_1263,In_1581);
xor U3299 (N_3299,In_2310,In_1169);
nor U3300 (N_3300,In_2073,In_994);
xnor U3301 (N_3301,In_1909,In_1793);
and U3302 (N_3302,In_1042,In_1871);
nor U3303 (N_3303,In_1714,In_394);
and U3304 (N_3304,In_1403,In_22);
and U3305 (N_3305,In_1687,In_824);
and U3306 (N_3306,In_1703,In_1245);
or U3307 (N_3307,In_576,In_1825);
xnor U3308 (N_3308,In_1582,In_1850);
and U3309 (N_3309,In_379,In_512);
nand U3310 (N_3310,In_648,In_534);
nand U3311 (N_3311,In_467,In_1361);
and U3312 (N_3312,In_182,In_908);
or U3313 (N_3313,In_1627,In_1596);
and U3314 (N_3314,In_2328,In_2453);
nand U3315 (N_3315,In_1550,In_799);
and U3316 (N_3316,In_1472,In_1040);
nor U3317 (N_3317,In_1431,In_2318);
nor U3318 (N_3318,In_2010,In_1738);
nand U3319 (N_3319,In_2189,In_1361);
and U3320 (N_3320,In_1749,In_914);
and U3321 (N_3321,In_2461,In_1489);
xor U3322 (N_3322,In_765,In_2412);
nor U3323 (N_3323,In_2452,In_2097);
or U3324 (N_3324,In_1723,In_342);
nor U3325 (N_3325,In_1002,In_768);
nor U3326 (N_3326,In_1289,In_562);
nor U3327 (N_3327,In_1107,In_1047);
and U3328 (N_3328,In_319,In_650);
nor U3329 (N_3329,In_741,In_303);
nor U3330 (N_3330,In_185,In_1703);
xnor U3331 (N_3331,In_2232,In_485);
xor U3332 (N_3332,In_308,In_171);
and U3333 (N_3333,In_1650,In_878);
nand U3334 (N_3334,In_143,In_1156);
or U3335 (N_3335,In_945,In_2171);
or U3336 (N_3336,In_1873,In_415);
nand U3337 (N_3337,In_721,In_1542);
xnor U3338 (N_3338,In_2096,In_2474);
xor U3339 (N_3339,In_1844,In_1718);
nand U3340 (N_3340,In_1584,In_2122);
and U3341 (N_3341,In_2100,In_894);
nor U3342 (N_3342,In_1774,In_1473);
nand U3343 (N_3343,In_1232,In_78);
nor U3344 (N_3344,In_2485,In_1267);
nand U3345 (N_3345,In_268,In_2143);
nand U3346 (N_3346,In_284,In_100);
nor U3347 (N_3347,In_1868,In_1789);
and U3348 (N_3348,In_1619,In_1485);
nor U3349 (N_3349,In_2225,In_2237);
nand U3350 (N_3350,In_2087,In_340);
or U3351 (N_3351,In_2393,In_2246);
and U3352 (N_3352,In_1343,In_89);
and U3353 (N_3353,In_380,In_410);
nand U3354 (N_3354,In_1175,In_2123);
or U3355 (N_3355,In_1302,In_1663);
nor U3356 (N_3356,In_1724,In_1691);
and U3357 (N_3357,In_1551,In_1422);
or U3358 (N_3358,In_1535,In_143);
and U3359 (N_3359,In_384,In_776);
and U3360 (N_3360,In_87,In_2225);
and U3361 (N_3361,In_856,In_1829);
and U3362 (N_3362,In_1541,In_614);
nor U3363 (N_3363,In_341,In_771);
nand U3364 (N_3364,In_21,In_296);
nand U3365 (N_3365,In_1817,In_503);
and U3366 (N_3366,In_2474,In_1396);
and U3367 (N_3367,In_1623,In_771);
xor U3368 (N_3368,In_925,In_1222);
or U3369 (N_3369,In_2482,In_593);
nand U3370 (N_3370,In_85,In_1797);
xnor U3371 (N_3371,In_2165,In_1228);
nand U3372 (N_3372,In_2411,In_615);
nand U3373 (N_3373,In_1794,In_1981);
nor U3374 (N_3374,In_27,In_2231);
xnor U3375 (N_3375,In_1451,In_1281);
and U3376 (N_3376,In_1564,In_972);
and U3377 (N_3377,In_1460,In_1696);
nand U3378 (N_3378,In_780,In_743);
xor U3379 (N_3379,In_1441,In_3);
and U3380 (N_3380,In_2133,In_1630);
nand U3381 (N_3381,In_1912,In_945);
nand U3382 (N_3382,In_1447,In_2417);
xor U3383 (N_3383,In_2011,In_1623);
xnor U3384 (N_3384,In_2044,In_776);
nor U3385 (N_3385,In_1271,In_317);
or U3386 (N_3386,In_36,In_209);
nand U3387 (N_3387,In_180,In_1133);
nand U3388 (N_3388,In_1577,In_2331);
nor U3389 (N_3389,In_1898,In_2485);
xnor U3390 (N_3390,In_417,In_959);
nand U3391 (N_3391,In_497,In_1780);
nand U3392 (N_3392,In_499,In_2469);
nand U3393 (N_3393,In_1402,In_678);
or U3394 (N_3394,In_345,In_1590);
or U3395 (N_3395,In_777,In_755);
nor U3396 (N_3396,In_1745,In_1325);
or U3397 (N_3397,In_715,In_2041);
or U3398 (N_3398,In_1238,In_1662);
xnor U3399 (N_3399,In_1864,In_1726);
xor U3400 (N_3400,In_1279,In_2424);
nor U3401 (N_3401,In_1600,In_1141);
nor U3402 (N_3402,In_1603,In_2351);
xor U3403 (N_3403,In_1746,In_1616);
nand U3404 (N_3404,In_1869,In_30);
nand U3405 (N_3405,In_1153,In_688);
or U3406 (N_3406,In_1772,In_2414);
or U3407 (N_3407,In_1404,In_338);
and U3408 (N_3408,In_145,In_1964);
nand U3409 (N_3409,In_1378,In_515);
nand U3410 (N_3410,In_1504,In_739);
nor U3411 (N_3411,In_860,In_421);
and U3412 (N_3412,In_719,In_2168);
or U3413 (N_3413,In_211,In_403);
xor U3414 (N_3414,In_829,In_1480);
nand U3415 (N_3415,In_2209,In_39);
or U3416 (N_3416,In_1268,In_838);
nand U3417 (N_3417,In_819,In_509);
or U3418 (N_3418,In_2172,In_1773);
nand U3419 (N_3419,In_713,In_2054);
nor U3420 (N_3420,In_1245,In_294);
nand U3421 (N_3421,In_1942,In_1510);
and U3422 (N_3422,In_953,In_477);
or U3423 (N_3423,In_443,In_2216);
xnor U3424 (N_3424,In_2362,In_368);
or U3425 (N_3425,In_1308,In_1575);
nor U3426 (N_3426,In_304,In_892);
and U3427 (N_3427,In_1875,In_214);
and U3428 (N_3428,In_349,In_931);
or U3429 (N_3429,In_312,In_494);
xnor U3430 (N_3430,In_2382,In_2215);
or U3431 (N_3431,In_2030,In_2186);
nand U3432 (N_3432,In_1339,In_714);
or U3433 (N_3433,In_695,In_2158);
xor U3434 (N_3434,In_658,In_914);
and U3435 (N_3435,In_778,In_2446);
nand U3436 (N_3436,In_1160,In_634);
nand U3437 (N_3437,In_2347,In_234);
xnor U3438 (N_3438,In_1943,In_2149);
and U3439 (N_3439,In_2024,In_582);
or U3440 (N_3440,In_1151,In_1880);
or U3441 (N_3441,In_294,In_2229);
and U3442 (N_3442,In_547,In_714);
xor U3443 (N_3443,In_1096,In_1606);
nor U3444 (N_3444,In_2065,In_641);
or U3445 (N_3445,In_1849,In_347);
xnor U3446 (N_3446,In_2181,In_2022);
or U3447 (N_3447,In_1529,In_975);
nor U3448 (N_3448,In_954,In_1140);
and U3449 (N_3449,In_277,In_453);
nor U3450 (N_3450,In_1755,In_1180);
nor U3451 (N_3451,In_1295,In_2263);
or U3452 (N_3452,In_960,In_1806);
nand U3453 (N_3453,In_727,In_110);
nand U3454 (N_3454,In_811,In_1190);
nand U3455 (N_3455,In_693,In_2283);
or U3456 (N_3456,In_1893,In_1634);
nor U3457 (N_3457,In_1706,In_2135);
and U3458 (N_3458,In_1187,In_486);
nor U3459 (N_3459,In_947,In_2035);
nand U3460 (N_3460,In_155,In_2148);
nand U3461 (N_3461,In_2429,In_1691);
xnor U3462 (N_3462,In_1308,In_1585);
nand U3463 (N_3463,In_547,In_617);
nor U3464 (N_3464,In_1599,In_1352);
nor U3465 (N_3465,In_1778,In_1201);
nor U3466 (N_3466,In_739,In_2441);
nor U3467 (N_3467,In_1645,In_2381);
and U3468 (N_3468,In_1583,In_756);
nor U3469 (N_3469,In_1664,In_861);
nor U3470 (N_3470,In_1336,In_1366);
or U3471 (N_3471,In_3,In_2279);
nor U3472 (N_3472,In_1941,In_533);
or U3473 (N_3473,In_2269,In_1677);
xor U3474 (N_3474,In_2076,In_2027);
nor U3475 (N_3475,In_996,In_1264);
or U3476 (N_3476,In_2062,In_404);
nor U3477 (N_3477,In_1134,In_2395);
and U3478 (N_3478,In_893,In_279);
nor U3479 (N_3479,In_662,In_534);
nor U3480 (N_3480,In_1857,In_327);
xor U3481 (N_3481,In_2215,In_1920);
and U3482 (N_3482,In_2177,In_1151);
nand U3483 (N_3483,In_1061,In_625);
and U3484 (N_3484,In_167,In_59);
xnor U3485 (N_3485,In_2334,In_1546);
and U3486 (N_3486,In_1465,In_2140);
nand U3487 (N_3487,In_1746,In_1892);
nor U3488 (N_3488,In_1469,In_1375);
xnor U3489 (N_3489,In_884,In_1171);
nand U3490 (N_3490,In_483,In_1446);
nor U3491 (N_3491,In_1920,In_2220);
or U3492 (N_3492,In_2310,In_1748);
or U3493 (N_3493,In_2080,In_507);
nand U3494 (N_3494,In_1202,In_837);
and U3495 (N_3495,In_1955,In_547);
nand U3496 (N_3496,In_1216,In_963);
nand U3497 (N_3497,In_25,In_2176);
or U3498 (N_3498,In_1348,In_410);
nor U3499 (N_3499,In_402,In_21);
nand U3500 (N_3500,In_256,In_525);
and U3501 (N_3501,In_917,In_1684);
xor U3502 (N_3502,In_1773,In_1086);
or U3503 (N_3503,In_1935,In_117);
or U3504 (N_3504,In_1222,In_1155);
or U3505 (N_3505,In_462,In_1721);
and U3506 (N_3506,In_1104,In_375);
or U3507 (N_3507,In_1333,In_1449);
or U3508 (N_3508,In_1140,In_2461);
or U3509 (N_3509,In_84,In_102);
nand U3510 (N_3510,In_24,In_1945);
nor U3511 (N_3511,In_2015,In_191);
and U3512 (N_3512,In_1546,In_2439);
xnor U3513 (N_3513,In_1081,In_404);
nor U3514 (N_3514,In_81,In_106);
nand U3515 (N_3515,In_1803,In_489);
and U3516 (N_3516,In_829,In_245);
or U3517 (N_3517,In_522,In_529);
nand U3518 (N_3518,In_614,In_622);
xor U3519 (N_3519,In_642,In_2415);
xor U3520 (N_3520,In_2197,In_385);
or U3521 (N_3521,In_1795,In_2273);
and U3522 (N_3522,In_420,In_28);
nor U3523 (N_3523,In_158,In_1310);
nor U3524 (N_3524,In_1265,In_2000);
and U3525 (N_3525,In_2150,In_2199);
xnor U3526 (N_3526,In_1096,In_1477);
nor U3527 (N_3527,In_2443,In_1419);
xor U3528 (N_3528,In_594,In_1628);
and U3529 (N_3529,In_1330,In_635);
or U3530 (N_3530,In_273,In_1567);
xnor U3531 (N_3531,In_784,In_2486);
or U3532 (N_3532,In_286,In_553);
or U3533 (N_3533,In_1829,In_796);
xnor U3534 (N_3534,In_1276,In_2096);
or U3535 (N_3535,In_330,In_1094);
nor U3536 (N_3536,In_450,In_303);
nand U3537 (N_3537,In_1422,In_1227);
xnor U3538 (N_3538,In_1339,In_1003);
and U3539 (N_3539,In_1575,In_568);
nor U3540 (N_3540,In_1844,In_718);
and U3541 (N_3541,In_1000,In_1377);
nor U3542 (N_3542,In_1034,In_468);
nand U3543 (N_3543,In_2359,In_1714);
xnor U3544 (N_3544,In_1705,In_1907);
nor U3545 (N_3545,In_1654,In_997);
nand U3546 (N_3546,In_758,In_916);
or U3547 (N_3547,In_1681,In_1102);
nor U3548 (N_3548,In_9,In_1063);
or U3549 (N_3549,In_608,In_462);
or U3550 (N_3550,In_1952,In_2234);
nand U3551 (N_3551,In_1790,In_1599);
nor U3552 (N_3552,In_311,In_2365);
or U3553 (N_3553,In_1915,In_86);
or U3554 (N_3554,In_2365,In_132);
and U3555 (N_3555,In_1753,In_1555);
xnor U3556 (N_3556,In_1464,In_1669);
and U3557 (N_3557,In_75,In_167);
nand U3558 (N_3558,In_711,In_1450);
xor U3559 (N_3559,In_839,In_1143);
nand U3560 (N_3560,In_1013,In_1925);
and U3561 (N_3561,In_2417,In_175);
nor U3562 (N_3562,In_1729,In_1385);
nand U3563 (N_3563,In_1364,In_2254);
nand U3564 (N_3564,In_1572,In_1372);
or U3565 (N_3565,In_2050,In_2203);
or U3566 (N_3566,In_379,In_191);
and U3567 (N_3567,In_1518,In_855);
and U3568 (N_3568,In_1041,In_674);
and U3569 (N_3569,In_892,In_718);
and U3570 (N_3570,In_1383,In_280);
and U3571 (N_3571,In_2114,In_1490);
nor U3572 (N_3572,In_832,In_352);
nor U3573 (N_3573,In_1724,In_1283);
and U3574 (N_3574,In_1447,In_1422);
xor U3575 (N_3575,In_721,In_910);
or U3576 (N_3576,In_1868,In_1758);
nand U3577 (N_3577,In_1985,In_870);
xnor U3578 (N_3578,In_367,In_1044);
or U3579 (N_3579,In_1528,In_1261);
nor U3580 (N_3580,In_2122,In_465);
or U3581 (N_3581,In_335,In_682);
nor U3582 (N_3582,In_60,In_1630);
and U3583 (N_3583,In_50,In_1182);
xnor U3584 (N_3584,In_1166,In_275);
xor U3585 (N_3585,In_1302,In_1257);
or U3586 (N_3586,In_1141,In_1642);
nor U3587 (N_3587,In_2132,In_37);
xnor U3588 (N_3588,In_372,In_1543);
xnor U3589 (N_3589,In_2133,In_236);
and U3590 (N_3590,In_1561,In_1225);
nand U3591 (N_3591,In_989,In_2361);
and U3592 (N_3592,In_675,In_1559);
xnor U3593 (N_3593,In_313,In_2472);
nor U3594 (N_3594,In_942,In_999);
and U3595 (N_3595,In_616,In_2419);
or U3596 (N_3596,In_1326,In_609);
or U3597 (N_3597,In_1958,In_206);
xnor U3598 (N_3598,In_1934,In_868);
nand U3599 (N_3599,In_1321,In_207);
xor U3600 (N_3600,In_904,In_1493);
xnor U3601 (N_3601,In_1903,In_1472);
nor U3602 (N_3602,In_1304,In_255);
and U3603 (N_3603,In_877,In_450);
xnor U3604 (N_3604,In_1942,In_1695);
xnor U3605 (N_3605,In_1197,In_1968);
or U3606 (N_3606,In_1108,In_1154);
and U3607 (N_3607,In_274,In_1173);
and U3608 (N_3608,In_366,In_1648);
nand U3609 (N_3609,In_1900,In_426);
or U3610 (N_3610,In_2246,In_1113);
and U3611 (N_3611,In_1144,In_14);
or U3612 (N_3612,In_1627,In_1162);
and U3613 (N_3613,In_909,In_1938);
nand U3614 (N_3614,In_329,In_341);
or U3615 (N_3615,In_620,In_2399);
nor U3616 (N_3616,In_2003,In_383);
xor U3617 (N_3617,In_1791,In_939);
xnor U3618 (N_3618,In_2072,In_1933);
nor U3619 (N_3619,In_1234,In_448);
or U3620 (N_3620,In_666,In_14);
nand U3621 (N_3621,In_1821,In_2236);
xor U3622 (N_3622,In_116,In_1756);
xnor U3623 (N_3623,In_1948,In_19);
xnor U3624 (N_3624,In_2470,In_2451);
xnor U3625 (N_3625,In_865,In_887);
or U3626 (N_3626,In_1211,In_1630);
nor U3627 (N_3627,In_2118,In_1980);
nand U3628 (N_3628,In_2086,In_689);
or U3629 (N_3629,In_2406,In_402);
and U3630 (N_3630,In_1628,In_1429);
or U3631 (N_3631,In_1233,In_1826);
and U3632 (N_3632,In_1818,In_303);
xnor U3633 (N_3633,In_588,In_986);
and U3634 (N_3634,In_1853,In_906);
nor U3635 (N_3635,In_1927,In_148);
xor U3636 (N_3636,In_846,In_465);
nor U3637 (N_3637,In_1460,In_1062);
or U3638 (N_3638,In_1683,In_2157);
nor U3639 (N_3639,In_622,In_1577);
nand U3640 (N_3640,In_2479,In_57);
or U3641 (N_3641,In_1777,In_66);
and U3642 (N_3642,In_862,In_1673);
nand U3643 (N_3643,In_1946,In_408);
nor U3644 (N_3644,In_1027,In_2203);
nor U3645 (N_3645,In_240,In_2141);
and U3646 (N_3646,In_526,In_2309);
or U3647 (N_3647,In_1503,In_1983);
nand U3648 (N_3648,In_829,In_2485);
nand U3649 (N_3649,In_22,In_1254);
or U3650 (N_3650,In_622,In_148);
nor U3651 (N_3651,In_1364,In_814);
xor U3652 (N_3652,In_1806,In_1720);
or U3653 (N_3653,In_1608,In_1138);
or U3654 (N_3654,In_207,In_805);
nand U3655 (N_3655,In_1276,In_849);
nand U3656 (N_3656,In_2443,In_2294);
xnor U3657 (N_3657,In_595,In_1305);
and U3658 (N_3658,In_886,In_429);
xor U3659 (N_3659,In_2257,In_2256);
or U3660 (N_3660,In_2318,In_855);
xnor U3661 (N_3661,In_1135,In_1625);
nand U3662 (N_3662,In_422,In_1681);
xor U3663 (N_3663,In_410,In_2097);
nand U3664 (N_3664,In_2229,In_23);
or U3665 (N_3665,In_1806,In_2184);
or U3666 (N_3666,In_865,In_475);
xor U3667 (N_3667,In_59,In_2004);
and U3668 (N_3668,In_248,In_1712);
xor U3669 (N_3669,In_1911,In_1641);
nor U3670 (N_3670,In_668,In_1741);
nor U3671 (N_3671,In_2478,In_2351);
or U3672 (N_3672,In_2214,In_1685);
xor U3673 (N_3673,In_576,In_1514);
or U3674 (N_3674,In_1547,In_2279);
xor U3675 (N_3675,In_923,In_1306);
nand U3676 (N_3676,In_1524,In_1509);
and U3677 (N_3677,In_2210,In_1941);
nor U3678 (N_3678,In_334,In_722);
or U3679 (N_3679,In_96,In_2485);
nor U3680 (N_3680,In_1135,In_287);
and U3681 (N_3681,In_2078,In_241);
nand U3682 (N_3682,In_1932,In_304);
xor U3683 (N_3683,In_1861,In_1822);
or U3684 (N_3684,In_2214,In_1236);
or U3685 (N_3685,In_163,In_2016);
xor U3686 (N_3686,In_341,In_2385);
nand U3687 (N_3687,In_2190,In_1085);
nand U3688 (N_3688,In_827,In_2497);
or U3689 (N_3689,In_1168,In_451);
and U3690 (N_3690,In_993,In_1082);
nor U3691 (N_3691,In_1561,In_1728);
or U3692 (N_3692,In_2171,In_1055);
and U3693 (N_3693,In_564,In_276);
and U3694 (N_3694,In_568,In_1640);
xnor U3695 (N_3695,In_1563,In_132);
or U3696 (N_3696,In_582,In_2159);
nand U3697 (N_3697,In_2110,In_1443);
and U3698 (N_3698,In_1663,In_1267);
and U3699 (N_3699,In_181,In_763);
nor U3700 (N_3700,In_1275,In_569);
or U3701 (N_3701,In_966,In_225);
nor U3702 (N_3702,In_1341,In_538);
or U3703 (N_3703,In_17,In_1297);
and U3704 (N_3704,In_696,In_712);
nor U3705 (N_3705,In_96,In_238);
xor U3706 (N_3706,In_435,In_362);
and U3707 (N_3707,In_1315,In_2204);
xor U3708 (N_3708,In_585,In_2261);
xnor U3709 (N_3709,In_368,In_868);
or U3710 (N_3710,In_595,In_1600);
nand U3711 (N_3711,In_2279,In_2491);
nand U3712 (N_3712,In_274,In_2485);
xnor U3713 (N_3713,In_2404,In_1513);
nand U3714 (N_3714,In_303,In_2033);
nor U3715 (N_3715,In_1624,In_1007);
or U3716 (N_3716,In_247,In_1015);
and U3717 (N_3717,In_1562,In_1531);
and U3718 (N_3718,In_147,In_661);
xor U3719 (N_3719,In_173,In_2322);
or U3720 (N_3720,In_1592,In_1738);
nand U3721 (N_3721,In_1811,In_2437);
nor U3722 (N_3722,In_763,In_1000);
xnor U3723 (N_3723,In_2349,In_2241);
nand U3724 (N_3724,In_1241,In_1494);
xnor U3725 (N_3725,In_174,In_1251);
or U3726 (N_3726,In_1185,In_879);
nand U3727 (N_3727,In_2114,In_270);
nand U3728 (N_3728,In_970,In_1874);
xnor U3729 (N_3729,In_1576,In_2284);
xnor U3730 (N_3730,In_541,In_1013);
or U3731 (N_3731,In_1175,In_886);
xnor U3732 (N_3732,In_1071,In_100);
or U3733 (N_3733,In_1436,In_1189);
or U3734 (N_3734,In_381,In_1408);
xnor U3735 (N_3735,In_2166,In_1261);
nand U3736 (N_3736,In_952,In_2032);
and U3737 (N_3737,In_1856,In_1973);
nand U3738 (N_3738,In_1605,In_1969);
xnor U3739 (N_3739,In_802,In_470);
and U3740 (N_3740,In_2134,In_2366);
and U3741 (N_3741,In_1164,In_1886);
nor U3742 (N_3742,In_1180,In_1058);
nand U3743 (N_3743,In_580,In_1953);
xor U3744 (N_3744,In_932,In_1103);
or U3745 (N_3745,In_599,In_1323);
xor U3746 (N_3746,In_1627,In_1333);
xor U3747 (N_3747,In_1178,In_2269);
nand U3748 (N_3748,In_2192,In_1135);
and U3749 (N_3749,In_2069,In_1199);
nor U3750 (N_3750,In_293,In_1261);
nor U3751 (N_3751,In_1209,In_2095);
or U3752 (N_3752,In_168,In_124);
or U3753 (N_3753,In_2321,In_1219);
xnor U3754 (N_3754,In_1715,In_71);
and U3755 (N_3755,In_2377,In_2476);
xor U3756 (N_3756,In_921,In_845);
and U3757 (N_3757,In_363,In_517);
nor U3758 (N_3758,In_9,In_137);
xor U3759 (N_3759,In_1836,In_2415);
or U3760 (N_3760,In_1906,In_456);
xor U3761 (N_3761,In_1663,In_1967);
nand U3762 (N_3762,In_1440,In_1086);
and U3763 (N_3763,In_763,In_2052);
and U3764 (N_3764,In_1023,In_1897);
xnor U3765 (N_3765,In_195,In_1492);
nor U3766 (N_3766,In_938,In_766);
or U3767 (N_3767,In_2391,In_519);
xor U3768 (N_3768,In_2369,In_1387);
and U3769 (N_3769,In_2130,In_2352);
xor U3770 (N_3770,In_2241,In_2283);
or U3771 (N_3771,In_860,In_2026);
and U3772 (N_3772,In_1188,In_804);
nor U3773 (N_3773,In_1485,In_1978);
or U3774 (N_3774,In_2092,In_680);
xnor U3775 (N_3775,In_802,In_513);
or U3776 (N_3776,In_1597,In_822);
or U3777 (N_3777,In_856,In_2247);
xnor U3778 (N_3778,In_1737,In_2367);
nand U3779 (N_3779,In_1817,In_270);
or U3780 (N_3780,In_2020,In_81);
nand U3781 (N_3781,In_2180,In_2440);
or U3782 (N_3782,In_413,In_1043);
nor U3783 (N_3783,In_2232,In_363);
or U3784 (N_3784,In_1789,In_1338);
nand U3785 (N_3785,In_4,In_404);
nand U3786 (N_3786,In_587,In_396);
xor U3787 (N_3787,In_1989,In_1930);
and U3788 (N_3788,In_2433,In_110);
or U3789 (N_3789,In_847,In_2386);
and U3790 (N_3790,In_1824,In_413);
and U3791 (N_3791,In_1295,In_1415);
or U3792 (N_3792,In_2251,In_693);
or U3793 (N_3793,In_1590,In_769);
nor U3794 (N_3794,In_836,In_1591);
nor U3795 (N_3795,In_421,In_1702);
or U3796 (N_3796,In_1462,In_1764);
nor U3797 (N_3797,In_991,In_2157);
nor U3798 (N_3798,In_1457,In_2195);
and U3799 (N_3799,In_1885,In_998);
nand U3800 (N_3800,In_2146,In_687);
or U3801 (N_3801,In_848,In_283);
and U3802 (N_3802,In_1491,In_972);
and U3803 (N_3803,In_2114,In_1415);
or U3804 (N_3804,In_2034,In_2125);
nor U3805 (N_3805,In_705,In_1038);
nand U3806 (N_3806,In_1502,In_2277);
or U3807 (N_3807,In_2423,In_1973);
and U3808 (N_3808,In_1930,In_1126);
xnor U3809 (N_3809,In_490,In_2247);
nand U3810 (N_3810,In_1535,In_552);
xnor U3811 (N_3811,In_1732,In_337);
nor U3812 (N_3812,In_1126,In_1700);
nor U3813 (N_3813,In_1139,In_1711);
nand U3814 (N_3814,In_1161,In_1116);
nor U3815 (N_3815,In_1005,In_2261);
nor U3816 (N_3816,In_477,In_1176);
nor U3817 (N_3817,In_730,In_2318);
nor U3818 (N_3818,In_1978,In_1896);
xnor U3819 (N_3819,In_474,In_1561);
or U3820 (N_3820,In_920,In_75);
nand U3821 (N_3821,In_498,In_494);
and U3822 (N_3822,In_1084,In_1422);
xnor U3823 (N_3823,In_168,In_1556);
and U3824 (N_3824,In_1182,In_1409);
xnor U3825 (N_3825,In_752,In_1104);
nand U3826 (N_3826,In_549,In_111);
nand U3827 (N_3827,In_689,In_558);
xnor U3828 (N_3828,In_1464,In_1565);
nand U3829 (N_3829,In_263,In_1131);
nand U3830 (N_3830,In_63,In_709);
nand U3831 (N_3831,In_1431,In_1109);
or U3832 (N_3832,In_1289,In_2206);
and U3833 (N_3833,In_474,In_1500);
nor U3834 (N_3834,In_1955,In_1819);
nor U3835 (N_3835,In_1431,In_446);
nor U3836 (N_3836,In_2420,In_862);
nand U3837 (N_3837,In_271,In_2497);
and U3838 (N_3838,In_68,In_1531);
nor U3839 (N_3839,In_1561,In_772);
nor U3840 (N_3840,In_702,In_1223);
and U3841 (N_3841,In_1613,In_327);
xnor U3842 (N_3842,In_517,In_1358);
nor U3843 (N_3843,In_717,In_358);
and U3844 (N_3844,In_2472,In_967);
or U3845 (N_3845,In_1750,In_1120);
xor U3846 (N_3846,In_896,In_1217);
and U3847 (N_3847,In_479,In_1537);
xor U3848 (N_3848,In_180,In_3);
and U3849 (N_3849,In_2101,In_1560);
or U3850 (N_3850,In_1438,In_1960);
xor U3851 (N_3851,In_1000,In_1988);
xor U3852 (N_3852,In_1548,In_1952);
and U3853 (N_3853,In_1684,In_15);
xnor U3854 (N_3854,In_151,In_263);
nand U3855 (N_3855,In_1620,In_2244);
nand U3856 (N_3856,In_521,In_1162);
xor U3857 (N_3857,In_2212,In_1778);
nand U3858 (N_3858,In_2313,In_1177);
nor U3859 (N_3859,In_1957,In_2415);
nand U3860 (N_3860,In_1442,In_1253);
or U3861 (N_3861,In_2350,In_778);
nand U3862 (N_3862,In_594,In_2378);
nor U3863 (N_3863,In_156,In_1852);
nor U3864 (N_3864,In_1044,In_1760);
or U3865 (N_3865,In_1088,In_2486);
and U3866 (N_3866,In_1210,In_807);
and U3867 (N_3867,In_663,In_1758);
xnor U3868 (N_3868,In_1456,In_1855);
nand U3869 (N_3869,In_2212,In_1232);
and U3870 (N_3870,In_872,In_1200);
or U3871 (N_3871,In_1877,In_134);
or U3872 (N_3872,In_389,In_1431);
nand U3873 (N_3873,In_1137,In_1710);
or U3874 (N_3874,In_1978,In_1394);
and U3875 (N_3875,In_1453,In_1732);
and U3876 (N_3876,In_190,In_2273);
nand U3877 (N_3877,In_2207,In_2452);
nand U3878 (N_3878,In_169,In_1196);
or U3879 (N_3879,In_2459,In_668);
and U3880 (N_3880,In_2455,In_1789);
and U3881 (N_3881,In_2188,In_886);
nand U3882 (N_3882,In_396,In_1388);
nor U3883 (N_3883,In_1976,In_1360);
nand U3884 (N_3884,In_2022,In_1672);
and U3885 (N_3885,In_2188,In_2320);
nand U3886 (N_3886,In_486,In_1165);
xnor U3887 (N_3887,In_1233,In_2365);
nand U3888 (N_3888,In_757,In_427);
and U3889 (N_3889,In_1236,In_1319);
nor U3890 (N_3890,In_643,In_2420);
nand U3891 (N_3891,In_1134,In_1873);
xor U3892 (N_3892,In_1624,In_2421);
nor U3893 (N_3893,In_1719,In_1915);
nand U3894 (N_3894,In_1397,In_1543);
xnor U3895 (N_3895,In_497,In_1580);
xor U3896 (N_3896,In_1899,In_1562);
xor U3897 (N_3897,In_2118,In_2198);
and U3898 (N_3898,In_865,In_192);
or U3899 (N_3899,In_62,In_243);
nand U3900 (N_3900,In_2035,In_2066);
and U3901 (N_3901,In_601,In_1873);
nor U3902 (N_3902,In_965,In_1125);
xor U3903 (N_3903,In_1974,In_45);
and U3904 (N_3904,In_2246,In_916);
or U3905 (N_3905,In_2021,In_2040);
nand U3906 (N_3906,In_1126,In_1262);
nor U3907 (N_3907,In_1101,In_666);
xor U3908 (N_3908,In_1678,In_1285);
nand U3909 (N_3909,In_2006,In_1255);
xor U3910 (N_3910,In_246,In_44);
nand U3911 (N_3911,In_603,In_1691);
or U3912 (N_3912,In_164,In_1789);
nor U3913 (N_3913,In_1132,In_1982);
nand U3914 (N_3914,In_2349,In_1979);
xnor U3915 (N_3915,In_1439,In_1261);
nor U3916 (N_3916,In_2359,In_1272);
nor U3917 (N_3917,In_2362,In_1577);
xnor U3918 (N_3918,In_2079,In_779);
nor U3919 (N_3919,In_51,In_1714);
nor U3920 (N_3920,In_1121,In_173);
xnor U3921 (N_3921,In_2385,In_1702);
nand U3922 (N_3922,In_457,In_2064);
nor U3923 (N_3923,In_1428,In_614);
nor U3924 (N_3924,In_2297,In_210);
nor U3925 (N_3925,In_2076,In_2152);
and U3926 (N_3926,In_205,In_569);
nor U3927 (N_3927,In_2474,In_1390);
nand U3928 (N_3928,In_648,In_241);
and U3929 (N_3929,In_1729,In_1840);
nand U3930 (N_3930,In_1184,In_2353);
and U3931 (N_3931,In_1888,In_661);
or U3932 (N_3932,In_1599,In_1251);
nand U3933 (N_3933,In_1929,In_1780);
and U3934 (N_3934,In_2462,In_1619);
nor U3935 (N_3935,In_1128,In_2219);
or U3936 (N_3936,In_532,In_1395);
or U3937 (N_3937,In_886,In_1494);
nand U3938 (N_3938,In_1077,In_2100);
nand U3939 (N_3939,In_2073,In_1125);
xnor U3940 (N_3940,In_1691,In_2116);
and U3941 (N_3941,In_2178,In_1487);
and U3942 (N_3942,In_27,In_1638);
and U3943 (N_3943,In_2395,In_2036);
nand U3944 (N_3944,In_1763,In_1534);
nor U3945 (N_3945,In_604,In_1072);
or U3946 (N_3946,In_879,In_1134);
nor U3947 (N_3947,In_887,In_1859);
xnor U3948 (N_3948,In_1607,In_365);
nor U3949 (N_3949,In_1730,In_820);
xnor U3950 (N_3950,In_1720,In_983);
nor U3951 (N_3951,In_2308,In_1406);
or U3952 (N_3952,In_464,In_2230);
or U3953 (N_3953,In_2053,In_1402);
or U3954 (N_3954,In_563,In_7);
or U3955 (N_3955,In_1496,In_236);
xnor U3956 (N_3956,In_1409,In_2315);
xnor U3957 (N_3957,In_996,In_1190);
and U3958 (N_3958,In_2338,In_101);
nand U3959 (N_3959,In_1168,In_1493);
or U3960 (N_3960,In_98,In_1839);
and U3961 (N_3961,In_1053,In_1184);
nor U3962 (N_3962,In_375,In_1140);
xor U3963 (N_3963,In_1008,In_430);
or U3964 (N_3964,In_407,In_229);
xor U3965 (N_3965,In_903,In_1590);
xnor U3966 (N_3966,In_1052,In_1173);
xnor U3967 (N_3967,In_1467,In_2208);
nor U3968 (N_3968,In_762,In_1208);
nor U3969 (N_3969,In_1085,In_957);
or U3970 (N_3970,In_1175,In_953);
and U3971 (N_3971,In_660,In_590);
xnor U3972 (N_3972,In_2345,In_1118);
xor U3973 (N_3973,In_2394,In_2357);
xor U3974 (N_3974,In_1406,In_1560);
nand U3975 (N_3975,In_1217,In_86);
or U3976 (N_3976,In_105,In_496);
or U3977 (N_3977,In_2157,In_419);
and U3978 (N_3978,In_261,In_166);
nor U3979 (N_3979,In_1232,In_903);
xor U3980 (N_3980,In_1660,In_661);
nor U3981 (N_3981,In_1707,In_444);
or U3982 (N_3982,In_947,In_2461);
xor U3983 (N_3983,In_678,In_815);
nand U3984 (N_3984,In_1597,In_1751);
nand U3985 (N_3985,In_2449,In_924);
nor U3986 (N_3986,In_2411,In_1391);
nor U3987 (N_3987,In_2185,In_1479);
nand U3988 (N_3988,In_2091,In_2131);
or U3989 (N_3989,In_1497,In_1434);
nor U3990 (N_3990,In_397,In_1600);
nor U3991 (N_3991,In_1076,In_128);
nor U3992 (N_3992,In_1054,In_855);
nand U3993 (N_3993,In_2068,In_1044);
nor U3994 (N_3994,In_1286,In_823);
and U3995 (N_3995,In_423,In_1616);
nand U3996 (N_3996,In_1073,In_1844);
xor U3997 (N_3997,In_134,In_2315);
nor U3998 (N_3998,In_767,In_1470);
nand U3999 (N_3999,In_2453,In_631);
nor U4000 (N_4000,In_1939,In_2338);
and U4001 (N_4001,In_80,In_1687);
or U4002 (N_4002,In_584,In_1928);
or U4003 (N_4003,In_2261,In_170);
nand U4004 (N_4004,In_1993,In_586);
xnor U4005 (N_4005,In_293,In_756);
nand U4006 (N_4006,In_1462,In_192);
xor U4007 (N_4007,In_1666,In_2430);
nor U4008 (N_4008,In_1567,In_636);
nand U4009 (N_4009,In_857,In_1807);
and U4010 (N_4010,In_562,In_375);
nor U4011 (N_4011,In_1368,In_1619);
xor U4012 (N_4012,In_1081,In_907);
xor U4013 (N_4013,In_713,In_1736);
xor U4014 (N_4014,In_1919,In_172);
nand U4015 (N_4015,In_492,In_1518);
nand U4016 (N_4016,In_929,In_590);
nor U4017 (N_4017,In_27,In_2258);
xnor U4018 (N_4018,In_923,In_1251);
and U4019 (N_4019,In_1791,In_1694);
xor U4020 (N_4020,In_1775,In_2286);
xor U4021 (N_4021,In_2128,In_1913);
xnor U4022 (N_4022,In_391,In_1304);
nor U4023 (N_4023,In_1357,In_2354);
and U4024 (N_4024,In_1891,In_492);
and U4025 (N_4025,In_1064,In_1945);
or U4026 (N_4026,In_476,In_1158);
xnor U4027 (N_4027,In_806,In_2323);
and U4028 (N_4028,In_2005,In_2327);
xor U4029 (N_4029,In_205,In_1328);
or U4030 (N_4030,In_1485,In_1740);
nand U4031 (N_4031,In_88,In_2458);
nor U4032 (N_4032,In_934,In_2191);
and U4033 (N_4033,In_872,In_1923);
nand U4034 (N_4034,In_2446,In_2340);
xor U4035 (N_4035,In_296,In_1991);
and U4036 (N_4036,In_2084,In_194);
xnor U4037 (N_4037,In_687,In_852);
nor U4038 (N_4038,In_2456,In_816);
nand U4039 (N_4039,In_1274,In_1653);
or U4040 (N_4040,In_2441,In_1326);
or U4041 (N_4041,In_1854,In_2340);
nor U4042 (N_4042,In_1398,In_2248);
and U4043 (N_4043,In_609,In_2480);
or U4044 (N_4044,In_1191,In_2462);
and U4045 (N_4045,In_2259,In_1261);
nor U4046 (N_4046,In_1269,In_743);
nor U4047 (N_4047,In_96,In_1911);
nand U4048 (N_4048,In_161,In_1336);
xnor U4049 (N_4049,In_922,In_2340);
nor U4050 (N_4050,In_37,In_1656);
and U4051 (N_4051,In_2324,In_1828);
xor U4052 (N_4052,In_241,In_1686);
xnor U4053 (N_4053,In_2176,In_2181);
or U4054 (N_4054,In_1701,In_225);
or U4055 (N_4055,In_2131,In_686);
xor U4056 (N_4056,In_1831,In_1581);
or U4057 (N_4057,In_1360,In_2282);
and U4058 (N_4058,In_343,In_376);
nand U4059 (N_4059,In_650,In_809);
nor U4060 (N_4060,In_1754,In_1924);
or U4061 (N_4061,In_1639,In_1902);
and U4062 (N_4062,In_503,In_1242);
nand U4063 (N_4063,In_423,In_359);
xor U4064 (N_4064,In_768,In_879);
nand U4065 (N_4065,In_1607,In_169);
nand U4066 (N_4066,In_152,In_2306);
xor U4067 (N_4067,In_1809,In_1656);
nand U4068 (N_4068,In_1997,In_27);
xor U4069 (N_4069,In_2009,In_1944);
or U4070 (N_4070,In_2466,In_126);
xnor U4071 (N_4071,In_1861,In_1693);
or U4072 (N_4072,In_2288,In_1417);
and U4073 (N_4073,In_678,In_1599);
or U4074 (N_4074,In_363,In_1138);
nand U4075 (N_4075,In_99,In_2226);
nand U4076 (N_4076,In_2457,In_480);
nand U4077 (N_4077,In_1565,In_2080);
or U4078 (N_4078,In_1813,In_414);
nor U4079 (N_4079,In_2129,In_346);
or U4080 (N_4080,In_419,In_2148);
or U4081 (N_4081,In_702,In_113);
and U4082 (N_4082,In_2064,In_691);
or U4083 (N_4083,In_1717,In_876);
and U4084 (N_4084,In_809,In_740);
xnor U4085 (N_4085,In_1060,In_2189);
and U4086 (N_4086,In_1262,In_1228);
xor U4087 (N_4087,In_902,In_479);
or U4088 (N_4088,In_1586,In_762);
nand U4089 (N_4089,In_250,In_1503);
nor U4090 (N_4090,In_1804,In_577);
and U4091 (N_4091,In_303,In_1430);
nand U4092 (N_4092,In_523,In_2410);
nor U4093 (N_4093,In_2097,In_637);
nor U4094 (N_4094,In_1168,In_1431);
or U4095 (N_4095,In_200,In_1595);
and U4096 (N_4096,In_2139,In_1158);
nand U4097 (N_4097,In_710,In_97);
xor U4098 (N_4098,In_646,In_115);
xnor U4099 (N_4099,In_1623,In_568);
nand U4100 (N_4100,In_65,In_2473);
nand U4101 (N_4101,In_1282,In_602);
or U4102 (N_4102,In_568,In_3);
or U4103 (N_4103,In_1239,In_2188);
and U4104 (N_4104,In_787,In_1344);
nor U4105 (N_4105,In_1287,In_950);
nand U4106 (N_4106,In_2299,In_2376);
nand U4107 (N_4107,In_1692,In_2448);
and U4108 (N_4108,In_776,In_1124);
or U4109 (N_4109,In_895,In_2285);
nor U4110 (N_4110,In_2383,In_944);
and U4111 (N_4111,In_1946,In_2164);
nand U4112 (N_4112,In_2441,In_1714);
nor U4113 (N_4113,In_2017,In_2019);
nand U4114 (N_4114,In_1985,In_1615);
xor U4115 (N_4115,In_159,In_1077);
nor U4116 (N_4116,In_671,In_2024);
nor U4117 (N_4117,In_969,In_1553);
nor U4118 (N_4118,In_1075,In_1935);
nand U4119 (N_4119,In_1336,In_1750);
or U4120 (N_4120,In_2496,In_1950);
or U4121 (N_4121,In_2010,In_1793);
or U4122 (N_4122,In_814,In_233);
and U4123 (N_4123,In_367,In_363);
or U4124 (N_4124,In_151,In_1917);
xnor U4125 (N_4125,In_744,In_2084);
or U4126 (N_4126,In_1262,In_810);
xnor U4127 (N_4127,In_428,In_171);
nand U4128 (N_4128,In_617,In_1527);
nand U4129 (N_4129,In_1473,In_1897);
xnor U4130 (N_4130,In_1656,In_675);
nor U4131 (N_4131,In_0,In_185);
xnor U4132 (N_4132,In_571,In_2076);
xnor U4133 (N_4133,In_1020,In_2432);
xor U4134 (N_4134,In_11,In_43);
or U4135 (N_4135,In_519,In_2131);
and U4136 (N_4136,In_1714,In_2318);
nor U4137 (N_4137,In_316,In_1208);
xor U4138 (N_4138,In_1744,In_1201);
nand U4139 (N_4139,In_2159,In_454);
and U4140 (N_4140,In_1228,In_999);
xnor U4141 (N_4141,In_780,In_673);
or U4142 (N_4142,In_2127,In_283);
xor U4143 (N_4143,In_1158,In_2310);
and U4144 (N_4144,In_1100,In_471);
nand U4145 (N_4145,In_1023,In_2055);
and U4146 (N_4146,In_2183,In_779);
nand U4147 (N_4147,In_1596,In_961);
nor U4148 (N_4148,In_1291,In_1688);
or U4149 (N_4149,In_981,In_528);
nor U4150 (N_4150,In_1582,In_569);
nand U4151 (N_4151,In_1230,In_2360);
xnor U4152 (N_4152,In_780,In_1888);
xor U4153 (N_4153,In_1261,In_1513);
and U4154 (N_4154,In_1278,In_2486);
xnor U4155 (N_4155,In_2374,In_2395);
and U4156 (N_4156,In_1153,In_1979);
or U4157 (N_4157,In_1151,In_1379);
or U4158 (N_4158,In_1243,In_562);
nand U4159 (N_4159,In_658,In_949);
xnor U4160 (N_4160,In_2209,In_1860);
nor U4161 (N_4161,In_1155,In_2047);
xnor U4162 (N_4162,In_991,In_1488);
and U4163 (N_4163,In_2153,In_304);
nand U4164 (N_4164,In_2351,In_245);
xnor U4165 (N_4165,In_500,In_779);
xor U4166 (N_4166,In_1085,In_1354);
or U4167 (N_4167,In_2423,In_216);
and U4168 (N_4168,In_770,In_2050);
nor U4169 (N_4169,In_1507,In_463);
and U4170 (N_4170,In_1649,In_1433);
or U4171 (N_4171,In_2044,In_413);
nor U4172 (N_4172,In_110,In_961);
nand U4173 (N_4173,In_13,In_1784);
nand U4174 (N_4174,In_188,In_575);
xnor U4175 (N_4175,In_919,In_347);
nor U4176 (N_4176,In_1906,In_243);
nand U4177 (N_4177,In_75,In_1584);
or U4178 (N_4178,In_16,In_238);
nor U4179 (N_4179,In_2497,In_155);
or U4180 (N_4180,In_1077,In_563);
or U4181 (N_4181,In_1604,In_2233);
nor U4182 (N_4182,In_461,In_610);
nor U4183 (N_4183,In_1486,In_1888);
or U4184 (N_4184,In_1357,In_730);
nor U4185 (N_4185,In_1524,In_2249);
nand U4186 (N_4186,In_1540,In_335);
xnor U4187 (N_4187,In_913,In_1811);
nor U4188 (N_4188,In_2391,In_2299);
and U4189 (N_4189,In_1272,In_1864);
nor U4190 (N_4190,In_1105,In_2371);
nand U4191 (N_4191,In_762,In_1485);
or U4192 (N_4192,In_160,In_1823);
and U4193 (N_4193,In_2057,In_193);
nor U4194 (N_4194,In_890,In_246);
xor U4195 (N_4195,In_1826,In_222);
nand U4196 (N_4196,In_2497,In_2003);
xor U4197 (N_4197,In_2088,In_2232);
and U4198 (N_4198,In_394,In_2461);
or U4199 (N_4199,In_1716,In_514);
and U4200 (N_4200,In_142,In_323);
nand U4201 (N_4201,In_200,In_504);
nand U4202 (N_4202,In_601,In_45);
nor U4203 (N_4203,In_1696,In_329);
and U4204 (N_4204,In_986,In_1547);
nand U4205 (N_4205,In_870,In_1173);
xor U4206 (N_4206,In_2092,In_2009);
and U4207 (N_4207,In_2428,In_2406);
and U4208 (N_4208,In_2417,In_1908);
xnor U4209 (N_4209,In_2189,In_1004);
and U4210 (N_4210,In_1779,In_2163);
nor U4211 (N_4211,In_300,In_1447);
nor U4212 (N_4212,In_322,In_529);
and U4213 (N_4213,In_307,In_1796);
nor U4214 (N_4214,In_1795,In_2304);
or U4215 (N_4215,In_1866,In_2467);
or U4216 (N_4216,In_1677,In_2127);
nor U4217 (N_4217,In_2490,In_74);
or U4218 (N_4218,In_2483,In_1712);
or U4219 (N_4219,In_1674,In_883);
nor U4220 (N_4220,In_1076,In_478);
or U4221 (N_4221,In_505,In_1783);
xnor U4222 (N_4222,In_2405,In_2481);
nor U4223 (N_4223,In_1180,In_2444);
nor U4224 (N_4224,In_1617,In_1431);
nand U4225 (N_4225,In_894,In_2133);
or U4226 (N_4226,In_1862,In_2322);
nand U4227 (N_4227,In_92,In_678);
nand U4228 (N_4228,In_836,In_2204);
and U4229 (N_4229,In_364,In_735);
or U4230 (N_4230,In_1075,In_657);
or U4231 (N_4231,In_717,In_1798);
xnor U4232 (N_4232,In_1829,In_725);
xor U4233 (N_4233,In_129,In_568);
and U4234 (N_4234,In_900,In_739);
xor U4235 (N_4235,In_1656,In_411);
xnor U4236 (N_4236,In_1319,In_2493);
and U4237 (N_4237,In_621,In_1912);
xnor U4238 (N_4238,In_1890,In_1610);
xnor U4239 (N_4239,In_805,In_415);
xnor U4240 (N_4240,In_1213,In_1670);
nand U4241 (N_4241,In_1000,In_1025);
and U4242 (N_4242,In_2367,In_278);
nand U4243 (N_4243,In_749,In_911);
nor U4244 (N_4244,In_868,In_504);
nand U4245 (N_4245,In_628,In_2090);
nand U4246 (N_4246,In_452,In_2375);
or U4247 (N_4247,In_1769,In_2101);
xor U4248 (N_4248,In_988,In_2237);
and U4249 (N_4249,In_706,In_1414);
and U4250 (N_4250,In_1559,In_1890);
or U4251 (N_4251,In_1641,In_1037);
nor U4252 (N_4252,In_252,In_57);
nor U4253 (N_4253,In_1613,In_2315);
nand U4254 (N_4254,In_249,In_2491);
and U4255 (N_4255,In_544,In_537);
nor U4256 (N_4256,In_1668,In_1650);
and U4257 (N_4257,In_1929,In_386);
or U4258 (N_4258,In_2186,In_900);
nor U4259 (N_4259,In_116,In_35);
and U4260 (N_4260,In_245,In_933);
nand U4261 (N_4261,In_382,In_1038);
nor U4262 (N_4262,In_1665,In_2092);
and U4263 (N_4263,In_1649,In_1673);
or U4264 (N_4264,In_1801,In_1549);
or U4265 (N_4265,In_1597,In_759);
and U4266 (N_4266,In_836,In_1948);
and U4267 (N_4267,In_1074,In_905);
or U4268 (N_4268,In_669,In_894);
or U4269 (N_4269,In_1929,In_2442);
and U4270 (N_4270,In_211,In_747);
or U4271 (N_4271,In_593,In_772);
and U4272 (N_4272,In_2195,In_1808);
nand U4273 (N_4273,In_908,In_384);
xor U4274 (N_4274,In_143,In_1434);
nor U4275 (N_4275,In_1813,In_667);
nor U4276 (N_4276,In_129,In_669);
nand U4277 (N_4277,In_1086,In_2243);
nand U4278 (N_4278,In_1179,In_1621);
and U4279 (N_4279,In_1575,In_792);
and U4280 (N_4280,In_1558,In_827);
xnor U4281 (N_4281,In_1961,In_699);
or U4282 (N_4282,In_249,In_1697);
or U4283 (N_4283,In_613,In_1766);
xor U4284 (N_4284,In_35,In_1838);
or U4285 (N_4285,In_2217,In_1307);
nor U4286 (N_4286,In_2443,In_915);
and U4287 (N_4287,In_574,In_23);
and U4288 (N_4288,In_416,In_1664);
nor U4289 (N_4289,In_1322,In_2263);
and U4290 (N_4290,In_1236,In_113);
or U4291 (N_4291,In_2367,In_649);
xnor U4292 (N_4292,In_66,In_378);
xor U4293 (N_4293,In_2304,In_1659);
nor U4294 (N_4294,In_70,In_559);
xnor U4295 (N_4295,In_1699,In_1937);
or U4296 (N_4296,In_162,In_2105);
and U4297 (N_4297,In_534,In_2028);
nor U4298 (N_4298,In_741,In_1116);
nor U4299 (N_4299,In_454,In_69);
xnor U4300 (N_4300,In_1670,In_2293);
and U4301 (N_4301,In_1856,In_1640);
and U4302 (N_4302,In_1371,In_1733);
nand U4303 (N_4303,In_2495,In_847);
nand U4304 (N_4304,In_119,In_2208);
nand U4305 (N_4305,In_480,In_1208);
nand U4306 (N_4306,In_1242,In_1727);
nor U4307 (N_4307,In_993,In_2117);
xor U4308 (N_4308,In_34,In_1145);
or U4309 (N_4309,In_230,In_191);
or U4310 (N_4310,In_1614,In_39);
xor U4311 (N_4311,In_508,In_789);
xor U4312 (N_4312,In_2112,In_43);
nand U4313 (N_4313,In_504,In_382);
nor U4314 (N_4314,In_2050,In_1283);
nor U4315 (N_4315,In_1076,In_2345);
xor U4316 (N_4316,In_1470,In_1953);
nor U4317 (N_4317,In_384,In_2298);
xor U4318 (N_4318,In_1087,In_782);
and U4319 (N_4319,In_734,In_514);
and U4320 (N_4320,In_2448,In_2121);
and U4321 (N_4321,In_1513,In_1106);
or U4322 (N_4322,In_569,In_1749);
nand U4323 (N_4323,In_171,In_1996);
nor U4324 (N_4324,In_1681,In_288);
xor U4325 (N_4325,In_969,In_2113);
xnor U4326 (N_4326,In_925,In_1276);
or U4327 (N_4327,In_1859,In_1842);
nand U4328 (N_4328,In_1489,In_1208);
and U4329 (N_4329,In_1223,In_2218);
or U4330 (N_4330,In_519,In_590);
nand U4331 (N_4331,In_471,In_1538);
and U4332 (N_4332,In_1887,In_40);
nor U4333 (N_4333,In_1046,In_1974);
and U4334 (N_4334,In_658,In_1201);
and U4335 (N_4335,In_1040,In_1286);
xnor U4336 (N_4336,In_1946,In_901);
xor U4337 (N_4337,In_1576,In_1656);
and U4338 (N_4338,In_1979,In_1074);
or U4339 (N_4339,In_1541,In_1128);
xor U4340 (N_4340,In_398,In_1237);
and U4341 (N_4341,In_2458,In_2354);
nor U4342 (N_4342,In_1137,In_1543);
nor U4343 (N_4343,In_1004,In_1173);
nand U4344 (N_4344,In_1255,In_857);
nand U4345 (N_4345,In_826,In_353);
or U4346 (N_4346,In_978,In_693);
and U4347 (N_4347,In_1964,In_2476);
and U4348 (N_4348,In_1037,In_871);
or U4349 (N_4349,In_880,In_302);
or U4350 (N_4350,In_1278,In_954);
nand U4351 (N_4351,In_372,In_723);
nor U4352 (N_4352,In_1468,In_1792);
nor U4353 (N_4353,In_304,In_120);
and U4354 (N_4354,In_2345,In_312);
xor U4355 (N_4355,In_196,In_496);
and U4356 (N_4356,In_208,In_1004);
nand U4357 (N_4357,In_1250,In_468);
nor U4358 (N_4358,In_1192,In_2226);
nor U4359 (N_4359,In_275,In_78);
and U4360 (N_4360,In_2231,In_1018);
or U4361 (N_4361,In_1704,In_1987);
nor U4362 (N_4362,In_474,In_2257);
xnor U4363 (N_4363,In_1787,In_2353);
nand U4364 (N_4364,In_1810,In_2311);
or U4365 (N_4365,In_2367,In_1481);
xor U4366 (N_4366,In_1741,In_1077);
or U4367 (N_4367,In_1591,In_110);
xnor U4368 (N_4368,In_1317,In_125);
nand U4369 (N_4369,In_1545,In_965);
xor U4370 (N_4370,In_107,In_301);
nand U4371 (N_4371,In_1913,In_511);
and U4372 (N_4372,In_2211,In_1809);
or U4373 (N_4373,In_1851,In_374);
or U4374 (N_4374,In_1437,In_1040);
xnor U4375 (N_4375,In_858,In_1943);
or U4376 (N_4376,In_1217,In_1155);
or U4377 (N_4377,In_1834,In_514);
or U4378 (N_4378,In_1154,In_1610);
and U4379 (N_4379,In_594,In_2022);
or U4380 (N_4380,In_2380,In_1406);
nand U4381 (N_4381,In_1608,In_412);
nand U4382 (N_4382,In_1931,In_426);
or U4383 (N_4383,In_403,In_780);
nand U4384 (N_4384,In_977,In_1486);
or U4385 (N_4385,In_2093,In_2157);
xor U4386 (N_4386,In_508,In_973);
or U4387 (N_4387,In_2032,In_1595);
nand U4388 (N_4388,In_1006,In_563);
nand U4389 (N_4389,In_1785,In_1480);
xnor U4390 (N_4390,In_613,In_1350);
nand U4391 (N_4391,In_1227,In_1433);
or U4392 (N_4392,In_220,In_1653);
and U4393 (N_4393,In_212,In_136);
nor U4394 (N_4394,In_1463,In_808);
nor U4395 (N_4395,In_545,In_2165);
xor U4396 (N_4396,In_1791,In_1803);
nand U4397 (N_4397,In_650,In_1455);
and U4398 (N_4398,In_1565,In_1416);
xor U4399 (N_4399,In_2493,In_1976);
nor U4400 (N_4400,In_1275,In_371);
nand U4401 (N_4401,In_875,In_1813);
nor U4402 (N_4402,In_1148,In_250);
xnor U4403 (N_4403,In_846,In_2236);
nand U4404 (N_4404,In_890,In_1276);
nor U4405 (N_4405,In_223,In_1512);
nand U4406 (N_4406,In_472,In_1301);
and U4407 (N_4407,In_524,In_281);
or U4408 (N_4408,In_313,In_2308);
xnor U4409 (N_4409,In_864,In_2493);
nand U4410 (N_4410,In_610,In_1297);
or U4411 (N_4411,In_978,In_171);
xnor U4412 (N_4412,In_2091,In_2230);
nor U4413 (N_4413,In_666,In_1386);
nor U4414 (N_4414,In_1483,In_906);
or U4415 (N_4415,In_704,In_1719);
or U4416 (N_4416,In_2487,In_988);
or U4417 (N_4417,In_417,In_1773);
nor U4418 (N_4418,In_1535,In_764);
or U4419 (N_4419,In_1197,In_1220);
nor U4420 (N_4420,In_618,In_1874);
and U4421 (N_4421,In_192,In_272);
or U4422 (N_4422,In_1527,In_1663);
nor U4423 (N_4423,In_1397,In_582);
or U4424 (N_4424,In_1194,In_599);
nand U4425 (N_4425,In_1418,In_206);
nand U4426 (N_4426,In_2048,In_309);
or U4427 (N_4427,In_1265,In_1061);
nand U4428 (N_4428,In_1280,In_1006);
nand U4429 (N_4429,In_1416,In_132);
nand U4430 (N_4430,In_2083,In_155);
or U4431 (N_4431,In_361,In_1425);
or U4432 (N_4432,In_93,In_1834);
nor U4433 (N_4433,In_2262,In_1943);
or U4434 (N_4434,In_674,In_846);
nand U4435 (N_4435,In_2462,In_1570);
nand U4436 (N_4436,In_1677,In_964);
nor U4437 (N_4437,In_924,In_862);
xor U4438 (N_4438,In_2186,In_1218);
xor U4439 (N_4439,In_1275,In_2463);
nor U4440 (N_4440,In_1480,In_2171);
nor U4441 (N_4441,In_2361,In_2471);
xnor U4442 (N_4442,In_30,In_666);
nor U4443 (N_4443,In_52,In_191);
nor U4444 (N_4444,In_2310,In_583);
xor U4445 (N_4445,In_1036,In_1139);
and U4446 (N_4446,In_859,In_2121);
or U4447 (N_4447,In_814,In_2457);
nand U4448 (N_4448,In_1727,In_177);
nor U4449 (N_4449,In_517,In_422);
xor U4450 (N_4450,In_1129,In_52);
xor U4451 (N_4451,In_184,In_1295);
nor U4452 (N_4452,In_1112,In_109);
nand U4453 (N_4453,In_710,In_2309);
nand U4454 (N_4454,In_1286,In_1485);
and U4455 (N_4455,In_2224,In_500);
nand U4456 (N_4456,In_323,In_2123);
xor U4457 (N_4457,In_1622,In_1879);
nand U4458 (N_4458,In_2384,In_2020);
xor U4459 (N_4459,In_1324,In_296);
and U4460 (N_4460,In_364,In_845);
and U4461 (N_4461,In_1948,In_319);
or U4462 (N_4462,In_2123,In_792);
xor U4463 (N_4463,In_2396,In_129);
and U4464 (N_4464,In_1666,In_1965);
and U4465 (N_4465,In_1035,In_205);
and U4466 (N_4466,In_2392,In_1751);
nor U4467 (N_4467,In_1201,In_2199);
and U4468 (N_4468,In_234,In_1835);
nor U4469 (N_4469,In_310,In_1725);
xnor U4470 (N_4470,In_2195,In_31);
nand U4471 (N_4471,In_2184,In_478);
xor U4472 (N_4472,In_1318,In_1251);
and U4473 (N_4473,In_2119,In_456);
nor U4474 (N_4474,In_1218,In_1874);
xor U4475 (N_4475,In_424,In_2120);
or U4476 (N_4476,In_1879,In_438);
nor U4477 (N_4477,In_1598,In_2455);
xnor U4478 (N_4478,In_138,In_760);
xnor U4479 (N_4479,In_1694,In_2044);
nor U4480 (N_4480,In_1503,In_912);
or U4481 (N_4481,In_1741,In_1796);
xnor U4482 (N_4482,In_477,In_1061);
xnor U4483 (N_4483,In_1115,In_1374);
nand U4484 (N_4484,In_2269,In_2387);
nor U4485 (N_4485,In_83,In_38);
xnor U4486 (N_4486,In_2366,In_657);
nand U4487 (N_4487,In_602,In_299);
and U4488 (N_4488,In_1638,In_227);
and U4489 (N_4489,In_2232,In_873);
nand U4490 (N_4490,In_1809,In_2402);
nand U4491 (N_4491,In_1851,In_1012);
nor U4492 (N_4492,In_2022,In_47);
and U4493 (N_4493,In_1592,In_2145);
and U4494 (N_4494,In_1433,In_2399);
xor U4495 (N_4495,In_1648,In_1036);
xnor U4496 (N_4496,In_2067,In_4);
and U4497 (N_4497,In_495,In_1659);
and U4498 (N_4498,In_1192,In_1734);
and U4499 (N_4499,In_248,In_1707);
and U4500 (N_4500,In_1047,In_819);
xnor U4501 (N_4501,In_1973,In_1195);
xor U4502 (N_4502,In_1826,In_1595);
nor U4503 (N_4503,In_1663,In_372);
nor U4504 (N_4504,In_34,In_2073);
nand U4505 (N_4505,In_1688,In_1878);
xnor U4506 (N_4506,In_2281,In_1150);
nand U4507 (N_4507,In_1610,In_2313);
or U4508 (N_4508,In_370,In_1640);
nand U4509 (N_4509,In_304,In_1131);
nor U4510 (N_4510,In_362,In_1000);
nand U4511 (N_4511,In_222,In_1029);
xor U4512 (N_4512,In_1033,In_582);
xor U4513 (N_4513,In_2050,In_143);
and U4514 (N_4514,In_1583,In_1593);
xnor U4515 (N_4515,In_1944,In_2079);
xnor U4516 (N_4516,In_2084,In_636);
xor U4517 (N_4517,In_2166,In_452);
or U4518 (N_4518,In_399,In_288);
nor U4519 (N_4519,In_880,In_225);
nand U4520 (N_4520,In_899,In_2464);
nand U4521 (N_4521,In_1774,In_2220);
nand U4522 (N_4522,In_1918,In_664);
nand U4523 (N_4523,In_999,In_773);
xnor U4524 (N_4524,In_493,In_822);
or U4525 (N_4525,In_975,In_1019);
or U4526 (N_4526,In_1524,In_1462);
nand U4527 (N_4527,In_2428,In_1950);
and U4528 (N_4528,In_1817,In_1605);
nand U4529 (N_4529,In_195,In_846);
and U4530 (N_4530,In_1243,In_882);
nor U4531 (N_4531,In_2031,In_2140);
xnor U4532 (N_4532,In_336,In_99);
and U4533 (N_4533,In_2158,In_632);
nand U4534 (N_4534,In_1336,In_962);
or U4535 (N_4535,In_1257,In_1764);
nor U4536 (N_4536,In_539,In_1609);
or U4537 (N_4537,In_593,In_1004);
and U4538 (N_4538,In_499,In_1301);
nor U4539 (N_4539,In_2057,In_242);
nand U4540 (N_4540,In_1803,In_692);
and U4541 (N_4541,In_1436,In_381);
xor U4542 (N_4542,In_1958,In_2498);
nor U4543 (N_4543,In_879,In_2176);
xor U4544 (N_4544,In_2203,In_1140);
or U4545 (N_4545,In_1929,In_1886);
nor U4546 (N_4546,In_2365,In_218);
nand U4547 (N_4547,In_1704,In_28);
or U4548 (N_4548,In_1997,In_1148);
nand U4549 (N_4549,In_840,In_490);
nor U4550 (N_4550,In_1803,In_1743);
or U4551 (N_4551,In_1398,In_745);
xor U4552 (N_4552,In_1257,In_808);
nor U4553 (N_4553,In_647,In_2110);
nand U4554 (N_4554,In_811,In_439);
nand U4555 (N_4555,In_330,In_928);
nand U4556 (N_4556,In_588,In_308);
nor U4557 (N_4557,In_1553,In_2244);
nand U4558 (N_4558,In_705,In_2371);
nor U4559 (N_4559,In_287,In_2429);
or U4560 (N_4560,In_1853,In_2424);
nand U4561 (N_4561,In_904,In_1047);
and U4562 (N_4562,In_1467,In_1351);
nor U4563 (N_4563,In_2330,In_821);
xor U4564 (N_4564,In_237,In_2156);
nand U4565 (N_4565,In_578,In_1287);
nand U4566 (N_4566,In_2223,In_144);
xor U4567 (N_4567,In_145,In_2227);
or U4568 (N_4568,In_1790,In_536);
nor U4569 (N_4569,In_226,In_1264);
nand U4570 (N_4570,In_426,In_549);
or U4571 (N_4571,In_1752,In_300);
and U4572 (N_4572,In_1367,In_221);
or U4573 (N_4573,In_1157,In_2007);
and U4574 (N_4574,In_216,In_2445);
and U4575 (N_4575,In_1945,In_2188);
nand U4576 (N_4576,In_1280,In_715);
xor U4577 (N_4577,In_797,In_714);
nor U4578 (N_4578,In_132,In_1695);
or U4579 (N_4579,In_290,In_2006);
or U4580 (N_4580,In_1777,In_1132);
nand U4581 (N_4581,In_1288,In_1550);
or U4582 (N_4582,In_639,In_1563);
nor U4583 (N_4583,In_127,In_1893);
or U4584 (N_4584,In_423,In_649);
or U4585 (N_4585,In_1129,In_2387);
nand U4586 (N_4586,In_462,In_178);
nor U4587 (N_4587,In_1764,In_1995);
nor U4588 (N_4588,In_1771,In_2173);
or U4589 (N_4589,In_975,In_1337);
nor U4590 (N_4590,In_1404,In_1189);
nor U4591 (N_4591,In_1275,In_1795);
and U4592 (N_4592,In_1814,In_1685);
or U4593 (N_4593,In_1316,In_1406);
and U4594 (N_4594,In_292,In_1389);
xnor U4595 (N_4595,In_1880,In_813);
or U4596 (N_4596,In_749,In_871);
nand U4597 (N_4597,In_187,In_2244);
or U4598 (N_4598,In_2491,In_224);
and U4599 (N_4599,In_1261,In_1963);
nand U4600 (N_4600,In_2076,In_1279);
xnor U4601 (N_4601,In_2174,In_1981);
or U4602 (N_4602,In_446,In_1219);
or U4603 (N_4603,In_2490,In_2427);
and U4604 (N_4604,In_291,In_140);
xor U4605 (N_4605,In_453,In_1998);
nand U4606 (N_4606,In_672,In_1717);
or U4607 (N_4607,In_460,In_2235);
and U4608 (N_4608,In_2315,In_1384);
nand U4609 (N_4609,In_13,In_761);
nand U4610 (N_4610,In_382,In_88);
nand U4611 (N_4611,In_392,In_275);
or U4612 (N_4612,In_2280,In_476);
nor U4613 (N_4613,In_1522,In_2146);
or U4614 (N_4614,In_1060,In_2408);
and U4615 (N_4615,In_1698,In_2491);
nand U4616 (N_4616,In_1271,In_608);
xnor U4617 (N_4617,In_35,In_2481);
nor U4618 (N_4618,In_156,In_1009);
nand U4619 (N_4619,In_1398,In_1308);
or U4620 (N_4620,In_1264,In_1611);
or U4621 (N_4621,In_1208,In_1269);
or U4622 (N_4622,In_2366,In_2031);
xnor U4623 (N_4623,In_1868,In_2050);
nand U4624 (N_4624,In_927,In_577);
nand U4625 (N_4625,In_1377,In_359);
xnor U4626 (N_4626,In_1221,In_915);
and U4627 (N_4627,In_1560,In_1282);
xnor U4628 (N_4628,In_2424,In_2265);
xor U4629 (N_4629,In_283,In_539);
or U4630 (N_4630,In_1354,In_2242);
or U4631 (N_4631,In_925,In_1571);
xor U4632 (N_4632,In_1272,In_2386);
xor U4633 (N_4633,In_940,In_1420);
nor U4634 (N_4634,In_99,In_1555);
nand U4635 (N_4635,In_1959,In_618);
and U4636 (N_4636,In_2210,In_857);
and U4637 (N_4637,In_994,In_680);
xor U4638 (N_4638,In_1907,In_1893);
or U4639 (N_4639,In_234,In_2182);
xnor U4640 (N_4640,In_1615,In_1240);
xnor U4641 (N_4641,In_1892,In_1919);
nor U4642 (N_4642,In_1131,In_557);
or U4643 (N_4643,In_813,In_1774);
and U4644 (N_4644,In_1625,In_235);
or U4645 (N_4645,In_119,In_2244);
nand U4646 (N_4646,In_1069,In_714);
nor U4647 (N_4647,In_81,In_294);
nand U4648 (N_4648,In_1870,In_1579);
or U4649 (N_4649,In_734,In_1051);
and U4650 (N_4650,In_986,In_2363);
nor U4651 (N_4651,In_768,In_789);
xnor U4652 (N_4652,In_613,In_1586);
and U4653 (N_4653,In_351,In_1964);
or U4654 (N_4654,In_2189,In_62);
nor U4655 (N_4655,In_2401,In_755);
and U4656 (N_4656,In_2318,In_1812);
nor U4657 (N_4657,In_1730,In_1053);
nand U4658 (N_4658,In_1073,In_79);
nand U4659 (N_4659,In_657,In_54);
xnor U4660 (N_4660,In_1869,In_153);
or U4661 (N_4661,In_981,In_1739);
or U4662 (N_4662,In_2345,In_1269);
or U4663 (N_4663,In_2090,In_2387);
nor U4664 (N_4664,In_2056,In_1440);
nand U4665 (N_4665,In_452,In_219);
nor U4666 (N_4666,In_336,In_1441);
nand U4667 (N_4667,In_2453,In_1234);
or U4668 (N_4668,In_484,In_1198);
nand U4669 (N_4669,In_1469,In_1453);
xor U4670 (N_4670,In_1332,In_658);
xnor U4671 (N_4671,In_526,In_2225);
nor U4672 (N_4672,In_584,In_1672);
and U4673 (N_4673,In_1310,In_1631);
xor U4674 (N_4674,In_2348,In_123);
nor U4675 (N_4675,In_1643,In_180);
and U4676 (N_4676,In_1100,In_1629);
xnor U4677 (N_4677,In_525,In_2466);
or U4678 (N_4678,In_73,In_370);
and U4679 (N_4679,In_1829,In_632);
or U4680 (N_4680,In_1985,In_828);
xnor U4681 (N_4681,In_2426,In_685);
xor U4682 (N_4682,In_1559,In_1282);
or U4683 (N_4683,In_1699,In_803);
nand U4684 (N_4684,In_2398,In_2209);
nor U4685 (N_4685,In_362,In_2363);
or U4686 (N_4686,In_152,In_2243);
nand U4687 (N_4687,In_279,In_1260);
xor U4688 (N_4688,In_1849,In_2185);
nor U4689 (N_4689,In_1986,In_790);
nand U4690 (N_4690,In_1221,In_1439);
nor U4691 (N_4691,In_2346,In_761);
xor U4692 (N_4692,In_93,In_1720);
and U4693 (N_4693,In_1409,In_784);
nor U4694 (N_4694,In_1172,In_186);
nand U4695 (N_4695,In_2407,In_2266);
nor U4696 (N_4696,In_508,In_2119);
nand U4697 (N_4697,In_2141,In_1453);
xnor U4698 (N_4698,In_1865,In_1015);
or U4699 (N_4699,In_2364,In_360);
nand U4700 (N_4700,In_1362,In_484);
or U4701 (N_4701,In_1475,In_859);
nand U4702 (N_4702,In_1240,In_1634);
nand U4703 (N_4703,In_1864,In_1224);
or U4704 (N_4704,In_1323,In_222);
nand U4705 (N_4705,In_1047,In_2178);
xnor U4706 (N_4706,In_1628,In_828);
or U4707 (N_4707,In_2016,In_1670);
nand U4708 (N_4708,In_2170,In_1008);
nand U4709 (N_4709,In_176,In_703);
or U4710 (N_4710,In_1048,In_234);
xnor U4711 (N_4711,In_555,In_905);
nor U4712 (N_4712,In_292,In_787);
nor U4713 (N_4713,In_373,In_477);
nand U4714 (N_4714,In_1336,In_937);
and U4715 (N_4715,In_891,In_1682);
or U4716 (N_4716,In_220,In_1507);
nor U4717 (N_4717,In_2312,In_798);
nor U4718 (N_4718,In_2459,In_509);
nor U4719 (N_4719,In_1751,In_1384);
nor U4720 (N_4720,In_1352,In_873);
and U4721 (N_4721,In_982,In_2336);
and U4722 (N_4722,In_845,In_1509);
xor U4723 (N_4723,In_2222,In_105);
nor U4724 (N_4724,In_76,In_1257);
or U4725 (N_4725,In_180,In_554);
and U4726 (N_4726,In_2145,In_1121);
nand U4727 (N_4727,In_2116,In_344);
nand U4728 (N_4728,In_571,In_1084);
xor U4729 (N_4729,In_1255,In_1899);
and U4730 (N_4730,In_404,In_151);
nor U4731 (N_4731,In_1473,In_658);
and U4732 (N_4732,In_2205,In_1786);
and U4733 (N_4733,In_1649,In_1774);
nand U4734 (N_4734,In_1890,In_2465);
or U4735 (N_4735,In_77,In_434);
or U4736 (N_4736,In_1845,In_1963);
xor U4737 (N_4737,In_1189,In_366);
or U4738 (N_4738,In_445,In_46);
nand U4739 (N_4739,In_221,In_376);
and U4740 (N_4740,In_1993,In_1454);
xnor U4741 (N_4741,In_1459,In_407);
xor U4742 (N_4742,In_176,In_260);
or U4743 (N_4743,In_903,In_601);
and U4744 (N_4744,In_1383,In_1802);
or U4745 (N_4745,In_554,In_2357);
xor U4746 (N_4746,In_1704,In_1576);
nand U4747 (N_4747,In_1484,In_2004);
or U4748 (N_4748,In_2312,In_677);
or U4749 (N_4749,In_29,In_1057);
nand U4750 (N_4750,In_1167,In_1230);
or U4751 (N_4751,In_1849,In_2340);
nor U4752 (N_4752,In_784,In_1083);
or U4753 (N_4753,In_1097,In_2161);
nand U4754 (N_4754,In_459,In_1421);
nand U4755 (N_4755,In_797,In_1358);
xor U4756 (N_4756,In_650,In_1678);
xor U4757 (N_4757,In_2356,In_1339);
and U4758 (N_4758,In_1790,In_902);
xnor U4759 (N_4759,In_2282,In_2158);
or U4760 (N_4760,In_431,In_1142);
nor U4761 (N_4761,In_2071,In_2312);
and U4762 (N_4762,In_1033,In_1895);
and U4763 (N_4763,In_2478,In_2401);
nand U4764 (N_4764,In_226,In_1111);
and U4765 (N_4765,In_1055,In_1162);
or U4766 (N_4766,In_1134,In_1428);
nor U4767 (N_4767,In_987,In_109);
xnor U4768 (N_4768,In_969,In_37);
or U4769 (N_4769,In_1929,In_968);
nand U4770 (N_4770,In_1455,In_227);
and U4771 (N_4771,In_2369,In_2042);
xnor U4772 (N_4772,In_1887,In_1214);
and U4773 (N_4773,In_1580,In_655);
and U4774 (N_4774,In_139,In_1641);
or U4775 (N_4775,In_704,In_1042);
nand U4776 (N_4776,In_446,In_587);
xnor U4777 (N_4777,In_1500,In_208);
or U4778 (N_4778,In_2050,In_1460);
nand U4779 (N_4779,In_1129,In_13);
nand U4780 (N_4780,In_1150,In_2343);
xor U4781 (N_4781,In_1182,In_122);
or U4782 (N_4782,In_18,In_2132);
or U4783 (N_4783,In_678,In_1017);
nor U4784 (N_4784,In_1182,In_1372);
nand U4785 (N_4785,In_1023,In_612);
and U4786 (N_4786,In_1557,In_1903);
nor U4787 (N_4787,In_91,In_2226);
and U4788 (N_4788,In_607,In_1246);
and U4789 (N_4789,In_1118,In_222);
nor U4790 (N_4790,In_932,In_1);
nand U4791 (N_4791,In_425,In_347);
or U4792 (N_4792,In_2205,In_1557);
or U4793 (N_4793,In_1254,In_189);
nor U4794 (N_4794,In_2103,In_1072);
nor U4795 (N_4795,In_2417,In_1716);
nor U4796 (N_4796,In_541,In_2393);
or U4797 (N_4797,In_1388,In_2303);
xnor U4798 (N_4798,In_293,In_2480);
or U4799 (N_4799,In_2258,In_735);
xnor U4800 (N_4800,In_1492,In_1213);
or U4801 (N_4801,In_576,In_958);
and U4802 (N_4802,In_2042,In_1279);
and U4803 (N_4803,In_2016,In_144);
nand U4804 (N_4804,In_2006,In_1321);
nor U4805 (N_4805,In_2154,In_1879);
nor U4806 (N_4806,In_1916,In_357);
nor U4807 (N_4807,In_1871,In_1448);
nor U4808 (N_4808,In_2116,In_155);
or U4809 (N_4809,In_1183,In_2109);
xor U4810 (N_4810,In_601,In_2474);
or U4811 (N_4811,In_616,In_1357);
nand U4812 (N_4812,In_139,In_694);
xor U4813 (N_4813,In_485,In_2170);
nor U4814 (N_4814,In_255,In_1134);
nand U4815 (N_4815,In_2354,In_881);
nor U4816 (N_4816,In_2199,In_1045);
or U4817 (N_4817,In_770,In_2268);
nand U4818 (N_4818,In_1540,In_1613);
or U4819 (N_4819,In_1702,In_1805);
nand U4820 (N_4820,In_589,In_2309);
nor U4821 (N_4821,In_1773,In_1982);
nor U4822 (N_4822,In_1059,In_794);
nand U4823 (N_4823,In_1414,In_1395);
or U4824 (N_4824,In_2206,In_1890);
or U4825 (N_4825,In_1299,In_1418);
and U4826 (N_4826,In_2215,In_1165);
and U4827 (N_4827,In_2305,In_982);
or U4828 (N_4828,In_1354,In_235);
nand U4829 (N_4829,In_157,In_1826);
nand U4830 (N_4830,In_2297,In_813);
nand U4831 (N_4831,In_21,In_158);
nand U4832 (N_4832,In_262,In_1169);
and U4833 (N_4833,In_1611,In_232);
nand U4834 (N_4834,In_2102,In_736);
xor U4835 (N_4835,In_678,In_1028);
and U4836 (N_4836,In_1679,In_1516);
xor U4837 (N_4837,In_269,In_1242);
and U4838 (N_4838,In_467,In_424);
or U4839 (N_4839,In_2458,In_2497);
nor U4840 (N_4840,In_768,In_1523);
nand U4841 (N_4841,In_1890,In_2493);
xor U4842 (N_4842,In_496,In_1154);
nor U4843 (N_4843,In_1793,In_1950);
nand U4844 (N_4844,In_2157,In_2253);
and U4845 (N_4845,In_1708,In_775);
and U4846 (N_4846,In_793,In_92);
and U4847 (N_4847,In_2356,In_2219);
nor U4848 (N_4848,In_1263,In_1780);
xor U4849 (N_4849,In_1602,In_507);
nor U4850 (N_4850,In_128,In_1986);
xor U4851 (N_4851,In_1649,In_409);
nand U4852 (N_4852,In_715,In_1062);
nor U4853 (N_4853,In_52,In_2179);
or U4854 (N_4854,In_1995,In_2293);
and U4855 (N_4855,In_1274,In_1359);
nand U4856 (N_4856,In_1789,In_1179);
xnor U4857 (N_4857,In_654,In_2078);
nand U4858 (N_4858,In_1443,In_2216);
nand U4859 (N_4859,In_2377,In_2211);
or U4860 (N_4860,In_1096,In_2303);
nand U4861 (N_4861,In_1590,In_1874);
nor U4862 (N_4862,In_1311,In_1930);
xnor U4863 (N_4863,In_1135,In_289);
nand U4864 (N_4864,In_858,In_1649);
and U4865 (N_4865,In_1723,In_1596);
nor U4866 (N_4866,In_1087,In_2440);
nor U4867 (N_4867,In_659,In_1330);
nor U4868 (N_4868,In_903,In_1723);
nor U4869 (N_4869,In_403,In_351);
or U4870 (N_4870,In_2005,In_1630);
and U4871 (N_4871,In_1153,In_1831);
and U4872 (N_4872,In_2178,In_971);
or U4873 (N_4873,In_819,In_1435);
and U4874 (N_4874,In_1224,In_299);
nor U4875 (N_4875,In_802,In_1782);
xnor U4876 (N_4876,In_1726,In_1592);
nand U4877 (N_4877,In_1430,In_893);
nor U4878 (N_4878,In_889,In_1842);
and U4879 (N_4879,In_1387,In_863);
and U4880 (N_4880,In_1255,In_983);
nor U4881 (N_4881,In_735,In_2344);
and U4882 (N_4882,In_174,In_1694);
nand U4883 (N_4883,In_937,In_577);
nand U4884 (N_4884,In_1022,In_130);
nand U4885 (N_4885,In_487,In_171);
nor U4886 (N_4886,In_2236,In_1519);
nor U4887 (N_4887,In_207,In_1487);
nand U4888 (N_4888,In_91,In_295);
nor U4889 (N_4889,In_848,In_2360);
or U4890 (N_4890,In_1428,In_153);
and U4891 (N_4891,In_1724,In_504);
nor U4892 (N_4892,In_2195,In_848);
and U4893 (N_4893,In_327,In_675);
and U4894 (N_4894,In_948,In_891);
or U4895 (N_4895,In_2205,In_172);
nor U4896 (N_4896,In_321,In_2427);
nor U4897 (N_4897,In_1080,In_483);
nand U4898 (N_4898,In_1522,In_811);
nor U4899 (N_4899,In_518,In_1852);
nor U4900 (N_4900,In_1082,In_676);
nand U4901 (N_4901,In_2400,In_818);
and U4902 (N_4902,In_686,In_1838);
and U4903 (N_4903,In_122,In_1909);
nor U4904 (N_4904,In_172,In_2094);
or U4905 (N_4905,In_1553,In_1265);
nor U4906 (N_4906,In_1479,In_1498);
nand U4907 (N_4907,In_2046,In_2032);
nand U4908 (N_4908,In_1441,In_1212);
or U4909 (N_4909,In_2489,In_96);
nand U4910 (N_4910,In_1960,In_347);
or U4911 (N_4911,In_2248,In_1860);
and U4912 (N_4912,In_1082,In_1926);
or U4913 (N_4913,In_517,In_1769);
and U4914 (N_4914,In_1313,In_398);
xor U4915 (N_4915,In_2444,In_2110);
xor U4916 (N_4916,In_803,In_1915);
or U4917 (N_4917,In_1090,In_1041);
or U4918 (N_4918,In_564,In_459);
nor U4919 (N_4919,In_666,In_2362);
nor U4920 (N_4920,In_850,In_810);
nor U4921 (N_4921,In_2421,In_1860);
xnor U4922 (N_4922,In_558,In_358);
nand U4923 (N_4923,In_1223,In_2227);
and U4924 (N_4924,In_175,In_1879);
nand U4925 (N_4925,In_2010,In_1378);
nor U4926 (N_4926,In_1209,In_2343);
nor U4927 (N_4927,In_2208,In_128);
nand U4928 (N_4928,In_2438,In_1453);
or U4929 (N_4929,In_2174,In_745);
and U4930 (N_4930,In_896,In_246);
nand U4931 (N_4931,In_1402,In_1849);
nor U4932 (N_4932,In_2445,In_969);
nand U4933 (N_4933,In_305,In_2160);
and U4934 (N_4934,In_1867,In_458);
and U4935 (N_4935,In_2317,In_242);
xor U4936 (N_4936,In_951,In_1491);
xnor U4937 (N_4937,In_2115,In_605);
nand U4938 (N_4938,In_1329,In_488);
nand U4939 (N_4939,In_200,In_1187);
nor U4940 (N_4940,In_2164,In_561);
and U4941 (N_4941,In_404,In_1026);
and U4942 (N_4942,In_2304,In_846);
nor U4943 (N_4943,In_2075,In_1266);
xor U4944 (N_4944,In_2071,In_1865);
nor U4945 (N_4945,In_1416,In_2015);
or U4946 (N_4946,In_1939,In_389);
xnor U4947 (N_4947,In_1696,In_421);
nand U4948 (N_4948,In_1169,In_2017);
xnor U4949 (N_4949,In_854,In_467);
xnor U4950 (N_4950,In_642,In_1895);
nand U4951 (N_4951,In_1906,In_1303);
and U4952 (N_4952,In_863,In_1061);
nor U4953 (N_4953,In_1120,In_1782);
or U4954 (N_4954,In_1047,In_811);
xnor U4955 (N_4955,In_905,In_391);
nor U4956 (N_4956,In_1233,In_1346);
xnor U4957 (N_4957,In_787,In_2309);
and U4958 (N_4958,In_1702,In_1620);
xor U4959 (N_4959,In_1856,In_1937);
nand U4960 (N_4960,In_2089,In_2296);
or U4961 (N_4961,In_627,In_957);
or U4962 (N_4962,In_601,In_924);
nand U4963 (N_4963,In_217,In_877);
nor U4964 (N_4964,In_2119,In_947);
and U4965 (N_4965,In_1290,In_1429);
nand U4966 (N_4966,In_2155,In_750);
xnor U4967 (N_4967,In_1041,In_1889);
and U4968 (N_4968,In_2194,In_1708);
or U4969 (N_4969,In_1958,In_1747);
xnor U4970 (N_4970,In_376,In_996);
or U4971 (N_4971,In_1020,In_1670);
xnor U4972 (N_4972,In_1929,In_1250);
and U4973 (N_4973,In_904,In_281);
nand U4974 (N_4974,In_857,In_1373);
and U4975 (N_4975,In_11,In_377);
or U4976 (N_4976,In_1027,In_1539);
nor U4977 (N_4977,In_2175,In_1804);
xor U4978 (N_4978,In_2417,In_2020);
nand U4979 (N_4979,In_722,In_279);
nand U4980 (N_4980,In_626,In_794);
nor U4981 (N_4981,In_2436,In_1231);
or U4982 (N_4982,In_159,In_209);
xor U4983 (N_4983,In_1837,In_181);
nand U4984 (N_4984,In_1686,In_1459);
nand U4985 (N_4985,In_436,In_1688);
xor U4986 (N_4986,In_1145,In_1776);
nand U4987 (N_4987,In_892,In_585);
or U4988 (N_4988,In_1302,In_2213);
nor U4989 (N_4989,In_853,In_587);
nand U4990 (N_4990,In_2313,In_342);
and U4991 (N_4991,In_1804,In_2439);
nand U4992 (N_4992,In_1168,In_2395);
or U4993 (N_4993,In_2399,In_1579);
nand U4994 (N_4994,In_1284,In_1697);
or U4995 (N_4995,In_1212,In_714);
nand U4996 (N_4996,In_1135,In_710);
nor U4997 (N_4997,In_1931,In_834);
nand U4998 (N_4998,In_1124,In_144);
and U4999 (N_4999,In_468,In_2116);
nand U5000 (N_5000,In_1803,In_1274);
nand U5001 (N_5001,In_891,In_358);
nand U5002 (N_5002,In_1525,In_1445);
or U5003 (N_5003,In_1317,In_898);
xor U5004 (N_5004,In_120,In_1098);
or U5005 (N_5005,In_685,In_1142);
nor U5006 (N_5006,In_940,In_62);
xor U5007 (N_5007,In_963,In_1293);
nand U5008 (N_5008,In_556,In_1796);
nor U5009 (N_5009,In_1139,In_1257);
nor U5010 (N_5010,In_2297,In_1852);
and U5011 (N_5011,In_2080,In_1611);
nor U5012 (N_5012,In_984,In_660);
nor U5013 (N_5013,In_735,In_1579);
nand U5014 (N_5014,In_1895,In_104);
nand U5015 (N_5015,In_899,In_1083);
nand U5016 (N_5016,In_932,In_1477);
xor U5017 (N_5017,In_1103,In_2354);
nor U5018 (N_5018,In_616,In_1660);
nand U5019 (N_5019,In_2233,In_1248);
nor U5020 (N_5020,In_457,In_410);
nor U5021 (N_5021,In_1078,In_1917);
and U5022 (N_5022,In_1051,In_2058);
or U5023 (N_5023,In_228,In_1919);
or U5024 (N_5024,In_645,In_2023);
nor U5025 (N_5025,In_89,In_1940);
nand U5026 (N_5026,In_350,In_321);
nor U5027 (N_5027,In_742,In_171);
or U5028 (N_5028,In_1282,In_87);
xor U5029 (N_5029,In_857,In_2154);
or U5030 (N_5030,In_1030,In_1285);
nor U5031 (N_5031,In_235,In_2102);
nand U5032 (N_5032,In_1156,In_1877);
or U5033 (N_5033,In_40,In_1154);
or U5034 (N_5034,In_327,In_1560);
or U5035 (N_5035,In_1036,In_15);
or U5036 (N_5036,In_777,In_1676);
or U5037 (N_5037,In_626,In_2471);
nand U5038 (N_5038,In_1797,In_1973);
or U5039 (N_5039,In_727,In_2296);
nor U5040 (N_5040,In_147,In_1120);
xnor U5041 (N_5041,In_2070,In_2317);
xnor U5042 (N_5042,In_2443,In_1828);
and U5043 (N_5043,In_444,In_2411);
and U5044 (N_5044,In_2273,In_1353);
nor U5045 (N_5045,In_1269,In_645);
xnor U5046 (N_5046,In_2010,In_1125);
and U5047 (N_5047,In_921,In_593);
or U5048 (N_5048,In_1736,In_637);
and U5049 (N_5049,In_1008,In_52);
nor U5050 (N_5050,In_2155,In_1488);
nor U5051 (N_5051,In_545,In_2359);
and U5052 (N_5052,In_1886,In_334);
xor U5053 (N_5053,In_2127,In_1863);
and U5054 (N_5054,In_247,In_768);
nand U5055 (N_5055,In_1251,In_1477);
nand U5056 (N_5056,In_30,In_2473);
xnor U5057 (N_5057,In_2332,In_1201);
xnor U5058 (N_5058,In_2354,In_205);
and U5059 (N_5059,In_445,In_2490);
and U5060 (N_5060,In_715,In_94);
xor U5061 (N_5061,In_1406,In_593);
nand U5062 (N_5062,In_925,In_491);
xnor U5063 (N_5063,In_549,In_661);
xnor U5064 (N_5064,In_693,In_1272);
or U5065 (N_5065,In_531,In_1304);
nor U5066 (N_5066,In_652,In_1614);
and U5067 (N_5067,In_1926,In_1958);
and U5068 (N_5068,In_1479,In_331);
nor U5069 (N_5069,In_646,In_2476);
nand U5070 (N_5070,In_796,In_1214);
and U5071 (N_5071,In_1336,In_1526);
or U5072 (N_5072,In_16,In_655);
nand U5073 (N_5073,In_1920,In_169);
or U5074 (N_5074,In_924,In_2137);
nand U5075 (N_5075,In_413,In_2140);
nand U5076 (N_5076,In_1012,In_1818);
xor U5077 (N_5077,In_1496,In_346);
or U5078 (N_5078,In_512,In_1780);
xor U5079 (N_5079,In_1983,In_2492);
and U5080 (N_5080,In_1932,In_1943);
and U5081 (N_5081,In_2033,In_2416);
or U5082 (N_5082,In_1841,In_1990);
or U5083 (N_5083,In_678,In_1962);
nand U5084 (N_5084,In_942,In_2365);
and U5085 (N_5085,In_317,In_488);
and U5086 (N_5086,In_744,In_682);
or U5087 (N_5087,In_1486,In_1835);
and U5088 (N_5088,In_2448,In_1415);
xor U5089 (N_5089,In_1901,In_864);
or U5090 (N_5090,In_1168,In_1916);
nor U5091 (N_5091,In_2234,In_2147);
and U5092 (N_5092,In_1723,In_455);
xor U5093 (N_5093,In_183,In_369);
or U5094 (N_5094,In_2102,In_147);
nand U5095 (N_5095,In_215,In_779);
or U5096 (N_5096,In_722,In_441);
nand U5097 (N_5097,In_2307,In_2137);
nand U5098 (N_5098,In_216,In_818);
nor U5099 (N_5099,In_1617,In_1327);
and U5100 (N_5100,In_1715,In_459);
xor U5101 (N_5101,In_1521,In_2086);
and U5102 (N_5102,In_34,In_1242);
nand U5103 (N_5103,In_948,In_2486);
nor U5104 (N_5104,In_149,In_2299);
and U5105 (N_5105,In_744,In_508);
xor U5106 (N_5106,In_140,In_2465);
nor U5107 (N_5107,In_1793,In_1244);
or U5108 (N_5108,In_659,In_494);
or U5109 (N_5109,In_2026,In_923);
xor U5110 (N_5110,In_1051,In_614);
nor U5111 (N_5111,In_1034,In_437);
nand U5112 (N_5112,In_2338,In_2288);
nor U5113 (N_5113,In_2311,In_164);
nand U5114 (N_5114,In_2496,In_1764);
and U5115 (N_5115,In_903,In_633);
and U5116 (N_5116,In_280,In_1308);
xor U5117 (N_5117,In_1192,In_1077);
or U5118 (N_5118,In_1051,In_1917);
or U5119 (N_5119,In_365,In_1533);
xnor U5120 (N_5120,In_910,In_2023);
nor U5121 (N_5121,In_1571,In_899);
nor U5122 (N_5122,In_1746,In_649);
xnor U5123 (N_5123,In_1063,In_199);
or U5124 (N_5124,In_1511,In_683);
and U5125 (N_5125,In_786,In_929);
and U5126 (N_5126,In_207,In_2228);
nor U5127 (N_5127,In_792,In_165);
or U5128 (N_5128,In_940,In_445);
nor U5129 (N_5129,In_1708,In_980);
nand U5130 (N_5130,In_1785,In_600);
nor U5131 (N_5131,In_224,In_54);
nand U5132 (N_5132,In_2224,In_1884);
or U5133 (N_5133,In_1770,In_68);
and U5134 (N_5134,In_2351,In_1744);
xnor U5135 (N_5135,In_993,In_1717);
nand U5136 (N_5136,In_385,In_538);
or U5137 (N_5137,In_985,In_1026);
xnor U5138 (N_5138,In_1090,In_984);
xnor U5139 (N_5139,In_2065,In_1789);
or U5140 (N_5140,In_102,In_2351);
xor U5141 (N_5141,In_790,In_1076);
nor U5142 (N_5142,In_354,In_2310);
or U5143 (N_5143,In_189,In_167);
nor U5144 (N_5144,In_2165,In_1731);
and U5145 (N_5145,In_2215,In_611);
or U5146 (N_5146,In_1044,In_2226);
nand U5147 (N_5147,In_1462,In_810);
or U5148 (N_5148,In_1205,In_2184);
or U5149 (N_5149,In_43,In_764);
nand U5150 (N_5150,In_2496,In_1499);
or U5151 (N_5151,In_1603,In_1422);
nor U5152 (N_5152,In_835,In_955);
or U5153 (N_5153,In_1867,In_2453);
or U5154 (N_5154,In_2423,In_1445);
xor U5155 (N_5155,In_290,In_498);
nor U5156 (N_5156,In_2090,In_2494);
xor U5157 (N_5157,In_709,In_877);
or U5158 (N_5158,In_899,In_671);
xor U5159 (N_5159,In_367,In_2061);
and U5160 (N_5160,In_1922,In_990);
and U5161 (N_5161,In_1804,In_214);
nand U5162 (N_5162,In_1357,In_879);
and U5163 (N_5163,In_1784,In_1030);
nand U5164 (N_5164,In_979,In_1249);
or U5165 (N_5165,In_2250,In_1763);
and U5166 (N_5166,In_318,In_40);
and U5167 (N_5167,In_1987,In_198);
nand U5168 (N_5168,In_1599,In_117);
nor U5169 (N_5169,In_1311,In_1621);
xnor U5170 (N_5170,In_2441,In_1763);
nand U5171 (N_5171,In_1595,In_322);
nor U5172 (N_5172,In_171,In_1263);
nor U5173 (N_5173,In_173,In_2193);
nand U5174 (N_5174,In_2167,In_1356);
nand U5175 (N_5175,In_9,In_1534);
nand U5176 (N_5176,In_1228,In_141);
xnor U5177 (N_5177,In_704,In_680);
nor U5178 (N_5178,In_2130,In_1817);
and U5179 (N_5179,In_2454,In_2070);
nand U5180 (N_5180,In_2067,In_573);
nor U5181 (N_5181,In_426,In_1903);
and U5182 (N_5182,In_1900,In_696);
xnor U5183 (N_5183,In_2008,In_667);
xor U5184 (N_5184,In_921,In_941);
and U5185 (N_5185,In_767,In_1171);
nand U5186 (N_5186,In_2427,In_1019);
nand U5187 (N_5187,In_589,In_1924);
nand U5188 (N_5188,In_325,In_1513);
and U5189 (N_5189,In_992,In_1274);
nand U5190 (N_5190,In_358,In_909);
nor U5191 (N_5191,In_2242,In_1934);
nor U5192 (N_5192,In_129,In_2259);
nand U5193 (N_5193,In_2134,In_1034);
nor U5194 (N_5194,In_2168,In_1402);
xor U5195 (N_5195,In_1010,In_787);
nor U5196 (N_5196,In_2456,In_2091);
xor U5197 (N_5197,In_2475,In_1848);
nand U5198 (N_5198,In_557,In_1902);
nand U5199 (N_5199,In_1726,In_1445);
or U5200 (N_5200,In_1320,In_1687);
nor U5201 (N_5201,In_250,In_43);
nor U5202 (N_5202,In_1648,In_1744);
or U5203 (N_5203,In_1766,In_532);
nand U5204 (N_5204,In_2327,In_2091);
nand U5205 (N_5205,In_2216,In_2488);
or U5206 (N_5206,In_2224,In_1478);
nor U5207 (N_5207,In_1213,In_2323);
or U5208 (N_5208,In_411,In_1759);
nand U5209 (N_5209,In_2436,In_1834);
and U5210 (N_5210,In_782,In_1626);
nor U5211 (N_5211,In_1133,In_70);
nor U5212 (N_5212,In_1987,In_438);
nand U5213 (N_5213,In_57,In_1275);
nand U5214 (N_5214,In_1363,In_1188);
nand U5215 (N_5215,In_1071,In_1496);
nor U5216 (N_5216,In_1769,In_1225);
xor U5217 (N_5217,In_1928,In_1373);
or U5218 (N_5218,In_2350,In_2192);
and U5219 (N_5219,In_540,In_747);
or U5220 (N_5220,In_2414,In_1864);
nor U5221 (N_5221,In_1682,In_2226);
or U5222 (N_5222,In_1008,In_2378);
nand U5223 (N_5223,In_11,In_576);
nand U5224 (N_5224,In_1176,In_1112);
nor U5225 (N_5225,In_2008,In_209);
nor U5226 (N_5226,In_1310,In_2257);
or U5227 (N_5227,In_109,In_1018);
and U5228 (N_5228,In_982,In_734);
and U5229 (N_5229,In_975,In_2055);
nor U5230 (N_5230,In_469,In_510);
nor U5231 (N_5231,In_282,In_1026);
nand U5232 (N_5232,In_1174,In_513);
nand U5233 (N_5233,In_928,In_2062);
nor U5234 (N_5234,In_404,In_1519);
nand U5235 (N_5235,In_218,In_1171);
xnor U5236 (N_5236,In_2290,In_654);
nand U5237 (N_5237,In_1351,In_37);
nor U5238 (N_5238,In_1314,In_1464);
and U5239 (N_5239,In_4,In_2010);
or U5240 (N_5240,In_232,In_1592);
xnor U5241 (N_5241,In_992,In_1592);
or U5242 (N_5242,In_1108,In_2448);
nor U5243 (N_5243,In_1759,In_1635);
or U5244 (N_5244,In_2398,In_1566);
nand U5245 (N_5245,In_944,In_1905);
and U5246 (N_5246,In_627,In_2065);
and U5247 (N_5247,In_612,In_540);
and U5248 (N_5248,In_767,In_2177);
or U5249 (N_5249,In_2134,In_429);
and U5250 (N_5250,In_2494,In_729);
nand U5251 (N_5251,In_1730,In_1628);
nor U5252 (N_5252,In_117,In_937);
and U5253 (N_5253,In_1264,In_103);
nor U5254 (N_5254,In_1455,In_1031);
nand U5255 (N_5255,In_603,In_736);
nor U5256 (N_5256,In_2074,In_1352);
xnor U5257 (N_5257,In_1602,In_1734);
nand U5258 (N_5258,In_970,In_2496);
nand U5259 (N_5259,In_1781,In_1682);
nor U5260 (N_5260,In_1245,In_180);
nor U5261 (N_5261,In_934,In_608);
nor U5262 (N_5262,In_162,In_619);
xnor U5263 (N_5263,In_2074,In_2193);
xnor U5264 (N_5264,In_2074,In_1032);
nand U5265 (N_5265,In_1461,In_1512);
xnor U5266 (N_5266,In_794,In_240);
nor U5267 (N_5267,In_485,In_1501);
xor U5268 (N_5268,In_1825,In_1036);
xnor U5269 (N_5269,In_228,In_818);
or U5270 (N_5270,In_1025,In_979);
nand U5271 (N_5271,In_2274,In_2402);
xor U5272 (N_5272,In_1411,In_100);
or U5273 (N_5273,In_1528,In_2436);
xnor U5274 (N_5274,In_1946,In_1528);
nor U5275 (N_5275,In_495,In_2286);
nand U5276 (N_5276,In_663,In_682);
xnor U5277 (N_5277,In_1922,In_2288);
xnor U5278 (N_5278,In_403,In_20);
and U5279 (N_5279,In_1514,In_1042);
xnor U5280 (N_5280,In_1800,In_428);
nand U5281 (N_5281,In_963,In_2316);
nand U5282 (N_5282,In_1880,In_1012);
nor U5283 (N_5283,In_1991,In_1427);
and U5284 (N_5284,In_960,In_1894);
nand U5285 (N_5285,In_1333,In_979);
and U5286 (N_5286,In_2410,In_1299);
nor U5287 (N_5287,In_1654,In_1460);
nor U5288 (N_5288,In_2051,In_1623);
and U5289 (N_5289,In_1932,In_1666);
nand U5290 (N_5290,In_1056,In_967);
xor U5291 (N_5291,In_1729,In_1666);
and U5292 (N_5292,In_1719,In_874);
nand U5293 (N_5293,In_588,In_750);
nand U5294 (N_5294,In_336,In_924);
xor U5295 (N_5295,In_807,In_2241);
xnor U5296 (N_5296,In_1685,In_1304);
xor U5297 (N_5297,In_672,In_1075);
and U5298 (N_5298,In_227,In_742);
and U5299 (N_5299,In_644,In_1000);
xnor U5300 (N_5300,In_1197,In_741);
nor U5301 (N_5301,In_2416,In_1938);
or U5302 (N_5302,In_2208,In_350);
or U5303 (N_5303,In_691,In_931);
or U5304 (N_5304,In_1733,In_217);
and U5305 (N_5305,In_144,In_1380);
nand U5306 (N_5306,In_1196,In_2442);
nand U5307 (N_5307,In_1425,In_285);
and U5308 (N_5308,In_2292,In_961);
nand U5309 (N_5309,In_1876,In_1845);
nand U5310 (N_5310,In_726,In_1588);
xnor U5311 (N_5311,In_1822,In_1559);
and U5312 (N_5312,In_1802,In_1795);
nor U5313 (N_5313,In_803,In_569);
xor U5314 (N_5314,In_218,In_784);
xnor U5315 (N_5315,In_65,In_2080);
nor U5316 (N_5316,In_1509,In_533);
nand U5317 (N_5317,In_563,In_2320);
nor U5318 (N_5318,In_1104,In_217);
nor U5319 (N_5319,In_226,In_1950);
xnor U5320 (N_5320,In_1135,In_2305);
or U5321 (N_5321,In_3,In_1413);
nor U5322 (N_5322,In_664,In_137);
and U5323 (N_5323,In_2266,In_641);
and U5324 (N_5324,In_86,In_2368);
or U5325 (N_5325,In_2441,In_168);
nor U5326 (N_5326,In_937,In_369);
and U5327 (N_5327,In_2148,In_1951);
or U5328 (N_5328,In_1474,In_1433);
nor U5329 (N_5329,In_1513,In_1439);
xor U5330 (N_5330,In_1301,In_2365);
or U5331 (N_5331,In_1988,In_1305);
or U5332 (N_5332,In_2062,In_2);
xnor U5333 (N_5333,In_1938,In_1960);
nand U5334 (N_5334,In_1250,In_1846);
or U5335 (N_5335,In_1468,In_826);
and U5336 (N_5336,In_941,In_2288);
xnor U5337 (N_5337,In_977,In_201);
or U5338 (N_5338,In_1431,In_505);
nor U5339 (N_5339,In_699,In_70);
and U5340 (N_5340,In_362,In_1998);
xnor U5341 (N_5341,In_491,In_1509);
nor U5342 (N_5342,In_646,In_1942);
and U5343 (N_5343,In_1852,In_437);
and U5344 (N_5344,In_2001,In_545);
or U5345 (N_5345,In_2106,In_1066);
or U5346 (N_5346,In_840,In_179);
nand U5347 (N_5347,In_1933,In_1610);
xor U5348 (N_5348,In_964,In_245);
or U5349 (N_5349,In_1904,In_1063);
xnor U5350 (N_5350,In_1626,In_441);
or U5351 (N_5351,In_1653,In_1088);
and U5352 (N_5352,In_1233,In_700);
nand U5353 (N_5353,In_1414,In_1458);
xor U5354 (N_5354,In_85,In_1823);
xor U5355 (N_5355,In_1917,In_1624);
or U5356 (N_5356,In_2207,In_737);
nor U5357 (N_5357,In_1941,In_1853);
and U5358 (N_5358,In_2100,In_195);
or U5359 (N_5359,In_2229,In_2398);
nand U5360 (N_5360,In_191,In_451);
and U5361 (N_5361,In_2204,In_505);
nor U5362 (N_5362,In_707,In_1084);
nand U5363 (N_5363,In_1202,In_1435);
nor U5364 (N_5364,In_2060,In_2370);
nand U5365 (N_5365,In_714,In_455);
nand U5366 (N_5366,In_1215,In_711);
and U5367 (N_5367,In_1050,In_2133);
or U5368 (N_5368,In_1842,In_1486);
xnor U5369 (N_5369,In_1566,In_620);
xor U5370 (N_5370,In_335,In_2151);
nor U5371 (N_5371,In_1306,In_1634);
xor U5372 (N_5372,In_2297,In_287);
and U5373 (N_5373,In_1164,In_908);
or U5374 (N_5374,In_1711,In_474);
nand U5375 (N_5375,In_2,In_2359);
or U5376 (N_5376,In_789,In_828);
nand U5377 (N_5377,In_1094,In_660);
nor U5378 (N_5378,In_253,In_1724);
or U5379 (N_5379,In_1653,In_1624);
xnor U5380 (N_5380,In_2405,In_1875);
nand U5381 (N_5381,In_589,In_1158);
and U5382 (N_5382,In_1129,In_945);
nand U5383 (N_5383,In_2062,In_1153);
nand U5384 (N_5384,In_815,In_1210);
nor U5385 (N_5385,In_2278,In_290);
xor U5386 (N_5386,In_1805,In_273);
xnor U5387 (N_5387,In_1224,In_1127);
and U5388 (N_5388,In_316,In_2229);
xnor U5389 (N_5389,In_100,In_1227);
nor U5390 (N_5390,In_423,In_832);
nor U5391 (N_5391,In_261,In_1756);
and U5392 (N_5392,In_1341,In_1006);
nor U5393 (N_5393,In_639,In_2189);
xor U5394 (N_5394,In_1985,In_1251);
xor U5395 (N_5395,In_577,In_1847);
and U5396 (N_5396,In_2008,In_1465);
and U5397 (N_5397,In_1740,In_2187);
nand U5398 (N_5398,In_534,In_586);
nand U5399 (N_5399,In_514,In_2113);
and U5400 (N_5400,In_527,In_776);
nand U5401 (N_5401,In_1861,In_2163);
nor U5402 (N_5402,In_192,In_427);
or U5403 (N_5403,In_2354,In_1997);
and U5404 (N_5404,In_2281,In_2014);
and U5405 (N_5405,In_102,In_2025);
nor U5406 (N_5406,In_288,In_498);
nand U5407 (N_5407,In_656,In_139);
or U5408 (N_5408,In_1032,In_281);
and U5409 (N_5409,In_2033,In_1814);
or U5410 (N_5410,In_15,In_2126);
xnor U5411 (N_5411,In_1745,In_1680);
or U5412 (N_5412,In_1718,In_2113);
nand U5413 (N_5413,In_710,In_1597);
xnor U5414 (N_5414,In_1187,In_1277);
xor U5415 (N_5415,In_1139,In_564);
and U5416 (N_5416,In_2452,In_739);
nand U5417 (N_5417,In_1868,In_2262);
nor U5418 (N_5418,In_1558,In_650);
nand U5419 (N_5419,In_459,In_1522);
nor U5420 (N_5420,In_325,In_827);
nand U5421 (N_5421,In_1831,In_1572);
or U5422 (N_5422,In_1657,In_1416);
or U5423 (N_5423,In_429,In_2037);
nand U5424 (N_5424,In_2224,In_857);
nor U5425 (N_5425,In_713,In_1900);
nand U5426 (N_5426,In_980,In_1816);
xnor U5427 (N_5427,In_975,In_1252);
and U5428 (N_5428,In_1484,In_2452);
or U5429 (N_5429,In_1045,In_2456);
nor U5430 (N_5430,In_1950,In_795);
and U5431 (N_5431,In_1000,In_575);
xor U5432 (N_5432,In_1221,In_979);
nor U5433 (N_5433,In_2340,In_1939);
nand U5434 (N_5434,In_1825,In_672);
and U5435 (N_5435,In_1914,In_453);
nand U5436 (N_5436,In_474,In_2354);
xnor U5437 (N_5437,In_125,In_1562);
and U5438 (N_5438,In_1078,In_801);
or U5439 (N_5439,In_1941,In_2437);
xor U5440 (N_5440,In_734,In_399);
nand U5441 (N_5441,In_240,In_638);
and U5442 (N_5442,In_204,In_188);
nor U5443 (N_5443,In_2306,In_543);
nand U5444 (N_5444,In_1601,In_2380);
nor U5445 (N_5445,In_2362,In_2377);
and U5446 (N_5446,In_849,In_1968);
xor U5447 (N_5447,In_2463,In_2212);
and U5448 (N_5448,In_1094,In_1140);
nand U5449 (N_5449,In_1864,In_1472);
or U5450 (N_5450,In_406,In_2140);
or U5451 (N_5451,In_1560,In_1164);
xnor U5452 (N_5452,In_1306,In_1643);
and U5453 (N_5453,In_1567,In_1340);
nand U5454 (N_5454,In_2001,In_437);
and U5455 (N_5455,In_307,In_2397);
or U5456 (N_5456,In_492,In_556);
and U5457 (N_5457,In_651,In_285);
nor U5458 (N_5458,In_375,In_1915);
xor U5459 (N_5459,In_2067,In_53);
nor U5460 (N_5460,In_1955,In_2336);
nor U5461 (N_5461,In_2287,In_2358);
or U5462 (N_5462,In_1766,In_2424);
nor U5463 (N_5463,In_2310,In_823);
nand U5464 (N_5464,In_1634,In_1929);
or U5465 (N_5465,In_1532,In_2332);
xor U5466 (N_5466,In_959,In_291);
nor U5467 (N_5467,In_384,In_576);
nand U5468 (N_5468,In_228,In_1241);
xnor U5469 (N_5469,In_1017,In_737);
xor U5470 (N_5470,In_1882,In_154);
nor U5471 (N_5471,In_321,In_1623);
or U5472 (N_5472,In_596,In_2353);
or U5473 (N_5473,In_55,In_183);
xor U5474 (N_5474,In_453,In_520);
or U5475 (N_5475,In_60,In_400);
xnor U5476 (N_5476,In_1978,In_1543);
or U5477 (N_5477,In_1539,In_1560);
xnor U5478 (N_5478,In_21,In_2356);
and U5479 (N_5479,In_467,In_407);
or U5480 (N_5480,In_2147,In_1764);
xor U5481 (N_5481,In_2426,In_1093);
and U5482 (N_5482,In_899,In_845);
nand U5483 (N_5483,In_1635,In_1910);
xnor U5484 (N_5484,In_1695,In_1203);
nand U5485 (N_5485,In_1350,In_88);
or U5486 (N_5486,In_492,In_98);
or U5487 (N_5487,In_868,In_2467);
nor U5488 (N_5488,In_1359,In_989);
nor U5489 (N_5489,In_1525,In_2393);
or U5490 (N_5490,In_1480,In_1759);
nand U5491 (N_5491,In_1479,In_719);
nor U5492 (N_5492,In_1048,In_1989);
or U5493 (N_5493,In_1302,In_2082);
and U5494 (N_5494,In_1659,In_817);
nand U5495 (N_5495,In_1136,In_1562);
or U5496 (N_5496,In_735,In_1383);
and U5497 (N_5497,In_416,In_1933);
xnor U5498 (N_5498,In_2136,In_1236);
nand U5499 (N_5499,In_1018,In_292);
and U5500 (N_5500,In_2245,In_1339);
nand U5501 (N_5501,In_1900,In_159);
and U5502 (N_5502,In_1372,In_1757);
nand U5503 (N_5503,In_1758,In_1342);
xor U5504 (N_5504,In_907,In_1943);
nor U5505 (N_5505,In_1745,In_2370);
or U5506 (N_5506,In_2133,In_2278);
nand U5507 (N_5507,In_2367,In_785);
nand U5508 (N_5508,In_344,In_1935);
nand U5509 (N_5509,In_264,In_1895);
xnor U5510 (N_5510,In_732,In_1754);
nand U5511 (N_5511,In_164,In_1378);
nand U5512 (N_5512,In_476,In_2371);
nor U5513 (N_5513,In_1566,In_464);
and U5514 (N_5514,In_1869,In_468);
nor U5515 (N_5515,In_2476,In_2260);
nand U5516 (N_5516,In_1281,In_1067);
or U5517 (N_5517,In_2473,In_1731);
and U5518 (N_5518,In_1107,In_1285);
nor U5519 (N_5519,In_1360,In_2450);
xnor U5520 (N_5520,In_988,In_7);
and U5521 (N_5521,In_1688,In_2042);
xnor U5522 (N_5522,In_1891,In_1617);
nor U5523 (N_5523,In_40,In_1425);
xor U5524 (N_5524,In_1811,In_2094);
nor U5525 (N_5525,In_953,In_499);
nand U5526 (N_5526,In_1697,In_1567);
nor U5527 (N_5527,In_1822,In_751);
xnor U5528 (N_5528,In_2072,In_1188);
nand U5529 (N_5529,In_2346,In_2493);
nand U5530 (N_5530,In_2367,In_1025);
nand U5531 (N_5531,In_2341,In_850);
nand U5532 (N_5532,In_1251,In_2480);
xnor U5533 (N_5533,In_770,In_1668);
or U5534 (N_5534,In_52,In_1669);
nor U5535 (N_5535,In_1989,In_392);
and U5536 (N_5536,In_1822,In_1989);
xnor U5537 (N_5537,In_1404,In_213);
nor U5538 (N_5538,In_1817,In_573);
xor U5539 (N_5539,In_193,In_2334);
nand U5540 (N_5540,In_2104,In_2065);
and U5541 (N_5541,In_677,In_987);
nand U5542 (N_5542,In_88,In_1610);
and U5543 (N_5543,In_644,In_1443);
nor U5544 (N_5544,In_1637,In_589);
nand U5545 (N_5545,In_1364,In_793);
and U5546 (N_5546,In_1172,In_1885);
and U5547 (N_5547,In_1966,In_1249);
xor U5548 (N_5548,In_1642,In_396);
nor U5549 (N_5549,In_817,In_218);
nand U5550 (N_5550,In_2393,In_387);
nor U5551 (N_5551,In_636,In_692);
nor U5552 (N_5552,In_2003,In_2252);
or U5553 (N_5553,In_743,In_2049);
xor U5554 (N_5554,In_511,In_1474);
nor U5555 (N_5555,In_2258,In_758);
xnor U5556 (N_5556,In_2390,In_1180);
nor U5557 (N_5557,In_1408,In_629);
xor U5558 (N_5558,In_2006,In_1111);
nor U5559 (N_5559,In_25,In_756);
and U5560 (N_5560,In_2472,In_857);
xnor U5561 (N_5561,In_128,In_98);
nor U5562 (N_5562,In_1738,In_2304);
nand U5563 (N_5563,In_1350,In_959);
nor U5564 (N_5564,In_522,In_1897);
or U5565 (N_5565,In_1217,In_803);
or U5566 (N_5566,In_1380,In_148);
and U5567 (N_5567,In_1682,In_487);
or U5568 (N_5568,In_1791,In_691);
nand U5569 (N_5569,In_1736,In_1004);
and U5570 (N_5570,In_2321,In_2248);
nor U5571 (N_5571,In_1172,In_1691);
nor U5572 (N_5572,In_2207,In_458);
nor U5573 (N_5573,In_885,In_1241);
and U5574 (N_5574,In_98,In_2272);
nand U5575 (N_5575,In_2246,In_106);
nand U5576 (N_5576,In_2231,In_58);
and U5577 (N_5577,In_1688,In_1226);
nand U5578 (N_5578,In_458,In_2214);
or U5579 (N_5579,In_1461,In_930);
nand U5580 (N_5580,In_2059,In_282);
nor U5581 (N_5581,In_472,In_22);
nor U5582 (N_5582,In_477,In_406);
nor U5583 (N_5583,In_964,In_1238);
or U5584 (N_5584,In_580,In_1546);
xor U5585 (N_5585,In_2035,In_1177);
xor U5586 (N_5586,In_1509,In_877);
nand U5587 (N_5587,In_222,In_1727);
nor U5588 (N_5588,In_73,In_1134);
and U5589 (N_5589,In_1308,In_1703);
nor U5590 (N_5590,In_73,In_1213);
or U5591 (N_5591,In_2476,In_477);
and U5592 (N_5592,In_1844,In_1792);
or U5593 (N_5593,In_1045,In_1031);
xor U5594 (N_5594,In_984,In_1661);
xnor U5595 (N_5595,In_2389,In_1331);
nand U5596 (N_5596,In_1191,In_467);
xnor U5597 (N_5597,In_2490,In_1427);
or U5598 (N_5598,In_959,In_2302);
and U5599 (N_5599,In_629,In_1212);
and U5600 (N_5600,In_1310,In_2035);
and U5601 (N_5601,In_2433,In_1546);
or U5602 (N_5602,In_1716,In_650);
and U5603 (N_5603,In_1340,In_904);
nand U5604 (N_5604,In_1845,In_1264);
nor U5605 (N_5605,In_350,In_1741);
and U5606 (N_5606,In_885,In_1319);
nand U5607 (N_5607,In_1345,In_1905);
or U5608 (N_5608,In_1848,In_444);
xor U5609 (N_5609,In_991,In_1427);
xor U5610 (N_5610,In_1888,In_1104);
nand U5611 (N_5611,In_876,In_205);
nand U5612 (N_5612,In_132,In_1370);
nand U5613 (N_5613,In_2480,In_147);
nand U5614 (N_5614,In_229,In_2227);
nand U5615 (N_5615,In_1108,In_1462);
or U5616 (N_5616,In_247,In_1873);
nor U5617 (N_5617,In_1959,In_1470);
xor U5618 (N_5618,In_2383,In_2422);
nand U5619 (N_5619,In_344,In_869);
nor U5620 (N_5620,In_1235,In_959);
xnor U5621 (N_5621,In_251,In_2330);
xor U5622 (N_5622,In_1014,In_1310);
nor U5623 (N_5623,In_1940,In_1298);
or U5624 (N_5624,In_2072,In_52);
xnor U5625 (N_5625,In_1343,In_2256);
nor U5626 (N_5626,In_1777,In_1431);
nor U5627 (N_5627,In_2454,In_1871);
nor U5628 (N_5628,In_281,In_405);
nor U5629 (N_5629,In_1716,In_2338);
nand U5630 (N_5630,In_444,In_1870);
nor U5631 (N_5631,In_778,In_1463);
nand U5632 (N_5632,In_2360,In_314);
nand U5633 (N_5633,In_2142,In_1833);
nand U5634 (N_5634,In_1405,In_521);
nand U5635 (N_5635,In_613,In_2060);
nand U5636 (N_5636,In_1971,In_1840);
xor U5637 (N_5637,In_1093,In_306);
or U5638 (N_5638,In_108,In_1664);
and U5639 (N_5639,In_172,In_495);
nor U5640 (N_5640,In_2255,In_1935);
xnor U5641 (N_5641,In_1492,In_1342);
and U5642 (N_5642,In_1889,In_1757);
or U5643 (N_5643,In_189,In_606);
or U5644 (N_5644,In_2225,In_1424);
nand U5645 (N_5645,In_891,In_250);
nand U5646 (N_5646,In_1155,In_2279);
nor U5647 (N_5647,In_300,In_223);
or U5648 (N_5648,In_392,In_1307);
or U5649 (N_5649,In_1743,In_1046);
nand U5650 (N_5650,In_1231,In_1415);
or U5651 (N_5651,In_1533,In_1097);
or U5652 (N_5652,In_491,In_1737);
xor U5653 (N_5653,In_2002,In_5);
nand U5654 (N_5654,In_933,In_1065);
nor U5655 (N_5655,In_904,In_802);
and U5656 (N_5656,In_334,In_464);
and U5657 (N_5657,In_190,In_1854);
and U5658 (N_5658,In_2274,In_61);
or U5659 (N_5659,In_1336,In_1917);
xor U5660 (N_5660,In_1271,In_2133);
and U5661 (N_5661,In_145,In_1322);
xor U5662 (N_5662,In_369,In_1755);
or U5663 (N_5663,In_1888,In_1996);
nand U5664 (N_5664,In_500,In_538);
or U5665 (N_5665,In_1163,In_644);
nand U5666 (N_5666,In_1423,In_168);
xnor U5667 (N_5667,In_913,In_1883);
and U5668 (N_5668,In_1154,In_1014);
or U5669 (N_5669,In_1214,In_1984);
xnor U5670 (N_5670,In_1500,In_1431);
xnor U5671 (N_5671,In_830,In_176);
nor U5672 (N_5672,In_368,In_1581);
and U5673 (N_5673,In_1957,In_939);
nand U5674 (N_5674,In_191,In_1706);
and U5675 (N_5675,In_578,In_124);
or U5676 (N_5676,In_1493,In_1402);
nor U5677 (N_5677,In_1349,In_1984);
nand U5678 (N_5678,In_1444,In_144);
nor U5679 (N_5679,In_461,In_1635);
nor U5680 (N_5680,In_988,In_659);
xor U5681 (N_5681,In_2116,In_478);
or U5682 (N_5682,In_436,In_432);
and U5683 (N_5683,In_809,In_220);
xnor U5684 (N_5684,In_2355,In_932);
and U5685 (N_5685,In_2382,In_2019);
nor U5686 (N_5686,In_542,In_1148);
nand U5687 (N_5687,In_1149,In_884);
or U5688 (N_5688,In_1791,In_99);
and U5689 (N_5689,In_1336,In_1131);
and U5690 (N_5690,In_2168,In_908);
nand U5691 (N_5691,In_628,In_2102);
nand U5692 (N_5692,In_1372,In_2236);
nor U5693 (N_5693,In_2180,In_1526);
or U5694 (N_5694,In_2349,In_1039);
nand U5695 (N_5695,In_1762,In_1602);
and U5696 (N_5696,In_289,In_1633);
or U5697 (N_5697,In_1310,In_2219);
or U5698 (N_5698,In_1625,In_1179);
nand U5699 (N_5699,In_1067,In_1815);
or U5700 (N_5700,In_91,In_1032);
nor U5701 (N_5701,In_2179,In_1679);
or U5702 (N_5702,In_920,In_630);
nor U5703 (N_5703,In_1977,In_1463);
or U5704 (N_5704,In_839,In_1917);
nand U5705 (N_5705,In_1173,In_2279);
nand U5706 (N_5706,In_717,In_924);
nand U5707 (N_5707,In_496,In_681);
xnor U5708 (N_5708,In_2114,In_967);
xor U5709 (N_5709,In_405,In_808);
nand U5710 (N_5710,In_1492,In_1276);
nor U5711 (N_5711,In_1868,In_2090);
nor U5712 (N_5712,In_305,In_1177);
nor U5713 (N_5713,In_557,In_1451);
nand U5714 (N_5714,In_2324,In_581);
nand U5715 (N_5715,In_2279,In_835);
nand U5716 (N_5716,In_1450,In_957);
xnor U5717 (N_5717,In_2260,In_2105);
xnor U5718 (N_5718,In_678,In_757);
nand U5719 (N_5719,In_2200,In_1584);
or U5720 (N_5720,In_1128,In_2148);
nand U5721 (N_5721,In_839,In_67);
xor U5722 (N_5722,In_480,In_2175);
xor U5723 (N_5723,In_1040,In_1329);
or U5724 (N_5724,In_1891,In_870);
nand U5725 (N_5725,In_1264,In_1950);
nor U5726 (N_5726,In_1514,In_591);
nor U5727 (N_5727,In_2176,In_2084);
and U5728 (N_5728,In_180,In_980);
nand U5729 (N_5729,In_2278,In_2248);
nor U5730 (N_5730,In_2198,In_1917);
nand U5731 (N_5731,In_625,In_1376);
nor U5732 (N_5732,In_74,In_1982);
nor U5733 (N_5733,In_1507,In_1379);
or U5734 (N_5734,In_1562,In_1778);
nand U5735 (N_5735,In_2393,In_485);
nor U5736 (N_5736,In_2486,In_1103);
nor U5737 (N_5737,In_276,In_1876);
or U5738 (N_5738,In_828,In_1838);
nand U5739 (N_5739,In_1444,In_15);
or U5740 (N_5740,In_671,In_2059);
or U5741 (N_5741,In_16,In_907);
and U5742 (N_5742,In_691,In_1322);
nor U5743 (N_5743,In_2221,In_312);
or U5744 (N_5744,In_244,In_587);
xnor U5745 (N_5745,In_526,In_1927);
and U5746 (N_5746,In_1077,In_240);
xor U5747 (N_5747,In_1723,In_2294);
xnor U5748 (N_5748,In_261,In_913);
or U5749 (N_5749,In_2436,In_1415);
nand U5750 (N_5750,In_2021,In_1457);
nand U5751 (N_5751,In_1033,In_116);
and U5752 (N_5752,In_421,In_2411);
nor U5753 (N_5753,In_2056,In_1978);
or U5754 (N_5754,In_280,In_849);
xnor U5755 (N_5755,In_731,In_1000);
nor U5756 (N_5756,In_1952,In_184);
nor U5757 (N_5757,In_1567,In_421);
nor U5758 (N_5758,In_1680,In_2017);
nand U5759 (N_5759,In_36,In_1409);
or U5760 (N_5760,In_119,In_292);
and U5761 (N_5761,In_57,In_1072);
nor U5762 (N_5762,In_1604,In_1195);
xnor U5763 (N_5763,In_1667,In_1727);
nor U5764 (N_5764,In_1955,In_1564);
or U5765 (N_5765,In_549,In_1612);
nand U5766 (N_5766,In_1747,In_26);
nand U5767 (N_5767,In_2457,In_484);
and U5768 (N_5768,In_2299,In_1533);
xnor U5769 (N_5769,In_777,In_2272);
nor U5770 (N_5770,In_268,In_1200);
nor U5771 (N_5771,In_1165,In_1719);
xnor U5772 (N_5772,In_725,In_1804);
nand U5773 (N_5773,In_1748,In_1872);
nand U5774 (N_5774,In_1226,In_140);
nand U5775 (N_5775,In_408,In_265);
nor U5776 (N_5776,In_1705,In_2215);
xor U5777 (N_5777,In_2025,In_2009);
and U5778 (N_5778,In_855,In_2475);
and U5779 (N_5779,In_1863,In_580);
or U5780 (N_5780,In_2424,In_1979);
xor U5781 (N_5781,In_1659,In_821);
xnor U5782 (N_5782,In_1864,In_880);
or U5783 (N_5783,In_96,In_189);
nand U5784 (N_5784,In_1248,In_1331);
xor U5785 (N_5785,In_29,In_2304);
nand U5786 (N_5786,In_1077,In_174);
nand U5787 (N_5787,In_60,In_1638);
xor U5788 (N_5788,In_767,In_1830);
nand U5789 (N_5789,In_1912,In_2259);
nor U5790 (N_5790,In_1971,In_2358);
nor U5791 (N_5791,In_1884,In_2176);
nor U5792 (N_5792,In_2109,In_1596);
xor U5793 (N_5793,In_2450,In_570);
or U5794 (N_5794,In_1455,In_617);
nand U5795 (N_5795,In_1846,In_1258);
and U5796 (N_5796,In_1305,In_13);
and U5797 (N_5797,In_810,In_2277);
nor U5798 (N_5798,In_2307,In_2256);
nor U5799 (N_5799,In_1669,In_1158);
nand U5800 (N_5800,In_1905,In_956);
and U5801 (N_5801,In_2496,In_1968);
or U5802 (N_5802,In_2029,In_2118);
or U5803 (N_5803,In_682,In_904);
nand U5804 (N_5804,In_246,In_241);
and U5805 (N_5805,In_725,In_2393);
nand U5806 (N_5806,In_1521,In_2260);
xnor U5807 (N_5807,In_1645,In_178);
nand U5808 (N_5808,In_744,In_336);
and U5809 (N_5809,In_1489,In_1649);
and U5810 (N_5810,In_1789,In_74);
and U5811 (N_5811,In_1823,In_1049);
nor U5812 (N_5812,In_1930,In_1388);
and U5813 (N_5813,In_286,In_2327);
nor U5814 (N_5814,In_56,In_2222);
or U5815 (N_5815,In_986,In_1301);
xor U5816 (N_5816,In_2406,In_1646);
and U5817 (N_5817,In_1380,In_2003);
or U5818 (N_5818,In_240,In_1985);
nor U5819 (N_5819,In_392,In_321);
or U5820 (N_5820,In_1494,In_1534);
or U5821 (N_5821,In_451,In_707);
nor U5822 (N_5822,In_2375,In_193);
nor U5823 (N_5823,In_1779,In_2353);
and U5824 (N_5824,In_1874,In_1105);
and U5825 (N_5825,In_1896,In_717);
or U5826 (N_5826,In_1055,In_188);
and U5827 (N_5827,In_650,In_617);
and U5828 (N_5828,In_1482,In_1714);
xor U5829 (N_5829,In_1427,In_2066);
nand U5830 (N_5830,In_2196,In_2233);
nand U5831 (N_5831,In_696,In_562);
nor U5832 (N_5832,In_1706,In_1728);
or U5833 (N_5833,In_1473,In_799);
nand U5834 (N_5834,In_2385,In_1895);
nand U5835 (N_5835,In_2076,In_1817);
or U5836 (N_5836,In_2459,In_1724);
or U5837 (N_5837,In_1626,In_550);
or U5838 (N_5838,In_1939,In_2031);
nand U5839 (N_5839,In_2127,In_75);
nor U5840 (N_5840,In_30,In_2184);
or U5841 (N_5841,In_609,In_1332);
xnor U5842 (N_5842,In_1219,In_2259);
and U5843 (N_5843,In_2444,In_1909);
xor U5844 (N_5844,In_2174,In_552);
or U5845 (N_5845,In_1419,In_1704);
xnor U5846 (N_5846,In_1186,In_653);
nor U5847 (N_5847,In_1801,In_2379);
or U5848 (N_5848,In_980,In_2157);
nor U5849 (N_5849,In_655,In_1179);
and U5850 (N_5850,In_1091,In_2027);
or U5851 (N_5851,In_1809,In_2226);
xor U5852 (N_5852,In_1161,In_2330);
and U5853 (N_5853,In_592,In_1813);
xnor U5854 (N_5854,In_1828,In_1687);
nand U5855 (N_5855,In_2162,In_2247);
or U5856 (N_5856,In_2263,In_90);
and U5857 (N_5857,In_1870,In_456);
xnor U5858 (N_5858,In_1236,In_2372);
xnor U5859 (N_5859,In_2115,In_2078);
or U5860 (N_5860,In_2042,In_77);
xnor U5861 (N_5861,In_70,In_2436);
or U5862 (N_5862,In_239,In_2352);
nand U5863 (N_5863,In_1530,In_121);
nand U5864 (N_5864,In_1895,In_2207);
nand U5865 (N_5865,In_196,In_2476);
and U5866 (N_5866,In_582,In_1660);
nand U5867 (N_5867,In_2006,In_2201);
xor U5868 (N_5868,In_2419,In_1248);
nand U5869 (N_5869,In_107,In_1556);
nand U5870 (N_5870,In_125,In_1454);
nor U5871 (N_5871,In_223,In_1865);
nand U5872 (N_5872,In_964,In_2131);
or U5873 (N_5873,In_2254,In_1728);
or U5874 (N_5874,In_646,In_915);
nor U5875 (N_5875,In_1992,In_827);
and U5876 (N_5876,In_2462,In_1166);
and U5877 (N_5877,In_312,In_413);
nor U5878 (N_5878,In_1451,In_1100);
and U5879 (N_5879,In_1101,In_475);
or U5880 (N_5880,In_2267,In_1437);
or U5881 (N_5881,In_592,In_153);
nand U5882 (N_5882,In_1762,In_1636);
xnor U5883 (N_5883,In_1966,In_497);
xnor U5884 (N_5884,In_552,In_1884);
xor U5885 (N_5885,In_1898,In_1525);
and U5886 (N_5886,In_1147,In_1190);
nor U5887 (N_5887,In_2010,In_99);
nor U5888 (N_5888,In_1392,In_2248);
nand U5889 (N_5889,In_1070,In_1171);
xnor U5890 (N_5890,In_956,In_2025);
xnor U5891 (N_5891,In_1919,In_1415);
nor U5892 (N_5892,In_404,In_1526);
nand U5893 (N_5893,In_2412,In_1580);
nand U5894 (N_5894,In_820,In_1875);
xor U5895 (N_5895,In_1103,In_1742);
and U5896 (N_5896,In_1245,In_319);
nor U5897 (N_5897,In_2382,In_1648);
and U5898 (N_5898,In_1537,In_1701);
nand U5899 (N_5899,In_1650,In_667);
or U5900 (N_5900,In_144,In_127);
nor U5901 (N_5901,In_756,In_587);
or U5902 (N_5902,In_1195,In_1255);
and U5903 (N_5903,In_987,In_46);
nand U5904 (N_5904,In_1678,In_1471);
nor U5905 (N_5905,In_44,In_711);
xnor U5906 (N_5906,In_760,In_656);
or U5907 (N_5907,In_2135,In_1321);
nand U5908 (N_5908,In_2396,In_578);
or U5909 (N_5909,In_1525,In_2027);
xor U5910 (N_5910,In_1962,In_2005);
nand U5911 (N_5911,In_462,In_6);
nand U5912 (N_5912,In_1916,In_2428);
nor U5913 (N_5913,In_2098,In_938);
nor U5914 (N_5914,In_847,In_845);
or U5915 (N_5915,In_2488,In_791);
nor U5916 (N_5916,In_1736,In_2143);
xor U5917 (N_5917,In_2212,In_1537);
and U5918 (N_5918,In_94,In_698);
xor U5919 (N_5919,In_1608,In_555);
nand U5920 (N_5920,In_389,In_589);
xor U5921 (N_5921,In_1887,In_397);
nand U5922 (N_5922,In_1948,In_1676);
xor U5923 (N_5923,In_748,In_1416);
or U5924 (N_5924,In_553,In_2217);
xor U5925 (N_5925,In_2227,In_1743);
nor U5926 (N_5926,In_2029,In_251);
xnor U5927 (N_5927,In_1334,In_857);
nor U5928 (N_5928,In_379,In_390);
and U5929 (N_5929,In_617,In_351);
and U5930 (N_5930,In_1571,In_1035);
or U5931 (N_5931,In_1337,In_256);
nor U5932 (N_5932,In_2186,In_2348);
xor U5933 (N_5933,In_420,In_1304);
and U5934 (N_5934,In_158,In_1625);
and U5935 (N_5935,In_1062,In_1539);
nor U5936 (N_5936,In_1246,In_1856);
xor U5937 (N_5937,In_2228,In_2398);
nor U5938 (N_5938,In_1218,In_411);
xor U5939 (N_5939,In_2036,In_1648);
nor U5940 (N_5940,In_1143,In_2488);
nor U5941 (N_5941,In_804,In_867);
nor U5942 (N_5942,In_129,In_1851);
nor U5943 (N_5943,In_978,In_440);
nand U5944 (N_5944,In_409,In_290);
nor U5945 (N_5945,In_162,In_113);
nand U5946 (N_5946,In_2012,In_2107);
and U5947 (N_5947,In_1030,In_408);
and U5948 (N_5948,In_2479,In_1660);
xnor U5949 (N_5949,In_2313,In_2306);
and U5950 (N_5950,In_512,In_2193);
or U5951 (N_5951,In_1468,In_1781);
and U5952 (N_5952,In_1476,In_283);
nand U5953 (N_5953,In_1000,In_1794);
nand U5954 (N_5954,In_1999,In_845);
nand U5955 (N_5955,In_2301,In_567);
nor U5956 (N_5956,In_2091,In_1565);
nand U5957 (N_5957,In_1551,In_2140);
nand U5958 (N_5958,In_2186,In_1671);
or U5959 (N_5959,In_2308,In_2353);
and U5960 (N_5960,In_662,In_170);
nor U5961 (N_5961,In_227,In_135);
xnor U5962 (N_5962,In_2432,In_699);
nor U5963 (N_5963,In_1116,In_135);
or U5964 (N_5964,In_2235,In_1);
nand U5965 (N_5965,In_1356,In_1911);
xor U5966 (N_5966,In_806,In_1235);
xnor U5967 (N_5967,In_1299,In_556);
xor U5968 (N_5968,In_1299,In_967);
xnor U5969 (N_5969,In_326,In_265);
xnor U5970 (N_5970,In_515,In_1143);
and U5971 (N_5971,In_549,In_271);
nand U5972 (N_5972,In_1341,In_977);
and U5973 (N_5973,In_147,In_2280);
nand U5974 (N_5974,In_634,In_421);
or U5975 (N_5975,In_190,In_1655);
xor U5976 (N_5976,In_1541,In_2387);
nor U5977 (N_5977,In_1715,In_757);
and U5978 (N_5978,In_2354,In_573);
nand U5979 (N_5979,In_196,In_1428);
and U5980 (N_5980,In_2052,In_456);
nand U5981 (N_5981,In_365,In_1853);
and U5982 (N_5982,In_131,In_1682);
nand U5983 (N_5983,In_420,In_1547);
or U5984 (N_5984,In_1164,In_1534);
nor U5985 (N_5985,In_1106,In_1726);
nor U5986 (N_5986,In_636,In_753);
nand U5987 (N_5987,In_1967,In_538);
nor U5988 (N_5988,In_933,In_572);
and U5989 (N_5989,In_1950,In_1398);
nor U5990 (N_5990,In_433,In_1614);
nor U5991 (N_5991,In_1520,In_1999);
xnor U5992 (N_5992,In_874,In_469);
and U5993 (N_5993,In_1027,In_2496);
nand U5994 (N_5994,In_698,In_1480);
or U5995 (N_5995,In_1257,In_757);
nand U5996 (N_5996,In_1849,In_431);
nor U5997 (N_5997,In_341,In_44);
and U5998 (N_5998,In_1314,In_1539);
xnor U5999 (N_5999,In_125,In_2027);
or U6000 (N_6000,In_399,In_1760);
xor U6001 (N_6001,In_397,In_1363);
and U6002 (N_6002,In_1512,In_1901);
nand U6003 (N_6003,In_954,In_553);
nor U6004 (N_6004,In_973,In_2373);
nor U6005 (N_6005,In_1452,In_2139);
xnor U6006 (N_6006,In_1020,In_1133);
xor U6007 (N_6007,In_1196,In_1030);
and U6008 (N_6008,In_1788,In_165);
or U6009 (N_6009,In_1727,In_1757);
and U6010 (N_6010,In_445,In_1256);
and U6011 (N_6011,In_1537,In_650);
xnor U6012 (N_6012,In_1335,In_340);
xnor U6013 (N_6013,In_1255,In_571);
or U6014 (N_6014,In_1412,In_515);
and U6015 (N_6015,In_2391,In_509);
nand U6016 (N_6016,In_1832,In_2334);
or U6017 (N_6017,In_1698,In_1659);
nand U6018 (N_6018,In_2098,In_1446);
nand U6019 (N_6019,In_275,In_2139);
nand U6020 (N_6020,In_120,In_1867);
nor U6021 (N_6021,In_320,In_1288);
and U6022 (N_6022,In_653,In_2108);
nand U6023 (N_6023,In_2477,In_1291);
and U6024 (N_6024,In_920,In_1143);
nor U6025 (N_6025,In_639,In_1266);
or U6026 (N_6026,In_1595,In_593);
and U6027 (N_6027,In_526,In_1133);
nand U6028 (N_6028,In_966,In_1486);
nand U6029 (N_6029,In_1143,In_148);
xnor U6030 (N_6030,In_1661,In_1857);
nor U6031 (N_6031,In_1463,In_677);
and U6032 (N_6032,In_2059,In_1261);
xnor U6033 (N_6033,In_448,In_2061);
nand U6034 (N_6034,In_241,In_1151);
nand U6035 (N_6035,In_163,In_1949);
or U6036 (N_6036,In_261,In_92);
nor U6037 (N_6037,In_720,In_671);
nand U6038 (N_6038,In_2194,In_2499);
or U6039 (N_6039,In_2163,In_1505);
or U6040 (N_6040,In_1787,In_1740);
and U6041 (N_6041,In_2059,In_270);
nor U6042 (N_6042,In_2386,In_104);
or U6043 (N_6043,In_242,In_374);
and U6044 (N_6044,In_2119,In_667);
nand U6045 (N_6045,In_902,In_2230);
nor U6046 (N_6046,In_2042,In_1008);
nor U6047 (N_6047,In_456,In_46);
nor U6048 (N_6048,In_485,In_1286);
xnor U6049 (N_6049,In_2417,In_1856);
and U6050 (N_6050,In_547,In_1657);
nand U6051 (N_6051,In_2114,In_2407);
or U6052 (N_6052,In_2110,In_2057);
and U6053 (N_6053,In_1887,In_1851);
and U6054 (N_6054,In_2150,In_1645);
and U6055 (N_6055,In_722,In_1037);
xor U6056 (N_6056,In_743,In_94);
nor U6057 (N_6057,In_912,In_1492);
and U6058 (N_6058,In_782,In_2392);
and U6059 (N_6059,In_1820,In_238);
nor U6060 (N_6060,In_1821,In_981);
and U6061 (N_6061,In_1763,In_2104);
or U6062 (N_6062,In_593,In_2495);
and U6063 (N_6063,In_2484,In_1236);
nor U6064 (N_6064,In_446,In_313);
nor U6065 (N_6065,In_1638,In_737);
and U6066 (N_6066,In_2320,In_1283);
and U6067 (N_6067,In_1866,In_928);
or U6068 (N_6068,In_714,In_1735);
or U6069 (N_6069,In_536,In_1587);
xnor U6070 (N_6070,In_1086,In_1349);
nand U6071 (N_6071,In_240,In_634);
xnor U6072 (N_6072,In_164,In_304);
nand U6073 (N_6073,In_1767,In_527);
and U6074 (N_6074,In_1880,In_2494);
nor U6075 (N_6075,In_1812,In_104);
or U6076 (N_6076,In_2202,In_2186);
xnor U6077 (N_6077,In_1963,In_2228);
nor U6078 (N_6078,In_181,In_822);
nand U6079 (N_6079,In_1634,In_2346);
nor U6080 (N_6080,In_2445,In_2232);
and U6081 (N_6081,In_1272,In_2121);
nor U6082 (N_6082,In_1354,In_2067);
and U6083 (N_6083,In_2260,In_2306);
or U6084 (N_6084,In_269,In_116);
or U6085 (N_6085,In_146,In_1130);
or U6086 (N_6086,In_2246,In_1105);
and U6087 (N_6087,In_2455,In_1635);
nor U6088 (N_6088,In_381,In_1316);
nor U6089 (N_6089,In_1265,In_2302);
xor U6090 (N_6090,In_552,In_1832);
and U6091 (N_6091,In_1706,In_2116);
xor U6092 (N_6092,In_2359,In_1082);
xnor U6093 (N_6093,In_438,In_2264);
or U6094 (N_6094,In_1536,In_439);
xnor U6095 (N_6095,In_1279,In_1894);
nand U6096 (N_6096,In_1752,In_1608);
nor U6097 (N_6097,In_959,In_2368);
xor U6098 (N_6098,In_160,In_829);
xnor U6099 (N_6099,In_575,In_1204);
and U6100 (N_6100,In_186,In_397);
and U6101 (N_6101,In_2103,In_1346);
nor U6102 (N_6102,In_2003,In_1089);
nand U6103 (N_6103,In_1759,In_1212);
and U6104 (N_6104,In_1960,In_1682);
and U6105 (N_6105,In_1344,In_1520);
or U6106 (N_6106,In_1401,In_1223);
xor U6107 (N_6107,In_417,In_2021);
or U6108 (N_6108,In_1771,In_2032);
nor U6109 (N_6109,In_93,In_175);
or U6110 (N_6110,In_1104,In_1895);
xnor U6111 (N_6111,In_431,In_164);
and U6112 (N_6112,In_968,In_857);
xor U6113 (N_6113,In_1394,In_460);
or U6114 (N_6114,In_485,In_606);
xor U6115 (N_6115,In_1103,In_1979);
nand U6116 (N_6116,In_2169,In_234);
nor U6117 (N_6117,In_1090,In_170);
and U6118 (N_6118,In_1306,In_799);
or U6119 (N_6119,In_1875,In_642);
nor U6120 (N_6120,In_2052,In_1860);
or U6121 (N_6121,In_698,In_839);
nor U6122 (N_6122,In_2181,In_643);
nor U6123 (N_6123,In_1306,In_1365);
and U6124 (N_6124,In_584,In_2437);
or U6125 (N_6125,In_1884,In_1209);
or U6126 (N_6126,In_139,In_1320);
or U6127 (N_6127,In_2226,In_468);
xor U6128 (N_6128,In_2195,In_1317);
xnor U6129 (N_6129,In_320,In_1348);
and U6130 (N_6130,In_1480,In_2462);
and U6131 (N_6131,In_1477,In_303);
nor U6132 (N_6132,In_1038,In_2420);
xnor U6133 (N_6133,In_463,In_632);
nand U6134 (N_6134,In_1741,In_1412);
and U6135 (N_6135,In_2277,In_1338);
xor U6136 (N_6136,In_69,In_1740);
nor U6137 (N_6137,In_239,In_2176);
xor U6138 (N_6138,In_2280,In_1091);
nor U6139 (N_6139,In_1214,In_845);
and U6140 (N_6140,In_2031,In_465);
and U6141 (N_6141,In_616,In_1619);
and U6142 (N_6142,In_1225,In_2000);
nor U6143 (N_6143,In_2023,In_1130);
or U6144 (N_6144,In_1806,In_1762);
nor U6145 (N_6145,In_2391,In_1510);
xnor U6146 (N_6146,In_1323,In_2445);
nand U6147 (N_6147,In_597,In_1191);
nor U6148 (N_6148,In_482,In_48);
nor U6149 (N_6149,In_1209,In_1373);
xnor U6150 (N_6150,In_273,In_1118);
nor U6151 (N_6151,In_1399,In_480);
or U6152 (N_6152,In_2425,In_2189);
nand U6153 (N_6153,In_1070,In_49);
or U6154 (N_6154,In_1715,In_2085);
nand U6155 (N_6155,In_1442,In_558);
and U6156 (N_6156,In_1440,In_353);
and U6157 (N_6157,In_958,In_95);
or U6158 (N_6158,In_794,In_2491);
nand U6159 (N_6159,In_221,In_8);
or U6160 (N_6160,In_1514,In_592);
nand U6161 (N_6161,In_1606,In_1990);
or U6162 (N_6162,In_1698,In_210);
nand U6163 (N_6163,In_1095,In_1241);
and U6164 (N_6164,In_2083,In_1724);
and U6165 (N_6165,In_2064,In_904);
xnor U6166 (N_6166,In_1221,In_337);
nand U6167 (N_6167,In_2214,In_337);
or U6168 (N_6168,In_1937,In_315);
nor U6169 (N_6169,In_2397,In_1208);
or U6170 (N_6170,In_949,In_1124);
nor U6171 (N_6171,In_2242,In_140);
nand U6172 (N_6172,In_2350,In_1297);
nor U6173 (N_6173,In_5,In_732);
or U6174 (N_6174,In_304,In_1758);
nor U6175 (N_6175,In_1753,In_2349);
xnor U6176 (N_6176,In_86,In_2269);
nor U6177 (N_6177,In_1022,In_1073);
nor U6178 (N_6178,In_1019,In_1464);
or U6179 (N_6179,In_2167,In_138);
nand U6180 (N_6180,In_26,In_2203);
or U6181 (N_6181,In_856,In_911);
nand U6182 (N_6182,In_2372,In_2478);
or U6183 (N_6183,In_299,In_1261);
or U6184 (N_6184,In_2316,In_2136);
xnor U6185 (N_6185,In_2225,In_1515);
or U6186 (N_6186,In_1832,In_758);
nor U6187 (N_6187,In_2040,In_2023);
xor U6188 (N_6188,In_1675,In_1680);
nand U6189 (N_6189,In_979,In_250);
or U6190 (N_6190,In_863,In_1975);
xnor U6191 (N_6191,In_1710,In_2177);
nor U6192 (N_6192,In_600,In_1290);
nor U6193 (N_6193,In_259,In_337);
nor U6194 (N_6194,In_1452,In_2288);
nand U6195 (N_6195,In_1685,In_2116);
xor U6196 (N_6196,In_117,In_838);
and U6197 (N_6197,In_1102,In_1935);
nor U6198 (N_6198,In_614,In_1210);
xor U6199 (N_6199,In_1792,In_1095);
nand U6200 (N_6200,In_2037,In_2363);
nor U6201 (N_6201,In_2298,In_2138);
and U6202 (N_6202,In_1396,In_872);
and U6203 (N_6203,In_1988,In_706);
xor U6204 (N_6204,In_2214,In_439);
or U6205 (N_6205,In_1632,In_2376);
nor U6206 (N_6206,In_817,In_2104);
nand U6207 (N_6207,In_993,In_1410);
or U6208 (N_6208,In_600,In_1940);
and U6209 (N_6209,In_138,In_747);
and U6210 (N_6210,In_1216,In_1786);
or U6211 (N_6211,In_1258,In_367);
nand U6212 (N_6212,In_1962,In_2234);
and U6213 (N_6213,In_1230,In_2120);
nand U6214 (N_6214,In_1399,In_1578);
nand U6215 (N_6215,In_616,In_1924);
xnor U6216 (N_6216,In_1803,In_1805);
and U6217 (N_6217,In_1119,In_1140);
nand U6218 (N_6218,In_576,In_241);
xnor U6219 (N_6219,In_490,In_2284);
xnor U6220 (N_6220,In_1074,In_1442);
xor U6221 (N_6221,In_35,In_1014);
and U6222 (N_6222,In_798,In_103);
and U6223 (N_6223,In_1200,In_2468);
and U6224 (N_6224,In_397,In_22);
nand U6225 (N_6225,In_2420,In_517);
and U6226 (N_6226,In_2341,In_467);
and U6227 (N_6227,In_166,In_1594);
and U6228 (N_6228,In_2325,In_2488);
and U6229 (N_6229,In_587,In_1245);
or U6230 (N_6230,In_2255,In_492);
and U6231 (N_6231,In_1761,In_988);
or U6232 (N_6232,In_2161,In_1970);
nand U6233 (N_6233,In_975,In_1567);
and U6234 (N_6234,In_586,In_1928);
or U6235 (N_6235,In_2158,In_1771);
nand U6236 (N_6236,In_1326,In_641);
nand U6237 (N_6237,In_943,In_143);
and U6238 (N_6238,In_1516,In_1181);
and U6239 (N_6239,In_1565,In_1843);
nor U6240 (N_6240,In_1319,In_2093);
nor U6241 (N_6241,In_2402,In_25);
nand U6242 (N_6242,In_1780,In_205);
or U6243 (N_6243,In_2147,In_2323);
nor U6244 (N_6244,In_1949,In_1234);
and U6245 (N_6245,In_1780,In_472);
and U6246 (N_6246,In_1464,In_441);
xor U6247 (N_6247,In_1383,In_489);
nand U6248 (N_6248,In_1212,In_1674);
xor U6249 (N_6249,In_1540,In_1819);
nand U6250 (N_6250,N_3252,N_952);
xnor U6251 (N_6251,N_3166,N_1475);
nor U6252 (N_6252,N_3930,N_2378);
nor U6253 (N_6253,N_4259,N_3381);
and U6254 (N_6254,N_1637,N_2973);
nor U6255 (N_6255,N_3987,N_994);
nand U6256 (N_6256,N_2521,N_5396);
nor U6257 (N_6257,N_1548,N_5758);
or U6258 (N_6258,N_2392,N_1380);
nand U6259 (N_6259,N_5838,N_1541);
nand U6260 (N_6260,N_1418,N_3031);
and U6261 (N_6261,N_2632,N_2465);
nand U6262 (N_6262,N_4734,N_2488);
nand U6263 (N_6263,N_5503,N_2054);
or U6264 (N_6264,N_2737,N_1274);
or U6265 (N_6265,N_2736,N_2027);
xnor U6266 (N_6266,N_944,N_428);
nor U6267 (N_6267,N_3374,N_103);
xnor U6268 (N_6268,N_1812,N_392);
nor U6269 (N_6269,N_1436,N_4179);
nand U6270 (N_6270,N_5827,N_4502);
and U6271 (N_6271,N_52,N_610);
and U6272 (N_6272,N_1137,N_4196);
and U6273 (N_6273,N_5303,N_1211);
xnor U6274 (N_6274,N_2038,N_55);
nand U6275 (N_6275,N_5772,N_3118);
and U6276 (N_6276,N_5698,N_1372);
nand U6277 (N_6277,N_5674,N_4093);
nor U6278 (N_6278,N_6167,N_3288);
nand U6279 (N_6279,N_1725,N_5451);
xnor U6280 (N_6280,N_4319,N_140);
or U6281 (N_6281,N_5891,N_4631);
xor U6282 (N_6282,N_2367,N_1545);
or U6283 (N_6283,N_3552,N_3078);
nand U6284 (N_6284,N_1588,N_5138);
xor U6285 (N_6285,N_808,N_5593);
xnor U6286 (N_6286,N_426,N_4853);
xor U6287 (N_6287,N_720,N_3097);
or U6288 (N_6288,N_1697,N_4885);
nand U6289 (N_6289,N_3316,N_2881);
or U6290 (N_6290,N_3787,N_1653);
xnor U6291 (N_6291,N_1673,N_3223);
nand U6292 (N_6292,N_3085,N_2398);
and U6293 (N_6293,N_6068,N_2251);
nand U6294 (N_6294,N_911,N_1424);
nor U6295 (N_6295,N_2074,N_6165);
nor U6296 (N_6296,N_413,N_5455);
xnor U6297 (N_6297,N_2180,N_3041);
and U6298 (N_6298,N_3120,N_4967);
or U6299 (N_6299,N_675,N_4619);
and U6300 (N_6300,N_3944,N_5633);
or U6301 (N_6301,N_4186,N_4121);
nand U6302 (N_6302,N_3047,N_4690);
and U6303 (N_6303,N_1707,N_3848);
nand U6304 (N_6304,N_327,N_3111);
or U6305 (N_6305,N_3654,N_954);
and U6306 (N_6306,N_5897,N_2695);
nor U6307 (N_6307,N_772,N_4830);
nand U6308 (N_6308,N_2536,N_2133);
nand U6309 (N_6309,N_1285,N_1013);
nand U6310 (N_6310,N_975,N_1757);
or U6311 (N_6311,N_4035,N_3967);
or U6312 (N_6312,N_5843,N_831);
or U6313 (N_6313,N_4531,N_3940);
nor U6314 (N_6314,N_5069,N_1605);
nor U6315 (N_6315,N_1534,N_2086);
and U6316 (N_6316,N_4114,N_3007);
nor U6317 (N_6317,N_167,N_4626);
nand U6318 (N_6318,N_5850,N_5228);
and U6319 (N_6319,N_3346,N_1549);
or U6320 (N_6320,N_1472,N_1406);
or U6321 (N_6321,N_5510,N_1983);
and U6322 (N_6322,N_5444,N_264);
nand U6323 (N_6323,N_3715,N_955);
xor U6324 (N_6324,N_3331,N_483);
or U6325 (N_6325,N_1842,N_3501);
or U6326 (N_6326,N_3993,N_3470);
and U6327 (N_6327,N_2933,N_4071);
xor U6328 (N_6328,N_1815,N_4863);
nor U6329 (N_6329,N_2958,N_1802);
nor U6330 (N_6330,N_2419,N_2513);
nor U6331 (N_6331,N_2360,N_5501);
or U6332 (N_6332,N_3990,N_5290);
xor U6333 (N_6333,N_2350,N_94);
nor U6334 (N_6334,N_5149,N_2598);
nor U6335 (N_6335,N_280,N_4498);
xnor U6336 (N_6336,N_539,N_3774);
or U6337 (N_6337,N_4563,N_524);
nor U6338 (N_6338,N_5110,N_1691);
and U6339 (N_6339,N_1165,N_4209);
and U6340 (N_6340,N_3587,N_4416);
or U6341 (N_6341,N_2742,N_5447);
nand U6342 (N_6342,N_613,N_1682);
or U6343 (N_6343,N_1944,N_1112);
nor U6344 (N_6344,N_5515,N_2222);
nand U6345 (N_6345,N_836,N_6189);
or U6346 (N_6346,N_4595,N_3926);
or U6347 (N_6347,N_5944,N_521);
nand U6348 (N_6348,N_4906,N_602);
nor U6349 (N_6349,N_4581,N_5927);
xor U6350 (N_6350,N_4213,N_5158);
nand U6351 (N_6351,N_69,N_3126);
xnor U6352 (N_6352,N_845,N_5459);
nand U6353 (N_6353,N_5300,N_5872);
or U6354 (N_6354,N_3415,N_2238);
or U6355 (N_6355,N_1024,N_4777);
and U6356 (N_6356,N_1870,N_1781);
nor U6357 (N_6357,N_2965,N_3686);
nor U6358 (N_6358,N_3218,N_396);
or U6359 (N_6359,N_395,N_1578);
or U6360 (N_6360,N_3991,N_697);
or U6361 (N_6361,N_3543,N_3580);
nor U6362 (N_6362,N_1095,N_25);
nand U6363 (N_6363,N_699,N_484);
and U6364 (N_6364,N_2905,N_3358);
xor U6365 (N_6365,N_4408,N_1338);
nor U6366 (N_6366,N_5449,N_3469);
nand U6367 (N_6367,N_1369,N_3795);
nand U6368 (N_6368,N_4284,N_5619);
and U6369 (N_6369,N_3095,N_1083);
xor U6370 (N_6370,N_3464,N_4986);
and U6371 (N_6371,N_4676,N_1167);
xor U6372 (N_6372,N_4660,N_4288);
xnor U6373 (N_6373,N_862,N_3716);
xnor U6374 (N_6374,N_3196,N_5097);
xnor U6375 (N_6375,N_3780,N_329);
or U6376 (N_6376,N_4350,N_4265);
and U6377 (N_6377,N_544,N_3411);
or U6378 (N_6378,N_1645,N_1303);
and U6379 (N_6379,N_4696,N_3599);
or U6380 (N_6380,N_5614,N_4098);
or U6381 (N_6381,N_3348,N_13);
and U6382 (N_6382,N_4804,N_3513);
nand U6383 (N_6383,N_4836,N_3073);
or U6384 (N_6384,N_734,N_3856);
and U6385 (N_6385,N_3386,N_2387);
or U6386 (N_6386,N_4720,N_1867);
or U6387 (N_6387,N_4026,N_5150);
and U6388 (N_6388,N_3682,N_3149);
or U6389 (N_6389,N_3375,N_3801);
nor U6390 (N_6390,N_2593,N_5479);
nor U6391 (N_6391,N_4282,N_5932);
xnor U6392 (N_6392,N_4617,N_2672);
nand U6393 (N_6393,N_4647,N_515);
nand U6394 (N_6394,N_5775,N_894);
nand U6395 (N_6395,N_5175,N_4207);
or U6396 (N_6396,N_1041,N_3495);
or U6397 (N_6397,N_2008,N_2418);
nor U6398 (N_6398,N_3498,N_382);
xor U6399 (N_6399,N_243,N_5737);
or U6400 (N_6400,N_2166,N_2297);
and U6401 (N_6401,N_2040,N_3918);
and U6402 (N_6402,N_3760,N_4464);
nand U6403 (N_6403,N_670,N_5880);
and U6404 (N_6404,N_1473,N_3979);
nand U6405 (N_6405,N_2510,N_4642);
and U6406 (N_6406,N_3623,N_3924);
nor U6407 (N_6407,N_2799,N_3763);
xor U6408 (N_6408,N_2315,N_673);
xor U6409 (N_6409,N_709,N_5728);
nand U6410 (N_6410,N_5990,N_2275);
nand U6411 (N_6411,N_784,N_4216);
nor U6412 (N_6412,N_5969,N_3185);
nor U6413 (N_6413,N_199,N_4152);
or U6414 (N_6414,N_5180,N_1139);
or U6415 (N_6415,N_4362,N_3884);
and U6416 (N_6416,N_1513,N_5974);
or U6417 (N_6417,N_525,N_4226);
nor U6418 (N_6418,N_4508,N_852);
nand U6419 (N_6419,N_2030,N_2851);
nor U6420 (N_6420,N_2191,N_2997);
xnor U6421 (N_6421,N_171,N_3536);
xnor U6422 (N_6422,N_393,N_5387);
xnor U6423 (N_6423,N_6040,N_3515);
xnor U6424 (N_6424,N_989,N_795);
and U6425 (N_6425,N_586,N_5170);
and U6426 (N_6426,N_2753,N_3402);
or U6427 (N_6427,N_5031,N_5399);
or U6428 (N_6428,N_3932,N_109);
xnor U6429 (N_6429,N_82,N_702);
and U6430 (N_6430,N_998,N_3838);
or U6431 (N_6431,N_4477,N_6194);
xnor U6432 (N_6432,N_1016,N_4033);
xnor U6433 (N_6433,N_4238,N_2535);
and U6434 (N_6434,N_3131,N_481);
or U6435 (N_6435,N_4530,N_3002);
nor U6436 (N_6436,N_3224,N_2940);
nor U6437 (N_6437,N_5469,N_1808);
and U6438 (N_6438,N_4818,N_6172);
xor U6439 (N_6439,N_7,N_3836);
and U6440 (N_6440,N_5032,N_3009);
xor U6441 (N_6441,N_3459,N_5085);
nor U6442 (N_6442,N_2670,N_2969);
xor U6443 (N_6443,N_4515,N_3554);
nor U6444 (N_6444,N_4507,N_21);
xnor U6445 (N_6445,N_1442,N_1845);
or U6446 (N_6446,N_2490,N_1580);
nand U6447 (N_6447,N_3326,N_2199);
xor U6448 (N_6448,N_4178,N_2907);
nand U6449 (N_6449,N_4234,N_1130);
and U6450 (N_6450,N_4333,N_3973);
nor U6451 (N_6451,N_1576,N_4633);
nand U6452 (N_6452,N_4680,N_3395);
nand U6453 (N_6453,N_3817,N_4841);
nand U6454 (N_6454,N_3075,N_5721);
and U6455 (N_6455,N_4629,N_3440);
and U6456 (N_6456,N_1689,N_3865);
and U6457 (N_6457,N_2331,N_5505);
and U6458 (N_6458,N_6170,N_5687);
or U6459 (N_6459,N_4048,N_2452);
and U6460 (N_6460,N_1203,N_2896);
and U6461 (N_6461,N_148,N_1055);
nand U6462 (N_6462,N_1098,N_1765);
or U6463 (N_6463,N_6162,N_5006);
and U6464 (N_6464,N_4052,N_5136);
and U6465 (N_6465,N_2467,N_2366);
nand U6466 (N_6466,N_569,N_498);
xnor U6467 (N_6467,N_5200,N_2173);
nand U6468 (N_6468,N_839,N_2639);
nor U6469 (N_6469,N_5125,N_3363);
xnor U6470 (N_6470,N_1672,N_686);
xnor U6471 (N_6471,N_3544,N_4274);
xnor U6472 (N_6472,N_4666,N_2286);
or U6473 (N_6473,N_2211,N_2061);
nor U6474 (N_6474,N_4322,N_600);
nor U6475 (N_6475,N_5852,N_1492);
and U6476 (N_6476,N_4807,N_5021);
xor U6477 (N_6477,N_1684,N_1599);
nand U6478 (N_6478,N_2414,N_4711);
or U6479 (N_6479,N_3471,N_1351);
and U6480 (N_6480,N_1556,N_6073);
or U6481 (N_6481,N_6206,N_2287);
nor U6482 (N_6482,N_508,N_2270);
or U6483 (N_6483,N_4598,N_32);
or U6484 (N_6484,N_3908,N_2817);
nand U6485 (N_6485,N_1177,N_4871);
nor U6486 (N_6486,N_4227,N_472);
nand U6487 (N_6487,N_5322,N_864);
or U6488 (N_6488,N_2487,N_3455);
nand U6489 (N_6489,N_186,N_3614);
xor U6490 (N_6490,N_651,N_2635);
nor U6491 (N_6491,N_5934,N_5871);
nand U6492 (N_6492,N_2236,N_5168);
xnor U6493 (N_6493,N_448,N_5608);
xor U6494 (N_6494,N_3633,N_231);
nand U6495 (N_6495,N_2206,N_5511);
nand U6496 (N_6496,N_5744,N_5845);
nor U6497 (N_6497,N_242,N_4966);
nand U6498 (N_6498,N_4389,N_5561);
and U6499 (N_6499,N_1195,N_4602);
xnor U6500 (N_6500,N_4937,N_3273);
xnor U6501 (N_6501,N_3893,N_3858);
xor U6502 (N_6502,N_2468,N_6061);
or U6503 (N_6503,N_464,N_2356);
and U6504 (N_6504,N_6174,N_3508);
and U6505 (N_6505,N_2050,N_5718);
xnor U6506 (N_6506,N_885,N_2200);
and U6507 (N_6507,N_6004,N_5206);
and U6508 (N_6508,N_5128,N_5916);
nand U6509 (N_6509,N_5063,N_2391);
or U6510 (N_6510,N_3767,N_169);
or U6511 (N_6511,N_1454,N_1566);
nand U6512 (N_6512,N_5985,N_4092);
nor U6513 (N_6513,N_3753,N_5724);
and U6514 (N_6514,N_603,N_4870);
xor U6515 (N_6515,N_1451,N_5693);
and U6516 (N_6516,N_6136,N_5950);
and U6517 (N_6517,N_4821,N_283);
or U6518 (N_6518,N_5291,N_833);
nand U6519 (N_6519,N_2539,N_3122);
and U6520 (N_6520,N_4010,N_3425);
nand U6521 (N_6521,N_3779,N_4847);
nand U6522 (N_6522,N_4089,N_2728);
and U6523 (N_6523,N_793,N_4131);
or U6524 (N_6524,N_114,N_3006);
or U6525 (N_6525,N_3446,N_4269);
or U6526 (N_6526,N_3844,N_5304);
nand U6527 (N_6527,N_4180,N_4046);
or U6528 (N_6528,N_4969,N_0);
or U6529 (N_6529,N_553,N_1897);
or U6530 (N_6530,N_2085,N_1886);
or U6531 (N_6531,N_3190,N_5155);
nor U6532 (N_6532,N_1124,N_2461);
xnor U6533 (N_6533,N_1467,N_1106);
or U6534 (N_6534,N_6173,N_1419);
xor U6535 (N_6535,N_2897,N_5904);
nand U6536 (N_6536,N_4536,N_4618);
nor U6537 (N_6537,N_6044,N_2503);
or U6538 (N_6538,N_6049,N_3879);
and U6539 (N_6539,N_1660,N_5480);
nor U6540 (N_6540,N_5671,N_5745);
nor U6541 (N_6541,N_732,N_3866);
or U6542 (N_6542,N_1162,N_4560);
and U6543 (N_6543,N_1706,N_5377);
xnor U6544 (N_6544,N_1030,N_4055);
and U6545 (N_6545,N_1289,N_3448);
xor U6546 (N_6546,N_1594,N_2454);
or U6547 (N_6547,N_2499,N_4215);
or U6548 (N_6548,N_3917,N_5878);
nor U6549 (N_6549,N_764,N_1178);
nand U6550 (N_6550,N_4294,N_3761);
xnor U6551 (N_6551,N_4997,N_2372);
and U6552 (N_6552,N_6090,N_5263);
nand U6553 (N_6553,N_4625,N_2921);
nand U6554 (N_6554,N_678,N_93);
nand U6555 (N_6555,N_3164,N_1053);
nand U6556 (N_6556,N_2502,N_3782);
and U6557 (N_6557,N_3839,N_2956);
nand U6558 (N_6558,N_4047,N_2150);
nand U6559 (N_6559,N_1817,N_2244);
nor U6560 (N_6560,N_5363,N_4231);
nand U6561 (N_6561,N_829,N_2225);
or U6562 (N_6562,N_2435,N_4664);
or U6563 (N_6563,N_2332,N_6159);
or U6564 (N_6564,N_6239,N_4535);
or U6565 (N_6565,N_1528,N_5317);
nand U6566 (N_6566,N_1266,N_2272);
nor U6567 (N_6567,N_3328,N_1611);
and U6568 (N_6568,N_4988,N_3796);
xnor U6569 (N_6569,N_3758,N_3127);
xnor U6570 (N_6570,N_837,N_1606);
xor U6571 (N_6571,N_3863,N_1969);
nand U6572 (N_6572,N_917,N_5389);
xor U6573 (N_6573,N_306,N_4669);
nand U6574 (N_6574,N_791,N_1929);
nand U6575 (N_6575,N_2010,N_2328);
xor U6576 (N_6576,N_644,N_715);
nand U6577 (N_6577,N_3886,N_1771);
nor U6578 (N_6578,N_5244,N_4246);
nor U6579 (N_6579,N_4199,N_2748);
xnor U6580 (N_6580,N_5338,N_6130);
nand U6581 (N_6581,N_4099,N_2966);
nand U6582 (N_6582,N_3861,N_10);
nor U6583 (N_6583,N_2928,N_2051);
nor U6584 (N_6584,N_981,N_5020);
and U6585 (N_6585,N_4165,N_680);
nor U6586 (N_6586,N_4414,N_2589);
xor U6587 (N_6587,N_4214,N_3750);
xnor U6588 (N_6588,N_1311,N_4557);
or U6589 (N_6589,N_1242,N_3809);
nand U6590 (N_6590,N_147,N_1168);
and U6591 (N_6591,N_3862,N_4205);
nor U6592 (N_6592,N_1950,N_2285);
or U6593 (N_6593,N_4086,N_2101);
and U6594 (N_6594,N_2570,N_1038);
and U6595 (N_6595,N_3921,N_2825);
xnor U6596 (N_6596,N_6238,N_5009);
xnor U6597 (N_6597,N_3671,N_984);
nor U6598 (N_6598,N_26,N_1820);
nand U6599 (N_6599,N_2919,N_5776);
nand U6600 (N_6600,N_1863,N_3632);
xor U6601 (N_6601,N_5905,N_5488);
and U6602 (N_6602,N_4174,N_4481);
xor U6603 (N_6603,N_3260,N_2738);
nand U6604 (N_6604,N_698,N_2479);
nand U6605 (N_6605,N_3933,N_4400);
and U6606 (N_6606,N_3883,N_3871);
nor U6607 (N_6607,N_4023,N_1364);
xor U6608 (N_6608,N_3029,N_1490);
xor U6609 (N_6609,N_3188,N_3216);
and U6610 (N_6610,N_260,N_3390);
nand U6611 (N_6611,N_3821,N_4074);
and U6612 (N_6612,N_466,N_6135);
nor U6613 (N_6613,N_6151,N_1826);
or U6614 (N_6614,N_6228,N_4298);
nor U6615 (N_6615,N_3627,N_3345);
and U6616 (N_6616,N_558,N_3657);
nand U6617 (N_6617,N_1743,N_5749);
or U6618 (N_6618,N_2795,N_1184);
or U6619 (N_6619,N_3943,N_2469);
or U6620 (N_6620,N_2717,N_3562);
and U6621 (N_6621,N_5961,N_1382);
and U6622 (N_6622,N_4411,N_2384);
and U6623 (N_6623,N_359,N_1110);
nand U6624 (N_6624,N_5086,N_5729);
or U6625 (N_6625,N_5275,N_6028);
nor U6626 (N_6626,N_5082,N_1517);
or U6627 (N_6627,N_3229,N_499);
xnor U6628 (N_6628,N_5997,N_619);
or U6629 (N_6629,N_2797,N_4903);
nor U6630 (N_6630,N_1542,N_5507);
nor U6631 (N_6631,N_163,N_691);
nor U6632 (N_6632,N_5349,N_1667);
nor U6633 (N_6633,N_1994,N_3946);
and U6634 (N_6634,N_253,N_1670);
and U6635 (N_6635,N_439,N_2478);
nor U6636 (N_6636,N_3749,N_5050);
xor U6637 (N_6637,N_876,N_4687);
and U6638 (N_6638,N_6193,N_3892);
and U6639 (N_6639,N_5662,N_2209);
nor U6640 (N_6640,N_4422,N_3820);
xnor U6641 (N_6641,N_2868,N_4615);
nand U6642 (N_6642,N_4859,N_1368);
nand U6643 (N_6643,N_5770,N_6096);
nor U6644 (N_6644,N_6066,N_5120);
or U6645 (N_6645,N_4980,N_3430);
xnor U6646 (N_6646,N_4483,N_2380);
nor U6647 (N_6647,N_2250,N_5115);
nand U6648 (N_6648,N_3373,N_2088);
nor U6649 (N_6649,N_1734,N_4081);
or U6650 (N_6650,N_6153,N_6025);
xnor U6651 (N_6651,N_5637,N_1704);
nor U6652 (N_6652,N_1275,N_388);
and U6653 (N_6653,N_4424,N_4589);
or U6654 (N_6654,N_2137,N_2397);
and U6655 (N_6655,N_2645,N_3368);
or U6656 (N_6656,N_1828,N_5277);
or U6657 (N_6657,N_235,N_2215);
nand U6658 (N_6658,N_298,N_5955);
nand U6659 (N_6659,N_3619,N_4307);
nor U6660 (N_6660,N_4183,N_1361);
xnor U6661 (N_6661,N_1679,N_5070);
or U6662 (N_6662,N_2876,N_4438);
nand U6663 (N_6663,N_3981,N_5741);
nand U6664 (N_6664,N_4244,N_3797);
xor U6665 (N_6665,N_2960,N_3663);
nand U6666 (N_6666,N_655,N_225);
or U6667 (N_6667,N_4159,N_2949);
and U6668 (N_6668,N_446,N_1224);
and U6669 (N_6669,N_2679,N_1348);
and U6670 (N_6670,N_3702,N_4806);
xnor U6671 (N_6671,N_102,N_1352);
or U6672 (N_6672,N_4930,N_4194);
or U6673 (N_6673,N_6052,N_4463);
or U6674 (N_6674,N_3474,N_585);
nand U6675 (N_6675,N_5330,N_942);
and U6676 (N_6676,N_36,N_581);
xnor U6677 (N_6677,N_3148,N_125);
xor U6678 (N_6678,N_1161,N_690);
and U6679 (N_6679,N_887,N_1919);
nor U6680 (N_6680,N_4292,N_5407);
nor U6681 (N_6681,N_632,N_5759);
or U6682 (N_6682,N_3355,N_5272);
xnor U6683 (N_6683,N_1587,N_2127);
nor U6684 (N_6684,N_2779,N_323);
and U6685 (N_6685,N_2401,N_4223);
nor U6686 (N_6686,N_1811,N_297);
nand U6687 (N_6687,N_4978,N_1304);
nand U6688 (N_6688,N_3499,N_2266);
nand U6689 (N_6689,N_206,N_4802);
nand U6690 (N_6690,N_867,N_2388);
nand U6691 (N_6691,N_4418,N_1231);
xnor U6692 (N_6692,N_4908,N_2048);
or U6693 (N_6693,N_4295,N_4432);
nor U6694 (N_6694,N_4782,N_948);
and U6695 (N_6695,N_6002,N_4719);
xnor U6696 (N_6696,N_433,N_6192);
and U6697 (N_6697,N_5460,N_4439);
and U6698 (N_6698,N_2545,N_2385);
and U6699 (N_6699,N_4702,N_849);
and U6700 (N_6700,N_2996,N_4798);
nand U6701 (N_6701,N_1748,N_4191);
nand U6702 (N_6702,N_5378,N_1849);
nor U6703 (N_6703,N_5340,N_5919);
and U6704 (N_6704,N_4797,N_1480);
nand U6705 (N_6705,N_2951,N_5984);
xnor U6706 (N_6706,N_6001,N_3174);
xnor U6707 (N_6707,N_1952,N_1292);
nor U6708 (N_6708,N_92,N_1785);
nand U6709 (N_6709,N_4313,N_3666);
nand U6710 (N_6710,N_5999,N_2967);
or U6711 (N_6711,N_3503,N_3530);
or U6712 (N_6712,N_1049,N_4017);
nor U6713 (N_6713,N_2389,N_932);
and U6714 (N_6714,N_3613,N_561);
xnor U6715 (N_6715,N_2616,N_4467);
or U6716 (N_6716,N_3603,N_374);
nand U6717 (N_6717,N_834,N_4013);
and U6718 (N_6718,N_946,N_4684);
nand U6719 (N_6719,N_355,N_4904);
and U6720 (N_6720,N_441,N_5035);
nor U6721 (N_6721,N_4545,N_3044);
nand U6722 (N_6722,N_4534,N_6190);
xor U6723 (N_6723,N_1313,N_6069);
or U6724 (N_6724,N_5692,N_4869);
nor U6725 (N_6725,N_6099,N_2543);
nand U6726 (N_6726,N_4459,N_1029);
nand U6727 (N_6727,N_4565,N_5145);
xnor U6728 (N_6728,N_5941,N_5201);
xor U6729 (N_6729,N_3594,N_4367);
xnor U6730 (N_6730,N_5172,N_3644);
and U6731 (N_6731,N_2647,N_3408);
or U6732 (N_6732,N_4861,N_1946);
nor U6733 (N_6733,N_1892,N_4656);
and U6734 (N_6734,N_3874,N_1477);
nand U6735 (N_6735,N_997,N_5975);
nand U6736 (N_6736,N_5610,N_3232);
nand U6737 (N_6737,N_5787,N_4096);
xor U6738 (N_6738,N_5016,N_5234);
nand U6739 (N_6739,N_5079,N_1977);
nor U6740 (N_6740,N_2318,N_1180);
nor U6741 (N_6741,N_1744,N_2711);
and U6742 (N_6742,N_1898,N_4587);
nand U6743 (N_6743,N_1685,N_4549);
nand U6744 (N_6744,N_4140,N_2256);
or U6745 (N_6745,N_5325,N_3894);
nor U6746 (N_6746,N_2693,N_3621);
xor U6747 (N_6747,N_3432,N_3692);
and U6748 (N_6748,N_3816,N_2508);
or U6749 (N_6749,N_2504,N_5736);
or U6750 (N_6750,N_308,N_4774);
nand U6751 (N_6751,N_418,N_4015);
nand U6752 (N_6752,N_2562,N_1516);
nand U6753 (N_6753,N_531,N_1150);
nand U6754 (N_6754,N_1708,N_2611);
xor U6755 (N_6755,N_2124,N_5939);
or U6756 (N_6756,N_2114,N_3451);
nand U6757 (N_6757,N_1630,N_3719);
or U6758 (N_6758,N_5575,N_390);
nand U6759 (N_6759,N_840,N_6163);
and U6760 (N_6760,N_4714,N_3151);
xnor U6761 (N_6761,N_4648,N_3112);
xor U6762 (N_6762,N_5229,N_2754);
nand U6763 (N_6763,N_506,N_1108);
nand U6764 (N_6764,N_1495,N_6220);
xor U6765 (N_6765,N_3276,N_1398);
nor U6766 (N_6766,N_1321,N_1739);
xor U6767 (N_6767,N_1479,N_1573);
and U6768 (N_6768,N_1414,N_5651);
and U6769 (N_6769,N_3852,N_2682);
or U6770 (N_6770,N_4956,N_4065);
nand U6771 (N_6771,N_267,N_3482);
or U6772 (N_6772,N_716,N_2120);
xor U6773 (N_6773,N_1432,N_5732);
xor U6774 (N_6774,N_662,N_5945);
xor U6775 (N_6775,N_58,N_1862);
nand U6776 (N_6776,N_2507,N_4917);
nand U6777 (N_6777,N_1856,N_1683);
nand U6778 (N_6778,N_6199,N_2660);
nand U6779 (N_6779,N_5113,N_57);
nor U6780 (N_6780,N_957,N_559);
and U6781 (N_6781,N_4068,N_679);
and U6782 (N_6782,N_6188,N_2920);
and U6783 (N_6783,N_2617,N_883);
nand U6784 (N_6784,N_1081,N_1973);
or U6785 (N_6785,N_1301,N_1962);
nor U6786 (N_6786,N_3189,N_4723);
xnor U6787 (N_6787,N_4588,N_4844);
nor U6788 (N_6788,N_4996,N_3800);
or U6789 (N_6789,N_4755,N_1752);
xor U6790 (N_6790,N_3955,N_3602);
or U6791 (N_6791,N_2802,N_2948);
nand U6792 (N_6792,N_5635,N_1251);
nor U6793 (N_6793,N_2156,N_1172);
nor U6794 (N_6794,N_3339,N_5419);
xnor U6795 (N_6795,N_6133,N_5788);
xor U6796 (N_6796,N_853,N_2678);
nor U6797 (N_6797,N_2080,N_202);
xor U6798 (N_6798,N_5509,N_674);
nor U6799 (N_6799,N_647,N_5047);
xor U6800 (N_6800,N_4591,N_3099);
nand U6801 (N_6801,N_340,N_4654);
or U6802 (N_6802,N_5646,N_3915);
or U6803 (N_6803,N_919,N_3690);
nor U6804 (N_6804,N_4877,N_659);
nand U6805 (N_6805,N_480,N_2629);
nand U6806 (N_6806,N_1032,N_627);
nor U6807 (N_6807,N_4163,N_1766);
xor U6808 (N_6808,N_6166,N_4809);
and U6809 (N_6809,N_5562,N_4128);
nand U6810 (N_6810,N_1487,N_1850);
and U6811 (N_6811,N_6055,N_1887);
nand U6812 (N_6812,N_787,N_4960);
nor U6813 (N_6813,N_5026,N_2175);
xor U6814 (N_6814,N_2929,N_232);
or U6815 (N_6815,N_4965,N_658);
nor U6816 (N_6816,N_666,N_2149);
or U6817 (N_6817,N_3937,N_4758);
xnor U6818 (N_6818,N_3896,N_6129);
nor U6819 (N_6819,N_1738,N_2406);
nand U6820 (N_6820,N_2201,N_3192);
nor U6821 (N_6821,N_3776,N_5221);
xnor U6822 (N_6822,N_205,N_2276);
or U6823 (N_6823,N_4590,N_5544);
nor U6824 (N_6824,N_2816,N_5475);
or U6825 (N_6825,N_792,N_3383);
or U6826 (N_6826,N_6160,N_3555);
nor U6827 (N_6827,N_4646,N_3028);
nand U6828 (N_6828,N_881,N_830);
or U6829 (N_6829,N_41,N_1427);
or U6830 (N_6830,N_1724,N_1363);
xnor U6831 (N_6831,N_5179,N_2155);
xor U6832 (N_6832,N_6232,N_5036);
xor U6833 (N_6833,N_2067,N_2382);
xnor U6834 (N_6834,N_4767,N_4526);
and U6835 (N_6835,N_4914,N_2702);
nand U6836 (N_6836,N_353,N_6223);
xnor U6837 (N_6837,N_3799,N_2564);
xnor U6838 (N_6838,N_5811,N_2495);
or U6839 (N_6839,N_2446,N_279);
and U6840 (N_6840,N_2935,N_99);
and U6841 (N_6841,N_5186,N_5345);
xnor U6842 (N_6842,N_312,N_3040);
xnor U6843 (N_6843,N_157,N_1909);
or U6844 (N_6844,N_5487,N_244);
nand U6845 (N_6845,N_2152,N_1241);
nor U6846 (N_6846,N_2190,N_1459);
nor U6847 (N_6847,N_5220,N_5907);
nand U6848 (N_6848,N_2001,N_3072);
and U6849 (N_6849,N_780,N_6011);
nand U6850 (N_6850,N_423,N_2198);
and U6851 (N_6851,N_4668,N_1772);
xnor U6852 (N_6852,N_3558,N_387);
xor U6853 (N_6853,N_3532,N_2815);
or U6854 (N_6854,N_3133,N_5301);
nor U6855 (N_6855,N_5080,N_3406);
xor U6856 (N_6856,N_4658,N_4799);
nor U6857 (N_6857,N_5881,N_2530);
or U6858 (N_6858,N_4036,N_1132);
or U6859 (N_6859,N_719,N_4118);
nor U6860 (N_6860,N_3583,N_3280);
xnor U6861 (N_6861,N_1669,N_2281);
xor U6862 (N_6862,N_497,N_3803);
nor U6863 (N_6863,N_220,N_2375);
nor U6864 (N_6864,N_3,N_4726);
xnor U6865 (N_6865,N_3016,N_1591);
or U6866 (N_6866,N_1246,N_2301);
nand U6867 (N_6867,N_995,N_124);
and U6868 (N_6868,N_4287,N_2761);
or U6869 (N_6869,N_5152,N_4553);
xnor U6870 (N_6870,N_4444,N_1116);
or U6871 (N_6871,N_3285,N_3030);
nand U6872 (N_6872,N_5485,N_4088);
or U6873 (N_6873,N_180,N_1563);
and U6874 (N_6874,N_2857,N_4107);
and U6875 (N_6875,N_6161,N_5521);
and U6876 (N_6876,N_2873,N_1700);
or U6877 (N_6877,N_1259,N_4950);
and U6878 (N_6878,N_5554,N_520);
nand U6879 (N_6879,N_1435,N_2216);
and U6880 (N_6880,N_4097,N_5081);
or U6881 (N_6881,N_5748,N_1468);
and U6882 (N_6882,N_6183,N_3172);
and U6883 (N_6883,N_5392,N_964);
nand U6884 (N_6884,N_4880,N_5307);
or U6885 (N_6885,N_4510,N_113);
or U6886 (N_6886,N_4446,N_5461);
xor U6887 (N_6887,N_1899,N_2942);
nor U6888 (N_6888,N_3225,N_6184);
nand U6889 (N_6889,N_5441,N_1215);
or U6890 (N_6890,N_5083,N_5243);
nand U6891 (N_6891,N_4681,N_4354);
nand U6892 (N_6892,N_5923,N_4532);
and U6893 (N_6893,N_4117,N_5926);
or U6894 (N_6894,N_3652,N_6179);
nand U6895 (N_6895,N_4923,N_583);
or U6896 (N_6896,N_2810,N_2601);
and U6897 (N_6897,N_4445,N_2771);
nand U6898 (N_6898,N_5060,N_3018);
or U6899 (N_6899,N_4795,N_3854);
or U6900 (N_6900,N_1113,N_3650);
and U6901 (N_6901,N_908,N_5699);
nand U6902 (N_6902,N_3160,N_452);
xnor U6903 (N_6903,N_3813,N_3060);
nand U6904 (N_6904,N_4805,N_5426);
xnor U6905 (N_6905,N_105,N_4193);
or U6906 (N_6906,N_3258,N_516);
xor U6907 (N_6907,N_4902,N_579);
nand U6908 (N_6908,N_3359,N_1750);
nor U6909 (N_6909,N_3518,N_4387);
nor U6910 (N_6910,N_3457,N_174);
nor U6911 (N_6911,N_4360,N_4357);
and U6912 (N_6912,N_5824,N_2514);
and U6913 (N_6913,N_1263,N_1176);
nand U6914 (N_6914,N_2070,N_5684);
or U6915 (N_6915,N_1701,N_5796);
or U6916 (N_6916,N_4607,N_5596);
and U6917 (N_6917,N_2987,N_2903);
nand U6918 (N_6918,N_2122,N_1054);
or U6919 (N_6919,N_73,N_3920);
nor U6920 (N_6920,N_5847,N_636);
nand U6921 (N_6921,N_5896,N_1570);
nand U6922 (N_6922,N_855,N_4161);
nand U6923 (N_6923,N_4729,N_5952);
nand U6924 (N_6924,N_3207,N_1721);
nand U6925 (N_6925,N_3141,N_302);
nor U6926 (N_6926,N_996,N_1062);
and U6927 (N_6927,N_5333,N_3615);
xnor U6928 (N_6928,N_2062,N_20);
and U6929 (N_6929,N_5943,N_3591);
and U6930 (N_6930,N_168,N_3837);
nor U6931 (N_6931,N_1853,N_291);
or U6932 (N_6932,N_5682,N_3642);
and U6933 (N_6933,N_4621,N_3278);
nor U6934 (N_6934,N_177,N_4399);
or U6935 (N_6935,N_5482,N_4139);
nor U6936 (N_6936,N_6063,N_1373);
nor U6937 (N_6937,N_5281,N_5278);
xnor U6938 (N_6938,N_1656,N_2829);
or U6939 (N_6939,N_3960,N_5920);
xor U6940 (N_6940,N_535,N_1770);
or U6941 (N_6941,N_2565,N_2213);
xor U6942 (N_6942,N_589,N_181);
nor U6943 (N_6943,N_3497,N_1377);
or U6944 (N_6944,N_5523,N_4576);
xnor U6945 (N_6945,N_2079,N_2773);
nor U6946 (N_6946,N_4067,N_1733);
xor U6947 (N_6947,N_4455,N_5413);
nor U6948 (N_6948,N_3542,N_5191);
nand U6949 (N_6949,N_1904,N_5252);
xnor U6950 (N_6950,N_4484,N_759);
nand U6951 (N_6951,N_6078,N_2999);
xor U6952 (N_6952,N_1598,N_5620);
nor U6953 (N_6953,N_1034,N_436);
and U6954 (N_6954,N_1960,N_1210);
or U6955 (N_6955,N_1126,N_3640);
and U6956 (N_6956,N_5954,N_391);
or U6957 (N_6957,N_3829,N_5395);
xnor U6958 (N_6958,N_2426,N_4392);
or U6959 (N_6959,N_305,N_5052);
nand U6960 (N_6960,N_1918,N_467);
and U6961 (N_6961,N_599,N_3294);
nand U6962 (N_6962,N_3941,N_324);
or U6963 (N_6963,N_3687,N_1383);
nor U6964 (N_6964,N_1417,N_5644);
or U6965 (N_6965,N_5098,N_4944);
or U6966 (N_6966,N_1827,N_963);
and U6967 (N_6967,N_4240,N_1128);
and U6968 (N_6968,N_1732,N_4162);
and U6969 (N_6969,N_1339,N_4016);
or U6970 (N_6970,N_3608,N_4456);
xor U6971 (N_6971,N_5490,N_3220);
or U6972 (N_6972,N_3400,N_961);
xnor U6973 (N_6973,N_462,N_5343);
or U6974 (N_6974,N_5473,N_2671);
nand U6975 (N_6975,N_5341,N_657);
or U6976 (N_6976,N_4744,N_4958);
nor U6977 (N_6977,N_6013,N_4867);
and U6978 (N_6978,N_2060,N_2612);
or U6979 (N_6979,N_4103,N_1244);
or U6980 (N_6980,N_427,N_95);
or U6981 (N_6981,N_4539,N_2394);
and U6982 (N_6982,N_3113,N_1327);
xor U6983 (N_6983,N_5893,N_2864);
and U6984 (N_6984,N_4523,N_4820);
nand U6985 (N_6985,N_5779,N_385);
or U6986 (N_6986,N_1520,N_3864);
xnor U6987 (N_6987,N_929,N_4593);
nand U6988 (N_6988,N_573,N_5743);
nand U6989 (N_6989,N_5359,N_4524);
nand U6990 (N_6990,N_1175,N_3165);
and U6991 (N_6991,N_4394,N_6128);
nor U6992 (N_6992,N_218,N_6106);
or U6993 (N_6993,N_4731,N_5851);
nor U6994 (N_6994,N_419,N_770);
or U6995 (N_6995,N_1810,N_4538);
nor U6996 (N_6996,N_5382,N_4109);
and U6997 (N_6997,N_1813,N_3020);
and U6998 (N_6998,N_5717,N_2073);
or U6999 (N_6999,N_5369,N_1900);
or U7000 (N_7000,N_3277,N_3401);
and U7001 (N_7001,N_3638,N_3354);
and U7002 (N_7002,N_4789,N_1965);
xor U7003 (N_7003,N_2986,N_2763);
xor U7004 (N_7004,N_5001,N_4281);
nand U7005 (N_7005,N_2634,N_2578);
and U7006 (N_7006,N_4769,N_1430);
or U7007 (N_7007,N_4941,N_2805);
xor U7008 (N_7008,N_2368,N_4918);
nor U7009 (N_7009,N_5027,N_3504);
and U7010 (N_7010,N_3202,N_4989);
or U7011 (N_7011,N_5948,N_5045);
or U7012 (N_7012,N_5074,N_4447);
xor U7013 (N_7013,N_2900,N_6100);
and U7014 (N_7014,N_1974,N_847);
xnor U7015 (N_7015,N_5142,N_5664);
nand U7016 (N_7016,N_2746,N_4453);
nand U7017 (N_7017,N_1336,N_2934);
or U7018 (N_7018,N_5383,N_6201);
or U7019 (N_7019,N_1501,N_4651);
nor U7020 (N_7020,N_4053,N_546);
nor U7021 (N_7021,N_3259,N_5262);
or U7022 (N_7022,N_14,N_4204);
nor U7023 (N_7023,N_1753,N_2944);
and U7024 (N_7024,N_3091,N_2780);
and U7025 (N_7025,N_1681,N_2845);
nor U7026 (N_7026,N_5305,N_1801);
and U7027 (N_7027,N_1015,N_5236);
and U7028 (N_7028,N_6114,N_3335);
nand U7029 (N_7029,N_629,N_5335);
nand U7030 (N_7030,N_1121,N_5273);
or U7031 (N_7031,N_1025,N_3805);
xnor U7032 (N_7032,N_3807,N_2355);
nor U7033 (N_7033,N_5938,N_3616);
nor U7034 (N_7034,N_5512,N_5078);
xnor U7035 (N_7035,N_5462,N_724);
xor U7036 (N_7036,N_5889,N_149);
nor U7037 (N_7037,N_4406,N_1388);
nor U7038 (N_7038,N_2072,N_5421);
xor U7039 (N_7039,N_5616,N_5265);
nor U7040 (N_7040,N_238,N_931);
or U7041 (N_7041,N_4404,N_6217);
nor U7042 (N_7042,N_5607,N_844);
nor U7043 (N_7043,N_221,N_2163);
nand U7044 (N_7044,N_5622,N_2625);
nor U7045 (N_7045,N_1655,N_5185);
nor U7046 (N_7046,N_3352,N_5464);
nor U7047 (N_7047,N_71,N_3902);
nand U7048 (N_7048,N_2316,N_5527);
or U7049 (N_7049,N_5247,N_3840);
xnor U7050 (N_7050,N_5643,N_4316);
or U7051 (N_7051,N_2442,N_1500);
nor U7052 (N_7052,N_3535,N_2640);
or U7053 (N_7053,N_1258,N_4529);
and U7054 (N_7054,N_4202,N_4084);
nor U7055 (N_7055,N_5547,N_744);
nor U7056 (N_7056,N_1792,N_2219);
nand U7057 (N_7057,N_1011,N_2861);
nand U7058 (N_7058,N_5883,N_652);
or U7059 (N_7059,N_2195,N_2044);
and U7060 (N_7060,N_4982,N_3789);
or U7061 (N_7061,N_5066,N_3551);
nand U7062 (N_7062,N_1229,N_4559);
xnor U7063 (N_7063,N_47,N_733);
nand U7064 (N_7064,N_2836,N_3098);
nor U7065 (N_7065,N_2624,N_1370);
xnor U7066 (N_7066,N_1868,N_3298);
and U7067 (N_7067,N_1934,N_331);
and U7068 (N_7068,N_5552,N_2520);
nand U7069 (N_7069,N_3819,N_2186);
nor U7070 (N_7070,N_819,N_3319);
nand U7071 (N_7071,N_2729,N_3063);
or U7072 (N_7072,N_4352,N_5707);
nor U7073 (N_7073,N_4341,N_3956);
nor U7074 (N_7074,N_3520,N_5119);
nor U7075 (N_7075,N_1858,N_2874);
or U7076 (N_7076,N_4386,N_3887);
xor U7077 (N_7077,N_3450,N_409);
or U7078 (N_7078,N_3814,N_607);
or U7079 (N_7079,N_892,N_411);
or U7080 (N_7080,N_1607,N_4243);
or U7081 (N_7081,N_5738,N_1179);
nand U7082 (N_7082,N_5902,N_5364);
nor U7083 (N_7083,N_3635,N_2794);
nor U7084 (N_7084,N_3435,N_4949);
and U7085 (N_7085,N_2649,N_6244);
and U7086 (N_7086,N_6097,N_3978);
or U7087 (N_7087,N_2400,N_2126);
nor U7088 (N_7088,N_5000,N_2686);
and U7089 (N_7089,N_2220,N_5495);
xor U7090 (N_7090,N_1485,N_1160);
or U7091 (N_7091,N_3788,N_1759);
or U7092 (N_7092,N_1079,N_1941);
nor U7093 (N_7093,N_3938,N_3005);
and U7094 (N_7094,N_4976,N_3756);
nand U7095 (N_7095,N_4649,N_5762);
or U7096 (N_7096,N_2681,N_4076);
and U7097 (N_7097,N_3773,N_2091);
nand U7098 (N_7098,N_1021,N_6016);
nand U7099 (N_7099,N_5795,N_4911);
xor U7100 (N_7100,N_4892,N_1186);
nor U7101 (N_7101,N_1234,N_2026);
xor U7102 (N_7102,N_3349,N_1581);
or U7103 (N_7103,N_739,N_40);
and U7104 (N_7104,N_2991,N_5807);
nand U7105 (N_7105,N_672,N_5287);
or U7106 (N_7106,N_5733,N_259);
nand U7107 (N_7107,N_1117,N_2710);
and U7108 (N_7108,N_5673,N_5887);
and U7109 (N_7109,N_5794,N_3881);
or U7110 (N_7110,N_1375,N_3397);
nor U7111 (N_7111,N_4558,N_4878);
xor U7112 (N_7112,N_4919,N_1271);
nor U7113 (N_7113,N_332,N_735);
and U7114 (N_7114,N_2012,N_3730);
and U7115 (N_7115,N_596,N_333);
or U7116 (N_7116,N_5618,N_2292);
nand U7117 (N_7117,N_4764,N_1575);
nor U7118 (N_7118,N_2343,N_3391);
nor U7119 (N_7119,N_3061,N_5854);
or U7120 (N_7120,N_1536,N_3625);
nor U7121 (N_7121,N_3631,N_4388);
nand U7122 (N_7122,N_2533,N_3958);
and U7123 (N_7123,N_2259,N_2567);
nand U7124 (N_7124,N_858,N_1914);
nand U7125 (N_7125,N_1014,N_4461);
xnor U7126 (N_7126,N_1426,N_1197);
and U7127 (N_7127,N_2842,N_1264);
nand U7128 (N_7128,N_5471,N_1547);
xor U7129 (N_7129,N_5790,N_1963);
or U7130 (N_7130,N_4051,N_5202);
nor U7131 (N_7131,N_993,N_5519);
nor U7132 (N_7132,N_4336,N_2458);
xnor U7133 (N_7133,N_4567,N_4138);
or U7134 (N_7134,N_88,N_3472);
or U7135 (N_7135,N_1825,N_445);
and U7136 (N_7136,N_5192,N_3522);
nor U7137 (N_7137,N_661,N_5321);
xnor U7138 (N_7138,N_2814,N_4898);
nor U7139 (N_7139,N_2045,N_4008);
and U7140 (N_7140,N_5853,N_1360);
xnor U7141 (N_7141,N_3088,N_4382);
or U7142 (N_7142,N_4736,N_626);
xor U7143 (N_7143,N_2354,N_3538);
nand U7144 (N_7144,N_6240,N_4620);
or U7145 (N_7145,N_5866,N_4662);
nand U7146 (N_7146,N_2882,N_3612);
or U7147 (N_7147,N_4741,N_5496);
nor U7148 (N_7148,N_5508,N_2274);
nor U7149 (N_7149,N_5127,N_5018);
nand U7150 (N_7150,N_3846,N_3664);
xor U7151 (N_7151,N_1455,N_2428);
nand U7152 (N_7152,N_3283,N_2859);
nor U7153 (N_7153,N_5055,N_87);
nand U7154 (N_7154,N_2136,N_2888);
and U7155 (N_7155,N_3102,N_1999);
nand U7156 (N_7156,N_4959,N_4210);
nand U7157 (N_7157,N_1256,N_2092);
or U7158 (N_7158,N_2020,N_1933);
or U7159 (N_7159,N_6222,N_219);
or U7160 (N_7160,N_843,N_3264);
or U7161 (N_7161,N_3004,N_1959);
nand U7162 (N_7162,N_5025,N_2572);
nor U7163 (N_7163,N_3011,N_6126);
and U7164 (N_7164,N_3154,N_4934);
xnor U7165 (N_7165,N_1429,N_5675);
and U7166 (N_7166,N_4585,N_4427);
nand U7167 (N_7167,N_5132,N_2807);
nor U7168 (N_7168,N_2855,N_4258);
or U7169 (N_7169,N_1439,N_3826);
or U7170 (N_7170,N_5367,N_1216);
and U7171 (N_7171,N_2883,N_4324);
or U7172 (N_7172,N_352,N_638);
nand U7173 (N_7173,N_4754,N_2110);
nor U7174 (N_7174,N_1071,N_2837);
nor U7175 (N_7175,N_757,N_5169);
or U7176 (N_7176,N_4482,N_342);
nand U7177 (N_7177,N_4768,N_5751);
nor U7178 (N_7178,N_886,N_5443);
and U7179 (N_7179,N_4599,N_2800);
xnor U7180 (N_7180,N_320,N_170);
or U7181 (N_7181,N_3089,N_2303);
nand U7182 (N_7182,N_3317,N_3201);
and U7183 (N_7183,N_1836,N_2922);
xnor U7184 (N_7184,N_2466,N_6023);
xor U7185 (N_7185,N_4555,N_5640);
xnor U7186 (N_7186,N_289,N_5870);
xor U7187 (N_7187,N_4751,N_682);
and U7188 (N_7188,N_5437,N_5877);
nand U7189 (N_7189,N_5256,N_4564);
nor U7190 (N_7190,N_6045,N_2396);
and U7191 (N_7191,N_2526,N_6020);
nand U7192 (N_7192,N_5995,N_2963);
and U7193 (N_7193,N_1553,N_1561);
and U7194 (N_7194,N_1324,N_4454);
xor U7195 (N_7195,N_5534,N_937);
nor U7196 (N_7196,N_3665,N_3968);
and U7197 (N_7197,N_3985,N_1389);
or U7198 (N_7198,N_2984,N_4957);
nand U7199 (N_7199,N_5068,N_5123);
xor U7200 (N_7200,N_4169,N_488);
nand U7201 (N_7201,N_4166,N_89);
and U7202 (N_7202,N_5261,N_2579);
and U7203 (N_7203,N_1428,N_294);
nand U7204 (N_7204,N_3828,N_2894);
or U7205 (N_7205,N_746,N_921);
and U7206 (N_7206,N_2840,N_5100);
or U7207 (N_7207,N_1498,N_4745);
or U7208 (N_7208,N_5008,N_5284);
and U7209 (N_7209,N_947,N_3167);
xnor U7210 (N_7210,N_1247,N_2534);
nor U7211 (N_7211,N_991,N_1308);
xnor U7212 (N_7212,N_4188,N_2619);
nor U7213 (N_7213,N_3272,N_3215);
or U7214 (N_7214,N_269,N_5558);
nand U7215 (N_7215,N_5809,N_1319);
nor U7216 (N_7216,N_6168,N_2901);
or U7217 (N_7217,N_4353,N_4512);
nand U7218 (N_7218,N_3867,N_2972);
nor U7219 (N_7219,N_2643,N_1237);
and U7220 (N_7220,N_530,N_1539);
nand U7221 (N_7221,N_4112,N_3117);
xnor U7222 (N_7222,N_2221,N_3812);
nor U7223 (N_7223,N_2809,N_3751);
nand U7224 (N_7224,N_5194,N_5960);
xnor U7225 (N_7225,N_5656,N_3618);
nor U7226 (N_7226,N_582,N_3302);
xor U7227 (N_7227,N_1090,N_376);
xor U7228 (N_7228,N_3153,N_3722);
nor U7229 (N_7229,N_5310,N_5800);
xor U7230 (N_7230,N_2130,N_2189);
nor U7231 (N_7231,N_3162,N_53);
xnor U7232 (N_7232,N_857,N_5597);
and U7233 (N_7233,N_4855,N_4475);
and U7234 (N_7234,N_3290,N_3027);
and U7235 (N_7235,N_778,N_4866);
xnor U7236 (N_7236,N_2978,N_5294);
and U7237 (N_7237,N_3975,N_1557);
or U7238 (N_7238,N_2359,N_1746);
and U7239 (N_7239,N_3096,N_2713);
nand U7240 (N_7240,N_6147,N_222);
or U7241 (N_7241,N_5015,N_5468);
xor U7242 (N_7242,N_5579,N_406);
nor U7243 (N_7243,N_916,N_4369);
nor U7244 (N_7244,N_303,N_408);
nand U7245 (N_7245,N_3263,N_1996);
nand U7246 (N_7246,N_2801,N_1005);
nand U7247 (N_7247,N_17,N_1751);
and U7248 (N_7248,N_6000,N_1092);
or U7249 (N_7249,N_4127,N_2788);
nand U7250 (N_7250,N_4592,N_59);
nand U7251 (N_7251,N_1796,N_4671);
nand U7252 (N_7252,N_3516,N_2571);
or U7253 (N_7253,N_2464,N_4794);
xor U7254 (N_7254,N_5603,N_3466);
and U7255 (N_7255,N_549,N_3916);
and U7256 (N_7256,N_2657,N_2000);
nand U7257 (N_7257,N_2735,N_3394);
xnor U7258 (N_7258,N_2953,N_5826);
or U7259 (N_7259,N_3835,N_902);
nor U7260 (N_7260,N_54,N_2932);
and U7261 (N_7261,N_6191,N_5722);
or U7262 (N_7262,N_4999,N_4920);
nand U7263 (N_7263,N_5013,N_2214);
nor U7264 (N_7264,N_3017,N_956);
nand U7265 (N_7265,N_4577,N_4014);
xnor U7266 (N_7266,N_4685,N_4594);
or U7267 (N_7267,N_1876,N_978);
and U7268 (N_7268,N_2381,N_6156);
or U7269 (N_7269,N_2411,N_2650);
nand U7270 (N_7270,N_3706,N_3745);
nor U7271 (N_7271,N_6158,N_5159);
nor U7272 (N_7272,N_5702,N_4962);
xnor U7273 (N_7273,N_42,N_1555);
nor U7274 (N_7274,N_37,N_6064);
nand U7275 (N_7275,N_1694,N_5255);
nand U7276 (N_7276,N_1891,N_1395);
or U7277 (N_7277,N_4426,N_5312);
xnor U7278 (N_7278,N_46,N_166);
nor U7279 (N_7279,N_1196,N_5884);
nor U7280 (N_7280,N_3300,N_3158);
nor U7281 (N_7281,N_2097,N_1280);
or U7282 (N_7282,N_3626,N_3114);
and U7283 (N_7283,N_5761,N_3505);
nand U7284 (N_7284,N_3711,N_2687);
and U7285 (N_7285,N_5658,N_434);
nor U7286 (N_7286,N_4358,N_1065);
and U7287 (N_7287,N_3934,N_3159);
or U7288 (N_7288,N_1416,N_3053);
xnor U7289 (N_7289,N_1958,N_3903);
or U7290 (N_7290,N_3152,N_310);
xnor U7291 (N_7291,N_2095,N_2558);
nand U7292 (N_7292,N_5555,N_2423);
and U7293 (N_7293,N_1144,N_368);
nor U7294 (N_7294,N_421,N_5559);
or U7295 (N_7295,N_4317,N_4985);
nand U7296 (N_7296,N_1794,N_1783);
and U7297 (N_7297,N_577,N_6057);
or U7298 (N_7298,N_4170,N_2577);
xnor U7299 (N_7299,N_2586,N_4042);
nor U7300 (N_7300,N_3748,N_4544);
nor U7301 (N_7301,N_3834,N_4875);
nor U7302 (N_7302,N_4314,N_4421);
and U7303 (N_7303,N_3356,N_2480);
nor U7304 (N_7304,N_2444,N_198);
xor U7305 (N_7305,N_3766,N_5320);
xnor U7306 (N_7306,N_2714,N_2115);
nor U7307 (N_7307,N_2013,N_6221);
nor U7308 (N_7308,N_83,N_2684);
xor U7309 (N_7309,N_5427,N_1061);
nand U7310 (N_7310,N_1445,N_3342);
xnor U7311 (N_7311,N_5792,N_4891);
nand U7312 (N_7312,N_3299,N_5248);
or U7313 (N_7313,N_4309,N_5869);
nand U7314 (N_7314,N_3262,N_139);
nand U7315 (N_7315,N_5266,N_151);
nand U7316 (N_7316,N_1273,N_1985);
nand U7317 (N_7317,N_6046,N_3524);
or U7318 (N_7318,N_4826,N_2069);
nand U7319 (N_7319,N_3912,N_1756);
nor U7320 (N_7320,N_1951,N_2856);
nand U7321 (N_7321,N_5213,N_2153);
xor U7322 (N_7322,N_1728,N_1926);
xor U7323 (N_7323,N_763,N_960);
or U7324 (N_7324,N_112,N_1020);
nor U7325 (N_7325,N_6245,N_741);
xnor U7326 (N_7326,N_5797,N_6085);
or U7327 (N_7327,N_4643,N_2789);
xor U7328 (N_7328,N_5844,N_3743);
nor U7329 (N_7329,N_3701,N_6177);
or U7330 (N_7330,N_2358,N_4003);
xnor U7331 (N_7331,N_3344,N_3436);
and U7332 (N_7332,N_2116,N_3191);
xor U7333 (N_7333,N_137,N_1306);
or U7334 (N_7334,N_2704,N_4616);
or U7335 (N_7335,N_3703,N_1290);
xnor U7336 (N_7336,N_476,N_6150);
or U7337 (N_7337,N_3001,N_4948);
xor U7338 (N_7338,N_1627,N_478);
nand U7339 (N_7339,N_3909,N_5104);
xor U7340 (N_7340,N_3054,N_4677);
nand U7341 (N_7341,N_4813,N_4361);
nor U7342 (N_7342,N_4040,N_6053);
nor U7343 (N_7343,N_3669,N_4974);
or U7344 (N_7344,N_6241,N_4873);
nand U7345 (N_7345,N_4277,N_1719);
xor U7346 (N_7346,N_493,N_5388);
nor U7347 (N_7347,N_3693,N_4846);
nand U7348 (N_7348,N_3895,N_2192);
xnor U7349 (N_7349,N_2171,N_615);
and U7350 (N_7350,N_775,N_4435);
xnor U7351 (N_7351,N_1478,N_4951);
nand U7352 (N_7352,N_4372,N_2913);
nand U7353 (N_7353,N_5264,N_1915);
or U7354 (N_7354,N_4568,N_5829);
or U7355 (N_7355,N_5146,N_3238);
xnor U7356 (N_7356,N_5631,N_4760);
and U7357 (N_7357,N_1943,N_4570);
and U7358 (N_7358,N_742,N_3714);
or U7359 (N_7359,N_668,N_3013);
nand U7360 (N_7360,N_4743,N_3398);
nand U7361 (N_7361,N_1662,N_4449);
nor U7362 (N_7362,N_4710,N_965);
and U7363 (N_7363,N_4270,N_4116);
and U7364 (N_7364,N_1202,N_416);
and U7365 (N_7365,N_3849,N_5780);
nor U7366 (N_7366,N_2813,N_4695);
and U7367 (N_7367,N_261,N_5940);
and U7368 (N_7368,N_4737,N_3843);
nand U7369 (N_7369,N_1971,N_2708);
xor U7370 (N_7370,N_1819,N_4776);
or U7371 (N_7371,N_2962,N_1924);
or U7372 (N_7372,N_2295,N_4407);
xnor U7373 (N_7373,N_2049,N_2719);
nor U7374 (N_7374,N_5022,N_2053);
and U7375 (N_7375,N_3995,N_2680);
or U7376 (N_7376,N_5043,N_60);
nand U7377 (N_7377,N_4490,N_1767);
nor U7378 (N_7378,N_2347,N_1158);
nand U7379 (N_7379,N_4267,N_4145);
nand U7380 (N_7380,N_803,N_5578);
and U7381 (N_7381,N_970,N_3574);
and U7382 (N_7382,N_3145,N_1343);
or U7383 (N_7383,N_2500,N_5802);
or U7384 (N_7384,N_1069,N_614);
xnor U7385 (N_7385,N_3295,N_1902);
nor U7386 (N_7386,N_850,N_3170);
nor U7387 (N_7387,N_5196,N_4132);
nor U7388 (N_7388,N_48,N_2090);
xnor U7389 (N_7389,N_6149,N_722);
nand U7390 (N_7390,N_5242,N_1671);
or U7391 (N_7391,N_4251,N_1968);
nor U7392 (N_7392,N_2784,N_1884);
nor U7393 (N_7393,N_5129,N_4971);
and U7394 (N_7394,N_5306,N_1374);
nand U7395 (N_7395,N_2099,N_2353);
nor U7396 (N_7396,N_4037,N_4500);
or U7397 (N_7397,N_3270,N_1677);
or U7398 (N_7398,N_5966,N_4122);
and U7399 (N_7399,N_2925,N_1874);
xnor U7400 (N_7400,N_782,N_4686);
nor U7401 (N_7401,N_1415,N_4610);
nand U7402 (N_7402,N_362,N_4264);
and U7403 (N_7403,N_2774,N_4709);
or U7404 (N_7404,N_3249,N_245);
nor U7405 (N_7405,N_717,N_4983);
or U7406 (N_7406,N_85,N_5591);
xnor U7407 (N_7407,N_4895,N_1666);
and U7408 (N_7408,N_3493,N_2260);
xnor U7409 (N_7409,N_4907,N_1136);
xor U7410 (N_7410,N_1822,N_5010);
xor U7411 (N_7411,N_5962,N_4704);
nor U7412 (N_7412,N_4395,N_2218);
nand U7413 (N_7413,N_4102,N_3059);
xnor U7414 (N_7414,N_2185,N_4419);
or U7415 (N_7415,N_1720,N_6032);
nand U7416 (N_7416,N_4229,N_5816);
nand U7417 (N_7417,N_1381,N_5901);
or U7418 (N_7418,N_3194,N_3851);
nor U7419 (N_7419,N_491,N_1795);
xor U7420 (N_7420,N_4689,N_4573);
nor U7421 (N_7421,N_2914,N_1505);
nand U7422 (N_7422,N_5094,N_4724);
xnor U7423 (N_7423,N_510,N_1847);
and U7424 (N_7424,N_1446,N_1976);
or U7425 (N_7425,N_2974,N_5681);
or U7426 (N_7426,N_6079,N_748);
nand U7427 (N_7427,N_2765,N_2501);
nand U7428 (N_7428,N_1755,N_2352);
or U7429 (N_7429,N_1975,N_2111);
nand U7430 (N_7430,N_2648,N_2838);
or U7431 (N_7431,N_776,N_1527);
nand U7432 (N_7432,N_159,N_545);
and U7433 (N_7433,N_2689,N_5730);
nand U7434 (N_7434,N_4597,N_175);
xnor U7435 (N_7435,N_3420,N_2786);
and U7436 (N_7436,N_1741,N_4019);
or U7437 (N_7437,N_4217,N_3876);
nand U7438 (N_7438,N_1329,N_2493);
or U7439 (N_7439,N_5630,N_216);
nand U7440 (N_7440,N_2506,N_2420);
nand U7441 (N_7441,N_4955,N_1149);
nor U7442 (N_7442,N_3372,N_5655);
or U7443 (N_7443,N_2147,N_924);
and U7444 (N_7444,N_5542,N_2664);
or U7445 (N_7445,N_3974,N_3000);
or U7446 (N_7446,N_5914,N_5108);
or U7447 (N_7447,N_6033,N_4245);
and U7448 (N_7448,N_4562,N_2118);
xor U7449 (N_7449,N_788,N_5187);
xnor U7450 (N_7450,N_5925,N_1543);
or U7451 (N_7451,N_5167,N_4466);
xnor U7452 (N_7452,N_3179,N_5704);
or U7453 (N_7453,N_2312,N_3697);
xor U7454 (N_7454,N_3700,N_4208);
nor U7455 (N_7455,N_435,N_5143);
or U7456 (N_7456,N_5472,N_2203);
nand U7457 (N_7457,N_6027,N_5546);
nor U7458 (N_7458,N_1949,N_5917);
nor U7459 (N_7459,N_2596,N_4034);
or U7460 (N_7460,N_2369,N_6047);
and U7461 (N_7461,N_3739,N_5292);
nor U7462 (N_7462,N_1615,N_3168);
xor U7463 (N_7463,N_485,N_2781);
nor U7464 (N_7464,N_648,N_1068);
nor U7465 (N_7465,N_2265,N_4059);
nor U7466 (N_7466,N_4887,N_3645);
and U7467 (N_7467,N_5756,N_2104);
xor U7468 (N_7468,N_1191,N_6012);
xor U7469 (N_7469,N_2968,N_2324);
and U7470 (N_7470,N_3248,N_1268);
nor U7471 (N_7471,N_3695,N_2065);
or U7472 (N_7472,N_191,N_6209);
and U7473 (N_7473,N_2018,N_410);
or U7474 (N_7474,N_3136,N_2743);
and U7475 (N_7475,N_4004,N_3875);
and U7476 (N_7476,N_4682,N_796);
nand U7477 (N_7477,N_1462,N_5048);
nand U7478 (N_7478,N_5386,N_2429);
or U7479 (N_7479,N_2123,N_5937);
nand U7480 (N_7480,N_5139,N_204);
nor U7481 (N_7481,N_4108,N_2390);
nand U7482 (N_7482,N_6227,N_1984);
nand U7483 (N_7483,N_2496,N_2237);
or U7484 (N_7484,N_4441,N_5648);
or U7485 (N_7485,N_3247,N_262);
and U7486 (N_7486,N_2591,N_3193);
and U7487 (N_7487,N_1776,N_1642);
nand U7488 (N_7488,N_5690,N_5814);
nor U7489 (N_7489,N_437,N_6182);
nand U7490 (N_7490,N_5428,N_5453);
nand U7491 (N_7491,N_681,N_1192);
and U7492 (N_7492,N_5134,N_5223);
and U7493 (N_7493,N_3200,N_5373);
xnor U7494 (N_7494,N_5697,N_2033);
nand U7495 (N_7495,N_2141,N_2204);
nand U7496 (N_7496,N_135,N_1410);
or U7497 (N_7497,N_3433,N_5536);
xor U7498 (N_7498,N_1359,N_3197);
nor U7499 (N_7499,N_2703,N_2498);
nand U7500 (N_7500,N_1797,N_3233);
xnor U7501 (N_7501,N_2964,N_4874);
nor U7502 (N_7502,N_2003,N_1009);
and U7503 (N_7503,N_617,N_6207);
or U7504 (N_7504,N_2884,N_1333);
or U7505 (N_7505,N_5111,N_5786);
and U7506 (N_7506,N_2046,N_1371);
or U7507 (N_7507,N_3957,N_121);
or U7508 (N_7508,N_1636,N_5283);
nand U7509 (N_7509,N_412,N_4520);
nand U7510 (N_7510,N_3129,N_3679);
or U7511 (N_7511,N_384,N_557);
or U7512 (N_7512,N_5911,N_4070);
nor U7513 (N_7513,N_1298,N_35);
and U7514 (N_7514,N_3775,N_5712);
xnor U7515 (N_7515,N_511,N_5668);
xnor U7516 (N_7516,N_2035,N_4177);
or U7517 (N_7517,N_6109,N_1779);
xnor U7518 (N_7518,N_692,N_1228);
and U7519 (N_7519,N_3125,N_1687);
xor U7520 (N_7520,N_4136,N_2676);
xnor U7521 (N_7521,N_1070,N_976);
or U7522 (N_7522,N_3084,N_1182);
nand U7523 (N_7523,N_3315,N_3674);
nand U7524 (N_7524,N_5886,N_4271);
xor U7525 (N_7525,N_3304,N_1101);
xor U7526 (N_7526,N_361,N_1288);
xnor U7527 (N_7527,N_2344,N_4020);
nor U7528 (N_7528,N_5246,N_1066);
and U7529 (N_7529,N_2132,N_3906);
nand U7530 (N_7530,N_1905,N_339);
and U7531 (N_7531,N_5406,N_5535);
xor U7532 (N_7532,N_2235,N_3577);
or U7533 (N_7533,N_1107,N_1613);
and U7534 (N_7534,N_3929,N_5506);
nor U7535 (N_7535,N_420,N_4796);
or U7536 (N_7536,N_1270,N_3942);
nand U7537 (N_7537,N_2580,N_5981);
or U7538 (N_7538,N_2376,N_3649);
nand U7539 (N_7539,N_2696,N_1717);
xor U7540 (N_7540,N_1491,N_1624);
nand U7541 (N_7541,N_2224,N_766);
xnor U7542 (N_7542,N_3855,N_1051);
xor U7543 (N_7543,N_1077,N_1608);
and U7544 (N_7544,N_4837,N_567);
or U7545 (N_7545,N_1661,N_3721);
nor U7546 (N_7546,N_5817,N_564);
and U7547 (N_7547,N_1332,N_3405);
nand U7548 (N_7548,N_3293,N_5638);
or U7549 (N_7549,N_3463,N_3279);
and U7550 (N_7550,N_3178,N_2154);
nand U7551 (N_7551,N_4742,N_5653);
and U7552 (N_7552,N_4889,N_5101);
or U7553 (N_7553,N_6005,N_3236);
nor U7554 (N_7554,N_5573,N_901);
xor U7555 (N_7555,N_2371,N_707);
nor U7556 (N_7556,N_251,N_5967);
nor U7557 (N_7557,N_4256,N_4224);
nand U7558 (N_7558,N_2712,N_2683);
xor U7559 (N_7559,N_3539,N_5408);
and U7560 (N_7560,N_4628,N_2548);
and U7561 (N_7561,N_133,N_1104);
and U7562 (N_7562,N_896,N_3035);
or U7563 (N_7563,N_4143,N_5898);
or U7564 (N_7564,N_1940,N_609);
xor U7565 (N_7565,N_3370,N_5813);
nor U7566 (N_7566,N_2459,N_5374);
nand U7567 (N_7567,N_1518,N_5822);
or U7568 (N_7568,N_1052,N_5289);
or U7569 (N_7569,N_504,N_1230);
nand U7570 (N_7570,N_1493,N_1790);
and U7571 (N_7571,N_1986,N_3048);
nor U7572 (N_7572,N_3559,N_3492);
or U7573 (N_7573,N_5627,N_2818);
or U7574 (N_7574,N_2898,N_5267);
and U7575 (N_7575,N_379,N_2205);
xor U7576 (N_7576,N_6098,N_3999);
or U7577 (N_7577,N_4972,N_5588);
and U7578 (N_7578,N_5833,N_5014);
nand U7579 (N_7579,N_282,N_4377);
nor U7580 (N_7580,N_44,N_3746);
and U7581 (N_7581,N_2827,N_519);
nor U7582 (N_7582,N_318,N_344);
and U7583 (N_7583,N_2791,N_4032);
and U7584 (N_7584,N_1702,N_6056);
nor U7585 (N_7585,N_3556,N_4409);
nor U7586 (N_7586,N_2540,N_3596);
or U7587 (N_7587,N_141,N_4761);
xor U7588 (N_7588,N_835,N_832);
nand U7589 (N_7589,N_3529,N_2971);
or U7590 (N_7590,N_3155,N_1396);
nor U7591 (N_7591,N_4425,N_1800);
xnor U7592 (N_7592,N_6048,N_723);
nand U7593 (N_7593,N_4321,N_1204);
nand U7594 (N_7594,N_2421,N_4203);
or U7595 (N_7595,N_4080,N_2869);
xor U7596 (N_7596,N_6213,N_3598);
and U7597 (N_7597,N_643,N_489);
nor U7598 (N_7598,N_2937,N_246);
xor U7599 (N_7599,N_5834,N_2119);
nor U7600 (N_7600,N_3637,N_1727);
xor U7601 (N_7601,N_1037,N_3936);
xnor U7602 (N_7602,N_3510,N_2872);
nor U7603 (N_7603,N_2299,N_6196);
xnor U7604 (N_7604,N_4938,N_2273);
xor U7605 (N_7605,N_532,N_953);
or U7606 (N_7606,N_3847,N_774);
xnor U7607 (N_7607,N_4471,N_2379);
xor U7608 (N_7608,N_4085,N_2289);
or U7609 (N_7609,N_6205,N_1296);
xor U7610 (N_7610,N_4296,N_6131);
or U7611 (N_7611,N_2701,N_4572);
nand U7612 (N_7612,N_2066,N_1565);
and U7613 (N_7613,N_2853,N_3081);
nor U7614 (N_7614,N_982,N_3092);
and U7615 (N_7615,N_1532,N_6110);
xor U7616 (N_7616,N_256,N_1341);
xor U7617 (N_7617,N_263,N_5879);
nand U7618 (N_7618,N_1012,N_5);
and U7619 (N_7619,N_6230,N_1620);
nand U7620 (N_7620,N_3514,N_130);
nor U7621 (N_7621,N_5282,N_2839);
nor U7622 (N_7622,N_4623,N_5041);
xor U7623 (N_7623,N_2174,N_1590);
or U7624 (N_7624,N_3144,N_1143);
nand U7625 (N_7625,N_4828,N_3764);
and U7626 (N_7626,N_5423,N_4673);
nor U7627 (N_7627,N_1220,N_2112);
nand U7628 (N_7628,N_1,N_108);
nand U7629 (N_7629,N_2556,N_2194);
xnor U7630 (N_7630,N_6062,N_3928);
nor U7631 (N_7631,N_4342,N_5715);
nand U7632 (N_7632,N_1399,N_5773);
xor U7633 (N_7633,N_5203,N_5942);
xor U7634 (N_7634,N_1775,N_1675);
xnor U7635 (N_7635,N_4890,N_5765);
and U7636 (N_7636,N_5157,N_2718);
xor U7637 (N_7637,N_5695,N_3589);
or U7638 (N_7638,N_4750,N_2587);
or U7639 (N_7639,N_2769,N_4635);
or U7640 (N_7640,N_6071,N_2076);
or U7641 (N_7641,N_4728,N_880);
and U7642 (N_7642,N_2731,N_5924);
xnor U7643 (N_7643,N_6072,N_4024);
or U7644 (N_7644,N_1240,N_4733);
or U7645 (N_7645,N_1354,N_2109);
and U7646 (N_7646,N_538,N_5076);
nand U7647 (N_7647,N_4995,N_1585);
and U7648 (N_7648,N_3039,N_3323);
and U7649 (N_7649,N_292,N_4824);
nor U7650 (N_7650,N_927,N_5106);
nand U7651 (N_7651,N_3234,N_6164);
nor U7652 (N_7652,N_347,N_2184);
nand U7653 (N_7653,N_1658,N_1407);
nand U7654 (N_7654,N_3550,N_5465);
nand U7655 (N_7655,N_4351,N_842);
or U7656 (N_7656,N_3772,N_541);
nor U7657 (N_7657,N_5841,N_3336);
and U7658 (N_7658,N_1413,N_5531);
or U7659 (N_7659,N_711,N_6070);
or U7660 (N_7660,N_6101,N_97);
or U7661 (N_7661,N_4120,N_2846);
xor U7662 (N_7662,N_5319,N_2162);
nand U7663 (N_7663,N_2726,N_4050);
or U7664 (N_7664,N_750,N_5727);
and U7665 (N_7665,N_2720,N_2477);
and U7666 (N_7666,N_3329,N_120);
and U7667 (N_7667,N_1443,N_879);
or U7668 (N_7668,N_162,N_3382);
and U7669 (N_7669,N_625,N_80);
or U7670 (N_7670,N_3741,N_3090);
nand U7671 (N_7671,N_5381,N_2100);
nand U7672 (N_7672,N_4434,N_4785);
xnor U7673 (N_7673,N_3221,N_1737);
xor U7674 (N_7674,N_1913,N_1039);
and U7675 (N_7675,N_241,N_2093);
nor U7676 (N_7676,N_938,N_2923);
nand U7677 (N_7677,N_254,N_3523);
nand U7678 (N_7678,N_769,N_5639);
nor U7679 (N_7679,N_4916,N_1036);
and U7680 (N_7680,N_3033,N_6175);
nor U7681 (N_7681,N_5764,N_1384);
xor U7682 (N_7682,N_6118,N_1703);
nand U7683 (N_7683,N_29,N_4977);
or U7684 (N_7684,N_6102,N_5084);
xor U7685 (N_7685,N_2305,N_2157);
or U7686 (N_7686,N_2019,N_1003);
and U7687 (N_7687,N_533,N_2497);
and U7688 (N_7688,N_197,N_2293);
and U7689 (N_7689,N_5825,N_3327);
nand U7690 (N_7690,N_319,N_1120);
nor U7691 (N_7691,N_315,N_2437);
or U7692 (N_7692,N_3563,N_2139);
or U7693 (N_7693,N_6077,N_593);
and U7694 (N_7694,N_3718,N_1678);
nand U7695 (N_7695,N_1957,N_5711);
nor U7696 (N_7696,N_4582,N_3297);
and U7697 (N_7697,N_5582,N_756);
and U7698 (N_7698,N_4452,N_865);
xor U7699 (N_7699,N_1616,N_1647);
nand U7700 (N_7700,N_1378,N_184);
nor U7701 (N_7701,N_3802,N_5516);
nor U7702 (N_7702,N_5393,N_1448);
xor U7703 (N_7703,N_3334,N_4542);
or U7704 (N_7704,N_75,N_2917);
nand U7705 (N_7705,N_6181,N_1972);
or U7706 (N_7706,N_4220,N_5046);
and U7707 (N_7707,N_4325,N_5998);
xnor U7708 (N_7708,N_1535,N_4678);
or U7709 (N_7709,N_3460,N_3980);
nand U7710 (N_7710,N_1091,N_5983);
or U7711 (N_7711,N_2582,N_2512);
or U7712 (N_7712,N_5171,N_758);
xnor U7713 (N_7713,N_3476,N_4412);
or U7714 (N_7714,N_4814,N_1893);
or U7715 (N_7715,N_4273,N_1552);
or U7716 (N_7716,N_1879,N_1460);
nand U7717 (N_7717,N_5953,N_4184);
nor U7718 (N_7718,N_6202,N_2879);
xor U7719 (N_7719,N_1595,N_1747);
and U7720 (N_7720,N_2131,N_2407);
xor U7721 (N_7721,N_2523,N_1115);
xor U7722 (N_7722,N_5288,N_5219);
xor U7723 (N_7723,N_6215,N_1236);
xor U7724 (N_7724,N_5805,N_918);
nor U7725 (N_7725,N_2904,N_1046);
or U7726 (N_7726,N_3804,N_5760);
nand U7727 (N_7727,N_4130,N_4713);
or U7728 (N_7728,N_2722,N_4420);
nand U7729 (N_7729,N_1183,N_2707);
and U7730 (N_7730,N_2597,N_223);
or U7731 (N_7731,N_5092,N_3791);
or U7732 (N_7732,N_3698,N_4513);
nor U7733 (N_7733,N_4235,N_3709);
xor U7734 (N_7734,N_3988,N_2758);
or U7735 (N_7735,N_824,N_5892);
nand U7736 (N_7736,N_4390,N_2697);
xnor U7737 (N_7737,N_534,N_2438);
nand U7738 (N_7738,N_1896,N_5771);
nand U7739 (N_7739,N_1831,N_2654);
xnor U7740 (N_7740,N_501,N_4237);
nor U7741 (N_7741,N_2552,N_2715);
and U7742 (N_7742,N_1059,N_1609);
nor U7743 (N_7743,N_2336,N_1988);
or U7744 (N_7744,N_2644,N_5663);
or U7745 (N_7745,N_3253,N_1218);
nand U7746 (N_7746,N_4627,N_5326);
nor U7747 (N_7747,N_2170,N_2187);
and U7748 (N_7748,N_5567,N_247);
nor U7749 (N_7749,N_2566,N_5379);
xnor U7750 (N_7750,N_574,N_2604);
xor U7751 (N_7751,N_1989,N_185);
nand U7752 (N_7752,N_5133,N_940);
nor U7753 (N_7753,N_2431,N_183);
and U7754 (N_7754,N_4499,N_2561);
xnor U7755 (N_7755,N_2308,N_31);
or U7756 (N_7756,N_5545,N_4571);
or U7757 (N_7757,N_604,N_646);
or U7758 (N_7758,N_4283,N_3853);
xor U7759 (N_7759,N_2734,N_217);
nand U7760 (N_7760,N_2608,N_1105);
xor U7761 (N_7761,N_1676,N_3553);
and U7762 (N_7762,N_2992,N_3842);
or U7763 (N_7763,N_1173,N_3590);
and U7764 (N_7764,N_1768,N_2875);
or U7765 (N_7765,N_6091,N_2931);
or U7766 (N_7766,N_5863,N_2024);
and U7767 (N_7767,N_2357,N_5271);
nor U7768 (N_7768,N_3410,N_3068);
nor U7769 (N_7769,N_5215,N_372);
xnor U7770 (N_7770,N_401,N_227);
nand U7771 (N_7771,N_812,N_429);
nor U7772 (N_7772,N_4077,N_618);
nand U7773 (N_7773,N_3055,N_2415);
or U7774 (N_7774,N_4337,N_1235);
nand U7775 (N_7775,N_3570,N_3898);
or U7776 (N_7776,N_4149,N_2592);
or U7777 (N_7777,N_2638,N_1469);
and U7778 (N_7778,N_2916,N_5037);
nor U7779 (N_7779,N_2954,N_5334);
or U7780 (N_7780,N_86,N_4257);
or U7781 (N_7781,N_4575,N_2820);
xor U7782 (N_7782,N_3086,N_375);
nor U7783 (N_7783,N_4636,N_3494);
and U7784 (N_7784,N_1328,N_161);
and U7785 (N_7785,N_1698,N_4105);
or U7786 (N_7786,N_5207,N_4727);
xor U7787 (N_7787,N_5831,N_6146);
nand U7788 (N_7788,N_293,N_4504);
or U7789 (N_7789,N_4708,N_386);
nand U7790 (N_7790,N_2549,N_2595);
nand U7791 (N_7791,N_4451,N_5354);
and U7792 (N_7792,N_2739,N_4225);
nor U7793 (N_7793,N_5053,N_278);
nor U7794 (N_7794,N_4706,N_1449);
nand U7795 (N_7795,N_4655,N_4604);
and U7796 (N_7796,N_4218,N_1742);
nand U7797 (N_7797,N_5250,N_888);
nand U7798 (N_7798,N_5494,N_2662);
nor U7799 (N_7799,N_3458,N_4659);
nor U7800 (N_7800,N_1521,N_2255);
or U7801 (N_7801,N_4860,N_848);
xnor U7802 (N_7802,N_1855,N_370);
nor U7803 (N_7803,N_209,N_348);
or U7804 (N_7804,N_3325,N_3074);
nand U7805 (N_7805,N_3140,N_4770);
nor U7806 (N_7806,N_3963,N_1194);
and U7807 (N_7807,N_2107,N_2427);
or U7808 (N_7808,N_2522,N_3885);
xor U7809 (N_7809,N_3266,N_1930);
and U7810 (N_7810,N_1291,N_3181);
xnor U7811 (N_7811,N_5979,N_765);
nor U7812 (N_7812,N_490,N_2298);
or U7813 (N_7813,N_1100,N_1367);
or U7814 (N_7814,N_2528,N_2599);
or U7815 (N_7815,N_3309,N_3251);
nor U7816 (N_7816,N_4882,N_6185);
or U7817 (N_7817,N_1138,N_5989);
and U7818 (N_7818,N_3519,N_4190);
nor U7819 (N_7819,N_3239,N_1441);
nand U7820 (N_7820,N_5112,N_2057);
xnor U7821 (N_7821,N_2317,N_2899);
xor U7822 (N_7822,N_4694,N_513);
or U7823 (N_7823,N_2007,N_1133);
xor U7824 (N_7824,N_1362,N_802);
and U7825 (N_7825,N_5781,N_806);
xnor U7826 (N_7826,N_4840,N_3412);
nand U7827 (N_7827,N_3783,N_4603);
nand U7828 (N_7828,N_3736,N_3311);
or U7829 (N_7829,N_6198,N_3891);
and U7830 (N_7830,N_4263,N_4991);
xor U7831 (N_7831,N_1600,N_943);
xnor U7832 (N_7832,N_317,N_189);
nor U7833 (N_7833,N_762,N_3119);
and U7834 (N_7834,N_1154,N_4106);
xor U7835 (N_7835,N_5072,N_1869);
and U7836 (N_7836,N_4331,N_3609);
or U7837 (N_7837,N_3904,N_3431);
nand U7838 (N_7838,N_4356,N_3139);
nand U7839 (N_7839,N_6094,N_773);
nand U7840 (N_7840,N_1562,N_5217);
and U7841 (N_7841,N_1572,N_365);
and U7842 (N_7842,N_1040,N_2450);
and U7843 (N_7843,N_258,N_2823);
xor U7844 (N_7844,N_6037,N_3560);
nor U7845 (N_7845,N_620,N_5042);
or U7846 (N_7846,N_2952,N_394);
or U7847 (N_7847,N_4072,N_1227);
nand U7848 (N_7848,N_2063,N_164);
and U7849 (N_7849,N_4371,N_129);
or U7850 (N_7850,N_330,N_1047);
xor U7851 (N_7851,N_5064,N_4083);
xor U7852 (N_7852,N_117,N_3371);
nor U7853 (N_7853,N_1882,N_4168);
xnor U7854 (N_7854,N_1711,N_588);
and U7855 (N_7855,N_4791,N_371);
or U7856 (N_7856,N_474,N_1403);
and U7857 (N_7857,N_3977,N_563);
xor U7858 (N_7858,N_4000,N_1589);
xor U7859 (N_7859,N_3105,N_27);
nand U7860 (N_7860,N_5164,N_67);
and U7861 (N_7861,N_4022,N_4212);
xor U7862 (N_7862,N_1159,N_4487);
nor U7863 (N_7863,N_2588,N_190);
and U7864 (N_7864,N_1420,N_2042);
nor U7865 (N_7865,N_5577,N_3806);
xnor U7866 (N_7866,N_2568,N_645);
xor U7867 (N_7867,N_4448,N_5295);
xnor U7868 (N_7868,N_2087,N_3322);
nor U7869 (N_7869,N_5992,N_3025);
nand U7870 (N_7870,N_3689,N_2574);
and U7871 (N_7871,N_248,N_3362);
xnor U7872 (N_7872,N_5478,N_1279);
and U7873 (N_7873,N_6200,N_3150);
nand U7874 (N_7874,N_718,N_5371);
xnor U7875 (N_7875,N_5867,N_1567);
and U7876 (N_7876,N_277,N_3417);
and U7877 (N_7877,N_4038,N_4612);
nor U7878 (N_7878,N_5719,N_3389);
and U7879 (N_7879,N_1103,N_1315);
nand U7880 (N_7880,N_2618,N_1434);
and U7881 (N_7881,N_5676,N_453);
or U7882 (N_7882,N_2792,N_1504);
and U7883 (N_7883,N_357,N_5433);
xor U7884 (N_7884,N_358,N_1961);
xnor U7885 (N_7885,N_4403,N_3043);
or U7886 (N_7886,N_4528,N_4868);
or U7887 (N_7887,N_3882,N_527);
xor U7888 (N_7888,N_4126,N_3245);
or U7889 (N_7889,N_5560,N_1835);
nand U7890 (N_7890,N_4285,N_5963);
and U7891 (N_7891,N_3762,N_196);
and U7892 (N_7892,N_6125,N_905);
nor U7893 (N_7893,N_6242,N_2641);
nor U7894 (N_7894,N_1928,N_1232);
nand U7895 (N_7895,N_4872,N_3971);
nand U7896 (N_7896,N_1023,N_606);
xnor U7897 (N_7897,N_3008,N_465);
and U7898 (N_7898,N_4410,N_4547);
and U7899 (N_7899,N_4320,N_1000);
and U7900 (N_7900,N_2787,N_1550);
nand U7901 (N_7901,N_1073,N_2021);
and U7902 (N_7902,N_4845,N_1334);
nand U7903 (N_7903,N_2257,N_2160);
xor U7904 (N_7904,N_2602,N_1992);
nor U7905 (N_7905,N_5030,N_90);
xor U7906 (N_7906,N_1248,N_5348);
and U7907 (N_7907,N_1890,N_4747);
xnor U7908 (N_7908,N_5073,N_2106);
xor U7909 (N_7909,N_3246,N_4221);
xnor U7910 (N_7910,N_5980,N_2575);
nor U7911 (N_7911,N_4195,N_4346);
xor U7912 (N_7912,N_2143,N_2636);
nand U7913 (N_7913,N_5174,N_2752);
xor U7914 (N_7914,N_6115,N_3620);
or U7915 (N_7915,N_3857,N_922);
nand U7916 (N_7916,N_383,N_2291);
or U7917 (N_7917,N_5051,N_2694);
xor U7918 (N_7918,N_5298,N_1206);
nor U7919 (N_7919,N_4373,N_811);
nor U7920 (N_7920,N_3651,N_5700);
nor U7921 (N_7921,N_6218,N_3377);
nor U7922 (N_7922,N_4370,N_3094);
nor U7923 (N_7923,N_4883,N_56);
nand U7924 (N_7924,N_2491,N_275);
or U7925 (N_7925,N_575,N_3347);
xnor U7926 (N_7926,N_2666,N_4738);
nand U7927 (N_7927,N_4815,N_1546);
nor U7928 (N_7928,N_1626,N_5930);
nand U7929 (N_7929,N_5121,N_6112);
or U7930 (N_7930,N_2706,N_4087);
nand U7931 (N_7931,N_4423,N_1709);
nand U7932 (N_7932,N_5476,N_5208);
or U7933 (N_7933,N_781,N_2483);
xnor U7934 (N_7934,N_5065,N_5949);
xor U7935 (N_7935,N_2620,N_3019);
and U7936 (N_7936,N_3138,N_4075);
or U7937 (N_7937,N_4101,N_4436);
nand U7938 (N_7938,N_1761,N_2077);
nor U7939 (N_7939,N_4300,N_1109);
nand U7940 (N_7940,N_3781,N_3228);
or U7941 (N_7941,N_3445,N_517);
and U7942 (N_7942,N_4913,N_969);
nor U7943 (N_7943,N_5368,N_4927);
and U7944 (N_7944,N_210,N_2436);
xnor U7945 (N_7945,N_4380,N_2125);
nor U7946 (N_7946,N_624,N_5600);
and U7947 (N_7947,N_3489,N_4189);
or U7948 (N_7948,N_677,N_5380);
nor U7949 (N_7949,N_6216,N_898);
nor U7950 (N_7950,N_3547,N_846);
and U7951 (N_7951,N_188,N_5894);
xnor U7952 (N_7952,N_1514,N_281);
nor U7953 (N_7953,N_1088,N_5336);
nand U7954 (N_7954,N_284,N_6086);
nand U7955 (N_7955,N_5316,N_1335);
nor U7956 (N_7956,N_3284,N_4862);
or U7957 (N_7957,N_3877,N_2017);
nor U7958 (N_7958,N_6089,N_854);
xnor U7959 (N_7959,N_3388,N_1894);
and U7960 (N_7960,N_903,N_4222);
nor U7961 (N_7961,N_1001,N_1169);
nand U7962 (N_7962,N_933,N_5951);
and U7963 (N_7963,N_2254,N_1238);
xnor U7964 (N_7964,N_2277,N_962);
xnor U7965 (N_7965,N_6082,N_1953);
xnor U7966 (N_7966,N_2098,N_2023);
and U7967 (N_7967,N_1715,N_2068);
or U7968 (N_7968,N_442,N_4850);
nand U7969 (N_7969,N_2764,N_800);
and U7970 (N_7970,N_5483,N_874);
nor U7971 (N_7971,N_6187,N_5783);
and U7972 (N_7972,N_334,N_495);
nand U7973 (N_7973,N_5454,N_6229);
xnor U7974 (N_7974,N_590,N_3275);
xnor U7975 (N_7975,N_451,N_5029);
nand U7976 (N_7976,N_5533,N_5302);
nand U7977 (N_7977,N_4473,N_3403);
and U7978 (N_7978,N_1638,N_3521);
nand U7979 (N_7979,N_2229,N_4366);
nand U7980 (N_7980,N_1805,N_5057);
nor U7981 (N_7981,N_512,N_4514);
nand U7982 (N_7982,N_3301,N_3340);
nor U7983 (N_7983,N_6117,N_5965);
nand U7984 (N_7984,N_988,N_3357);
xnor U7985 (N_7985,N_4497,N_6231);
and U7986 (N_7986,N_39,N_4848);
xnor U7987 (N_7987,N_1010,N_4929);
xor U7988 (N_7988,N_1111,N_5107);
nand U7989 (N_7989,N_5154,N_696);
or U7990 (N_7990,N_568,N_3353);
and U7991 (N_7991,N_3305,N_5922);
nand U7992 (N_7992,N_2167,N_1431);
xnor U7993 (N_7993,N_3222,N_2663);
or U7994 (N_7994,N_2453,N_1146);
xor U7995 (N_7995,N_2179,N_4580);
and U7996 (N_7996,N_727,N_641);
nor U7997 (N_7997,N_1777,N_2628);
and U7998 (N_7998,N_107,N_2891);
nand U7999 (N_7999,N_5007,N_2349);
and U8000 (N_8000,N_5091,N_4624);
xnor U8001 (N_8001,N_3606,N_4397);
or U8002 (N_8002,N_1044,N_3592);
and U8003 (N_8003,N_900,N_3925);
xor U8004 (N_8004,N_2607,N_753);
nand U8005 (N_8005,N_621,N_3676);
nand U8006 (N_8006,N_2655,N_1632);
nand U8007 (N_8007,N_5988,N_1936);
and U8008 (N_8008,N_2989,N_5609);
or U8009 (N_8009,N_2455,N_62);
or U8010 (N_8010,N_5463,N_3961);
xor U8011 (N_8011,N_5232,N_1114);
and U8012 (N_8012,N_1523,N_2314);
and U8013 (N_8013,N_494,N_3217);
or U8014 (N_8014,N_3684,N_5611);
and U8015 (N_8015,N_5908,N_1821);
and U8016 (N_8016,N_268,N_3341);
nand U8017 (N_8017,N_3108,N_321);
xor U8018 (N_8018,N_966,N_337);
and U8019 (N_8019,N_1789,N_631);
nand U8020 (N_8020,N_878,N_4586);
xor U8021 (N_8021,N_5739,N_5735);
nand U8022 (N_8022,N_2841,N_1652);
xnor U8023 (N_8023,N_4975,N_4543);
and U8024 (N_8024,N_4305,N_550);
and U8025 (N_8025,N_4665,N_3379);
or U8026 (N_8026,N_4073,N_3827);
or U8027 (N_8027,N_4993,N_2824);
or U8028 (N_8028,N_3992,N_400);
nor U8029 (N_8029,N_6214,N_2821);
and U8030 (N_8030,N_2207,N_1617);
xnor U8031 (N_8031,N_415,N_5594);
nand U8032 (N_8032,N_777,N_3424);
and U8033 (N_8033,N_5323,N_4979);
or U8034 (N_8034,N_3421,N_838);
nand U8035 (N_8035,N_2329,N_2014);
or U8036 (N_8036,N_1450,N_6030);
and U8037 (N_8037,N_1654,N_2995);
xnor U8038 (N_8038,N_6054,N_4347);
xor U8039 (N_8039,N_1089,N_208);
xor U8040 (N_8040,N_2862,N_6019);
or U8041 (N_8041,N_3042,N_5204);
nand U8042 (N_8042,N_4609,N_3488);
nor U8043 (N_8043,N_4622,N_5411);
nor U8044 (N_8044,N_4584,N_4291);
nand U8045 (N_8045,N_1297,N_2309);
and U8046 (N_8046,N_1649,N_5580);
and U8047 (N_8047,N_813,N_96);
xnor U8048 (N_8048,N_2370,N_4569);
nand U8049 (N_8049,N_5160,N_4254);
nand U8050 (N_8050,N_2541,N_4302);
nand U8051 (N_8051,N_1830,N_5875);
xnor U8052 (N_8052,N_5747,N_5436);
nor U8053 (N_8053,N_2878,N_912);
xnor U8054 (N_8054,N_2918,N_3486);
or U8055 (N_8055,N_1464,N_5587);
xor U8056 (N_8056,N_1931,N_1481);
and U8057 (N_8057,N_2408,N_1483);
or U8058 (N_8058,N_925,N_1840);
xnor U8059 (N_8059,N_366,N_1564);
nand U8060 (N_8060,N_4817,N_1713);
and U8061 (N_8061,N_5874,N_5178);
or U8062 (N_8062,N_3393,N_4344);
nor U8063 (N_8063,N_2140,N_2011);
and U8064 (N_8064,N_3177,N_5857);
nand U8065 (N_8065,N_642,N_920);
nor U8066 (N_8066,N_4478,N_3051);
xnor U8067 (N_8067,N_4940,N_5017);
nor U8068 (N_8068,N_4469,N_2569);
or U8069 (N_8069,N_1316,N_2058);
and U8070 (N_8070,N_3274,N_5493);
and U8071 (N_8071,N_899,N_4819);
or U8072 (N_8072,N_1349,N_4005);
nand U8073 (N_8073,N_4111,N_4771);
and U8074 (N_8074,N_5666,N_1722);
or U8075 (N_8075,N_1644,N_3206);
nor U8076 (N_8076,N_3500,N_1207);
nor U8077 (N_8077,N_3868,N_5198);
nand U8078 (N_8078,N_1509,N_611);
nor U8079 (N_8079,N_4472,N_1099);
and U8080 (N_8080,N_2462,N_2094);
nand U8081 (N_8081,N_1060,N_1287);
nand U8082 (N_8082,N_1394,N_1916);
or U8083 (N_8083,N_1979,N_1657);
and U8084 (N_8084,N_4012,N_873);
nand U8085 (N_8085,N_522,N_5457);
xor U8086 (N_8086,N_6050,N_1033);
or U8087 (N_8087,N_4428,N_28);
nor U8088 (N_8088,N_4181,N_4233);
nor U8089 (N_8089,N_5401,N_601);
and U8090 (N_8090,N_1042,N_4376);
or U8091 (N_8091,N_16,N_5331);
xnor U8092 (N_8092,N_5502,N_5474);
or U8093 (N_8093,N_1199,N_923);
nor U8094 (N_8094,N_1942,N_1674);
nand U8095 (N_8095,N_4328,N_5403);
and U8096 (N_8096,N_2665,N_2283);
nand U8097 (N_8097,N_4125,N_1889);
xor U8098 (N_8098,N_3012,N_5163);
and U8099 (N_8099,N_5677,N_5222);
xnor U8100 (N_8100,N_122,N_6009);
xnor U8101 (N_8101,N_3822,N_3710);
nor U8102 (N_8102,N_1282,N_2323);
nor U8103 (N_8103,N_3478,N_4293);
or U8104 (N_8104,N_249,N_5672);
and U8105 (N_8105,N_4506,N_2002);
xor U8106 (N_8106,N_4803,N_1402);
nand U8107 (N_8107,N_2025,N_4402);
nor U8108 (N_8108,N_2700,N_5093);
xor U8109 (N_8109,N_5543,N_4900);
xor U8110 (N_8110,N_1391,N_444);
xnor U8111 (N_8111,N_5947,N_1875);
nand U8112 (N_8112,N_2252,N_999);
xor U8113 (N_8113,N_5686,N_350);
xor U8114 (N_8114,N_5297,N_4129);
xnor U8115 (N_8115,N_5657,N_2441);
nor U8116 (N_8116,N_4700,N_81);
xor U8117 (N_8117,N_4801,N_110);
nor U8118 (N_8118,N_2646,N_6148);
nor U8119 (N_8119,N_1618,N_3872);
nand U8120 (N_8120,N_338,N_2059);
xor U8121 (N_8121,N_119,N_3897);
and U8122 (N_8122,N_2227,N_1860);
or U8123 (N_8123,N_5450,N_4275);
nor U8124 (N_8124,N_1260,N_5253);
and U8125 (N_8125,N_4197,N_4041);
nand U8126 (N_8126,N_5873,N_2296);
or U8127 (N_8127,N_5819,N_5189);
nor U8128 (N_8128,N_1852,N_2325);
or U8129 (N_8129,N_2756,N_3404);
xnor U8130 (N_8130,N_2028,N_4675);
nor U8131 (N_8131,N_5909,N_2165);
nand U8132 (N_8132,N_771,N_3286);
or U8133 (N_8133,N_66,N_2262);
and U8134 (N_8134,N_5270,N_2744);
nand U8135 (N_8135,N_799,N_3667);
xnor U8136 (N_8136,N_1579,N_4290);
nand U8137 (N_8137,N_1222,N_5846);
nand U8138 (N_8138,N_3250,N_1641);
nor U8139 (N_8139,N_2108,N_4018);
xnor U8140 (N_8140,N_5972,N_5931);
and U8141 (N_8141,N_2911,N_2908);
xor U8142 (N_8142,N_2351,N_1085);
nand U8143 (N_8143,N_165,N_3367);
nor U8144 (N_8144,N_2688,N_5176);
and U8145 (N_8145,N_3023,N_945);
and U8146 (N_8146,N_4606,N_2979);
nor U8147 (N_8147,N_1762,N_1233);
nor U8148 (N_8148,N_726,N_461);
and U8149 (N_8149,N_572,N_4757);
or U8150 (N_8150,N_4856,N_4110);
and U8151 (N_8151,N_1002,N_299);
and U8152 (N_8152,N_4440,N_4158);
nor U8153 (N_8153,N_1300,N_178);
and U8154 (N_8154,N_487,N_5708);
xnor U8155 (N_8155,N_554,N_5865);
nand U8156 (N_8156,N_1982,N_6140);
nand U8157 (N_8157,N_1558,N_2716);
nor U8158 (N_8158,N_5793,N_2361);
and U8159 (N_8159,N_5410,N_132);
or U8160 (N_8160,N_3213,N_2290);
or U8161 (N_8161,N_142,N_3658);
nand U8162 (N_8162,N_4692,N_500);
and U8163 (N_8163,N_6243,N_4579);
xnor U8164 (N_8164,N_3994,N_2113);
or U8165 (N_8165,N_4182,N_2342);
xor U8166 (N_8166,N_2550,N_3728);
and U8167 (N_8167,N_3271,N_459);
nand U8168 (N_8168,N_5599,N_910);
or U8169 (N_8169,N_8,N_314);
and U8170 (N_8170,N_276,N_1187);
nor U8171 (N_8171,N_6186,N_2181);
nor U8172 (N_8172,N_3575,N_3396);
or U8173 (N_8173,N_685,N_5714);
nor U8174 (N_8174,N_4601,N_3948);
nor U8175 (N_8175,N_4548,N_440);
nand U8176 (N_8176,N_1740,N_5650);
nand U8177 (N_8177,N_4104,N_3668);
nand U8178 (N_8178,N_555,N_126);
and U8179 (N_8179,N_2015,N_4773);
and U8180 (N_8180,N_4787,N_1412);
and U8181 (N_8181,N_2554,N_2741);
nand U8182 (N_8182,N_3123,N_738);
xnor U8183 (N_8183,N_1956,N_1026);
nor U8184 (N_8184,N_2770,N_5376);
or U8185 (N_8185,N_4011,N_3211);
xnor U8186 (N_8186,N_3324,N_4672);
xnor U8187 (N_8187,N_5311,N_2975);
and U8188 (N_8188,N_5725,N_2808);
nor U8189 (N_8189,N_2833,N_817);
nand U8190 (N_8190,N_5970,N_1799);
nand U8191 (N_8191,N_977,N_4433);
and U8192 (N_8192,N_4683,N_1438);
or U8193 (N_8193,N_4879,N_3537);
and U8194 (N_8194,N_1939,N_4952);
or U8195 (N_8195,N_3825,N_3254);
xnor U8196 (N_8196,N_4330,N_5659);
and U8197 (N_8197,N_3291,N_3269);
nor U8198 (N_8198,N_1692,N_979);
nor U8199 (N_8199,N_5569,N_2749);
xnor U8200 (N_8200,N_959,N_5785);
nand U8201 (N_8201,N_301,N_3959);
or U8202 (N_8202,N_3534,N_5188);
xnor U8203 (N_8203,N_2782,N_4082);
and U8204 (N_8204,N_4632,N_3951);
and U8205 (N_8205,N_3428,N_377);
nor U8206 (N_8206,N_4417,N_5568);
and U8207 (N_8207,N_3103,N_1824);
or U8208 (N_8208,N_1094,N_3256);
nand U8209 (N_8209,N_1482,N_4248);
xor U8210 (N_8210,N_1006,N_5404);
or U8211 (N_8211,N_4323,N_3312);
nor U8212 (N_8212,N_1730,N_3032);
nand U8213 (N_8213,N_5929,N_1458);
or U8214 (N_8214,N_4886,N_5058);
nor U8215 (N_8215,N_797,N_2311);
and U8216 (N_8216,N_3135,N_6237);
nand U8217 (N_8217,N_23,N_3531);
nand U8218 (N_8218,N_224,N_5124);
xor U8219 (N_8219,N_4922,N_950);
xor U8220 (N_8220,N_2217,N_414);
or U8221 (N_8221,N_1086,N_307);
or U8222 (N_8222,N_4064,N_4006);
or U8223 (N_8223,N_4349,N_2138);
nand U8224 (N_8224,N_2333,N_2976);
and U8225 (N_8225,N_5696,N_2268);
xnor U8226 (N_8226,N_5071,N_2867);
nor U8227 (N_8227,N_5241,N_5647);
nand U8228 (N_8228,N_2247,N_5260);
and U8229 (N_8229,N_1345,N_5144);
and U8230 (N_8230,N_578,N_477);
nor U8231 (N_8231,N_3966,N_3901);
xnor U8232 (N_8232,N_1166,N_77);
or U8233 (N_8233,N_6169,N_116);
or U8234 (N_8234,N_1980,N_2866);
or U8235 (N_8235,N_2034,N_4304);
and U8236 (N_8236,N_2142,N_822);
nor U8237 (N_8237,N_5861,N_4715);
xor U8238 (N_8238,N_868,N_1217);
nand U8239 (N_8239,N_3636,N_3914);
xnor U8240 (N_8240,N_4175,N_616);
nor U8241 (N_8241,N_2006,N_3079);
xor U8242 (N_8242,N_4740,N_4550);
nand U8243 (N_8243,N_904,N_4703);
xor U8244 (N_8244,N_3050,N_1045);
or U8245 (N_8245,N_6171,N_730);
xor U8246 (N_8246,N_3124,N_3422);
and U8247 (N_8247,N_1695,N_2621);
and U8248 (N_8248,N_2804,N_2651);
or U8249 (N_8249,N_5498,N_705);
and U8250 (N_8250,N_2383,N_2239);
nor U8251 (N_8251,N_252,N_2887);
nor U8252 (N_8252,N_3996,N_3142);
or U8253 (N_8253,N_3418,N_2778);
nor U8254 (N_8254,N_6247,N_2208);
or U8255 (N_8255,N_2732,N_4968);
nand U8256 (N_8256,N_1387,N_2081);
xnor U8257 (N_8257,N_5118,N_4468);
nand U8258 (N_8258,N_1181,N_3737);
nand U8259 (N_8259,N_6235,N_5424);
and U8260 (N_8260,N_1295,N_514);
xor U8261 (N_8261,N_767,N_4574);
nor U8262 (N_8262,N_2,N_5665);
xor U8263 (N_8263,N_3581,N_4359);
xnor U8264 (N_8264,N_1401,N_4759);
nor U8265 (N_8265,N_100,N_4289);
nand U8266 (N_8266,N_2460,N_5860);
xor U8267 (N_8267,N_5977,N_335);
nand U8268 (N_8268,N_1209,N_3109);
and U8269 (N_8269,N_4732,N_2961);
nand U8270 (N_8270,N_1322,N_328);
nor U8271 (N_8271,N_2585,N_4790);
nand U8272 (N_8272,N_432,N_656);
and U8273 (N_8273,N_4299,N_6119);
nor U8274 (N_8274,N_5466,N_4705);
nand U8275 (N_8275,N_3241,N_4541);
and U8276 (N_8276,N_155,N_5683);
or U8277 (N_8277,N_389,N_5299);
or U8278 (N_8278,N_296,N_1277);
or U8279 (N_8279,N_1265,N_968);
xnor U8280 (N_8280,N_4718,N_311);
nor U8281 (N_8281,N_3656,N_861);
and U8282 (N_8282,N_5504,N_2750);
nor U8283 (N_8283,N_6041,N_6088);
or U8284 (N_8284,N_6035,N_5586);
and U8285 (N_8285,N_2910,N_9);
nor U8286 (N_8286,N_5214,N_2489);
nor U8287 (N_8287,N_523,N_1705);
nand U8288 (N_8288,N_6211,N_721);
or U8289 (N_8289,N_381,N_1664);
nor U8290 (N_8290,N_5804,N_3771);
nand U8291 (N_8291,N_424,N_5754);
nor U8292 (N_8292,N_172,N_4230);
xor U8293 (N_8293,N_4378,N_2740);
or U8294 (N_8294,N_1157,N_5405);
or U8295 (N_8295,N_1508,N_5821);
and U8296 (N_8296,N_4437,N_737);
xor U8297 (N_8297,N_4044,N_4219);
nand U8298 (N_8298,N_1007,N_5440);
nor U8299 (N_8299,N_2242,N_1923);
or U8300 (N_8300,N_2492,N_4276);
xor U8301 (N_8301,N_4693,N_4173);
nor U8302 (N_8302,N_3830,N_5642);
or U8303 (N_8303,N_1307,N_2377);
or U8304 (N_8304,N_2022,N_4981);
or U8305 (N_8305,N_1809,N_1198);
xnor U8306 (N_8306,N_3203,N_6234);
nand U8307 (N_8307,N_1190,N_1818);
and U8308 (N_8308,N_2404,N_3456);
and U8309 (N_8309,N_1693,N_2476);
and U8310 (N_8310,N_5438,N_3350);
and U8311 (N_8311,N_1603,N_1122);
and U8312 (N_8312,N_4537,N_1219);
or U8313 (N_8313,N_740,N_815);
or U8314 (N_8314,N_5040,N_2745);
or U8315 (N_8315,N_1650,N_3729);
or U8316 (N_8316,N_3287,N_5061);
nand U8317 (N_8317,N_587,N_2083);
nor U8318 (N_8318,N_4614,N_1568);
xor U8319 (N_8319,N_176,N_3673);
and U8320 (N_8320,N_1861,N_1993);
xor U8321 (N_8321,N_4031,N_3939);
xor U8322 (N_8322,N_2983,N_3409);
nand U8323 (N_8323,N_1533,N_2525);
xnor U8324 (N_8324,N_1995,N_1205);
nor U8325 (N_8325,N_3610,N_5661);
or U8326 (N_8326,N_1393,N_5358);
nor U8327 (N_8327,N_5520,N_1063);
nand U8328 (N_8328,N_3364,N_1400);
nand U8329 (N_8329,N_4340,N_1057);
and U8330 (N_8330,N_2912,N_5835);
or U8331 (N_8331,N_5563,N_447);
nand U8332 (N_8332,N_3824,N_3597);
and U8333 (N_8333,N_5088,N_2902);
or U8334 (N_8334,N_5385,N_4485);
nor U8335 (N_8335,N_1773,N_1577);
and U8336 (N_8336,N_2330,N_3694);
xnor U8337 (N_8337,N_3900,N_4007);
or U8338 (N_8338,N_2691,N_752);
and U8339 (N_8339,N_4928,N_2485);
nor U8340 (N_8340,N_2231,N_1365);
and U8341 (N_8341,N_591,N_6180);
nand U8342 (N_8342,N_5240,N_2519);
and U8343 (N_8343,N_4925,N_3677);
and U8344 (N_8344,N_1668,N_1625);
and U8345 (N_8345,N_1723,N_2320);
or U8346 (N_8346,N_5890,N_5087);
xnor U8347 (N_8347,N_2481,N_1621);
xor U8348 (N_8348,N_4429,N_751);
and U8349 (N_8349,N_3100,N_2340);
and U8350 (N_8350,N_4119,N_5318);
or U8351 (N_8351,N_6142,N_823);
nand U8352 (N_8352,N_537,N_3540);
and U8353 (N_8353,N_5529,N_3147);
or U8354 (N_8354,N_6083,N_5497);
nor U8355 (N_8355,N_805,N_3707);
and U8356 (N_8356,N_2005,N_1245);
nor U8357 (N_8357,N_1433,N_704);
nand U8358 (N_8358,N_3754,N_1885);
xor U8359 (N_8359,N_3205,N_6007);
and U8360 (N_8360,N_1998,N_6224);
nor U8361 (N_8361,N_316,N_2843);
nor U8362 (N_8362,N_5612,N_2410);
nand U8363 (N_8363,N_6034,N_3187);
or U8364 (N_8364,N_1782,N_6143);
nor U8365 (N_8365,N_5964,N_5752);
nand U8366 (N_8366,N_356,N_650);
nand U8367 (N_8367,N_5274,N_138);
nand U8368 (N_8368,N_1035,N_5584);
and U8369 (N_8369,N_2193,N_4232);
nand U8370 (N_8370,N_4200,N_1864);
nor U8371 (N_8371,N_745,N_1622);
and U8372 (N_8372,N_3137,N_2685);
nor U8373 (N_8373,N_761,N_45);
nor U8374 (N_8374,N_3244,N_1718);
and U8375 (N_8375,N_5806,N_4091);
nand U8376 (N_8376,N_5767,N_1076);
nand U8377 (N_8377,N_2826,N_3725);
nand U8378 (N_8378,N_1278,N_1140);
or U8379 (N_8379,N_3541,N_3815);
and U8380 (N_8380,N_106,N_4752);
and U8381 (N_8381,N_5141,N_3634);
nand U8382 (N_8382,N_5446,N_2584);
nor U8383 (N_8383,N_4688,N_5257);
and U8384 (N_8384,N_987,N_1312);
nand U8385 (N_8385,N_640,N_1043);
nor U8386 (N_8386,N_2402,N_1764);
nand U8387 (N_8387,N_1938,N_2844);
nand U8388 (N_8388,N_2946,N_986);
nand U8389 (N_8389,N_5352,N_5417);
nor U8390 (N_8390,N_4310,N_3913);
nor U8391 (N_8391,N_5706,N_3015);
nand U8392 (N_8392,N_3705,N_3572);
nor U8393 (N_8393,N_3680,N_3624);
or U8394 (N_8394,N_1937,N_1955);
nor U8395 (N_8395,N_2084,N_1350);
or U8396 (N_8396,N_5211,N_5604);
nand U8397 (N_8397,N_4691,N_5470);
xnor U8398 (N_8398,N_3647,N_3209);
nand U8399 (N_8399,N_6093,N_4383);
nand U8400 (N_8400,N_153,N_1048);
or U8401 (N_8401,N_3949,N_906);
nor U8402 (N_8402,N_1686,N_3380);
xor U8403 (N_8403,N_3911,N_2232);
nor U8404 (N_8404,N_5105,N_3306);
xor U8405 (N_8405,N_3919,N_3077);
or U8406 (N_8406,N_5685,N_3143);
nor U8407 (N_8407,N_4881,N_1816);
xor U8408 (N_8408,N_4894,N_3720);
or U8409 (N_8409,N_265,N_1610);
nand U8410 (N_8410,N_5912,N_4842);
nor U8411 (N_8411,N_6155,N_5422);
or U8412 (N_8412,N_2440,N_454);
nor U8413 (N_8413,N_1663,N_425);
nor U8414 (N_8414,N_5173,N_1284);
xnor U8415 (N_8415,N_5344,N_2631);
xnor U8416 (N_8416,N_3171,N_3585);
and U8417 (N_8417,N_5731,N_1859);
nor U8418 (N_8418,N_5233,N_1476);
nand U8419 (N_8419,N_4113,N_664);
or U8420 (N_8420,N_3986,N_6075);
or U8421 (N_8421,N_1851,N_2169);
or U8422 (N_8422,N_4657,N_5442);
nor U8423 (N_8423,N_4674,N_1760);
xor U8424 (N_8424,N_2475,N_3731);
and U8425 (N_8425,N_4315,N_5766);
nand U8426 (N_8426,N_3447,N_5004);
or U8427 (N_8427,N_1397,N_2004);
and U8428 (N_8428,N_4793,N_3204);
nor U8429 (N_8429,N_4987,N_1474);
xor U8430 (N_8430,N_570,N_4779);
xor U8431 (N_8431,N_2417,N_2482);
nand U8432 (N_8432,N_3953,N_2871);
xnor U8433 (N_8433,N_4897,N_5430);
nand U8434 (N_8434,N_2877,N_2172);
and U8435 (N_8435,N_5679,N_3427);
nor U8436 (N_8436,N_4124,N_1337);
or U8437 (N_8437,N_4505,N_552);
or U8438 (N_8438,N_3998,N_5431);
nand U8439 (N_8439,N_4822,N_2730);
nand U8440 (N_8440,N_623,N_1854);
or U8441 (N_8441,N_5632,N_4551);
xnor U8442 (N_8442,N_2576,N_1778);
and U8443 (N_8443,N_4533,N_1262);
nor U8444 (N_8444,N_1908,N_2486);
nor U8445 (N_8445,N_3064,N_856);
xnor U8446 (N_8446,N_3333,N_74);
nor U8447 (N_8447,N_3607,N_6137);
xor U8448 (N_8448,N_5486,N_2447);
xor U8449 (N_8449,N_11,N_2434);
nand U8450 (N_8450,N_1791,N_2302);
nand U8451 (N_8451,N_3880,N_5254);
nand U8452 (N_8452,N_1530,N_907);
nand U8453 (N_8453,N_669,N_4470);
and U8454 (N_8454,N_3475,N_2812);
or U8455 (N_8455,N_4479,N_3629);
and U8456 (N_8456,N_3416,N_3392);
or U8457 (N_8457,N_5350,N_700);
xor U8458 (N_8458,N_4835,N_5332);
xor U8459 (N_8459,N_4147,N_492);
xor U8460 (N_8460,N_1583,N_271);
xor U8461 (N_8461,N_2448,N_5959);
xnor U8462 (N_8462,N_6092,N_6018);
nand U8463 (N_8463,N_785,N_5140);
and U8464 (N_8464,N_3661,N_1763);
and U8465 (N_8465,N_4,N_3437);
nand U8466 (N_8466,N_5583,N_4253);
or U8467 (N_8467,N_2642,N_5868);
nor U8468 (N_8468,N_2321,N_1155);
and U8469 (N_8469,N_941,N_2699);
nand U8470 (N_8470,N_5239,N_4457);
or U8471 (N_8471,N_708,N_1510);
or U8472 (N_8472,N_287,N_1787);
or U8473 (N_8473,N_2263,N_3873);
or U8474 (N_8474,N_1135,N_5445);
nor U8475 (N_8475,N_2559,N_2471);
xor U8476 (N_8476,N_2755,N_2970);
and U8477 (N_8477,N_4142,N_2304);
nor U8478 (N_8478,N_5978,N_2096);
xnor U8479 (N_8479,N_5197,N_4062);
nand U8480 (N_8480,N_4153,N_3180);
nor U8481 (N_8481,N_4748,N_4893);
xor U8482 (N_8482,N_2776,N_4511);
nand U8483 (N_8483,N_3407,N_5789);
nor U8484 (N_8484,N_754,N_6138);
nand U8485 (N_8485,N_4613,N_1226);
and U8486 (N_8486,N_4272,N_841);
or U8487 (N_8487,N_3732,N_3964);
nor U8488 (N_8488,N_1456,N_4638);
and U8489 (N_8489,N_5691,N_2727);
and U8490 (N_8490,N_1152,N_701);
xnor U8491 (N_8491,N_182,N_1320);
nor U8492 (N_8492,N_5212,N_2653);
nor U8493 (N_8493,N_5425,N_4334);
xor U8494 (N_8494,N_1208,N_4043);
nor U8495 (N_8495,N_5537,N_3163);
nand U8496 (N_8496,N_4255,N_5709);
or U8497 (N_8497,N_594,N_3226);
or U8498 (N_8498,N_4912,N_4079);
nor U8499 (N_8499,N_671,N_2659);
nor U8500 (N_8500,N_5660,N_3983);
xor U8501 (N_8501,N_2338,N_2909);
and U8502 (N_8502,N_2339,N_3970);
nor U8503 (N_8503,N_1084,N_2064);
nor U8504 (N_8504,N_3833,N_4527);
or U8505 (N_8505,N_402,N_5958);
nor U8506 (N_8506,N_5626,N_5720);
or U8507 (N_8507,N_6026,N_1878);
or U8508 (N_8508,N_4552,N_2433);
xor U8509 (N_8509,N_5038,N_5353);
or U8510 (N_8510,N_1680,N_3744);
nor U8511 (N_8511,N_309,N_4778);
nand U8512 (N_8512,N_143,N_3752);
and U8513 (N_8513,N_1634,N_2957);
and U8514 (N_8514,N_2551,N_4398);
xor U8515 (N_8515,N_5903,N_2422);
nor U8516 (N_8516,N_6043,N_2927);
nor U8517 (N_8517,N_1651,N_5566);
or U8518 (N_8518,N_3365,N_1425);
or U8519 (N_8519,N_5993,N_1502);
or U8520 (N_8520,N_4228,N_4493);
and U8521 (N_8521,N_939,N_215);
and U8522 (N_8522,N_5678,N_1272);
and U8523 (N_8523,N_2248,N_1807);
nand U8524 (N_8524,N_4339,N_5309);
xor U8525 (N_8525,N_893,N_6084);
nand U8526 (N_8526,N_1560,N_5565);
or U8527 (N_8527,N_1423,N_2581);
or U8528 (N_8528,N_5836,N_2733);
xor U8529 (N_8529,N_891,N_4644);
and U8530 (N_8530,N_3441,N_2234);
or U8531 (N_8531,N_4249,N_3582);
or U8532 (N_8532,N_3230,N_2600);
nand U8533 (N_8533,N_3793,N_1404);
xor U8534 (N_8534,N_3548,N_3442);
nand U8535 (N_8535,N_5224,N_5996);
and U8536 (N_8536,N_70,N_3685);
and U8537 (N_8537,N_2403,N_5238);
and U8538 (N_8538,N_5513,N_203);
xor U8539 (N_8539,N_285,N_2294);
and U8540 (N_8540,N_1519,N_4909);
xor U8541 (N_8541,N_713,N_5342);
or U8542 (N_8542,N_1499,N_2673);
or U8543 (N_8543,N_4303,N_2848);
and U8544 (N_8544,N_1286,N_5528);
and U8545 (N_8545,N_3888,N_1910);
and U8546 (N_8546,N_2470,N_3502);
nand U8547 (N_8547,N_3890,N_118);
and U8548 (N_8548,N_5090,N_1780);
and U8549 (N_8549,N_1355,N_1200);
nand U8550 (N_8550,N_6120,N_5541);
xnor U8551 (N_8551,N_4931,N_3571);
or U8552 (N_8552,N_456,N_1736);
and U8553 (N_8553,N_3360,N_684);
nor U8554 (N_8554,N_6014,N_3116);
nand U8555 (N_8555,N_237,N_6058);
nand U8556 (N_8556,N_1170,N_3212);
nor U8557 (N_8557,N_4964,N_2544);
nand U8558 (N_8558,N_5109,N_6127);
xor U8559 (N_8559,N_1901,N_5837);
and U8560 (N_8560,N_195,N_4144);
or U8561 (N_8561,N_3314,N_5492);
nor U8562 (N_8562,N_1497,N_1212);
and U8563 (N_8563,N_2860,N_4509);
and U8564 (N_8564,N_4057,N_2849);
nand U8565 (N_8565,N_5365,N_1559);
or U8566 (N_8566,N_5799,N_4661);
nor U8567 (N_8567,N_2669,N_4849);
or U8568 (N_8568,N_5481,N_5296);
or U8569 (N_8569,N_2159,N_1318);
xor U8570 (N_8570,N_3491,N_4381);
nor U8571 (N_8571,N_3444,N_2555);
nor U8572 (N_8572,N_4823,N_5526);
nand U8573 (N_8573,N_3870,N_1392);
nand U8574 (N_8574,N_4943,N_5906);
xnor U8575 (N_8575,N_1596,N_1134);
and U8576 (N_8576,N_4832,N_4739);
nor U8577 (N_8577,N_5398,N_1970);
and U8578 (N_8578,N_6141,N_3065);
and U8579 (N_8579,N_1640,N_4150);
nor U8580 (N_8580,N_6076,N_4663);
xnor U8581 (N_8581,N_3332,N_6203);
or U8582 (N_8582,N_2517,N_2348);
nand U8583 (N_8583,N_4308,N_5329);
nor U8584 (N_8584,N_1405,N_479);
xnor U8585 (N_8585,N_3605,N_286);
or U8586 (N_8586,N_1305,N_405);
nor U8587 (N_8587,N_1294,N_2032);
or U8588 (N_8588,N_3506,N_3461);
xor U8589 (N_8589,N_5921,N_2463);
or U8590 (N_8590,N_5782,N_4596);
xor U8591 (N_8591,N_6152,N_5351);
nand U8592 (N_8592,N_449,N_1629);
xor U8593 (N_8593,N_1261,N_5231);
and U8594 (N_8594,N_5624,N_5858);
nor U8595 (N_8595,N_3104,N_913);
and U8596 (N_8596,N_5339,N_2594);
nand U8597 (N_8597,N_4630,N_486);
nor U8598 (N_8598,N_3601,N_2553);
and U8599 (N_8599,N_972,N_5670);
or U8600 (N_8600,N_5023,N_1602);
nand U8601 (N_8601,N_2747,N_5581);
and U8602 (N_8602,N_4546,N_635);
nand U8603 (N_8603,N_2346,N_4385);
xor U8604 (N_8604,N_2267,N_1340);
and U8605 (N_8605,N_226,N_5629);
nand U8606 (N_8606,N_2386,N_2484);
nand U8607 (N_8607,N_2393,N_5184);
nand U8608 (N_8608,N_3369,N_2269);
nor U8609 (N_8609,N_3385,N_5859);
or U8610 (N_8610,N_5598,N_6103);
nor U8611 (N_8611,N_6195,N_1421);
nor U8612 (N_8612,N_5356,N_1635);
xnor U8613 (N_8613,N_5011,N_2798);
or U8614 (N_8614,N_2395,N_2724);
and U8615 (N_8615,N_2811,N_2128);
and U8616 (N_8616,N_6210,N_236);
nor U8617 (N_8617,N_5613,N_4450);
and U8618 (N_8618,N_2212,N_2939);
and U8619 (N_8619,N_2796,N_3734);
nand U8620 (N_8620,N_4712,N_1823);
nor U8621 (N_8621,N_4192,N_4100);
xnor U8622 (N_8622,N_79,N_3923);
and U8623 (N_8623,N_683,N_6029);
nor U8624 (N_8624,N_3818,N_3036);
nand U8625 (N_8625,N_2036,N_6021);
nor U8626 (N_8626,N_3045,N_4176);
xnor U8627 (N_8627,N_5209,N_5162);
nor U8628 (N_8628,N_4211,N_1153);
and U8629 (N_8629,N_3210,N_3281);
nor U8630 (N_8630,N_1376,N_1631);
and U8631 (N_8631,N_2319,N_4786);
xor U8632 (N_8632,N_5991,N_5570);
and U8633 (N_8633,N_233,N_2279);
nor U8634 (N_8634,N_4458,N_2337);
xor U8635 (N_8635,N_663,N_18);
nand U8636 (N_8636,N_5840,N_5864);
or U8637 (N_8637,N_4393,N_49);
or U8638 (N_8638,N_3198,N_1921);
xnor U8639 (N_8639,N_556,N_1064);
xor U8640 (N_8640,N_3261,N_4489);
nor U8641 (N_8641,N_2886,N_4201);
or U8642 (N_8642,N_983,N_1325);
or U8643 (N_8643,N_5968,N_4280);
nor U8644 (N_8644,N_1058,N_580);
xnor U8645 (N_8645,N_5148,N_3525);
and U8646 (N_8646,N_2990,N_4474);
and U8647 (N_8647,N_4775,N_860);
nand U8648 (N_8648,N_649,N_343);
nand U8649 (N_8649,N_4343,N_1877);
nor U8650 (N_8650,N_2307,N_5862);
nor U8651 (N_8651,N_3037,N_5226);
and U8652 (N_8652,N_6036,N_825);
nor U8653 (N_8653,N_5416,N_5746);
nor U8654 (N_8654,N_3128,N_4002);
xor U8655 (N_8655,N_710,N_1346);
and U8656 (N_8656,N_6104,N_4753);
nor U8657 (N_8657,N_187,N_5553);
and U8658 (N_8658,N_6108,N_3653);
nor U8659 (N_8659,N_2725,N_1714);
xnor U8660 (N_8660,N_5315,N_3338);
nor U8661 (N_8661,N_1214,N_2326);
nor U8662 (N_8662,N_5710,N_5855);
nor U8663 (N_8663,N_3860,N_6226);
nor U8664 (N_8664,N_6017,N_1895);
nor U8665 (N_8665,N_4311,N_926);
or U8666 (N_8666,N_1524,N_2981);
and U8667 (N_8667,N_1018,N_1866);
and U8668 (N_8668,N_4781,N_4133);
nor U8669 (N_8669,N_404,N_5432);
and U8670 (N_8670,N_3738,N_786);
nor U8671 (N_8671,N_2161,N_4556);
and U8672 (N_8672,N_2474,N_4028);
or U8673 (N_8673,N_2158,N_173);
nor U8674 (N_8674,N_4554,N_6139);
nand U8675 (N_8675,N_4998,N_5227);
nand U8676 (N_8676,N_1593,N_5370);
nor U8677 (N_8677,N_3429,N_5763);
xor U8678 (N_8678,N_4061,N_1283);
and U8679 (N_8679,N_3296,N_3082);
or U8680 (N_8680,N_3972,N_2041);
and U8681 (N_8681,N_3010,N_1250);
or U8682 (N_8682,N_1185,N_1873);
and U8683 (N_8683,N_2668,N_5808);
and U8684 (N_8684,N_870,N_5418);
or U8685 (N_8685,N_3564,N_1592);
or U8686 (N_8686,N_4954,N_2993);
nor U8687 (N_8687,N_4540,N_2906);
xor U8688 (N_8688,N_584,N_1769);
and U8689 (N_8689,N_194,N_2945);
and U8690 (N_8690,N_4746,N_760);
or U8691 (N_8691,N_1072,N_3083);
xnor U8692 (N_8692,N_4355,N_3014);
xnor U8693 (N_8693,N_5054,N_4141);
and U8694 (N_8694,N_5986,N_5987);
nor U8695 (N_8695,N_354,N_240);
xor U8696 (N_8696,N_2345,N_1422);
nand U8697 (N_8697,N_3330,N_3257);
nor U8698 (N_8698,N_4329,N_5973);
or U8699 (N_8699,N_2542,N_6003);
nor U8700 (N_8700,N_4839,N_2327);
xnor U8701 (N_8701,N_4707,N_5876);
or U8702 (N_8702,N_810,N_2210);
nor U8703 (N_8703,N_1317,N_971);
and U8704 (N_8704,N_2674,N_4241);
or U8705 (N_8705,N_6113,N_2573);
or U8706 (N_8706,N_5669,N_5918);
nand U8707 (N_8707,N_595,N_605);
and U8708 (N_8708,N_4583,N_3093);
nor U8709 (N_8709,N_3569,N_5957);
nor U8710 (N_8710,N_637,N_2151);
and U8711 (N_8711,N_3561,N_2055);
or U8712 (N_8712,N_2609,N_6123);
xnor U8713 (N_8713,N_566,N_725);
and U8714 (N_8714,N_3186,N_1189);
and U8715 (N_8715,N_5218,N_72);
or U8716 (N_8716,N_3878,N_3907);
xor U8717 (N_8717,N_5701,N_5156);
xor U8718 (N_8718,N_1833,N_3512);
nor U8719 (N_8719,N_2182,N_4924);
and U8720 (N_8720,N_5625,N_1512);
and U8721 (N_8721,N_228,N_3982);
or U8722 (N_8722,N_4172,N_2148);
and U8723 (N_8723,N_4401,N_4816);
xnor U8724 (N_8724,N_1846,N_43);
and U8725 (N_8725,N_3604,N_1302);
and U8726 (N_8726,N_714,N_639);
or U8727 (N_8727,N_4730,N_341);
nor U8728 (N_8728,N_3641,N_1408);
nor U8729 (N_8729,N_3303,N_1803);
or U8730 (N_8730,N_3622,N_2547);
nand U8731 (N_8731,N_5177,N_1293);
or U8732 (N_8732,N_1537,N_5688);
and U8733 (N_8733,N_2762,N_4268);
xor U8734 (N_8734,N_3208,N_3378);
nor U8735 (N_8735,N_4896,N_3683);
xnor U8736 (N_8736,N_1093,N_3794);
and U8737 (N_8737,N_1028,N_3989);
xnor U8738 (N_8738,N_325,N_422);
or U8739 (N_8739,N_3465,N_3351);
or U8740 (N_8740,N_4025,N_3584);
or U8741 (N_8741,N_1193,N_2334);
or U8742 (N_8742,N_5328,N_144);
or U8743 (N_8743,N_980,N_1174);
nor U8744 (N_8744,N_2834,N_3704);
nor U8745 (N_8745,N_4327,N_2516);
nand U8746 (N_8746,N_5161,N_5394);
or U8747 (N_8747,N_1784,N_2806);
nand U8748 (N_8748,N_3659,N_1749);
and U8749 (N_8749,N_5077,N_5249);
nor U8750 (N_8750,N_2439,N_1253);
xor U8751 (N_8751,N_5193,N_4476);
or U8752 (N_8752,N_4698,N_1127);
nor U8753 (N_8753,N_540,N_3808);
or U8754 (N_8754,N_3038,N_2082);
and U8755 (N_8755,N_4491,N_4501);
and U8756 (N_8756,N_1119,N_4492);
xor U8757 (N_8757,N_2456,N_5400);
or U8758 (N_8758,N_5946,N_2980);
nand U8759 (N_8759,N_5634,N_3115);
and U8760 (N_8760,N_4829,N_380);
nand U8761 (N_8761,N_5933,N_4725);
nand U8762 (N_8762,N_455,N_3462);
nor U8763 (N_8763,N_1142,N_3052);
and U8764 (N_8764,N_2416,N_1967);
nor U8765 (N_8765,N_4961,N_5590);
nand U8766 (N_8766,N_1544,N_935);
nand U8767 (N_8767,N_3481,N_5645);
nor U8768 (N_8768,N_4851,N_505);
xnor U8769 (N_8769,N_213,N_4364);
xor U8770 (N_8770,N_2282,N_1156);
xor U8771 (N_8771,N_4946,N_6095);
or U8772 (N_8772,N_5585,N_634);
nand U8773 (N_8773,N_1281,N_818);
nand U8774 (N_8774,N_1188,N_1793);
nand U8775 (N_8775,N_5280,N_5915);
xor U8776 (N_8776,N_1437,N_909);
nor U8777 (N_8777,N_2692,N_3199);
nor U8778 (N_8778,N_1067,N_2399);
nor U8779 (N_8779,N_3242,N_3067);
nand U8780 (N_8780,N_1954,N_373);
or U8781 (N_8781,N_5689,N_5096);
and U8782 (N_8782,N_4151,N_798);
xnor U8783 (N_8783,N_3231,N_4653);
nand U8784 (N_8784,N_5285,N_872);
nand U8785 (N_8785,N_1964,N_1299);
or U8786 (N_8786,N_2852,N_2760);
nand U8787 (N_8787,N_4134,N_5572);
xor U8788 (N_8788,N_84,N_1366);
or U8789 (N_8789,N_91,N_4021);
and U8790 (N_8790,N_367,N_2537);
nand U8791 (N_8791,N_2374,N_2075);
or U8792 (N_8792,N_6225,N_1571);
or U8793 (N_8793,N_1888,N_5680);
nand U8794 (N_8794,N_1201,N_2613);
nand U8795 (N_8795,N_1525,N_1832);
nand U8796 (N_8796,N_693,N_1754);
nand U8797 (N_8797,N_134,N_2188);
xnor U8798 (N_8798,N_1735,N_4854);
xnor U8799 (N_8799,N_1463,N_3726);
nand U8800 (N_8800,N_1252,N_5602);
nand U8801 (N_8801,N_5477,N_4864);
nand U8802 (N_8802,N_1907,N_5936);
and U8803 (N_8803,N_4722,N_364);
nor U8804 (N_8804,N_6208,N_5801);
xor U8805 (N_8805,N_2144,N_2052);
or U8806 (N_8806,N_1597,N_4430);
xor U8807 (N_8807,N_2892,N_1731);
nand U8808 (N_8808,N_990,N_4066);
nor U8809 (N_8809,N_5439,N_2494);
nor U8810 (N_8810,N_3648,N_2938);
and U8811 (N_8811,N_4009,N_2605);
nand U8812 (N_8812,N_5491,N_5012);
nor U8813 (N_8813,N_3708,N_4443);
or U8814 (N_8814,N_1987,N_3176);
xnor U8815 (N_8815,N_5615,N_1358);
nor U8816 (N_8816,N_2950,N_4637);
nor U8817 (N_8817,N_5205,N_2870);
and U8818 (N_8818,N_1522,N_431);
nand U8819 (N_8819,N_3426,N_4365);
xnor U8820 (N_8820,N_958,N_3182);
nor U8821 (N_8821,N_866,N_5269);
xnor U8822 (N_8822,N_3869,N_4252);
xnor U8823 (N_8823,N_2943,N_4312);
xor U8824 (N_8824,N_4679,N_460);
xor U8825 (N_8825,N_5815,N_2930);
or U8826 (N_8826,N_597,N_3976);
and U8827 (N_8827,N_5830,N_2341);
and U8828 (N_8828,N_3910,N_2777);
nor U8829 (N_8829,N_2606,N_4156);
nor U8830 (N_8830,N_3639,N_5694);
or U8831 (N_8831,N_5623,N_2766);
xor U8832 (N_8832,N_98,N_1574);
xnor U8833 (N_8833,N_4762,N_2793);
or U8834 (N_8834,N_4279,N_104);
nor U8835 (N_8835,N_688,N_6134);
nand U8836 (N_8836,N_1712,N_1788);
nand U8837 (N_8837,N_2078,N_150);
and U8838 (N_8838,N_930,N_3507);
nand U8839 (N_8839,N_3161,N_5210);
nor U8840 (N_8840,N_1804,N_5982);
or U8841 (N_8841,N_6081,N_363);
nor U8842 (N_8842,N_6051,N_3798);
and U8843 (N_8843,N_4932,N_3484);
or U8844 (N_8844,N_5391,N_2121);
and U8845 (N_8845,N_2511,N_3467);
xnor U8846 (N_8846,N_1129,N_4521);
xnor U8847 (N_8847,N_1347,N_3387);
nand U8848 (N_8848,N_4578,N_288);
xor U8849 (N_8849,N_2029,N_2261);
nand U8850 (N_8850,N_859,N_1922);
xor U8851 (N_8851,N_1257,N_828);
or U8852 (N_8852,N_654,N_5089);
and U8853 (N_8853,N_5538,N_5888);
and U8854 (N_8854,N_4525,N_290);
and U8855 (N_8855,N_3935,N_2858);
or U8856 (N_8856,N_4800,N_1633);
or U8857 (N_8857,N_1470,N_1096);
xnor U8858 (N_8858,N_2432,N_2630);
and U8859 (N_8859,N_5530,N_24);
and U8860 (N_8860,N_3453,N_2518);
xor U8861 (N_8861,N_5654,N_3905);
nor U8862 (N_8862,N_2926,N_3268);
nor U8863 (N_8863,N_2865,N_789);
nor U8864 (N_8864,N_2258,N_4936);
nor U8865 (N_8865,N_542,N_2819);
nand U8866 (N_8866,N_5067,N_304);
nand U8867 (N_8867,N_5856,N_5409);
or U8868 (N_8868,N_2982,N_1357);
or U8869 (N_8869,N_1276,N_3588);
xor U8870 (N_8870,N_1239,N_6219);
or U8871 (N_8871,N_3496,N_3255);
or U8872 (N_8872,N_4167,N_543);
and U8873 (N_8873,N_2300,N_4338);
nor U8874 (N_8874,N_4260,N_4838);
xor U8875 (N_8875,N_747,N_4945);
nor U8876 (N_8876,N_2775,N_1843);
and U8877 (N_8877,N_4094,N_2709);
or U8878 (N_8878,N_5402,N_12);
nand U8879 (N_8879,N_2031,N_565);
xnor U8880 (N_8880,N_4518,N_5589);
nor U8881 (N_8881,N_5448,N_5181);
xnor U8882 (N_8882,N_3173,N_2284);
xor U8883 (N_8883,N_3384,N_3423);
and U8884 (N_8884,N_3672,N_1102);
xnor U8885 (N_8885,N_3240,N_2264);
or U8886 (N_8886,N_1331,N_5539);
and U8887 (N_8887,N_3713,N_274);
nand U8888 (N_8888,N_3696,N_1554);
and U8889 (N_8889,N_3003,N_5895);
xnor U8890 (N_8890,N_5812,N_6015);
nor U8891 (N_8891,N_3134,N_192);
nor U8892 (N_8892,N_131,N_3321);
nor U8893 (N_8893,N_2785,N_5742);
nor U8894 (N_8894,N_457,N_1628);
or U8895 (N_8895,N_3080,N_2335);
nand U8896 (N_8896,N_4833,N_5532);
nand U8897 (N_8897,N_2449,N_3026);
nand U8898 (N_8898,N_6,N_1659);
or U8899 (N_8899,N_473,N_877);
xnor U8900 (N_8900,N_6008,N_3184);
and U8901 (N_8901,N_895,N_3183);
nand U8902 (N_8902,N_755,N_4780);
nor U8903 (N_8903,N_2129,N_4984);
or U8904 (N_8904,N_398,N_4935);
and U8905 (N_8905,N_2637,N_4374);
xnor U8906 (N_8906,N_4852,N_4465);
and U8907 (N_8907,N_3646,N_3343);
or U8908 (N_8908,N_3786,N_50);
xor U8909 (N_8909,N_4650,N_3070);
nor U8910 (N_8910,N_1486,N_313);
nor U8911 (N_8911,N_193,N_4645);
nor U8912 (N_8912,N_1409,N_653);
nor U8913 (N_8913,N_5757,N_526);
or U8914 (N_8914,N_266,N_2445);
xnor U8915 (N_8915,N_3282,N_1344);
nor U8916 (N_8916,N_1118,N_6122);
nor U8917 (N_8917,N_871,N_4495);
or U8918 (N_8918,N_6065,N_2310);
or U8919 (N_8919,N_2243,N_3969);
nand U8920 (N_8920,N_2245,N_2768);
or U8921 (N_8921,N_2603,N_4600);
or U8922 (N_8922,N_3477,N_1511);
or U8923 (N_8923,N_4858,N_3021);
nand U8924 (N_8924,N_4486,N_3630);
nor U8925 (N_8925,N_2039,N_496);
xor U8926 (N_8926,N_736,N_4326);
nand U8927 (N_8927,N_4634,N_3107);
xnor U8928 (N_8928,N_6067,N_2164);
and U8929 (N_8929,N_1314,N_5628);
or U8930 (N_8930,N_5182,N_3528);
and U8931 (N_8931,N_3792,N_5117);
and U8932 (N_8932,N_5034,N_5024);
nand U8933 (N_8933,N_4827,N_807);
or U8934 (N_8934,N_4090,N_3024);
and U8935 (N_8935,N_3452,N_5514);
nand U8936 (N_8936,N_6124,N_5723);
nand U8937 (N_8937,N_5062,N_1639);
xor U8938 (N_8938,N_1774,N_3307);
and U8939 (N_8939,N_5571,N_3984);
nor U8940 (N_8940,N_2994,N_4335);
xor U8941 (N_8941,N_3931,N_1865);
and U8942 (N_8942,N_743,N_407);
xor U8943 (N_8943,N_1643,N_5375);
nor U8944 (N_8944,N_3434,N_3509);
and U8945 (N_8945,N_1716,N_3952);
xnor U8946 (N_8946,N_2505,N_5279);
nor U8947 (N_8947,N_5414,N_1494);
and U8948 (N_8948,N_5190,N_5803);
and U8949 (N_8949,N_783,N_951);
and U8950 (N_8950,N_5956,N_397);
or U8951 (N_8951,N_3567,N_4442);
and U8952 (N_8952,N_4171,N_5003);
or U8953 (N_8953,N_403,N_152);
nor U8954 (N_8954,N_5810,N_1022);
nor U8955 (N_8955,N_2998,N_695);
and U8956 (N_8956,N_160,N_4480);
nand U8957 (N_8957,N_2790,N_1489);
and U8958 (N_8958,N_2893,N_3643);
nor U8959 (N_8959,N_1148,N_2560);
xor U8960 (N_8960,N_146,N_15);
nor U8961 (N_8961,N_5147,N_4160);
nor U8962 (N_8962,N_1506,N_5550);
and U8963 (N_8963,N_19,N_1912);
and U8964 (N_8964,N_2145,N_5778);
nor U8965 (N_8965,N_3576,N_5703);
xnor U8966 (N_8966,N_1056,N_5075);
xor U8967 (N_8967,N_4063,N_5372);
or U8968 (N_8968,N_608,N_78);
or U8969 (N_8969,N_1844,N_1806);
nor U8970 (N_8970,N_3778,N_1342);
nand U8971 (N_8971,N_1078,N_2667);
or U8972 (N_8972,N_3101,N_4717);
nand U8973 (N_8973,N_3832,N_5337);
and U8974 (N_8974,N_2889,N_3058);
nand U8975 (N_8975,N_3545,N_814);
and U8976 (N_8976,N_2177,N_5820);
or U8977 (N_8977,N_5357,N_2690);
nand U8978 (N_8978,N_1496,N_4749);
xnor U8979 (N_8979,N_1452,N_5456);
nand U8980 (N_8980,N_3747,N_1309);
and U8981 (N_8981,N_1786,N_3487);
and U8982 (N_8982,N_123,N_5126);
nand U8983 (N_8983,N_322,N_5429);
or U8984 (N_8984,N_3600,N_4857);
xor U8985 (N_8985,N_4670,N_914);
or U8986 (N_8986,N_2767,N_336);
nand U8987 (N_8987,N_2627,N_6249);
nand U8988 (N_8988,N_2135,N_2016);
nand U8989 (N_8989,N_2583,N_3628);
and U8990 (N_8990,N_2532,N_2622);
nor U8991 (N_8991,N_1466,N_1906);
or U8992 (N_8992,N_6038,N_61);
xor U8993 (N_8993,N_4198,N_5842);
xor U8994 (N_8994,N_3831,N_1841);
xor U8995 (N_8995,N_1920,N_1326);
nor U8996 (N_8996,N_300,N_1696);
nor U8997 (N_8997,N_2202,N_5183);
xnor U8998 (N_8998,N_1379,N_4901);
xnor U8999 (N_8999,N_1935,N_4262);
and U9000 (N_9000,N_346,N_3483);
nor U9001 (N_9001,N_2515,N_1269);
nand U9002 (N_9002,N_4030,N_1471);
nor U9003 (N_9003,N_4721,N_127);
xnor U9004 (N_9004,N_2863,N_5151);
nand U9005 (N_9005,N_2365,N_3057);
xnor U9006 (N_9006,N_1688,N_3811);
nor U9007 (N_9007,N_5740,N_3784);
nand U9008 (N_9008,N_536,N_1911);
nor U9009 (N_9009,N_5499,N_6154);
xnor U9010 (N_9010,N_2009,N_4396);
nand U9011 (N_9011,N_482,N_6144);
and U9012 (N_9012,N_1880,N_4905);
xnor U9013 (N_9013,N_1531,N_3046);
nand U9014 (N_9014,N_5774,N_5849);
or U9015 (N_9015,N_4286,N_1848);
or U9016 (N_9016,N_3069,N_5452);
nor U9017 (N_9017,N_4561,N_6236);
xnor U9018 (N_9018,N_985,N_3414);
and U9019 (N_9019,N_3578,N_547);
nor U9020 (N_9020,N_4519,N_1829);
and U9021 (N_9021,N_890,N_4926);
or U9022 (N_9022,N_2675,N_6111);
nor U9023 (N_9023,N_295,N_4766);
nand U9024 (N_9024,N_4164,N_4915);
nor U9025 (N_9025,N_179,N_463);
and U9026 (N_9026,N_592,N_4431);
and U9027 (N_9027,N_1123,N_4876);
nor U9028 (N_9028,N_5601,N_4792);
or U9029 (N_9029,N_5900,N_1453);
nand U9030 (N_9030,N_790,N_2524);
and U9031 (N_9031,N_4735,N_136);
nor U9032 (N_9032,N_2196,N_2705);
xnor U9033 (N_9033,N_345,N_5667);
xor U9034 (N_9034,N_1213,N_1147);
nand U9035 (N_9035,N_974,N_4756);
nor U9036 (N_9036,N_2531,N_2457);
xor U9037 (N_9037,N_4301,N_3841);
nand U9038 (N_9038,N_5913,N_4834);
nor U9039 (N_9039,N_1758,N_1925);
or U9040 (N_9040,N_360,N_417);
or U9041 (N_9041,N_3511,N_1584);
and U9042 (N_9042,N_430,N_3733);
nand U9043 (N_9043,N_1330,N_2364);
and U9044 (N_9044,N_1699,N_1646);
nor U9045 (N_9045,N_4069,N_3227);
and U9046 (N_9046,N_1540,N_6178);
and U9047 (N_9047,N_1385,N_2280);
nand U9048 (N_9048,N_3195,N_1981);
and U9049 (N_9049,N_1966,N_2721);
or U9050 (N_9050,N_5195,N_5556);
and U9051 (N_9051,N_5540,N_2723);
xor U9052 (N_9052,N_4494,N_502);
nor U9053 (N_9053,N_1990,N_5049);
or U9054 (N_9054,N_3413,N_4332);
nand U9055 (N_9055,N_4611,N_6087);
or U9056 (N_9056,N_3611,N_5649);
nor U9057 (N_9057,N_5524,N_1838);
xor U9058 (N_9058,N_2056,N_201);
xnor U9059 (N_9059,N_706,N_4318);
and U9060 (N_9060,N_5114,N_3219);
nand U9061 (N_9061,N_1648,N_4865);
nand U9062 (N_9062,N_5346,N_5095);
and U9063 (N_9063,N_4155,N_5019);
nand U9064 (N_9064,N_6246,N_1444);
xnor U9065 (N_9065,N_4415,N_5549);
nor U9066 (N_9066,N_2557,N_4250);
or U9067 (N_9067,N_2430,N_507);
and U9068 (N_9068,N_2443,N_6212);
or U9069 (N_9069,N_5768,N_1871);
or U9070 (N_9070,N_1080,N_949);
and U9071 (N_9071,N_5726,N_5595);
xnor U9072 (N_9072,N_1074,N_2246);
or U9073 (N_9073,N_3678,N_2850);
and U9074 (N_9074,N_4078,N_3565);
and U9075 (N_9075,N_4763,N_2835);
xnor U9076 (N_9076,N_3927,N_4379);
or U9077 (N_9077,N_5268,N_5308);
or U9078 (N_9078,N_349,N_2472);
and U9079 (N_9079,N_145,N_5885);
nor U9080 (N_9080,N_4994,N_3419);
nand U9081 (N_9081,N_3549,N_250);
xor U9082 (N_9082,N_4970,N_438);
nand U9083 (N_9083,N_469,N_3655);
and U9084 (N_9084,N_4148,N_5434);
and U9085 (N_9085,N_2241,N_3076);
and U9086 (N_9086,N_214,N_4247);
or U9087 (N_9087,N_4187,N_3965);
and U9088 (N_9088,N_3062,N_5489);
xnor U9089 (N_9089,N_369,N_63);
and U9090 (N_9090,N_5362,N_3755);
xor U9091 (N_9091,N_2425,N_3922);
or U9092 (N_9092,N_6059,N_2614);
nor U9093 (N_9093,N_4054,N_1488);
or U9094 (N_9094,N_5102,N_200);
or U9095 (N_9095,N_2313,N_5361);
nor U9096 (N_9096,N_3485,N_76);
xor U9097 (N_9097,N_2047,N_6248);
and U9098 (N_9098,N_5705,N_4808);
nor U9099 (N_9099,N_212,N_5517);
nand U9100 (N_9100,N_5467,N_4716);
xnor U9101 (N_9101,N_5548,N_816);
nor U9102 (N_9102,N_1837,N_2362);
xnor U9103 (N_9103,N_1903,N_3675);
nand U9104 (N_9104,N_5910,N_1465);
and U9105 (N_9105,N_665,N_5033);
or U9106 (N_9106,N_6006,N_1927);
nor U9107 (N_9107,N_5574,N_3777);
nand U9108 (N_9108,N_768,N_1503);
xor U9109 (N_9109,N_2847,N_5225);
nor U9110 (N_9110,N_2134,N_628);
and U9111 (N_9111,N_22,N_1411);
xnor U9112 (N_9112,N_4363,N_2253);
xor U9113 (N_9113,N_1834,N_399);
xnor U9114 (N_9114,N_3214,N_660);
xnor U9115 (N_9115,N_5777,N_2880);
and U9116 (N_9116,N_827,N_38);
nand U9117 (N_9117,N_2102,N_3479);
nor U9118 (N_9118,N_6116,N_468);
xnor U9119 (N_9119,N_5153,N_2828);
or U9120 (N_9120,N_5324,N_4345);
nand U9121 (N_9121,N_3727,N_5576);
nor U9122 (N_9122,N_5564,N_471);
nand U9123 (N_9123,N_5039,N_3376);
nand U9124 (N_9124,N_2249,N_5103);
nand U9125 (N_9125,N_2226,N_571);
nor U9126 (N_9126,N_804,N_2178);
xor U9127 (N_9127,N_3337,N_5551);
nand U9128 (N_9128,N_1141,N_5420);
xor U9129 (N_9129,N_5237,N_6157);
nor U9130 (N_9130,N_1798,N_915);
nand U9131 (N_9131,N_1614,N_2890);
nand U9132 (N_9132,N_4639,N_1461);
and U9133 (N_9133,N_973,N_3071);
nor U9134 (N_9134,N_5397,N_4236);
xnor U9135 (N_9135,N_1225,N_4027);
nor U9136 (N_9136,N_257,N_3308);
and U9137 (N_9137,N_3473,N_211);
or U9138 (N_9138,N_1947,N_5216);
or U9139 (N_9139,N_4029,N_1745);
xnor U9140 (N_9140,N_1551,N_3757);
xor U9141 (N_9141,N_3810,N_3066);
and U9142 (N_9142,N_3454,N_2271);
nand U9143 (N_9143,N_3517,N_6022);
xor U9144 (N_9144,N_4123,N_2529);
or U9145 (N_9145,N_4522,N_4185);
or U9146 (N_9146,N_1529,N_4261);
or U9147 (N_9147,N_5755,N_1223);
nor U9148 (N_9148,N_4831,N_4135);
or U9149 (N_9149,N_5716,N_882);
nand U9150 (N_9150,N_4115,N_2424);
or U9151 (N_9151,N_548,N_2509);
and U9152 (N_9152,N_3681,N_239);
xnor U9153 (N_9153,N_4391,N_612);
xnor U9154 (N_9154,N_4640,N_2661);
xnor U9155 (N_9155,N_3449,N_794);
or U9156 (N_9156,N_2168,N_2677);
and U9157 (N_9157,N_3740,N_3850);
nand U9158 (N_9158,N_2105,N_1586);
xor U9159 (N_9159,N_5355,N_4460);
xor U9160 (N_9160,N_528,N_128);
xor U9161 (N_9161,N_1171,N_5641);
xnor U9162 (N_9162,N_928,N_2615);
nand U9163 (N_9163,N_509,N_3087);
nor U9164 (N_9164,N_728,N_2089);
and U9165 (N_9165,N_2955,N_1310);
xor U9166 (N_9166,N_5899,N_4266);
nor U9167 (N_9167,N_1457,N_3121);
or U9168 (N_9168,N_1484,N_3770);
nand U9169 (N_9169,N_4608,N_5384);
nand U9170 (N_9170,N_5823,N_4405);
and U9171 (N_9171,N_5606,N_2751);
or U9172 (N_9172,N_5818,N_3318);
nor U9173 (N_9173,N_5116,N_4306);
nand U9174 (N_9174,N_3785,N_4652);
nor U9175 (N_9175,N_3468,N_3947);
nand U9176 (N_9176,N_230,N_2757);
and U9177 (N_9177,N_6132,N_4278);
nor U9178 (N_9178,N_4517,N_1163);
or U9179 (N_9179,N_4697,N_5882);
or U9180 (N_9180,N_3670,N_2783);
nor U9181 (N_9181,N_2197,N_4297);
nor U9182 (N_9182,N_2223,N_3292);
xnor U9183 (N_9183,N_2959,N_875);
nor U9184 (N_9184,N_1145,N_4049);
xnor U9185 (N_9185,N_5848,N_503);
and U9186 (N_9186,N_3175,N_6204);
nor U9187 (N_9187,N_3790,N_3438);
or U9188 (N_9188,N_3366,N_6233);
or U9189 (N_9189,N_6145,N_4947);
or U9190 (N_9190,N_4503,N_3156);
or U9191 (N_9191,N_3595,N_4413);
and U9192 (N_9192,N_3617,N_4810);
or U9193 (N_9193,N_1356,N_5784);
xor U9194 (N_9194,N_801,N_2412);
xnor U9195 (N_9195,N_5832,N_5313);
xor U9196 (N_9196,N_156,N_5130);
and U9197 (N_9197,N_3573,N_4496);
xor U9198 (N_9198,N_1353,N_5592);
nand U9199 (N_9199,N_3443,N_3243);
nor U9200 (N_9200,N_4784,N_4239);
nor U9201 (N_9201,N_5605,N_6176);
xor U9202 (N_9202,N_229,N_4146);
nor U9203 (N_9203,N_4772,N_687);
xnor U9204 (N_9204,N_5415,N_2413);
nor U9205 (N_9205,N_5199,N_4566);
nand U9206 (N_9206,N_5131,N_4843);
nand U9207 (N_9207,N_3765,N_4783);
xnor U9208 (N_9208,N_2473,N_676);
and U9209 (N_9209,N_1131,N_1019);
nand U9210 (N_9210,N_3533,N_6080);
nand U9211 (N_9211,N_5258,N_5518);
nor U9212 (N_9212,N_576,N_4953);
and U9213 (N_9213,N_5617,N_1726);
and U9214 (N_9214,N_3320,N_1221);
or U9215 (N_9215,N_3267,N_2538);
xnor U9216 (N_9216,N_4157,N_470);
xor U9217 (N_9217,N_2988,N_551);
nor U9218 (N_9218,N_529,N_936);
nor U9219 (N_9219,N_4701,N_6039);
and U9220 (N_9220,N_2947,N_1526);
and U9221 (N_9221,N_5137,N_4384);
nand U9222 (N_9222,N_4963,N_3132);
xor U9223 (N_9223,N_1323,N_51);
and U9224 (N_9224,N_2832,N_5713);
or U9225 (N_9225,N_2772,N_3712);
and U9226 (N_9226,N_4095,N_5839);
nor U9227 (N_9227,N_1814,N_5286);
nand U9228 (N_9228,N_3265,N_3310);
nand U9229 (N_9229,N_1623,N_6105);
xnor U9230 (N_9230,N_3688,N_3237);
xor U9231 (N_9231,N_115,N_3110);
nor U9232 (N_9232,N_3049,N_2831);
xor U9233 (N_9233,N_3557,N_1515);
xnor U9234 (N_9234,N_4056,N_443);
nand U9235 (N_9235,N_2977,N_1267);
nand U9236 (N_9236,N_2915,N_2183);
nand U9237 (N_9237,N_2527,N_5314);
nand U9238 (N_9238,N_2451,N_1872);
xor U9239 (N_9239,N_5750,N_2563);
or U9240 (N_9240,N_5525,N_3490);
xor U9241 (N_9241,N_689,N_4973);
or U9242 (N_9242,N_1390,N_2941);
nor U9243 (N_9243,N_2037,N_1857);
or U9244 (N_9244,N_33,N_3735);
nor U9245 (N_9245,N_1075,N_326);
or U9246 (N_9246,N_4605,N_6197);
or U9247 (N_9247,N_3568,N_34);
and U9248 (N_9248,N_2658,N_3691);
xnor U9249 (N_9249,N_1665,N_5245);
nand U9250 (N_9250,N_5734,N_4910);
xor U9251 (N_9251,N_3566,N_5366);
or U9252 (N_9252,N_5002,N_1619);
and U9253 (N_9253,N_3717,N_1883);
and U9254 (N_9254,N_3546,N_2043);
and U9255 (N_9255,N_3945,N_779);
or U9256 (N_9256,N_3439,N_729);
nand U9257 (N_9257,N_4899,N_270);
nor U9258 (N_9258,N_2117,N_154);
or U9259 (N_9259,N_5500,N_5028);
xnor U9260 (N_9260,N_3823,N_5166);
nor U9261 (N_9261,N_234,N_731);
nor U9262 (N_9262,N_809,N_1027);
or U9263 (N_9263,N_712,N_6024);
nor U9264 (N_9264,N_2233,N_5251);
xor U9265 (N_9265,N_1538,N_5935);
xor U9266 (N_9266,N_450,N_2623);
nand U9267 (N_9267,N_2985,N_5971);
xnor U9268 (N_9268,N_3759,N_5621);
nand U9269 (N_9269,N_272,N_3660);
or U9270 (N_9270,N_4884,N_5099);
or U9271 (N_9271,N_4368,N_2822);
nand U9272 (N_9272,N_4348,N_273);
and U9273 (N_9273,N_2363,N_2854);
nor U9274 (N_9274,N_4812,N_5276);
or U9275 (N_9275,N_3724,N_4206);
xor U9276 (N_9276,N_3768,N_5165);
or U9277 (N_9277,N_5005,N_1569);
xor U9278 (N_9278,N_378,N_6031);
or U9279 (N_9279,N_5412,N_1729);
nand U9280 (N_9280,N_5994,N_5135);
and U9281 (N_9281,N_3289,N_1997);
or U9282 (N_9282,N_4039,N_4060);
xor U9283 (N_9283,N_3235,N_863);
nor U9284 (N_9284,N_2322,N_3769);
nand U9285 (N_9285,N_6074,N_6121);
nor U9286 (N_9286,N_2546,N_884);
xnor U9287 (N_9287,N_821,N_4765);
nor U9288 (N_9288,N_560,N_5435);
nor U9289 (N_9289,N_5484,N_2759);
xnor U9290 (N_9290,N_3845,N_869);
nand U9291 (N_9291,N_967,N_1004);
nor U9292 (N_9292,N_5522,N_1601);
xnor U9293 (N_9293,N_3859,N_1151);
and U9294 (N_9294,N_3899,N_633);
and U9295 (N_9295,N_518,N_5056);
or U9296 (N_9296,N_4488,N_5652);
nor U9297 (N_9297,N_111,N_4154);
xnor U9298 (N_9298,N_897,N_1507);
or U9299 (N_9299,N_3313,N_2830);
or U9300 (N_9300,N_2409,N_1582);
xor U9301 (N_9301,N_3579,N_3157);
nor U9302 (N_9302,N_2176,N_2803);
or U9303 (N_9303,N_889,N_5122);
nand U9304 (N_9304,N_5798,N_2610);
nor U9305 (N_9305,N_4001,N_6042);
nand U9306 (N_9306,N_3954,N_1447);
and U9307 (N_9307,N_4137,N_5230);
nand U9308 (N_9308,N_4888,N_6060);
or U9309 (N_9309,N_820,N_2278);
and U9310 (N_9310,N_475,N_3742);
nor U9311 (N_9311,N_2936,N_5259);
nor U9312 (N_9312,N_5928,N_4825);
nand U9313 (N_9313,N_4462,N_101);
or U9314 (N_9314,N_3106,N_65);
or U9315 (N_9315,N_5059,N_694);
or U9316 (N_9316,N_1991,N_1839);
or U9317 (N_9317,N_1249,N_5636);
or U9318 (N_9318,N_3723,N_5791);
nor U9319 (N_9319,N_4045,N_1164);
nand U9320 (N_9320,N_2288,N_2230);
xor U9321 (N_9321,N_1948,N_1440);
nand U9322 (N_9322,N_3056,N_5557);
and U9323 (N_9323,N_3662,N_4942);
and U9324 (N_9324,N_207,N_5458);
and U9325 (N_9325,N_2373,N_3962);
nor U9326 (N_9326,N_1243,N_2103);
nand U9327 (N_9327,N_5327,N_1690);
nor U9328 (N_9328,N_5390,N_2626);
nor U9329 (N_9329,N_2698,N_4375);
or U9330 (N_9330,N_3593,N_30);
nor U9331 (N_9331,N_4921,N_826);
xor U9332 (N_9332,N_4058,N_5753);
and U9333 (N_9333,N_1017,N_4667);
xor U9334 (N_9334,N_68,N_667);
and U9335 (N_9335,N_4811,N_6107);
or U9336 (N_9336,N_4939,N_351);
nand U9337 (N_9337,N_458,N_2656);
or U9338 (N_9338,N_3950,N_3399);
nand U9339 (N_9339,N_2146,N_1008);
xor U9340 (N_9340,N_4641,N_598);
and U9341 (N_9341,N_562,N_3526);
and U9342 (N_9342,N_3034,N_2228);
nor U9343 (N_9343,N_5347,N_3480);
xor U9344 (N_9344,N_5293,N_255);
xor U9345 (N_9345,N_1097,N_622);
or U9346 (N_9346,N_5828,N_1917);
or U9347 (N_9347,N_1710,N_630);
and U9348 (N_9348,N_1604,N_2071);
nand U9349 (N_9349,N_1932,N_1254);
nor U9350 (N_9350,N_1386,N_2652);
and U9351 (N_9351,N_2924,N_4788);
nand U9352 (N_9352,N_3889,N_4242);
nor U9353 (N_9353,N_1082,N_1612);
or U9354 (N_9354,N_3169,N_1978);
nand U9355 (N_9355,N_2895,N_1125);
and U9356 (N_9356,N_3997,N_1031);
and U9357 (N_9357,N_1945,N_703);
nor U9358 (N_9358,N_6010,N_158);
xnor U9359 (N_9359,N_1087,N_3130);
xnor U9360 (N_9360,N_3022,N_1881);
xnor U9361 (N_9361,N_1255,N_4933);
nand U9362 (N_9362,N_934,N_5769);
xor U9363 (N_9363,N_5044,N_992);
nor U9364 (N_9364,N_2306,N_749);
xor U9365 (N_9365,N_4516,N_4990);
or U9366 (N_9366,N_3361,N_5976);
nor U9367 (N_9367,N_3699,N_2885);
or U9368 (N_9368,N_851,N_5235);
nor U9369 (N_9369,N_2240,N_3586);
nand U9370 (N_9370,N_1050,N_3146);
xnor U9371 (N_9371,N_5360,N_2590);
nor U9372 (N_9372,N_4699,N_2405);
nand U9373 (N_9373,N_4992,N_64);
or U9374 (N_9374,N_2633,N_3527);
nand U9375 (N_9375,N_833,N_4581);
nand U9376 (N_9376,N_5736,N_5781);
nor U9377 (N_9377,N_2467,N_1504);
and U9378 (N_9378,N_50,N_2781);
nor U9379 (N_9379,N_5933,N_2639);
nand U9380 (N_9380,N_3574,N_4112);
nand U9381 (N_9381,N_1132,N_758);
and U9382 (N_9382,N_3507,N_1949);
xor U9383 (N_9383,N_1649,N_5209);
or U9384 (N_9384,N_4117,N_4026);
nor U9385 (N_9385,N_129,N_2562);
xor U9386 (N_9386,N_5606,N_1386);
xor U9387 (N_9387,N_2751,N_6154);
or U9388 (N_9388,N_1936,N_1976);
or U9389 (N_9389,N_2424,N_5601);
nor U9390 (N_9390,N_5512,N_3258);
nand U9391 (N_9391,N_3465,N_1192);
and U9392 (N_9392,N_1838,N_2531);
nor U9393 (N_9393,N_4223,N_622);
nor U9394 (N_9394,N_2289,N_3596);
nand U9395 (N_9395,N_5276,N_642);
or U9396 (N_9396,N_2304,N_3820);
xor U9397 (N_9397,N_796,N_3135);
xnor U9398 (N_9398,N_1427,N_968);
and U9399 (N_9399,N_1987,N_3679);
xnor U9400 (N_9400,N_5942,N_6227);
nand U9401 (N_9401,N_2524,N_5984);
nand U9402 (N_9402,N_5770,N_2526);
xnor U9403 (N_9403,N_4834,N_3496);
nor U9404 (N_9404,N_5765,N_4591);
nor U9405 (N_9405,N_1777,N_3720);
or U9406 (N_9406,N_2958,N_1338);
nor U9407 (N_9407,N_3323,N_1362);
nand U9408 (N_9408,N_2479,N_742);
xor U9409 (N_9409,N_3384,N_1101);
nand U9410 (N_9410,N_1919,N_1495);
nor U9411 (N_9411,N_5426,N_1223);
xnor U9412 (N_9412,N_2860,N_2087);
xnor U9413 (N_9413,N_3141,N_1978);
and U9414 (N_9414,N_2287,N_2832);
nand U9415 (N_9415,N_4852,N_4275);
nor U9416 (N_9416,N_4716,N_4093);
nand U9417 (N_9417,N_4787,N_3595);
and U9418 (N_9418,N_4164,N_1147);
or U9419 (N_9419,N_4014,N_5748);
xnor U9420 (N_9420,N_4764,N_2755);
nor U9421 (N_9421,N_2569,N_1598);
nor U9422 (N_9422,N_1115,N_710);
nand U9423 (N_9423,N_3961,N_1843);
and U9424 (N_9424,N_2293,N_4489);
nor U9425 (N_9425,N_4602,N_3491);
xnor U9426 (N_9426,N_3014,N_2160);
nand U9427 (N_9427,N_2397,N_4468);
or U9428 (N_9428,N_861,N_5278);
nor U9429 (N_9429,N_1291,N_727);
or U9430 (N_9430,N_1587,N_6164);
or U9431 (N_9431,N_1706,N_5211);
xor U9432 (N_9432,N_5710,N_3787);
nand U9433 (N_9433,N_2670,N_350);
or U9434 (N_9434,N_5967,N_4680);
nor U9435 (N_9435,N_593,N_5334);
and U9436 (N_9436,N_2814,N_4775);
or U9437 (N_9437,N_6168,N_3639);
or U9438 (N_9438,N_5732,N_4027);
xnor U9439 (N_9439,N_4182,N_4922);
or U9440 (N_9440,N_5253,N_1064);
nand U9441 (N_9441,N_939,N_2067);
and U9442 (N_9442,N_674,N_4132);
nand U9443 (N_9443,N_1336,N_5101);
xnor U9444 (N_9444,N_4785,N_3121);
and U9445 (N_9445,N_887,N_4673);
nor U9446 (N_9446,N_4066,N_1813);
or U9447 (N_9447,N_3307,N_5809);
and U9448 (N_9448,N_4776,N_5632);
nor U9449 (N_9449,N_3164,N_5683);
xnor U9450 (N_9450,N_203,N_1231);
nand U9451 (N_9451,N_4382,N_5601);
xor U9452 (N_9452,N_776,N_2634);
nand U9453 (N_9453,N_706,N_3865);
or U9454 (N_9454,N_2960,N_178);
and U9455 (N_9455,N_2690,N_4044);
and U9456 (N_9456,N_3291,N_6118);
nor U9457 (N_9457,N_2785,N_1472);
nand U9458 (N_9458,N_3667,N_4862);
and U9459 (N_9459,N_28,N_5267);
or U9460 (N_9460,N_2437,N_5788);
xor U9461 (N_9461,N_4748,N_1419);
xnor U9462 (N_9462,N_132,N_3135);
nor U9463 (N_9463,N_1733,N_4892);
nand U9464 (N_9464,N_3011,N_1209);
or U9465 (N_9465,N_1825,N_3059);
nor U9466 (N_9466,N_4617,N_4757);
nor U9467 (N_9467,N_2471,N_2991);
and U9468 (N_9468,N_3496,N_4538);
nand U9469 (N_9469,N_1060,N_1717);
and U9470 (N_9470,N_143,N_1605);
or U9471 (N_9471,N_1393,N_782);
nor U9472 (N_9472,N_5523,N_518);
nand U9473 (N_9473,N_5660,N_1880);
nor U9474 (N_9474,N_80,N_3731);
nor U9475 (N_9475,N_4018,N_6008);
nor U9476 (N_9476,N_4934,N_4821);
and U9477 (N_9477,N_3284,N_5623);
nand U9478 (N_9478,N_4512,N_25);
xor U9479 (N_9479,N_2274,N_1621);
or U9480 (N_9480,N_3035,N_1671);
xnor U9481 (N_9481,N_3016,N_5650);
or U9482 (N_9482,N_4191,N_3371);
nand U9483 (N_9483,N_574,N_1506);
nor U9484 (N_9484,N_475,N_1274);
or U9485 (N_9485,N_5981,N_808);
xor U9486 (N_9486,N_5524,N_573);
xnor U9487 (N_9487,N_2876,N_2197);
or U9488 (N_9488,N_165,N_4596);
nand U9489 (N_9489,N_3253,N_3872);
or U9490 (N_9490,N_2020,N_2878);
nand U9491 (N_9491,N_5731,N_4230);
and U9492 (N_9492,N_4760,N_1141);
xor U9493 (N_9493,N_1235,N_2853);
nor U9494 (N_9494,N_2753,N_6113);
xor U9495 (N_9495,N_1653,N_4400);
xnor U9496 (N_9496,N_4015,N_1662);
and U9497 (N_9497,N_5161,N_156);
nand U9498 (N_9498,N_711,N_1032);
nand U9499 (N_9499,N_5015,N_1048);
nor U9500 (N_9500,N_942,N_4411);
nand U9501 (N_9501,N_457,N_3839);
xor U9502 (N_9502,N_48,N_3097);
nor U9503 (N_9503,N_5662,N_5440);
nor U9504 (N_9504,N_2402,N_2431);
or U9505 (N_9505,N_5533,N_1421);
xor U9506 (N_9506,N_4257,N_6116);
nor U9507 (N_9507,N_1540,N_5136);
xor U9508 (N_9508,N_154,N_1584);
and U9509 (N_9509,N_1180,N_5414);
or U9510 (N_9510,N_1935,N_1767);
nand U9511 (N_9511,N_4548,N_5656);
nor U9512 (N_9512,N_1057,N_4465);
nand U9513 (N_9513,N_2395,N_5829);
or U9514 (N_9514,N_6105,N_1045);
or U9515 (N_9515,N_3433,N_3330);
xnor U9516 (N_9516,N_5076,N_115);
or U9517 (N_9517,N_5178,N_2677);
and U9518 (N_9518,N_1239,N_1132);
xnor U9519 (N_9519,N_4979,N_2789);
xnor U9520 (N_9520,N_2135,N_597);
xor U9521 (N_9521,N_5792,N_5040);
xor U9522 (N_9522,N_1697,N_1030);
xnor U9523 (N_9523,N_5333,N_4634);
nor U9524 (N_9524,N_399,N_5284);
xnor U9525 (N_9525,N_1796,N_5821);
xnor U9526 (N_9526,N_1905,N_4542);
and U9527 (N_9527,N_1956,N_958);
or U9528 (N_9528,N_5890,N_4015);
nor U9529 (N_9529,N_3881,N_3968);
xor U9530 (N_9530,N_4135,N_3872);
nor U9531 (N_9531,N_4772,N_5120);
nor U9532 (N_9532,N_6028,N_1296);
and U9533 (N_9533,N_977,N_447);
or U9534 (N_9534,N_6181,N_2878);
nand U9535 (N_9535,N_4551,N_4096);
xnor U9536 (N_9536,N_2454,N_1714);
and U9537 (N_9537,N_4411,N_771);
or U9538 (N_9538,N_1339,N_5034);
xor U9539 (N_9539,N_3384,N_5607);
or U9540 (N_9540,N_1690,N_2992);
or U9541 (N_9541,N_2864,N_5005);
and U9542 (N_9542,N_3532,N_4576);
xnor U9543 (N_9543,N_4048,N_2911);
xor U9544 (N_9544,N_5466,N_115);
or U9545 (N_9545,N_3457,N_2246);
and U9546 (N_9546,N_1230,N_4345);
or U9547 (N_9547,N_3753,N_1651);
nor U9548 (N_9548,N_772,N_2226);
or U9549 (N_9549,N_4103,N_442);
nand U9550 (N_9550,N_6165,N_4583);
nand U9551 (N_9551,N_5534,N_3552);
xor U9552 (N_9552,N_2897,N_328);
nand U9553 (N_9553,N_4105,N_2792);
nand U9554 (N_9554,N_2196,N_2327);
nor U9555 (N_9555,N_4409,N_5481);
nand U9556 (N_9556,N_4305,N_4347);
nand U9557 (N_9557,N_955,N_819);
xnor U9558 (N_9558,N_843,N_3741);
nand U9559 (N_9559,N_3205,N_3432);
or U9560 (N_9560,N_731,N_1680);
nor U9561 (N_9561,N_1181,N_2560);
xor U9562 (N_9562,N_5069,N_2229);
or U9563 (N_9563,N_6148,N_284);
nand U9564 (N_9564,N_2569,N_5026);
xnor U9565 (N_9565,N_4756,N_1726);
xor U9566 (N_9566,N_503,N_105);
xor U9567 (N_9567,N_4342,N_2619);
nor U9568 (N_9568,N_2272,N_4868);
xor U9569 (N_9569,N_580,N_4234);
or U9570 (N_9570,N_2181,N_2476);
nor U9571 (N_9571,N_4693,N_4953);
or U9572 (N_9572,N_2527,N_4575);
or U9573 (N_9573,N_1236,N_777);
and U9574 (N_9574,N_5351,N_291);
nand U9575 (N_9575,N_3350,N_1982);
xor U9576 (N_9576,N_1065,N_3869);
nor U9577 (N_9577,N_3142,N_3602);
nand U9578 (N_9578,N_760,N_4333);
or U9579 (N_9579,N_5692,N_1181);
nor U9580 (N_9580,N_5402,N_1157);
nand U9581 (N_9581,N_3705,N_1867);
xor U9582 (N_9582,N_2662,N_3704);
and U9583 (N_9583,N_4286,N_3497);
nor U9584 (N_9584,N_3473,N_2098);
nand U9585 (N_9585,N_5150,N_15);
xnor U9586 (N_9586,N_4149,N_5351);
nand U9587 (N_9587,N_3004,N_699);
nand U9588 (N_9588,N_2398,N_692);
nand U9589 (N_9589,N_6175,N_1844);
and U9590 (N_9590,N_1980,N_1687);
nor U9591 (N_9591,N_1021,N_2706);
xor U9592 (N_9592,N_3067,N_4508);
xor U9593 (N_9593,N_5970,N_2561);
or U9594 (N_9594,N_3618,N_3422);
and U9595 (N_9595,N_4776,N_3361);
and U9596 (N_9596,N_6174,N_5029);
or U9597 (N_9597,N_180,N_453);
and U9598 (N_9598,N_1655,N_3861);
xnor U9599 (N_9599,N_1351,N_5526);
and U9600 (N_9600,N_2531,N_3769);
nand U9601 (N_9601,N_3883,N_2984);
nand U9602 (N_9602,N_445,N_5459);
nor U9603 (N_9603,N_1325,N_692);
nand U9604 (N_9604,N_1541,N_6232);
xor U9605 (N_9605,N_4479,N_103);
or U9606 (N_9606,N_2507,N_5503);
nor U9607 (N_9607,N_5511,N_524);
or U9608 (N_9608,N_2869,N_2964);
nor U9609 (N_9609,N_5599,N_5371);
xnor U9610 (N_9610,N_5645,N_2120);
or U9611 (N_9611,N_6031,N_1532);
nor U9612 (N_9612,N_3825,N_5732);
nor U9613 (N_9613,N_5488,N_3069);
and U9614 (N_9614,N_4445,N_3346);
xor U9615 (N_9615,N_684,N_1775);
or U9616 (N_9616,N_3625,N_3029);
nor U9617 (N_9617,N_4409,N_2807);
or U9618 (N_9618,N_5098,N_3551);
or U9619 (N_9619,N_3660,N_2382);
nand U9620 (N_9620,N_5704,N_1023);
xor U9621 (N_9621,N_2031,N_2764);
nor U9622 (N_9622,N_2470,N_2697);
and U9623 (N_9623,N_5282,N_2608);
nand U9624 (N_9624,N_866,N_5979);
nand U9625 (N_9625,N_4677,N_1354);
and U9626 (N_9626,N_1478,N_257);
nand U9627 (N_9627,N_2990,N_4435);
nor U9628 (N_9628,N_1063,N_5116);
nand U9629 (N_9629,N_884,N_1425);
nor U9630 (N_9630,N_5439,N_3714);
or U9631 (N_9631,N_4810,N_1033);
or U9632 (N_9632,N_1935,N_3617);
xor U9633 (N_9633,N_2428,N_4012);
and U9634 (N_9634,N_61,N_1489);
and U9635 (N_9635,N_5975,N_5340);
or U9636 (N_9636,N_1501,N_2496);
and U9637 (N_9637,N_4684,N_5817);
or U9638 (N_9638,N_1306,N_1458);
nor U9639 (N_9639,N_5222,N_1883);
xnor U9640 (N_9640,N_2958,N_5923);
xnor U9641 (N_9641,N_944,N_5232);
or U9642 (N_9642,N_5367,N_4880);
nand U9643 (N_9643,N_636,N_973);
nand U9644 (N_9644,N_4519,N_1809);
xnor U9645 (N_9645,N_2246,N_4450);
nor U9646 (N_9646,N_6030,N_3563);
nor U9647 (N_9647,N_6053,N_3783);
and U9648 (N_9648,N_5075,N_1035);
or U9649 (N_9649,N_6208,N_5033);
nand U9650 (N_9650,N_181,N_4182);
xnor U9651 (N_9651,N_5205,N_2018);
xor U9652 (N_9652,N_226,N_5936);
nand U9653 (N_9653,N_6176,N_6091);
and U9654 (N_9654,N_3863,N_5256);
or U9655 (N_9655,N_4774,N_4539);
xnor U9656 (N_9656,N_1976,N_2908);
nor U9657 (N_9657,N_5738,N_5399);
nor U9658 (N_9658,N_5788,N_5749);
nor U9659 (N_9659,N_3240,N_5373);
and U9660 (N_9660,N_4686,N_3128);
and U9661 (N_9661,N_939,N_3437);
nand U9662 (N_9662,N_4902,N_3952);
and U9663 (N_9663,N_5337,N_4228);
nand U9664 (N_9664,N_410,N_6243);
nand U9665 (N_9665,N_5006,N_6076);
xor U9666 (N_9666,N_5796,N_1081);
xnor U9667 (N_9667,N_972,N_254);
nand U9668 (N_9668,N_2702,N_4388);
nand U9669 (N_9669,N_1975,N_4677);
xnor U9670 (N_9670,N_1077,N_4677);
nor U9671 (N_9671,N_4579,N_1455);
xnor U9672 (N_9672,N_5790,N_1145);
and U9673 (N_9673,N_1608,N_116);
xor U9674 (N_9674,N_1394,N_2403);
or U9675 (N_9675,N_4752,N_5414);
xnor U9676 (N_9676,N_5805,N_3111);
or U9677 (N_9677,N_4655,N_646);
xor U9678 (N_9678,N_2674,N_105);
and U9679 (N_9679,N_4215,N_1959);
xnor U9680 (N_9680,N_5886,N_2346);
nor U9681 (N_9681,N_2372,N_1577);
nand U9682 (N_9682,N_1190,N_2471);
nor U9683 (N_9683,N_1803,N_581);
or U9684 (N_9684,N_1042,N_5088);
and U9685 (N_9685,N_5302,N_3553);
or U9686 (N_9686,N_387,N_3418);
and U9687 (N_9687,N_2701,N_3046);
nor U9688 (N_9688,N_1989,N_363);
and U9689 (N_9689,N_1227,N_4803);
and U9690 (N_9690,N_3294,N_4522);
or U9691 (N_9691,N_2038,N_2913);
nand U9692 (N_9692,N_5109,N_5587);
or U9693 (N_9693,N_1403,N_989);
nor U9694 (N_9694,N_5226,N_4728);
and U9695 (N_9695,N_5503,N_3187);
or U9696 (N_9696,N_1334,N_1685);
xor U9697 (N_9697,N_6201,N_1731);
or U9698 (N_9698,N_2067,N_1245);
nand U9699 (N_9699,N_4901,N_3393);
xnor U9700 (N_9700,N_890,N_2077);
nand U9701 (N_9701,N_2408,N_1820);
xnor U9702 (N_9702,N_3995,N_5139);
nor U9703 (N_9703,N_3050,N_758);
nand U9704 (N_9704,N_4508,N_76);
nor U9705 (N_9705,N_341,N_3518);
nand U9706 (N_9706,N_3983,N_3156);
nor U9707 (N_9707,N_5383,N_977);
xnor U9708 (N_9708,N_1527,N_4972);
or U9709 (N_9709,N_3398,N_5223);
or U9710 (N_9710,N_1519,N_1288);
or U9711 (N_9711,N_5585,N_3942);
and U9712 (N_9712,N_2033,N_1566);
or U9713 (N_9713,N_2225,N_4211);
nand U9714 (N_9714,N_5897,N_414);
and U9715 (N_9715,N_4500,N_1816);
xnor U9716 (N_9716,N_107,N_5791);
nor U9717 (N_9717,N_4825,N_4309);
nor U9718 (N_9718,N_406,N_4107);
nor U9719 (N_9719,N_4557,N_5909);
or U9720 (N_9720,N_1806,N_2751);
nand U9721 (N_9721,N_2947,N_1558);
or U9722 (N_9722,N_4815,N_3625);
nand U9723 (N_9723,N_3497,N_2685);
or U9724 (N_9724,N_5864,N_5754);
xor U9725 (N_9725,N_5663,N_3519);
or U9726 (N_9726,N_4032,N_1487);
nor U9727 (N_9727,N_3799,N_3597);
nand U9728 (N_9728,N_4243,N_3960);
nor U9729 (N_9729,N_353,N_511);
nor U9730 (N_9730,N_6055,N_4099);
or U9731 (N_9731,N_2533,N_3612);
nor U9732 (N_9732,N_2414,N_2485);
and U9733 (N_9733,N_2123,N_3792);
xor U9734 (N_9734,N_4756,N_3239);
nand U9735 (N_9735,N_3503,N_4323);
xnor U9736 (N_9736,N_3346,N_4651);
or U9737 (N_9737,N_174,N_1368);
and U9738 (N_9738,N_570,N_4975);
nor U9739 (N_9739,N_5625,N_3817);
or U9740 (N_9740,N_1714,N_1737);
and U9741 (N_9741,N_4191,N_3775);
nor U9742 (N_9742,N_3041,N_1296);
or U9743 (N_9743,N_2807,N_3651);
and U9744 (N_9744,N_1198,N_1629);
nand U9745 (N_9745,N_2191,N_2639);
nor U9746 (N_9746,N_3046,N_4063);
nand U9747 (N_9747,N_3201,N_5229);
or U9748 (N_9748,N_2191,N_122);
nand U9749 (N_9749,N_1085,N_3112);
nand U9750 (N_9750,N_2164,N_4118);
nand U9751 (N_9751,N_5454,N_1712);
or U9752 (N_9752,N_654,N_57);
nand U9753 (N_9753,N_6238,N_2810);
nor U9754 (N_9754,N_1484,N_2128);
nand U9755 (N_9755,N_398,N_2417);
xnor U9756 (N_9756,N_5956,N_3532);
nand U9757 (N_9757,N_5618,N_259);
xor U9758 (N_9758,N_2380,N_3682);
and U9759 (N_9759,N_2514,N_1543);
and U9760 (N_9760,N_1779,N_2695);
or U9761 (N_9761,N_2001,N_1732);
and U9762 (N_9762,N_5472,N_509);
xnor U9763 (N_9763,N_1149,N_3478);
or U9764 (N_9764,N_246,N_2726);
and U9765 (N_9765,N_4034,N_4604);
nand U9766 (N_9766,N_1509,N_5211);
and U9767 (N_9767,N_5464,N_2162);
and U9768 (N_9768,N_643,N_4050);
nand U9769 (N_9769,N_5405,N_3677);
and U9770 (N_9770,N_3363,N_5268);
nand U9771 (N_9771,N_5352,N_6147);
and U9772 (N_9772,N_5923,N_3106);
nor U9773 (N_9773,N_3378,N_4137);
or U9774 (N_9774,N_5573,N_5101);
nor U9775 (N_9775,N_577,N_3650);
and U9776 (N_9776,N_2428,N_863);
or U9777 (N_9777,N_1270,N_5502);
and U9778 (N_9778,N_2738,N_153);
or U9779 (N_9779,N_2540,N_3237);
or U9780 (N_9780,N_1791,N_3872);
xor U9781 (N_9781,N_1859,N_4728);
nand U9782 (N_9782,N_2847,N_5638);
nor U9783 (N_9783,N_4087,N_4103);
nand U9784 (N_9784,N_3398,N_2794);
and U9785 (N_9785,N_882,N_4926);
or U9786 (N_9786,N_1792,N_5174);
and U9787 (N_9787,N_5175,N_178);
and U9788 (N_9788,N_4824,N_5271);
and U9789 (N_9789,N_319,N_4494);
nand U9790 (N_9790,N_2233,N_4006);
nand U9791 (N_9791,N_3047,N_6152);
xnor U9792 (N_9792,N_2235,N_2787);
nand U9793 (N_9793,N_5759,N_5031);
xor U9794 (N_9794,N_404,N_1817);
and U9795 (N_9795,N_3913,N_2253);
xor U9796 (N_9796,N_2420,N_1056);
nor U9797 (N_9797,N_5324,N_336);
xnor U9798 (N_9798,N_2415,N_5580);
nand U9799 (N_9799,N_86,N_5160);
nor U9800 (N_9800,N_3689,N_4455);
nand U9801 (N_9801,N_5273,N_721);
nand U9802 (N_9802,N_1661,N_2682);
or U9803 (N_9803,N_171,N_1769);
nand U9804 (N_9804,N_586,N_6111);
and U9805 (N_9805,N_3765,N_5885);
nand U9806 (N_9806,N_3028,N_4694);
nor U9807 (N_9807,N_5161,N_3147);
and U9808 (N_9808,N_1495,N_387);
and U9809 (N_9809,N_4687,N_3086);
or U9810 (N_9810,N_688,N_2287);
and U9811 (N_9811,N_3470,N_63);
nand U9812 (N_9812,N_1041,N_3726);
xor U9813 (N_9813,N_2577,N_1635);
xnor U9814 (N_9814,N_2226,N_4850);
xnor U9815 (N_9815,N_752,N_1180);
or U9816 (N_9816,N_3704,N_3345);
nor U9817 (N_9817,N_6190,N_3916);
nor U9818 (N_9818,N_5309,N_5042);
nand U9819 (N_9819,N_275,N_5194);
nor U9820 (N_9820,N_6157,N_1830);
nor U9821 (N_9821,N_6137,N_1751);
or U9822 (N_9822,N_6008,N_4643);
nor U9823 (N_9823,N_1831,N_3637);
xor U9824 (N_9824,N_2804,N_3130);
xor U9825 (N_9825,N_4752,N_5042);
or U9826 (N_9826,N_3864,N_5157);
or U9827 (N_9827,N_3540,N_2662);
or U9828 (N_9828,N_4642,N_5769);
xnor U9829 (N_9829,N_2654,N_1661);
xnor U9830 (N_9830,N_1489,N_3024);
nor U9831 (N_9831,N_4049,N_4177);
nand U9832 (N_9832,N_4067,N_2951);
or U9833 (N_9833,N_5815,N_1211);
or U9834 (N_9834,N_3682,N_5482);
or U9835 (N_9835,N_3024,N_1798);
xnor U9836 (N_9836,N_2311,N_5530);
or U9837 (N_9837,N_3373,N_2334);
xor U9838 (N_9838,N_3630,N_4944);
or U9839 (N_9839,N_5856,N_1289);
nand U9840 (N_9840,N_5453,N_293);
and U9841 (N_9841,N_2435,N_5388);
or U9842 (N_9842,N_3442,N_5352);
and U9843 (N_9843,N_5373,N_4397);
xor U9844 (N_9844,N_3736,N_2810);
nand U9845 (N_9845,N_5971,N_6180);
or U9846 (N_9846,N_2601,N_2559);
and U9847 (N_9847,N_4123,N_4961);
and U9848 (N_9848,N_3368,N_4976);
nor U9849 (N_9849,N_2188,N_5786);
nand U9850 (N_9850,N_1502,N_5065);
and U9851 (N_9851,N_2078,N_6003);
or U9852 (N_9852,N_2614,N_4730);
nand U9853 (N_9853,N_1130,N_1145);
or U9854 (N_9854,N_5045,N_4498);
or U9855 (N_9855,N_67,N_2085);
and U9856 (N_9856,N_5768,N_3771);
xnor U9857 (N_9857,N_5843,N_4925);
or U9858 (N_9858,N_107,N_6133);
xor U9859 (N_9859,N_2353,N_5245);
or U9860 (N_9860,N_5583,N_5637);
nor U9861 (N_9861,N_3563,N_5085);
and U9862 (N_9862,N_5770,N_281);
or U9863 (N_9863,N_1159,N_4497);
or U9864 (N_9864,N_6101,N_1681);
or U9865 (N_9865,N_3976,N_3024);
or U9866 (N_9866,N_296,N_4634);
xnor U9867 (N_9867,N_6056,N_92);
nor U9868 (N_9868,N_2284,N_3669);
and U9869 (N_9869,N_1272,N_1003);
nor U9870 (N_9870,N_5251,N_127);
or U9871 (N_9871,N_5974,N_5571);
xnor U9872 (N_9872,N_1647,N_1515);
nor U9873 (N_9873,N_3954,N_4588);
nor U9874 (N_9874,N_3897,N_3375);
xor U9875 (N_9875,N_4166,N_983);
nor U9876 (N_9876,N_124,N_1984);
and U9877 (N_9877,N_2346,N_2605);
and U9878 (N_9878,N_6056,N_5839);
nand U9879 (N_9879,N_1616,N_147);
and U9880 (N_9880,N_844,N_1866);
or U9881 (N_9881,N_3643,N_774);
nor U9882 (N_9882,N_4448,N_2286);
and U9883 (N_9883,N_6153,N_141);
and U9884 (N_9884,N_1832,N_3610);
nand U9885 (N_9885,N_3518,N_5710);
and U9886 (N_9886,N_3304,N_4637);
nand U9887 (N_9887,N_4519,N_2358);
or U9888 (N_9888,N_5235,N_6136);
nand U9889 (N_9889,N_979,N_6067);
and U9890 (N_9890,N_3229,N_2982);
and U9891 (N_9891,N_1195,N_5618);
nand U9892 (N_9892,N_6195,N_5791);
or U9893 (N_9893,N_1635,N_1751);
and U9894 (N_9894,N_4887,N_2215);
nand U9895 (N_9895,N_5185,N_3080);
and U9896 (N_9896,N_5701,N_3763);
and U9897 (N_9897,N_3664,N_6152);
nand U9898 (N_9898,N_2425,N_1486);
or U9899 (N_9899,N_4666,N_1946);
nor U9900 (N_9900,N_739,N_3611);
xnor U9901 (N_9901,N_4788,N_4133);
and U9902 (N_9902,N_3801,N_4786);
nor U9903 (N_9903,N_1292,N_1716);
nor U9904 (N_9904,N_4604,N_3101);
xnor U9905 (N_9905,N_5732,N_5084);
nor U9906 (N_9906,N_4155,N_4593);
xnor U9907 (N_9907,N_1301,N_5425);
xnor U9908 (N_9908,N_425,N_470);
nand U9909 (N_9909,N_3174,N_1737);
and U9910 (N_9910,N_5097,N_2595);
and U9911 (N_9911,N_1100,N_6167);
or U9912 (N_9912,N_5395,N_1436);
and U9913 (N_9913,N_2030,N_2638);
nor U9914 (N_9914,N_3073,N_1006);
nand U9915 (N_9915,N_4372,N_5786);
xor U9916 (N_9916,N_3389,N_5552);
xnor U9917 (N_9917,N_3294,N_5137);
nor U9918 (N_9918,N_2539,N_4799);
and U9919 (N_9919,N_3542,N_3468);
xnor U9920 (N_9920,N_2616,N_284);
xnor U9921 (N_9921,N_606,N_5135);
nor U9922 (N_9922,N_864,N_3473);
nor U9923 (N_9923,N_4914,N_902);
xnor U9924 (N_9924,N_2843,N_3463);
nor U9925 (N_9925,N_996,N_5963);
nand U9926 (N_9926,N_3062,N_3070);
xor U9927 (N_9927,N_1729,N_4614);
or U9928 (N_9928,N_1463,N_1392);
or U9929 (N_9929,N_1100,N_4889);
xor U9930 (N_9930,N_3025,N_1006);
and U9931 (N_9931,N_5390,N_3527);
nor U9932 (N_9932,N_3435,N_3904);
or U9933 (N_9933,N_5221,N_227);
or U9934 (N_9934,N_2099,N_2704);
or U9935 (N_9935,N_5457,N_2115);
nand U9936 (N_9936,N_4629,N_5265);
nor U9937 (N_9937,N_5186,N_1791);
and U9938 (N_9938,N_6047,N_5653);
nand U9939 (N_9939,N_1092,N_353);
and U9940 (N_9940,N_1964,N_3340);
nor U9941 (N_9941,N_2979,N_1428);
xor U9942 (N_9942,N_3311,N_2768);
and U9943 (N_9943,N_6231,N_2764);
and U9944 (N_9944,N_3659,N_3887);
xor U9945 (N_9945,N_5045,N_3677);
nand U9946 (N_9946,N_2051,N_2488);
nor U9947 (N_9947,N_1214,N_797);
or U9948 (N_9948,N_1773,N_427);
xnor U9949 (N_9949,N_1313,N_3182);
or U9950 (N_9950,N_4541,N_1382);
or U9951 (N_9951,N_921,N_221);
or U9952 (N_9952,N_2667,N_4352);
nand U9953 (N_9953,N_617,N_1106);
or U9954 (N_9954,N_814,N_3044);
nand U9955 (N_9955,N_5033,N_4140);
nor U9956 (N_9956,N_837,N_5855);
xnor U9957 (N_9957,N_2406,N_1621);
nor U9958 (N_9958,N_902,N_4098);
xor U9959 (N_9959,N_1782,N_5369);
xor U9960 (N_9960,N_2625,N_3010);
nand U9961 (N_9961,N_2978,N_892);
or U9962 (N_9962,N_327,N_2585);
and U9963 (N_9963,N_2286,N_1794);
and U9964 (N_9964,N_3364,N_4648);
nand U9965 (N_9965,N_3619,N_5303);
and U9966 (N_9966,N_3367,N_406);
xnor U9967 (N_9967,N_982,N_3864);
and U9968 (N_9968,N_3859,N_5326);
nand U9969 (N_9969,N_523,N_1279);
nor U9970 (N_9970,N_4344,N_412);
and U9971 (N_9971,N_3353,N_1107);
or U9972 (N_9972,N_658,N_4318);
nor U9973 (N_9973,N_312,N_4809);
nor U9974 (N_9974,N_4393,N_629);
nor U9975 (N_9975,N_6092,N_616);
and U9976 (N_9976,N_4164,N_2695);
nand U9977 (N_9977,N_6166,N_3877);
nor U9978 (N_9978,N_4657,N_895);
or U9979 (N_9979,N_709,N_2506);
or U9980 (N_9980,N_4458,N_6247);
or U9981 (N_9981,N_4968,N_3246);
and U9982 (N_9982,N_1567,N_2171);
or U9983 (N_9983,N_4148,N_5118);
and U9984 (N_9984,N_4773,N_763);
and U9985 (N_9985,N_3849,N_867);
nor U9986 (N_9986,N_2337,N_8);
xnor U9987 (N_9987,N_5367,N_6191);
and U9988 (N_9988,N_5263,N_5625);
nand U9989 (N_9989,N_4747,N_3036);
nand U9990 (N_9990,N_774,N_1342);
nand U9991 (N_9991,N_1482,N_1796);
xor U9992 (N_9992,N_3514,N_3583);
nor U9993 (N_9993,N_3519,N_1827);
nand U9994 (N_9994,N_1327,N_1511);
and U9995 (N_9995,N_251,N_3663);
xnor U9996 (N_9996,N_5892,N_1738);
xnor U9997 (N_9997,N_2918,N_3006);
and U9998 (N_9998,N_3266,N_5875);
nor U9999 (N_9999,N_5431,N_3665);
and U10000 (N_10000,N_6138,N_3633);
xor U10001 (N_10001,N_6232,N_1998);
nand U10002 (N_10002,N_4088,N_5106);
nor U10003 (N_10003,N_277,N_1042);
nor U10004 (N_10004,N_4462,N_1569);
nand U10005 (N_10005,N_3381,N_3396);
nand U10006 (N_10006,N_4358,N_4837);
or U10007 (N_10007,N_2517,N_623);
nand U10008 (N_10008,N_1064,N_2852);
and U10009 (N_10009,N_4992,N_3894);
and U10010 (N_10010,N_5843,N_3391);
and U10011 (N_10011,N_4360,N_1916);
nor U10012 (N_10012,N_5189,N_6016);
nand U10013 (N_10013,N_2421,N_3564);
and U10014 (N_10014,N_52,N_4317);
and U10015 (N_10015,N_5005,N_3304);
xnor U10016 (N_10016,N_2068,N_754);
or U10017 (N_10017,N_1776,N_4824);
xor U10018 (N_10018,N_506,N_2122);
nor U10019 (N_10019,N_1287,N_1895);
nand U10020 (N_10020,N_5021,N_4537);
and U10021 (N_10021,N_1458,N_2815);
and U10022 (N_10022,N_5353,N_1605);
xor U10023 (N_10023,N_2843,N_1493);
or U10024 (N_10024,N_6073,N_1912);
and U10025 (N_10025,N_155,N_3767);
xor U10026 (N_10026,N_4358,N_4228);
and U10027 (N_10027,N_5533,N_2352);
xnor U10028 (N_10028,N_140,N_32);
and U10029 (N_10029,N_1987,N_3859);
or U10030 (N_10030,N_4807,N_3539);
or U10031 (N_10031,N_887,N_3959);
nand U10032 (N_10032,N_5908,N_3522);
and U10033 (N_10033,N_4482,N_4045);
and U10034 (N_10034,N_4348,N_3266);
or U10035 (N_10035,N_1949,N_2610);
xor U10036 (N_10036,N_2702,N_193);
nor U10037 (N_10037,N_256,N_4336);
nand U10038 (N_10038,N_5648,N_1959);
nand U10039 (N_10039,N_1052,N_2869);
or U10040 (N_10040,N_4411,N_4529);
and U10041 (N_10041,N_3057,N_2222);
or U10042 (N_10042,N_6138,N_1126);
nand U10043 (N_10043,N_4723,N_5640);
xnor U10044 (N_10044,N_5676,N_1961);
nor U10045 (N_10045,N_2320,N_2438);
nand U10046 (N_10046,N_1980,N_3742);
xnor U10047 (N_10047,N_1566,N_4372);
nor U10048 (N_10048,N_1439,N_4756);
and U10049 (N_10049,N_5227,N_849);
nand U10050 (N_10050,N_5237,N_4511);
nor U10051 (N_10051,N_4296,N_5148);
xor U10052 (N_10052,N_5460,N_351);
nand U10053 (N_10053,N_237,N_246);
and U10054 (N_10054,N_4069,N_5055);
and U10055 (N_10055,N_4475,N_4519);
or U10056 (N_10056,N_6246,N_2981);
nand U10057 (N_10057,N_3899,N_5220);
and U10058 (N_10058,N_2055,N_1065);
or U10059 (N_10059,N_1023,N_4527);
xnor U10060 (N_10060,N_2719,N_2228);
nand U10061 (N_10061,N_2728,N_4824);
nand U10062 (N_10062,N_3500,N_4462);
and U10063 (N_10063,N_3708,N_4179);
nor U10064 (N_10064,N_5323,N_5052);
nand U10065 (N_10065,N_5442,N_4935);
nand U10066 (N_10066,N_4437,N_2455);
xnor U10067 (N_10067,N_653,N_2863);
and U10068 (N_10068,N_6075,N_2780);
and U10069 (N_10069,N_1235,N_3122);
and U10070 (N_10070,N_4284,N_4625);
nand U10071 (N_10071,N_4911,N_1988);
xnor U10072 (N_10072,N_1997,N_4916);
or U10073 (N_10073,N_3696,N_2450);
and U10074 (N_10074,N_655,N_5716);
and U10075 (N_10075,N_2815,N_1495);
nor U10076 (N_10076,N_4640,N_2044);
xor U10077 (N_10077,N_2291,N_4475);
nand U10078 (N_10078,N_2465,N_1995);
nand U10079 (N_10079,N_3478,N_127);
nand U10080 (N_10080,N_512,N_2502);
or U10081 (N_10081,N_4777,N_4327);
xor U10082 (N_10082,N_6098,N_747);
nand U10083 (N_10083,N_880,N_2727);
or U10084 (N_10084,N_2752,N_6191);
nand U10085 (N_10085,N_1615,N_376);
or U10086 (N_10086,N_5442,N_447);
nand U10087 (N_10087,N_3123,N_3756);
nand U10088 (N_10088,N_2272,N_162);
nand U10089 (N_10089,N_270,N_754);
nor U10090 (N_10090,N_1481,N_2457);
nor U10091 (N_10091,N_4515,N_998);
or U10092 (N_10092,N_5380,N_3846);
nand U10093 (N_10093,N_6219,N_3488);
xnor U10094 (N_10094,N_806,N_1654);
nand U10095 (N_10095,N_3015,N_2430);
or U10096 (N_10096,N_3694,N_2130);
or U10097 (N_10097,N_4908,N_1461);
and U10098 (N_10098,N_4805,N_5971);
or U10099 (N_10099,N_119,N_2976);
xor U10100 (N_10100,N_1511,N_3108);
or U10101 (N_10101,N_417,N_5682);
xor U10102 (N_10102,N_2340,N_2670);
or U10103 (N_10103,N_2114,N_618);
or U10104 (N_10104,N_2937,N_3048);
xor U10105 (N_10105,N_2999,N_5690);
nor U10106 (N_10106,N_3577,N_5965);
xnor U10107 (N_10107,N_565,N_5855);
xor U10108 (N_10108,N_5027,N_1596);
or U10109 (N_10109,N_3703,N_609);
nor U10110 (N_10110,N_3722,N_712);
or U10111 (N_10111,N_4722,N_1546);
nor U10112 (N_10112,N_2265,N_113);
or U10113 (N_10113,N_4432,N_379);
or U10114 (N_10114,N_3568,N_2283);
and U10115 (N_10115,N_6058,N_3282);
or U10116 (N_10116,N_4495,N_1600);
or U10117 (N_10117,N_3501,N_929);
nand U10118 (N_10118,N_4008,N_6226);
nand U10119 (N_10119,N_145,N_3654);
nand U10120 (N_10120,N_4159,N_6121);
xnor U10121 (N_10121,N_3697,N_163);
and U10122 (N_10122,N_1,N_6173);
and U10123 (N_10123,N_250,N_3573);
or U10124 (N_10124,N_3710,N_5585);
xnor U10125 (N_10125,N_4844,N_6168);
nand U10126 (N_10126,N_2927,N_591);
or U10127 (N_10127,N_1585,N_2921);
and U10128 (N_10128,N_1649,N_2911);
nor U10129 (N_10129,N_3387,N_5611);
nand U10130 (N_10130,N_5802,N_4935);
xor U10131 (N_10131,N_5877,N_4933);
and U10132 (N_10132,N_3769,N_2559);
nand U10133 (N_10133,N_4962,N_2741);
xor U10134 (N_10134,N_6232,N_2795);
nor U10135 (N_10135,N_5482,N_3287);
nor U10136 (N_10136,N_4772,N_1571);
nor U10137 (N_10137,N_2824,N_4642);
xor U10138 (N_10138,N_1768,N_1656);
and U10139 (N_10139,N_1524,N_5636);
and U10140 (N_10140,N_4887,N_149);
nor U10141 (N_10141,N_1487,N_694);
and U10142 (N_10142,N_5607,N_5995);
nor U10143 (N_10143,N_1896,N_5012);
and U10144 (N_10144,N_855,N_5105);
or U10145 (N_10145,N_3253,N_6178);
nand U10146 (N_10146,N_185,N_237);
and U10147 (N_10147,N_4031,N_2440);
nand U10148 (N_10148,N_2292,N_3909);
and U10149 (N_10149,N_5688,N_4471);
nand U10150 (N_10150,N_3414,N_5696);
xor U10151 (N_10151,N_293,N_266);
xor U10152 (N_10152,N_3952,N_1626);
and U10153 (N_10153,N_1134,N_5117);
nor U10154 (N_10154,N_5178,N_396);
nor U10155 (N_10155,N_4192,N_2435);
nor U10156 (N_10156,N_827,N_5849);
nor U10157 (N_10157,N_2495,N_4343);
nor U10158 (N_10158,N_2924,N_2330);
and U10159 (N_10159,N_703,N_4538);
nor U10160 (N_10160,N_143,N_648);
and U10161 (N_10161,N_5769,N_3437);
xnor U10162 (N_10162,N_5801,N_3775);
xnor U10163 (N_10163,N_4977,N_3554);
and U10164 (N_10164,N_1761,N_2446);
nor U10165 (N_10165,N_5177,N_3891);
xnor U10166 (N_10166,N_764,N_5246);
nand U10167 (N_10167,N_2909,N_6198);
and U10168 (N_10168,N_1375,N_2460);
xnor U10169 (N_10169,N_5156,N_3091);
nand U10170 (N_10170,N_314,N_1732);
or U10171 (N_10171,N_3009,N_4764);
and U10172 (N_10172,N_152,N_2246);
and U10173 (N_10173,N_519,N_3414);
and U10174 (N_10174,N_2854,N_2866);
and U10175 (N_10175,N_5412,N_6233);
nand U10176 (N_10176,N_4977,N_3954);
nor U10177 (N_10177,N_1749,N_4544);
or U10178 (N_10178,N_4478,N_3253);
xnor U10179 (N_10179,N_4928,N_3214);
nor U10180 (N_10180,N_4977,N_4222);
or U10181 (N_10181,N_3339,N_2383);
or U10182 (N_10182,N_1285,N_764);
nand U10183 (N_10183,N_717,N_4007);
and U10184 (N_10184,N_4176,N_5452);
and U10185 (N_10185,N_5261,N_208);
xor U10186 (N_10186,N_5398,N_23);
nor U10187 (N_10187,N_3744,N_4638);
and U10188 (N_10188,N_4208,N_2748);
nand U10189 (N_10189,N_729,N_5522);
nand U10190 (N_10190,N_4326,N_85);
nor U10191 (N_10191,N_2018,N_3411);
or U10192 (N_10192,N_2898,N_5684);
nand U10193 (N_10193,N_4762,N_1797);
or U10194 (N_10194,N_824,N_6146);
nor U10195 (N_10195,N_3695,N_1733);
or U10196 (N_10196,N_5618,N_1087);
nor U10197 (N_10197,N_5626,N_1505);
xor U10198 (N_10198,N_4920,N_5223);
and U10199 (N_10199,N_528,N_1286);
nor U10200 (N_10200,N_837,N_2694);
and U10201 (N_10201,N_5174,N_3838);
nor U10202 (N_10202,N_5195,N_1380);
or U10203 (N_10203,N_443,N_5330);
nand U10204 (N_10204,N_78,N_346);
nand U10205 (N_10205,N_6044,N_4410);
nor U10206 (N_10206,N_569,N_5696);
nand U10207 (N_10207,N_3858,N_2758);
and U10208 (N_10208,N_3577,N_3912);
nor U10209 (N_10209,N_6130,N_3983);
nor U10210 (N_10210,N_251,N_992);
nand U10211 (N_10211,N_4353,N_4217);
and U10212 (N_10212,N_1228,N_5091);
nand U10213 (N_10213,N_900,N_2280);
and U10214 (N_10214,N_3474,N_3964);
and U10215 (N_10215,N_2265,N_61);
xnor U10216 (N_10216,N_3009,N_5418);
or U10217 (N_10217,N_1334,N_3610);
and U10218 (N_10218,N_3506,N_4479);
and U10219 (N_10219,N_5529,N_4573);
xnor U10220 (N_10220,N_5476,N_3059);
or U10221 (N_10221,N_4625,N_4989);
nor U10222 (N_10222,N_1468,N_3324);
and U10223 (N_10223,N_5111,N_1406);
nor U10224 (N_10224,N_4436,N_3028);
nor U10225 (N_10225,N_5134,N_1847);
xnor U10226 (N_10226,N_499,N_6227);
and U10227 (N_10227,N_556,N_1150);
or U10228 (N_10228,N_3416,N_5656);
or U10229 (N_10229,N_3769,N_1633);
nand U10230 (N_10230,N_101,N_5024);
or U10231 (N_10231,N_4438,N_2545);
or U10232 (N_10232,N_4600,N_3689);
nand U10233 (N_10233,N_2628,N_5537);
or U10234 (N_10234,N_3368,N_4301);
or U10235 (N_10235,N_4944,N_2971);
and U10236 (N_10236,N_6037,N_4262);
or U10237 (N_10237,N_6164,N_4130);
and U10238 (N_10238,N_1910,N_1006);
xor U10239 (N_10239,N_5497,N_3726);
and U10240 (N_10240,N_647,N_5536);
xnor U10241 (N_10241,N_6176,N_5791);
and U10242 (N_10242,N_5962,N_4196);
xnor U10243 (N_10243,N_5347,N_5556);
nand U10244 (N_10244,N_2385,N_5732);
nand U10245 (N_10245,N_5058,N_3612);
and U10246 (N_10246,N_808,N_5251);
xnor U10247 (N_10247,N_3820,N_3823);
nand U10248 (N_10248,N_679,N_3670);
nor U10249 (N_10249,N_1272,N_131);
and U10250 (N_10250,N_2527,N_4745);
or U10251 (N_10251,N_6098,N_5527);
nand U10252 (N_10252,N_6159,N_973);
or U10253 (N_10253,N_3423,N_1131);
nand U10254 (N_10254,N_3744,N_252);
nor U10255 (N_10255,N_3560,N_1630);
xor U10256 (N_10256,N_2726,N_3530);
and U10257 (N_10257,N_2125,N_918);
and U10258 (N_10258,N_2582,N_3061);
nor U10259 (N_10259,N_6223,N_6175);
nor U10260 (N_10260,N_5587,N_5669);
xnor U10261 (N_10261,N_5947,N_4632);
xnor U10262 (N_10262,N_3553,N_3687);
nor U10263 (N_10263,N_1633,N_5889);
or U10264 (N_10264,N_2948,N_1452);
xor U10265 (N_10265,N_1387,N_1069);
xnor U10266 (N_10266,N_1905,N_2935);
and U10267 (N_10267,N_3048,N_3498);
or U10268 (N_10268,N_502,N_432);
nor U10269 (N_10269,N_915,N_4720);
or U10270 (N_10270,N_4335,N_3345);
nand U10271 (N_10271,N_2448,N_3618);
nor U10272 (N_10272,N_3730,N_570);
or U10273 (N_10273,N_5007,N_4384);
and U10274 (N_10274,N_4717,N_3944);
or U10275 (N_10275,N_3246,N_5069);
nand U10276 (N_10276,N_1291,N_2630);
nor U10277 (N_10277,N_3013,N_874);
nor U10278 (N_10278,N_5029,N_5174);
or U10279 (N_10279,N_4673,N_500);
and U10280 (N_10280,N_5349,N_3211);
xor U10281 (N_10281,N_1937,N_1565);
xor U10282 (N_10282,N_4185,N_1392);
nand U10283 (N_10283,N_3323,N_907);
nor U10284 (N_10284,N_2848,N_3764);
and U10285 (N_10285,N_4821,N_4699);
nor U10286 (N_10286,N_1211,N_6149);
nor U10287 (N_10287,N_4840,N_3921);
or U10288 (N_10288,N_5811,N_2889);
xnor U10289 (N_10289,N_2524,N_4307);
xor U10290 (N_10290,N_830,N_5176);
nand U10291 (N_10291,N_2772,N_5813);
nor U10292 (N_10292,N_5651,N_2843);
nor U10293 (N_10293,N_4716,N_2883);
or U10294 (N_10294,N_5360,N_2787);
xnor U10295 (N_10295,N_104,N_410);
nor U10296 (N_10296,N_2238,N_842);
nand U10297 (N_10297,N_1170,N_769);
nor U10298 (N_10298,N_5739,N_2565);
nor U10299 (N_10299,N_6215,N_3830);
nand U10300 (N_10300,N_2269,N_4977);
nand U10301 (N_10301,N_4276,N_1419);
or U10302 (N_10302,N_3201,N_1166);
or U10303 (N_10303,N_1207,N_3630);
xnor U10304 (N_10304,N_618,N_3959);
and U10305 (N_10305,N_2709,N_4367);
xor U10306 (N_10306,N_4270,N_3582);
and U10307 (N_10307,N_1513,N_5814);
or U10308 (N_10308,N_3358,N_3513);
or U10309 (N_10309,N_4579,N_5299);
nand U10310 (N_10310,N_4670,N_5283);
nand U10311 (N_10311,N_5868,N_1266);
nand U10312 (N_10312,N_3283,N_2459);
and U10313 (N_10313,N_5069,N_4385);
nor U10314 (N_10314,N_583,N_2149);
or U10315 (N_10315,N_23,N_2490);
or U10316 (N_10316,N_2462,N_5262);
xnor U10317 (N_10317,N_1297,N_5736);
and U10318 (N_10318,N_2005,N_1706);
or U10319 (N_10319,N_316,N_5681);
nand U10320 (N_10320,N_5796,N_1977);
xor U10321 (N_10321,N_6050,N_536);
nand U10322 (N_10322,N_1209,N_3154);
or U10323 (N_10323,N_4519,N_2514);
nand U10324 (N_10324,N_4467,N_3113);
nor U10325 (N_10325,N_259,N_94);
and U10326 (N_10326,N_456,N_4613);
and U10327 (N_10327,N_2815,N_5714);
and U10328 (N_10328,N_4340,N_3778);
xor U10329 (N_10329,N_2521,N_1266);
nor U10330 (N_10330,N_4533,N_97);
nand U10331 (N_10331,N_5747,N_3773);
nand U10332 (N_10332,N_5952,N_3939);
or U10333 (N_10333,N_917,N_2732);
or U10334 (N_10334,N_5858,N_3950);
xnor U10335 (N_10335,N_4273,N_5279);
and U10336 (N_10336,N_5592,N_4642);
nand U10337 (N_10337,N_3601,N_5671);
and U10338 (N_10338,N_5275,N_2239);
or U10339 (N_10339,N_3341,N_1317);
and U10340 (N_10340,N_4666,N_152);
xor U10341 (N_10341,N_224,N_1867);
nor U10342 (N_10342,N_2028,N_860);
nand U10343 (N_10343,N_4742,N_5196);
nor U10344 (N_10344,N_3004,N_285);
xor U10345 (N_10345,N_1424,N_4719);
or U10346 (N_10346,N_5433,N_1096);
and U10347 (N_10347,N_723,N_191);
nor U10348 (N_10348,N_3771,N_6048);
xor U10349 (N_10349,N_1816,N_4351);
or U10350 (N_10350,N_4653,N_5006);
or U10351 (N_10351,N_4648,N_1960);
or U10352 (N_10352,N_4766,N_551);
nor U10353 (N_10353,N_2782,N_4773);
and U10354 (N_10354,N_3960,N_3254);
and U10355 (N_10355,N_2837,N_5046);
nor U10356 (N_10356,N_1258,N_6129);
nand U10357 (N_10357,N_5373,N_5239);
or U10358 (N_10358,N_1136,N_4065);
and U10359 (N_10359,N_1021,N_422);
or U10360 (N_10360,N_1281,N_4104);
or U10361 (N_10361,N_3338,N_767);
xor U10362 (N_10362,N_2531,N_1544);
or U10363 (N_10363,N_2830,N_4628);
xnor U10364 (N_10364,N_6224,N_3191);
or U10365 (N_10365,N_3059,N_2611);
nand U10366 (N_10366,N_4119,N_6244);
or U10367 (N_10367,N_5996,N_3089);
nand U10368 (N_10368,N_2545,N_3579);
or U10369 (N_10369,N_2534,N_133);
nand U10370 (N_10370,N_1872,N_4401);
nand U10371 (N_10371,N_2585,N_987);
nor U10372 (N_10372,N_998,N_3762);
nor U10373 (N_10373,N_2188,N_4668);
nand U10374 (N_10374,N_757,N_2621);
nand U10375 (N_10375,N_3587,N_5159);
nor U10376 (N_10376,N_3694,N_2125);
nand U10377 (N_10377,N_1973,N_2303);
xor U10378 (N_10378,N_5424,N_3780);
nand U10379 (N_10379,N_1503,N_3058);
or U10380 (N_10380,N_3823,N_581);
or U10381 (N_10381,N_2763,N_189);
nor U10382 (N_10382,N_3974,N_2302);
and U10383 (N_10383,N_4667,N_5171);
nor U10384 (N_10384,N_2877,N_4974);
or U10385 (N_10385,N_4321,N_4159);
or U10386 (N_10386,N_2884,N_5520);
nor U10387 (N_10387,N_5509,N_978);
and U10388 (N_10388,N_2724,N_5621);
nand U10389 (N_10389,N_2482,N_3233);
xor U10390 (N_10390,N_1985,N_1060);
and U10391 (N_10391,N_5187,N_118);
or U10392 (N_10392,N_1122,N_4478);
or U10393 (N_10393,N_4510,N_4362);
or U10394 (N_10394,N_5855,N_6013);
or U10395 (N_10395,N_4449,N_109);
nand U10396 (N_10396,N_2722,N_14);
and U10397 (N_10397,N_3648,N_98);
or U10398 (N_10398,N_224,N_4676);
nand U10399 (N_10399,N_5541,N_1489);
nand U10400 (N_10400,N_5080,N_4232);
or U10401 (N_10401,N_5264,N_3783);
nor U10402 (N_10402,N_2184,N_1468);
nor U10403 (N_10403,N_5004,N_1382);
xnor U10404 (N_10404,N_4727,N_523);
nor U10405 (N_10405,N_3441,N_3210);
and U10406 (N_10406,N_3351,N_4393);
nand U10407 (N_10407,N_5791,N_4780);
nor U10408 (N_10408,N_1503,N_2112);
or U10409 (N_10409,N_6217,N_2637);
xnor U10410 (N_10410,N_2701,N_672);
nand U10411 (N_10411,N_4928,N_5418);
or U10412 (N_10412,N_551,N_929);
nor U10413 (N_10413,N_2932,N_4005);
nor U10414 (N_10414,N_3411,N_4324);
xnor U10415 (N_10415,N_199,N_3415);
nor U10416 (N_10416,N_49,N_3283);
nor U10417 (N_10417,N_2006,N_2506);
and U10418 (N_10418,N_4374,N_1942);
and U10419 (N_10419,N_6247,N_3870);
nor U10420 (N_10420,N_663,N_3214);
xor U10421 (N_10421,N_505,N_3374);
or U10422 (N_10422,N_385,N_2935);
xnor U10423 (N_10423,N_2456,N_5787);
or U10424 (N_10424,N_5402,N_5419);
nand U10425 (N_10425,N_1393,N_2264);
xnor U10426 (N_10426,N_5892,N_1234);
nand U10427 (N_10427,N_5780,N_2819);
and U10428 (N_10428,N_398,N_3152);
nand U10429 (N_10429,N_575,N_5188);
nor U10430 (N_10430,N_2625,N_2792);
nand U10431 (N_10431,N_5776,N_1163);
nor U10432 (N_10432,N_1834,N_3666);
and U10433 (N_10433,N_5627,N_2182);
or U10434 (N_10434,N_5068,N_5110);
and U10435 (N_10435,N_5119,N_5776);
nor U10436 (N_10436,N_3247,N_4613);
and U10437 (N_10437,N_679,N_5714);
nor U10438 (N_10438,N_2514,N_585);
nand U10439 (N_10439,N_727,N_1344);
nor U10440 (N_10440,N_1329,N_2667);
nand U10441 (N_10441,N_5759,N_3897);
or U10442 (N_10442,N_1988,N_3966);
xnor U10443 (N_10443,N_944,N_19);
nand U10444 (N_10444,N_2197,N_3415);
nor U10445 (N_10445,N_6013,N_995);
xnor U10446 (N_10446,N_6225,N_5216);
nand U10447 (N_10447,N_4615,N_2875);
nor U10448 (N_10448,N_2531,N_5234);
xnor U10449 (N_10449,N_3089,N_2016);
or U10450 (N_10450,N_5266,N_3633);
nor U10451 (N_10451,N_2138,N_5991);
and U10452 (N_10452,N_1387,N_4065);
nor U10453 (N_10453,N_117,N_4748);
or U10454 (N_10454,N_3914,N_1796);
nor U10455 (N_10455,N_1663,N_6003);
xor U10456 (N_10456,N_5834,N_1997);
xnor U10457 (N_10457,N_2850,N_3469);
nor U10458 (N_10458,N_3989,N_4312);
xor U10459 (N_10459,N_3863,N_1861);
xor U10460 (N_10460,N_5845,N_3901);
xnor U10461 (N_10461,N_2839,N_2415);
nor U10462 (N_10462,N_6182,N_2827);
nor U10463 (N_10463,N_3718,N_3160);
and U10464 (N_10464,N_3849,N_646);
nand U10465 (N_10465,N_2496,N_610);
nand U10466 (N_10466,N_1462,N_6202);
and U10467 (N_10467,N_4269,N_1500);
xor U10468 (N_10468,N_1693,N_5745);
and U10469 (N_10469,N_81,N_3451);
and U10470 (N_10470,N_3190,N_2605);
nor U10471 (N_10471,N_3853,N_3507);
xor U10472 (N_10472,N_5052,N_2437);
nand U10473 (N_10473,N_4625,N_5914);
nor U10474 (N_10474,N_4399,N_1449);
or U10475 (N_10475,N_5219,N_5169);
nand U10476 (N_10476,N_2961,N_3964);
and U10477 (N_10477,N_3781,N_5124);
nand U10478 (N_10478,N_6035,N_3310);
xnor U10479 (N_10479,N_2928,N_3312);
nor U10480 (N_10480,N_4512,N_1895);
and U10481 (N_10481,N_1228,N_447);
xor U10482 (N_10482,N_5389,N_1129);
nand U10483 (N_10483,N_1711,N_1984);
nand U10484 (N_10484,N_1359,N_5519);
and U10485 (N_10485,N_4128,N_4216);
or U10486 (N_10486,N_1063,N_5047);
nand U10487 (N_10487,N_623,N_1065);
and U10488 (N_10488,N_1162,N_625);
nand U10489 (N_10489,N_5798,N_2292);
or U10490 (N_10490,N_4386,N_784);
nand U10491 (N_10491,N_2993,N_1385);
xor U10492 (N_10492,N_6110,N_3456);
nand U10493 (N_10493,N_2261,N_4924);
xnor U10494 (N_10494,N_420,N_5817);
or U10495 (N_10495,N_1202,N_5947);
xor U10496 (N_10496,N_5115,N_6196);
and U10497 (N_10497,N_3170,N_2213);
or U10498 (N_10498,N_3410,N_3438);
xnor U10499 (N_10499,N_3177,N_4484);
xor U10500 (N_10500,N_4927,N_5118);
nand U10501 (N_10501,N_3935,N_4759);
and U10502 (N_10502,N_33,N_4214);
and U10503 (N_10503,N_5602,N_3102);
or U10504 (N_10504,N_4834,N_2016);
nor U10505 (N_10505,N_1844,N_1911);
nor U10506 (N_10506,N_5348,N_2400);
xor U10507 (N_10507,N_1431,N_1744);
or U10508 (N_10508,N_5600,N_3221);
or U10509 (N_10509,N_1042,N_3518);
and U10510 (N_10510,N_5123,N_3753);
xnor U10511 (N_10511,N_675,N_2975);
or U10512 (N_10512,N_5050,N_4517);
nor U10513 (N_10513,N_4335,N_1035);
nand U10514 (N_10514,N_4170,N_4112);
or U10515 (N_10515,N_4325,N_152);
xor U10516 (N_10516,N_1548,N_2256);
nor U10517 (N_10517,N_3442,N_307);
and U10518 (N_10518,N_5391,N_3427);
and U10519 (N_10519,N_2170,N_4015);
or U10520 (N_10520,N_3559,N_5765);
nor U10521 (N_10521,N_3458,N_4244);
and U10522 (N_10522,N_1177,N_4410);
xnor U10523 (N_10523,N_4774,N_4353);
or U10524 (N_10524,N_1389,N_1619);
nor U10525 (N_10525,N_1345,N_3194);
and U10526 (N_10526,N_2415,N_2350);
nand U10527 (N_10527,N_6000,N_1089);
nor U10528 (N_10528,N_6129,N_3816);
or U10529 (N_10529,N_5638,N_1319);
or U10530 (N_10530,N_80,N_2551);
or U10531 (N_10531,N_1166,N_5615);
and U10532 (N_10532,N_1423,N_6135);
nand U10533 (N_10533,N_5323,N_1415);
xor U10534 (N_10534,N_712,N_1173);
or U10535 (N_10535,N_2358,N_2534);
xor U10536 (N_10536,N_4496,N_441);
xnor U10537 (N_10537,N_950,N_4347);
or U10538 (N_10538,N_3303,N_3112);
and U10539 (N_10539,N_2968,N_4586);
nand U10540 (N_10540,N_5553,N_3206);
nand U10541 (N_10541,N_899,N_2212);
nand U10542 (N_10542,N_3228,N_3575);
nand U10543 (N_10543,N_5205,N_2097);
nor U10544 (N_10544,N_3871,N_4963);
nand U10545 (N_10545,N_3729,N_653);
xor U10546 (N_10546,N_1770,N_2771);
nor U10547 (N_10547,N_5046,N_2388);
nand U10548 (N_10548,N_104,N_2965);
nand U10549 (N_10549,N_1054,N_193);
nor U10550 (N_10550,N_3664,N_339);
xnor U10551 (N_10551,N_5095,N_2601);
nor U10552 (N_10552,N_2915,N_2440);
nand U10553 (N_10553,N_5133,N_5485);
xnor U10554 (N_10554,N_4272,N_3357);
or U10555 (N_10555,N_547,N_1824);
xnor U10556 (N_10556,N_2581,N_1847);
nor U10557 (N_10557,N_1515,N_5550);
nand U10558 (N_10558,N_198,N_893);
nand U10559 (N_10559,N_2695,N_73);
xor U10560 (N_10560,N_2935,N_206);
or U10561 (N_10561,N_3782,N_4757);
or U10562 (N_10562,N_3616,N_279);
and U10563 (N_10563,N_383,N_3174);
nor U10564 (N_10564,N_2706,N_2018);
and U10565 (N_10565,N_4993,N_4494);
nand U10566 (N_10566,N_6231,N_5667);
nand U10567 (N_10567,N_3391,N_5178);
or U10568 (N_10568,N_5622,N_2402);
nor U10569 (N_10569,N_2345,N_4923);
nand U10570 (N_10570,N_3103,N_694);
nand U10571 (N_10571,N_2227,N_672);
and U10572 (N_10572,N_3959,N_5681);
nor U10573 (N_10573,N_5201,N_3896);
xnor U10574 (N_10574,N_638,N_5497);
or U10575 (N_10575,N_2019,N_1363);
nor U10576 (N_10576,N_282,N_4429);
or U10577 (N_10577,N_3272,N_410);
nor U10578 (N_10578,N_5580,N_4332);
or U10579 (N_10579,N_2827,N_2313);
nand U10580 (N_10580,N_5093,N_1636);
nor U10581 (N_10581,N_562,N_1968);
nor U10582 (N_10582,N_5213,N_4386);
nand U10583 (N_10583,N_783,N_4950);
xnor U10584 (N_10584,N_5763,N_1562);
nand U10585 (N_10585,N_1294,N_5579);
or U10586 (N_10586,N_2081,N_340);
nand U10587 (N_10587,N_4603,N_5093);
and U10588 (N_10588,N_5074,N_4174);
and U10589 (N_10589,N_721,N_1794);
nor U10590 (N_10590,N_1552,N_3932);
nand U10591 (N_10591,N_4429,N_5035);
nor U10592 (N_10592,N_6041,N_584);
or U10593 (N_10593,N_672,N_3864);
xor U10594 (N_10594,N_3368,N_2418);
and U10595 (N_10595,N_3084,N_1766);
xor U10596 (N_10596,N_745,N_5996);
nand U10597 (N_10597,N_144,N_5804);
and U10598 (N_10598,N_5978,N_2487);
or U10599 (N_10599,N_1723,N_2018);
nand U10600 (N_10600,N_2940,N_3850);
xnor U10601 (N_10601,N_2727,N_2013);
nor U10602 (N_10602,N_3458,N_4886);
nand U10603 (N_10603,N_5978,N_5883);
nor U10604 (N_10604,N_1016,N_3315);
nand U10605 (N_10605,N_5479,N_5853);
or U10606 (N_10606,N_2641,N_682);
nor U10607 (N_10607,N_613,N_3688);
and U10608 (N_10608,N_2893,N_1469);
xor U10609 (N_10609,N_4505,N_6184);
nand U10610 (N_10610,N_3509,N_2472);
nand U10611 (N_10611,N_1625,N_2257);
nand U10612 (N_10612,N_3986,N_5784);
nor U10613 (N_10613,N_3622,N_3020);
and U10614 (N_10614,N_3694,N_3856);
or U10615 (N_10615,N_1059,N_5615);
and U10616 (N_10616,N_3061,N_2021);
nor U10617 (N_10617,N_533,N_1253);
nor U10618 (N_10618,N_1714,N_156);
or U10619 (N_10619,N_2935,N_227);
and U10620 (N_10620,N_375,N_488);
or U10621 (N_10621,N_3926,N_1037);
and U10622 (N_10622,N_2650,N_1726);
xor U10623 (N_10623,N_3793,N_3790);
nand U10624 (N_10624,N_5548,N_1317);
or U10625 (N_10625,N_5883,N_612);
xnor U10626 (N_10626,N_3367,N_5172);
nor U10627 (N_10627,N_5287,N_3174);
xor U10628 (N_10628,N_4275,N_3770);
xnor U10629 (N_10629,N_2341,N_2089);
or U10630 (N_10630,N_2919,N_2582);
nand U10631 (N_10631,N_3363,N_3466);
xnor U10632 (N_10632,N_5079,N_2771);
xor U10633 (N_10633,N_4526,N_1502);
or U10634 (N_10634,N_518,N_206);
and U10635 (N_10635,N_1376,N_1063);
xor U10636 (N_10636,N_3358,N_5616);
xor U10637 (N_10637,N_1475,N_942);
nand U10638 (N_10638,N_1968,N_5517);
nor U10639 (N_10639,N_359,N_3687);
or U10640 (N_10640,N_4994,N_4762);
or U10641 (N_10641,N_2583,N_624);
nor U10642 (N_10642,N_1060,N_3941);
nor U10643 (N_10643,N_34,N_3626);
nand U10644 (N_10644,N_741,N_4646);
nor U10645 (N_10645,N_4505,N_1688);
or U10646 (N_10646,N_5042,N_3902);
or U10647 (N_10647,N_1030,N_935);
nor U10648 (N_10648,N_3075,N_2028);
xnor U10649 (N_10649,N_4058,N_18);
or U10650 (N_10650,N_5704,N_2236);
and U10651 (N_10651,N_4071,N_1442);
nor U10652 (N_10652,N_2883,N_1412);
xor U10653 (N_10653,N_3588,N_5123);
xnor U10654 (N_10654,N_2066,N_5844);
and U10655 (N_10655,N_4965,N_3228);
nand U10656 (N_10656,N_6034,N_5854);
or U10657 (N_10657,N_2036,N_347);
xor U10658 (N_10658,N_1808,N_3456);
and U10659 (N_10659,N_5350,N_3040);
and U10660 (N_10660,N_2665,N_3846);
nand U10661 (N_10661,N_4438,N_2228);
xnor U10662 (N_10662,N_2150,N_1746);
nor U10663 (N_10663,N_1694,N_268);
or U10664 (N_10664,N_3600,N_3192);
or U10665 (N_10665,N_3688,N_2680);
and U10666 (N_10666,N_5383,N_4848);
xor U10667 (N_10667,N_955,N_2334);
and U10668 (N_10668,N_2039,N_4241);
and U10669 (N_10669,N_3767,N_1686);
xor U10670 (N_10670,N_922,N_4058);
nor U10671 (N_10671,N_4681,N_488);
xor U10672 (N_10672,N_5216,N_5378);
xnor U10673 (N_10673,N_2747,N_1551);
and U10674 (N_10674,N_1453,N_4569);
nor U10675 (N_10675,N_2322,N_2539);
or U10676 (N_10676,N_3374,N_1656);
xor U10677 (N_10677,N_4997,N_5140);
or U10678 (N_10678,N_828,N_206);
nand U10679 (N_10679,N_2337,N_4063);
and U10680 (N_10680,N_2516,N_5991);
nor U10681 (N_10681,N_4979,N_5863);
nor U10682 (N_10682,N_1677,N_4152);
nand U10683 (N_10683,N_3662,N_3619);
and U10684 (N_10684,N_1822,N_5714);
xnor U10685 (N_10685,N_2759,N_2669);
nor U10686 (N_10686,N_124,N_2238);
nor U10687 (N_10687,N_2966,N_2558);
nor U10688 (N_10688,N_5621,N_4163);
nor U10689 (N_10689,N_3825,N_4540);
xor U10690 (N_10690,N_1146,N_1259);
nand U10691 (N_10691,N_328,N_4809);
or U10692 (N_10692,N_3382,N_1580);
nand U10693 (N_10693,N_3920,N_1650);
nand U10694 (N_10694,N_2203,N_6085);
nor U10695 (N_10695,N_4077,N_3095);
nor U10696 (N_10696,N_2235,N_3708);
or U10697 (N_10697,N_4211,N_2216);
xor U10698 (N_10698,N_2351,N_3327);
nor U10699 (N_10699,N_4458,N_3178);
and U10700 (N_10700,N_2273,N_3495);
nor U10701 (N_10701,N_5799,N_2684);
nor U10702 (N_10702,N_5652,N_3573);
xnor U10703 (N_10703,N_2233,N_2591);
nand U10704 (N_10704,N_1910,N_1880);
or U10705 (N_10705,N_4730,N_4610);
and U10706 (N_10706,N_5809,N_3514);
nor U10707 (N_10707,N_241,N_1699);
xor U10708 (N_10708,N_1199,N_3725);
or U10709 (N_10709,N_5128,N_3198);
and U10710 (N_10710,N_5819,N_5015);
xnor U10711 (N_10711,N_338,N_1279);
or U10712 (N_10712,N_4933,N_1545);
nand U10713 (N_10713,N_913,N_2230);
xor U10714 (N_10714,N_1625,N_3853);
nand U10715 (N_10715,N_199,N_2933);
nor U10716 (N_10716,N_4814,N_967);
nand U10717 (N_10717,N_1136,N_3131);
nor U10718 (N_10718,N_4714,N_4952);
and U10719 (N_10719,N_5362,N_1390);
nand U10720 (N_10720,N_2908,N_4472);
nor U10721 (N_10721,N_3187,N_3449);
nand U10722 (N_10722,N_3892,N_2123);
nand U10723 (N_10723,N_4963,N_621);
nor U10724 (N_10724,N_3994,N_422);
nor U10725 (N_10725,N_2083,N_2408);
nand U10726 (N_10726,N_5751,N_5866);
nand U10727 (N_10727,N_4008,N_5660);
nand U10728 (N_10728,N_2137,N_4393);
nor U10729 (N_10729,N_4708,N_2481);
and U10730 (N_10730,N_5803,N_104);
and U10731 (N_10731,N_5677,N_2779);
or U10732 (N_10732,N_92,N_2669);
xor U10733 (N_10733,N_5453,N_5504);
nand U10734 (N_10734,N_3784,N_3340);
nor U10735 (N_10735,N_1073,N_4978);
xnor U10736 (N_10736,N_1968,N_3753);
and U10737 (N_10737,N_5263,N_5492);
and U10738 (N_10738,N_2503,N_2487);
nor U10739 (N_10739,N_3321,N_6033);
nor U10740 (N_10740,N_4393,N_237);
xor U10741 (N_10741,N_5643,N_3351);
or U10742 (N_10742,N_806,N_3512);
and U10743 (N_10743,N_1082,N_6098);
nand U10744 (N_10744,N_986,N_5595);
xnor U10745 (N_10745,N_3158,N_1233);
nor U10746 (N_10746,N_5852,N_4242);
and U10747 (N_10747,N_4269,N_3975);
or U10748 (N_10748,N_3289,N_152);
nor U10749 (N_10749,N_4932,N_3937);
xnor U10750 (N_10750,N_5564,N_3489);
or U10751 (N_10751,N_5256,N_3938);
nand U10752 (N_10752,N_4762,N_6179);
nand U10753 (N_10753,N_6164,N_141);
or U10754 (N_10754,N_4031,N_4996);
nor U10755 (N_10755,N_5234,N_2175);
nand U10756 (N_10756,N_5127,N_2412);
nand U10757 (N_10757,N_2252,N_2007);
nand U10758 (N_10758,N_2656,N_3315);
and U10759 (N_10759,N_3634,N_2426);
nand U10760 (N_10760,N_2900,N_4788);
nand U10761 (N_10761,N_997,N_5040);
nor U10762 (N_10762,N_3852,N_869);
and U10763 (N_10763,N_4952,N_1821);
xnor U10764 (N_10764,N_918,N_1515);
or U10765 (N_10765,N_1273,N_5107);
or U10766 (N_10766,N_3875,N_4519);
nand U10767 (N_10767,N_2478,N_193);
nand U10768 (N_10768,N_3406,N_710);
and U10769 (N_10769,N_1279,N_796);
nand U10770 (N_10770,N_4012,N_4143);
and U10771 (N_10771,N_544,N_5399);
nand U10772 (N_10772,N_1421,N_5261);
or U10773 (N_10773,N_2063,N_5634);
nand U10774 (N_10774,N_3843,N_2051);
and U10775 (N_10775,N_5480,N_337);
xor U10776 (N_10776,N_2263,N_2);
and U10777 (N_10777,N_5323,N_6242);
nor U10778 (N_10778,N_60,N_4180);
and U10779 (N_10779,N_947,N_1601);
nor U10780 (N_10780,N_4444,N_5964);
xnor U10781 (N_10781,N_4347,N_1611);
nand U10782 (N_10782,N_2692,N_3886);
or U10783 (N_10783,N_2532,N_4558);
xor U10784 (N_10784,N_2273,N_4730);
xnor U10785 (N_10785,N_690,N_6017);
nand U10786 (N_10786,N_255,N_3644);
or U10787 (N_10787,N_1289,N_2993);
or U10788 (N_10788,N_2978,N_3637);
xor U10789 (N_10789,N_4732,N_5738);
xor U10790 (N_10790,N_4293,N_3519);
nor U10791 (N_10791,N_4114,N_5613);
xnor U10792 (N_10792,N_873,N_2333);
or U10793 (N_10793,N_1550,N_839);
and U10794 (N_10794,N_336,N_3970);
xnor U10795 (N_10795,N_3059,N_609);
or U10796 (N_10796,N_893,N_4114);
nand U10797 (N_10797,N_5801,N_231);
nor U10798 (N_10798,N_1839,N_2503);
nand U10799 (N_10799,N_4076,N_2694);
nor U10800 (N_10800,N_833,N_2308);
nand U10801 (N_10801,N_3999,N_5771);
nand U10802 (N_10802,N_1817,N_282);
xnor U10803 (N_10803,N_182,N_881);
nand U10804 (N_10804,N_6140,N_4346);
and U10805 (N_10805,N_3446,N_1196);
xor U10806 (N_10806,N_6005,N_4368);
nor U10807 (N_10807,N_5512,N_3782);
nor U10808 (N_10808,N_413,N_183);
nor U10809 (N_10809,N_1188,N_5923);
or U10810 (N_10810,N_889,N_5253);
or U10811 (N_10811,N_5136,N_1383);
nor U10812 (N_10812,N_4959,N_799);
nand U10813 (N_10813,N_1767,N_2495);
or U10814 (N_10814,N_4646,N_2685);
nand U10815 (N_10815,N_5187,N_2272);
xnor U10816 (N_10816,N_6204,N_2533);
nand U10817 (N_10817,N_459,N_341);
nand U10818 (N_10818,N_4456,N_5910);
nand U10819 (N_10819,N_4407,N_878);
or U10820 (N_10820,N_2085,N_6072);
nand U10821 (N_10821,N_2240,N_3825);
nor U10822 (N_10822,N_5549,N_5615);
xor U10823 (N_10823,N_6149,N_3540);
nor U10824 (N_10824,N_4592,N_145);
xnor U10825 (N_10825,N_1550,N_3314);
and U10826 (N_10826,N_5540,N_2916);
or U10827 (N_10827,N_1942,N_2632);
and U10828 (N_10828,N_4309,N_425);
and U10829 (N_10829,N_893,N_4263);
or U10830 (N_10830,N_4731,N_5778);
xor U10831 (N_10831,N_4496,N_5024);
nand U10832 (N_10832,N_248,N_3142);
nor U10833 (N_10833,N_33,N_1290);
or U10834 (N_10834,N_3420,N_3435);
xnor U10835 (N_10835,N_2541,N_1474);
or U10836 (N_10836,N_4073,N_768);
nand U10837 (N_10837,N_2235,N_301);
and U10838 (N_10838,N_5346,N_1085);
nor U10839 (N_10839,N_4621,N_1038);
or U10840 (N_10840,N_3087,N_4311);
nor U10841 (N_10841,N_2772,N_64);
nor U10842 (N_10842,N_5009,N_1874);
nor U10843 (N_10843,N_4878,N_2332);
nor U10844 (N_10844,N_712,N_5423);
nand U10845 (N_10845,N_1028,N_3014);
xnor U10846 (N_10846,N_5553,N_2788);
or U10847 (N_10847,N_625,N_2366);
xor U10848 (N_10848,N_3162,N_3067);
and U10849 (N_10849,N_6161,N_4301);
nand U10850 (N_10850,N_5147,N_5091);
nor U10851 (N_10851,N_6222,N_2031);
and U10852 (N_10852,N_6006,N_4023);
xnor U10853 (N_10853,N_259,N_191);
nand U10854 (N_10854,N_344,N_3819);
xnor U10855 (N_10855,N_5898,N_5173);
and U10856 (N_10856,N_4976,N_6212);
and U10857 (N_10857,N_5089,N_4953);
xnor U10858 (N_10858,N_2748,N_1287);
or U10859 (N_10859,N_1163,N_3094);
and U10860 (N_10860,N_3693,N_3194);
and U10861 (N_10861,N_5229,N_5145);
nor U10862 (N_10862,N_3261,N_3206);
and U10863 (N_10863,N_4042,N_3227);
and U10864 (N_10864,N_4723,N_3943);
nand U10865 (N_10865,N_3657,N_4589);
or U10866 (N_10866,N_208,N_4062);
nand U10867 (N_10867,N_4489,N_2843);
nor U10868 (N_10868,N_6177,N_2656);
or U10869 (N_10869,N_453,N_4029);
nand U10870 (N_10870,N_3135,N_5446);
or U10871 (N_10871,N_4876,N_917);
nor U10872 (N_10872,N_3937,N_3972);
nor U10873 (N_10873,N_3814,N_4934);
and U10874 (N_10874,N_620,N_717);
nor U10875 (N_10875,N_3653,N_1125);
nor U10876 (N_10876,N_963,N_2817);
or U10877 (N_10877,N_2126,N_2641);
nand U10878 (N_10878,N_3600,N_303);
xnor U10879 (N_10879,N_1220,N_5627);
or U10880 (N_10880,N_2227,N_4172);
or U10881 (N_10881,N_992,N_5927);
nor U10882 (N_10882,N_1675,N_3529);
and U10883 (N_10883,N_936,N_710);
and U10884 (N_10884,N_2526,N_5754);
nor U10885 (N_10885,N_4596,N_3112);
xor U10886 (N_10886,N_2366,N_3128);
nor U10887 (N_10887,N_5516,N_2148);
nor U10888 (N_10888,N_2526,N_5089);
and U10889 (N_10889,N_6013,N_4282);
nand U10890 (N_10890,N_602,N_421);
or U10891 (N_10891,N_5270,N_4076);
nand U10892 (N_10892,N_3853,N_5453);
and U10893 (N_10893,N_3745,N_3899);
xnor U10894 (N_10894,N_1976,N_6042);
xnor U10895 (N_10895,N_4758,N_3650);
and U10896 (N_10896,N_2979,N_4145);
and U10897 (N_10897,N_2698,N_464);
or U10898 (N_10898,N_5154,N_4721);
nor U10899 (N_10899,N_2545,N_2082);
or U10900 (N_10900,N_817,N_3118);
xnor U10901 (N_10901,N_6123,N_5350);
nor U10902 (N_10902,N_1291,N_5081);
xnor U10903 (N_10903,N_5238,N_61);
nand U10904 (N_10904,N_216,N_2226);
xor U10905 (N_10905,N_804,N_6036);
xor U10906 (N_10906,N_807,N_3143);
nor U10907 (N_10907,N_4673,N_5102);
xor U10908 (N_10908,N_1591,N_2888);
and U10909 (N_10909,N_1423,N_4197);
or U10910 (N_10910,N_1426,N_1766);
xor U10911 (N_10911,N_2931,N_4772);
xor U10912 (N_10912,N_5130,N_982);
or U10913 (N_10913,N_5844,N_5388);
xor U10914 (N_10914,N_4599,N_4188);
nor U10915 (N_10915,N_1387,N_1193);
and U10916 (N_10916,N_700,N_3853);
nor U10917 (N_10917,N_964,N_443);
xor U10918 (N_10918,N_2615,N_4423);
or U10919 (N_10919,N_3618,N_1697);
xnor U10920 (N_10920,N_4535,N_905);
and U10921 (N_10921,N_2416,N_5819);
nor U10922 (N_10922,N_5895,N_5916);
or U10923 (N_10923,N_3125,N_607);
or U10924 (N_10924,N_4596,N_4776);
and U10925 (N_10925,N_4222,N_678);
xnor U10926 (N_10926,N_1283,N_2965);
and U10927 (N_10927,N_4736,N_5348);
and U10928 (N_10928,N_180,N_2731);
and U10929 (N_10929,N_2698,N_1480);
nor U10930 (N_10930,N_2112,N_1900);
xnor U10931 (N_10931,N_782,N_1975);
xor U10932 (N_10932,N_744,N_6083);
and U10933 (N_10933,N_4315,N_5623);
or U10934 (N_10934,N_1168,N_637);
and U10935 (N_10935,N_5890,N_3000);
or U10936 (N_10936,N_3542,N_817);
xor U10937 (N_10937,N_2882,N_1843);
xor U10938 (N_10938,N_3520,N_3517);
nand U10939 (N_10939,N_5461,N_2479);
nand U10940 (N_10940,N_4963,N_150);
nand U10941 (N_10941,N_4052,N_1186);
or U10942 (N_10942,N_303,N_5283);
nor U10943 (N_10943,N_2732,N_3263);
xor U10944 (N_10944,N_5896,N_4900);
xor U10945 (N_10945,N_328,N_2477);
or U10946 (N_10946,N_404,N_4965);
nor U10947 (N_10947,N_4256,N_543);
nand U10948 (N_10948,N_3711,N_3358);
nor U10949 (N_10949,N_4512,N_462);
and U10950 (N_10950,N_691,N_830);
or U10951 (N_10951,N_83,N_959);
nand U10952 (N_10952,N_1609,N_501);
nand U10953 (N_10953,N_3013,N_5352);
or U10954 (N_10954,N_785,N_6003);
or U10955 (N_10955,N_5917,N_1012);
nand U10956 (N_10956,N_2863,N_677);
nand U10957 (N_10957,N_5547,N_2364);
xnor U10958 (N_10958,N_4184,N_4448);
xor U10959 (N_10959,N_3738,N_3201);
xnor U10960 (N_10960,N_4941,N_6214);
and U10961 (N_10961,N_5590,N_2516);
nand U10962 (N_10962,N_5842,N_4666);
nand U10963 (N_10963,N_5610,N_1602);
nor U10964 (N_10964,N_1895,N_2235);
or U10965 (N_10965,N_3990,N_2614);
and U10966 (N_10966,N_3941,N_2557);
nand U10967 (N_10967,N_6044,N_1764);
xor U10968 (N_10968,N_3806,N_5977);
nand U10969 (N_10969,N_239,N_4782);
nor U10970 (N_10970,N_3165,N_5294);
and U10971 (N_10971,N_6206,N_2333);
nor U10972 (N_10972,N_2882,N_3383);
nand U10973 (N_10973,N_549,N_6139);
nor U10974 (N_10974,N_326,N_5879);
nor U10975 (N_10975,N_1120,N_505);
nor U10976 (N_10976,N_278,N_773);
nand U10977 (N_10977,N_3632,N_4923);
and U10978 (N_10978,N_5025,N_5432);
and U10979 (N_10979,N_233,N_3315);
and U10980 (N_10980,N_3457,N_4743);
xor U10981 (N_10981,N_5613,N_918);
and U10982 (N_10982,N_3924,N_3075);
nand U10983 (N_10983,N_2353,N_4933);
or U10984 (N_10984,N_5566,N_102);
or U10985 (N_10985,N_2104,N_2710);
nor U10986 (N_10986,N_4906,N_207);
or U10987 (N_10987,N_3213,N_5950);
xnor U10988 (N_10988,N_2505,N_1406);
xor U10989 (N_10989,N_3734,N_2654);
nand U10990 (N_10990,N_3053,N_4384);
and U10991 (N_10991,N_1244,N_1894);
nand U10992 (N_10992,N_2800,N_3013);
or U10993 (N_10993,N_2851,N_107);
xor U10994 (N_10994,N_4949,N_4409);
nand U10995 (N_10995,N_4518,N_2215);
nor U10996 (N_10996,N_628,N_2178);
or U10997 (N_10997,N_2761,N_1401);
nand U10998 (N_10998,N_5761,N_18);
xnor U10999 (N_10999,N_1516,N_4786);
nand U11000 (N_11000,N_2754,N_2545);
nand U11001 (N_11001,N_5933,N_5461);
nor U11002 (N_11002,N_5172,N_4794);
nor U11003 (N_11003,N_2846,N_3176);
or U11004 (N_11004,N_4916,N_4833);
nand U11005 (N_11005,N_5187,N_24);
or U11006 (N_11006,N_3104,N_3741);
nand U11007 (N_11007,N_1613,N_3316);
and U11008 (N_11008,N_3238,N_4366);
or U11009 (N_11009,N_1581,N_2932);
and U11010 (N_11010,N_1254,N_5534);
or U11011 (N_11011,N_1827,N_3305);
nor U11012 (N_11012,N_5469,N_1858);
and U11013 (N_11013,N_4091,N_2018);
nor U11014 (N_11014,N_4024,N_2020);
and U11015 (N_11015,N_1852,N_2485);
nor U11016 (N_11016,N_4419,N_4649);
nor U11017 (N_11017,N_2119,N_164);
nor U11018 (N_11018,N_748,N_5614);
nor U11019 (N_11019,N_5173,N_5425);
xnor U11020 (N_11020,N_4262,N_2640);
and U11021 (N_11021,N_1982,N_4709);
xnor U11022 (N_11022,N_6022,N_3625);
nor U11023 (N_11023,N_5978,N_5455);
nand U11024 (N_11024,N_5966,N_5405);
and U11025 (N_11025,N_4295,N_3408);
xnor U11026 (N_11026,N_2166,N_967);
or U11027 (N_11027,N_182,N_4435);
xor U11028 (N_11028,N_1607,N_3061);
nor U11029 (N_11029,N_1081,N_5860);
or U11030 (N_11030,N_3263,N_1962);
nand U11031 (N_11031,N_5276,N_3615);
or U11032 (N_11032,N_964,N_1302);
xor U11033 (N_11033,N_2306,N_5511);
and U11034 (N_11034,N_4693,N_3049);
or U11035 (N_11035,N_1664,N_2088);
nor U11036 (N_11036,N_4402,N_1337);
or U11037 (N_11037,N_670,N_4431);
or U11038 (N_11038,N_5906,N_6035);
nor U11039 (N_11039,N_2918,N_3589);
or U11040 (N_11040,N_5204,N_4982);
and U11041 (N_11041,N_1522,N_6070);
xnor U11042 (N_11042,N_4864,N_1697);
nand U11043 (N_11043,N_5827,N_4428);
or U11044 (N_11044,N_1492,N_2877);
nand U11045 (N_11045,N_1044,N_5174);
xnor U11046 (N_11046,N_2816,N_4672);
and U11047 (N_11047,N_4064,N_3998);
nand U11048 (N_11048,N_5575,N_1861);
nand U11049 (N_11049,N_3008,N_1737);
and U11050 (N_11050,N_6152,N_2802);
nor U11051 (N_11051,N_4872,N_5258);
xnor U11052 (N_11052,N_2280,N_895);
xor U11053 (N_11053,N_1072,N_128);
nand U11054 (N_11054,N_1568,N_4267);
and U11055 (N_11055,N_5181,N_5323);
xnor U11056 (N_11056,N_1455,N_3442);
nand U11057 (N_11057,N_2007,N_1471);
nor U11058 (N_11058,N_3119,N_1499);
nand U11059 (N_11059,N_5313,N_5325);
xor U11060 (N_11060,N_5346,N_3057);
or U11061 (N_11061,N_2225,N_4330);
nand U11062 (N_11062,N_3141,N_377);
or U11063 (N_11063,N_1194,N_143);
and U11064 (N_11064,N_2800,N_3116);
or U11065 (N_11065,N_4079,N_5063);
or U11066 (N_11066,N_680,N_1305);
and U11067 (N_11067,N_5886,N_5539);
nor U11068 (N_11068,N_3388,N_700);
nand U11069 (N_11069,N_4116,N_3711);
nand U11070 (N_11070,N_3631,N_326);
nor U11071 (N_11071,N_4068,N_372);
nand U11072 (N_11072,N_4420,N_5240);
xor U11073 (N_11073,N_5564,N_112);
and U11074 (N_11074,N_6015,N_3515);
nor U11075 (N_11075,N_1044,N_3635);
xnor U11076 (N_11076,N_5009,N_3344);
and U11077 (N_11077,N_2172,N_5941);
and U11078 (N_11078,N_60,N_4041);
and U11079 (N_11079,N_3559,N_2707);
or U11080 (N_11080,N_4493,N_5581);
nand U11081 (N_11081,N_2378,N_5964);
nand U11082 (N_11082,N_2396,N_5648);
and U11083 (N_11083,N_1934,N_1480);
and U11084 (N_11084,N_3376,N_3950);
nor U11085 (N_11085,N_4006,N_175);
or U11086 (N_11086,N_624,N_4270);
and U11087 (N_11087,N_1458,N_2851);
nand U11088 (N_11088,N_4457,N_1687);
xnor U11089 (N_11089,N_1531,N_3975);
xor U11090 (N_11090,N_2033,N_3009);
nand U11091 (N_11091,N_4872,N_3563);
nor U11092 (N_11092,N_394,N_3409);
nand U11093 (N_11093,N_154,N_1851);
or U11094 (N_11094,N_3408,N_2512);
and U11095 (N_11095,N_647,N_2319);
and U11096 (N_11096,N_1161,N_2079);
or U11097 (N_11097,N_1985,N_3829);
nand U11098 (N_11098,N_3728,N_4085);
xnor U11099 (N_11099,N_443,N_4499);
nand U11100 (N_11100,N_2947,N_3840);
nand U11101 (N_11101,N_5994,N_5031);
nand U11102 (N_11102,N_4900,N_1110);
nand U11103 (N_11103,N_2340,N_6056);
or U11104 (N_11104,N_1762,N_5357);
and U11105 (N_11105,N_4986,N_288);
and U11106 (N_11106,N_6090,N_3738);
and U11107 (N_11107,N_267,N_4042);
nand U11108 (N_11108,N_246,N_1044);
nor U11109 (N_11109,N_5860,N_3870);
and U11110 (N_11110,N_1864,N_941);
or U11111 (N_11111,N_1678,N_5033);
and U11112 (N_11112,N_946,N_5558);
nor U11113 (N_11113,N_915,N_5386);
or U11114 (N_11114,N_50,N_2235);
or U11115 (N_11115,N_448,N_998);
nand U11116 (N_11116,N_3747,N_1332);
nand U11117 (N_11117,N_5429,N_3676);
and U11118 (N_11118,N_2063,N_2226);
xnor U11119 (N_11119,N_4435,N_3415);
nand U11120 (N_11120,N_3865,N_5564);
xnor U11121 (N_11121,N_1024,N_2388);
nor U11122 (N_11122,N_4015,N_6139);
or U11123 (N_11123,N_5728,N_5676);
or U11124 (N_11124,N_2870,N_4912);
nand U11125 (N_11125,N_57,N_2604);
nand U11126 (N_11126,N_1985,N_1801);
xnor U11127 (N_11127,N_1476,N_1336);
or U11128 (N_11128,N_1734,N_778);
and U11129 (N_11129,N_5508,N_4393);
nor U11130 (N_11130,N_4290,N_4709);
nor U11131 (N_11131,N_4005,N_1345);
and U11132 (N_11132,N_4740,N_3248);
nor U11133 (N_11133,N_5810,N_5086);
nor U11134 (N_11134,N_1624,N_3456);
nand U11135 (N_11135,N_5836,N_323);
xor U11136 (N_11136,N_5199,N_3208);
nor U11137 (N_11137,N_2920,N_2657);
xor U11138 (N_11138,N_4267,N_5337);
nand U11139 (N_11139,N_1776,N_733);
nand U11140 (N_11140,N_744,N_1387);
nor U11141 (N_11141,N_4983,N_1750);
nand U11142 (N_11142,N_4444,N_1463);
and U11143 (N_11143,N_5584,N_166);
or U11144 (N_11144,N_4283,N_5485);
or U11145 (N_11145,N_2417,N_1960);
xnor U11146 (N_11146,N_405,N_5716);
nor U11147 (N_11147,N_2935,N_5136);
xor U11148 (N_11148,N_3440,N_5169);
and U11149 (N_11149,N_4275,N_651);
nor U11150 (N_11150,N_3363,N_348);
and U11151 (N_11151,N_1653,N_4087);
and U11152 (N_11152,N_4973,N_3834);
nand U11153 (N_11153,N_630,N_1312);
xnor U11154 (N_11154,N_1792,N_864);
and U11155 (N_11155,N_5769,N_4817);
and U11156 (N_11156,N_6146,N_5810);
xnor U11157 (N_11157,N_6014,N_2602);
nand U11158 (N_11158,N_1992,N_2928);
xor U11159 (N_11159,N_12,N_759);
nor U11160 (N_11160,N_2257,N_3370);
and U11161 (N_11161,N_3846,N_4636);
and U11162 (N_11162,N_4220,N_297);
or U11163 (N_11163,N_4471,N_3468);
or U11164 (N_11164,N_930,N_1475);
nor U11165 (N_11165,N_3410,N_5353);
and U11166 (N_11166,N_2589,N_1599);
and U11167 (N_11167,N_5576,N_2724);
nand U11168 (N_11168,N_1664,N_4371);
and U11169 (N_11169,N_3137,N_72);
and U11170 (N_11170,N_3272,N_1045);
or U11171 (N_11171,N_5376,N_721);
xor U11172 (N_11172,N_2535,N_1122);
and U11173 (N_11173,N_5635,N_4149);
nor U11174 (N_11174,N_2159,N_210);
and U11175 (N_11175,N_728,N_4218);
nand U11176 (N_11176,N_2571,N_4013);
xor U11177 (N_11177,N_5355,N_480);
nand U11178 (N_11178,N_2438,N_3198);
nor U11179 (N_11179,N_2054,N_2079);
nor U11180 (N_11180,N_2467,N_4944);
xnor U11181 (N_11181,N_5491,N_4815);
or U11182 (N_11182,N_5859,N_4201);
and U11183 (N_11183,N_1025,N_5369);
xnor U11184 (N_11184,N_2000,N_4699);
or U11185 (N_11185,N_6215,N_3237);
nand U11186 (N_11186,N_2208,N_2992);
nand U11187 (N_11187,N_4579,N_3064);
nand U11188 (N_11188,N_2913,N_1547);
xnor U11189 (N_11189,N_4775,N_2647);
xnor U11190 (N_11190,N_2238,N_81);
and U11191 (N_11191,N_3257,N_704);
or U11192 (N_11192,N_2462,N_1136);
or U11193 (N_11193,N_4128,N_5488);
nor U11194 (N_11194,N_2208,N_2191);
nor U11195 (N_11195,N_3531,N_393);
or U11196 (N_11196,N_2432,N_5283);
or U11197 (N_11197,N_3899,N_1747);
and U11198 (N_11198,N_3414,N_3965);
xnor U11199 (N_11199,N_1893,N_1259);
nor U11200 (N_11200,N_4649,N_2074);
nor U11201 (N_11201,N_866,N_5814);
nand U11202 (N_11202,N_684,N_3577);
or U11203 (N_11203,N_2921,N_4531);
nor U11204 (N_11204,N_3067,N_342);
and U11205 (N_11205,N_2609,N_6040);
nand U11206 (N_11206,N_4548,N_2594);
nand U11207 (N_11207,N_725,N_795);
or U11208 (N_11208,N_3594,N_4986);
nand U11209 (N_11209,N_668,N_5270);
and U11210 (N_11210,N_6188,N_3291);
xnor U11211 (N_11211,N_2614,N_3666);
nand U11212 (N_11212,N_1036,N_2161);
nor U11213 (N_11213,N_3695,N_1120);
nand U11214 (N_11214,N_4362,N_3617);
and U11215 (N_11215,N_4949,N_4125);
xnor U11216 (N_11216,N_3391,N_1688);
xor U11217 (N_11217,N_2857,N_4915);
and U11218 (N_11218,N_849,N_3352);
nand U11219 (N_11219,N_2160,N_2960);
and U11220 (N_11220,N_184,N_2110);
nor U11221 (N_11221,N_5745,N_4860);
and U11222 (N_11222,N_5235,N_3751);
nand U11223 (N_11223,N_2489,N_4451);
or U11224 (N_11224,N_1613,N_75);
or U11225 (N_11225,N_5005,N_2886);
xor U11226 (N_11226,N_1338,N_1763);
nor U11227 (N_11227,N_1996,N_4088);
nand U11228 (N_11228,N_5739,N_3451);
xor U11229 (N_11229,N_6229,N_6231);
nand U11230 (N_11230,N_928,N_5060);
and U11231 (N_11231,N_3932,N_5848);
or U11232 (N_11232,N_135,N_5162);
nand U11233 (N_11233,N_3718,N_4962);
nand U11234 (N_11234,N_3037,N_3171);
nor U11235 (N_11235,N_2071,N_731);
and U11236 (N_11236,N_1122,N_5294);
and U11237 (N_11237,N_282,N_5903);
or U11238 (N_11238,N_2203,N_4472);
or U11239 (N_11239,N_199,N_4006);
nor U11240 (N_11240,N_5237,N_4285);
nor U11241 (N_11241,N_4233,N_3133);
nor U11242 (N_11242,N_1519,N_1409);
nor U11243 (N_11243,N_124,N_3296);
and U11244 (N_11244,N_3282,N_2403);
nor U11245 (N_11245,N_1531,N_4141);
or U11246 (N_11246,N_2145,N_2926);
nand U11247 (N_11247,N_1184,N_6022);
and U11248 (N_11248,N_986,N_5783);
nor U11249 (N_11249,N_4957,N_3882);
nand U11250 (N_11250,N_1091,N_5549);
nor U11251 (N_11251,N_5005,N_1230);
nand U11252 (N_11252,N_5864,N_1000);
nor U11253 (N_11253,N_1475,N_239);
nor U11254 (N_11254,N_4722,N_3806);
and U11255 (N_11255,N_302,N_1392);
and U11256 (N_11256,N_4835,N_609);
or U11257 (N_11257,N_795,N_2503);
nand U11258 (N_11258,N_5156,N_955);
nand U11259 (N_11259,N_2393,N_2148);
xor U11260 (N_11260,N_2855,N_1795);
and U11261 (N_11261,N_1220,N_1847);
and U11262 (N_11262,N_4974,N_10);
nor U11263 (N_11263,N_6132,N_1321);
or U11264 (N_11264,N_3319,N_1891);
or U11265 (N_11265,N_3847,N_235);
nor U11266 (N_11266,N_123,N_6032);
and U11267 (N_11267,N_1406,N_1493);
nor U11268 (N_11268,N_169,N_1693);
and U11269 (N_11269,N_5522,N_2929);
nor U11270 (N_11270,N_5776,N_5424);
or U11271 (N_11271,N_6001,N_3908);
nand U11272 (N_11272,N_5999,N_1368);
or U11273 (N_11273,N_5013,N_2803);
and U11274 (N_11274,N_3276,N_1572);
and U11275 (N_11275,N_6004,N_5693);
and U11276 (N_11276,N_2480,N_3720);
and U11277 (N_11277,N_1727,N_571);
xnor U11278 (N_11278,N_4850,N_3827);
xnor U11279 (N_11279,N_2725,N_370);
xnor U11280 (N_11280,N_3243,N_719);
or U11281 (N_11281,N_3823,N_3896);
nor U11282 (N_11282,N_2798,N_1825);
xor U11283 (N_11283,N_1881,N_2419);
nand U11284 (N_11284,N_1021,N_5985);
nor U11285 (N_11285,N_6212,N_2592);
and U11286 (N_11286,N_1895,N_1346);
xor U11287 (N_11287,N_5827,N_4458);
and U11288 (N_11288,N_2039,N_4274);
nand U11289 (N_11289,N_1944,N_1850);
nand U11290 (N_11290,N_3007,N_1872);
and U11291 (N_11291,N_5142,N_2877);
nand U11292 (N_11292,N_3163,N_581);
or U11293 (N_11293,N_3847,N_3797);
or U11294 (N_11294,N_4715,N_392);
xnor U11295 (N_11295,N_5541,N_5876);
xor U11296 (N_11296,N_4912,N_4703);
nor U11297 (N_11297,N_1234,N_4283);
nand U11298 (N_11298,N_2668,N_1618);
nor U11299 (N_11299,N_4019,N_899);
and U11300 (N_11300,N_3867,N_1540);
nor U11301 (N_11301,N_6114,N_2873);
and U11302 (N_11302,N_5227,N_4477);
and U11303 (N_11303,N_1854,N_4188);
nor U11304 (N_11304,N_5490,N_1678);
nor U11305 (N_11305,N_245,N_3480);
xor U11306 (N_11306,N_2310,N_5602);
or U11307 (N_11307,N_1135,N_2820);
and U11308 (N_11308,N_4799,N_1853);
and U11309 (N_11309,N_3538,N_3380);
nor U11310 (N_11310,N_1905,N_4396);
or U11311 (N_11311,N_1746,N_5728);
nor U11312 (N_11312,N_1001,N_1951);
and U11313 (N_11313,N_2392,N_444);
or U11314 (N_11314,N_1920,N_127);
nand U11315 (N_11315,N_1123,N_3672);
and U11316 (N_11316,N_1713,N_2621);
and U11317 (N_11317,N_3250,N_5137);
xor U11318 (N_11318,N_4996,N_543);
and U11319 (N_11319,N_480,N_5431);
nand U11320 (N_11320,N_3344,N_1655);
and U11321 (N_11321,N_4577,N_738);
xnor U11322 (N_11322,N_3074,N_4188);
nor U11323 (N_11323,N_4249,N_4545);
nand U11324 (N_11324,N_1267,N_5520);
and U11325 (N_11325,N_5598,N_5587);
or U11326 (N_11326,N_3962,N_1183);
xor U11327 (N_11327,N_3747,N_3272);
and U11328 (N_11328,N_4129,N_2371);
and U11329 (N_11329,N_4688,N_5990);
nand U11330 (N_11330,N_2600,N_1854);
nor U11331 (N_11331,N_544,N_1545);
or U11332 (N_11332,N_5102,N_462);
nand U11333 (N_11333,N_3629,N_1249);
nor U11334 (N_11334,N_5317,N_4052);
xnor U11335 (N_11335,N_3762,N_1830);
and U11336 (N_11336,N_4341,N_5872);
and U11337 (N_11337,N_411,N_938);
xor U11338 (N_11338,N_4852,N_4371);
nand U11339 (N_11339,N_5010,N_3711);
and U11340 (N_11340,N_989,N_2265);
nand U11341 (N_11341,N_4859,N_4423);
nand U11342 (N_11342,N_4894,N_3911);
nand U11343 (N_11343,N_2296,N_5674);
nand U11344 (N_11344,N_6151,N_1336);
nor U11345 (N_11345,N_1760,N_4714);
and U11346 (N_11346,N_4386,N_2547);
and U11347 (N_11347,N_5559,N_3384);
and U11348 (N_11348,N_3498,N_3349);
or U11349 (N_11349,N_5463,N_1622);
nor U11350 (N_11350,N_4027,N_3025);
and U11351 (N_11351,N_1603,N_2773);
and U11352 (N_11352,N_108,N_931);
nand U11353 (N_11353,N_1921,N_1116);
nand U11354 (N_11354,N_1941,N_2709);
xnor U11355 (N_11355,N_5494,N_2649);
nor U11356 (N_11356,N_2521,N_5223);
or U11357 (N_11357,N_3942,N_356);
and U11358 (N_11358,N_2614,N_3418);
and U11359 (N_11359,N_628,N_792);
and U11360 (N_11360,N_2234,N_3492);
nor U11361 (N_11361,N_2051,N_2638);
or U11362 (N_11362,N_5067,N_2273);
or U11363 (N_11363,N_4021,N_5702);
or U11364 (N_11364,N_3271,N_3771);
nor U11365 (N_11365,N_2614,N_2716);
nor U11366 (N_11366,N_3082,N_2241);
and U11367 (N_11367,N_3275,N_5098);
nand U11368 (N_11368,N_4091,N_1420);
nand U11369 (N_11369,N_5177,N_444);
nand U11370 (N_11370,N_5192,N_3636);
nand U11371 (N_11371,N_2759,N_3501);
and U11372 (N_11372,N_2878,N_1364);
xnor U11373 (N_11373,N_5281,N_6038);
nor U11374 (N_11374,N_810,N_3116);
nor U11375 (N_11375,N_3612,N_2765);
xnor U11376 (N_11376,N_5671,N_5780);
nand U11377 (N_11377,N_5272,N_2450);
and U11378 (N_11378,N_3400,N_3194);
or U11379 (N_11379,N_5536,N_4349);
nor U11380 (N_11380,N_1452,N_1502);
or U11381 (N_11381,N_466,N_4353);
nor U11382 (N_11382,N_559,N_502);
nand U11383 (N_11383,N_4439,N_5295);
nand U11384 (N_11384,N_3243,N_1789);
nand U11385 (N_11385,N_2637,N_1711);
or U11386 (N_11386,N_4744,N_5241);
nor U11387 (N_11387,N_1551,N_1220);
xnor U11388 (N_11388,N_1521,N_5436);
nand U11389 (N_11389,N_1525,N_4796);
xnor U11390 (N_11390,N_879,N_2497);
xnor U11391 (N_11391,N_4295,N_3149);
nor U11392 (N_11392,N_100,N_5837);
xnor U11393 (N_11393,N_2500,N_968);
and U11394 (N_11394,N_2558,N_449);
nand U11395 (N_11395,N_4917,N_2648);
and U11396 (N_11396,N_2550,N_3171);
xor U11397 (N_11397,N_2138,N_4613);
nand U11398 (N_11398,N_4839,N_923);
and U11399 (N_11399,N_156,N_583);
nor U11400 (N_11400,N_4306,N_5180);
xnor U11401 (N_11401,N_2742,N_5675);
nor U11402 (N_11402,N_2068,N_3661);
or U11403 (N_11403,N_6180,N_4912);
and U11404 (N_11404,N_5139,N_2276);
nor U11405 (N_11405,N_1042,N_1661);
nand U11406 (N_11406,N_1682,N_5542);
nor U11407 (N_11407,N_2907,N_3018);
or U11408 (N_11408,N_4334,N_3820);
or U11409 (N_11409,N_553,N_1712);
and U11410 (N_11410,N_5310,N_492);
xor U11411 (N_11411,N_2176,N_506);
xnor U11412 (N_11412,N_5924,N_5923);
nand U11413 (N_11413,N_857,N_114);
nor U11414 (N_11414,N_4566,N_6078);
xnor U11415 (N_11415,N_2982,N_5358);
nand U11416 (N_11416,N_3087,N_4537);
nand U11417 (N_11417,N_3574,N_5638);
or U11418 (N_11418,N_5020,N_3666);
xnor U11419 (N_11419,N_4580,N_2801);
nand U11420 (N_11420,N_5299,N_1445);
nand U11421 (N_11421,N_5194,N_4193);
nand U11422 (N_11422,N_3396,N_6112);
xor U11423 (N_11423,N_5539,N_1537);
nor U11424 (N_11424,N_848,N_1776);
xnor U11425 (N_11425,N_2077,N_3787);
or U11426 (N_11426,N_2493,N_1640);
and U11427 (N_11427,N_4570,N_4839);
nor U11428 (N_11428,N_328,N_2558);
or U11429 (N_11429,N_3688,N_1325);
nor U11430 (N_11430,N_3506,N_1649);
or U11431 (N_11431,N_5755,N_30);
and U11432 (N_11432,N_753,N_1532);
nor U11433 (N_11433,N_2699,N_1446);
or U11434 (N_11434,N_4693,N_1302);
xor U11435 (N_11435,N_582,N_2006);
and U11436 (N_11436,N_3186,N_3801);
and U11437 (N_11437,N_3368,N_5616);
and U11438 (N_11438,N_2479,N_4161);
or U11439 (N_11439,N_1707,N_1174);
or U11440 (N_11440,N_389,N_3689);
xnor U11441 (N_11441,N_5642,N_4452);
and U11442 (N_11442,N_2735,N_5108);
or U11443 (N_11443,N_2884,N_5873);
and U11444 (N_11444,N_2514,N_1265);
nor U11445 (N_11445,N_1610,N_1052);
or U11446 (N_11446,N_3397,N_1379);
or U11447 (N_11447,N_2861,N_936);
nor U11448 (N_11448,N_2388,N_2605);
nand U11449 (N_11449,N_24,N_1748);
nand U11450 (N_11450,N_3576,N_5975);
nor U11451 (N_11451,N_3958,N_2387);
xor U11452 (N_11452,N_3676,N_319);
nor U11453 (N_11453,N_900,N_5716);
nor U11454 (N_11454,N_126,N_2845);
nand U11455 (N_11455,N_848,N_1356);
or U11456 (N_11456,N_2412,N_3302);
and U11457 (N_11457,N_1313,N_508);
xor U11458 (N_11458,N_5005,N_1625);
and U11459 (N_11459,N_1763,N_2536);
nand U11460 (N_11460,N_2042,N_3397);
and U11461 (N_11461,N_1551,N_2325);
or U11462 (N_11462,N_4855,N_5590);
or U11463 (N_11463,N_4966,N_3983);
or U11464 (N_11464,N_292,N_3353);
nor U11465 (N_11465,N_2198,N_4118);
or U11466 (N_11466,N_1624,N_4343);
or U11467 (N_11467,N_826,N_139);
xnor U11468 (N_11468,N_2572,N_5270);
nand U11469 (N_11469,N_6125,N_4086);
xnor U11470 (N_11470,N_3134,N_128);
nor U11471 (N_11471,N_987,N_4788);
nand U11472 (N_11472,N_1565,N_852);
xor U11473 (N_11473,N_865,N_4498);
and U11474 (N_11474,N_1264,N_2231);
nand U11475 (N_11475,N_2885,N_4953);
or U11476 (N_11476,N_892,N_2353);
and U11477 (N_11477,N_5146,N_2314);
and U11478 (N_11478,N_180,N_1551);
or U11479 (N_11479,N_1911,N_3475);
xnor U11480 (N_11480,N_3721,N_3486);
or U11481 (N_11481,N_5963,N_531);
nor U11482 (N_11482,N_3379,N_1569);
xor U11483 (N_11483,N_5929,N_5841);
xor U11484 (N_11484,N_5588,N_1896);
and U11485 (N_11485,N_2008,N_803);
nand U11486 (N_11486,N_4068,N_443);
nand U11487 (N_11487,N_33,N_1350);
xor U11488 (N_11488,N_2675,N_883);
nand U11489 (N_11489,N_3563,N_2555);
or U11490 (N_11490,N_441,N_2497);
nand U11491 (N_11491,N_4968,N_6038);
and U11492 (N_11492,N_1178,N_1782);
and U11493 (N_11493,N_1657,N_4819);
nor U11494 (N_11494,N_4056,N_6249);
nand U11495 (N_11495,N_4753,N_5415);
nor U11496 (N_11496,N_506,N_4713);
nor U11497 (N_11497,N_2608,N_1137);
nor U11498 (N_11498,N_999,N_2608);
and U11499 (N_11499,N_3196,N_3330);
nor U11500 (N_11500,N_3696,N_3852);
nand U11501 (N_11501,N_6164,N_2185);
xnor U11502 (N_11502,N_2307,N_3630);
nand U11503 (N_11503,N_844,N_6197);
and U11504 (N_11504,N_3623,N_2975);
nand U11505 (N_11505,N_1083,N_2911);
or U11506 (N_11506,N_1827,N_1079);
or U11507 (N_11507,N_5582,N_3661);
nor U11508 (N_11508,N_3035,N_1864);
or U11509 (N_11509,N_4148,N_524);
nand U11510 (N_11510,N_5729,N_3668);
xor U11511 (N_11511,N_3597,N_5154);
nand U11512 (N_11512,N_850,N_5197);
nor U11513 (N_11513,N_2028,N_1873);
xnor U11514 (N_11514,N_3204,N_3863);
nand U11515 (N_11515,N_755,N_3383);
and U11516 (N_11516,N_5629,N_1367);
and U11517 (N_11517,N_1812,N_4621);
nand U11518 (N_11518,N_1935,N_5207);
and U11519 (N_11519,N_6248,N_4063);
or U11520 (N_11520,N_5550,N_3178);
nand U11521 (N_11521,N_2373,N_2248);
xnor U11522 (N_11522,N_1435,N_5074);
nand U11523 (N_11523,N_953,N_1723);
and U11524 (N_11524,N_5594,N_2449);
nor U11525 (N_11525,N_1577,N_1256);
xnor U11526 (N_11526,N_3977,N_161);
xnor U11527 (N_11527,N_3014,N_4122);
nor U11528 (N_11528,N_2556,N_4945);
and U11529 (N_11529,N_5366,N_6028);
and U11530 (N_11530,N_146,N_2858);
and U11531 (N_11531,N_3667,N_6207);
or U11532 (N_11532,N_2469,N_3689);
or U11533 (N_11533,N_6172,N_112);
nand U11534 (N_11534,N_436,N_2186);
or U11535 (N_11535,N_1024,N_6211);
nand U11536 (N_11536,N_5126,N_4418);
nor U11537 (N_11537,N_1099,N_3526);
nand U11538 (N_11538,N_2571,N_2117);
and U11539 (N_11539,N_4070,N_4590);
xor U11540 (N_11540,N_3023,N_2925);
and U11541 (N_11541,N_1047,N_2590);
and U11542 (N_11542,N_2563,N_5139);
nor U11543 (N_11543,N_1376,N_2872);
xnor U11544 (N_11544,N_4603,N_250);
or U11545 (N_11545,N_1570,N_3711);
or U11546 (N_11546,N_5172,N_2439);
nand U11547 (N_11547,N_3434,N_5140);
or U11548 (N_11548,N_3373,N_4283);
xor U11549 (N_11549,N_3494,N_267);
and U11550 (N_11550,N_1370,N_969);
nor U11551 (N_11551,N_2573,N_6189);
and U11552 (N_11552,N_1961,N_3078);
or U11553 (N_11553,N_1388,N_4890);
xnor U11554 (N_11554,N_2956,N_1000);
nor U11555 (N_11555,N_4340,N_478);
xnor U11556 (N_11556,N_1482,N_903);
or U11557 (N_11557,N_2215,N_3559);
nor U11558 (N_11558,N_3538,N_3359);
and U11559 (N_11559,N_2230,N_288);
xor U11560 (N_11560,N_3881,N_4494);
and U11561 (N_11561,N_1616,N_2456);
or U11562 (N_11562,N_5538,N_1511);
and U11563 (N_11563,N_3332,N_2848);
xnor U11564 (N_11564,N_5491,N_2996);
xnor U11565 (N_11565,N_4767,N_6159);
nor U11566 (N_11566,N_1148,N_2082);
and U11567 (N_11567,N_5011,N_3900);
or U11568 (N_11568,N_4934,N_181);
nor U11569 (N_11569,N_2279,N_4918);
or U11570 (N_11570,N_3989,N_4738);
nand U11571 (N_11571,N_3498,N_3627);
nor U11572 (N_11572,N_3325,N_4149);
and U11573 (N_11573,N_2506,N_5916);
nand U11574 (N_11574,N_3296,N_4830);
nor U11575 (N_11575,N_2691,N_5942);
or U11576 (N_11576,N_2738,N_293);
and U11577 (N_11577,N_2649,N_2213);
and U11578 (N_11578,N_262,N_475);
and U11579 (N_11579,N_4890,N_5977);
and U11580 (N_11580,N_3703,N_4547);
or U11581 (N_11581,N_6017,N_3343);
and U11582 (N_11582,N_2274,N_4788);
nor U11583 (N_11583,N_2025,N_3905);
and U11584 (N_11584,N_1345,N_3639);
and U11585 (N_11585,N_595,N_877);
or U11586 (N_11586,N_3326,N_2407);
and U11587 (N_11587,N_5114,N_6030);
xnor U11588 (N_11588,N_520,N_5308);
nor U11589 (N_11589,N_121,N_3978);
or U11590 (N_11590,N_1543,N_3750);
or U11591 (N_11591,N_2186,N_1891);
nor U11592 (N_11592,N_4177,N_2590);
or U11593 (N_11593,N_58,N_5248);
and U11594 (N_11594,N_3371,N_1571);
xnor U11595 (N_11595,N_32,N_4758);
nand U11596 (N_11596,N_3700,N_180);
or U11597 (N_11597,N_3807,N_5522);
xor U11598 (N_11598,N_4714,N_2078);
nand U11599 (N_11599,N_4963,N_5582);
or U11600 (N_11600,N_3435,N_3615);
xor U11601 (N_11601,N_3059,N_3583);
or U11602 (N_11602,N_5716,N_3927);
nand U11603 (N_11603,N_2207,N_3105);
nand U11604 (N_11604,N_2857,N_690);
nor U11605 (N_11605,N_1832,N_908);
nand U11606 (N_11606,N_4302,N_71);
xor U11607 (N_11607,N_5996,N_4913);
or U11608 (N_11608,N_5305,N_3496);
or U11609 (N_11609,N_1292,N_688);
or U11610 (N_11610,N_5866,N_591);
nand U11611 (N_11611,N_3270,N_4002);
nand U11612 (N_11612,N_4654,N_5751);
or U11613 (N_11613,N_5527,N_1006);
xor U11614 (N_11614,N_4330,N_3374);
or U11615 (N_11615,N_4488,N_3670);
or U11616 (N_11616,N_502,N_1126);
and U11617 (N_11617,N_2647,N_5593);
nor U11618 (N_11618,N_3203,N_5488);
xor U11619 (N_11619,N_2365,N_2923);
xnor U11620 (N_11620,N_2494,N_2999);
or U11621 (N_11621,N_5818,N_2121);
nor U11622 (N_11622,N_3027,N_2549);
and U11623 (N_11623,N_253,N_4300);
or U11624 (N_11624,N_3704,N_2436);
or U11625 (N_11625,N_4956,N_2638);
xnor U11626 (N_11626,N_4265,N_899);
xnor U11627 (N_11627,N_595,N_5128);
and U11628 (N_11628,N_5021,N_515);
and U11629 (N_11629,N_2675,N_1761);
and U11630 (N_11630,N_5483,N_1651);
xnor U11631 (N_11631,N_1264,N_4838);
and U11632 (N_11632,N_6059,N_4539);
nor U11633 (N_11633,N_842,N_5958);
and U11634 (N_11634,N_3656,N_6188);
nor U11635 (N_11635,N_1117,N_2540);
and U11636 (N_11636,N_2619,N_6074);
nor U11637 (N_11637,N_4306,N_4173);
and U11638 (N_11638,N_947,N_1176);
or U11639 (N_11639,N_1387,N_4471);
or U11640 (N_11640,N_1996,N_4126);
nand U11641 (N_11641,N_1971,N_5191);
and U11642 (N_11642,N_2035,N_2826);
nand U11643 (N_11643,N_1292,N_2136);
nor U11644 (N_11644,N_1012,N_548);
nand U11645 (N_11645,N_1358,N_1236);
and U11646 (N_11646,N_4185,N_3978);
xnor U11647 (N_11647,N_744,N_5461);
xnor U11648 (N_11648,N_5123,N_5303);
and U11649 (N_11649,N_4878,N_1524);
or U11650 (N_11650,N_3718,N_5509);
nand U11651 (N_11651,N_5476,N_4527);
or U11652 (N_11652,N_2638,N_542);
and U11653 (N_11653,N_2205,N_5064);
and U11654 (N_11654,N_104,N_1713);
and U11655 (N_11655,N_948,N_2126);
or U11656 (N_11656,N_5525,N_5760);
nor U11657 (N_11657,N_5381,N_3832);
nand U11658 (N_11658,N_2800,N_2286);
nand U11659 (N_11659,N_1129,N_5513);
nand U11660 (N_11660,N_46,N_3335);
nor U11661 (N_11661,N_5752,N_3504);
nand U11662 (N_11662,N_1096,N_3597);
nand U11663 (N_11663,N_5674,N_4232);
xnor U11664 (N_11664,N_964,N_3854);
xor U11665 (N_11665,N_479,N_3906);
nor U11666 (N_11666,N_3914,N_6094);
nand U11667 (N_11667,N_3602,N_2665);
and U11668 (N_11668,N_3562,N_3510);
and U11669 (N_11669,N_4842,N_1107);
and U11670 (N_11670,N_265,N_1960);
or U11671 (N_11671,N_816,N_5182);
nand U11672 (N_11672,N_1895,N_1740);
xor U11673 (N_11673,N_773,N_3512);
nor U11674 (N_11674,N_2428,N_1182);
or U11675 (N_11675,N_4882,N_4900);
nand U11676 (N_11676,N_2374,N_5);
and U11677 (N_11677,N_3847,N_5070);
nand U11678 (N_11678,N_1513,N_817);
or U11679 (N_11679,N_4196,N_4799);
xnor U11680 (N_11680,N_2867,N_2683);
or U11681 (N_11681,N_1374,N_660);
nor U11682 (N_11682,N_3159,N_3957);
or U11683 (N_11683,N_4147,N_4652);
nor U11684 (N_11684,N_665,N_565);
or U11685 (N_11685,N_4681,N_3780);
nor U11686 (N_11686,N_601,N_3000);
xnor U11687 (N_11687,N_3669,N_4071);
and U11688 (N_11688,N_851,N_6238);
nand U11689 (N_11689,N_2931,N_790);
xnor U11690 (N_11690,N_6033,N_1663);
nand U11691 (N_11691,N_4856,N_4628);
nor U11692 (N_11692,N_5389,N_5944);
or U11693 (N_11693,N_3234,N_1375);
xor U11694 (N_11694,N_1128,N_1573);
nand U11695 (N_11695,N_59,N_467);
xnor U11696 (N_11696,N_961,N_4206);
nand U11697 (N_11697,N_4601,N_5019);
or U11698 (N_11698,N_3656,N_1220);
nand U11699 (N_11699,N_3874,N_2690);
or U11700 (N_11700,N_2064,N_3440);
nand U11701 (N_11701,N_274,N_2857);
nor U11702 (N_11702,N_3401,N_345);
nand U11703 (N_11703,N_1518,N_5470);
nor U11704 (N_11704,N_1280,N_1972);
or U11705 (N_11705,N_2339,N_6248);
nand U11706 (N_11706,N_2834,N_717);
nor U11707 (N_11707,N_672,N_2017);
xor U11708 (N_11708,N_5518,N_3358);
xnor U11709 (N_11709,N_4799,N_5018);
nand U11710 (N_11710,N_4638,N_1837);
xor U11711 (N_11711,N_1499,N_3048);
nand U11712 (N_11712,N_613,N_3133);
nor U11713 (N_11713,N_2569,N_2570);
or U11714 (N_11714,N_1674,N_4445);
and U11715 (N_11715,N_2270,N_1733);
or U11716 (N_11716,N_5920,N_5880);
nand U11717 (N_11717,N_4549,N_5023);
or U11718 (N_11718,N_2433,N_3081);
or U11719 (N_11719,N_332,N_2107);
nor U11720 (N_11720,N_3595,N_2066);
or U11721 (N_11721,N_1626,N_4838);
and U11722 (N_11722,N_1209,N_1459);
or U11723 (N_11723,N_705,N_4109);
nor U11724 (N_11724,N_907,N_2371);
and U11725 (N_11725,N_2657,N_5658);
or U11726 (N_11726,N_2127,N_1431);
xnor U11727 (N_11727,N_3975,N_724);
xnor U11728 (N_11728,N_5572,N_1582);
nand U11729 (N_11729,N_6205,N_803);
or U11730 (N_11730,N_5967,N_5238);
xor U11731 (N_11731,N_1415,N_5984);
nand U11732 (N_11732,N_26,N_4062);
or U11733 (N_11733,N_3320,N_2842);
xor U11734 (N_11734,N_2933,N_5729);
nand U11735 (N_11735,N_4438,N_3265);
xor U11736 (N_11736,N_4737,N_1236);
or U11737 (N_11737,N_5993,N_4596);
nand U11738 (N_11738,N_1287,N_2784);
nor U11739 (N_11739,N_2152,N_273);
or U11740 (N_11740,N_2466,N_749);
and U11741 (N_11741,N_1121,N_4751);
xnor U11742 (N_11742,N_317,N_5416);
or U11743 (N_11743,N_4721,N_477);
nor U11744 (N_11744,N_6195,N_4461);
nand U11745 (N_11745,N_2148,N_718);
nand U11746 (N_11746,N_1256,N_6221);
xor U11747 (N_11747,N_86,N_5145);
xor U11748 (N_11748,N_5780,N_5606);
xor U11749 (N_11749,N_794,N_3897);
xnor U11750 (N_11750,N_806,N_4779);
or U11751 (N_11751,N_4472,N_1085);
nor U11752 (N_11752,N_589,N_2392);
nor U11753 (N_11753,N_1933,N_5196);
nand U11754 (N_11754,N_5721,N_5338);
and U11755 (N_11755,N_4302,N_1405);
or U11756 (N_11756,N_4748,N_2145);
or U11757 (N_11757,N_1170,N_1038);
or U11758 (N_11758,N_5911,N_3872);
or U11759 (N_11759,N_1507,N_3914);
or U11760 (N_11760,N_5379,N_6182);
nand U11761 (N_11761,N_2214,N_709);
and U11762 (N_11762,N_5138,N_565);
or U11763 (N_11763,N_2163,N_884);
xnor U11764 (N_11764,N_2650,N_3977);
and U11765 (N_11765,N_3846,N_3377);
nand U11766 (N_11766,N_4655,N_1324);
xnor U11767 (N_11767,N_5393,N_1087);
or U11768 (N_11768,N_3334,N_4509);
or U11769 (N_11769,N_2090,N_288);
and U11770 (N_11770,N_5258,N_557);
xnor U11771 (N_11771,N_980,N_6182);
nand U11772 (N_11772,N_4369,N_2540);
and U11773 (N_11773,N_677,N_5297);
or U11774 (N_11774,N_5092,N_3293);
or U11775 (N_11775,N_3444,N_517);
nand U11776 (N_11776,N_1437,N_459);
nor U11777 (N_11777,N_5287,N_1730);
or U11778 (N_11778,N_3604,N_4379);
nand U11779 (N_11779,N_2946,N_858);
nand U11780 (N_11780,N_369,N_5830);
and U11781 (N_11781,N_4528,N_761);
nor U11782 (N_11782,N_284,N_3017);
or U11783 (N_11783,N_4382,N_2238);
and U11784 (N_11784,N_3689,N_3560);
or U11785 (N_11785,N_311,N_3168);
nor U11786 (N_11786,N_4733,N_5340);
nor U11787 (N_11787,N_1919,N_92);
nand U11788 (N_11788,N_457,N_1991);
nor U11789 (N_11789,N_6185,N_5976);
nor U11790 (N_11790,N_4589,N_107);
nor U11791 (N_11791,N_5672,N_4481);
and U11792 (N_11792,N_1529,N_5679);
nand U11793 (N_11793,N_5925,N_4252);
and U11794 (N_11794,N_4541,N_1464);
or U11795 (N_11795,N_3956,N_4203);
and U11796 (N_11796,N_263,N_4898);
xnor U11797 (N_11797,N_5556,N_5323);
xnor U11798 (N_11798,N_2533,N_2662);
nand U11799 (N_11799,N_2281,N_4946);
nor U11800 (N_11800,N_4223,N_5761);
xnor U11801 (N_11801,N_4263,N_4289);
or U11802 (N_11802,N_4467,N_4924);
xor U11803 (N_11803,N_477,N_5156);
or U11804 (N_11804,N_3341,N_5736);
nor U11805 (N_11805,N_2679,N_1419);
nor U11806 (N_11806,N_3712,N_3976);
nor U11807 (N_11807,N_3074,N_125);
and U11808 (N_11808,N_115,N_1393);
or U11809 (N_11809,N_5280,N_1246);
and U11810 (N_11810,N_2860,N_249);
xor U11811 (N_11811,N_1498,N_3393);
nor U11812 (N_11812,N_4627,N_4471);
or U11813 (N_11813,N_5923,N_1171);
xor U11814 (N_11814,N_2239,N_4183);
nand U11815 (N_11815,N_2713,N_5613);
and U11816 (N_11816,N_808,N_4248);
or U11817 (N_11817,N_3205,N_5614);
xnor U11818 (N_11818,N_4270,N_5292);
or U11819 (N_11819,N_4530,N_5674);
xor U11820 (N_11820,N_2652,N_1409);
and U11821 (N_11821,N_3581,N_2456);
nor U11822 (N_11822,N_2148,N_2128);
nand U11823 (N_11823,N_4108,N_620);
nand U11824 (N_11824,N_1508,N_2523);
xnor U11825 (N_11825,N_525,N_5695);
nand U11826 (N_11826,N_3074,N_2333);
nand U11827 (N_11827,N_3116,N_3109);
nand U11828 (N_11828,N_5394,N_1400);
xor U11829 (N_11829,N_2933,N_169);
and U11830 (N_11830,N_5626,N_3058);
nand U11831 (N_11831,N_4000,N_3280);
and U11832 (N_11832,N_5360,N_210);
xor U11833 (N_11833,N_5607,N_5337);
xor U11834 (N_11834,N_843,N_2190);
and U11835 (N_11835,N_5793,N_5223);
and U11836 (N_11836,N_558,N_33);
xor U11837 (N_11837,N_2466,N_3458);
xnor U11838 (N_11838,N_120,N_3312);
nor U11839 (N_11839,N_2629,N_4105);
and U11840 (N_11840,N_5589,N_4455);
xnor U11841 (N_11841,N_1254,N_3070);
and U11842 (N_11842,N_1918,N_4347);
xnor U11843 (N_11843,N_343,N_2158);
and U11844 (N_11844,N_2905,N_3068);
xnor U11845 (N_11845,N_4541,N_4319);
and U11846 (N_11846,N_2559,N_4809);
xor U11847 (N_11847,N_5145,N_4643);
nor U11848 (N_11848,N_6219,N_1299);
and U11849 (N_11849,N_3458,N_1345);
xor U11850 (N_11850,N_673,N_257);
nor U11851 (N_11851,N_4507,N_1458);
and U11852 (N_11852,N_5367,N_3825);
nor U11853 (N_11853,N_370,N_3161);
xor U11854 (N_11854,N_5014,N_973);
nor U11855 (N_11855,N_1934,N_3131);
xnor U11856 (N_11856,N_2530,N_5391);
nand U11857 (N_11857,N_2741,N_3932);
nor U11858 (N_11858,N_4664,N_1607);
or U11859 (N_11859,N_3042,N_4826);
nand U11860 (N_11860,N_3394,N_5760);
and U11861 (N_11861,N_2264,N_4521);
xnor U11862 (N_11862,N_3301,N_202);
nand U11863 (N_11863,N_1910,N_2587);
xor U11864 (N_11864,N_402,N_4787);
nand U11865 (N_11865,N_3608,N_2721);
and U11866 (N_11866,N_1199,N_614);
xor U11867 (N_11867,N_1219,N_6141);
xnor U11868 (N_11868,N_5403,N_1529);
or U11869 (N_11869,N_2215,N_2308);
nand U11870 (N_11870,N_2303,N_3303);
nand U11871 (N_11871,N_543,N_932);
nand U11872 (N_11872,N_2610,N_2982);
or U11873 (N_11873,N_588,N_4470);
xnor U11874 (N_11874,N_4999,N_2536);
and U11875 (N_11875,N_2586,N_2454);
nand U11876 (N_11876,N_1019,N_790);
xnor U11877 (N_11877,N_2513,N_2382);
or U11878 (N_11878,N_155,N_5713);
xor U11879 (N_11879,N_2796,N_1092);
and U11880 (N_11880,N_2374,N_2567);
nand U11881 (N_11881,N_5792,N_5577);
xnor U11882 (N_11882,N_2193,N_2297);
and U11883 (N_11883,N_352,N_5573);
or U11884 (N_11884,N_5389,N_3784);
nand U11885 (N_11885,N_4313,N_1404);
nor U11886 (N_11886,N_5945,N_92);
nand U11887 (N_11887,N_1741,N_3592);
or U11888 (N_11888,N_5933,N_4797);
and U11889 (N_11889,N_1492,N_3007);
or U11890 (N_11890,N_1323,N_3204);
or U11891 (N_11891,N_1108,N_2514);
and U11892 (N_11892,N_4874,N_3645);
or U11893 (N_11893,N_4977,N_5274);
or U11894 (N_11894,N_1439,N_4500);
nor U11895 (N_11895,N_320,N_5646);
xor U11896 (N_11896,N_1781,N_4579);
nand U11897 (N_11897,N_79,N_1438);
nor U11898 (N_11898,N_879,N_5049);
nand U11899 (N_11899,N_3803,N_1543);
xnor U11900 (N_11900,N_4322,N_6071);
xnor U11901 (N_11901,N_1659,N_547);
or U11902 (N_11902,N_4843,N_1497);
or U11903 (N_11903,N_4078,N_481);
nand U11904 (N_11904,N_521,N_3681);
nand U11905 (N_11905,N_482,N_3815);
nor U11906 (N_11906,N_4289,N_4012);
nor U11907 (N_11907,N_3259,N_2997);
nor U11908 (N_11908,N_4475,N_3712);
nand U11909 (N_11909,N_497,N_460);
xnor U11910 (N_11910,N_4501,N_3845);
xor U11911 (N_11911,N_301,N_3496);
xnor U11912 (N_11912,N_3074,N_3084);
and U11913 (N_11913,N_2339,N_149);
or U11914 (N_11914,N_3753,N_96);
nand U11915 (N_11915,N_5504,N_2246);
or U11916 (N_11916,N_3896,N_3474);
nand U11917 (N_11917,N_4322,N_3243);
xnor U11918 (N_11918,N_2638,N_5999);
and U11919 (N_11919,N_2791,N_1133);
nand U11920 (N_11920,N_4019,N_1195);
xnor U11921 (N_11921,N_3589,N_872);
and U11922 (N_11922,N_5309,N_3927);
xor U11923 (N_11923,N_6094,N_4554);
and U11924 (N_11924,N_1374,N_2004);
nor U11925 (N_11925,N_2659,N_1164);
or U11926 (N_11926,N_1331,N_5292);
and U11927 (N_11927,N_4509,N_4917);
xor U11928 (N_11928,N_381,N_3990);
nor U11929 (N_11929,N_188,N_335);
and U11930 (N_11930,N_2023,N_3034);
xnor U11931 (N_11931,N_4853,N_5037);
and U11932 (N_11932,N_1630,N_3488);
nand U11933 (N_11933,N_5400,N_4915);
or U11934 (N_11934,N_202,N_3102);
nand U11935 (N_11935,N_2078,N_2250);
or U11936 (N_11936,N_5096,N_4911);
nor U11937 (N_11937,N_5598,N_5896);
and U11938 (N_11938,N_5029,N_4352);
or U11939 (N_11939,N_5904,N_5396);
nor U11940 (N_11940,N_2392,N_5604);
nand U11941 (N_11941,N_89,N_2114);
and U11942 (N_11942,N_49,N_5985);
nor U11943 (N_11943,N_3237,N_383);
xnor U11944 (N_11944,N_4180,N_287);
or U11945 (N_11945,N_1097,N_1722);
nand U11946 (N_11946,N_4878,N_3221);
xnor U11947 (N_11947,N_4776,N_3193);
nand U11948 (N_11948,N_5765,N_2599);
nand U11949 (N_11949,N_2940,N_3071);
and U11950 (N_11950,N_5234,N_2149);
and U11951 (N_11951,N_1781,N_5219);
or U11952 (N_11952,N_1778,N_5365);
nand U11953 (N_11953,N_5507,N_5550);
or U11954 (N_11954,N_2714,N_2370);
or U11955 (N_11955,N_1323,N_2582);
or U11956 (N_11956,N_3984,N_5455);
nand U11957 (N_11957,N_956,N_6155);
nor U11958 (N_11958,N_4755,N_305);
and U11959 (N_11959,N_1419,N_104);
or U11960 (N_11960,N_5262,N_4573);
or U11961 (N_11961,N_2992,N_619);
nor U11962 (N_11962,N_4343,N_928);
and U11963 (N_11963,N_5533,N_4602);
xor U11964 (N_11964,N_50,N_1267);
nor U11965 (N_11965,N_4631,N_418);
and U11966 (N_11966,N_2547,N_59);
nand U11967 (N_11967,N_5599,N_122);
nor U11968 (N_11968,N_36,N_3546);
and U11969 (N_11969,N_292,N_5814);
xnor U11970 (N_11970,N_3740,N_5417);
or U11971 (N_11971,N_3459,N_989);
nand U11972 (N_11972,N_6013,N_1050);
nor U11973 (N_11973,N_1293,N_1414);
nor U11974 (N_11974,N_1842,N_1699);
xnor U11975 (N_11975,N_3616,N_2860);
or U11976 (N_11976,N_5015,N_1101);
and U11977 (N_11977,N_1216,N_5191);
and U11978 (N_11978,N_5852,N_4385);
xnor U11979 (N_11979,N_4504,N_264);
nand U11980 (N_11980,N_2716,N_2148);
and U11981 (N_11981,N_1768,N_1451);
xnor U11982 (N_11982,N_772,N_1102);
nor U11983 (N_11983,N_4541,N_5475);
nor U11984 (N_11984,N_4150,N_3354);
and U11985 (N_11985,N_5311,N_2309);
xor U11986 (N_11986,N_1812,N_6163);
and U11987 (N_11987,N_1538,N_3744);
xnor U11988 (N_11988,N_4214,N_1345);
xnor U11989 (N_11989,N_9,N_103);
and U11990 (N_11990,N_6198,N_5421);
nor U11991 (N_11991,N_2795,N_5770);
nor U11992 (N_11992,N_5908,N_6123);
xnor U11993 (N_11993,N_16,N_3985);
or U11994 (N_11994,N_2445,N_4838);
xnor U11995 (N_11995,N_101,N_5253);
xnor U11996 (N_11996,N_2662,N_1687);
xnor U11997 (N_11997,N_5434,N_27);
nand U11998 (N_11998,N_2877,N_4044);
nand U11999 (N_11999,N_267,N_143);
xnor U12000 (N_12000,N_4716,N_3457);
xnor U12001 (N_12001,N_5636,N_4587);
xor U12002 (N_12002,N_372,N_2576);
or U12003 (N_12003,N_283,N_1166);
nand U12004 (N_12004,N_3494,N_1386);
or U12005 (N_12005,N_4714,N_2588);
and U12006 (N_12006,N_2155,N_1928);
nand U12007 (N_12007,N_1084,N_1961);
xor U12008 (N_12008,N_2803,N_4750);
nand U12009 (N_12009,N_3325,N_5015);
and U12010 (N_12010,N_126,N_5490);
and U12011 (N_12011,N_3419,N_5819);
nand U12012 (N_12012,N_4794,N_6242);
xor U12013 (N_12013,N_875,N_5670);
nand U12014 (N_12014,N_2078,N_1479);
nor U12015 (N_12015,N_1652,N_5119);
and U12016 (N_12016,N_2614,N_1972);
xor U12017 (N_12017,N_4555,N_2509);
and U12018 (N_12018,N_3983,N_5557);
or U12019 (N_12019,N_5108,N_538);
nand U12020 (N_12020,N_3213,N_2460);
nor U12021 (N_12021,N_637,N_3178);
and U12022 (N_12022,N_3487,N_1717);
xnor U12023 (N_12023,N_5862,N_2280);
xnor U12024 (N_12024,N_5528,N_3212);
nand U12025 (N_12025,N_112,N_5651);
and U12026 (N_12026,N_2252,N_2331);
nor U12027 (N_12027,N_2877,N_6134);
and U12028 (N_12028,N_1545,N_1918);
xor U12029 (N_12029,N_384,N_5260);
nand U12030 (N_12030,N_722,N_70);
nand U12031 (N_12031,N_2707,N_1466);
nand U12032 (N_12032,N_2801,N_4285);
or U12033 (N_12033,N_722,N_1294);
nor U12034 (N_12034,N_476,N_3865);
nand U12035 (N_12035,N_1505,N_142);
or U12036 (N_12036,N_4283,N_2334);
or U12037 (N_12037,N_4749,N_2867);
or U12038 (N_12038,N_2552,N_477);
nand U12039 (N_12039,N_455,N_5005);
nand U12040 (N_12040,N_3846,N_4100);
or U12041 (N_12041,N_179,N_791);
nand U12042 (N_12042,N_3715,N_3944);
xor U12043 (N_12043,N_893,N_2856);
or U12044 (N_12044,N_695,N_1778);
and U12045 (N_12045,N_969,N_4120);
or U12046 (N_12046,N_2622,N_111);
nand U12047 (N_12047,N_3795,N_3567);
xnor U12048 (N_12048,N_1908,N_2154);
or U12049 (N_12049,N_5385,N_3458);
or U12050 (N_12050,N_5933,N_1632);
and U12051 (N_12051,N_2657,N_890);
nor U12052 (N_12052,N_5852,N_1185);
or U12053 (N_12053,N_835,N_1851);
and U12054 (N_12054,N_1384,N_5019);
or U12055 (N_12055,N_2545,N_1532);
and U12056 (N_12056,N_2737,N_5965);
nand U12057 (N_12057,N_4146,N_1656);
nor U12058 (N_12058,N_4287,N_3762);
and U12059 (N_12059,N_5743,N_1789);
or U12060 (N_12060,N_945,N_1957);
nor U12061 (N_12061,N_2482,N_2609);
nand U12062 (N_12062,N_4453,N_5768);
and U12063 (N_12063,N_2365,N_601);
nand U12064 (N_12064,N_5291,N_4328);
or U12065 (N_12065,N_137,N_1899);
xnor U12066 (N_12066,N_4185,N_3226);
and U12067 (N_12067,N_5896,N_4865);
nand U12068 (N_12068,N_5111,N_5213);
nor U12069 (N_12069,N_3874,N_1521);
nor U12070 (N_12070,N_1528,N_4569);
or U12071 (N_12071,N_1701,N_5259);
nand U12072 (N_12072,N_5570,N_436);
or U12073 (N_12073,N_2472,N_5352);
or U12074 (N_12074,N_1024,N_2405);
nor U12075 (N_12075,N_1,N_5901);
or U12076 (N_12076,N_1426,N_2362);
or U12077 (N_12077,N_1004,N_1153);
and U12078 (N_12078,N_2332,N_1199);
or U12079 (N_12079,N_5595,N_1867);
nor U12080 (N_12080,N_2471,N_2725);
and U12081 (N_12081,N_3331,N_2213);
nor U12082 (N_12082,N_697,N_2228);
nand U12083 (N_12083,N_1055,N_2406);
nor U12084 (N_12084,N_704,N_2362);
xnor U12085 (N_12085,N_2117,N_5953);
xnor U12086 (N_12086,N_3742,N_2286);
nor U12087 (N_12087,N_3380,N_3548);
xor U12088 (N_12088,N_5686,N_65);
or U12089 (N_12089,N_5268,N_4799);
nand U12090 (N_12090,N_2870,N_0);
nor U12091 (N_12091,N_4657,N_2810);
and U12092 (N_12092,N_5331,N_525);
or U12093 (N_12093,N_5028,N_4747);
nand U12094 (N_12094,N_559,N_5707);
and U12095 (N_12095,N_1399,N_1456);
and U12096 (N_12096,N_1363,N_1462);
nand U12097 (N_12097,N_151,N_5269);
xnor U12098 (N_12098,N_2367,N_2954);
and U12099 (N_12099,N_3650,N_5369);
or U12100 (N_12100,N_1743,N_1336);
xor U12101 (N_12101,N_2685,N_78);
or U12102 (N_12102,N_1328,N_129);
nor U12103 (N_12103,N_3570,N_6045);
nand U12104 (N_12104,N_4077,N_3293);
or U12105 (N_12105,N_3546,N_6086);
or U12106 (N_12106,N_2049,N_2716);
and U12107 (N_12107,N_3247,N_1503);
xor U12108 (N_12108,N_1787,N_4956);
nand U12109 (N_12109,N_101,N_4604);
xor U12110 (N_12110,N_634,N_5589);
or U12111 (N_12111,N_3993,N_393);
xnor U12112 (N_12112,N_2225,N_1399);
or U12113 (N_12113,N_3337,N_5994);
nand U12114 (N_12114,N_501,N_466);
or U12115 (N_12115,N_3428,N_4517);
nand U12116 (N_12116,N_1698,N_5065);
xnor U12117 (N_12117,N_5317,N_1022);
or U12118 (N_12118,N_4349,N_6141);
and U12119 (N_12119,N_1598,N_4725);
or U12120 (N_12120,N_1483,N_6053);
or U12121 (N_12121,N_2414,N_158);
and U12122 (N_12122,N_6062,N_370);
nor U12123 (N_12123,N_5912,N_3862);
nand U12124 (N_12124,N_4335,N_2446);
nor U12125 (N_12125,N_1295,N_4058);
and U12126 (N_12126,N_2912,N_5518);
xnor U12127 (N_12127,N_4178,N_7);
nand U12128 (N_12128,N_3818,N_5863);
nor U12129 (N_12129,N_2323,N_4501);
xnor U12130 (N_12130,N_5739,N_1435);
and U12131 (N_12131,N_2077,N_620);
or U12132 (N_12132,N_235,N_3979);
nand U12133 (N_12133,N_4945,N_2501);
or U12134 (N_12134,N_836,N_1830);
or U12135 (N_12135,N_2889,N_1980);
or U12136 (N_12136,N_5639,N_1167);
xnor U12137 (N_12137,N_3035,N_495);
or U12138 (N_12138,N_47,N_3505);
nand U12139 (N_12139,N_4577,N_254);
nand U12140 (N_12140,N_6171,N_885);
nand U12141 (N_12141,N_5681,N_3609);
and U12142 (N_12142,N_3000,N_3011);
nand U12143 (N_12143,N_1250,N_559);
nand U12144 (N_12144,N_5403,N_6148);
nand U12145 (N_12145,N_3593,N_5416);
xnor U12146 (N_12146,N_5605,N_1010);
xor U12147 (N_12147,N_2515,N_3522);
xnor U12148 (N_12148,N_2754,N_3293);
and U12149 (N_12149,N_4291,N_3808);
xnor U12150 (N_12150,N_5211,N_1129);
or U12151 (N_12151,N_5487,N_4551);
or U12152 (N_12152,N_1522,N_3086);
or U12153 (N_12153,N_5918,N_5808);
or U12154 (N_12154,N_4468,N_3022);
nand U12155 (N_12155,N_1146,N_4270);
nor U12156 (N_12156,N_3239,N_3586);
nor U12157 (N_12157,N_1892,N_1499);
or U12158 (N_12158,N_3921,N_2004);
nand U12159 (N_12159,N_5860,N_5859);
and U12160 (N_12160,N_150,N_255);
and U12161 (N_12161,N_2122,N_5380);
and U12162 (N_12162,N_179,N_5498);
nor U12163 (N_12163,N_2869,N_4351);
or U12164 (N_12164,N_5927,N_3311);
xnor U12165 (N_12165,N_2613,N_4850);
nand U12166 (N_12166,N_2117,N_857);
xor U12167 (N_12167,N_2733,N_3342);
nand U12168 (N_12168,N_4915,N_1340);
or U12169 (N_12169,N_958,N_5856);
nand U12170 (N_12170,N_5835,N_3312);
nor U12171 (N_12171,N_1253,N_4837);
and U12172 (N_12172,N_4787,N_5781);
nand U12173 (N_12173,N_653,N_4793);
or U12174 (N_12174,N_4190,N_1720);
xnor U12175 (N_12175,N_1517,N_704);
nor U12176 (N_12176,N_3474,N_3402);
xnor U12177 (N_12177,N_4169,N_4181);
nor U12178 (N_12178,N_2610,N_2803);
nand U12179 (N_12179,N_2648,N_4808);
nor U12180 (N_12180,N_6186,N_3414);
nor U12181 (N_12181,N_2208,N_4620);
or U12182 (N_12182,N_2196,N_4435);
xor U12183 (N_12183,N_6023,N_5677);
or U12184 (N_12184,N_6087,N_3633);
nand U12185 (N_12185,N_1850,N_4985);
nand U12186 (N_12186,N_1415,N_1326);
nor U12187 (N_12187,N_844,N_251);
or U12188 (N_12188,N_2880,N_1310);
nor U12189 (N_12189,N_338,N_5740);
nor U12190 (N_12190,N_3009,N_4480);
or U12191 (N_12191,N_4078,N_1179);
and U12192 (N_12192,N_73,N_3438);
nand U12193 (N_12193,N_3648,N_4630);
nand U12194 (N_12194,N_417,N_4885);
nand U12195 (N_12195,N_4189,N_2968);
nand U12196 (N_12196,N_3182,N_847);
nor U12197 (N_12197,N_5485,N_4535);
or U12198 (N_12198,N_2857,N_3212);
nor U12199 (N_12199,N_2531,N_2774);
and U12200 (N_12200,N_2607,N_2673);
or U12201 (N_12201,N_1129,N_225);
xnor U12202 (N_12202,N_5768,N_4851);
nand U12203 (N_12203,N_2187,N_674);
nand U12204 (N_12204,N_3880,N_3504);
and U12205 (N_12205,N_2396,N_657);
nor U12206 (N_12206,N_5598,N_5093);
xor U12207 (N_12207,N_4010,N_2336);
xnor U12208 (N_12208,N_3950,N_5376);
nand U12209 (N_12209,N_4223,N_5046);
nor U12210 (N_12210,N_527,N_361);
xnor U12211 (N_12211,N_2965,N_2375);
nand U12212 (N_12212,N_1354,N_4631);
or U12213 (N_12213,N_1067,N_2165);
and U12214 (N_12214,N_3503,N_2108);
or U12215 (N_12215,N_5992,N_4686);
xor U12216 (N_12216,N_4314,N_6242);
and U12217 (N_12217,N_1977,N_2043);
xor U12218 (N_12218,N_4166,N_5975);
xor U12219 (N_12219,N_3807,N_2618);
nor U12220 (N_12220,N_3092,N_1561);
xnor U12221 (N_12221,N_4608,N_5853);
xor U12222 (N_12222,N_3911,N_4518);
nand U12223 (N_12223,N_3525,N_2176);
xnor U12224 (N_12224,N_369,N_2675);
and U12225 (N_12225,N_186,N_5955);
and U12226 (N_12226,N_5119,N_6162);
or U12227 (N_12227,N_1243,N_2626);
or U12228 (N_12228,N_5308,N_506);
and U12229 (N_12229,N_1299,N_5795);
and U12230 (N_12230,N_325,N_5993);
and U12231 (N_12231,N_5738,N_3126);
and U12232 (N_12232,N_1235,N_5692);
or U12233 (N_12233,N_3922,N_6089);
nor U12234 (N_12234,N_1902,N_1019);
nand U12235 (N_12235,N_3766,N_1679);
nand U12236 (N_12236,N_5654,N_4132);
and U12237 (N_12237,N_4790,N_4297);
and U12238 (N_12238,N_3985,N_2944);
and U12239 (N_12239,N_918,N_3995);
nor U12240 (N_12240,N_2963,N_5784);
nand U12241 (N_12241,N_3131,N_2886);
nor U12242 (N_12242,N_3661,N_2462);
and U12243 (N_12243,N_5786,N_6209);
nand U12244 (N_12244,N_4307,N_4348);
and U12245 (N_12245,N_5811,N_6109);
nor U12246 (N_12246,N_5658,N_349);
or U12247 (N_12247,N_4405,N_5988);
xnor U12248 (N_12248,N_4370,N_4909);
nand U12249 (N_12249,N_812,N_5931);
and U12250 (N_12250,N_4246,N_2204);
and U12251 (N_12251,N_1580,N_5315);
xor U12252 (N_12252,N_1745,N_3635);
nand U12253 (N_12253,N_60,N_2493);
and U12254 (N_12254,N_5051,N_62);
or U12255 (N_12255,N_3718,N_5806);
nor U12256 (N_12256,N_2664,N_2851);
or U12257 (N_12257,N_424,N_4401);
xor U12258 (N_12258,N_5530,N_6062);
or U12259 (N_12259,N_1733,N_1608);
nor U12260 (N_12260,N_6121,N_4138);
xnor U12261 (N_12261,N_1589,N_5158);
or U12262 (N_12262,N_2981,N_2364);
xor U12263 (N_12263,N_4591,N_4081);
or U12264 (N_12264,N_1414,N_880);
and U12265 (N_12265,N_934,N_3250);
nand U12266 (N_12266,N_5966,N_730);
or U12267 (N_12267,N_5981,N_5516);
nor U12268 (N_12268,N_3552,N_3028);
and U12269 (N_12269,N_4050,N_3479);
and U12270 (N_12270,N_849,N_5152);
nand U12271 (N_12271,N_1783,N_2924);
or U12272 (N_12272,N_2962,N_5110);
or U12273 (N_12273,N_5461,N_2395);
or U12274 (N_12274,N_4385,N_426);
and U12275 (N_12275,N_4306,N_2286);
or U12276 (N_12276,N_4226,N_703);
nand U12277 (N_12277,N_2411,N_6217);
nand U12278 (N_12278,N_5145,N_3099);
and U12279 (N_12279,N_1661,N_6113);
and U12280 (N_12280,N_4409,N_513);
xnor U12281 (N_12281,N_5790,N_661);
xnor U12282 (N_12282,N_4822,N_4874);
and U12283 (N_12283,N_4794,N_1037);
nor U12284 (N_12284,N_3241,N_1387);
and U12285 (N_12285,N_3694,N_2231);
or U12286 (N_12286,N_3768,N_1222);
xor U12287 (N_12287,N_1100,N_3222);
nand U12288 (N_12288,N_2103,N_5333);
xnor U12289 (N_12289,N_4138,N_4622);
or U12290 (N_12290,N_3523,N_1937);
and U12291 (N_12291,N_4335,N_5347);
xor U12292 (N_12292,N_4729,N_5940);
xor U12293 (N_12293,N_477,N_1619);
nor U12294 (N_12294,N_4276,N_4790);
nor U12295 (N_12295,N_2821,N_5157);
and U12296 (N_12296,N_1857,N_1786);
nand U12297 (N_12297,N_6204,N_2935);
nand U12298 (N_12298,N_2992,N_875);
xor U12299 (N_12299,N_1808,N_4867);
and U12300 (N_12300,N_5224,N_4085);
and U12301 (N_12301,N_2837,N_2069);
nor U12302 (N_12302,N_1219,N_5835);
nor U12303 (N_12303,N_4143,N_2254);
nor U12304 (N_12304,N_241,N_2298);
and U12305 (N_12305,N_813,N_5446);
or U12306 (N_12306,N_175,N_4097);
nand U12307 (N_12307,N_3640,N_109);
xnor U12308 (N_12308,N_6237,N_1690);
or U12309 (N_12309,N_594,N_4188);
and U12310 (N_12310,N_1027,N_3684);
and U12311 (N_12311,N_5889,N_5542);
or U12312 (N_12312,N_3070,N_3296);
nand U12313 (N_12313,N_1783,N_2437);
or U12314 (N_12314,N_519,N_5198);
nand U12315 (N_12315,N_1416,N_216);
nand U12316 (N_12316,N_1899,N_5872);
nor U12317 (N_12317,N_4521,N_6145);
nor U12318 (N_12318,N_2957,N_3754);
and U12319 (N_12319,N_2887,N_3381);
xnor U12320 (N_12320,N_2605,N_134);
nor U12321 (N_12321,N_6213,N_6111);
nand U12322 (N_12322,N_5134,N_4118);
and U12323 (N_12323,N_1592,N_4418);
or U12324 (N_12324,N_6041,N_3864);
nor U12325 (N_12325,N_5759,N_1160);
xor U12326 (N_12326,N_2298,N_2518);
nand U12327 (N_12327,N_458,N_1230);
or U12328 (N_12328,N_5004,N_2741);
and U12329 (N_12329,N_6214,N_2409);
xor U12330 (N_12330,N_1515,N_3989);
xnor U12331 (N_12331,N_1992,N_6020);
xor U12332 (N_12332,N_2406,N_4355);
nand U12333 (N_12333,N_5629,N_604);
or U12334 (N_12334,N_2651,N_711);
nor U12335 (N_12335,N_2778,N_5360);
and U12336 (N_12336,N_6060,N_4371);
and U12337 (N_12337,N_2581,N_895);
nand U12338 (N_12338,N_5842,N_2606);
xnor U12339 (N_12339,N_2516,N_6112);
nor U12340 (N_12340,N_1883,N_4219);
nand U12341 (N_12341,N_4859,N_4188);
or U12342 (N_12342,N_4859,N_3466);
and U12343 (N_12343,N_5428,N_2964);
nand U12344 (N_12344,N_1089,N_2184);
and U12345 (N_12345,N_5337,N_5050);
xor U12346 (N_12346,N_5953,N_4147);
nand U12347 (N_12347,N_2680,N_3402);
xor U12348 (N_12348,N_6073,N_5744);
nor U12349 (N_12349,N_2691,N_5917);
nand U12350 (N_12350,N_1350,N_4051);
xnor U12351 (N_12351,N_4287,N_3208);
or U12352 (N_12352,N_2682,N_2436);
and U12353 (N_12353,N_4492,N_792);
xnor U12354 (N_12354,N_6194,N_5963);
xor U12355 (N_12355,N_74,N_5423);
or U12356 (N_12356,N_309,N_5127);
or U12357 (N_12357,N_4157,N_6230);
nor U12358 (N_12358,N_4501,N_1758);
nor U12359 (N_12359,N_4597,N_5361);
nor U12360 (N_12360,N_2901,N_5864);
xnor U12361 (N_12361,N_183,N_2019);
nand U12362 (N_12362,N_5809,N_4245);
nand U12363 (N_12363,N_3942,N_1448);
nand U12364 (N_12364,N_1122,N_2766);
nor U12365 (N_12365,N_31,N_1891);
or U12366 (N_12366,N_5164,N_260);
xor U12367 (N_12367,N_6144,N_679);
nor U12368 (N_12368,N_3127,N_2817);
xor U12369 (N_12369,N_2850,N_23);
nor U12370 (N_12370,N_473,N_6235);
or U12371 (N_12371,N_5678,N_5205);
nor U12372 (N_12372,N_6132,N_4228);
xnor U12373 (N_12373,N_829,N_4609);
nand U12374 (N_12374,N_6181,N_5800);
and U12375 (N_12375,N_3371,N_5803);
or U12376 (N_12376,N_4053,N_879);
xnor U12377 (N_12377,N_5793,N_3986);
or U12378 (N_12378,N_2609,N_4495);
xor U12379 (N_12379,N_2660,N_43);
nor U12380 (N_12380,N_2052,N_4853);
and U12381 (N_12381,N_3628,N_4450);
nand U12382 (N_12382,N_3811,N_3217);
and U12383 (N_12383,N_5199,N_4882);
xnor U12384 (N_12384,N_5228,N_3322);
and U12385 (N_12385,N_3798,N_680);
or U12386 (N_12386,N_3590,N_2765);
nor U12387 (N_12387,N_480,N_4376);
xnor U12388 (N_12388,N_4706,N_404);
nand U12389 (N_12389,N_1561,N_1884);
nand U12390 (N_12390,N_3737,N_748);
xor U12391 (N_12391,N_1529,N_242);
nor U12392 (N_12392,N_1013,N_4687);
nor U12393 (N_12393,N_3231,N_1014);
and U12394 (N_12394,N_3069,N_3267);
nand U12395 (N_12395,N_5691,N_2287);
xnor U12396 (N_12396,N_5710,N_6214);
or U12397 (N_12397,N_4941,N_1352);
nand U12398 (N_12398,N_4307,N_911);
nor U12399 (N_12399,N_6017,N_3428);
or U12400 (N_12400,N_1323,N_2359);
or U12401 (N_12401,N_3654,N_2270);
xnor U12402 (N_12402,N_2378,N_2508);
or U12403 (N_12403,N_5497,N_1517);
xor U12404 (N_12404,N_1821,N_317);
nor U12405 (N_12405,N_6061,N_3253);
or U12406 (N_12406,N_5405,N_3717);
or U12407 (N_12407,N_968,N_3065);
or U12408 (N_12408,N_4884,N_1393);
nor U12409 (N_12409,N_1151,N_4896);
nor U12410 (N_12410,N_2334,N_1880);
nand U12411 (N_12411,N_4315,N_2819);
nor U12412 (N_12412,N_668,N_441);
and U12413 (N_12413,N_2147,N_3121);
and U12414 (N_12414,N_5593,N_1007);
nand U12415 (N_12415,N_948,N_3467);
nor U12416 (N_12416,N_5801,N_1073);
and U12417 (N_12417,N_4987,N_3594);
or U12418 (N_12418,N_610,N_1995);
and U12419 (N_12419,N_5501,N_5570);
xor U12420 (N_12420,N_4942,N_481);
and U12421 (N_12421,N_4836,N_2493);
xnor U12422 (N_12422,N_3548,N_1926);
nor U12423 (N_12423,N_2445,N_485);
or U12424 (N_12424,N_2973,N_4710);
or U12425 (N_12425,N_3972,N_4654);
and U12426 (N_12426,N_1252,N_4820);
xor U12427 (N_12427,N_5074,N_1113);
nor U12428 (N_12428,N_1504,N_1635);
nor U12429 (N_12429,N_5896,N_4852);
or U12430 (N_12430,N_396,N_5619);
nand U12431 (N_12431,N_2565,N_1421);
nor U12432 (N_12432,N_1942,N_4138);
nand U12433 (N_12433,N_3768,N_1450);
and U12434 (N_12434,N_4002,N_823);
nand U12435 (N_12435,N_1930,N_987);
or U12436 (N_12436,N_1207,N_3374);
or U12437 (N_12437,N_5391,N_3952);
or U12438 (N_12438,N_564,N_971);
nand U12439 (N_12439,N_2698,N_5433);
or U12440 (N_12440,N_3689,N_891);
nand U12441 (N_12441,N_3819,N_3679);
nand U12442 (N_12442,N_2446,N_5140);
nor U12443 (N_12443,N_2850,N_1346);
or U12444 (N_12444,N_6186,N_808);
or U12445 (N_12445,N_5253,N_5339);
or U12446 (N_12446,N_1016,N_3257);
or U12447 (N_12447,N_3230,N_3324);
nor U12448 (N_12448,N_4284,N_1112);
nand U12449 (N_12449,N_2838,N_3414);
and U12450 (N_12450,N_3066,N_2898);
and U12451 (N_12451,N_3781,N_2975);
or U12452 (N_12452,N_368,N_4971);
nand U12453 (N_12453,N_4266,N_1555);
or U12454 (N_12454,N_5825,N_1668);
nor U12455 (N_12455,N_1330,N_3958);
xnor U12456 (N_12456,N_2326,N_5809);
or U12457 (N_12457,N_3944,N_1177);
and U12458 (N_12458,N_4291,N_775);
nor U12459 (N_12459,N_2134,N_1528);
nand U12460 (N_12460,N_5341,N_2986);
nor U12461 (N_12461,N_5117,N_2702);
xnor U12462 (N_12462,N_4207,N_6123);
nor U12463 (N_12463,N_327,N_5374);
nand U12464 (N_12464,N_3534,N_1407);
nand U12465 (N_12465,N_3665,N_1267);
xnor U12466 (N_12466,N_4903,N_2823);
nor U12467 (N_12467,N_4843,N_172);
nand U12468 (N_12468,N_4942,N_1303);
nor U12469 (N_12469,N_3829,N_5151);
nand U12470 (N_12470,N_4494,N_2946);
nand U12471 (N_12471,N_133,N_512);
nor U12472 (N_12472,N_848,N_961);
nor U12473 (N_12473,N_2131,N_5574);
xnor U12474 (N_12474,N_3514,N_3406);
xor U12475 (N_12475,N_4915,N_1928);
or U12476 (N_12476,N_3418,N_4168);
and U12477 (N_12477,N_2140,N_2088);
nor U12478 (N_12478,N_5779,N_5266);
nand U12479 (N_12479,N_1270,N_2875);
nand U12480 (N_12480,N_6014,N_3787);
and U12481 (N_12481,N_342,N_4706);
nand U12482 (N_12482,N_1052,N_778);
nor U12483 (N_12483,N_3843,N_4640);
xor U12484 (N_12484,N_404,N_603);
xnor U12485 (N_12485,N_4821,N_2952);
and U12486 (N_12486,N_4493,N_4189);
or U12487 (N_12487,N_3625,N_77);
or U12488 (N_12488,N_4970,N_1301);
and U12489 (N_12489,N_1961,N_5650);
or U12490 (N_12490,N_2861,N_5177);
nand U12491 (N_12491,N_4852,N_1076);
xor U12492 (N_12492,N_2646,N_110);
xor U12493 (N_12493,N_5701,N_573);
xnor U12494 (N_12494,N_3289,N_5238);
or U12495 (N_12495,N_14,N_514);
and U12496 (N_12496,N_2146,N_3664);
xnor U12497 (N_12497,N_1210,N_4308);
nand U12498 (N_12498,N_2812,N_2667);
nand U12499 (N_12499,N_5746,N_1305);
xnor U12500 (N_12500,N_6797,N_12266);
nand U12501 (N_12501,N_9340,N_6668);
or U12502 (N_12502,N_11534,N_10735);
nor U12503 (N_12503,N_10015,N_10853);
and U12504 (N_12504,N_7074,N_6834);
nand U12505 (N_12505,N_7711,N_9974);
and U12506 (N_12506,N_11135,N_10510);
and U12507 (N_12507,N_7991,N_9207);
nand U12508 (N_12508,N_6357,N_10725);
and U12509 (N_12509,N_7143,N_7402);
nand U12510 (N_12510,N_7150,N_12179);
nand U12511 (N_12511,N_12484,N_12254);
nor U12512 (N_12512,N_9664,N_12250);
and U12513 (N_12513,N_6833,N_6636);
xor U12514 (N_12514,N_11013,N_8166);
or U12515 (N_12515,N_7736,N_10347);
and U12516 (N_12516,N_9169,N_11225);
xnor U12517 (N_12517,N_11442,N_11128);
and U12518 (N_12518,N_8077,N_10927);
nand U12519 (N_12519,N_11792,N_8573);
or U12520 (N_12520,N_11168,N_9021);
or U12521 (N_12521,N_10301,N_9161);
nor U12522 (N_12522,N_9280,N_9709);
nor U12523 (N_12523,N_11720,N_11704);
or U12524 (N_12524,N_11217,N_12190);
nor U12525 (N_12525,N_12495,N_10990);
nor U12526 (N_12526,N_7213,N_11468);
nor U12527 (N_12527,N_9850,N_10863);
and U12528 (N_12528,N_11830,N_6708);
xnor U12529 (N_12529,N_10078,N_8822);
and U12530 (N_12530,N_9486,N_11173);
xnor U12531 (N_12531,N_11444,N_8564);
or U12532 (N_12532,N_11141,N_8603);
nand U12533 (N_12533,N_8454,N_8031);
and U12534 (N_12534,N_8843,N_11210);
nand U12535 (N_12535,N_6404,N_6896);
or U12536 (N_12536,N_6395,N_9581);
and U12537 (N_12537,N_12413,N_10213);
nand U12538 (N_12538,N_11417,N_8037);
nand U12539 (N_12539,N_6702,N_9611);
and U12540 (N_12540,N_11240,N_12186);
nor U12541 (N_12541,N_9313,N_10586);
or U12542 (N_12542,N_9227,N_11449);
nand U12543 (N_12543,N_10470,N_8882);
nor U12544 (N_12544,N_10421,N_8247);
and U12545 (N_12545,N_6898,N_6371);
and U12546 (N_12546,N_9725,N_10490);
nor U12547 (N_12547,N_8890,N_11418);
xor U12548 (N_12548,N_6270,N_10223);
and U12549 (N_12549,N_7082,N_12074);
xor U12550 (N_12550,N_10198,N_7425);
and U12551 (N_12551,N_11668,N_9790);
nand U12552 (N_12552,N_8589,N_9091);
xor U12553 (N_12553,N_8266,N_9258);
nor U12554 (N_12554,N_11954,N_12176);
nor U12555 (N_12555,N_12294,N_9605);
or U12556 (N_12556,N_7359,N_12381);
xor U12557 (N_12557,N_8296,N_10189);
xnor U12558 (N_12558,N_9650,N_8088);
nand U12559 (N_12559,N_12349,N_6997);
or U12560 (N_12560,N_12209,N_10958);
xor U12561 (N_12561,N_8445,N_11184);
xor U12562 (N_12562,N_10133,N_10203);
or U12563 (N_12563,N_12088,N_10807);
or U12564 (N_12564,N_11707,N_10914);
xor U12565 (N_12565,N_7782,N_11764);
nand U12566 (N_12566,N_9440,N_11018);
nor U12567 (N_12567,N_8932,N_6418);
xnor U12568 (N_12568,N_6544,N_9439);
xnor U12569 (N_12569,N_8778,N_9515);
nand U12570 (N_12570,N_10062,N_8139);
and U12571 (N_12571,N_8257,N_11475);
nor U12572 (N_12572,N_7266,N_9622);
xor U12573 (N_12573,N_11885,N_9388);
xor U12574 (N_12574,N_10453,N_7668);
xor U12575 (N_12575,N_11189,N_8938);
nand U12576 (N_12576,N_11835,N_8268);
or U12577 (N_12577,N_11087,N_10911);
nand U12578 (N_12578,N_6654,N_10605);
nor U12579 (N_12579,N_11608,N_6366);
nand U12580 (N_12580,N_10960,N_8873);
nor U12581 (N_12581,N_11714,N_7181);
or U12582 (N_12582,N_6323,N_10538);
xnor U12583 (N_12583,N_7217,N_12280);
or U12584 (N_12584,N_11179,N_12299);
and U12585 (N_12585,N_11022,N_9076);
or U12586 (N_12586,N_6575,N_11043);
nor U12587 (N_12587,N_10776,N_7506);
or U12588 (N_12588,N_10265,N_11749);
xor U12589 (N_12589,N_12168,N_8020);
or U12590 (N_12590,N_8983,N_10098);
nand U12591 (N_12591,N_10868,N_6559);
nor U12592 (N_12592,N_10022,N_11049);
and U12593 (N_12593,N_12105,N_9818);
nand U12594 (N_12594,N_10786,N_11302);
nor U12595 (N_12595,N_9051,N_7903);
nand U12596 (N_12596,N_9792,N_8342);
nand U12597 (N_12597,N_9306,N_8903);
xor U12598 (N_12598,N_11702,N_8340);
nor U12599 (N_12599,N_10076,N_9585);
and U12600 (N_12600,N_8710,N_9367);
xnor U12601 (N_12601,N_7588,N_7803);
nor U12602 (N_12602,N_11530,N_8200);
nor U12603 (N_12603,N_10152,N_6503);
xnor U12604 (N_12604,N_11322,N_7199);
or U12605 (N_12605,N_8465,N_8863);
xnor U12606 (N_12606,N_11224,N_6713);
nand U12607 (N_12607,N_7378,N_8324);
nor U12608 (N_12608,N_8473,N_12406);
nand U12609 (N_12609,N_8093,N_11577);
nor U12610 (N_12610,N_8336,N_10548);
nand U12611 (N_12611,N_7839,N_6510);
xor U12612 (N_12612,N_9404,N_11933);
or U12613 (N_12613,N_11039,N_9008);
nor U12614 (N_12614,N_10057,N_8131);
nand U12615 (N_12615,N_6916,N_9814);
nor U12616 (N_12616,N_6359,N_8785);
xnor U12617 (N_12617,N_9208,N_8495);
and U12618 (N_12618,N_8854,N_7988);
and U12619 (N_12619,N_6677,N_9748);
nand U12620 (N_12620,N_6354,N_8199);
and U12621 (N_12621,N_10650,N_7067);
xor U12622 (N_12622,N_11843,N_7428);
or U12623 (N_12623,N_8004,N_9590);
xor U12624 (N_12624,N_12323,N_6878);
nand U12625 (N_12625,N_7384,N_7544);
xnor U12626 (N_12626,N_8711,N_6365);
and U12627 (N_12627,N_7034,N_10254);
and U12628 (N_12628,N_11185,N_9211);
nand U12629 (N_12629,N_8745,N_8192);
or U12630 (N_12630,N_10436,N_11560);
nand U12631 (N_12631,N_10321,N_10410);
or U12632 (N_12632,N_8563,N_6574);
or U12633 (N_12633,N_11641,N_9411);
nand U12634 (N_12634,N_7805,N_8323);
xor U12635 (N_12635,N_9341,N_8069);
xor U12636 (N_12636,N_8285,N_9631);
nor U12637 (N_12637,N_11640,N_10405);
nand U12638 (N_12638,N_10329,N_11724);
xor U12639 (N_12639,N_12379,N_7685);
nand U12640 (N_12640,N_9506,N_6719);
xor U12641 (N_12641,N_9846,N_10626);
nand U12642 (N_12642,N_7447,N_8698);
xnor U12643 (N_12643,N_8365,N_8759);
xor U12644 (N_12644,N_8018,N_6267);
or U12645 (N_12645,N_8218,N_12213);
nand U12646 (N_12646,N_10357,N_9653);
nand U12647 (N_12647,N_6488,N_7243);
or U12648 (N_12648,N_7460,N_8942);
nor U12649 (N_12649,N_8674,N_7438);
or U12650 (N_12650,N_8439,N_6567);
xor U12651 (N_12651,N_7886,N_11464);
or U12652 (N_12652,N_11545,N_9349);
or U12653 (N_12653,N_10147,N_12479);
or U12654 (N_12654,N_6942,N_9312);
nor U12655 (N_12655,N_7442,N_8726);
and U12656 (N_12656,N_8065,N_11425);
or U12657 (N_12657,N_9285,N_6547);
nor U12658 (N_12658,N_12214,N_7969);
nor U12659 (N_12659,N_6373,N_7024);
xnor U12660 (N_12660,N_9327,N_7472);
nand U12661 (N_12661,N_10514,N_7806);
nand U12662 (N_12662,N_11887,N_12155);
and U12663 (N_12663,N_10408,N_12210);
xnor U12664 (N_12664,N_11732,N_9261);
nor U12665 (N_12665,N_9243,N_6954);
and U12666 (N_12666,N_7222,N_6434);
nor U12667 (N_12667,N_8629,N_7424);
nor U12668 (N_12668,N_9444,N_8697);
or U12669 (N_12669,N_11871,N_12346);
or U12670 (N_12670,N_12255,N_11664);
nand U12671 (N_12671,N_11784,N_11351);
xnor U12672 (N_12672,N_7382,N_11307);
or U12673 (N_12673,N_12410,N_8703);
or U12674 (N_12674,N_10156,N_10957);
and U12675 (N_12675,N_9045,N_9830);
and U12676 (N_12676,N_8043,N_7648);
and U12677 (N_12677,N_8352,N_9625);
nand U12678 (N_12678,N_9635,N_7502);
nand U12679 (N_12679,N_9975,N_6608);
and U12680 (N_12680,N_10272,N_7151);
nand U12681 (N_12681,N_10689,N_11708);
or U12682 (N_12682,N_9598,N_6429);
nand U12683 (N_12683,N_8681,N_9481);
or U12684 (N_12684,N_8633,N_6659);
nor U12685 (N_12685,N_7889,N_8859);
or U12686 (N_12686,N_6733,N_9568);
nand U12687 (N_12687,N_12496,N_6825);
nand U12688 (N_12688,N_9134,N_7778);
nand U12689 (N_12689,N_7927,N_7929);
nor U12690 (N_12690,N_9869,N_11804);
nor U12691 (N_12691,N_8164,N_9263);
or U12692 (N_12692,N_10093,N_11350);
or U12693 (N_12693,N_7342,N_8271);
xor U12694 (N_12694,N_11609,N_10847);
nand U12695 (N_12695,N_11359,N_9401);
or U12696 (N_12696,N_6947,N_11544);
xnor U12697 (N_12697,N_10296,N_11884);
nor U12698 (N_12698,N_12145,N_11424);
or U12699 (N_12699,N_6963,N_11414);
nor U12700 (N_12700,N_8419,N_9746);
or U12701 (N_12701,N_6331,N_7632);
and U12702 (N_12702,N_9474,N_11689);
nor U12703 (N_12703,N_6690,N_11421);
xor U12704 (N_12704,N_8202,N_7374);
xor U12705 (N_12705,N_6975,N_7968);
nor U12706 (N_12706,N_12051,N_9954);
and U12707 (N_12707,N_10867,N_9656);
nand U12708 (N_12708,N_8382,N_8949);
or U12709 (N_12709,N_9373,N_11542);
or U12710 (N_12710,N_10407,N_8328);
or U12711 (N_12711,N_11983,N_10909);
and U12712 (N_12712,N_8229,N_12384);
xnor U12713 (N_12713,N_11139,N_9289);
or U12714 (N_12714,N_7494,N_9291);
nand U12715 (N_12715,N_10117,N_10440);
and U12716 (N_12716,N_10602,N_12199);
nand U12717 (N_12717,N_8689,N_10392);
xnor U12718 (N_12718,N_10527,N_12258);
nand U12719 (N_12719,N_8637,N_9383);
or U12720 (N_12720,N_6277,N_10517);
and U12721 (N_12721,N_8567,N_10525);
nor U12722 (N_12722,N_11723,N_11762);
nand U12723 (N_12723,N_6743,N_8104);
and U12724 (N_12724,N_9087,N_7844);
nand U12725 (N_12725,N_8203,N_10435);
nor U12726 (N_12726,N_7670,N_7023);
and U12727 (N_12727,N_10509,N_7339);
and U12728 (N_12728,N_7423,N_8046);
or U12729 (N_12729,N_9777,N_7992);
xor U12730 (N_12730,N_10688,N_8855);
or U12731 (N_12731,N_7452,N_8406);
and U12732 (N_12732,N_8420,N_10524);
nand U12733 (N_12733,N_8702,N_8925);
nor U12734 (N_12734,N_10830,N_11977);
xor U12735 (N_12735,N_8278,N_8511);
or U12736 (N_12736,N_11950,N_7247);
xor U12737 (N_12737,N_9923,N_9187);
or U12738 (N_12738,N_9623,N_7086);
nand U12739 (N_12739,N_12437,N_8213);
nor U12740 (N_12740,N_10639,N_6647);
xor U12741 (N_12741,N_12197,N_6800);
nor U12742 (N_12742,N_11842,N_12350);
xnor U12743 (N_12743,N_9062,N_6319);
xor U12744 (N_12744,N_6250,N_7906);
nor U12745 (N_12745,N_8103,N_7441);
and U12746 (N_12746,N_8971,N_8728);
nand U12747 (N_12747,N_12004,N_12243);
and U12748 (N_12748,N_12154,N_9819);
nor U12749 (N_12749,N_8430,N_12124);
nand U12750 (N_12750,N_12412,N_8198);
or U12751 (N_12751,N_11131,N_11344);
xor U12752 (N_12752,N_10401,N_10917);
nor U12753 (N_12753,N_11581,N_11208);
or U12754 (N_12754,N_7864,N_11891);
nand U12755 (N_12755,N_6338,N_7935);
or U12756 (N_12756,N_10445,N_10291);
nand U12757 (N_12757,N_9673,N_7451);
or U12758 (N_12758,N_9249,N_8753);
nor U12759 (N_12759,N_7930,N_12314);
nand U12760 (N_12760,N_9115,N_10027);
nor U12761 (N_12761,N_11023,N_8006);
nand U12762 (N_12762,N_12083,N_9994);
nor U12763 (N_12763,N_11747,N_9736);
or U12764 (N_12764,N_8927,N_11484);
xnor U12765 (N_12765,N_6731,N_7265);
nand U12766 (N_12766,N_10233,N_10131);
nor U12767 (N_12767,N_10207,N_8919);
and U12768 (N_12768,N_9145,N_11953);
xnor U12769 (N_12769,N_10590,N_10141);
nand U12770 (N_12770,N_7307,N_9095);
nor U12771 (N_12771,N_7413,N_8312);
xor U12772 (N_12772,N_10817,N_10986);
nand U12773 (N_12773,N_11080,N_12364);
or U12774 (N_12774,N_12371,N_11527);
and U12775 (N_12775,N_11625,N_9668);
or U12776 (N_12776,N_10297,N_11451);
nand U12777 (N_12777,N_7667,N_9562);
or U12778 (N_12778,N_7841,N_8708);
xor U12779 (N_12779,N_10876,N_9414);
and U12780 (N_12780,N_6516,N_9260);
xor U12781 (N_12781,N_7884,N_9437);
and U12782 (N_12782,N_11693,N_7394);
nand U12783 (N_12783,N_9752,N_6257);
nor U12784 (N_12784,N_7322,N_9442);
xnor U12785 (N_12785,N_9152,N_6817);
nand U12786 (N_12786,N_8254,N_12191);
nor U12787 (N_12787,N_11275,N_7691);
and U12788 (N_12788,N_6540,N_11183);
nor U12789 (N_12789,N_7784,N_10221);
nand U12790 (N_12790,N_7986,N_6394);
or U12791 (N_12791,N_11261,N_7408);
xnor U12792 (N_12792,N_6579,N_9302);
nor U12793 (N_12793,N_7120,N_11236);
nor U12794 (N_12794,N_8349,N_11161);
or U12795 (N_12795,N_6557,N_10919);
nand U12796 (N_12796,N_10243,N_9505);
and U12797 (N_12797,N_6915,N_10733);
xnor U12798 (N_12798,N_8738,N_10275);
xor U12799 (N_12799,N_8764,N_10034);
xnor U12800 (N_12800,N_9155,N_9485);
nand U12801 (N_12801,N_10926,N_11011);
and U12802 (N_12802,N_8668,N_10678);
nand U12803 (N_12803,N_10754,N_8294);
or U12804 (N_12804,N_9049,N_11800);
and U12805 (N_12805,N_8542,N_9894);
and U12806 (N_12806,N_8048,N_10481);
xor U12807 (N_12807,N_9405,N_6470);
or U12808 (N_12808,N_9473,N_11398);
and U12809 (N_12809,N_10163,N_10944);
and U12810 (N_12810,N_9047,N_9331);
xor U12811 (N_12811,N_7657,N_10751);
and U12812 (N_12812,N_10516,N_8013);
or U12813 (N_12813,N_7586,N_7688);
and U12814 (N_12814,N_11684,N_9369);
and U12815 (N_12815,N_12400,N_7054);
nor U12816 (N_12816,N_8087,N_9362);
nor U12817 (N_12817,N_6391,N_9947);
nand U12818 (N_12818,N_8232,N_10448);
nand U12819 (N_12819,N_12234,N_10671);
nor U12820 (N_12820,N_8049,N_9137);
and U12821 (N_12821,N_6598,N_8106);
nor U12822 (N_12822,N_8251,N_11604);
nor U12823 (N_12823,N_11061,N_11150);
xor U12824 (N_12824,N_11405,N_11159);
and U12825 (N_12825,N_12049,N_10838);
or U12826 (N_12826,N_11134,N_10928);
nor U12827 (N_12827,N_12293,N_11892);
xor U12828 (N_12828,N_10942,N_11375);
nand U12829 (N_12829,N_7654,N_10779);
xor U12830 (N_12830,N_11448,N_11976);
and U12831 (N_12831,N_7798,N_11157);
xnor U12832 (N_12832,N_10464,N_11591);
and U12833 (N_12833,N_8146,N_6742);
xor U12834 (N_12834,N_9205,N_8116);
and U12835 (N_12835,N_9825,N_9416);
nor U12836 (N_12836,N_9520,N_8391);
or U12837 (N_12837,N_6988,N_6845);
or U12838 (N_12838,N_10149,N_8731);
nor U12839 (N_12839,N_7952,N_9379);
and U12840 (N_12840,N_11868,N_9560);
xnor U12841 (N_12841,N_11403,N_10961);
nor U12842 (N_12842,N_7231,N_12080);
nor U12843 (N_12843,N_11774,N_6284);
or U12844 (N_12844,N_11423,N_7118);
nor U12845 (N_12845,N_10587,N_8153);
or U12846 (N_12846,N_10573,N_6973);
xnor U12847 (N_12847,N_6486,N_9057);
and U12848 (N_12848,N_10628,N_10334);
and U12849 (N_12849,N_6259,N_11223);
nor U12850 (N_12850,N_6970,N_7198);
nor U12851 (N_12851,N_8063,N_7899);
nor U12852 (N_12852,N_7341,N_9834);
and U12853 (N_12853,N_11777,N_8516);
xor U12854 (N_12854,N_6414,N_9633);
or U12855 (N_12855,N_7715,N_8579);
xnor U12856 (N_12856,N_7720,N_7562);
nor U12857 (N_12857,N_11955,N_11199);
xnor U12858 (N_12858,N_10319,N_7958);
nand U12859 (N_12859,N_8421,N_10624);
xnor U12860 (N_12860,N_12386,N_12283);
xor U12861 (N_12861,N_8304,N_9604);
nand U12862 (N_12862,N_8231,N_9122);
xor U12863 (N_12863,N_10571,N_7095);
xnor U12864 (N_12864,N_8970,N_11276);
nand U12865 (N_12865,N_10806,N_9538);
xnor U12866 (N_12866,N_11929,N_6587);
nand U12867 (N_12867,N_11323,N_8791);
and U12868 (N_12868,N_7960,N_8246);
nor U12869 (N_12869,N_7953,N_6506);
or U12870 (N_12870,N_9268,N_8794);
nand U12871 (N_12871,N_8144,N_9649);
xor U12872 (N_12872,N_10783,N_12095);
or U12873 (N_12873,N_6465,N_10480);
xnor U12874 (N_12874,N_8094,N_9529);
or U12875 (N_12875,N_8551,N_6716);
nor U12876 (N_12876,N_6995,N_12041);
xor U12877 (N_12877,N_8409,N_11400);
xnor U12878 (N_12878,N_10528,N_12081);
or U12879 (N_12879,N_6646,N_10603);
nor U12880 (N_12880,N_11343,N_9204);
or U12881 (N_12881,N_11593,N_8606);
xor U12882 (N_12882,N_10711,N_11738);
nor U12883 (N_12883,N_12481,N_8112);
and U12884 (N_12884,N_11863,N_9901);
nand U12885 (N_12885,N_6867,N_11197);
xor U12886 (N_12886,N_8662,N_10075);
nor U12887 (N_12887,N_10187,N_9662);
and U12888 (N_12888,N_9575,N_8168);
nand U12889 (N_12889,N_7616,N_10483);
nand U12890 (N_12890,N_7827,N_12402);
and U12891 (N_12891,N_11748,N_6645);
or U12892 (N_12892,N_11721,N_9813);
nor U12893 (N_12893,N_12423,N_10774);
or U12894 (N_12894,N_8652,N_9443);
xor U12895 (N_12895,N_11558,N_7980);
or U12896 (N_12896,N_6344,N_7318);
and U12897 (N_12897,N_11687,N_7268);
nand U12898 (N_12898,N_8646,N_8626);
xnor U12899 (N_12899,N_10870,N_10413);
or U12900 (N_12900,N_7192,N_8317);
xor U12901 (N_12901,N_6489,N_8835);
nand U12902 (N_12902,N_10307,N_7730);
and U12903 (N_12903,N_8379,N_11396);
or U12904 (N_12904,N_7161,N_12007);
nor U12905 (N_12905,N_10941,N_11540);
nor U12906 (N_12906,N_10353,N_10292);
xor U12907 (N_12907,N_7454,N_8634);
and U12908 (N_12908,N_8081,N_8082);
nand U12909 (N_12909,N_8747,N_11531);
and U12910 (N_12910,N_8776,N_6548);
nand U12911 (N_12911,N_10971,N_10261);
nand U12912 (N_12912,N_11921,N_11420);
or U12913 (N_12913,N_6798,N_8872);
and U12914 (N_12914,N_8366,N_8201);
and U12915 (N_12915,N_10600,N_6499);
xnor U12916 (N_12916,N_10106,N_9909);
nand U12917 (N_12917,N_11840,N_12089);
xnor U12918 (N_12918,N_7195,N_6508);
nor U12919 (N_12919,N_8401,N_10616);
or U12920 (N_12920,N_6826,N_6409);
nand U12921 (N_12921,N_7241,N_10797);
and U12922 (N_12922,N_6529,N_6669);
xor U12923 (N_12923,N_9472,N_6333);
xor U12924 (N_12924,N_8783,N_9743);
nor U12925 (N_12925,N_6885,N_11971);
and U12926 (N_12926,N_11551,N_6736);
xnor U12927 (N_12927,N_6334,N_11074);
and U12928 (N_12928,N_11710,N_11112);
nand U12929 (N_12929,N_7395,N_7155);
or U12930 (N_12930,N_6408,N_10750);
nor U12931 (N_12931,N_8376,N_9262);
nor U12932 (N_12932,N_8513,N_11858);
or U12933 (N_12933,N_12042,N_7761);
and U12934 (N_12934,N_9824,N_11127);
and U12935 (N_12935,N_11637,N_9963);
and U12936 (N_12936,N_11172,N_9763);
or U12937 (N_12937,N_10818,N_8057);
nor U12938 (N_12938,N_10286,N_8865);
nand U12939 (N_12939,N_9429,N_10002);
and U12940 (N_12940,N_10976,N_9328);
nor U12941 (N_12941,N_12491,N_9804);
nand U12942 (N_12942,N_11142,N_6657);
or U12943 (N_12943,N_10798,N_9671);
and U12944 (N_12944,N_9352,N_11780);
or U12945 (N_12945,N_6724,N_8457);
nand U12946 (N_12946,N_10757,N_8779);
xnor U12947 (N_12947,N_10881,N_11911);
and U12948 (N_12948,N_11057,N_7001);
or U12949 (N_12949,N_7252,N_8559);
or U12950 (N_12950,N_7430,N_10036);
xnor U12951 (N_12951,N_8905,N_7661);
and U12952 (N_12952,N_7727,N_11501);
xnor U12953 (N_12953,N_11395,N_7933);
nor U12954 (N_12954,N_6445,N_7713);
and U12955 (N_12955,N_10135,N_7234);
and U12956 (N_12956,N_7587,N_9501);
nor U12957 (N_12957,N_11355,N_11821);
nor U12958 (N_12958,N_11368,N_9252);
and U12959 (N_12959,N_7115,N_9663);
xor U12960 (N_12960,N_7399,N_9791);
or U12961 (N_12961,N_12478,N_10165);
nand U12962 (N_12962,N_9168,N_12061);
xnor U12963 (N_12963,N_11460,N_9292);
nand U12964 (N_12964,N_11736,N_8607);
and U12965 (N_12965,N_6820,N_11988);
xnor U12966 (N_12966,N_10840,N_9167);
and U12967 (N_12967,N_11873,N_6770);
nand U12968 (N_12968,N_7053,N_9800);
or U12969 (N_12969,N_7066,N_8984);
and U12970 (N_12970,N_8456,N_9866);
xnor U12971 (N_12971,N_6431,N_10235);
or U12972 (N_12972,N_6895,N_6869);
nand U12973 (N_12973,N_11329,N_12445);
nand U12974 (N_12974,N_12029,N_12008);
or U12975 (N_12975,N_10855,N_12269);
nand U12976 (N_12976,N_10655,N_9097);
xor U12977 (N_12977,N_7182,N_8138);
and U12978 (N_12978,N_9288,N_12417);
or U12979 (N_12979,N_9461,N_6872);
nand U12980 (N_12980,N_10253,N_6313);
nor U12981 (N_12981,N_9096,N_11825);
nor U12982 (N_12982,N_8749,N_6693);
nor U12983 (N_12983,N_11627,N_8152);
nor U12984 (N_12984,N_8499,N_8907);
and U12985 (N_12985,N_8986,N_7117);
xnor U12986 (N_12986,N_7434,N_8191);
and U12987 (N_12987,N_8469,N_10895);
nor U12988 (N_12988,N_12367,N_10745);
nand U12989 (N_12989,N_8884,N_9696);
xor U12990 (N_12990,N_10420,N_8870);
nand U12991 (N_12991,N_8472,N_7219);
xor U12992 (N_12992,N_10816,N_9674);
or U12993 (N_12993,N_9679,N_6282);
or U12994 (N_12994,N_10859,N_11700);
and U12995 (N_12995,N_8461,N_7305);
xnor U12996 (N_12996,N_9274,N_11441);
nand U12997 (N_12997,N_7824,N_11568);
or U12998 (N_12998,N_11940,N_8347);
or U12999 (N_12999,N_7205,N_7361);
or U13000 (N_13000,N_8255,N_7724);
and U13001 (N_13001,N_6629,N_10844);
or U13002 (N_13002,N_11052,N_10260);
and U13003 (N_13003,N_8475,N_9140);
or U13004 (N_13004,N_10866,N_10282);
and U13005 (N_13005,N_11562,N_7700);
and U13006 (N_13006,N_9223,N_8714);
nor U13007 (N_13007,N_9835,N_11848);
nand U13008 (N_13008,N_11603,N_8692);
and U13009 (N_13009,N_8667,N_6278);
or U13010 (N_13010,N_9059,N_9949);
nand U13011 (N_13011,N_7156,N_12161);
or U13012 (N_13012,N_11045,N_10736);
and U13013 (N_13013,N_11430,N_12221);
and U13014 (N_13014,N_7317,N_8127);
and U13015 (N_13015,N_11260,N_9582);
nand U13016 (N_13016,N_6305,N_11681);
nor U13017 (N_13017,N_6822,N_9802);
or U13018 (N_13018,N_9574,N_6612);
nor U13019 (N_13019,N_6387,N_10641);
nor U13020 (N_13020,N_6462,N_10674);
nand U13021 (N_13021,N_11918,N_8679);
and U13022 (N_13022,N_9394,N_8619);
and U13023 (N_13023,N_10373,N_11075);
and U13024 (N_13024,N_7170,N_9082);
nand U13025 (N_13025,N_6907,N_8742);
nand U13026 (N_13026,N_11415,N_8771);
nor U13027 (N_13027,N_8375,N_6618);
and U13028 (N_13028,N_10263,N_8761);
xnor U13029 (N_13029,N_7592,N_8631);
nand U13030 (N_13030,N_11133,N_7403);
and U13031 (N_13031,N_11657,N_6712);
xnor U13032 (N_13032,N_10326,N_8937);
and U13033 (N_13033,N_6673,N_7649);
nor U13034 (N_13034,N_9110,N_10549);
and U13035 (N_13035,N_6564,N_6407);
xnor U13036 (N_13036,N_9170,N_10432);
and U13037 (N_13037,N_8586,N_9005);
and U13038 (N_13038,N_6309,N_11959);
or U13039 (N_13039,N_11097,N_7582);
xor U13040 (N_13040,N_7471,N_11214);
xnor U13041 (N_13041,N_6467,N_8616);
or U13042 (N_13042,N_9364,N_7790);
nand U13043 (N_13043,N_6982,N_6533);
and U13044 (N_13044,N_12375,N_8068);
nor U13045 (N_13045,N_7235,N_9221);
or U13046 (N_13046,N_9993,N_12188);
xor U13047 (N_13047,N_6591,N_11033);
xor U13048 (N_13048,N_7267,N_7100);
nor U13049 (N_13049,N_6265,N_9991);
xor U13050 (N_13050,N_10300,N_11229);
nand U13051 (N_13051,N_9877,N_12228);
or U13052 (N_13052,N_11931,N_9517);
xor U13053 (N_13053,N_12482,N_12211);
and U13054 (N_13054,N_6509,N_11869);
xnor U13055 (N_13055,N_8774,N_7414);
or U13056 (N_13056,N_8125,N_8211);
or U13057 (N_13057,N_9479,N_10284);
and U13058 (N_13058,N_9962,N_8120);
xnor U13059 (N_13059,N_12429,N_7308);
nor U13060 (N_13060,N_11026,N_12475);
xnor U13061 (N_13061,N_8723,N_12057);
xnor U13062 (N_13062,N_7041,N_7936);
or U13063 (N_13063,N_7660,N_6556);
or U13064 (N_13064,N_6477,N_6589);
or U13065 (N_13065,N_9875,N_7042);
and U13066 (N_13066,N_10028,N_11968);
nand U13067 (N_13067,N_8943,N_11740);
nor U13068 (N_13068,N_8122,N_9918);
nor U13069 (N_13069,N_7142,N_10534);
nand U13070 (N_13070,N_7578,N_9406);
xnor U13071 (N_13071,N_8351,N_10621);
or U13072 (N_13072,N_7343,N_9713);
or U13073 (N_13073,N_10544,N_7171);
nand U13074 (N_13074,N_8163,N_7084);
nand U13075 (N_13075,N_11099,N_12169);
nand U13076 (N_13076,N_12117,N_11510);
nor U13077 (N_13077,N_10108,N_6739);
nor U13078 (N_13078,N_9693,N_6390);
or U13079 (N_13079,N_11914,N_9295);
xnor U13080 (N_13080,N_8186,N_10072);
nor U13081 (N_13081,N_8130,N_10580);
nand U13082 (N_13082,N_6992,N_8842);
nand U13083 (N_13083,N_7716,N_11727);
nor U13084 (N_13084,N_11653,N_9214);
xor U13085 (N_13085,N_6772,N_11538);
nand U13086 (N_13086,N_7125,N_9024);
xnor U13087 (N_13087,N_8383,N_6914);
xnor U13088 (N_13088,N_12356,N_11882);
or U13089 (N_13089,N_11956,N_10891);
xor U13090 (N_13090,N_7098,N_11994);
xnor U13091 (N_13091,N_7951,N_10657);
or U13092 (N_13092,N_9242,N_11245);
xnor U13093 (N_13093,N_9248,N_11101);
nand U13094 (N_13094,N_7303,N_6550);
nand U13095 (N_13095,N_7534,N_8493);
or U13096 (N_13096,N_9768,N_12206);
and U13097 (N_13097,N_8160,N_7554);
nand U13098 (N_13098,N_10511,N_11638);
xnor U13099 (N_13099,N_11810,N_8248);
nand U13100 (N_13100,N_11237,N_11472);
nor U13101 (N_13101,N_12262,N_11345);
and U13102 (N_13102,N_11406,N_9175);
or U13103 (N_13103,N_6738,N_8170);
and U13104 (N_13104,N_6287,N_7271);
or U13105 (N_13105,N_7102,N_11447);
xnor U13106 (N_13106,N_11270,N_8844);
nor U13107 (N_13107,N_8346,N_11090);
or U13108 (N_13108,N_9028,N_8250);
nand U13109 (N_13109,N_12151,N_11650);
or U13110 (N_13110,N_11200,N_11187);
or U13111 (N_13111,N_10682,N_8496);
xor U13112 (N_13112,N_8719,N_9648);
nor U13113 (N_13113,N_12162,N_10998);
and U13114 (N_13114,N_8480,N_11408);
nor U13115 (N_13115,N_9283,N_9320);
xor U13116 (N_13116,N_9733,N_10893);
nor U13117 (N_13117,N_8074,N_12164);
or U13118 (N_13118,N_10618,N_6505);
nor U13119 (N_13119,N_9789,N_7484);
nand U13120 (N_13120,N_11985,N_11239);
and U13121 (N_13121,N_9985,N_7977);
nand U13122 (N_13122,N_9425,N_12227);
nand U13123 (N_13123,N_9457,N_6952);
and U13124 (N_13124,N_11487,N_7464);
or U13125 (N_13125,N_11317,N_11813);
xnor U13126 (N_13126,N_7981,N_12337);
nand U13127 (N_13127,N_7223,N_6380);
xor U13128 (N_13128,N_11969,N_8293);
nor U13129 (N_13129,N_7325,N_7916);
nor U13130 (N_13130,N_8284,N_7278);
or U13131 (N_13131,N_12342,N_9946);
xnor U13132 (N_13132,N_6352,N_12338);
nand U13133 (N_13133,N_10679,N_7911);
nor U13134 (N_13134,N_6403,N_8962);
xor U13135 (N_13135,N_6522,N_8002);
and U13136 (N_13136,N_7467,N_8236);
xnor U13137 (N_13137,N_12411,N_7897);
nor U13138 (N_13138,N_9900,N_6857);
xnor U13139 (N_13139,N_10719,N_7802);
nand U13140 (N_13140,N_9978,N_9956);
or U13141 (N_13141,N_8389,N_6964);
and U13142 (N_13142,N_6602,N_9321);
and U13143 (N_13143,N_8330,N_10788);
xnor U13144 (N_13144,N_9921,N_12407);
and U13145 (N_13145,N_11919,N_12014);
and U13146 (N_13146,N_8209,N_11817);
nand U13147 (N_13147,N_12278,N_10972);
or U13148 (N_13148,N_8810,N_7801);
or U13149 (N_13149,N_10380,N_9491);
xor U13150 (N_13150,N_9346,N_10277);
and U13151 (N_13151,N_7218,N_11942);
xnor U13152 (N_13152,N_9722,N_9178);
and U13153 (N_13153,N_8451,N_7851);
xnor U13154 (N_13154,N_11907,N_12391);
nand U13155 (N_13155,N_11335,N_9914);
or U13156 (N_13156,N_7867,N_12312);
nor U13157 (N_13157,N_12260,N_7870);
or U13158 (N_13158,N_12353,N_10963);
xnor U13159 (N_13159,N_9400,N_6643);
and U13160 (N_13160,N_8022,N_12467);
and U13161 (N_13161,N_7291,N_8400);
nor U13162 (N_13162,N_10608,N_7449);
nand U13163 (N_13163,N_9309,N_7532);
nand U13164 (N_13164,N_12052,N_11808);
and U13165 (N_13165,N_9469,N_11232);
nor U13166 (N_13166,N_11294,N_11180);
nor U13167 (N_13167,N_8060,N_11121);
nor U13168 (N_13168,N_12160,N_7352);
nor U13169 (N_13169,N_8045,N_6881);
or U13170 (N_13170,N_8580,N_9727);
or U13171 (N_13171,N_9530,N_8238);
and U13172 (N_13172,N_10644,N_6806);
or U13173 (N_13173,N_9463,N_11926);
or U13174 (N_13174,N_9783,N_7285);
or U13175 (N_13175,N_11575,N_11937);
nand U13176 (N_13176,N_12322,N_8987);
xor U13177 (N_13177,N_8267,N_10966);
nand U13178 (N_13178,N_10215,N_7470);
nand U13179 (N_13179,N_11596,N_6890);
nand U13180 (N_13180,N_10025,N_9988);
nor U13181 (N_13181,N_9010,N_11987);
and U13182 (N_13182,N_6433,N_10563);
or U13183 (N_13183,N_8038,N_11014);
nor U13184 (N_13184,N_9403,N_11741);
or U13185 (N_13185,N_6483,N_10100);
nand U13186 (N_13186,N_7009,N_11474);
nor U13187 (N_13187,N_8041,N_10447);
nand U13188 (N_13188,N_7796,N_11255);
nor U13189 (N_13189,N_10982,N_9548);
nand U13190 (N_13190,N_10793,N_8670);
and U13191 (N_13191,N_11630,N_9334);
and U13192 (N_13192,N_9464,N_11006);
nor U13193 (N_13193,N_10346,N_9606);
or U13194 (N_13194,N_9182,N_8282);
and U13195 (N_13195,N_8428,N_8438);
and U13196 (N_13196,N_11119,N_9614);
and U13197 (N_13197,N_7902,N_11431);
or U13198 (N_13198,N_10955,N_9054);
nor U13199 (N_13199,N_9157,N_7894);
or U13200 (N_13200,N_7245,N_10166);
nor U13201 (N_13201,N_11193,N_10128);
or U13202 (N_13202,N_11570,N_11373);
nand U13203 (N_13203,N_7242,N_12094);
or U13204 (N_13204,N_11896,N_7949);
xor U13205 (N_13205,N_12224,N_11490);
nor U13206 (N_13206,N_9452,N_10675);
nand U13207 (N_13207,N_10438,N_9587);
or U13208 (N_13208,N_7196,N_7371);
nor U13209 (N_13209,N_7584,N_12419);
xor U13210 (N_13210,N_6581,N_11691);
nand U13211 (N_13211,N_11543,N_8239);
nand U13212 (N_13212,N_8974,N_6435);
nor U13213 (N_13213,N_9381,N_9200);
and U13214 (N_13214,N_7704,N_9127);
nor U13215 (N_13215,N_6424,N_7274);
nor U13216 (N_13216,N_11037,N_10367);
xnor U13217 (N_13217,N_7931,N_11822);
nand U13218 (N_13218,N_6372,N_10529);
nor U13219 (N_13219,N_11928,N_11151);
nor U13220 (N_13220,N_10546,N_9930);
or U13221 (N_13221,N_11073,N_11009);
nor U13222 (N_13222,N_11154,N_7388);
or U13223 (N_13223,N_12448,N_11145);
nand U13224 (N_13224,N_9025,N_6779);
nor U13225 (N_13225,N_10023,N_9276);
or U13226 (N_13226,N_7029,N_6474);
nor U13227 (N_13227,N_9004,N_8653);
nor U13228 (N_13228,N_11759,N_12165);
nor U13229 (N_13229,N_7407,N_11965);
nand U13230 (N_13230,N_12090,N_7473);
xnor U13231 (N_13231,N_8721,N_10704);
nor U13232 (N_13232,N_11089,N_9944);
xnor U13233 (N_13233,N_11773,N_9508);
and U13234 (N_13234,N_6584,N_6796);
nor U13235 (N_13235,N_7895,N_10570);
or U13236 (N_13236,N_8033,N_8596);
xnor U13237 (N_13237,N_11654,N_9339);
and U13238 (N_13238,N_10836,N_10946);
and U13239 (N_13239,N_9983,N_6537);
or U13240 (N_13240,N_12135,N_11281);
nand U13241 (N_13241,N_12134,N_8169);
nor U13242 (N_13242,N_12152,N_7204);
xnor U13243 (N_13243,N_6595,N_11113);
or U13244 (N_13244,N_6866,N_9188);
or U13245 (N_13245,N_7611,N_10138);
nor U13246 (N_13246,N_9512,N_11372);
nor U13247 (N_13247,N_7847,N_8780);
and U13248 (N_13248,N_9762,N_11587);
or U13249 (N_13249,N_8228,N_9510);
and U13250 (N_13250,N_7116,N_10981);
or U13251 (N_13251,N_10032,N_11434);
nand U13252 (N_13252,N_11055,N_9691);
nor U13253 (N_13253,N_10795,N_8645);
xor U13254 (N_13254,N_10137,N_6804);
and U13255 (N_13255,N_12104,N_9594);
nand U13256 (N_13256,N_12247,N_8867);
or U13257 (N_13257,N_8371,N_11124);
nor U13258 (N_13258,N_9540,N_8541);
and U13259 (N_13259,N_9667,N_9470);
or U13260 (N_13260,N_10229,N_11718);
xnor U13261 (N_13261,N_7499,N_9820);
or U13262 (N_13262,N_6325,N_10662);
and U13263 (N_13263,N_10249,N_11231);
and U13264 (N_13264,N_7915,N_11658);
or U13265 (N_13265,N_7961,N_8314);
and U13266 (N_13266,N_6805,N_9646);
and U13267 (N_13267,N_9544,N_9710);
xor U13268 (N_13268,N_10121,N_7599);
nor U13269 (N_13269,N_12193,N_8385);
nor U13270 (N_13270,N_11692,N_7077);
nand U13271 (N_13271,N_11213,N_6969);
or U13272 (N_13272,N_9281,N_8518);
and U13273 (N_13273,N_11470,N_8830);
and U13274 (N_13274,N_11556,N_6484);
xor U13275 (N_13275,N_6936,N_6398);
nor U13276 (N_13276,N_10107,N_11512);
nor U13277 (N_13277,N_11917,N_7292);
and U13278 (N_13278,N_12201,N_10953);
nor U13279 (N_13279,N_6546,N_11794);
and U13280 (N_13280,N_11506,N_7404);
or U13281 (N_13281,N_8571,N_9566);
nand U13282 (N_13282,N_10991,N_10386);
nand U13283 (N_13283,N_9387,N_6285);
xnor U13284 (N_13284,N_8154,N_11592);
xnor U13285 (N_13285,N_9799,N_10827);
or U13286 (N_13286,N_8588,N_11000);
or U13287 (N_13287,N_11274,N_11859);
xor U13288 (N_13288,N_9643,N_8709);
or U13289 (N_13289,N_9011,N_12216);
or U13290 (N_13290,N_9114,N_7417);
or U13291 (N_13291,N_11387,N_8627);
xnor U13292 (N_13292,N_7975,N_9459);
and U13293 (N_13293,N_9603,N_8275);
and U13294 (N_13294,N_8819,N_9591);
xnor U13295 (N_13295,N_7512,N_9366);
nor U13296 (N_13296,N_9488,N_6882);
nor U13297 (N_13297,N_7823,N_10742);
or U13298 (N_13298,N_9852,N_7869);
nand U13299 (N_13299,N_11429,N_9573);
xor U13300 (N_13300,N_8233,N_6521);
nor U13301 (N_13301,N_7739,N_10973);
nand U13302 (N_13302,N_7344,N_8951);
or U13303 (N_13303,N_9989,N_6900);
and U13304 (N_13304,N_12215,N_11238);
xnor U13305 (N_13305,N_9504,N_10068);
or U13306 (N_13306,N_9843,N_10670);
nand U13307 (N_13307,N_11832,N_7463);
and U13308 (N_13308,N_11035,N_12010);
nor U13309 (N_13309,N_8833,N_9948);
nor U13310 (N_13310,N_11767,N_7063);
xnor U13311 (N_13311,N_10904,N_11801);
or U13312 (N_13312,N_6468,N_11249);
or U13313 (N_13313,N_10829,N_10055);
nand U13314 (N_13314,N_7174,N_11469);
nor U13315 (N_13315,N_9029,N_10680);
nand U13316 (N_13316,N_8497,N_10331);
nand U13317 (N_13317,N_8622,N_10912);
nor U13318 (N_13318,N_6298,N_7746);
xnor U13319 (N_13319,N_6455,N_11471);
nor U13320 (N_13320,N_8838,N_7346);
nor U13321 (N_13321,N_10728,N_10404);
or U13322 (N_13322,N_8308,N_11095);
nor U13323 (N_13323,N_8666,N_7832);
nor U13324 (N_13324,N_7837,N_6439);
or U13325 (N_13325,N_9480,N_9602);
or U13326 (N_13326,N_6402,N_12399);
or U13327 (N_13327,N_6355,N_11573);
nor U13328 (N_13328,N_7405,N_8825);
xnor U13329 (N_13329,N_6861,N_7491);
nand U13330 (N_13330,N_6616,N_10439);
nand U13331 (N_13331,N_8602,N_7129);
or U13332 (N_13332,N_10564,N_12150);
nand U13333 (N_13333,N_9094,N_7113);
or U13334 (N_13334,N_10094,N_8724);
nand U13335 (N_13335,N_12351,N_12330);
nand U13336 (N_13336,N_12466,N_9056);
and U13337 (N_13337,N_10395,N_10299);
or U13338 (N_13338,N_9741,N_6686);
nand U13339 (N_13339,N_7776,N_8217);
and U13340 (N_13340,N_6655,N_11314);
xnor U13341 (N_13341,N_7964,N_8184);
nand U13342 (N_13342,N_9636,N_11820);
nor U13343 (N_13343,N_8494,N_10820);
nor U13344 (N_13344,N_7881,N_12016);
xnor U13345 (N_13345,N_8829,N_11362);
nand U13346 (N_13346,N_8762,N_10018);
nor U13347 (N_13347,N_9721,N_9545);
nand U13348 (N_13348,N_6894,N_10666);
or U13349 (N_13349,N_7883,N_12053);
xor U13350 (N_13350,N_8115,N_6795);
xor U13351 (N_13351,N_10375,N_6363);
or U13352 (N_13352,N_10635,N_8176);
and U13353 (N_13353,N_7448,N_6945);
and U13354 (N_13354,N_8334,N_7697);
xor U13355 (N_13355,N_11459,N_6960);
nor U13356 (N_13356,N_8556,N_7760);
xnor U13357 (N_13357,N_11520,N_7623);
xor U13358 (N_13358,N_7364,N_7335);
and U13359 (N_13359,N_8568,N_12229);
nand U13360 (N_13360,N_9100,N_7925);
nor U13361 (N_13361,N_7787,N_10755);
or U13362 (N_13362,N_7080,N_9335);
and U13363 (N_13363,N_10889,N_10984);
or U13364 (N_13364,N_9968,N_10482);
or U13365 (N_13365,N_8159,N_8922);
or U13366 (N_13366,N_8011,N_12111);
xor U13367 (N_13367,N_6703,N_9307);
nor U13368 (N_13368,N_10278,N_9588);
nor U13369 (N_13369,N_9020,N_9130);
nand U13370 (N_13370,N_6569,N_12290);
and U13371 (N_13371,N_9784,N_7890);
nor U13372 (N_13372,N_10305,N_9973);
xor U13373 (N_13373,N_6721,N_10532);
and U13374 (N_13374,N_12282,N_8145);
nor U13375 (N_13375,N_7031,N_6704);
xnor U13376 (N_13376,N_8536,N_10737);
nor U13377 (N_13377,N_9220,N_7855);
xor U13378 (N_13378,N_10484,N_12098);
nor U13379 (N_13379,N_9899,N_10939);
nand U13380 (N_13380,N_10058,N_7947);
and U13381 (N_13381,N_6858,N_8322);
nand U13382 (N_13382,N_7842,N_11656);
nand U13383 (N_13383,N_8526,N_7495);
and U13384 (N_13384,N_9150,N_11480);
and U13385 (N_13385,N_10611,N_9184);
or U13386 (N_13386,N_11614,N_7091);
and U13387 (N_13387,N_11318,N_7269);
nor U13388 (N_13388,N_9769,N_11452);
and U13389 (N_13389,N_12056,N_11060);
nor U13390 (N_13390,N_8078,N_10938);
nor U13391 (N_13391,N_7328,N_10040);
and U13392 (N_13392,N_10161,N_8394);
xor U13393 (N_13393,N_9642,N_8527);
nand U13394 (N_13394,N_9698,N_7825);
and U13395 (N_13395,N_6951,N_9098);
or U13396 (N_13396,N_9191,N_10042);
or U13397 (N_13397,N_9549,N_11047);
xor U13398 (N_13398,N_6990,N_7744);
nand U13399 (N_13399,N_9092,N_11002);
nor U13400 (N_13400,N_8793,N_8860);
xnor U13401 (N_13401,N_11256,N_10964);
nor U13402 (N_13402,N_11320,N_9185);
nand U13403 (N_13403,N_6846,N_10916);
nand U13404 (N_13404,N_9392,N_8183);
nor U13405 (N_13405,N_9785,N_11982);
nor U13406 (N_13406,N_8455,N_10425);
nand U13407 (N_13407,N_11137,N_12313);
nand U13408 (N_13408,N_12476,N_9965);
nand U13409 (N_13409,N_10937,N_9013);
nor U13410 (N_13410,N_7277,N_11171);
nor U13411 (N_13411,N_6700,N_8452);
and U13412 (N_13412,N_6531,N_11174);
and U13413 (N_13413,N_6920,N_8392);
nor U13414 (N_13414,N_12189,N_6695);
nor U13415 (N_13415,N_10097,N_7400);
or U13416 (N_13416,N_6451,N_9787);
and U13417 (N_13417,N_11786,N_9938);
nor U13418 (N_13418,N_11579,N_10390);
nor U13419 (N_13419,N_11802,N_11446);
nor U13420 (N_13420,N_11612,N_11624);
nand U13421 (N_13421,N_11912,N_8000);
nand U13422 (N_13422,N_9570,N_11086);
or U13423 (N_13423,N_6460,N_11103);
nand U13424 (N_13424,N_8206,N_7878);
nor U13425 (N_13425,N_12458,N_11504);
nor U13426 (N_13426,N_9754,N_10746);
nor U13427 (N_13427,N_10775,N_10066);
nor U13428 (N_13428,N_10902,N_12037);
nand U13429 (N_13429,N_8848,N_7148);
xnor U13430 (N_13430,N_12236,N_12086);
xor U13431 (N_13431,N_12108,N_7908);
nor U13432 (N_13432,N_11296,N_6294);
and U13433 (N_13433,N_9880,N_9936);
and U13434 (N_13434,N_7071,N_8758);
nor U13435 (N_13435,N_10363,N_8877);
nand U13436 (N_13436,N_7251,N_9066);
or U13437 (N_13437,N_7176,N_9050);
or U13438 (N_13438,N_7373,N_9413);
xor U13439 (N_13439,N_10760,N_10101);
nor U13440 (N_13440,N_6339,N_8182);
xnor U13441 (N_13441,N_8677,N_7780);
and U13442 (N_13442,N_12102,N_11526);
and U13443 (N_13443,N_6764,N_8064);
nor U13444 (N_13444,N_9109,N_7107);
nor U13445 (N_13445,N_8478,N_6778);
nand U13446 (N_13446,N_6692,N_7078);
nand U13447 (N_13447,N_8237,N_7600);
or U13448 (N_13448,N_12018,N_8367);
nor U13449 (N_13449,N_9652,N_12082);
nor U13450 (N_13450,N_11876,N_11574);
and U13451 (N_13451,N_9971,N_11943);
or U13452 (N_13452,N_11282,N_7543);
xnor U13453 (N_13453,N_10540,N_7879);
nand U13454 (N_13454,N_9969,N_11327);
and U13455 (N_13455,N_11160,N_9149);
and U13456 (N_13456,N_11763,N_7457);
xor U13457 (N_13457,N_10332,N_8875);
and U13458 (N_13458,N_7162,N_7759);
nand U13459 (N_13459,N_7239,N_8868);
and U13460 (N_13460,N_6854,N_9500);
xor U13461 (N_13461,N_10923,N_8715);
xor U13462 (N_13462,N_9970,N_12493);
nor U13463 (N_13463,N_11514,N_10472);
xor U13464 (N_13464,N_11264,N_8885);
or U13465 (N_13465,N_10740,N_11298);
nor U13466 (N_13466,N_8917,N_6670);
or U13467 (N_13467,N_11861,N_10637);
xor U13468 (N_13468,N_8009,N_12398);
or U13469 (N_13469,N_7560,N_10398);
xnor U13470 (N_13470,N_9456,N_9359);
xnor U13471 (N_13471,N_8972,N_11149);
xnor U13472 (N_13472,N_12069,N_12220);
nand U13473 (N_13473,N_9478,N_8643);
nor U13474 (N_13474,N_10690,N_6459);
or U13475 (N_13475,N_11063,N_10593);
nor U13476 (N_13476,N_6625,N_8335);
or U13477 (N_13477,N_7396,N_7357);
nand U13478 (N_13478,N_11622,N_10466);
or U13479 (N_13479,N_7984,N_7225);
nand U13480 (N_13480,N_7602,N_9599);
and U13481 (N_13481,N_7987,N_8886);
nor U13482 (N_13482,N_8861,N_8671);
xnor U13483 (N_13483,N_7781,N_10185);
xnor U13484 (N_13484,N_7989,N_9915);
nand U13485 (N_13485,N_11713,N_8333);
xnor U13486 (N_13486,N_8701,N_6874);
nor U13487 (N_13487,N_10053,N_10553);
or U13488 (N_13488,N_11079,N_6717);
nand U13489 (N_13489,N_10208,N_6706);
nor U13490 (N_13490,N_9123,N_10530);
nand U13491 (N_13491,N_7997,N_6300);
nor U13492 (N_13492,N_6553,N_8429);
or U13493 (N_13493,N_11004,N_8359);
or U13494 (N_13494,N_10808,N_6777);
and U13495 (N_13495,N_9498,N_8318);
or U13496 (N_13496,N_10592,N_6347);
nor U13497 (N_13497,N_11250,N_6923);
nor U13498 (N_13498,N_10289,N_12288);
nor U13499 (N_13499,N_12040,N_8402);
and U13500 (N_13500,N_11897,N_8707);
or U13501 (N_13501,N_9358,N_8109);
xnor U13502 (N_13502,N_7607,N_10705);
and U13503 (N_13503,N_6985,N_7422);
or U13504 (N_13504,N_12141,N_10262);
nor U13505 (N_13505,N_7690,N_9837);
nand U13506 (N_13506,N_8613,N_11341);
or U13507 (N_13507,N_7030,N_11743);
xor U13508 (N_13508,N_7003,N_9660);
nor U13509 (N_13509,N_7458,N_8460);
or U13510 (N_13510,N_6276,N_9697);
nor U13511 (N_13511,N_10877,N_6283);
or U13512 (N_13512,N_11554,N_8058);
or U13513 (N_13513,N_10070,N_8124);
nand U13514 (N_13514,N_9147,N_9845);
xnor U13515 (N_13515,N_12231,N_8770);
and U13516 (N_13516,N_11176,N_10747);
and U13517 (N_13517,N_10701,N_12257);
xnor U13518 (N_13518,N_11999,N_8975);
or U13519 (N_13519,N_12238,N_8459);
xnor U13520 (N_13520,N_12013,N_12170);
xor U13521 (N_13521,N_10967,N_6379);
xnor U13522 (N_13522,N_11029,N_7416);
nor U13523 (N_13523,N_7809,N_6940);
nor U13524 (N_13524,N_12024,N_10789);
xor U13525 (N_13525,N_7057,N_7293);
nor U13526 (N_13526,N_11576,N_10812);
nor U13527 (N_13527,N_7167,N_12119);
xnor U13528 (N_13528,N_9704,N_8789);
nor U13529 (N_13529,N_10809,N_12109);
nand U13530 (N_13530,N_7141,N_8390);
nand U13531 (N_13531,N_8934,N_10999);
or U13532 (N_13532,N_11319,N_7189);
and U13533 (N_13533,N_6295,N_6776);
and U13534 (N_13534,N_8215,N_7348);
or U13535 (N_13535,N_8105,N_11855);
xnor U13536 (N_13536,N_11787,N_10399);
nand U13537 (N_13537,N_8864,N_7835);
nor U13538 (N_13538,N_6621,N_10948);
xor U13539 (N_13539,N_9490,N_11838);
and U13540 (N_13540,N_7510,N_8023);
nor U13541 (N_13541,N_7163,N_9090);
nand U13542 (N_13542,N_8509,N_10560);
nor U13543 (N_13543,N_8767,N_12459);
and U13544 (N_13544,N_11555,N_10312);
nand U13545 (N_13545,N_10154,N_12273);
xor U13546 (N_13546,N_8448,N_11034);
or U13547 (N_13547,N_10476,N_8286);
nor U13548 (N_13548,N_9782,N_7368);
xnor U13549 (N_13549,N_10551,N_11153);
or U13550 (N_13550,N_8341,N_8565);
nor U13551 (N_13551,N_10124,N_10171);
and U13552 (N_13552,N_8486,N_6382);
and U13553 (N_13553,N_7468,N_12114);
nand U13554 (N_13554,N_11336,N_7893);
or U13555 (N_13555,N_8740,N_12363);
or U13556 (N_13556,N_7190,N_11332);
and U13557 (N_13557,N_9868,N_10591);
nand U13558 (N_13558,N_10298,N_11202);
nand U13559 (N_13559,N_10713,N_7628);
nor U13560 (N_13560,N_11201,N_9058);
nor U13561 (N_13561,N_6989,N_7445);
xor U13562 (N_13562,N_8244,N_7946);
and U13563 (N_13563,N_10105,N_7409);
and U13564 (N_13564,N_7865,N_8187);
and U13565 (N_13565,N_9890,N_8175);
or U13566 (N_13566,N_10669,N_9932);
or U13567 (N_13567,N_7733,N_8338);
and U13568 (N_13568,N_6741,N_9475);
xnor U13569 (N_13569,N_10411,N_10875);
or U13570 (N_13570,N_7556,N_7302);
and U13571 (N_13571,N_10266,N_6836);
and U13572 (N_13572,N_10873,N_9589);
xnor U13573 (N_13573,N_9889,N_6681);
xnor U13574 (N_13574,N_11021,N_11705);
and U13575 (N_13575,N_9726,N_11138);
or U13576 (N_13576,N_9493,N_12063);
or U13577 (N_13577,N_10801,N_12405);
nand U13578 (N_13578,N_11666,N_7500);
nor U13579 (N_13579,N_7202,N_12103);
or U13580 (N_13580,N_9390,N_11163);
xor U13581 (N_13581,N_9729,N_10777);
or U13582 (N_13582,N_9032,N_7896);
nor U13583 (N_13583,N_7530,N_7135);
and U13584 (N_13584,N_11258,N_9101);
nand U13585 (N_13585,N_8896,N_9857);
xor U13586 (N_13586,N_11979,N_7914);
xnor U13587 (N_13587,N_6734,N_11539);
nor U13588 (N_13588,N_8440,N_11148);
nor U13589 (N_13589,N_7019,N_11701);
or U13590 (N_13590,N_11357,N_10355);
nor U13591 (N_13591,N_6384,N_11849);
and U13592 (N_13592,N_11020,N_8718);
xnor U13593 (N_13593,N_11984,N_8208);
xor U13594 (N_13594,N_11027,N_7617);
nor U13595 (N_13595,N_11750,N_11078);
nor U13596 (N_13596,N_12489,N_12357);
xnor U13597 (N_13597,N_6273,N_9299);
or U13598 (N_13598,N_10954,N_6761);
nand U13599 (N_13599,N_12309,N_7701);
or U13600 (N_13600,N_6694,N_11036);
or U13601 (N_13601,N_7596,N_9984);
or U13602 (N_13602,N_9026,N_9081);
nand U13603 (N_13603,N_9009,N_10547);
xor U13604 (N_13604,N_10174,N_11288);
xor U13605 (N_13605,N_8150,N_9408);
or U13606 (N_13606,N_11532,N_11170);
and U13607 (N_13607,N_6675,N_8878);
or U13608 (N_13608,N_11872,N_7389);
and U13609 (N_13609,N_8085,N_6956);
nand U13610 (N_13610,N_9559,N_11334);
and U13611 (N_13611,N_12368,N_8210);
and U13612 (N_13612,N_7917,N_12110);
and U13613 (N_13613,N_9347,N_10416);
nand U13614 (N_13614,N_8797,N_10824);
xnor U13615 (N_13615,N_9886,N_8091);
nand U13616 (N_13616,N_12159,N_10159);
nor U13617 (N_13617,N_11098,N_7619);
nand U13618 (N_13618,N_7016,N_7319);
and U13619 (N_13619,N_7555,N_8224);
and U13620 (N_13620,N_6737,N_10031);
nand U13621 (N_13621,N_7820,N_10246);
nor U13622 (N_13622,N_6441,N_9647);
or U13623 (N_13623,N_12468,N_11974);
and U13624 (N_13624,N_9446,N_6593);
nor U13625 (N_13625,N_8490,N_7940);
nand U13626 (N_13626,N_11203,N_10024);
nand U13627 (N_13627,N_10843,N_7264);
xnor U13628 (N_13628,N_6684,N_11130);
nor U13629 (N_13629,N_10559,N_11453);
nor U13630 (N_13630,N_8801,N_10748);
nand U13631 (N_13631,N_8630,N_7963);
xor U13632 (N_13632,N_6256,N_7301);
and U13633 (N_13633,N_8360,N_7297);
xor U13634 (N_13634,N_6839,N_9450);
nand U13635 (N_13635,N_11381,N_8837);
xnor U13636 (N_13636,N_7840,N_11651);
nor U13637 (N_13637,N_8487,N_6517);
nor U13638 (N_13638,N_6534,N_6909);
xor U13639 (N_13639,N_6928,N_10431);
nor U13640 (N_13640,N_9487,N_10245);
or U13641 (N_13641,N_6824,N_11432);
xnor U13642 (N_13642,N_10047,N_8792);
and U13643 (N_13643,N_8503,N_8955);
and U13644 (N_13644,N_6793,N_10696);
and U13645 (N_13645,N_7055,N_10280);
nor U13646 (N_13646,N_12025,N_10583);
or U13647 (N_13647,N_8162,N_9063);
or U13648 (N_13648,N_9353,N_11326);
xor U13649 (N_13649,N_7816,N_8909);
xor U13650 (N_13650,N_6281,N_7791);
xnor U13651 (N_13651,N_7996,N_9164);
nand U13652 (N_13652,N_10318,N_12079);
nand U13653 (N_13653,N_8117,N_8977);
and U13654 (N_13654,N_12256,N_10850);
or U13655 (N_13655,N_9584,N_7418);
xnor U13656 (N_13656,N_9146,N_10364);
or U13657 (N_13657,N_10309,N_9620);
and U13658 (N_13658,N_8012,N_6383);
or U13659 (N_13659,N_12378,N_7153);
nor U13660 (N_13660,N_12490,N_12499);
nand U13661 (N_13661,N_8549,N_8507);
or U13662 (N_13662,N_7743,N_7631);
nor U13663 (N_13663,N_9705,N_9465);
and U13664 (N_13664,N_9148,N_11537);
and U13665 (N_13665,N_11678,N_11870);
xor U13666 (N_13666,N_12455,N_9788);
xnor U13667 (N_13667,N_12065,N_10200);
or U13668 (N_13668,N_12071,N_10442);
and U13669 (N_13669,N_10947,N_10020);
nand U13670 (N_13670,N_11378,N_8477);
nand U13671 (N_13671,N_10722,N_8858);
or U13672 (N_13672,N_12070,N_11807);
xnor U13673 (N_13673,N_10977,N_7508);
nand U13674 (N_13674,N_9861,N_10677);
and U13675 (N_13675,N_9987,N_11115);
nand U13676 (N_13676,N_8869,N_6527);
xnor U13677 (N_13677,N_10767,N_6539);
nand U13678 (N_13678,N_7035,N_9273);
nor U13679 (N_13679,N_7002,N_12480);
or U13680 (N_13680,N_6370,N_11050);
or U13681 (N_13681,N_10691,N_10610);
or U13682 (N_13682,N_7255,N_7942);
xnor U13683 (N_13683,N_10005,N_11785);
and U13684 (N_13684,N_6860,N_11618);
and U13685 (N_13685,N_10727,N_7794);
nor U13686 (N_13686,N_10417,N_7651);
nand U13687 (N_13687,N_7489,N_8887);
and U13688 (N_13688,N_8649,N_11454);
xor U13689 (N_13689,N_8730,N_8750);
or U13690 (N_13690,N_7183,N_8221);
nor U13691 (N_13691,N_10684,N_10522);
nand U13692 (N_13692,N_6310,N_11390);
nor U13693 (N_13693,N_9739,N_10115);
nor U13694 (N_13694,N_11619,N_10656);
nand U13695 (N_13695,N_8831,N_10218);
and U13696 (N_13696,N_6427,N_10649);
nor U13697 (N_13697,N_8034,N_11393);
nor U13698 (N_13698,N_7876,N_10090);
xnor U13699 (N_13699,N_10340,N_11505);
xnor U13700 (N_13700,N_10488,N_8437);
nand U13701 (N_13701,N_10306,N_9197);
and U13702 (N_13702,N_8901,N_12146);
nor U13703 (N_13703,N_7106,N_6794);
and U13704 (N_13704,N_8500,N_12446);
nor U13705 (N_13705,N_11790,N_12112);
xnor U13706 (N_13706,N_7324,N_12291);
nand U13707 (N_13707,N_9419,N_6565);
xnor U13708 (N_13708,N_10647,N_7561);
xor U13709 (N_13709,N_10033,N_11467);
nor U13710 (N_13710,N_6938,N_7520);
or U13711 (N_13711,N_12030,N_7943);
nor U13712 (N_13712,N_11306,N_6590);
nor U13713 (N_13713,N_8958,N_6925);
xor U13714 (N_13714,N_12183,N_11437);
xnor U13715 (N_13715,N_11853,N_10391);
nand U13716 (N_13716,N_12470,N_10006);
and U13717 (N_13717,N_6688,N_7998);
nand U13718 (N_13718,N_9986,N_8281);
nand U13719 (N_13719,N_11655,N_8966);
nand U13720 (N_13720,N_6634,N_7574);
nand U13721 (N_13721,N_12422,N_12218);
or U13722 (N_13722,N_9141,N_10183);
or U13723 (N_13723,N_6732,N_12054);
nor U13724 (N_13724,N_9682,N_11951);
nand U13725 (N_13725,N_11712,N_12366);
nor U13726 (N_13726,N_8952,N_9712);
or U13727 (N_13727,N_11065,N_6381);
and U13728 (N_13728,N_7634,N_6707);
or U13729 (N_13729,N_11915,N_6876);
or U13730 (N_13730,N_9972,N_8519);
or U13731 (N_13731,N_8821,N_11088);
xnor U13732 (N_13732,N_10044,N_12142);
xnor U13733 (N_13733,N_8137,N_12307);
nor U13734 (N_13734,N_9807,N_11455);
nand U13735 (N_13735,N_9596,N_7721);
xnor U13736 (N_13736,N_11594,N_8914);
xnor U13737 (N_13737,N_8019,N_11466);
and U13738 (N_13738,N_6606,N_10773);
or U13739 (N_13739,N_10567,N_9234);
nor U13740 (N_13740,N_8550,N_6607);
or U13741 (N_13741,N_11305,N_12409);
nor U13742 (N_13742,N_10192,N_8601);
nor U13743 (N_13743,N_8387,N_7036);
nand U13744 (N_13744,N_12383,N_7296);
and U13745 (N_13745,N_8683,N_8193);
and U13746 (N_13746,N_8099,N_7097);
or U13747 (N_13747,N_10320,N_6369);
nor U13748 (N_13748,N_10883,N_10730);
and U13749 (N_13749,N_9831,N_6637);
and U13750 (N_13750,N_10426,N_12432);
or U13751 (N_13751,N_7748,N_8540);
or U13752 (N_13752,N_10485,N_7995);
nor U13753 (N_13753,N_8298,N_10144);
xor U13754 (N_13754,N_7377,N_12263);
xnor U13755 (N_13755,N_9849,N_12456);
nor U13756 (N_13756,N_8757,N_10857);
nand U13757 (N_13757,N_10935,N_11646);
or U13758 (N_13758,N_8585,N_8891);
nor U13759 (N_13759,N_7612,N_12431);
or U13760 (N_13760,N_8343,N_11064);
and U13761 (N_13761,N_8468,N_10555);
nand U13762 (N_13762,N_7647,N_8569);
nor U13763 (N_13763,N_10835,N_10302);
nor U13764 (N_13764,N_10248,N_7232);
and U13765 (N_13765,N_7609,N_11012);
nand U13766 (N_13766,N_7858,N_8599);
nand U13767 (N_13767,N_8930,N_9162);
and U13768 (N_13768,N_6630,N_11280);
nor U13769 (N_13769,N_12452,N_11990);
xor U13770 (N_13770,N_10226,N_9509);
nand U13771 (N_13771,N_8433,N_10452);
and U13772 (N_13772,N_12149,N_9080);
or U13773 (N_13773,N_6663,N_8453);
nand U13774 (N_13774,N_9927,N_7913);
nor U13775 (N_13775,N_9719,N_9135);
or U13776 (N_13776,N_9499,N_10945);
and U13777 (N_13777,N_7764,N_12096);
nor U13778 (N_13778,N_9776,N_7519);
or U13779 (N_13779,N_12382,N_6320);
nor U13780 (N_13780,N_7493,N_8070);
xor U13781 (N_13781,N_7683,N_7527);
or U13782 (N_13782,N_12122,N_9068);
xnor U13783 (N_13783,N_9483,N_9898);
and U13784 (N_13784,N_10209,N_9937);
or U13785 (N_13785,N_10557,N_9892);
or U13786 (N_13786,N_9678,N_7676);
and U13787 (N_13787,N_7626,N_12373);
or U13788 (N_13788,N_11519,N_9174);
and U13789 (N_13789,N_8227,N_7070);
or U13790 (N_13790,N_12329,N_12249);
or U13791 (N_13791,N_11782,N_6784);
or U13792 (N_13792,N_11699,N_7814);
xor U13793 (N_13793,N_8806,N_12158);
nand U13794 (N_13794,N_6399,N_6912);
nor U13795 (N_13795,N_9074,N_7830);
and U13796 (N_13796,N_10285,N_10575);
nor U13797 (N_13797,N_11567,N_11198);
or U13798 (N_13798,N_9073,N_9567);
and U13799 (N_13799,N_10129,N_7754);
nand U13800 (N_13800,N_7004,N_9841);
nor U13801 (N_13801,N_9202,N_9422);
nor U13802 (N_13802,N_11755,N_6308);
or U13803 (N_13803,N_10374,N_6397);
xor U13804 (N_13804,N_9298,N_9022);
and U13805 (N_13805,N_12245,N_6752);
xor U13806 (N_13806,N_12058,N_8968);
xor U13807 (N_13807,N_10763,N_8126);
nor U13808 (N_13808,N_10180,N_7773);
or U13809 (N_13809,N_9235,N_8449);
nand U13810 (N_13810,N_11024,N_10825);
and U13811 (N_13811,N_6288,N_9224);
xnor U13812 (N_13812,N_12387,N_9929);
and U13813 (N_13813,N_7164,N_10011);
or U13814 (N_13814,N_10569,N_10846);
nor U13815 (N_13815,N_12325,N_11435);
xnor U13816 (N_13816,N_6921,N_11679);
and U13817 (N_13817,N_8641,N_6635);
and U13818 (N_13818,N_10433,N_6530);
or U13819 (N_13819,N_8856,N_12361);
and U13820 (N_13820,N_11816,N_10787);
nand U13821 (N_13821,N_12465,N_9412);
nand U13822 (N_13822,N_11243,N_11793);
nor U13823 (N_13823,N_12438,N_9126);
or U13824 (N_13824,N_12344,N_11093);
or U13825 (N_13825,N_7763,N_9531);
nand U13826 (N_13826,N_7516,N_11234);
and U13827 (N_13827,N_9724,N_6811);
or U13828 (N_13828,N_9069,N_8824);
nand U13829 (N_13829,N_12107,N_10441);
nor U13830 (N_13830,N_9925,N_9750);
nor U13831 (N_13831,N_8688,N_6306);
nor U13832 (N_13832,N_10310,N_6726);
or U13833 (N_13833,N_8356,N_8651);
xor U13834 (N_13834,N_6532,N_6554);
nand U13835 (N_13835,N_9629,N_11144);
nor U13836 (N_13836,N_11175,N_9610);
and U13837 (N_13837,N_11660,N_6649);
or U13838 (N_13838,N_8381,N_10460);
or U13839 (N_13839,N_8025,N_10337);
or U13840 (N_13840,N_11242,N_8817);
or U13841 (N_13841,N_9913,N_11397);
and U13842 (N_13842,N_6955,N_8158);
nand U13843 (N_13843,N_9270,N_11025);
or U13844 (N_13844,N_9541,N_10381);
nor U13845 (N_13845,N_9317,N_7011);
xnor U13846 (N_13846,N_6326,N_10155);
or U13847 (N_13847,N_10578,N_10338);
nor U13848 (N_13848,N_11152,N_11631);
xor U13849 (N_13849,N_8990,N_7332);
and U13850 (N_13850,N_11629,N_7531);
and U13851 (N_13851,N_10354,N_7551);
xor U13852 (N_13852,N_7138,N_8913);
and U13853 (N_13853,N_7972,N_9502);
xor U13854 (N_13854,N_7538,N_8739);
and U13855 (N_13855,N_12457,N_11077);
xnor U13856 (N_13856,N_12120,N_8999);
and U13857 (N_13857,N_6345,N_9264);
nor U13858 (N_13858,N_11775,N_8820);
xor U13859 (N_13859,N_8042,N_10880);
xnor U13860 (N_13860,N_6749,N_11497);
nor U13861 (N_13861,N_9035,N_6588);
nand U13862 (N_13862,N_7406,N_10400);
or U13863 (N_13863,N_10059,N_6972);
and U13864 (N_13864,N_7238,N_8735);
nor U13865 (N_13865,N_12370,N_11263);
xor U13866 (N_13866,N_10369,N_6753);
or U13867 (N_13867,N_11998,N_8612);
and U13868 (N_13868,N_7567,N_6472);
nor U13869 (N_13869,N_7926,N_6336);
nor U13870 (N_13870,N_9595,N_11071);
xor U13871 (N_13871,N_7286,N_6877);
nand U13872 (N_13872,N_6321,N_11495);
xor U13873 (N_13873,N_11084,N_10377);
xnor U13874 (N_13874,N_10109,N_7639);
nand U13875 (N_13875,N_11935,N_9862);
nor U13876 (N_13876,N_12286,N_10606);
nand U13877 (N_13877,N_9982,N_9104);
xnor U13878 (N_13878,N_9657,N_7900);
or U13879 (N_13879,N_7090,N_7675);
and U13880 (N_13880,N_8010,N_8432);
nand U13881 (N_13881,N_7487,N_6599);
and U13882 (N_13882,N_11799,N_11597);
or U13883 (N_13883,N_10463,N_9815);
xnor U13884 (N_13884,N_7040,N_7032);
nand U13885 (N_13885,N_12272,N_9269);
nand U13886 (N_13886,N_8799,N_7498);
nor U13887 (N_13887,N_8777,N_9154);
or U13888 (N_13888,N_7227,N_9801);
nand U13889 (N_13889,N_9571,N_10060);
nand U13890 (N_13890,N_8171,N_11628);
and U13891 (N_13891,N_6922,N_11483);
or U13892 (N_13892,N_10237,N_9277);
nor U13893 (N_13893,N_9827,N_9878);
or U13894 (N_13894,N_7525,N_11757);
nor U13895 (N_13895,N_8264,N_6699);
nand U13896 (N_13896,N_7211,N_7800);
xnor U13897 (N_13897,N_9239,N_10845);
nor U13898 (N_13898,N_8295,N_7622);
xor U13899 (N_13899,N_8849,N_9521);
and U13900 (N_13900,N_7707,N_11092);
and U13901 (N_13901,N_6958,N_11966);
nand U13902 (N_13902,N_8321,N_10533);
xor U13903 (N_13903,N_10832,N_8751);
nor U13904 (N_13904,N_10089,N_6792);
xnor U13905 (N_13905,N_6862,N_9133);
nor U13906 (N_13906,N_10317,N_11132);
nor U13907 (N_13907,N_11569,N_7038);
or U13908 (N_13908,N_7797,N_9003);
nand U13909 (N_13909,N_12011,N_6889);
or U13910 (N_13910,N_12200,N_8574);
or U13911 (N_13911,N_11440,N_8752);
nor U13912 (N_13912,N_8538,N_9555);
xnor U13913 (N_13913,N_9447,N_8123);
nand U13914 (N_13914,N_11682,N_10839);
or U13915 (N_13915,N_8073,N_11602);
nand U13916 (N_13916,N_7819,N_10856);
or U13917 (N_13917,N_9976,N_9107);
nand U13918 (N_13918,N_11147,N_7546);
xnor U13919 (N_13919,N_12461,N_6971);
nor U13920 (N_13920,N_11360,N_11195);
nand U13921 (N_13921,N_11207,N_6624);
nor U13922 (N_13922,N_7420,N_7145);
nand U13923 (N_13923,N_11028,N_9286);
or U13924 (N_13924,N_10074,N_6786);
or U13925 (N_13925,N_9117,N_10136);
or U13926 (N_13926,N_9284,N_9744);
nand U13927 (N_13927,N_8220,N_9811);
xor U13928 (N_13928,N_10456,N_11363);
and U13929 (N_13929,N_8354,N_8947);
nor U13930 (N_13930,N_10734,N_12403);
or U13931 (N_13931,N_11489,N_12303);
xor U13932 (N_13932,N_6535,N_7044);
and U13933 (N_13933,N_6611,N_8422);
nand U13934 (N_13934,N_11053,N_8978);
nand U13935 (N_13935,N_11652,N_10496);
and U13936 (N_13936,N_10478,N_7859);
nand U13937 (N_13937,N_11717,N_12147);
and U13938 (N_13938,N_9860,N_6935);
nor U13939 (N_13939,N_11010,N_12270);
or U13940 (N_13940,N_11833,N_8980);
nand U13941 (N_13941,N_8462,N_8803);
or U13942 (N_13942,N_10102,N_8270);
and U13943 (N_13943,N_12241,N_10199);
nand U13944 (N_13944,N_6513,N_6837);
nand U13945 (N_13945,N_7103,N_7514);
and U13946 (N_13946,N_6765,N_12172);
nor U13947 (N_13947,N_10313,N_9887);
xnor U13948 (N_13948,N_7144,N_10118);
nor U13949 (N_13949,N_11392,N_11136);
and U13950 (N_13950,N_10989,N_6810);
or U13951 (N_13951,N_11427,N_7788);
nand U13952 (N_13952,N_7154,N_9431);
and U13953 (N_13953,N_7208,N_7392);
or U13954 (N_13954,N_7650,N_12390);
xor U13955 (N_13955,N_10543,N_11482);
nand U13956 (N_13956,N_12184,N_12334);
nand U13957 (N_13957,N_9655,N_10661);
nor U13958 (N_13958,N_8695,N_9891);
nand U13959 (N_13959,N_11899,N_6875);
and U13960 (N_13960,N_7547,N_7863);
xnor U13961 (N_13961,N_11711,N_11980);
nand U13962 (N_13962,N_8483,N_8450);
xor U13963 (N_13963,N_12181,N_12015);
nand U13964 (N_13964,N_7401,N_7340);
nor U13965 (N_13965,N_10157,N_7421);
nor U13966 (N_13966,N_11672,N_11923);
nand U13967 (N_13967,N_10394,N_8605);
nand U13968 (N_13968,N_10048,N_8180);
nor U13969 (N_13969,N_11901,N_11867);
or U13970 (N_13970,N_9451,N_10158);
nor U13971 (N_13971,N_11377,N_6883);
and U13972 (N_13972,N_10095,N_10451);
nand U13973 (N_13973,N_7210,N_6356);
and U13974 (N_13974,N_9190,N_6782);
nand U13975 (N_13975,N_11826,N_9016);
nor U13976 (N_13976,N_9356,N_7887);
and U13977 (N_13977,N_8826,N_8464);
or U13978 (N_13978,N_12073,N_8593);
or U13979 (N_13979,N_6816,N_9015);
nand U13980 (N_13980,N_7875,N_10550);
xnor U13981 (N_13981,N_7570,N_9305);
or U13982 (N_13982,N_9173,N_12317);
and U13983 (N_13983,N_7656,N_7331);
nor U13984 (N_13984,N_12440,N_10348);
and U13985 (N_13985,N_10362,N_8535);
or U13986 (N_13986,N_10716,N_6760);
nand U13987 (N_13987,N_10625,N_10762);
nor U13988 (N_13988,N_9139,N_9761);
and U13989 (N_13989,N_9342,N_7254);
nand U13990 (N_13990,N_10673,N_9967);
or U13991 (N_13991,N_7272,N_6892);
xnor U13992 (N_13992,N_10500,N_6421);
or U13993 (N_13993,N_6568,N_11244);
nand U13994 (N_13994,N_8680,N_8434);
xor U13995 (N_13995,N_9350,N_8700);
xnor U13996 (N_13996,N_6769,N_7186);
xor U13997 (N_13997,N_11273,N_10974);
and U13998 (N_13998,N_9617,N_10771);
and U13999 (N_13999,N_8916,N_9360);
or U14000 (N_14000,N_7258,N_6976);
nor U14001 (N_14001,N_9767,N_6631);
nor U14002 (N_14002,N_11783,N_11991);
nand U14003 (N_14003,N_7215,N_9565);
xnor U14004 (N_14004,N_9600,N_9060);
nand U14005 (N_14005,N_11216,N_7432);
xnor U14006 (N_14006,N_9393,N_11409);
or U14007 (N_14007,N_12497,N_8226);
and U14008 (N_14008,N_10471,N_6605);
nor U14009 (N_14009,N_6639,N_10010);
nand U14010 (N_14010,N_11371,N_11557);
nand U14011 (N_14011,N_10643,N_11595);
nor U14012 (N_14012,N_10491,N_8398);
and U14013 (N_14013,N_6859,N_6623);
and U14014 (N_14014,N_6924,N_9597);
nand U14015 (N_14015,N_9873,N_10085);
and U14016 (N_14016,N_12100,N_11507);
and U14017 (N_14017,N_9229,N_6480);
nor U14018 (N_14018,N_6937,N_7568);
and U14019 (N_14019,N_7712,N_9039);
nor U14020 (N_14020,N_10910,N_7479);
or U14021 (N_14021,N_11938,N_8095);
xor U14022 (N_14022,N_7708,N_11754);
nor U14023 (N_14023,N_8028,N_7985);
and U14024 (N_14024,N_7320,N_7719);
nand U14025 (N_14025,N_7962,N_10936);
nand U14026 (N_14026,N_10228,N_10083);
xor U14027 (N_14027,N_7909,N_9904);
nor U14028 (N_14028,N_8083,N_9266);
and U14029 (N_14029,N_11383,N_11529);
nor U14030 (N_14030,N_8142,N_6360);
or U14031 (N_14031,N_6957,N_9879);
nor U14032 (N_14032,N_6542,N_6927);
xnor U14033 (N_14033,N_6592,N_6893);
nand U14034 (N_14034,N_11165,N_7982);
nand U14035 (N_14035,N_7954,N_12301);
nand U14036 (N_14036,N_11473,N_7336);
nor U14037 (N_14037,N_11862,N_7240);
and U14038 (N_14038,N_12486,N_9507);
nor U14039 (N_14039,N_6656,N_10523);
nand U14040 (N_14040,N_8279,N_7671);
or U14041 (N_14041,N_10508,N_10241);
or U14042 (N_14042,N_8584,N_6727);
or U14043 (N_14043,N_6926,N_12287);
nor U14044 (N_14044,N_11809,N_8902);
or U14045 (N_14045,N_12275,N_8832);
xnor U14046 (N_14046,N_10739,N_6376);
xnor U14047 (N_14047,N_9781,N_9882);
nand U14048 (N_14048,N_9519,N_7505);
or U14049 (N_14049,N_11399,N_11753);
nor U14050 (N_14050,N_11048,N_12038);
nand U14051 (N_14051,N_8492,N_12235);
and U14052 (N_14052,N_11634,N_10339);
nand U14053 (N_14053,N_7644,N_7474);
and U14054 (N_14054,N_6831,N_11523);
nand U14055 (N_14055,N_8648,N_10890);
or U14056 (N_14056,N_11922,N_7014);
or U14057 (N_14057,N_7853,N_9666);
or U14058 (N_14058,N_7261,N_7740);
nor U14059 (N_14059,N_7515,N_6648);
nand U14060 (N_14060,N_12401,N_7093);
xor U14061 (N_14061,N_10765,N_6697);
nor U14062 (N_14062,N_7386,N_6570);
or U14063 (N_14063,N_10418,N_10041);
and U14064 (N_14064,N_6415,N_7076);
nor U14065 (N_14065,N_12194,N_12001);
and U14066 (N_14066,N_11358,N_11125);
nor U14067 (N_14067,N_11493,N_6849);
or U14068 (N_14068,N_9027,N_8044);
or U14069 (N_14069,N_12374,N_7015);
xnor U14070 (N_14070,N_9920,N_10894);
and U14071 (N_14071,N_8517,N_7337);
nor U14072 (N_14072,N_11382,N_8178);
and U14073 (N_14073,N_9322,N_8128);
or U14074 (N_14074,N_12460,N_8303);
and U14075 (N_14075,N_9370,N_11731);
nand U14076 (N_14076,N_10497,N_8241);
xor U14077 (N_14077,N_11673,N_9686);
and U14078 (N_14078,N_8485,N_11600);
or U14079 (N_14079,N_6386,N_8944);
or U14080 (N_14080,N_8712,N_9043);
or U14081 (N_14081,N_7601,N_11287);
and U14082 (N_14082,N_6615,N_10604);
or U14083 (N_14083,N_12418,N_6549);
xor U14084 (N_14084,N_12121,N_11946);
or U14085 (N_14085,N_10236,N_10487);
or U14086 (N_14086,N_12474,N_7101);
nand U14087 (N_14087,N_10311,N_6600);
nand U14088 (N_14088,N_6996,N_11312);
nor U14089 (N_14089,N_11443,N_8618);
nand U14090 (N_14090,N_12137,N_8948);
and U14091 (N_14091,N_10993,N_11339);
and U14092 (N_14092,N_8672,N_9552);
xor U14093 (N_14093,N_6303,N_8729);
or U14094 (N_14094,N_10615,N_11517);
and U14095 (N_14095,N_9720,N_11992);
nand U14096 (N_14096,N_12331,N_10216);
xnor U14097 (N_14097,N_9779,N_7083);
nand U14098 (N_14098,N_7768,N_7597);
nand U14099 (N_14099,N_10234,N_11662);
nand U14100 (N_14100,N_7259,N_11110);
or U14101 (N_14101,N_6791,N_6873);
nand U14102 (N_14102,N_7330,N_8617);
xor U14103 (N_14103,N_7669,N_8353);
and U14104 (N_14104,N_6755,N_10140);
or U14105 (N_14105,N_8741,N_12017);
and U14106 (N_14106,N_12408,N_10080);
or U14107 (N_14107,N_6562,N_10931);
xor U14108 (N_14108,N_9036,N_11709);
nor U14109 (N_14109,N_7059,N_11886);
and U14110 (N_14110,N_8604,N_7810);
xnor U14111 (N_14111,N_6775,N_8134);
nand U14112 (N_14112,N_12451,N_7537);
and U14113 (N_14113,N_6524,N_10104);
nor U14114 (N_14114,N_10996,N_11796);
and U14115 (N_14115,N_10654,N_10225);
nor U14116 (N_14116,N_7857,N_10710);
nor U14117 (N_14117,N_10139,N_7552);
or U14118 (N_14118,N_10257,N_10342);
nor U14119 (N_14119,N_7486,N_6979);
xor U14120 (N_14120,N_12271,N_11698);
or U14121 (N_14121,N_10240,N_11536);
and U14122 (N_14122,N_10805,N_12068);
xor U14123 (N_14123,N_11347,N_11779);
xnor U14124 (N_14124,N_8663,N_6832);
xor U14125 (N_14125,N_11111,N_12443);
or U14126 (N_14126,N_10325,N_7366);
nand U14127 (N_14127,N_9933,N_11330);
xnor U14128 (N_14128,N_11528,N_10270);
and U14129 (N_14129,N_11734,N_10176);
and U14130 (N_14130,N_8929,N_6641);
or U14131 (N_14131,N_8578,N_11865);
nor U14132 (N_14132,N_7233,N_9609);
xor U14133 (N_14133,N_12126,N_10495);
nor U14134 (N_14134,N_8524,N_6994);
nand U14135 (N_14135,N_6560,N_8418);
and U14136 (N_14136,N_10315,N_6661);
nand U14137 (N_14137,N_9151,N_12163);
and U14138 (N_14138,N_10073,N_6871);
and U14139 (N_14139,N_6664,N_11916);
nor U14140 (N_14140,N_11957,N_8331);
xnor U14141 (N_14141,N_12118,N_7922);
nand U14142 (N_14142,N_9085,N_10841);
or U14143 (N_14143,N_12488,N_10069);
or U14144 (N_14144,N_8108,N_8380);
xor U14145 (N_14145,N_12420,N_10799);
or U14146 (N_14146,N_11742,N_10371);
xnor U14147 (N_14147,N_10631,N_10029);
nand U14148 (N_14148,N_6425,N_11547);
nand U14149 (N_14149,N_9826,N_7085);
xor U14150 (N_14150,N_9033,N_7862);
nor U14151 (N_14151,N_9863,N_12277);
or U14152 (N_14152,N_10686,N_10014);
or U14153 (N_14153,N_11986,N_8661);
xnor U14154 (N_14154,N_8047,N_11607);
and U14155 (N_14155,N_10304,N_8393);
or U14156 (N_14156,N_12498,N_11481);
or U14157 (N_14157,N_7436,N_6667);
nand U14158 (N_14158,N_6946,N_8061);
or U14159 (N_14159,N_11272,N_9363);
and U14160 (N_14160,N_9438,N_9131);
xor U14161 (N_14161,N_10467,N_9423);
or U14162 (N_14162,N_8470,N_6619);
nor U14163 (N_14163,N_10151,N_8174);
xor U14164 (N_14164,N_6341,N_8302);
xnor U14165 (N_14165,N_8157,N_12222);
nor U14166 (N_14166,N_8364,N_10860);
and U14167 (N_14167,N_6868,N_7655);
or U14168 (N_14168,N_10194,N_7666);
xor U14169 (N_14169,N_8149,N_8148);
or U14170 (N_14170,N_10848,N_8704);
or U14171 (N_14171,N_8307,N_12115);
or U14172 (N_14172,N_10537,N_6447);
or U14173 (N_14173,N_7048,N_11722);
xnor U14174 (N_14174,N_8446,N_12244);
xor U14175 (N_14175,N_10001,N_8399);
or U14176 (N_14176,N_11535,N_9210);
nor U14177 (N_14177,N_12178,N_7334);
or U14178 (N_14178,N_9354,N_11874);
or U14179 (N_14179,N_10247,N_9672);
nand U14180 (N_14180,N_11814,N_8272);
xor U14181 (N_14181,N_9821,N_7027);
or U14182 (N_14182,N_7185,N_9084);
and U14183 (N_14183,N_10566,N_7589);
nand U14184 (N_14184,N_7821,N_10983);
nand U14185 (N_14185,N_9345,N_8811);
xnor U14186 (N_14186,N_9166,N_11309);
and U14187 (N_14187,N_11331,N_11930);
or U14188 (N_14188,N_8319,N_9012);
or U14189 (N_14189,N_10473,N_9300);
xor U14190 (N_14190,N_8092,N_6917);
nor U14191 (N_14191,N_9344,N_11190);
or U14192 (N_14192,N_10980,N_6296);
nor U14193 (N_14193,N_9766,N_6322);
xor U14194 (N_14194,N_7152,N_10778);
xnor U14195 (N_14195,N_10790,N_6604);
or U14196 (N_14196,N_11209,N_11941);
xnor U14197 (N_14197,N_10350,N_6475);
nor U14198 (N_14198,N_8545,N_9534);
xnor U14199 (N_14199,N_9896,N_8883);
nand U14200 (N_14200,N_8505,N_7168);
and U14201 (N_14201,N_12333,N_10933);
xor U14202 (N_14202,N_9189,N_10630);
xnor U14203 (N_14203,N_6941,N_9420);
xnor U14204 (N_14204,N_10091,N_9911);
or U14205 (N_14205,N_6729,N_11642);
and U14206 (N_14206,N_10929,N_8533);
and U14207 (N_14207,N_7959,N_6771);
xnor U14208 (N_14208,N_8924,N_11590);
or U14209 (N_14209,N_10459,N_6555);
nor U14210 (N_14210,N_7081,N_11385);
nor U14211 (N_14211,N_6813,N_9908);
nor U14212 (N_14212,N_7924,N_9232);
nor U14213 (N_14213,N_8577,N_7979);
nor U14214 (N_14214,N_6818,N_8994);
or U14215 (N_14215,N_6342,N_8039);
nor U14216 (N_14216,N_7203,N_7311);
nor U14217 (N_14217,N_8466,N_11516);
nor U14218 (N_14218,N_8532,N_10469);
nor U14219 (N_14219,N_12012,N_7483);
nand U14220 (N_14220,N_11389,N_6756);
xnor U14221 (N_14221,N_8189,N_8850);
xor U14222 (N_14222,N_8768,N_10344);
nand U14223 (N_14223,N_10685,N_7387);
or U14224 (N_14224,N_12297,N_8165);
xor U14225 (N_14225,N_9417,N_6423);
or U14226 (N_14226,N_7122,N_9203);
and U14227 (N_14227,N_10619,N_11164);
nor U14228 (N_14228,N_12050,N_12311);
nand U14229 (N_14229,N_11488,N_10099);
and U14230 (N_14230,N_6843,N_9701);
xor U14231 (N_14231,N_7426,N_11295);
nand U14232 (N_14232,N_11559,N_9747);
nor U14233 (N_14233,N_10356,N_11515);
nor U14234 (N_14234,N_10577,N_7734);
or U14235 (N_14235,N_8441,N_10756);
nand U14236 (N_14236,N_8973,N_7758);
and U14237 (N_14237,N_8659,N_6680);
xnor U14238 (N_14238,N_10693,N_9183);
nor U14239 (N_14239,N_12031,N_7838);
xor U14240 (N_14240,N_6787,N_12316);
nand U14241 (N_14241,N_7504,N_8960);
xor U14242 (N_14242,N_11903,N_7573);
nand U14243 (N_14243,N_9267,N_9740);
and U14244 (N_14244,N_7018,N_10123);
xnor U14245 (N_14245,N_8788,N_8912);
or U14246 (N_14246,N_6638,N_9030);
or U14247 (N_14247,N_10379,N_6389);
nand U14248 (N_14248,N_7465,N_7397);
and U14249 (N_14249,N_8615,N_8581);
xnor U14250 (N_14250,N_7723,N_6944);
nand U14251 (N_14251,N_6609,N_7087);
nor U14252 (N_14252,N_10328,N_11218);
or U14253 (N_14253,N_8007,N_7476);
and U14254 (N_14254,N_7868,N_11617);
nor U14255 (N_14255,N_11477,N_10026);
and U14256 (N_14256,N_10256,N_7146);
or U14257 (N_14257,N_8196,N_8242);
or U14258 (N_14258,N_12388,N_10968);
xnor U14259 (N_14259,N_9639,N_7725);
xnor U14260 (N_14260,N_9424,N_7873);
nand U14261 (N_14261,N_10724,N_10061);
nor U14262 (N_14262,N_10828,N_10622);
and U14263 (N_14263,N_11715,N_11995);
xor U14264 (N_14264,N_7742,N_9275);
or U14265 (N_14265,N_8554,N_11044);
and U14266 (N_14266,N_11391,N_10239);
nand U14267 (N_14267,N_9311,N_7094);
or U14268 (N_14268,N_6514,N_8945);
nor U14269 (N_14269,N_8179,N_8030);
and U14270 (N_14270,N_6835,N_7323);
xnor U14271 (N_14271,N_9695,N_9638);
nor U14272 (N_14272,N_7229,N_7777);
nor U14273 (N_14273,N_9215,N_7891);
or U14274 (N_14274,N_8444,N_7598);
and U14275 (N_14275,N_12462,N_8782);
nand U14276 (N_14276,N_6263,N_6790);
and U14277 (N_14277,N_8309,N_11623);
nand U14278 (N_14278,N_6986,N_11107);
or U14279 (N_14279,N_10134,N_9518);
and U14280 (N_14280,N_8676,N_7477);
or U14281 (N_14281,N_7350,N_11719);
xnor U14282 (N_14282,N_12078,N_6856);
nand U14283 (N_14283,N_10493,N_7284);
nand U14284 (N_14284,N_9511,N_9231);
nand U14285 (N_14285,N_12187,N_9738);
nor U14286 (N_14286,N_9661,N_6469);
nor U14287 (N_14287,N_7948,N_12248);
and U14288 (N_14288,N_6711,N_9089);
xnor U14289 (N_14289,N_10512,N_9040);
or U14290 (N_14290,N_10731,N_9613);
xor U14291 (N_14291,N_8818,N_6801);
and U14292 (N_14292,N_8529,N_8642);
xnor U14293 (N_14293,N_11108,N_9992);
nor U14294 (N_14294,N_12171,N_7774);
xor U14295 (N_14295,N_7049,N_9853);
nand U14296 (N_14296,N_12442,N_8993);
nand U14297 (N_14297,N_8181,N_7750);
and U14298 (N_14298,N_8915,N_11106);
or U14299 (N_14299,N_9796,N_12393);
nor U14300 (N_14300,N_11649,N_11669);
nand U14301 (N_14301,N_9484,N_7411);
nand U14302 (N_14302,N_10813,N_10393);
and U14303 (N_14303,N_9756,N_7312);
and U14304 (N_14304,N_8871,N_12292);
or U14305 (N_14305,N_8265,N_6393);
nor U14306 (N_14306,N_8156,N_12192);
and U14307 (N_14307,N_9550,N_8029);
nor U14308 (N_14308,N_9271,N_11665);
xnor U14309 (N_14309,N_6762,N_8283);
xnor U14310 (N_14310,N_9658,N_10462);
or U14311 (N_14311,N_11599,N_7603);
and U14312 (N_14312,N_11643,N_7326);
and U14313 (N_14313,N_12365,N_6728);
nand U14314 (N_14314,N_6910,N_9680);
and U14315 (N_14315,N_11831,N_9644);
nand U14316 (N_14316,N_10352,N_12032);
nor U14317 (N_14317,N_6597,N_8866);
nand U14318 (N_14318,N_10252,N_6807);
xnor U14319 (N_14319,N_8276,N_12175);
nand U14320 (N_14320,N_12033,N_6984);
or U14321 (N_14321,N_7627,N_9708);
nand U14322 (N_14322,N_8995,N_7475);
or U14323 (N_14323,N_7679,N_9964);
and U14324 (N_14324,N_8514,N_9308);
and U14325 (N_14325,N_8062,N_7620);
and U14326 (N_14326,N_8748,N_12085);
and U14327 (N_14327,N_6400,N_11878);
nor U14328 (N_14328,N_7184,N_11730);
xnor U14329 (N_14329,N_11266,N_10071);
and U14330 (N_14330,N_9707,N_7658);
xor U14331 (N_14331,N_9006,N_7444);
or U14332 (N_14332,N_10184,N_9218);
or U14333 (N_14333,N_11837,N_7524);
or U14334 (N_14334,N_10915,N_9734);
nor U14335 (N_14335,N_8292,N_10211);
xor U14336 (N_14336,N_10922,N_12047);
and U14337 (N_14337,N_10119,N_9282);
and U14338 (N_14338,N_7333,N_7010);
or U14339 (N_14339,N_11683,N_7583);
or U14340 (N_14340,N_11361,N_9859);
xnor U14341 (N_14341,N_12006,N_9053);
or U14342 (N_14342,N_10718,N_10627);
nand U14343 (N_14343,N_9333,N_7548);
xnor U14344 (N_14344,N_8119,N_8350);
and U14345 (N_14345,N_9676,N_7455);
nand U14346 (N_14346,N_6965,N_10267);
and U14347 (N_14347,N_7172,N_7478);
and U14348 (N_14348,N_10370,N_12485);
nor U14349 (N_14349,N_9907,N_7542);
nor U14350 (N_14350,N_10427,N_10732);
or U14351 (N_14351,N_8823,N_8967);
and U14352 (N_14352,N_6437,N_6520);
nor U14353 (N_14353,N_8512,N_7220);
xnor U14354 (N_14354,N_9775,N_9409);
and U14355 (N_14355,N_9093,N_9206);
xnor U14356 (N_14356,N_10264,N_7466);
nand U14357 (N_14357,N_6500,N_9872);
nand U14358 (N_14358,N_12059,N_8899);
nor U14359 (N_14359,N_10858,N_10699);
nand U14360 (N_14360,N_9547,N_8893);
nor U14361 (N_14361,N_10535,N_12097);
and U14362 (N_14362,N_10132,N_10892);
or U14363 (N_14363,N_11289,N_11143);
and U14364 (N_14364,N_12265,N_7945);
or U14365 (N_14365,N_6419,N_9421);
and U14366 (N_14366,N_7695,N_11007);
xor U14367 (N_14367,N_11829,N_6485);
xor U14368 (N_14368,N_9961,N_6754);
or U14369 (N_14369,N_10796,N_11299);
xnor U14370 (N_14370,N_10479,N_8590);
and U14371 (N_14371,N_11635,N_7329);
or U14372 (N_14372,N_8086,N_8675);
nand U14373 (N_14373,N_7026,N_11864);
and U14374 (N_14374,N_6558,N_11925);
xor U14375 (N_14375,N_7753,N_9395);
or U14376 (N_14376,N_8520,N_10250);
xor U14377 (N_14377,N_7017,N_9683);
and U14378 (N_14378,N_9120,N_7160);
nand U14379 (N_14379,N_8625,N_8240);
nor U14380 (N_14380,N_8327,N_7848);
nand U14381 (N_14381,N_10901,N_7246);
nand U14382 (N_14382,N_10378,N_11502);
or U14383 (N_14383,N_12125,N_9083);
nand U14384 (N_14384,N_11303,N_8348);
xnor U14385 (N_14385,N_8744,N_6658);
xnor U14386 (N_14386,N_12101,N_9237);
and U14387 (N_14387,N_9301,N_8531);
xor U14388 (N_14388,N_7818,N_9558);
xnor U14389 (N_14389,N_8471,N_8921);
xor U14390 (N_14390,N_7653,N_10687);
nand U14391 (N_14391,N_11509,N_9468);
and U14392 (N_14392,N_10652,N_6934);
nor U14393 (N_14393,N_10181,N_7496);
nor U14394 (N_14394,N_10585,N_6552);
nor U14395 (N_14395,N_8143,N_8769);
nor U14396 (N_14396,N_7287,N_11254);
or U14397 (N_14397,N_9681,N_6375);
and U14398 (N_14398,N_6950,N_8528);
and U14399 (N_14399,N_9436,N_11271);
and U14400 (N_14400,N_8981,N_8737);
xnor U14401 (N_14401,N_7008,N_8658);
nor U14402 (N_14402,N_9462,N_12483);
nor U14403 (N_14403,N_10148,N_7509);
xor U14404 (N_14404,N_8306,N_6518);
nor U14405 (N_14405,N_7593,N_11051);
or U14406 (N_14406,N_6768,N_7939);
xor U14407 (N_14407,N_11032,N_8853);
nand U14408 (N_14408,N_7158,N_7462);
xor U14409 (N_14409,N_8836,N_7169);
nand U14410 (N_14410,N_9103,N_12113);
xnor U14411 (N_14411,N_12425,N_8802);
or U14412 (N_14412,N_11422,N_8874);
or U14413 (N_14413,N_10276,N_9477);
xor U14414 (N_14414,N_10576,N_10043);
nor U14415 (N_14415,N_9471,N_8299);
or U14416 (N_14416,N_11401,N_8961);
or U14417 (N_14417,N_10046,N_8427);
and U14418 (N_14418,N_11615,N_6830);
xnor U14419 (N_14419,N_9780,N_10759);
and U14420 (N_14420,N_11961,N_7729);
nor U14421 (N_14421,N_11338,N_9430);
and U14422 (N_14422,N_9943,N_8713);
xnor U14423 (N_14423,N_8591,N_10330);
or U14424 (N_14424,N_10279,N_6456);
xor U14425 (N_14425,N_10717,N_11283);
nand U14426 (N_14426,N_7999,N_11352);
or U14427 (N_14427,N_6959,N_9542);
xnor U14428 (N_14428,N_6682,N_11498);
nand U14429 (N_14429,N_8816,N_10454);
nor U14430 (N_14430,N_11735,N_7693);
nor U14431 (N_14431,N_9786,N_10366);
nor U14432 (N_14432,N_9338,N_8954);
nand U14433 (N_14433,N_8543,N_11340);
nand U14434 (N_14434,N_7522,N_10651);
and U14435 (N_14435,N_10667,N_8252);
or U14436 (N_14436,N_10086,N_7672);
nor U14437 (N_14437,N_11192,N_7228);
or U14438 (N_14438,N_8795,N_9398);
nand U14439 (N_14439,N_10609,N_6642);
and U14440 (N_14440,N_8358,N_10052);
xnor U14441 (N_14441,N_10017,N_8055);
or U14442 (N_14442,N_12177,N_9864);
nand U14443 (N_14443,N_12377,N_11769);
or U14444 (N_14444,N_9822,N_11818);
xor U14445 (N_14445,N_8424,N_12473);
nor U14446 (N_14446,N_10004,N_8415);
nand U14447 (N_14447,N_8113,N_7061);
or U14448 (N_14448,N_7433,N_6478);
nand U14449 (N_14449,N_6457,N_11958);
xor U14450 (N_14450,N_12487,N_7262);
xnor U14451 (N_14451,N_8405,N_7224);
or U14452 (N_14452,N_6967,N_12492);
xnor U14453 (N_14453,N_9434,N_12385);
nand U14454 (N_14454,N_11269,N_11445);
and U14455 (N_14455,N_7253,N_8998);
or U14456 (N_14456,N_7880,N_9939);
or U14457 (N_14457,N_8548,N_7033);
xnor U14458 (N_14458,N_7765,N_7786);
or U14459 (N_14459,N_9836,N_12326);
nor U14460 (N_14460,N_8155,N_10653);
xnor U14461 (N_14461,N_10970,N_8172);
or U14462 (N_14462,N_6903,N_11781);
xor U14463 (N_14463,N_12341,N_9124);
xor U14464 (N_14464,N_6745,N_8904);
and U14465 (N_14465,N_9228,N_6613);
and U14466 (N_14466,N_6512,N_12324);
nand U14467 (N_14467,N_8263,N_10861);
nand U14468 (N_14468,N_8635,N_8807);
nor U14469 (N_14469,N_8561,N_7613);
or U14470 (N_14470,N_7689,N_7706);
xor U14471 (N_14471,N_6931,N_10565);
or U14472 (N_14472,N_10715,N_7191);
xnor U14473 (N_14473,N_8132,N_8691);
nor U14474 (N_14474,N_11927,N_9125);
nor U14475 (N_14475,N_11233,N_10126);
nand U14476 (N_14476,N_6594,N_11353);
nor U14477 (N_14477,N_9576,N_6511);
xor U14478 (N_14478,N_6617,N_10324);
nand U14479 (N_14479,N_6324,N_12352);
xor U14480 (N_14480,N_12173,N_12127);
nor U14481 (N_14481,N_11478,N_6458);
nand U14482 (N_14482,N_6367,N_6515);
nand U14483 (N_14483,N_8918,N_7638);
nand U14484 (N_14484,N_7133,N_7694);
nor U14485 (N_14485,N_9951,N_7854);
nor U14486 (N_14486,N_8552,N_12347);
and U14487 (N_14487,N_7892,N_10269);
nor U14488 (N_14488,N_11993,N_7714);
and U14489 (N_14489,N_11963,N_10012);
xnor U14490 (N_14490,N_9522,N_8611);
and U14491 (N_14491,N_9256,N_8488);
and U14492 (N_14492,N_6740,N_11324);
xor U14493 (N_14493,N_10224,N_6780);
nand U14494 (N_14494,N_10222,N_8114);
xnor U14495 (N_14495,N_8026,N_9225);
and U14496 (N_14496,N_7263,N_10021);
or U14497 (N_14497,N_9675,N_10811);
xnor U14498 (N_14498,N_10175,N_9569);
xor U14499 (N_14499,N_11644,N_12447);
xnor U14500 (N_14500,N_6577,N_8636);
and U14501 (N_14501,N_9829,N_7874);
and U14502 (N_14502,N_8939,N_6450);
and U14503 (N_14503,N_11285,N_10088);
xnor U14504 (N_14504,N_8243,N_7021);
nor U14505 (N_14505,N_9070,N_9593);
nor U14506 (N_14506,N_11694,N_10122);
nand U14507 (N_14507,N_12471,N_9496);
nor U14508 (N_14508,N_10242,N_9607);
nor U14509 (N_14509,N_12087,N_11354);
nor U14510 (N_14510,N_8979,N_8632);
or U14511 (N_14511,N_6479,N_11906);
and U14512 (N_14512,N_10195,N_9833);
nor U14513 (N_14513,N_7513,N_6980);
or U14514 (N_14514,N_12185,N_7480);
and U14515 (N_14515,N_10826,N_6289);
nand U14516 (N_14516,N_12392,N_10594);
and U14517 (N_14517,N_10064,N_11096);
and U14518 (N_14518,N_10492,N_9304);
and U14519 (N_14519,N_11851,N_9935);
and U14520 (N_14520,N_12424,N_6254);
nand U14521 (N_14521,N_12084,N_8888);
nand U14522 (N_14522,N_9632,N_6495);
nand U14523 (N_14523,N_11866,N_11589);
xnor U14524 (N_14524,N_12060,N_10013);
nor U14525 (N_14525,N_10468,N_8690);
and U14526 (N_14526,N_12204,N_9702);
xor U14527 (N_14527,N_10188,N_12464);
and U14528 (N_14528,N_9723,N_12305);
and U14529 (N_14529,N_6411,N_11582);
or U14530 (N_14530,N_11349,N_7565);
and U14531 (N_14531,N_9699,N_10646);
xor U14532 (N_14532,N_9718,N_11847);
xor U14533 (N_14533,N_11726,N_6438);
xor U14534 (N_14534,N_9330,N_9532);
and U14535 (N_14535,N_7826,N_11550);
or U14536 (N_14536,N_7633,N_11070);
or U14537 (N_14537,N_11436,N_7065);
or U14538 (N_14538,N_11008,N_10918);
and U14539 (N_14539,N_7976,N_8686);
nor U14540 (N_14540,N_8225,N_7846);
nor U14541 (N_14541,N_10170,N_10503);
and U14542 (N_14542,N_11042,N_6966);
or U14543 (N_14543,N_6343,N_6464);
and U14544 (N_14544,N_11364,N_7579);
or U14545 (N_14545,N_9445,N_11215);
nand U14546 (N_14546,N_11030,N_11297);
xnor U14547 (N_14547,N_8005,N_8076);
nand U14548 (N_14548,N_7793,N_11085);
nor U14549 (N_14549,N_11284,N_9172);
nor U14550 (N_14550,N_8280,N_8067);
xnor U14551 (N_14551,N_7216,N_8786);
and U14552 (N_14552,N_9193,N_7605);
or U14553 (N_14553,N_11806,N_8560);
nor U14554 (N_14554,N_12281,N_10365);
xor U14555 (N_14555,N_6932,N_9194);
or U14556 (N_14556,N_6904,N_10290);
nand U14557 (N_14557,N_10191,N_10045);
and U14558 (N_14558,N_7295,N_10116);
and U14559 (N_14559,N_10791,N_8809);
and U14560 (N_14560,N_10581,N_6981);
xnor U14561 (N_14561,N_10874,N_6497);
nor U14562 (N_14562,N_6340,N_8828);
nand U14563 (N_14563,N_8411,N_8717);
xnor U14564 (N_14564,N_6864,N_10268);
nand U14565 (N_14565,N_11674,N_6476);
nor U14566 (N_14566,N_7443,N_8315);
xnor U14567 (N_14567,N_7580,N_8188);
nand U14568 (N_14568,N_6851,N_6317);
xor U14569 (N_14569,N_12237,N_9368);
nor U14570 (N_14570,N_9372,N_10992);
nand U14571 (N_14571,N_6948,N_7710);
and U14572 (N_14572,N_6426,N_9893);
nor U14573 (N_14573,N_11328,N_11572);
or U14574 (N_14574,N_12348,N_7910);
nand U14575 (N_14575,N_6349,N_7905);
and U14576 (N_14576,N_7132,N_10288);
nor U14577 (N_14577,N_8052,N_6840);
nor U14578 (N_14578,N_10541,N_11744);
or U14579 (N_14579,N_10642,N_12217);
nor U14580 (N_14580,N_8287,N_9563);
nand U14581 (N_14581,N_6848,N_12043);
xor U14582 (N_14582,N_7705,N_11463);
and U14583 (N_14583,N_10572,N_7005);
nand U14584 (N_14584,N_6884,N_6962);
or U14585 (N_14585,N_9180,N_11286);
or U14586 (N_14586,N_11978,N_7367);
xnor U14587 (N_14587,N_7535,N_6850);
nor U14588 (N_14588,N_7159,N_10443);
xnor U14589 (N_14589,N_12140,N_10281);
nand U14590 (N_14590,N_11616,N_6436);
and U14591 (N_14591,N_8230,N_10906);
and U14592 (N_14592,N_11416,N_7795);
nor U14593 (N_14593,N_11292,N_11366);
nor U14594 (N_14594,N_9319,N_10920);
xor U14595 (N_14595,N_7270,N_11146);
xnor U14596 (N_14596,N_9454,N_9397);
or U14597 (N_14597,N_10130,N_11824);
and U14598 (N_14598,N_10212,N_6580);
nand U14599 (N_14599,N_10815,N_8897);
or U14600 (N_14600,N_11761,N_11670);
nor U14601 (N_14601,N_8277,N_8743);
or U14602 (N_14602,N_9526,N_8474);
or U14603 (N_14603,N_9945,N_12156);
xor U14604 (N_14604,N_6482,N_9844);
xor U14605 (N_14605,N_12055,N_9048);
xnor U14606 (N_14606,N_6808,N_10323);
xor U14607 (N_14607,N_11262,N_9315);
nand U14608 (N_14608,N_9007,N_10879);
or U14609 (N_14609,N_9684,N_6744);
or U14610 (N_14610,N_7299,N_11126);
xor U14611 (N_14611,N_9415,N_8413);
nor U14612 (N_14612,N_10614,N_6943);
xnor U14613 (N_14613,N_11068,N_11316);
xor U14614 (N_14614,N_8396,N_9758);
nor U14615 (N_14615,N_8931,N_10035);
nand U14616 (N_14616,N_8705,N_10552);
and U14617 (N_14617,N_7956,N_11685);
nand U14618 (N_14618,N_10494,N_9213);
or U14619 (N_14619,N_6498,N_11379);
xor U14620 (N_14620,N_7698,N_6410);
nor U14621 (N_14621,N_12106,N_6788);
or U14622 (N_14622,N_8190,N_7861);
or U14623 (N_14623,N_10743,N_9042);
nand U14624 (N_14624,N_6432,N_8827);
or U14625 (N_14625,N_9374,N_8310);
xnor U14626 (N_14626,N_8946,N_8136);
xor U14627 (N_14627,N_6855,N_8815);
nand U14628 (N_14628,N_11834,N_6368);
xnor U14629 (N_14629,N_12289,N_8582);
xnor U14630 (N_14630,N_7680,N_10554);
nor U14631 (N_14631,N_11279,N_7718);
nor U14632 (N_14632,N_8609,N_11325);
or U14633 (N_14633,N_9616,N_12414);
or U14634 (N_14634,N_6275,N_11308);
xnor U14635 (N_14635,N_10658,N_7836);
xor U14636 (N_14636,N_7276,N_8476);
nand U14637 (N_14637,N_9586,N_11648);
nor U14638 (N_14638,N_9128,N_12075);
xnor U14639 (N_14639,N_6891,N_6735);
nand U14640 (N_14640,N_9318,N_10000);
or U14641 (N_14641,N_10214,N_7928);
xnor U14642 (N_14642,N_7629,N_12143);
or U14643 (N_14643,N_10461,N_7459);
or U14644 (N_14644,N_9055,N_9337);
nor U14645 (N_14645,N_7728,N_8982);
nand U14646 (N_14646,N_8985,N_10384);
and U14647 (N_14647,N_9764,N_9858);
or U14648 (N_14648,N_8851,N_6723);
and U14649 (N_14649,N_8479,N_11017);
nand U14650 (N_14650,N_8212,N_6911);
xor U14651 (N_14651,N_8638,N_10885);
and U14652 (N_14652,N_6781,N_9865);
or U14653 (N_14653,N_7696,N_6523);
or U14654 (N_14654,N_10792,N_11268);
and U14655 (N_14655,N_8056,N_7585);
or U14656 (N_14656,N_7197,N_9343);
nor U14657 (N_14657,N_7137,N_10056);
xor U14658 (N_14658,N_11894,N_7507);
nor U14659 (N_14659,N_6266,N_10645);
and U14660 (N_14660,N_9177,N_9995);
xnor U14661 (N_14661,N_11696,N_9031);
and U14662 (N_14662,N_10457,N_9942);
or U14663 (N_14663,N_8790,N_10274);
and U14664 (N_14664,N_11756,N_10385);
or U14665 (N_14665,N_10785,N_7114);
xnor U14666 (N_14666,N_8834,N_11494);
and U14667 (N_14667,N_11875,N_10536);
and U14668 (N_14668,N_11503,N_11394);
and U14669 (N_14669,N_10595,N_10660);
and U14670 (N_14670,N_10142,N_7130);
nor U14671 (N_14671,N_8906,N_6536);
and U14672 (N_14672,N_7022,N_10659);
nor U14673 (N_14673,N_8256,N_6327);
xor U14674 (N_14674,N_6443,N_8852);
xor U14675 (N_14675,N_12046,N_10498);
and U14676 (N_14676,N_10349,N_11578);
nand U14677 (N_14677,N_9253,N_8734);
nor U14678 (N_14678,N_9765,N_11252);
or U14679 (N_14679,N_7741,N_8928);
and U14680 (N_14680,N_8953,N_7068);
nand U14681 (N_14681,N_7606,N_9427);
or U14682 (N_14682,N_9546,N_12205);
and U14683 (N_14683,N_7517,N_10359);
or U14684 (N_14684,N_9325,N_9759);
xor U14685 (N_14685,N_10539,N_12354);
nand U14686 (N_14686,N_6676,N_9159);
and U14687 (N_14687,N_9870,N_10900);
or U14688 (N_14688,N_9244,N_8510);
xor U14689 (N_14689,N_7136,N_8362);
and U14690 (N_14690,N_6644,N_9453);
xnor U14691 (N_14691,N_6685,N_10120);
xnor U14692 (N_14692,N_11182,N_8988);
or U14693 (N_14693,N_10238,N_10721);
or U14694 (N_14694,N_11038,N_6545);
or U14695 (N_14695,N_8684,N_10016);
and U14696 (N_14696,N_9751,N_10112);
nor U14697 (N_14697,N_9458,N_8547);
nand U14698 (N_14698,N_10414,N_9002);
xor U14699 (N_14699,N_6633,N_8066);
or U14700 (N_14700,N_8357,N_7877);
nor U14701 (N_14701,N_8760,N_7279);
or U14702 (N_14702,N_10205,N_11797);
xor U14703 (N_14703,N_11228,N_9823);
nand U14704 (N_14704,N_7481,N_8484);
or U14705 (N_14705,N_7757,N_8234);
nor U14706 (N_14706,N_10287,N_7557);
nor U14707 (N_14707,N_9980,N_7450);
or U14708 (N_14708,N_11100,N_9278);
or U14709 (N_14709,N_8595,N_10293);
nand U14710 (N_14710,N_10403,N_10823);
nor U14711 (N_14711,N_8040,N_8669);
and U14712 (N_14712,N_10663,N_9812);
xor U14713 (N_14713,N_7419,N_10636);
nand U14714 (N_14714,N_9176,N_7636);
xnor U14715 (N_14715,N_7571,N_12195);
nor U14716 (N_14716,N_11944,N_11585);
nor U14717 (N_14717,N_8766,N_8621);
nand U14718 (N_14718,N_9240,N_8051);
and U14719 (N_14719,N_7792,N_7766);
and U14720 (N_14720,N_6286,N_6448);
and U14721 (N_14721,N_6253,N_7747);
xnor U14722 (N_14722,N_12048,N_8839);
nand U14723 (N_14723,N_8725,N_10428);
and U14724 (N_14724,N_11521,N_11772);
or U14725 (N_14725,N_10087,N_6316);
nor U14726 (N_14726,N_7327,N_9966);
or U14727 (N_14727,N_11765,N_10505);
and U14728 (N_14728,N_12369,N_9941);
and U14729 (N_14729,N_12019,N_7944);
or U14730 (N_14730,N_9192,N_7347);
and U14731 (N_14731,N_10164,N_10173);
nor U14732 (N_14732,N_6652,N_9144);
and U14733 (N_14733,N_9828,N_9212);
nand U14734 (N_14734,N_11204,N_6785);
and U14735 (N_14735,N_7811,N_6750);
xor U14736 (N_14736,N_8313,N_11081);
xor U14737 (N_14737,N_9061,N_9953);
nand U14738 (N_14738,N_10913,N_8501);
nand U14739 (N_14739,N_7283,N_9105);
nand U14740 (N_14740,N_11015,N_7564);
nand U14741 (N_14741,N_7643,N_10899);
or U14742 (N_14742,N_11166,N_8733);
and U14743 (N_14743,N_12026,N_7200);
nand U14744 (N_14744,N_9247,N_12242);
nand U14745 (N_14745,N_7677,N_8027);
nand U14746 (N_14746,N_10327,N_6614);
and U14747 (N_14747,N_8097,N_8345);
nor U14748 (N_14748,N_8173,N_9881);
nand U14749 (N_14749,N_8845,N_12196);
and U14750 (N_14750,N_11117,N_9072);
or U14751 (N_14751,N_7932,N_11140);
nor U14752 (N_14752,N_12372,N_7437);
nor U14753 (N_14753,N_12067,N_6687);
and U14754 (N_14754,N_7260,N_10424);
or U14755 (N_14755,N_7536,N_8147);
and U14756 (N_14756,N_9580,N_6492);
or U14757 (N_14757,N_8423,N_6491);
xnor U14758 (N_14758,N_8699,N_9654);
xor U14759 (N_14759,N_9052,N_8862);
nand U14760 (N_14760,N_11606,N_10864);
and U14761 (N_14761,N_9847,N_8491);
xor U14762 (N_14762,N_11588,N_7020);
and U14763 (N_14763,N_8135,N_11902);
and U14764 (N_14764,N_7482,N_10700);
or U14765 (N_14765,N_7860,N_7109);
nand U14766 (N_14766,N_11500,N_10749);
or U14767 (N_14767,N_6374,N_9557);
nor U14768 (N_14768,N_6757,N_6396);
or U14769 (N_14769,N_11798,N_8644);
or U14770 (N_14770,N_8320,N_9615);
and U14771 (N_14771,N_9533,N_8015);
xor U14772 (N_14772,N_8660,N_10849);
and U14773 (N_14773,N_7971,N_9217);
or U14774 (N_14774,N_10501,N_12023);
or U14775 (N_14775,N_6525,N_11219);
nor U14776 (N_14776,N_10037,N_7415);
xnor U14777 (N_14777,N_8110,N_12132);
xor U14778 (N_14778,N_10096,N_9467);
nor U14779 (N_14779,N_9287,N_11251);
and U14780 (N_14780,N_10103,N_9355);
or U14781 (N_14781,N_11123,N_9670);
or U14782 (N_14782,N_9998,N_11058);
nor U14783 (N_14783,N_8374,N_9981);
and U14784 (N_14784,N_11860,N_7646);
nand U14785 (N_14785,N_6346,N_7640);
nand U14786 (N_14786,N_11823,N_11752);
and U14787 (N_14787,N_11766,N_9179);
nand U14788 (N_14788,N_7779,N_7994);
or U14789 (N_14789,N_10430,N_8100);
nor U14790 (N_14790,N_11584,N_11789);
nand U14791 (N_14791,N_8096,N_6802);
nor U14792 (N_14792,N_11889,N_7817);
or U14793 (N_14793,N_10423,N_8258);
nor U14794 (N_14794,N_10921,N_9357);
nor U14795 (N_14795,N_9316,N_10697);
nand U14796 (N_14796,N_9922,N_9856);
and U14797 (N_14797,N_9910,N_11105);
xor U14798 (N_14798,N_6998,N_8656);
and U14799 (N_14799,N_10620,N_11676);
or U14800 (N_14800,N_12039,N_9075);
nand U14801 (N_14801,N_11725,N_11247);
nand U14802 (N_14802,N_10932,N_9265);
nand U14803 (N_14803,N_10051,N_8442);
xor U14804 (N_14804,N_8008,N_6413);
or U14805 (N_14805,N_6888,N_8311);
xnor U14806 (N_14806,N_9628,N_6709);
and U14807 (N_14807,N_8102,N_12021);
and U14808 (N_14808,N_11226,N_7652);
and U14809 (N_14809,N_10168,N_6582);
and U14810 (N_14810,N_6696,N_6268);
xor U14811 (N_14811,N_9014,N_8425);
nor U14812 (N_14812,N_9163,N_11438);
nor U14813 (N_14813,N_8262,N_8436);
xor U14814 (N_14814,N_6766,N_11369);
and U14815 (N_14815,N_11001,N_9257);
xor U14816 (N_14816,N_10556,N_11005);
and U14817 (N_14817,N_6528,N_7360);
nand U14818 (N_14818,N_6853,N_9386);
or U14819 (N_14819,N_11220,N_6767);
nand U14820 (N_14820,N_9497,N_6819);
nor U14821 (N_14821,N_7594,N_6689);
or U14822 (N_14822,N_11565,N_8813);
nor U14823 (N_14823,N_6578,N_6332);
nand U14824 (N_14824,N_9119,N_9867);
or U14825 (N_14825,N_8397,N_11206);
and U14826 (N_14826,N_10193,N_6939);
nand U14827 (N_14827,N_9703,N_9482);
xor U14828 (N_14828,N_6953,N_9735);
nand U14829 (N_14829,N_8151,N_7088);
xnor U14830 (N_14830,N_8800,N_12219);
xor U14831 (N_14831,N_7257,N_10127);
or U14832 (N_14832,N_8222,N_11934);
or U14833 (N_14833,N_10387,N_10804);
and U14834 (N_14834,N_11259,N_10322);
xnor U14835 (N_14835,N_7663,N_8587);
nor U14836 (N_14836,N_10794,N_6803);
and U14837 (N_14837,N_6847,N_11811);
nor U14838 (N_14838,N_7012,N_6361);
nand U14839 (N_14839,N_11513,N_6586);
nand U14840 (N_14840,N_11677,N_7751);
and U14841 (N_14841,N_7345,N_7767);
nand U14842 (N_14842,N_8515,N_10230);
nand U14843 (N_14843,N_9455,N_11404);
nor U14844 (N_14844,N_7687,N_9000);
or U14845 (N_14845,N_7966,N_9917);
or U14846 (N_14846,N_7349,N_9495);
and U14847 (N_14847,N_7092,N_10908);
or U14848 (N_14848,N_10397,N_11945);
nand U14849 (N_14849,N_6991,N_10351);
and U14850 (N_14850,N_8544,N_10227);
nand U14851 (N_14851,N_11580,N_11496);
and U14852 (N_14852,N_8846,N_10629);
nor U14853 (N_14853,N_9230,N_11533);
nand U14854 (N_14854,N_6977,N_8003);
nand U14855 (N_14855,N_10803,N_10019);
and U14856 (N_14856,N_9551,N_6691);
or U14857 (N_14857,N_11611,N_12276);
or U14858 (N_14858,N_8194,N_11178);
xor U14859 (N_14859,N_8305,N_11456);
xor U14860 (N_14860,N_9618,N_6828);
xnor U14861 (N_14861,N_7119,N_6576);
or U14862 (N_14862,N_6487,N_6701);
or U14863 (N_14863,N_8036,N_9336);
or U14864 (N_14864,N_7381,N_7828);
nor U14865 (N_14865,N_10489,N_10258);
and U14866 (N_14866,N_8889,N_11828);
xor U14867 (N_14867,N_8316,N_7581);
or U14868 (N_14868,N_11486,N_6672);
or U14869 (N_14869,N_8521,N_6678);
nand U14870 (N_14870,N_9186,N_7918);
or U14871 (N_14871,N_9078,N_10665);
nor U14872 (N_14872,N_9692,N_7941);
or U14873 (N_14873,N_8879,N_6746);
and U14874 (N_14874,N_7775,N_8111);
or U14875 (N_14875,N_6269,N_10764);
and U14876 (N_14876,N_11059,N_7799);
nor U14877 (N_14877,N_10943,N_8329);
and U14878 (N_14878,N_8992,N_8772);
nand U14879 (N_14879,N_8195,N_8969);
xnor U14880 (N_14880,N_6863,N_11815);
nor U14881 (N_14881,N_11932,N_8079);
and U14882 (N_14882,N_9365,N_11293);
nand U14883 (N_14883,N_10518,N_10507);
and U14884 (N_14884,N_8910,N_7722);
nand U14885 (N_14885,N_10335,N_6603);
xor U14886 (N_14886,N_9142,N_10316);
or U14887 (N_14887,N_7563,N_7938);
nor U14888 (N_14888,N_8546,N_12202);
nor U14889 (N_14889,N_6852,N_6490);
nand U14890 (N_14890,N_8654,N_9426);
nor U14891 (N_14891,N_11546,N_7236);
xnor U14892 (N_14892,N_8288,N_10294);
or U14893 (N_14893,N_8458,N_8940);
xor U14894 (N_14894,N_7553,N_7511);
nand U14895 (N_14895,N_11613,N_8032);
and U14896 (N_14896,N_10896,N_11227);
nor U14897 (N_14897,N_6933,N_11522);
and U14898 (N_14898,N_9233,N_10884);
nand U14899 (N_14899,N_7112,N_9553);
xnor U14900 (N_14900,N_9771,N_11511);
or U14901 (N_14901,N_12494,N_7226);
nor U14902 (N_14902,N_7314,N_7139);
xor U14903 (N_14903,N_6968,N_10341);
and U14904 (N_14904,N_6304,N_12174);
and U14905 (N_14905,N_7393,N_7362);
xnor U14906 (N_14906,N_7369,N_9916);
and U14907 (N_14907,N_10499,N_7298);
or U14908 (N_14908,N_6406,N_12339);
nand U14909 (N_14909,N_10244,N_9294);
nand U14910 (N_14910,N_9960,N_7550);
or U14911 (N_14911,N_9774,N_11082);
nor U14912 (N_14912,N_10640,N_9466);
and U14913 (N_14913,N_7179,N_6377);
and U14914 (N_14914,N_9121,N_8694);
or U14915 (N_14915,N_7919,N_11850);
xor U14916 (N_14916,N_8129,N_9272);
or U14917 (N_14917,N_9245,N_6453);
nor U14918 (N_14918,N_10206,N_10217);
nor U14919 (N_14919,N_7099,N_8373);
nand U14920 (N_14920,N_7755,N_10409);
or U14921 (N_14921,N_10486,N_12003);
nor U14922 (N_14922,N_9608,N_7769);
and U14923 (N_14923,N_10145,N_7175);
or U14924 (N_14924,N_7313,N_10821);
nand U14925 (N_14925,N_11920,N_9805);
and U14926 (N_14926,N_6299,N_11880);
and U14927 (N_14927,N_9064,N_10562);
or U14928 (N_14928,N_9361,N_9250);
nor U14929 (N_14929,N_12318,N_9111);
or U14930 (N_14930,N_11120,N_8273);
or U14931 (N_14931,N_11888,N_7641);
xor U14932 (N_14932,N_10872,N_8506);
xor U14933 (N_14933,N_10862,N_6759);
nand U14934 (N_14934,N_6362,N_6290);
xnor U14935 (N_14935,N_10810,N_8235);
xnor U14936 (N_14936,N_9770,N_7461);
xor U14937 (N_14937,N_8417,N_6541);
nand U14938 (N_14938,N_10712,N_11304);
or U14939 (N_14939,N_10613,N_12300);
or U14940 (N_14940,N_10232,N_11686);
or U14941 (N_14941,N_11205,N_9323);
xor U14942 (N_14942,N_8935,N_9685);
nor U14943 (N_14943,N_10568,N_8141);
nor U14944 (N_14944,N_6454,N_10888);
nor U14945 (N_14945,N_7735,N_9885);
and U14946 (N_14946,N_8583,N_6870);
and U14947 (N_14947,N_11854,N_12264);
nor U14948 (N_14948,N_8463,N_10449);
nor U14949 (N_14949,N_7783,N_9816);
and U14950 (N_14950,N_7047,N_7709);
nand U14951 (N_14951,N_8361,N_8431);
nand U14952 (N_14952,N_6251,N_9809);
xor U14953 (N_14953,N_6258,N_7856);
nor U14954 (N_14954,N_7772,N_8991);
nor U14955 (N_14955,N_8167,N_8489);
xor U14956 (N_14956,N_9407,N_12345);
xnor U14957 (N_14957,N_6679,N_6722);
nor U14958 (N_14958,N_7726,N_11402);
nor U14959 (N_14959,N_11605,N_10477);
nor U14960 (N_14960,N_8911,N_9564);
nand U14961 (N_14961,N_9259,N_7123);
xor U14962 (N_14962,N_6815,N_11465);
or U14963 (N_14963,N_11967,N_8950);
or U14964 (N_14964,N_7852,N_9489);
or U14965 (N_14965,N_9688,N_11155);
or U14966 (N_14966,N_6961,N_11356);
and U14967 (N_14967,N_9926,N_12139);
xor U14968 (N_14968,N_12394,N_11076);
nor U14969 (N_14969,N_10589,N_7281);
nand U14970 (N_14970,N_11407,N_11895);
nor U14971 (N_14971,N_10579,N_8133);
xor U14972 (N_14972,N_12298,N_9556);
and U14973 (N_14973,N_7207,N_7904);
xor U14974 (N_14974,N_7684,N_10113);
xor U14975 (N_14975,N_6725,N_7108);
nor U14976 (N_14976,N_7177,N_10545);
xnor U14977 (N_14977,N_11788,N_7244);
and U14978 (N_14978,N_6420,N_10664);
and U14979 (N_14979,N_12226,N_9067);
nor U14980 (N_14980,N_10465,N_11386);
and U14981 (N_14981,N_11839,N_12332);
or U14982 (N_14982,N_7096,N_8050);
nand U14983 (N_14983,N_11221,N_11905);
and U14984 (N_14984,N_9940,N_9874);
nor U14985 (N_14985,N_6494,N_9201);
xor U14986 (N_14986,N_10709,N_10633);
or U14987 (N_14987,N_11253,N_6783);
nor U14988 (N_14988,N_7569,N_9677);
nor U14989 (N_14989,N_9181,N_12198);
or U14990 (N_14990,N_11639,N_6301);
xnor U14991 (N_14991,N_11989,N_8291);
nor U14992 (N_14992,N_8539,N_11191);
xor U14993 (N_14993,N_12203,N_6714);
nand U14994 (N_14994,N_10429,N_11621);
xor U14995 (N_14995,N_10729,N_12020);
nand U14996 (N_14996,N_6640,N_7526);
and U14997 (N_14997,N_7294,N_8687);
or U14998 (N_14998,N_8001,N_9919);
xnor U14999 (N_14999,N_8847,N_7872);
or U15000 (N_15000,N_8084,N_6493);
and U15001 (N_15001,N_11181,N_8207);
nor U15002 (N_15002,N_12434,N_10143);
xor U15003 (N_15003,N_12251,N_10360);
nor U15004 (N_15004,N_6466,N_7110);
nand U15005 (N_15005,N_11413,N_10871);
nor U15006 (N_15006,N_7485,N_9742);
or U15007 (N_15007,N_7290,N_9332);
nor U15008 (N_15008,N_9376,N_10668);
xor U15009 (N_15009,N_11290,N_9326);
xnor U15010 (N_15010,N_7385,N_8959);
and U15011 (N_15011,N_8059,N_9019);
and U15012 (N_15012,N_7576,N_12469);
and U15013 (N_15013,N_9561,N_7804);
nor U15014 (N_15014,N_10978,N_10415);
or U15015 (N_15015,N_10531,N_6666);
xnor U15016 (N_15016,N_8696,N_7351);
nand U15017 (N_15017,N_10802,N_9958);
nand U15018 (N_15018,N_12153,N_10588);
and U15019 (N_15019,N_9165,N_9730);
nor U15020 (N_15020,N_10219,N_6827);
or U15021 (N_15021,N_8498,N_11492);
nor U15022 (N_15022,N_9732,N_7104);
or U15023 (N_15023,N_7321,N_7072);
nor U15024 (N_15024,N_6271,N_9955);
xor U15025 (N_15025,N_9329,N_9924);
and U15026 (N_15026,N_10598,N_6978);
nor U15027 (N_15027,N_10167,N_8614);
or U15028 (N_15028,N_9433,N_8664);
nor U15029 (N_15029,N_7529,N_10574);
nand U15030 (N_15030,N_8900,N_9851);
and U15031 (N_15031,N_7518,N_11936);
xnor U15032 (N_15032,N_7127,N_10475);
nand U15033 (N_15033,N_6905,N_10940);
nand U15034 (N_15034,N_7815,N_6401);
and U15035 (N_15035,N_9492,N_10770);
or U15036 (N_15036,N_10706,N_11310);
or U15037 (N_15037,N_6773,N_6632);
xor U15038 (N_15038,N_9996,N_7674);
or U15039 (N_15039,N_10308,N_10526);
and U15040 (N_15040,N_8682,N_11910);
and U15041 (N_15041,N_11241,N_11016);
and U15042 (N_15042,N_11879,N_11962);
xor U15043 (N_15043,N_9516,N_11770);
nor U15044 (N_15044,N_6417,N_9665);
nand U15045 (N_15045,N_6730,N_9641);
nand U15046 (N_15046,N_10761,N_7822);
or U15047 (N_15047,N_9255,N_6297);
and U15048 (N_15048,N_10987,N_10766);
or U15049 (N_15049,N_7921,N_7273);
or U15050 (N_15050,N_11374,N_11632);
and U15051 (N_15051,N_8941,N_8575);
xnor U15052 (N_15052,N_9902,N_7439);
or U15053 (N_15053,N_7807,N_11675);
xor U15054 (N_15054,N_12285,N_9410);
or U15055 (N_15055,N_8530,N_11647);
nand U15056 (N_15056,N_7178,N_11003);
nand U15057 (N_15057,N_12336,N_7901);
nand U15058 (N_15058,N_10634,N_8673);
xor U15059 (N_15059,N_11158,N_9626);
xnor U15060 (N_15060,N_10814,N_9728);
or U15061 (N_15061,N_6481,N_7702);
and U15062 (N_15062,N_10878,N_8121);
and U15063 (N_15063,N_7957,N_7635);
xnor U15064 (N_15064,N_7866,N_10772);
nand U15065 (N_15065,N_12428,N_8796);
nand U15066 (N_15066,N_6561,N_7056);
nand U15067 (N_15067,N_6628,N_10784);
and U15068 (N_15068,N_8249,N_8685);
and U15069 (N_15069,N_10067,N_8555);
xor U15070 (N_15070,N_12136,N_9778);
or U15071 (N_15071,N_9156,N_6626);
nand U15072 (N_15072,N_6507,N_11541);
nor U15073 (N_15073,N_10050,N_7356);
or U15074 (N_15074,N_9226,N_8773);
xnor U15075 (N_15075,N_6430,N_6405);
nor U15076 (N_15076,N_7121,N_7745);
nor U15077 (N_15077,N_9112,N_8570);
and U15078 (N_15078,N_6307,N_7614);
and U15079 (N_15079,N_7625,N_9385);
or U15080 (N_15080,N_10681,N_12212);
or U15081 (N_15081,N_9088,N_10474);
xnor U15082 (N_15082,N_10146,N_10382);
xor U15083 (N_15083,N_9903,N_10698);
nor U15084 (N_15084,N_10008,N_9577);
xnor U15085 (N_15085,N_9375,N_6260);
xnor U15086 (N_15086,N_9554,N_6471);
nand U15087 (N_15087,N_7845,N_6763);
nand U15088 (N_15088,N_7256,N_11122);
nand U15089 (N_15089,N_6496,N_8118);
nor U15090 (N_15090,N_6842,N_11996);
or U15091 (N_15091,N_11973,N_6902);
nor U15092 (N_15092,N_9523,N_10202);
nor U15093 (N_15093,N_6715,N_10951);
or U15094 (N_15094,N_7052,N_8414);
xor U15095 (N_15095,N_10708,N_11908);
or U15096 (N_15096,N_10683,N_11795);
nand U15097 (N_15097,N_6264,N_9399);
nor U15098 (N_15098,N_9236,N_12077);
xnor U15099 (N_15099,N_9855,N_8640);
nand U15100 (N_15100,N_10975,N_7682);
nand U15101 (N_15101,N_11586,N_8021);
and U15102 (N_15102,N_10907,N_7456);
nor U15103 (N_15103,N_6929,N_11900);
or U15104 (N_15104,N_6351,N_12239);
nand U15105 (N_15105,N_11479,N_11365);
nor U15106 (N_15106,N_7541,N_11768);
or U15107 (N_15107,N_8300,N_7871);
and U15108 (N_15108,N_8089,N_12138);
xnor U15109 (N_15109,N_11461,N_8504);
xor U15110 (N_15110,N_7549,N_6446);
xnor U15111 (N_15111,N_11548,N_10897);
nand U15112 (N_15112,N_7355,N_8325);
xnor U15113 (N_15113,N_11411,N_9171);
and U15114 (N_15114,N_9449,N_6461);
and U15115 (N_15115,N_9290,N_12167);
nor U15116 (N_15116,N_7678,N_7789);
nand U15117 (N_15117,N_6302,N_10295);
or U15118 (N_15118,N_9351,N_8219);
xor U15119 (N_15119,N_7288,N_10852);
xor U15120 (N_15120,N_9832,N_11109);
or U15121 (N_15121,N_9757,N_6880);
and U15122 (N_15122,N_11836,N_7539);
xor U15123 (N_15123,N_8920,N_8647);
xor U15124 (N_15124,N_8481,N_12358);
nand U15125 (N_15125,N_10632,N_6280);
or U15126 (N_15126,N_9348,N_8537);
nor U15127 (N_15127,N_9928,N_8657);
and U15128 (N_15128,N_7558,N_11663);
nand U15129 (N_15129,N_10582,N_7111);
nor U15130 (N_15130,N_10905,N_7469);
nand U15131 (N_15131,N_7338,N_9099);
nand U15132 (N_15132,N_11952,N_12180);
or U15133 (N_15133,N_9716,N_9690);
nand U15134 (N_15134,N_10741,N_6519);
nand U15135 (N_15135,N_12076,N_8384);
or U15136 (N_15136,N_9934,N_12268);
nand U15137 (N_15137,N_11196,N_6348);
xnor U15138 (N_15138,N_7665,N_8177);
and U15139 (N_15139,N_11893,N_10752);
xnor U15140 (N_15140,N_9884,N_9848);
and U15141 (N_15141,N_6665,N_8678);
xor U15142 (N_15142,N_9795,N_8841);
or U15143 (N_15143,N_9448,N_11571);
or U15144 (N_15144,N_11975,N_7306);
or U15145 (N_15145,N_9990,N_9715);
nor U15146 (N_15146,N_8804,N_11690);
nor U15147 (N_15147,N_10419,N_8755);
and U15148 (N_15148,N_6705,N_10455);
nor U15149 (N_15149,N_11751,N_6526);
nor U15150 (N_15150,N_7831,N_10994);
nor U15151 (N_15151,N_9572,N_11321);
nand U15152 (N_15152,N_11384,N_7488);
xnor U15153 (N_15153,N_10831,N_10596);
nand U15154 (N_15154,N_10065,N_6291);
and U15155 (N_15155,N_11388,N_7637);
or U15156 (N_15156,N_7618,N_9525);
and U15157 (N_15157,N_9377,N_7907);
or U15158 (N_15158,N_8936,N_6543);
xnor U15159 (N_15159,N_7615,N_6364);
nor U15160 (N_15160,N_7134,N_9794);
and U15161 (N_15161,N_6416,N_10782);
xnor U15162 (N_15162,N_10930,N_11116);
and U15163 (N_15163,N_8572,N_8344);
xnor U15164 (N_15164,N_6660,N_12157);
nor U15165 (N_15165,N_9428,N_10584);
nor U15166 (N_15166,N_8892,N_8024);
and U15167 (N_15167,N_10196,N_9997);
xnor U15168 (N_15168,N_11311,N_10383);
xnor U15169 (N_15169,N_9241,N_7737);
and U15170 (N_15170,N_9539,N_10283);
and U15171 (N_15171,N_11525,N_9514);
or U15172 (N_15172,N_9838,N_7812);
xor U15173 (N_15173,N_8812,N_6504);
nand U15174 (N_15174,N_6596,N_10160);
xnor U15175 (N_15175,N_9895,N_6388);
xnor U15176 (N_15176,N_8876,N_10695);
or U15177 (N_15177,N_9537,N_11939);
and U15178 (N_15178,N_9209,N_11428);
nor U15179 (N_15179,N_11235,N_11031);
and U15180 (N_15180,N_9854,N_12233);
nand U15181 (N_15181,N_7410,N_12116);
nor U15182 (N_15182,N_7974,N_7390);
or U15183 (N_15183,N_6897,N_11791);
nor U15184 (N_15184,N_9640,N_8557);
or U15185 (N_15185,N_11856,N_10406);
or U15186 (N_15186,N_10504,N_10934);
xor U15187 (N_15187,N_8245,N_7045);
xor U15188 (N_15188,N_8370,N_11583);
xor U15189 (N_15189,N_10082,N_8808);
or U15190 (N_15190,N_11561,N_7064);
or U15191 (N_15191,N_10949,N_12360);
nand U15192 (N_15192,N_9883,N_11552);
or U15193 (N_15193,N_11177,N_9711);
nand U15194 (N_15194,N_8072,N_9106);
nand U15195 (N_15195,N_10720,N_7686);
nor U15196 (N_15196,N_11315,N_9216);
or U15197 (N_15197,N_12279,N_12380);
xor U15198 (N_15198,N_8261,N_7194);
nor U15199 (N_15199,N_9731,N_11852);
and U15200 (N_15200,N_8290,N_10781);
nor U15201 (N_15201,N_9840,N_10515);
and U15202 (N_15202,N_6610,N_7503);
and U15203 (N_15203,N_7173,N_6949);
xnor U15204 (N_15204,N_7380,N_11167);
nand U15205 (N_15205,N_8016,N_10969);
nand U15206 (N_15206,N_7000,N_11890);
xor U15207 (N_15207,N_11118,N_9999);
xor U15208 (N_15208,N_9314,N_9627);
and U15209 (N_15209,N_9023,N_6274);
nor U15210 (N_15210,N_10758,N_9755);
xor U15211 (N_15211,N_11278,N_7050);
nor U15212 (N_15212,N_11186,N_12230);
xnor U15213 (N_15213,N_7157,N_11563);
or U15214 (N_15214,N_10110,N_9871);
nand U15215 (N_15215,N_8624,N_7069);
xor U15216 (N_15216,N_8035,N_9876);
xor U15217 (N_15217,N_9717,N_7955);
or U15218 (N_15218,N_10376,N_8895);
or U15219 (N_15219,N_6622,N_11301);
xor U15220 (N_15220,N_11439,N_6919);
nand U15221 (N_15221,N_12035,N_8435);
and U15222 (N_15222,N_9038,N_10361);
and U15223 (N_15223,N_9753,N_7492);
nand U15224 (N_15224,N_7912,N_12328);
xnor U15225 (N_15225,N_6653,N_12166);
nand U15226 (N_15226,N_10768,N_12267);
and U15227 (N_15227,N_10597,N_11367);
nor U15228 (N_15228,N_7126,N_10231);
nor U15229 (N_15229,N_8600,N_10519);
or U15230 (N_15230,N_7105,N_12246);
nand U15231 (N_15231,N_6901,N_10822);
nand U15232 (N_15232,N_8592,N_9303);
or U15233 (N_15233,N_8185,N_9651);
nand U15234 (N_15234,N_8297,N_9619);
nor U15235 (N_15235,N_7595,N_10169);
and U15236 (N_15236,N_9199,N_9086);
nor U15237 (N_15237,N_7206,N_7391);
nor U15238 (N_15238,N_12240,N_11265);
nor U15239 (N_15239,N_9634,N_12252);
nand U15240 (N_15240,N_10950,N_8416);
and U15241 (N_15241,N_9583,N_8386);
or U15242 (N_15242,N_7566,N_9749);
xnor U15243 (N_15243,N_9251,N_10358);
or U15244 (N_15244,N_9160,N_12463);
nor U15245 (N_15245,N_7446,N_8576);
and U15246 (N_15246,N_10612,N_10049);
nor U15247 (N_15247,N_8403,N_10898);
xnor U15248 (N_15248,N_6974,N_6865);
nor U15249 (N_15249,N_11114,N_10177);
and U15250 (N_15250,N_10744,N_12397);
nor U15251 (N_15251,N_10434,N_10039);
xor U15252 (N_15252,N_9694,N_7060);
xnor U15253 (N_15253,N_9435,N_7039);
or U15254 (N_15254,N_11883,N_6748);
nand U15255 (N_15255,N_11745,N_12477);
nor U15256 (N_15256,N_8756,N_8965);
xor U15257 (N_15257,N_9293,N_12099);
nand U15258 (N_15258,N_10997,N_10197);
nor U15259 (N_15259,N_12315,N_8857);
xor U15260 (N_15260,N_6279,N_7850);
xnor U15261 (N_15261,N_8410,N_10063);
nand U15262 (N_15262,N_11877,N_7659);
or U15263 (N_15263,N_6886,N_6650);
xor U15264 (N_15264,N_12128,N_9952);
and U15265 (N_15265,N_12355,N_10800);
and U15266 (N_15266,N_6538,N_8377);
or U15267 (N_15267,N_10925,N_10886);
xnor U15268 (N_15268,N_10956,N_9195);
and U15269 (N_15269,N_10714,N_9246);
nand U15270 (N_15270,N_11706,N_12435);
or U15271 (N_15271,N_9396,N_7973);
or U15272 (N_15272,N_9839,N_8610);
or U15273 (N_15273,N_9535,N_9222);
or U15274 (N_15274,N_7834,N_11948);
and U15275 (N_15275,N_10753,N_10903);
nand U15276 (N_15276,N_6452,N_7249);
or U15277 (N_15277,N_9669,N_9034);
xor U15278 (N_15278,N_10125,N_6987);
nor U15279 (N_15279,N_11194,N_12232);
xor U15280 (N_15280,N_7370,N_6789);
or U15281 (N_15281,N_9441,N_11680);
nand U15282 (N_15282,N_9659,N_7193);
and U15283 (N_15283,N_11671,N_9897);
nor U15284 (N_15284,N_10692,N_6358);
or U15285 (N_15285,N_7572,N_11230);
nand U15286 (N_15286,N_11346,N_7923);
nor U15287 (N_15287,N_8525,N_7577);
nand U15288 (N_15288,N_7089,N_10599);
nor U15289 (N_15289,N_11333,N_8071);
and U15290 (N_15290,N_8107,N_11964);
or U15291 (N_15291,N_8289,N_12253);
nand U15292 (N_15292,N_11412,N_8775);
nand U15293 (N_15293,N_7699,N_7316);
nor U15294 (N_15294,N_7978,N_6993);
nor U15295 (N_15295,N_11827,N_11844);
nand U15296 (N_15296,N_9527,N_10952);
xnor U15297 (N_15297,N_9378,N_7950);
or U15298 (N_15298,N_6328,N_9108);
or U15299 (N_15299,N_8798,N_11248);
nand U15300 (N_15300,N_7624,N_8558);
and U15301 (N_15301,N_11881,N_8976);
nand U15302 (N_15302,N_7304,N_11610);
or U15303 (N_15303,N_6899,N_8727);
nor U15304 (N_15304,N_10388,N_7497);
nand U15305 (N_15305,N_11102,N_11633);
nand U15306 (N_15306,N_11462,N_7970);
or U15307 (N_15307,N_8926,N_12433);
nand U15308 (N_15308,N_7365,N_10819);
or U15309 (N_15309,N_6751,N_8443);
nand U15310 (N_15310,N_11267,N_7275);
nand U15311 (N_15311,N_10402,N_6428);
xor U15312 (N_15312,N_7785,N_7379);
nor U15313 (N_15313,N_11162,N_7703);
nor U15314 (N_15314,N_9494,N_10343);
nor U15315 (N_15315,N_7610,N_8597);
or U15316 (N_15316,N_8908,N_12066);
or U15317 (N_15317,N_7898,N_8372);
or U15318 (N_15318,N_7732,N_11433);
or U15319 (N_15319,N_9219,N_8706);
or U15320 (N_15320,N_10251,N_7165);
nand U15321 (N_15321,N_8407,N_8598);
xnor U15322 (N_15322,N_10995,N_6444);
nand U15323 (N_15323,N_7523,N_10617);
or U15324 (N_15324,N_7006,N_12044);
nand U15325 (N_15325,N_8623,N_7209);
and U15326 (N_15326,N_7604,N_8098);
xnor U15327 (N_15327,N_9745,N_6353);
nand U15328 (N_15328,N_6601,N_7731);
nand U15329 (N_15329,N_9979,N_7166);
nor U15330 (N_15330,N_8269,N_10702);
or U15331 (N_15331,N_11812,N_10081);
and U15332 (N_15332,N_11819,N_10648);
nand U15333 (N_15333,N_6718,N_10854);
and U15334 (N_15334,N_8805,N_11041);
xnor U15335 (N_15335,N_6983,N_11566);
and U15336 (N_15336,N_10372,N_12274);
and U15337 (N_15337,N_12389,N_7358);
nor U15338 (N_15338,N_7590,N_11277);
nor U15339 (N_15339,N_12427,N_8840);
or U15340 (N_15340,N_9196,N_12449);
xnor U15341 (N_15341,N_7934,N_10437);
nand U15342 (N_15342,N_11972,N_6908);
nand U15343 (N_15343,N_9687,N_12129);
and U15344 (N_15344,N_7028,N_12340);
nor U15345 (N_15345,N_10558,N_12395);
nor U15346 (N_15346,N_12426,N_7591);
xnor U15347 (N_15347,N_11476,N_9113);
nand U15348 (N_15348,N_9977,N_11458);
xnor U15349 (N_15349,N_12093,N_7383);
nor U15350 (N_15350,N_7882,N_11909);
or U15351 (N_15351,N_7309,N_7375);
nand U15352 (N_15352,N_8053,N_9905);
or U15353 (N_15353,N_6913,N_11667);
nand U15354 (N_15354,N_8956,N_9297);
and U15355 (N_15355,N_12415,N_9578);
and U15356 (N_15356,N_12223,N_8522);
nand U15357 (N_15357,N_11380,N_10186);
xor U15358 (N_15358,N_7533,N_9001);
or U15359 (N_15359,N_11211,N_11066);
and U15360 (N_15360,N_7642,N_10959);
or U15361 (N_15361,N_7289,N_11841);
nand U15362 (N_15362,N_7645,N_11091);
nand U15363 (N_15363,N_8332,N_10111);
nor U15364 (N_15364,N_11094,N_11524);
or U15365 (N_15365,N_8404,N_11981);
nor U15366 (N_15366,N_12436,N_8736);
or U15367 (N_15367,N_9153,N_9528);
xor U15368 (N_15368,N_8894,N_7983);
nand U15369 (N_15369,N_11129,N_11776);
xnor U15370 (N_15370,N_12261,N_6330);
and U15371 (N_15371,N_8746,N_11645);
or U15372 (N_15372,N_8378,N_7248);
nand U15373 (N_15373,N_11695,N_7250);
or U15374 (N_15374,N_7073,N_10769);
xor U15375 (N_15375,N_11046,N_8716);
and U15376 (N_15376,N_9238,N_10271);
xor U15377 (N_15377,N_8787,N_6585);
nand U15378 (N_15378,N_12028,N_10833);
xnor U15379 (N_15379,N_10389,N_8260);
xor U15380 (N_15380,N_8054,N_7376);
or U15381 (N_15381,N_12000,N_9077);
or U15382 (N_15382,N_7300,N_7230);
nor U15383 (N_15383,N_11508,N_11083);
nand U15384 (N_15384,N_7717,N_10703);
xnor U15385 (N_15385,N_8594,N_10520);
nand U15386 (N_15386,N_9773,N_6252);
xor U15387 (N_15387,N_7528,N_9380);
xnor U15388 (N_15388,N_8720,N_7046);
or U15389 (N_15389,N_10513,N_7025);
nor U15390 (N_15390,N_9389,N_11857);
nand U15391 (N_15391,N_8523,N_6674);
and U15392 (N_15392,N_7849,N_11222);
and U15393 (N_15393,N_6823,N_9645);
nor U15394 (N_15394,N_10150,N_11898);
or U15395 (N_15395,N_7681,N_10114);
nor U15396 (N_15396,N_12306,N_12308);
or U15397 (N_15397,N_8214,N_9888);
nor U15398 (N_15398,N_7310,N_9689);
and U15399 (N_15399,N_6350,N_7888);
xor U15400 (N_15400,N_10201,N_6442);
nor U15401 (N_15401,N_12416,N_11410);
and U15402 (N_15402,N_10333,N_7051);
and U15403 (N_15403,N_9046,N_12005);
nand U15404 (N_15404,N_7429,N_8355);
nand U15405 (N_15405,N_9592,N_6879);
or U15406 (N_15406,N_11056,N_8964);
nor U15407 (N_15407,N_7673,N_6662);
or U15408 (N_15408,N_6627,N_8205);
or U15409 (N_15409,N_7630,N_11728);
nand U15410 (N_15410,N_8412,N_8781);
nor U15411 (N_15411,N_9503,N_12034);
or U15412 (N_15412,N_6747,N_10623);
nor U15413 (N_15413,N_6315,N_7829);
and U15414 (N_15414,N_10153,N_10204);
or U15415 (N_15415,N_10985,N_10314);
or U15416 (N_15416,N_7128,N_7149);
nand U15417 (N_15417,N_10079,N_9772);
and U15418 (N_15418,N_10210,N_11342);
or U15419 (N_15419,N_9310,N_8301);
or U15420 (N_15420,N_6814,N_11450);
and U15421 (N_15421,N_8259,N_6930);
nor U15422 (N_15422,N_6501,N_11729);
nand U15423 (N_15423,N_12444,N_10837);
xnor U15424 (N_15424,N_10965,N_9760);
xor U15425 (N_15425,N_6583,N_11659);
and U15426 (N_15426,N_11485,N_9806);
xor U15427 (N_15427,N_10738,N_6261);
or U15428 (N_15428,N_11072,N_10220);
xnor U15429 (N_15429,N_12092,N_6378);
or U15430 (N_15430,N_9041,N_10502);
or U15431 (N_15431,N_6571,N_9797);
nor U15432 (N_15432,N_11313,N_10865);
xor U15433 (N_15433,N_10458,N_9382);
and U15434 (N_15434,N_12131,N_6906);
nand U15435 (N_15435,N_10003,N_10561);
and U15436 (N_15436,N_11960,N_11661);
xnor U15437 (N_15437,N_8408,N_8140);
and U15438 (N_15438,N_7575,N_11805);
xnor U15439 (N_15439,N_8080,N_10601);
or U15440 (N_15440,N_7965,N_11376);
and U15441 (N_15441,N_8502,N_9037);
nor U15442 (N_15442,N_10542,N_9071);
nor U15443 (N_15443,N_12430,N_9906);
or U15444 (N_15444,N_9637,N_7075);
or U15445 (N_15445,N_9803,N_11019);
nor U15446 (N_15446,N_9536,N_9132);
or U15447 (N_15447,N_12295,N_6671);
and U15448 (N_15448,N_12454,N_8534);
nor U15449 (N_15449,N_8997,N_6563);
nor U15450 (N_15450,N_12064,N_12072);
and U15451 (N_15451,N_6318,N_12327);
nor U15452 (N_15452,N_7762,N_8650);
nand U15453 (N_15453,N_11426,N_10303);
nand U15454 (N_15454,N_8363,N_12045);
or U15455 (N_15455,N_12123,N_7079);
nor U15456 (N_15456,N_6337,N_9950);
or U15457 (N_15457,N_9138,N_9842);
or U15458 (N_15458,N_11803,N_6312);
or U15459 (N_15459,N_11778,N_9601);
or U15460 (N_15460,N_9143,N_8957);
or U15461 (N_15461,N_7770,N_11746);
or U15462 (N_15462,N_8996,N_9017);
or U15463 (N_15463,N_6774,N_12022);
nor U15464 (N_15464,N_7501,N_12133);
or U15465 (N_15465,N_10851,N_11054);
nor U15466 (N_15466,N_8482,N_12439);
nand U15467 (N_15467,N_12130,N_11601);
xor U15468 (N_15468,N_9513,N_7440);
or U15469 (N_15469,N_6272,N_9714);
or U15470 (N_15470,N_8881,N_10077);
or U15471 (N_15471,N_9793,N_11499);
nand U15472 (N_15472,N_6572,N_8693);
nor U15473 (N_15473,N_8566,N_11518);
nor U15474 (N_15474,N_8197,N_11688);
nand U15475 (N_15475,N_12362,N_7062);
nand U15476 (N_15476,N_11846,N_8101);
nor U15477 (N_15477,N_11737,N_11758);
nand U15478 (N_15478,N_12441,N_11949);
and U15479 (N_15479,N_9158,N_7058);
xor U15480 (N_15480,N_9116,N_6262);
xnor U15481 (N_15481,N_8784,N_8426);
nand U15482 (N_15482,N_9044,N_10412);
or U15483 (N_15483,N_10869,N_10672);
and U15484 (N_15484,N_9384,N_10255);
or U15485 (N_15485,N_10092,N_7752);
nand U15486 (N_15486,N_6809,N_7140);
and U15487 (N_15487,N_9931,N_10038);
xnor U15488 (N_15488,N_6829,N_7990);
nand U15489 (N_15489,N_7353,N_7749);
and U15490 (N_15490,N_12320,N_7354);
xor U15491 (N_15491,N_6449,N_6758);
nor U15492 (N_15492,N_8368,N_10030);
or U15493 (N_15493,N_12225,N_12335);
nor U15494 (N_15494,N_12207,N_6385);
nand U15495 (N_15495,N_11620,N_6720);
and U15496 (N_15496,N_7237,N_7013);
nor U15497 (N_15497,N_7545,N_7937);
or U15498 (N_15498,N_8017,N_12321);
or U15499 (N_15499,N_10054,N_6422);
nand U15500 (N_15500,N_6918,N_8722);
or U15501 (N_15501,N_12450,N_6293);
nand U15502 (N_15502,N_6440,N_8388);
nor U15503 (N_15503,N_12472,N_10084);
nand U15504 (N_15504,N_7843,N_12453);
nand U15505 (N_15505,N_11913,N_9460);
or U15506 (N_15506,N_9432,N_12396);
and U15507 (N_15507,N_10676,N_12144);
or U15508 (N_15508,N_11760,N_9957);
nor U15509 (N_15509,N_10007,N_11733);
xor U15510 (N_15510,N_11291,N_10446);
nand U15511 (N_15511,N_10172,N_9079);
and U15512 (N_15512,N_7187,N_8339);
or U15513 (N_15513,N_10182,N_11997);
or U15514 (N_15514,N_7621,N_7490);
and U15515 (N_15515,N_8223,N_6329);
xnor U15516 (N_15516,N_9065,N_11104);
xor U15517 (N_15517,N_9624,N_8337);
or U15518 (N_15518,N_7131,N_12310);
nand U15519 (N_15519,N_11970,N_6799);
xor U15520 (N_15520,N_10259,N_9700);
nand U15521 (N_15521,N_11553,N_11337);
and U15522 (N_15522,N_7372,N_6473);
xnor U15523 (N_15523,N_9912,N_7363);
nand U15524 (N_15524,N_11564,N_11419);
nand U15525 (N_15525,N_7967,N_6566);
nor U15526 (N_15526,N_10273,N_8395);
nor U15527 (N_15527,N_7412,N_9817);
and U15528 (N_15528,N_11062,N_6311);
xnor U15529 (N_15529,N_9810,N_12404);
and U15530 (N_15530,N_11739,N_6651);
and U15531 (N_15531,N_8665,N_8075);
and U15532 (N_15532,N_6683,N_6710);
nor U15533 (N_15533,N_8274,N_8898);
or U15534 (N_15534,N_9798,N_11067);
or U15535 (N_15535,N_12284,N_9296);
and U15536 (N_15536,N_10834,N_9254);
and U15537 (N_15537,N_6573,N_6335);
nand U15538 (N_15538,N_12359,N_11947);
and U15539 (N_15539,N_7007,N_9621);
or U15540 (N_15540,N_12421,N_6841);
and U15541 (N_15541,N_12182,N_8204);
and U15542 (N_15542,N_11212,N_9118);
nor U15543 (N_15543,N_11457,N_9418);
nand U15544 (N_15544,N_10707,N_10726);
nor U15545 (N_15545,N_8963,N_8765);
or U15546 (N_15546,N_10607,N_9391);
xor U15547 (N_15547,N_7398,N_7771);
nor U15548 (N_15548,N_11845,N_8447);
xnor U15549 (N_15549,N_10694,N_7813);
or U15550 (N_15550,N_7885,N_6812);
or U15551 (N_15551,N_11904,N_11771);
xor U15552 (N_15552,N_10450,N_8369);
nand U15553 (N_15553,N_10780,N_7280);
nand U15554 (N_15554,N_8639,N_8553);
and U15555 (N_15555,N_7738,N_7180);
and U15556 (N_15556,N_10887,N_10336);
xor U15557 (N_15557,N_7920,N_11169);
xor U15558 (N_15558,N_10882,N_8014);
and U15559 (N_15559,N_7453,N_7315);
nand U15560 (N_15560,N_7124,N_10009);
nor U15561 (N_15561,N_7993,N_8989);
nand U15562 (N_15562,N_6887,N_6255);
xor U15563 (N_15563,N_9524,N_6314);
nand U15564 (N_15564,N_11626,N_12376);
nor U15565 (N_15565,N_11069,N_6502);
nor U15566 (N_15566,N_8754,N_9612);
and U15567 (N_15567,N_7664,N_6412);
or U15568 (N_15568,N_11703,N_8814);
nand U15569 (N_15569,N_11156,N_10962);
xnor U15570 (N_15570,N_8880,N_8253);
or U15571 (N_15571,N_7037,N_9129);
nand U15572 (N_15572,N_11697,N_10638);
and U15573 (N_15573,N_11598,N_9402);
and U15574 (N_15574,N_10979,N_12091);
xnor U15575 (N_15575,N_6620,N_10162);
or U15576 (N_15576,N_7559,N_12036);
nand U15577 (N_15577,N_9630,N_10368);
nor U15578 (N_15578,N_11491,N_7431);
and U15579 (N_15579,N_11188,N_12148);
nor U15580 (N_15580,N_10190,N_7435);
nor U15581 (N_15581,N_10842,N_6844);
or U15582 (N_15582,N_7221,N_6463);
and U15583 (N_15583,N_9959,N_9543);
nand U15584 (N_15584,N_11257,N_6838);
xnor U15585 (N_15585,N_9102,N_8216);
nand U15586 (N_15586,N_6821,N_12208);
nor U15587 (N_15587,N_8655,N_12343);
or U15588 (N_15588,N_6999,N_10988);
nor U15589 (N_15589,N_12296,N_12302);
xnor U15590 (N_15590,N_9476,N_7608);
xor U15591 (N_15591,N_6698,N_9371);
nand U15592 (N_15592,N_10924,N_6392);
nor U15593 (N_15593,N_8628,N_9706);
xnor U15594 (N_15594,N_12062,N_12304);
nor U15595 (N_15595,N_7188,N_9808);
or U15596 (N_15596,N_8923,N_9579);
nand U15597 (N_15597,N_11636,N_8933);
nor U15598 (N_15598,N_10179,N_11549);
nor U15599 (N_15599,N_7808,N_9324);
or U15600 (N_15600,N_12259,N_7201);
or U15601 (N_15601,N_10521,N_12009);
xor U15602 (N_15602,N_11300,N_8763);
nand U15603 (N_15603,N_8608,N_7756);
nor U15604 (N_15604,N_11246,N_10422);
or U15605 (N_15605,N_7147,N_6292);
or U15606 (N_15606,N_7427,N_10345);
nand U15607 (N_15607,N_7692,N_12002);
nand U15608 (N_15608,N_9279,N_10396);
nand U15609 (N_15609,N_8326,N_7282);
nand U15610 (N_15610,N_11348,N_8090);
and U15611 (N_15611,N_9198,N_8161);
xor U15612 (N_15612,N_8732,N_7214);
or U15613 (N_15613,N_8467,N_10178);
nand U15614 (N_15614,N_9136,N_11924);
xor U15615 (N_15615,N_7043,N_8620);
nor U15616 (N_15616,N_11716,N_9018);
xor U15617 (N_15617,N_7521,N_7833);
xor U15618 (N_15618,N_10506,N_11040);
nor U15619 (N_15619,N_12027,N_8562);
nand U15620 (N_15620,N_10444,N_7212);
xor U15621 (N_15621,N_8508,N_9737);
and U15622 (N_15622,N_11370,N_7540);
nor U15623 (N_15623,N_12319,N_10723);
nor U15624 (N_15624,N_6551,N_7662);
or U15625 (N_15625,N_11644,N_7167);
or U15626 (N_15626,N_10724,N_9258);
nand U15627 (N_15627,N_7864,N_12070);
nand U15628 (N_15628,N_9967,N_10947);
and U15629 (N_15629,N_8055,N_6769);
or U15630 (N_15630,N_8726,N_7666);
or U15631 (N_15631,N_8155,N_11473);
nand U15632 (N_15632,N_6279,N_8084);
nor U15633 (N_15633,N_8208,N_11319);
nor U15634 (N_15634,N_8202,N_9869);
nand U15635 (N_15635,N_12387,N_11637);
xnor U15636 (N_15636,N_8064,N_11571);
and U15637 (N_15637,N_7000,N_12146);
xnor U15638 (N_15638,N_11490,N_9520);
and U15639 (N_15639,N_8874,N_6267);
nand U15640 (N_15640,N_10653,N_8608);
and U15641 (N_15641,N_8496,N_10426);
and U15642 (N_15642,N_7351,N_8122);
or U15643 (N_15643,N_10516,N_10313);
or U15644 (N_15644,N_6427,N_9800);
nor U15645 (N_15645,N_9753,N_8782);
nand U15646 (N_15646,N_9618,N_8396);
and U15647 (N_15647,N_9813,N_7159);
or U15648 (N_15648,N_11684,N_7868);
and U15649 (N_15649,N_9201,N_8417);
xnor U15650 (N_15650,N_8339,N_8598);
xnor U15651 (N_15651,N_11808,N_10880);
nand U15652 (N_15652,N_6564,N_7755);
nand U15653 (N_15653,N_8631,N_9326);
and U15654 (N_15654,N_10403,N_6881);
or U15655 (N_15655,N_9043,N_7042);
xor U15656 (N_15656,N_12054,N_6904);
xor U15657 (N_15657,N_9004,N_11221);
or U15658 (N_15658,N_9248,N_11494);
nor U15659 (N_15659,N_10158,N_7923);
xnor U15660 (N_15660,N_11162,N_6692);
xor U15661 (N_15661,N_9948,N_10144);
or U15662 (N_15662,N_9754,N_7839);
and U15663 (N_15663,N_10135,N_7462);
and U15664 (N_15664,N_10692,N_12151);
nor U15665 (N_15665,N_9970,N_8294);
or U15666 (N_15666,N_11494,N_11774);
nor U15667 (N_15667,N_6499,N_9960);
nor U15668 (N_15668,N_11418,N_11859);
nor U15669 (N_15669,N_9857,N_10766);
xor U15670 (N_15670,N_11714,N_6538);
or U15671 (N_15671,N_9473,N_9064);
and U15672 (N_15672,N_8283,N_7683);
xor U15673 (N_15673,N_6848,N_9798);
or U15674 (N_15674,N_11171,N_8939);
or U15675 (N_15675,N_7857,N_6837);
and U15676 (N_15676,N_11070,N_11853);
and U15677 (N_15677,N_7457,N_10238);
or U15678 (N_15678,N_7593,N_9301);
or U15679 (N_15679,N_7163,N_11429);
nand U15680 (N_15680,N_6420,N_7022);
and U15681 (N_15681,N_9838,N_6361);
xnor U15682 (N_15682,N_6839,N_6307);
nand U15683 (N_15683,N_12412,N_9204);
or U15684 (N_15684,N_7931,N_7975);
nand U15685 (N_15685,N_10008,N_7134);
and U15686 (N_15686,N_9233,N_11679);
or U15687 (N_15687,N_9289,N_9029);
nand U15688 (N_15688,N_9846,N_7246);
xor U15689 (N_15689,N_7499,N_9809);
nor U15690 (N_15690,N_8155,N_11335);
nand U15691 (N_15691,N_12463,N_7664);
and U15692 (N_15692,N_9041,N_10662);
xor U15693 (N_15693,N_11891,N_9134);
and U15694 (N_15694,N_9443,N_12344);
nor U15695 (N_15695,N_7598,N_8646);
and U15696 (N_15696,N_9018,N_11316);
nand U15697 (N_15697,N_6449,N_10934);
xor U15698 (N_15698,N_6363,N_11752);
nor U15699 (N_15699,N_7786,N_8953);
or U15700 (N_15700,N_7573,N_9144);
and U15701 (N_15701,N_11798,N_10105);
xnor U15702 (N_15702,N_7059,N_9011);
xnor U15703 (N_15703,N_10890,N_7116);
nand U15704 (N_15704,N_11212,N_10147);
xor U15705 (N_15705,N_7294,N_9801);
nand U15706 (N_15706,N_8704,N_7478);
nor U15707 (N_15707,N_9301,N_11008);
and U15708 (N_15708,N_10787,N_11978);
nor U15709 (N_15709,N_9514,N_11907);
nand U15710 (N_15710,N_8362,N_9904);
nand U15711 (N_15711,N_7460,N_8746);
nor U15712 (N_15712,N_6726,N_9529);
nor U15713 (N_15713,N_10882,N_12407);
nand U15714 (N_15714,N_12266,N_9162);
and U15715 (N_15715,N_12285,N_9199);
nor U15716 (N_15716,N_6913,N_10572);
nor U15717 (N_15717,N_8978,N_6807);
and U15718 (N_15718,N_9077,N_6986);
and U15719 (N_15719,N_9840,N_9537);
and U15720 (N_15720,N_7167,N_6645);
and U15721 (N_15721,N_6319,N_8682);
or U15722 (N_15722,N_7261,N_11877);
nand U15723 (N_15723,N_8819,N_9051);
and U15724 (N_15724,N_11662,N_10939);
xnor U15725 (N_15725,N_9116,N_10003);
xor U15726 (N_15726,N_7963,N_7957);
nor U15727 (N_15727,N_7339,N_7512);
or U15728 (N_15728,N_6945,N_7196);
nor U15729 (N_15729,N_12144,N_12477);
xnor U15730 (N_15730,N_12125,N_10748);
or U15731 (N_15731,N_7433,N_9392);
and U15732 (N_15732,N_8729,N_12049);
and U15733 (N_15733,N_8139,N_9507);
and U15734 (N_15734,N_6275,N_11730);
nand U15735 (N_15735,N_10305,N_8932);
nor U15736 (N_15736,N_10318,N_11324);
nand U15737 (N_15737,N_6324,N_10967);
xnor U15738 (N_15738,N_9198,N_11787);
nor U15739 (N_15739,N_12455,N_9648);
and U15740 (N_15740,N_6564,N_8966);
nand U15741 (N_15741,N_12457,N_7644);
and U15742 (N_15742,N_12017,N_6679);
nor U15743 (N_15743,N_7151,N_7559);
and U15744 (N_15744,N_6781,N_7985);
nor U15745 (N_15745,N_10989,N_9045);
or U15746 (N_15746,N_9255,N_6535);
nor U15747 (N_15747,N_7603,N_6431);
nor U15748 (N_15748,N_6770,N_7667);
xnor U15749 (N_15749,N_7649,N_8395);
or U15750 (N_15750,N_6674,N_11929);
or U15751 (N_15751,N_7425,N_10201);
xor U15752 (N_15752,N_10521,N_8075);
xor U15753 (N_15753,N_9892,N_6830);
xnor U15754 (N_15754,N_9463,N_7703);
nor U15755 (N_15755,N_8529,N_12109);
nand U15756 (N_15756,N_7188,N_10214);
and U15757 (N_15757,N_6702,N_12358);
and U15758 (N_15758,N_10225,N_10860);
or U15759 (N_15759,N_7146,N_12313);
or U15760 (N_15760,N_6840,N_9955);
and U15761 (N_15761,N_10937,N_6566);
xor U15762 (N_15762,N_6907,N_8905);
xor U15763 (N_15763,N_11579,N_8923);
or U15764 (N_15764,N_12311,N_11144);
nand U15765 (N_15765,N_10864,N_10392);
nor U15766 (N_15766,N_7999,N_8056);
nand U15767 (N_15767,N_12351,N_9219);
nor U15768 (N_15768,N_10729,N_12434);
and U15769 (N_15769,N_11442,N_6432);
or U15770 (N_15770,N_7616,N_12428);
or U15771 (N_15771,N_8818,N_7443);
nand U15772 (N_15772,N_6894,N_9378);
nand U15773 (N_15773,N_12110,N_12188);
and U15774 (N_15774,N_10175,N_10758);
and U15775 (N_15775,N_7555,N_12143);
nor U15776 (N_15776,N_11684,N_12238);
nor U15777 (N_15777,N_11545,N_10731);
and U15778 (N_15778,N_7363,N_10624);
and U15779 (N_15779,N_7485,N_10241);
or U15780 (N_15780,N_7669,N_10538);
or U15781 (N_15781,N_11377,N_11995);
nor U15782 (N_15782,N_12282,N_10958);
and U15783 (N_15783,N_8635,N_6825);
nand U15784 (N_15784,N_7551,N_12368);
or U15785 (N_15785,N_12086,N_11142);
nor U15786 (N_15786,N_6269,N_7821);
or U15787 (N_15787,N_6405,N_12282);
and U15788 (N_15788,N_6594,N_7181);
and U15789 (N_15789,N_9896,N_7000);
and U15790 (N_15790,N_8078,N_8102);
xor U15791 (N_15791,N_8700,N_11133);
nand U15792 (N_15792,N_11759,N_10974);
nor U15793 (N_15793,N_12171,N_8075);
xor U15794 (N_15794,N_6388,N_6625);
and U15795 (N_15795,N_9896,N_11969);
nand U15796 (N_15796,N_7189,N_10937);
and U15797 (N_15797,N_8395,N_7661);
nor U15798 (N_15798,N_7484,N_11652);
or U15799 (N_15799,N_11437,N_10012);
nor U15800 (N_15800,N_7586,N_8472);
xnor U15801 (N_15801,N_9622,N_6289);
nor U15802 (N_15802,N_7653,N_7572);
nand U15803 (N_15803,N_10751,N_7902);
nand U15804 (N_15804,N_9306,N_7347);
nor U15805 (N_15805,N_12375,N_9660);
nor U15806 (N_15806,N_10023,N_12318);
or U15807 (N_15807,N_12042,N_10520);
and U15808 (N_15808,N_10664,N_9858);
or U15809 (N_15809,N_6820,N_8553);
and U15810 (N_15810,N_8957,N_9489);
nor U15811 (N_15811,N_8806,N_8507);
xnor U15812 (N_15812,N_6467,N_6643);
or U15813 (N_15813,N_7504,N_6873);
xor U15814 (N_15814,N_10076,N_7017);
or U15815 (N_15815,N_7027,N_6379);
nand U15816 (N_15816,N_10255,N_11651);
xor U15817 (N_15817,N_9569,N_9862);
nand U15818 (N_15818,N_9191,N_6573);
nor U15819 (N_15819,N_11947,N_10293);
or U15820 (N_15820,N_8934,N_12193);
and U15821 (N_15821,N_6926,N_7852);
nor U15822 (N_15822,N_8684,N_10177);
or U15823 (N_15823,N_8598,N_7160);
or U15824 (N_15824,N_9022,N_7024);
nand U15825 (N_15825,N_11528,N_11482);
and U15826 (N_15826,N_9451,N_10801);
nor U15827 (N_15827,N_8037,N_6786);
and U15828 (N_15828,N_8545,N_7990);
nand U15829 (N_15829,N_10937,N_9608);
or U15830 (N_15830,N_12450,N_12326);
nand U15831 (N_15831,N_8357,N_7744);
xnor U15832 (N_15832,N_11213,N_7198);
nor U15833 (N_15833,N_9504,N_9145);
nor U15834 (N_15834,N_11659,N_10961);
or U15835 (N_15835,N_7744,N_9038);
xnor U15836 (N_15836,N_7155,N_9277);
xnor U15837 (N_15837,N_8215,N_8329);
nor U15838 (N_15838,N_7114,N_9925);
nand U15839 (N_15839,N_12227,N_11179);
xor U15840 (N_15840,N_11468,N_6608);
and U15841 (N_15841,N_7271,N_10120);
and U15842 (N_15842,N_12240,N_10581);
or U15843 (N_15843,N_7413,N_12150);
nor U15844 (N_15844,N_11588,N_9555);
and U15845 (N_15845,N_7532,N_11530);
xnor U15846 (N_15846,N_7214,N_8611);
nand U15847 (N_15847,N_10504,N_11561);
or U15848 (N_15848,N_6614,N_10129);
and U15849 (N_15849,N_7723,N_6808);
nor U15850 (N_15850,N_10631,N_7193);
or U15851 (N_15851,N_12430,N_11201);
xor U15852 (N_15852,N_7750,N_8351);
or U15853 (N_15853,N_12119,N_8912);
xor U15854 (N_15854,N_11653,N_6687);
nor U15855 (N_15855,N_9262,N_10960);
nor U15856 (N_15856,N_8012,N_9052);
or U15857 (N_15857,N_12400,N_10997);
or U15858 (N_15858,N_9167,N_11391);
or U15859 (N_15859,N_10665,N_7297);
and U15860 (N_15860,N_7271,N_7813);
nor U15861 (N_15861,N_9265,N_11948);
or U15862 (N_15862,N_11392,N_10458);
nor U15863 (N_15863,N_9417,N_8594);
nand U15864 (N_15864,N_10619,N_10517);
or U15865 (N_15865,N_7739,N_8104);
nand U15866 (N_15866,N_11139,N_7590);
xor U15867 (N_15867,N_8273,N_11963);
or U15868 (N_15868,N_6854,N_10701);
nor U15869 (N_15869,N_11083,N_7234);
nand U15870 (N_15870,N_11001,N_7854);
and U15871 (N_15871,N_10058,N_9737);
and U15872 (N_15872,N_9886,N_7042);
nor U15873 (N_15873,N_6928,N_12059);
xnor U15874 (N_15874,N_10094,N_12061);
nor U15875 (N_15875,N_9157,N_7692);
nand U15876 (N_15876,N_12492,N_12052);
nand U15877 (N_15877,N_8592,N_10412);
nand U15878 (N_15878,N_7154,N_6613);
and U15879 (N_15879,N_7244,N_10254);
nor U15880 (N_15880,N_9815,N_11650);
or U15881 (N_15881,N_12046,N_10975);
and U15882 (N_15882,N_10495,N_10544);
nand U15883 (N_15883,N_11882,N_8530);
nor U15884 (N_15884,N_11885,N_9896);
xor U15885 (N_15885,N_11766,N_10174);
nor U15886 (N_15886,N_9704,N_11401);
and U15887 (N_15887,N_11283,N_7947);
nand U15888 (N_15888,N_9285,N_7244);
nand U15889 (N_15889,N_6356,N_6704);
nand U15890 (N_15890,N_11970,N_8110);
and U15891 (N_15891,N_8401,N_8966);
nor U15892 (N_15892,N_10036,N_7982);
or U15893 (N_15893,N_8147,N_10562);
or U15894 (N_15894,N_9124,N_6535);
and U15895 (N_15895,N_8057,N_9997);
nand U15896 (N_15896,N_9247,N_9003);
or U15897 (N_15897,N_10508,N_11054);
xnor U15898 (N_15898,N_11431,N_10369);
xor U15899 (N_15899,N_8641,N_7657);
or U15900 (N_15900,N_9390,N_8786);
and U15901 (N_15901,N_6870,N_7488);
nor U15902 (N_15902,N_9358,N_8889);
nor U15903 (N_15903,N_10204,N_7437);
and U15904 (N_15904,N_8107,N_10615);
nand U15905 (N_15905,N_12196,N_11718);
xor U15906 (N_15906,N_10575,N_9001);
xor U15907 (N_15907,N_6988,N_10043);
xnor U15908 (N_15908,N_6752,N_6490);
nor U15909 (N_15909,N_10408,N_7086);
xor U15910 (N_15910,N_7713,N_9957);
and U15911 (N_15911,N_9678,N_7901);
or U15912 (N_15912,N_10912,N_10555);
xnor U15913 (N_15913,N_11810,N_11200);
nand U15914 (N_15914,N_8522,N_8039);
nand U15915 (N_15915,N_10424,N_6795);
nor U15916 (N_15916,N_7713,N_10675);
and U15917 (N_15917,N_9413,N_12139);
xor U15918 (N_15918,N_11701,N_6829);
and U15919 (N_15919,N_11425,N_7706);
xor U15920 (N_15920,N_11909,N_9301);
or U15921 (N_15921,N_7692,N_12064);
or U15922 (N_15922,N_7606,N_6671);
or U15923 (N_15923,N_7292,N_7534);
or U15924 (N_15924,N_9983,N_6803);
nand U15925 (N_15925,N_6809,N_11175);
and U15926 (N_15926,N_11323,N_12204);
nand U15927 (N_15927,N_7029,N_7930);
xnor U15928 (N_15928,N_10008,N_9352);
or U15929 (N_15929,N_6591,N_8704);
nand U15930 (N_15930,N_9015,N_7192);
or U15931 (N_15931,N_8052,N_12476);
and U15932 (N_15932,N_8377,N_8257);
nor U15933 (N_15933,N_6737,N_8251);
nand U15934 (N_15934,N_10324,N_8178);
and U15935 (N_15935,N_8123,N_11860);
or U15936 (N_15936,N_6992,N_11247);
xnor U15937 (N_15937,N_12488,N_11412);
and U15938 (N_15938,N_7810,N_10724);
and U15939 (N_15939,N_12407,N_9802);
xor U15940 (N_15940,N_8702,N_9546);
nor U15941 (N_15941,N_6438,N_10399);
and U15942 (N_15942,N_9154,N_11974);
or U15943 (N_15943,N_9200,N_6902);
or U15944 (N_15944,N_7690,N_7807);
or U15945 (N_15945,N_9418,N_9712);
or U15946 (N_15946,N_6562,N_9192);
or U15947 (N_15947,N_9523,N_10288);
and U15948 (N_15948,N_10781,N_10266);
nand U15949 (N_15949,N_6495,N_7442);
xnor U15950 (N_15950,N_11554,N_8986);
xnor U15951 (N_15951,N_9495,N_9899);
or U15952 (N_15952,N_8060,N_7210);
or U15953 (N_15953,N_9985,N_9830);
xor U15954 (N_15954,N_8414,N_10351);
or U15955 (N_15955,N_8634,N_9050);
xor U15956 (N_15956,N_10297,N_11477);
and U15957 (N_15957,N_8894,N_7991);
and U15958 (N_15958,N_10285,N_12041);
nand U15959 (N_15959,N_7191,N_8056);
and U15960 (N_15960,N_7925,N_10501);
xnor U15961 (N_15961,N_8672,N_8591);
or U15962 (N_15962,N_11604,N_9810);
or U15963 (N_15963,N_8102,N_6904);
or U15964 (N_15964,N_12458,N_8352);
nor U15965 (N_15965,N_6299,N_11679);
nor U15966 (N_15966,N_9828,N_9262);
or U15967 (N_15967,N_8498,N_8039);
nor U15968 (N_15968,N_11367,N_11230);
nand U15969 (N_15969,N_12213,N_7657);
xor U15970 (N_15970,N_10490,N_7938);
nor U15971 (N_15971,N_9463,N_12232);
xor U15972 (N_15972,N_10053,N_10659);
nor U15973 (N_15973,N_7085,N_6677);
xor U15974 (N_15974,N_11943,N_12031);
or U15975 (N_15975,N_8640,N_10827);
and U15976 (N_15976,N_10780,N_12491);
xnor U15977 (N_15977,N_8446,N_6632);
xor U15978 (N_15978,N_11563,N_11237);
or U15979 (N_15979,N_8052,N_9751);
or U15980 (N_15980,N_10770,N_6990);
nor U15981 (N_15981,N_8421,N_6802);
and U15982 (N_15982,N_9081,N_12067);
and U15983 (N_15983,N_11342,N_8541);
and U15984 (N_15984,N_7080,N_12271);
and U15985 (N_15985,N_10542,N_6583);
xnor U15986 (N_15986,N_11488,N_11996);
xor U15987 (N_15987,N_9728,N_11989);
and U15988 (N_15988,N_9457,N_9218);
or U15989 (N_15989,N_7945,N_11620);
nor U15990 (N_15990,N_7797,N_9335);
nand U15991 (N_15991,N_8116,N_8146);
nor U15992 (N_15992,N_7513,N_6535);
xnor U15993 (N_15993,N_10263,N_11586);
and U15994 (N_15994,N_9001,N_7218);
nor U15995 (N_15995,N_7617,N_7607);
or U15996 (N_15996,N_11210,N_8694);
nor U15997 (N_15997,N_9623,N_8418);
nor U15998 (N_15998,N_6423,N_11611);
and U15999 (N_15999,N_7922,N_7466);
and U16000 (N_16000,N_9010,N_6363);
and U16001 (N_16001,N_11447,N_9743);
nor U16002 (N_16002,N_7726,N_11826);
nand U16003 (N_16003,N_10900,N_7486);
xnor U16004 (N_16004,N_6648,N_6377);
nor U16005 (N_16005,N_12213,N_11023);
or U16006 (N_16006,N_11756,N_7433);
nand U16007 (N_16007,N_6959,N_6877);
nor U16008 (N_16008,N_9956,N_9807);
nor U16009 (N_16009,N_9435,N_6907);
nor U16010 (N_16010,N_10078,N_9212);
nor U16011 (N_16011,N_12448,N_8667);
or U16012 (N_16012,N_8909,N_11523);
xnor U16013 (N_16013,N_7657,N_10590);
or U16014 (N_16014,N_8314,N_8784);
xnor U16015 (N_16015,N_11481,N_8284);
and U16016 (N_16016,N_6590,N_8845);
nand U16017 (N_16017,N_12028,N_11301);
or U16018 (N_16018,N_8764,N_8621);
and U16019 (N_16019,N_10230,N_10102);
or U16020 (N_16020,N_10078,N_10337);
or U16021 (N_16021,N_9281,N_9081);
xnor U16022 (N_16022,N_7423,N_9232);
nor U16023 (N_16023,N_8123,N_11659);
nor U16024 (N_16024,N_11996,N_8418);
nand U16025 (N_16025,N_9638,N_9641);
nand U16026 (N_16026,N_8030,N_12033);
and U16027 (N_16027,N_8871,N_9036);
or U16028 (N_16028,N_7993,N_10822);
xnor U16029 (N_16029,N_6864,N_11802);
nor U16030 (N_16030,N_11154,N_11915);
or U16031 (N_16031,N_11270,N_9709);
nand U16032 (N_16032,N_10167,N_9616);
nor U16033 (N_16033,N_9391,N_11164);
or U16034 (N_16034,N_10239,N_10351);
and U16035 (N_16035,N_12084,N_9109);
and U16036 (N_16036,N_8879,N_7678);
nand U16037 (N_16037,N_10501,N_11519);
and U16038 (N_16038,N_6844,N_10849);
and U16039 (N_16039,N_6364,N_8120);
nand U16040 (N_16040,N_8388,N_8519);
xnor U16041 (N_16041,N_10246,N_9319);
or U16042 (N_16042,N_11517,N_10625);
nand U16043 (N_16043,N_11890,N_12212);
nor U16044 (N_16044,N_11294,N_10365);
xnor U16045 (N_16045,N_11283,N_8230);
and U16046 (N_16046,N_6573,N_9098);
or U16047 (N_16047,N_10574,N_6252);
nand U16048 (N_16048,N_10759,N_8655);
xnor U16049 (N_16049,N_8046,N_7778);
nor U16050 (N_16050,N_6496,N_10331);
xnor U16051 (N_16051,N_10889,N_11781);
xor U16052 (N_16052,N_11158,N_12040);
and U16053 (N_16053,N_11743,N_8738);
xor U16054 (N_16054,N_7661,N_11496);
nor U16055 (N_16055,N_12172,N_9178);
and U16056 (N_16056,N_7744,N_7307);
and U16057 (N_16057,N_10708,N_10073);
or U16058 (N_16058,N_11129,N_6543);
nand U16059 (N_16059,N_7414,N_9210);
nand U16060 (N_16060,N_10121,N_8347);
or U16061 (N_16061,N_10811,N_7890);
xor U16062 (N_16062,N_8253,N_9582);
xor U16063 (N_16063,N_7511,N_10205);
xor U16064 (N_16064,N_10567,N_9555);
nor U16065 (N_16065,N_10317,N_11126);
nand U16066 (N_16066,N_10733,N_10839);
nand U16067 (N_16067,N_12245,N_9464);
xor U16068 (N_16068,N_7462,N_8901);
or U16069 (N_16069,N_12498,N_8747);
or U16070 (N_16070,N_10429,N_6865);
or U16071 (N_16071,N_8661,N_11529);
or U16072 (N_16072,N_10212,N_12319);
xor U16073 (N_16073,N_11768,N_11901);
nor U16074 (N_16074,N_11983,N_11973);
xnor U16075 (N_16075,N_9046,N_10262);
nand U16076 (N_16076,N_10292,N_6272);
nand U16077 (N_16077,N_7283,N_7490);
xnor U16078 (N_16078,N_11912,N_9272);
xnor U16079 (N_16079,N_7578,N_8852);
xor U16080 (N_16080,N_11986,N_9390);
or U16081 (N_16081,N_11191,N_9418);
and U16082 (N_16082,N_9301,N_10673);
nand U16083 (N_16083,N_11835,N_9125);
nor U16084 (N_16084,N_9692,N_7901);
nor U16085 (N_16085,N_7001,N_12104);
and U16086 (N_16086,N_9758,N_11414);
nand U16087 (N_16087,N_12111,N_7726);
and U16088 (N_16088,N_8906,N_9168);
nand U16089 (N_16089,N_12008,N_11197);
nor U16090 (N_16090,N_12066,N_12454);
or U16091 (N_16091,N_11327,N_7531);
xnor U16092 (N_16092,N_12374,N_7068);
nor U16093 (N_16093,N_8322,N_10805);
and U16094 (N_16094,N_10748,N_10501);
nand U16095 (N_16095,N_11136,N_10133);
and U16096 (N_16096,N_9564,N_7692);
and U16097 (N_16097,N_12010,N_7772);
nor U16098 (N_16098,N_11311,N_11069);
and U16099 (N_16099,N_9141,N_10847);
xor U16100 (N_16100,N_7310,N_8480);
and U16101 (N_16101,N_8873,N_11124);
nor U16102 (N_16102,N_7898,N_8680);
or U16103 (N_16103,N_6975,N_7290);
or U16104 (N_16104,N_6334,N_7617);
xnor U16105 (N_16105,N_6390,N_11037);
nor U16106 (N_16106,N_7566,N_8725);
nor U16107 (N_16107,N_6811,N_12013);
nand U16108 (N_16108,N_11871,N_9899);
nand U16109 (N_16109,N_7271,N_8590);
or U16110 (N_16110,N_7607,N_9861);
nor U16111 (N_16111,N_10938,N_11180);
or U16112 (N_16112,N_6939,N_9034);
nand U16113 (N_16113,N_6513,N_10585);
and U16114 (N_16114,N_12101,N_8345);
and U16115 (N_16115,N_7756,N_8635);
nand U16116 (N_16116,N_6259,N_9330);
and U16117 (N_16117,N_10343,N_6292);
nand U16118 (N_16118,N_10706,N_8178);
nand U16119 (N_16119,N_6980,N_8355);
nor U16120 (N_16120,N_11745,N_12492);
or U16121 (N_16121,N_11779,N_9369);
nor U16122 (N_16122,N_6395,N_8774);
nand U16123 (N_16123,N_12097,N_8386);
xnor U16124 (N_16124,N_10036,N_7736);
and U16125 (N_16125,N_8384,N_11393);
nor U16126 (N_16126,N_9480,N_10646);
or U16127 (N_16127,N_10518,N_12284);
nand U16128 (N_16128,N_10533,N_8365);
or U16129 (N_16129,N_11289,N_6352);
or U16130 (N_16130,N_10627,N_9408);
and U16131 (N_16131,N_8221,N_7263);
nor U16132 (N_16132,N_8785,N_9891);
nand U16133 (N_16133,N_7045,N_7870);
xnor U16134 (N_16134,N_7060,N_7650);
nand U16135 (N_16135,N_6459,N_12057);
nand U16136 (N_16136,N_11091,N_10407);
or U16137 (N_16137,N_10510,N_10719);
nor U16138 (N_16138,N_7818,N_9788);
and U16139 (N_16139,N_8668,N_10727);
and U16140 (N_16140,N_10760,N_8473);
or U16141 (N_16141,N_9796,N_7263);
nand U16142 (N_16142,N_8380,N_9468);
xnor U16143 (N_16143,N_12075,N_12268);
and U16144 (N_16144,N_12032,N_6880);
nor U16145 (N_16145,N_8657,N_8384);
or U16146 (N_16146,N_9111,N_8558);
xnor U16147 (N_16147,N_12375,N_9428);
and U16148 (N_16148,N_9082,N_6947);
and U16149 (N_16149,N_6377,N_11289);
nor U16150 (N_16150,N_7853,N_7456);
and U16151 (N_16151,N_9623,N_8089);
or U16152 (N_16152,N_12295,N_10807);
or U16153 (N_16153,N_6258,N_11093);
nand U16154 (N_16154,N_7339,N_8279);
nor U16155 (N_16155,N_10966,N_10213);
nor U16156 (N_16156,N_8466,N_9043);
nor U16157 (N_16157,N_12367,N_10496);
xnor U16158 (N_16158,N_9917,N_12339);
or U16159 (N_16159,N_6508,N_7711);
xnor U16160 (N_16160,N_8207,N_10852);
xor U16161 (N_16161,N_10406,N_6325);
or U16162 (N_16162,N_12388,N_9293);
xnor U16163 (N_16163,N_11371,N_7733);
xnor U16164 (N_16164,N_7929,N_12110);
nand U16165 (N_16165,N_10463,N_9257);
xor U16166 (N_16166,N_8262,N_11308);
nand U16167 (N_16167,N_7441,N_6705);
nand U16168 (N_16168,N_11089,N_12362);
or U16169 (N_16169,N_7315,N_12384);
xnor U16170 (N_16170,N_6381,N_11517);
or U16171 (N_16171,N_12470,N_11574);
xnor U16172 (N_16172,N_12283,N_10437);
and U16173 (N_16173,N_12013,N_8037);
nor U16174 (N_16174,N_10764,N_9510);
or U16175 (N_16175,N_6536,N_7415);
nor U16176 (N_16176,N_8375,N_6900);
or U16177 (N_16177,N_10282,N_9059);
and U16178 (N_16178,N_7821,N_9259);
and U16179 (N_16179,N_12244,N_8283);
or U16180 (N_16180,N_12236,N_11381);
and U16181 (N_16181,N_8220,N_12489);
nand U16182 (N_16182,N_11368,N_8440);
and U16183 (N_16183,N_9327,N_10900);
nand U16184 (N_16184,N_8003,N_11187);
xnor U16185 (N_16185,N_11738,N_11141);
xnor U16186 (N_16186,N_8511,N_9007);
and U16187 (N_16187,N_9652,N_8157);
xor U16188 (N_16188,N_6914,N_7480);
or U16189 (N_16189,N_7901,N_9399);
or U16190 (N_16190,N_10076,N_8758);
nor U16191 (N_16191,N_7551,N_9257);
xnor U16192 (N_16192,N_7757,N_6823);
nand U16193 (N_16193,N_10362,N_10776);
or U16194 (N_16194,N_6398,N_8422);
nand U16195 (N_16195,N_7123,N_8737);
xor U16196 (N_16196,N_10132,N_9045);
xor U16197 (N_16197,N_8036,N_8546);
nand U16198 (N_16198,N_10027,N_9111);
or U16199 (N_16199,N_8871,N_6691);
xor U16200 (N_16200,N_10450,N_9332);
xnor U16201 (N_16201,N_8935,N_10755);
nor U16202 (N_16202,N_11227,N_7539);
or U16203 (N_16203,N_8181,N_8677);
nor U16204 (N_16204,N_10098,N_6951);
xnor U16205 (N_16205,N_6981,N_10825);
nor U16206 (N_16206,N_10894,N_9282);
or U16207 (N_16207,N_8648,N_10165);
nand U16208 (N_16208,N_8562,N_8277);
nand U16209 (N_16209,N_7623,N_7474);
nand U16210 (N_16210,N_9840,N_12405);
nor U16211 (N_16211,N_7694,N_9627);
and U16212 (N_16212,N_11200,N_9243);
or U16213 (N_16213,N_12387,N_9680);
xor U16214 (N_16214,N_6965,N_9059);
nor U16215 (N_16215,N_7240,N_9831);
or U16216 (N_16216,N_6587,N_8660);
xor U16217 (N_16217,N_9302,N_8271);
nor U16218 (N_16218,N_7412,N_9017);
nor U16219 (N_16219,N_10815,N_8867);
nor U16220 (N_16220,N_11423,N_10263);
and U16221 (N_16221,N_8899,N_12390);
and U16222 (N_16222,N_11566,N_6849);
nand U16223 (N_16223,N_10060,N_12447);
nand U16224 (N_16224,N_11301,N_10104);
nand U16225 (N_16225,N_6819,N_9851);
xnor U16226 (N_16226,N_8597,N_7194);
and U16227 (N_16227,N_7230,N_6824);
and U16228 (N_16228,N_7879,N_11994);
and U16229 (N_16229,N_11337,N_7906);
and U16230 (N_16230,N_11721,N_9164);
or U16231 (N_16231,N_10336,N_9653);
xnor U16232 (N_16232,N_9669,N_8534);
xor U16233 (N_16233,N_7659,N_8104);
nand U16234 (N_16234,N_10493,N_8854);
nand U16235 (N_16235,N_10638,N_9380);
nor U16236 (N_16236,N_10700,N_7710);
xor U16237 (N_16237,N_6587,N_10193);
or U16238 (N_16238,N_10376,N_9470);
or U16239 (N_16239,N_10963,N_12474);
and U16240 (N_16240,N_9312,N_10226);
nor U16241 (N_16241,N_8425,N_10813);
or U16242 (N_16242,N_7970,N_11249);
or U16243 (N_16243,N_10931,N_10140);
xnor U16244 (N_16244,N_11138,N_10476);
and U16245 (N_16245,N_6825,N_12189);
and U16246 (N_16246,N_9470,N_9014);
or U16247 (N_16247,N_9403,N_8023);
and U16248 (N_16248,N_6330,N_11132);
nand U16249 (N_16249,N_11427,N_8286);
nand U16250 (N_16250,N_8704,N_6895);
xnor U16251 (N_16251,N_7751,N_12386);
nor U16252 (N_16252,N_8330,N_10714);
xor U16253 (N_16253,N_7824,N_7678);
nand U16254 (N_16254,N_8662,N_8705);
or U16255 (N_16255,N_11076,N_6676);
and U16256 (N_16256,N_10533,N_7665);
nand U16257 (N_16257,N_6318,N_10403);
nand U16258 (N_16258,N_12140,N_9201);
nor U16259 (N_16259,N_6960,N_7110);
and U16260 (N_16260,N_6797,N_7746);
or U16261 (N_16261,N_7240,N_7295);
nor U16262 (N_16262,N_9822,N_6552);
and U16263 (N_16263,N_9327,N_9044);
and U16264 (N_16264,N_11957,N_11683);
and U16265 (N_16265,N_10006,N_6476);
nor U16266 (N_16266,N_7714,N_7000);
xnor U16267 (N_16267,N_12357,N_8941);
nor U16268 (N_16268,N_9413,N_12395);
xnor U16269 (N_16269,N_9571,N_6356);
nand U16270 (N_16270,N_12281,N_11731);
xnor U16271 (N_16271,N_7488,N_10589);
or U16272 (N_16272,N_11319,N_7195);
and U16273 (N_16273,N_11383,N_8868);
or U16274 (N_16274,N_11622,N_10080);
nor U16275 (N_16275,N_7821,N_11480);
nor U16276 (N_16276,N_10572,N_9361);
nor U16277 (N_16277,N_6854,N_10830);
nand U16278 (N_16278,N_12494,N_12386);
nor U16279 (N_16279,N_11076,N_11720);
or U16280 (N_16280,N_10587,N_9754);
xor U16281 (N_16281,N_8388,N_6802);
nor U16282 (N_16282,N_10505,N_6488);
and U16283 (N_16283,N_10500,N_11798);
nand U16284 (N_16284,N_7134,N_11389);
and U16285 (N_16285,N_10242,N_8044);
nor U16286 (N_16286,N_10147,N_9936);
and U16287 (N_16287,N_6836,N_6412);
nand U16288 (N_16288,N_12400,N_9470);
xor U16289 (N_16289,N_6545,N_8068);
nand U16290 (N_16290,N_12031,N_10171);
nor U16291 (N_16291,N_11948,N_10030);
and U16292 (N_16292,N_10665,N_7116);
nor U16293 (N_16293,N_9434,N_10366);
and U16294 (N_16294,N_11626,N_11067);
nor U16295 (N_16295,N_8412,N_8823);
or U16296 (N_16296,N_7973,N_9207);
nand U16297 (N_16297,N_11135,N_6312);
nor U16298 (N_16298,N_9032,N_11624);
and U16299 (N_16299,N_7878,N_8044);
xnor U16300 (N_16300,N_9842,N_9430);
xor U16301 (N_16301,N_7401,N_8576);
and U16302 (N_16302,N_10856,N_8516);
and U16303 (N_16303,N_9031,N_9345);
xnor U16304 (N_16304,N_7539,N_8085);
or U16305 (N_16305,N_10301,N_7790);
nand U16306 (N_16306,N_9715,N_9718);
or U16307 (N_16307,N_7250,N_10683);
nor U16308 (N_16308,N_9887,N_6484);
xnor U16309 (N_16309,N_6693,N_12372);
nor U16310 (N_16310,N_8708,N_6349);
nand U16311 (N_16311,N_12239,N_10234);
nand U16312 (N_16312,N_7712,N_10260);
or U16313 (N_16313,N_9970,N_10293);
nand U16314 (N_16314,N_11463,N_10011);
nor U16315 (N_16315,N_6868,N_7120);
xor U16316 (N_16316,N_7455,N_12091);
or U16317 (N_16317,N_9581,N_6908);
and U16318 (N_16318,N_10304,N_10952);
nand U16319 (N_16319,N_9716,N_11556);
nand U16320 (N_16320,N_7995,N_10842);
nand U16321 (N_16321,N_10493,N_10621);
and U16322 (N_16322,N_10514,N_8245);
xor U16323 (N_16323,N_8163,N_11084);
or U16324 (N_16324,N_6288,N_9185);
or U16325 (N_16325,N_8094,N_8038);
xor U16326 (N_16326,N_8051,N_8055);
xnor U16327 (N_16327,N_6616,N_11819);
nand U16328 (N_16328,N_11053,N_10706);
nor U16329 (N_16329,N_12413,N_8587);
nand U16330 (N_16330,N_7200,N_7272);
and U16331 (N_16331,N_7769,N_10747);
nand U16332 (N_16332,N_7179,N_7627);
or U16333 (N_16333,N_11394,N_10580);
nand U16334 (N_16334,N_10400,N_12338);
or U16335 (N_16335,N_11012,N_7406);
nand U16336 (N_16336,N_7864,N_8187);
and U16337 (N_16337,N_6641,N_6531);
or U16338 (N_16338,N_6376,N_11685);
nor U16339 (N_16339,N_10250,N_10987);
or U16340 (N_16340,N_9944,N_10716);
and U16341 (N_16341,N_12318,N_9700);
xor U16342 (N_16342,N_12338,N_7011);
and U16343 (N_16343,N_7086,N_11009);
nor U16344 (N_16344,N_9497,N_11012);
xnor U16345 (N_16345,N_9117,N_7712);
xnor U16346 (N_16346,N_9620,N_11358);
or U16347 (N_16347,N_10616,N_11917);
nor U16348 (N_16348,N_12299,N_9305);
and U16349 (N_16349,N_12067,N_8218);
nor U16350 (N_16350,N_11965,N_9035);
xnor U16351 (N_16351,N_10190,N_10561);
nand U16352 (N_16352,N_10694,N_10162);
xor U16353 (N_16353,N_12077,N_10700);
or U16354 (N_16354,N_10810,N_7311);
and U16355 (N_16355,N_11269,N_9822);
xnor U16356 (N_16356,N_11305,N_10885);
and U16357 (N_16357,N_8983,N_12443);
nand U16358 (N_16358,N_10120,N_11568);
xnor U16359 (N_16359,N_8944,N_10117);
nor U16360 (N_16360,N_8625,N_12352);
xnor U16361 (N_16361,N_9322,N_9918);
nor U16362 (N_16362,N_11697,N_8956);
and U16363 (N_16363,N_7936,N_7417);
xor U16364 (N_16364,N_8293,N_7680);
and U16365 (N_16365,N_9735,N_8670);
nor U16366 (N_16366,N_9011,N_10900);
and U16367 (N_16367,N_9544,N_10563);
or U16368 (N_16368,N_9045,N_12189);
or U16369 (N_16369,N_9398,N_6312);
nand U16370 (N_16370,N_8991,N_11704);
nand U16371 (N_16371,N_6532,N_9951);
and U16372 (N_16372,N_9961,N_8863);
xnor U16373 (N_16373,N_11075,N_11995);
or U16374 (N_16374,N_10049,N_10477);
nand U16375 (N_16375,N_7011,N_7818);
nand U16376 (N_16376,N_7537,N_8234);
nand U16377 (N_16377,N_11101,N_7531);
and U16378 (N_16378,N_8395,N_6661);
and U16379 (N_16379,N_11833,N_8953);
or U16380 (N_16380,N_8343,N_11595);
or U16381 (N_16381,N_6402,N_12496);
xor U16382 (N_16382,N_7175,N_9784);
xor U16383 (N_16383,N_9522,N_11888);
or U16384 (N_16384,N_12317,N_6985);
nand U16385 (N_16385,N_7012,N_10146);
nor U16386 (N_16386,N_11190,N_9315);
and U16387 (N_16387,N_10894,N_8306);
nand U16388 (N_16388,N_7377,N_10279);
or U16389 (N_16389,N_12181,N_9280);
and U16390 (N_16390,N_11624,N_12331);
or U16391 (N_16391,N_10182,N_7996);
or U16392 (N_16392,N_10140,N_12379);
or U16393 (N_16393,N_6553,N_10555);
and U16394 (N_16394,N_8749,N_6674);
nand U16395 (N_16395,N_9849,N_9762);
nand U16396 (N_16396,N_7814,N_7381);
nand U16397 (N_16397,N_11345,N_12420);
or U16398 (N_16398,N_9000,N_8518);
nand U16399 (N_16399,N_8626,N_7632);
or U16400 (N_16400,N_6708,N_10744);
xor U16401 (N_16401,N_8809,N_11938);
nor U16402 (N_16402,N_9582,N_10524);
and U16403 (N_16403,N_8218,N_12066);
nor U16404 (N_16404,N_9111,N_9610);
xor U16405 (N_16405,N_6758,N_10038);
nand U16406 (N_16406,N_12070,N_8753);
or U16407 (N_16407,N_12228,N_9233);
xor U16408 (N_16408,N_8577,N_10895);
or U16409 (N_16409,N_9486,N_6937);
or U16410 (N_16410,N_11989,N_9783);
xor U16411 (N_16411,N_9811,N_8842);
nand U16412 (N_16412,N_8573,N_12425);
nand U16413 (N_16413,N_7660,N_11056);
or U16414 (N_16414,N_8097,N_11757);
nand U16415 (N_16415,N_10675,N_8020);
and U16416 (N_16416,N_9247,N_7862);
or U16417 (N_16417,N_9807,N_8113);
nand U16418 (N_16418,N_8154,N_10281);
xor U16419 (N_16419,N_11430,N_9232);
nand U16420 (N_16420,N_11988,N_6532);
or U16421 (N_16421,N_11145,N_7926);
nand U16422 (N_16422,N_7145,N_9436);
xnor U16423 (N_16423,N_7091,N_9444);
and U16424 (N_16424,N_8307,N_12341);
nor U16425 (N_16425,N_9963,N_9728);
nor U16426 (N_16426,N_11491,N_10363);
and U16427 (N_16427,N_8398,N_7874);
or U16428 (N_16428,N_10015,N_11449);
xnor U16429 (N_16429,N_11749,N_9677);
nor U16430 (N_16430,N_10695,N_10521);
nand U16431 (N_16431,N_7462,N_7615);
or U16432 (N_16432,N_8814,N_11383);
nand U16433 (N_16433,N_10412,N_10682);
or U16434 (N_16434,N_8254,N_7111);
or U16435 (N_16435,N_9534,N_7104);
and U16436 (N_16436,N_10591,N_9175);
and U16437 (N_16437,N_11705,N_10261);
nor U16438 (N_16438,N_11855,N_7323);
or U16439 (N_16439,N_9863,N_9001);
nor U16440 (N_16440,N_11363,N_11097);
xnor U16441 (N_16441,N_7827,N_8887);
or U16442 (N_16442,N_8240,N_6536);
and U16443 (N_16443,N_7355,N_11518);
xnor U16444 (N_16444,N_6715,N_10662);
or U16445 (N_16445,N_11088,N_8487);
or U16446 (N_16446,N_8072,N_6605);
and U16447 (N_16447,N_6275,N_10752);
or U16448 (N_16448,N_10563,N_7977);
nor U16449 (N_16449,N_7979,N_11220);
and U16450 (N_16450,N_9474,N_7118);
nand U16451 (N_16451,N_11282,N_10388);
and U16452 (N_16452,N_9899,N_8226);
nand U16453 (N_16453,N_7469,N_12036);
nor U16454 (N_16454,N_7346,N_11902);
nor U16455 (N_16455,N_9287,N_7840);
nand U16456 (N_16456,N_12440,N_11196);
or U16457 (N_16457,N_12247,N_6380);
nor U16458 (N_16458,N_10487,N_9833);
nand U16459 (N_16459,N_8379,N_7089);
nor U16460 (N_16460,N_7284,N_10622);
nand U16461 (N_16461,N_10638,N_8449);
and U16462 (N_16462,N_9288,N_7013);
xor U16463 (N_16463,N_10200,N_9545);
and U16464 (N_16464,N_8980,N_11311);
nor U16465 (N_16465,N_9008,N_8841);
nor U16466 (N_16466,N_6590,N_11820);
nand U16467 (N_16467,N_11034,N_9652);
nand U16468 (N_16468,N_8917,N_7833);
nor U16469 (N_16469,N_10827,N_10423);
and U16470 (N_16470,N_7185,N_11934);
xnor U16471 (N_16471,N_10663,N_6614);
nor U16472 (N_16472,N_6688,N_6715);
xor U16473 (N_16473,N_7658,N_9738);
or U16474 (N_16474,N_11689,N_10912);
or U16475 (N_16475,N_8185,N_10805);
and U16476 (N_16476,N_9511,N_11860);
xnor U16477 (N_16477,N_6989,N_11967);
or U16478 (N_16478,N_8528,N_7120);
nor U16479 (N_16479,N_11230,N_10093);
xor U16480 (N_16480,N_11587,N_11675);
nand U16481 (N_16481,N_12348,N_10736);
and U16482 (N_16482,N_6696,N_7422);
nand U16483 (N_16483,N_10876,N_11716);
nor U16484 (N_16484,N_10160,N_7983);
nor U16485 (N_16485,N_10177,N_11291);
and U16486 (N_16486,N_11682,N_11685);
nor U16487 (N_16487,N_11503,N_10123);
or U16488 (N_16488,N_11282,N_7417);
or U16489 (N_16489,N_11948,N_10984);
nand U16490 (N_16490,N_10735,N_6385);
or U16491 (N_16491,N_11457,N_7976);
or U16492 (N_16492,N_6903,N_9720);
or U16493 (N_16493,N_10490,N_9157);
or U16494 (N_16494,N_9346,N_6254);
nand U16495 (N_16495,N_11757,N_12259);
nand U16496 (N_16496,N_11405,N_11926);
nand U16497 (N_16497,N_11270,N_8520);
nor U16498 (N_16498,N_10108,N_10018);
nand U16499 (N_16499,N_7175,N_8038);
xnor U16500 (N_16500,N_7031,N_11524);
nand U16501 (N_16501,N_8974,N_12266);
xnor U16502 (N_16502,N_9696,N_11402);
xnor U16503 (N_16503,N_11997,N_9707);
or U16504 (N_16504,N_6811,N_11352);
xor U16505 (N_16505,N_9986,N_6690);
nor U16506 (N_16506,N_10795,N_11306);
xnor U16507 (N_16507,N_6305,N_9024);
and U16508 (N_16508,N_11904,N_8940);
or U16509 (N_16509,N_10867,N_12478);
or U16510 (N_16510,N_9154,N_7619);
nor U16511 (N_16511,N_7159,N_9532);
nand U16512 (N_16512,N_7263,N_10461);
nor U16513 (N_16513,N_6363,N_8218);
xnor U16514 (N_16514,N_9342,N_10310);
and U16515 (N_16515,N_8163,N_10019);
xor U16516 (N_16516,N_8125,N_9281);
xnor U16517 (N_16517,N_11513,N_10494);
nand U16518 (N_16518,N_9146,N_8797);
nand U16519 (N_16519,N_11243,N_8439);
nand U16520 (N_16520,N_8771,N_8508);
or U16521 (N_16521,N_7663,N_8747);
xor U16522 (N_16522,N_8769,N_9011);
nor U16523 (N_16523,N_9948,N_8052);
nand U16524 (N_16524,N_7550,N_12085);
xor U16525 (N_16525,N_8778,N_9014);
nand U16526 (N_16526,N_12237,N_10115);
xor U16527 (N_16527,N_9546,N_7370);
nor U16528 (N_16528,N_10363,N_9026);
and U16529 (N_16529,N_12120,N_12434);
xor U16530 (N_16530,N_9511,N_7859);
nand U16531 (N_16531,N_12255,N_11677);
and U16532 (N_16532,N_10440,N_11723);
nand U16533 (N_16533,N_8181,N_8705);
nor U16534 (N_16534,N_8375,N_9241);
nor U16535 (N_16535,N_10241,N_10057);
and U16536 (N_16536,N_6844,N_11857);
xor U16537 (N_16537,N_9484,N_6700);
xnor U16538 (N_16538,N_11681,N_8620);
xor U16539 (N_16539,N_6717,N_6323);
and U16540 (N_16540,N_7540,N_11452);
nand U16541 (N_16541,N_11266,N_10029);
and U16542 (N_16542,N_9150,N_12233);
nor U16543 (N_16543,N_8850,N_9096);
nand U16544 (N_16544,N_9125,N_8204);
nor U16545 (N_16545,N_7184,N_6415);
nand U16546 (N_16546,N_10994,N_11499);
nor U16547 (N_16547,N_6487,N_6596);
xor U16548 (N_16548,N_7510,N_8489);
and U16549 (N_16549,N_9237,N_12473);
or U16550 (N_16550,N_10748,N_8062);
or U16551 (N_16551,N_10938,N_10506);
or U16552 (N_16552,N_6692,N_12238);
and U16553 (N_16553,N_10758,N_7028);
nand U16554 (N_16554,N_8742,N_8216);
xnor U16555 (N_16555,N_11966,N_7426);
and U16556 (N_16556,N_10513,N_7838);
xor U16557 (N_16557,N_10669,N_11825);
or U16558 (N_16558,N_12377,N_9675);
nor U16559 (N_16559,N_9214,N_10380);
xor U16560 (N_16560,N_10722,N_7314);
nand U16561 (N_16561,N_9169,N_9478);
xnor U16562 (N_16562,N_9800,N_8744);
xnor U16563 (N_16563,N_8145,N_9812);
nor U16564 (N_16564,N_9558,N_8870);
or U16565 (N_16565,N_10479,N_8102);
or U16566 (N_16566,N_10630,N_6500);
nand U16567 (N_16567,N_9917,N_6567);
or U16568 (N_16568,N_10689,N_9880);
or U16569 (N_16569,N_7960,N_9593);
or U16570 (N_16570,N_10001,N_9233);
or U16571 (N_16571,N_6551,N_8660);
and U16572 (N_16572,N_8242,N_9870);
nor U16573 (N_16573,N_9942,N_8430);
nand U16574 (N_16574,N_7878,N_12133);
nand U16575 (N_16575,N_8420,N_7536);
nor U16576 (N_16576,N_8787,N_11614);
xnor U16577 (N_16577,N_7829,N_6337);
nor U16578 (N_16578,N_11494,N_8572);
or U16579 (N_16579,N_8633,N_11826);
nor U16580 (N_16580,N_7140,N_10332);
nand U16581 (N_16581,N_6722,N_11983);
nand U16582 (N_16582,N_10087,N_6727);
nand U16583 (N_16583,N_9211,N_11369);
nand U16584 (N_16584,N_10511,N_10426);
xor U16585 (N_16585,N_6360,N_9859);
and U16586 (N_16586,N_9677,N_9754);
nand U16587 (N_16587,N_9477,N_7590);
or U16588 (N_16588,N_10501,N_8462);
or U16589 (N_16589,N_6858,N_9440);
xnor U16590 (N_16590,N_10456,N_8354);
xor U16591 (N_16591,N_7787,N_10370);
nor U16592 (N_16592,N_7305,N_9018);
xor U16593 (N_16593,N_11713,N_8734);
and U16594 (N_16594,N_6440,N_6760);
or U16595 (N_16595,N_8838,N_11555);
nand U16596 (N_16596,N_10223,N_9611);
and U16597 (N_16597,N_8740,N_6296);
nor U16598 (N_16598,N_8374,N_10851);
nand U16599 (N_16599,N_7396,N_9458);
nor U16600 (N_16600,N_10971,N_11522);
xnor U16601 (N_16601,N_10191,N_10715);
and U16602 (N_16602,N_9905,N_10079);
or U16603 (N_16603,N_9263,N_8609);
nand U16604 (N_16604,N_11966,N_11497);
nor U16605 (N_16605,N_6793,N_6995);
nor U16606 (N_16606,N_8017,N_12355);
nor U16607 (N_16607,N_8735,N_12452);
or U16608 (N_16608,N_9849,N_12111);
nor U16609 (N_16609,N_12440,N_6897);
or U16610 (N_16610,N_10726,N_8294);
or U16611 (N_16611,N_7334,N_11334);
nand U16612 (N_16612,N_7523,N_10544);
or U16613 (N_16613,N_6450,N_10419);
xnor U16614 (N_16614,N_10047,N_7879);
or U16615 (N_16615,N_10239,N_6505);
or U16616 (N_16616,N_7671,N_7861);
and U16617 (N_16617,N_9333,N_11004);
and U16618 (N_16618,N_11365,N_8977);
nor U16619 (N_16619,N_6528,N_9884);
or U16620 (N_16620,N_7772,N_8092);
nor U16621 (N_16621,N_7792,N_8019);
nor U16622 (N_16622,N_7382,N_9706);
xnor U16623 (N_16623,N_7092,N_10405);
nand U16624 (N_16624,N_10885,N_9175);
nor U16625 (N_16625,N_9709,N_11223);
nand U16626 (N_16626,N_11159,N_9764);
and U16627 (N_16627,N_7519,N_8292);
or U16628 (N_16628,N_8648,N_10720);
and U16629 (N_16629,N_7809,N_6710);
or U16630 (N_16630,N_9505,N_7713);
nand U16631 (N_16631,N_10808,N_10451);
nand U16632 (N_16632,N_10219,N_6262);
or U16633 (N_16633,N_11368,N_7721);
and U16634 (N_16634,N_9456,N_9075);
xnor U16635 (N_16635,N_8501,N_7945);
nor U16636 (N_16636,N_7835,N_7112);
nand U16637 (N_16637,N_12007,N_6681);
nor U16638 (N_16638,N_7136,N_9361);
xnor U16639 (N_16639,N_8092,N_10855);
nand U16640 (N_16640,N_9484,N_6304);
xnor U16641 (N_16641,N_10970,N_7370);
nor U16642 (N_16642,N_6508,N_6981);
or U16643 (N_16643,N_8558,N_8729);
nand U16644 (N_16644,N_12009,N_9917);
xor U16645 (N_16645,N_12391,N_9165);
and U16646 (N_16646,N_8724,N_8412);
nor U16647 (N_16647,N_10863,N_8061);
or U16648 (N_16648,N_12485,N_9344);
and U16649 (N_16649,N_6287,N_9205);
or U16650 (N_16650,N_8451,N_6653);
and U16651 (N_16651,N_11895,N_10775);
nor U16652 (N_16652,N_8803,N_9342);
and U16653 (N_16653,N_10470,N_10688);
nor U16654 (N_16654,N_7980,N_6461);
nor U16655 (N_16655,N_7545,N_9888);
nor U16656 (N_16656,N_7342,N_7200);
and U16657 (N_16657,N_8116,N_6902);
xnor U16658 (N_16658,N_7470,N_8432);
nand U16659 (N_16659,N_11209,N_9283);
nor U16660 (N_16660,N_11135,N_11120);
nor U16661 (N_16661,N_9387,N_9934);
or U16662 (N_16662,N_8730,N_9754);
nand U16663 (N_16663,N_10795,N_8759);
xnor U16664 (N_16664,N_9841,N_7140);
nor U16665 (N_16665,N_8935,N_8119);
nand U16666 (N_16666,N_8518,N_9562);
and U16667 (N_16667,N_9118,N_7112);
xnor U16668 (N_16668,N_9729,N_11460);
nor U16669 (N_16669,N_8814,N_6915);
nor U16670 (N_16670,N_7174,N_8541);
nand U16671 (N_16671,N_8365,N_11723);
nor U16672 (N_16672,N_6584,N_12355);
xnor U16673 (N_16673,N_12123,N_10668);
and U16674 (N_16674,N_12246,N_9847);
xnor U16675 (N_16675,N_7668,N_11968);
and U16676 (N_16676,N_6547,N_11591);
nand U16677 (N_16677,N_11322,N_9370);
or U16678 (N_16678,N_9992,N_6794);
and U16679 (N_16679,N_9601,N_10904);
nand U16680 (N_16680,N_10263,N_10395);
and U16681 (N_16681,N_10257,N_9832);
xor U16682 (N_16682,N_10302,N_7140);
xor U16683 (N_16683,N_8069,N_6855);
nor U16684 (N_16684,N_10244,N_10209);
and U16685 (N_16685,N_6495,N_8567);
and U16686 (N_16686,N_6912,N_7829);
nor U16687 (N_16687,N_10167,N_6862);
or U16688 (N_16688,N_9193,N_10210);
or U16689 (N_16689,N_10533,N_7580);
or U16690 (N_16690,N_7117,N_9079);
nand U16691 (N_16691,N_7487,N_10060);
and U16692 (N_16692,N_11155,N_9089);
nor U16693 (N_16693,N_6704,N_9715);
nand U16694 (N_16694,N_9855,N_12058);
nor U16695 (N_16695,N_11558,N_11945);
xor U16696 (N_16696,N_11787,N_9696);
nand U16697 (N_16697,N_8517,N_12009);
or U16698 (N_16698,N_8703,N_7391);
nand U16699 (N_16699,N_9863,N_9052);
and U16700 (N_16700,N_7326,N_6320);
or U16701 (N_16701,N_10485,N_12480);
nor U16702 (N_16702,N_9135,N_9158);
nand U16703 (N_16703,N_8723,N_8675);
and U16704 (N_16704,N_10942,N_7231);
and U16705 (N_16705,N_10705,N_9878);
and U16706 (N_16706,N_8610,N_9108);
or U16707 (N_16707,N_6498,N_12093);
nor U16708 (N_16708,N_7219,N_12464);
nand U16709 (N_16709,N_7811,N_7601);
or U16710 (N_16710,N_11322,N_9943);
xnor U16711 (N_16711,N_6767,N_8546);
xor U16712 (N_16712,N_11763,N_6909);
xor U16713 (N_16713,N_8272,N_10151);
nor U16714 (N_16714,N_12496,N_10711);
or U16715 (N_16715,N_6700,N_7680);
nand U16716 (N_16716,N_8400,N_9075);
or U16717 (N_16717,N_7040,N_10993);
nor U16718 (N_16718,N_8278,N_7500);
or U16719 (N_16719,N_9030,N_9345);
and U16720 (N_16720,N_8388,N_10560);
and U16721 (N_16721,N_10530,N_7083);
xor U16722 (N_16722,N_10060,N_12149);
or U16723 (N_16723,N_8168,N_7028);
nor U16724 (N_16724,N_11202,N_11515);
and U16725 (N_16725,N_10772,N_7400);
nor U16726 (N_16726,N_9710,N_6982);
and U16727 (N_16727,N_9861,N_8446);
nor U16728 (N_16728,N_7109,N_10666);
and U16729 (N_16729,N_7956,N_7885);
or U16730 (N_16730,N_12012,N_10078);
xor U16731 (N_16731,N_10849,N_6340);
xor U16732 (N_16732,N_10790,N_7594);
nor U16733 (N_16733,N_10271,N_10798);
nor U16734 (N_16734,N_9851,N_10608);
nand U16735 (N_16735,N_11941,N_6737);
nor U16736 (N_16736,N_8172,N_12385);
or U16737 (N_16737,N_7883,N_7177);
nor U16738 (N_16738,N_8271,N_6563);
nand U16739 (N_16739,N_8888,N_9288);
and U16740 (N_16740,N_7978,N_6748);
nor U16741 (N_16741,N_6287,N_11629);
nor U16742 (N_16742,N_11869,N_9233);
nor U16743 (N_16743,N_7006,N_11075);
nand U16744 (N_16744,N_6804,N_8191);
nor U16745 (N_16745,N_11151,N_9103);
or U16746 (N_16746,N_6773,N_8387);
xor U16747 (N_16747,N_9815,N_11402);
and U16748 (N_16748,N_8371,N_10153);
and U16749 (N_16749,N_9283,N_11373);
xnor U16750 (N_16750,N_9104,N_6557);
and U16751 (N_16751,N_6550,N_9871);
and U16752 (N_16752,N_6874,N_6379);
nor U16753 (N_16753,N_6572,N_11044);
nand U16754 (N_16754,N_7318,N_9561);
or U16755 (N_16755,N_10323,N_11435);
xor U16756 (N_16756,N_8878,N_10514);
nor U16757 (N_16757,N_12459,N_7528);
and U16758 (N_16758,N_10385,N_10807);
and U16759 (N_16759,N_11418,N_9815);
nand U16760 (N_16760,N_7722,N_9501);
xor U16761 (N_16761,N_7742,N_11637);
and U16762 (N_16762,N_12428,N_9621);
and U16763 (N_16763,N_11443,N_8011);
or U16764 (N_16764,N_8165,N_7441);
and U16765 (N_16765,N_6843,N_11744);
nor U16766 (N_16766,N_6453,N_12364);
and U16767 (N_16767,N_7544,N_11315);
xnor U16768 (N_16768,N_12034,N_6957);
xor U16769 (N_16769,N_10769,N_12051);
and U16770 (N_16770,N_10202,N_6375);
or U16771 (N_16771,N_11006,N_8767);
nand U16772 (N_16772,N_11424,N_8138);
and U16773 (N_16773,N_11087,N_10989);
nor U16774 (N_16774,N_11724,N_9547);
or U16775 (N_16775,N_6299,N_9633);
xnor U16776 (N_16776,N_7527,N_9693);
and U16777 (N_16777,N_11921,N_7186);
and U16778 (N_16778,N_12121,N_7195);
and U16779 (N_16779,N_9978,N_9602);
and U16780 (N_16780,N_7360,N_10090);
nand U16781 (N_16781,N_10789,N_12158);
or U16782 (N_16782,N_8208,N_8821);
or U16783 (N_16783,N_6440,N_10501);
nand U16784 (N_16784,N_9859,N_6631);
and U16785 (N_16785,N_7454,N_7921);
or U16786 (N_16786,N_10882,N_7039);
xnor U16787 (N_16787,N_12235,N_12448);
nand U16788 (N_16788,N_11272,N_9909);
xnor U16789 (N_16789,N_7848,N_8179);
nor U16790 (N_16790,N_7739,N_9725);
and U16791 (N_16791,N_7567,N_12333);
or U16792 (N_16792,N_10063,N_11268);
xnor U16793 (N_16793,N_8283,N_9463);
or U16794 (N_16794,N_11511,N_10653);
nor U16795 (N_16795,N_7344,N_10369);
nor U16796 (N_16796,N_10844,N_10503);
and U16797 (N_16797,N_9883,N_11188);
nand U16798 (N_16798,N_11605,N_6501);
xor U16799 (N_16799,N_10400,N_6976);
nand U16800 (N_16800,N_10550,N_7400);
nand U16801 (N_16801,N_9876,N_10909);
and U16802 (N_16802,N_11692,N_8840);
nor U16803 (N_16803,N_8185,N_10119);
or U16804 (N_16804,N_8898,N_10538);
or U16805 (N_16805,N_10274,N_8373);
nor U16806 (N_16806,N_12362,N_9218);
and U16807 (N_16807,N_10576,N_11545);
nor U16808 (N_16808,N_9177,N_8548);
or U16809 (N_16809,N_11636,N_8668);
nor U16810 (N_16810,N_11648,N_11069);
and U16811 (N_16811,N_7179,N_8708);
xor U16812 (N_16812,N_9435,N_10878);
or U16813 (N_16813,N_6561,N_11740);
xnor U16814 (N_16814,N_9015,N_8131);
xnor U16815 (N_16815,N_8681,N_6397);
and U16816 (N_16816,N_7507,N_11290);
xnor U16817 (N_16817,N_7839,N_11827);
and U16818 (N_16818,N_8239,N_10227);
and U16819 (N_16819,N_12262,N_8945);
nand U16820 (N_16820,N_8144,N_7419);
xor U16821 (N_16821,N_8789,N_11835);
and U16822 (N_16822,N_11462,N_8561);
nand U16823 (N_16823,N_9266,N_8458);
nand U16824 (N_16824,N_12467,N_9214);
and U16825 (N_16825,N_12171,N_6677);
and U16826 (N_16826,N_6633,N_11863);
or U16827 (N_16827,N_7461,N_8987);
nand U16828 (N_16828,N_8493,N_7319);
xnor U16829 (N_16829,N_7426,N_12377);
or U16830 (N_16830,N_11980,N_8134);
xor U16831 (N_16831,N_6991,N_10813);
or U16832 (N_16832,N_8944,N_9197);
xor U16833 (N_16833,N_7606,N_6838);
nand U16834 (N_16834,N_9015,N_10263);
nand U16835 (N_16835,N_8883,N_7678);
or U16836 (N_16836,N_9784,N_11764);
nand U16837 (N_16837,N_12342,N_10286);
or U16838 (N_16838,N_8073,N_12321);
and U16839 (N_16839,N_6275,N_10841);
or U16840 (N_16840,N_10704,N_7969);
or U16841 (N_16841,N_11801,N_7978);
nand U16842 (N_16842,N_6588,N_9612);
nor U16843 (N_16843,N_8903,N_9481);
nand U16844 (N_16844,N_7426,N_10938);
or U16845 (N_16845,N_12441,N_12019);
nor U16846 (N_16846,N_8127,N_8680);
nand U16847 (N_16847,N_11683,N_6872);
or U16848 (N_16848,N_10834,N_9378);
or U16849 (N_16849,N_6501,N_7971);
xnor U16850 (N_16850,N_8357,N_12142);
or U16851 (N_16851,N_7481,N_10482);
nand U16852 (N_16852,N_7074,N_6577);
nor U16853 (N_16853,N_10098,N_7045);
and U16854 (N_16854,N_6454,N_10388);
or U16855 (N_16855,N_10747,N_11707);
and U16856 (N_16856,N_8099,N_10438);
xnor U16857 (N_16857,N_6332,N_11655);
nor U16858 (N_16858,N_11431,N_12469);
nor U16859 (N_16859,N_10073,N_8802);
xnor U16860 (N_16860,N_10582,N_9338);
or U16861 (N_16861,N_12487,N_10468);
nand U16862 (N_16862,N_9675,N_12097);
or U16863 (N_16863,N_6961,N_10096);
or U16864 (N_16864,N_7340,N_11292);
or U16865 (N_16865,N_8162,N_9953);
nand U16866 (N_16866,N_11752,N_8271);
xor U16867 (N_16867,N_12214,N_7689);
nand U16868 (N_16868,N_12034,N_11759);
nor U16869 (N_16869,N_7576,N_7481);
xor U16870 (N_16870,N_10208,N_9737);
or U16871 (N_16871,N_6251,N_7139);
and U16872 (N_16872,N_6963,N_10248);
nand U16873 (N_16873,N_6625,N_7530);
nand U16874 (N_16874,N_8989,N_11992);
nor U16875 (N_16875,N_8345,N_7612);
nand U16876 (N_16876,N_11736,N_7022);
and U16877 (N_16877,N_7072,N_11736);
and U16878 (N_16878,N_9303,N_7386);
nand U16879 (N_16879,N_10065,N_12388);
and U16880 (N_16880,N_12241,N_9577);
nand U16881 (N_16881,N_9569,N_9433);
and U16882 (N_16882,N_11821,N_6493);
xnor U16883 (N_16883,N_11171,N_11524);
nand U16884 (N_16884,N_6844,N_9599);
nor U16885 (N_16885,N_10025,N_12050);
or U16886 (N_16886,N_12345,N_10673);
and U16887 (N_16887,N_10624,N_10384);
or U16888 (N_16888,N_6776,N_8155);
nand U16889 (N_16889,N_12433,N_11922);
nor U16890 (N_16890,N_6803,N_6417);
and U16891 (N_16891,N_10866,N_10857);
nor U16892 (N_16892,N_8549,N_11037);
nor U16893 (N_16893,N_6724,N_7143);
and U16894 (N_16894,N_6507,N_8375);
nand U16895 (N_16895,N_11685,N_11136);
nor U16896 (N_16896,N_11907,N_9738);
or U16897 (N_16897,N_9269,N_9133);
nor U16898 (N_16898,N_7827,N_10728);
nor U16899 (N_16899,N_10913,N_10060);
or U16900 (N_16900,N_10086,N_8226);
or U16901 (N_16901,N_10968,N_6425);
nand U16902 (N_16902,N_7938,N_12458);
nor U16903 (N_16903,N_9734,N_7626);
nand U16904 (N_16904,N_6436,N_10750);
and U16905 (N_16905,N_8204,N_7201);
or U16906 (N_16906,N_10312,N_6531);
nand U16907 (N_16907,N_6389,N_7082);
or U16908 (N_16908,N_12121,N_9090);
nand U16909 (N_16909,N_10819,N_7307);
nor U16910 (N_16910,N_10397,N_7163);
nor U16911 (N_16911,N_10893,N_10528);
or U16912 (N_16912,N_8724,N_6557);
nand U16913 (N_16913,N_10294,N_7460);
or U16914 (N_16914,N_6359,N_12192);
nand U16915 (N_16915,N_11315,N_11003);
xor U16916 (N_16916,N_9603,N_10968);
nand U16917 (N_16917,N_6379,N_9621);
xor U16918 (N_16918,N_10390,N_6628);
or U16919 (N_16919,N_8578,N_11050);
and U16920 (N_16920,N_10952,N_11582);
or U16921 (N_16921,N_6994,N_6871);
or U16922 (N_16922,N_7679,N_10470);
xor U16923 (N_16923,N_6467,N_7997);
nor U16924 (N_16924,N_10575,N_12082);
xor U16925 (N_16925,N_10100,N_9140);
and U16926 (N_16926,N_10378,N_7230);
or U16927 (N_16927,N_11029,N_6951);
or U16928 (N_16928,N_12041,N_9969);
or U16929 (N_16929,N_8743,N_12318);
xor U16930 (N_16930,N_8665,N_6325);
xnor U16931 (N_16931,N_7114,N_11070);
nand U16932 (N_16932,N_9287,N_7270);
and U16933 (N_16933,N_11918,N_11302);
nor U16934 (N_16934,N_11213,N_7352);
xor U16935 (N_16935,N_12191,N_7173);
and U16936 (N_16936,N_9912,N_9372);
nor U16937 (N_16937,N_6792,N_11815);
nand U16938 (N_16938,N_10891,N_7748);
nand U16939 (N_16939,N_8419,N_10474);
nand U16940 (N_16940,N_6997,N_11413);
or U16941 (N_16941,N_10160,N_11207);
nand U16942 (N_16942,N_11383,N_9037);
nand U16943 (N_16943,N_10838,N_10270);
nor U16944 (N_16944,N_7758,N_11766);
nor U16945 (N_16945,N_12484,N_7695);
and U16946 (N_16946,N_12141,N_7306);
xnor U16947 (N_16947,N_7881,N_11573);
nor U16948 (N_16948,N_7002,N_7255);
and U16949 (N_16949,N_8347,N_6692);
nor U16950 (N_16950,N_12044,N_9842);
nor U16951 (N_16951,N_10631,N_9120);
xnor U16952 (N_16952,N_7750,N_11327);
nand U16953 (N_16953,N_7160,N_8401);
nand U16954 (N_16954,N_6784,N_6513);
nor U16955 (N_16955,N_11790,N_8895);
nor U16956 (N_16956,N_11631,N_12043);
or U16957 (N_16957,N_9947,N_9820);
nand U16958 (N_16958,N_9540,N_11458);
nor U16959 (N_16959,N_11325,N_6252);
and U16960 (N_16960,N_8841,N_7783);
xnor U16961 (N_16961,N_10196,N_11878);
nand U16962 (N_16962,N_12312,N_8044);
or U16963 (N_16963,N_7263,N_10270);
or U16964 (N_16964,N_11847,N_6908);
xor U16965 (N_16965,N_8877,N_9616);
nor U16966 (N_16966,N_7251,N_7450);
nand U16967 (N_16967,N_7214,N_11860);
nor U16968 (N_16968,N_8149,N_9217);
or U16969 (N_16969,N_11261,N_7662);
and U16970 (N_16970,N_7612,N_11636);
nand U16971 (N_16971,N_8149,N_10496);
nand U16972 (N_16972,N_9328,N_12160);
xor U16973 (N_16973,N_11670,N_7763);
nor U16974 (N_16974,N_6281,N_6466);
xnor U16975 (N_16975,N_8168,N_10934);
and U16976 (N_16976,N_9975,N_6801);
nand U16977 (N_16977,N_8522,N_6329);
nand U16978 (N_16978,N_8053,N_9331);
and U16979 (N_16979,N_10231,N_6851);
and U16980 (N_16980,N_7781,N_9469);
nand U16981 (N_16981,N_10937,N_6309);
or U16982 (N_16982,N_8143,N_12258);
xor U16983 (N_16983,N_11430,N_11301);
nor U16984 (N_16984,N_11132,N_7233);
nand U16985 (N_16985,N_7369,N_11697);
and U16986 (N_16986,N_11927,N_7236);
nor U16987 (N_16987,N_8081,N_11473);
nand U16988 (N_16988,N_8124,N_6570);
nor U16989 (N_16989,N_11693,N_6676);
xnor U16990 (N_16990,N_6878,N_7844);
nor U16991 (N_16991,N_11928,N_9173);
and U16992 (N_16992,N_11564,N_10987);
nor U16993 (N_16993,N_10138,N_10778);
and U16994 (N_16994,N_10361,N_7111);
xnor U16995 (N_16995,N_11724,N_6300);
xor U16996 (N_16996,N_11484,N_7314);
nor U16997 (N_16997,N_10819,N_8444);
nor U16998 (N_16998,N_11810,N_12456);
nand U16999 (N_16999,N_8570,N_12019);
or U17000 (N_17000,N_11546,N_7674);
nand U17001 (N_17001,N_12162,N_12016);
and U17002 (N_17002,N_12464,N_9979);
or U17003 (N_17003,N_7648,N_10260);
and U17004 (N_17004,N_10304,N_8016);
xnor U17005 (N_17005,N_10510,N_11339);
nand U17006 (N_17006,N_9153,N_10725);
nor U17007 (N_17007,N_11486,N_10502);
nor U17008 (N_17008,N_9176,N_8143);
nor U17009 (N_17009,N_9737,N_8053);
or U17010 (N_17010,N_8437,N_6647);
and U17011 (N_17011,N_9411,N_7821);
nand U17012 (N_17012,N_6913,N_10784);
or U17013 (N_17013,N_8269,N_8725);
and U17014 (N_17014,N_8428,N_7453);
nor U17015 (N_17015,N_8299,N_8787);
nor U17016 (N_17016,N_6897,N_6422);
xor U17017 (N_17017,N_7224,N_8686);
and U17018 (N_17018,N_7251,N_8930);
and U17019 (N_17019,N_11613,N_9810);
nand U17020 (N_17020,N_11236,N_6313);
nand U17021 (N_17021,N_6777,N_7458);
xor U17022 (N_17022,N_8399,N_9999);
nor U17023 (N_17023,N_10839,N_8088);
or U17024 (N_17024,N_9830,N_10909);
nor U17025 (N_17025,N_9477,N_8649);
or U17026 (N_17026,N_8082,N_9340);
and U17027 (N_17027,N_11054,N_8024);
or U17028 (N_17028,N_9854,N_8583);
nand U17029 (N_17029,N_10691,N_8769);
nand U17030 (N_17030,N_11726,N_9073);
or U17031 (N_17031,N_9014,N_8060);
nand U17032 (N_17032,N_11642,N_11843);
or U17033 (N_17033,N_6946,N_9210);
nor U17034 (N_17034,N_10404,N_6825);
xor U17035 (N_17035,N_9664,N_6917);
nand U17036 (N_17036,N_11732,N_6544);
nand U17037 (N_17037,N_9550,N_9903);
and U17038 (N_17038,N_12022,N_6463);
nand U17039 (N_17039,N_7820,N_10172);
nand U17040 (N_17040,N_6398,N_9635);
or U17041 (N_17041,N_12237,N_11738);
xnor U17042 (N_17042,N_7256,N_8162);
nand U17043 (N_17043,N_10863,N_8482);
nand U17044 (N_17044,N_8156,N_6478);
nor U17045 (N_17045,N_12499,N_8634);
nand U17046 (N_17046,N_8923,N_12369);
nor U17047 (N_17047,N_8709,N_11106);
nor U17048 (N_17048,N_10018,N_7777);
or U17049 (N_17049,N_12043,N_6307);
nand U17050 (N_17050,N_9442,N_7775);
xor U17051 (N_17051,N_10304,N_10112);
and U17052 (N_17052,N_10370,N_8469);
xor U17053 (N_17053,N_9307,N_9313);
xor U17054 (N_17054,N_8326,N_6463);
or U17055 (N_17055,N_10978,N_6945);
or U17056 (N_17056,N_12217,N_9937);
or U17057 (N_17057,N_10747,N_8874);
xor U17058 (N_17058,N_10034,N_8616);
nand U17059 (N_17059,N_6680,N_7767);
and U17060 (N_17060,N_7386,N_8677);
nand U17061 (N_17061,N_9187,N_9176);
xnor U17062 (N_17062,N_6633,N_6738);
xor U17063 (N_17063,N_7665,N_12313);
and U17064 (N_17064,N_8050,N_10521);
xor U17065 (N_17065,N_7436,N_9377);
nor U17066 (N_17066,N_8234,N_7773);
nand U17067 (N_17067,N_6421,N_12393);
nor U17068 (N_17068,N_10665,N_9472);
and U17069 (N_17069,N_12158,N_9560);
and U17070 (N_17070,N_11594,N_7526);
xnor U17071 (N_17071,N_7818,N_11978);
xor U17072 (N_17072,N_7709,N_6332);
nand U17073 (N_17073,N_10383,N_7764);
xor U17074 (N_17074,N_11431,N_6681);
or U17075 (N_17075,N_8408,N_7804);
xnor U17076 (N_17076,N_8630,N_9093);
xnor U17077 (N_17077,N_10298,N_11446);
xnor U17078 (N_17078,N_6818,N_7728);
nand U17079 (N_17079,N_11218,N_6988);
nand U17080 (N_17080,N_12466,N_6655);
nand U17081 (N_17081,N_10409,N_9763);
and U17082 (N_17082,N_6912,N_6819);
and U17083 (N_17083,N_10700,N_10196);
or U17084 (N_17084,N_12054,N_12176);
xor U17085 (N_17085,N_9542,N_10281);
nand U17086 (N_17086,N_10471,N_6868);
and U17087 (N_17087,N_11964,N_8951);
nor U17088 (N_17088,N_10767,N_11599);
xnor U17089 (N_17089,N_7966,N_9113);
nand U17090 (N_17090,N_11295,N_9526);
or U17091 (N_17091,N_9931,N_7604);
or U17092 (N_17092,N_11785,N_7407);
and U17093 (N_17093,N_8683,N_8089);
nand U17094 (N_17094,N_9937,N_11266);
nand U17095 (N_17095,N_11006,N_7268);
or U17096 (N_17096,N_10954,N_7915);
and U17097 (N_17097,N_8265,N_7409);
xnor U17098 (N_17098,N_9842,N_9747);
and U17099 (N_17099,N_8220,N_12015);
xor U17100 (N_17100,N_9263,N_7568);
and U17101 (N_17101,N_6879,N_7608);
xnor U17102 (N_17102,N_8652,N_7425);
or U17103 (N_17103,N_9493,N_10885);
nand U17104 (N_17104,N_9514,N_9675);
nor U17105 (N_17105,N_9059,N_6715);
xor U17106 (N_17106,N_6941,N_9436);
and U17107 (N_17107,N_7424,N_11261);
nor U17108 (N_17108,N_10799,N_8696);
and U17109 (N_17109,N_11089,N_7509);
xnor U17110 (N_17110,N_10694,N_8676);
or U17111 (N_17111,N_7602,N_9787);
or U17112 (N_17112,N_7917,N_10090);
nor U17113 (N_17113,N_9856,N_6488);
nand U17114 (N_17114,N_8323,N_8363);
or U17115 (N_17115,N_9064,N_7781);
or U17116 (N_17116,N_7388,N_10827);
xnor U17117 (N_17117,N_9468,N_9375);
nand U17118 (N_17118,N_6354,N_8169);
nor U17119 (N_17119,N_10529,N_9464);
and U17120 (N_17120,N_6572,N_10557);
nor U17121 (N_17121,N_10402,N_10121);
or U17122 (N_17122,N_8986,N_8538);
or U17123 (N_17123,N_10596,N_11586);
xnor U17124 (N_17124,N_9837,N_6926);
or U17125 (N_17125,N_8932,N_10057);
nand U17126 (N_17126,N_6253,N_8037);
nor U17127 (N_17127,N_10921,N_9907);
or U17128 (N_17128,N_11204,N_6677);
nand U17129 (N_17129,N_12228,N_9370);
nand U17130 (N_17130,N_7375,N_11147);
xnor U17131 (N_17131,N_12012,N_9303);
xnor U17132 (N_17132,N_10617,N_10900);
xnor U17133 (N_17133,N_11040,N_6918);
or U17134 (N_17134,N_6848,N_8325);
and U17135 (N_17135,N_8787,N_9559);
and U17136 (N_17136,N_9652,N_7650);
nand U17137 (N_17137,N_7745,N_7558);
nor U17138 (N_17138,N_10358,N_10028);
and U17139 (N_17139,N_9867,N_7709);
nor U17140 (N_17140,N_10074,N_7216);
nor U17141 (N_17141,N_7761,N_9838);
xnor U17142 (N_17142,N_12407,N_11312);
xnor U17143 (N_17143,N_9559,N_11792);
or U17144 (N_17144,N_7633,N_10724);
or U17145 (N_17145,N_10368,N_8067);
and U17146 (N_17146,N_12296,N_9328);
xnor U17147 (N_17147,N_10859,N_8854);
nor U17148 (N_17148,N_6498,N_12475);
xnor U17149 (N_17149,N_10897,N_9429);
nor U17150 (N_17150,N_6333,N_9899);
nand U17151 (N_17151,N_10877,N_8537);
xnor U17152 (N_17152,N_9247,N_9170);
nand U17153 (N_17153,N_11598,N_10558);
and U17154 (N_17154,N_11019,N_12046);
or U17155 (N_17155,N_12018,N_9983);
and U17156 (N_17156,N_11224,N_11022);
nor U17157 (N_17157,N_9035,N_9140);
xor U17158 (N_17158,N_12227,N_6742);
and U17159 (N_17159,N_10291,N_8295);
and U17160 (N_17160,N_7730,N_6675);
or U17161 (N_17161,N_10846,N_7444);
nand U17162 (N_17162,N_9520,N_8510);
nand U17163 (N_17163,N_11620,N_7601);
or U17164 (N_17164,N_11985,N_10197);
nand U17165 (N_17165,N_8963,N_6895);
and U17166 (N_17166,N_8882,N_6854);
and U17167 (N_17167,N_9682,N_7024);
or U17168 (N_17168,N_12135,N_9312);
or U17169 (N_17169,N_10346,N_6936);
and U17170 (N_17170,N_8951,N_10838);
xor U17171 (N_17171,N_8597,N_7458);
nand U17172 (N_17172,N_8412,N_10837);
nand U17173 (N_17173,N_6330,N_11997);
and U17174 (N_17174,N_10980,N_9117);
nor U17175 (N_17175,N_8274,N_9324);
nand U17176 (N_17176,N_9421,N_8459);
or U17177 (N_17177,N_7302,N_7222);
nand U17178 (N_17178,N_7802,N_8953);
or U17179 (N_17179,N_10725,N_12248);
nor U17180 (N_17180,N_12167,N_11507);
nor U17181 (N_17181,N_10814,N_6251);
or U17182 (N_17182,N_8812,N_11775);
and U17183 (N_17183,N_9433,N_7140);
or U17184 (N_17184,N_7322,N_11018);
nor U17185 (N_17185,N_10189,N_9225);
xnor U17186 (N_17186,N_10480,N_8591);
or U17187 (N_17187,N_11528,N_7090);
or U17188 (N_17188,N_7030,N_11559);
or U17189 (N_17189,N_11546,N_9212);
xnor U17190 (N_17190,N_8895,N_11603);
nand U17191 (N_17191,N_7366,N_8573);
nand U17192 (N_17192,N_10322,N_6646);
nor U17193 (N_17193,N_9725,N_7514);
nand U17194 (N_17194,N_8993,N_7512);
and U17195 (N_17195,N_9214,N_8209);
xnor U17196 (N_17196,N_6567,N_10160);
nor U17197 (N_17197,N_8981,N_6824);
or U17198 (N_17198,N_9044,N_11642);
nor U17199 (N_17199,N_12114,N_11749);
xor U17200 (N_17200,N_7665,N_8654);
xnor U17201 (N_17201,N_7923,N_10370);
nor U17202 (N_17202,N_6664,N_7648);
and U17203 (N_17203,N_8358,N_6703);
and U17204 (N_17204,N_11622,N_10026);
nor U17205 (N_17205,N_6354,N_11492);
nor U17206 (N_17206,N_11074,N_11024);
nand U17207 (N_17207,N_7268,N_9035);
and U17208 (N_17208,N_6880,N_9266);
nor U17209 (N_17209,N_11200,N_10066);
nand U17210 (N_17210,N_7498,N_9060);
xor U17211 (N_17211,N_9303,N_8628);
nor U17212 (N_17212,N_8597,N_11329);
nand U17213 (N_17213,N_7319,N_12242);
or U17214 (N_17214,N_8457,N_9130);
and U17215 (N_17215,N_9705,N_7901);
xnor U17216 (N_17216,N_10601,N_11970);
nor U17217 (N_17217,N_10197,N_6280);
or U17218 (N_17218,N_8882,N_12320);
nand U17219 (N_17219,N_12094,N_9100);
or U17220 (N_17220,N_11178,N_7688);
nand U17221 (N_17221,N_9446,N_10776);
nor U17222 (N_17222,N_11038,N_6715);
nand U17223 (N_17223,N_12420,N_7709);
nand U17224 (N_17224,N_11657,N_10794);
xnor U17225 (N_17225,N_7782,N_8041);
and U17226 (N_17226,N_7923,N_11652);
nand U17227 (N_17227,N_12414,N_6409);
nor U17228 (N_17228,N_7756,N_11727);
nor U17229 (N_17229,N_9119,N_8080);
nand U17230 (N_17230,N_9510,N_9154);
nor U17231 (N_17231,N_10402,N_10149);
xnor U17232 (N_17232,N_11054,N_6710);
xor U17233 (N_17233,N_6803,N_7663);
and U17234 (N_17234,N_12428,N_9092);
nor U17235 (N_17235,N_9503,N_10181);
xnor U17236 (N_17236,N_10289,N_8415);
and U17237 (N_17237,N_11966,N_9037);
and U17238 (N_17238,N_10643,N_6473);
xor U17239 (N_17239,N_7311,N_9370);
xor U17240 (N_17240,N_10269,N_11176);
nand U17241 (N_17241,N_6715,N_8159);
nor U17242 (N_17242,N_11119,N_9529);
xor U17243 (N_17243,N_9748,N_9166);
and U17244 (N_17244,N_9902,N_8086);
or U17245 (N_17245,N_11205,N_8941);
or U17246 (N_17246,N_6431,N_8470);
or U17247 (N_17247,N_7286,N_7227);
and U17248 (N_17248,N_8576,N_12452);
and U17249 (N_17249,N_7757,N_10691);
or U17250 (N_17250,N_9437,N_12450);
nand U17251 (N_17251,N_7775,N_10570);
or U17252 (N_17252,N_9118,N_6857);
nor U17253 (N_17253,N_8524,N_12206);
nand U17254 (N_17254,N_7744,N_8619);
and U17255 (N_17255,N_6945,N_11630);
nand U17256 (N_17256,N_9665,N_11004);
and U17257 (N_17257,N_9326,N_6342);
nand U17258 (N_17258,N_10023,N_10102);
nand U17259 (N_17259,N_6437,N_7092);
and U17260 (N_17260,N_7197,N_11338);
nand U17261 (N_17261,N_9220,N_7183);
and U17262 (N_17262,N_10083,N_10202);
nor U17263 (N_17263,N_11520,N_7807);
or U17264 (N_17264,N_11584,N_8956);
nor U17265 (N_17265,N_9936,N_10686);
xnor U17266 (N_17266,N_6721,N_8373);
or U17267 (N_17267,N_6924,N_10643);
nand U17268 (N_17268,N_7511,N_11975);
nor U17269 (N_17269,N_7436,N_8491);
and U17270 (N_17270,N_6307,N_8211);
or U17271 (N_17271,N_7147,N_8256);
and U17272 (N_17272,N_9387,N_8835);
nor U17273 (N_17273,N_8939,N_7898);
xor U17274 (N_17274,N_9280,N_9593);
nand U17275 (N_17275,N_9324,N_12216);
and U17276 (N_17276,N_8567,N_6816);
xor U17277 (N_17277,N_10459,N_9596);
xnor U17278 (N_17278,N_7738,N_9558);
or U17279 (N_17279,N_9421,N_11122);
or U17280 (N_17280,N_6704,N_9652);
and U17281 (N_17281,N_8808,N_9559);
or U17282 (N_17282,N_11346,N_6878);
and U17283 (N_17283,N_10544,N_12477);
and U17284 (N_17284,N_6353,N_10115);
or U17285 (N_17285,N_11591,N_7697);
and U17286 (N_17286,N_6307,N_11318);
xnor U17287 (N_17287,N_8658,N_8761);
and U17288 (N_17288,N_8614,N_9346);
or U17289 (N_17289,N_6762,N_12177);
nor U17290 (N_17290,N_8410,N_7379);
or U17291 (N_17291,N_8972,N_9327);
or U17292 (N_17292,N_10230,N_11837);
xnor U17293 (N_17293,N_12030,N_11326);
nor U17294 (N_17294,N_10560,N_11493);
nor U17295 (N_17295,N_11452,N_7202);
or U17296 (N_17296,N_11467,N_6423);
xor U17297 (N_17297,N_11932,N_9279);
nand U17298 (N_17298,N_8723,N_9343);
and U17299 (N_17299,N_11656,N_12484);
nor U17300 (N_17300,N_8339,N_8574);
nor U17301 (N_17301,N_8665,N_11300);
nor U17302 (N_17302,N_9806,N_8036);
xor U17303 (N_17303,N_8063,N_10856);
xnor U17304 (N_17304,N_10976,N_11614);
and U17305 (N_17305,N_7928,N_8468);
nor U17306 (N_17306,N_10196,N_10455);
and U17307 (N_17307,N_11441,N_10603);
nand U17308 (N_17308,N_7108,N_7587);
and U17309 (N_17309,N_8210,N_6493);
nand U17310 (N_17310,N_9499,N_9883);
and U17311 (N_17311,N_7231,N_11601);
nor U17312 (N_17312,N_11424,N_8028);
and U17313 (N_17313,N_9913,N_10652);
and U17314 (N_17314,N_11864,N_12494);
nand U17315 (N_17315,N_6929,N_8627);
nand U17316 (N_17316,N_6719,N_9282);
nand U17317 (N_17317,N_7534,N_12346);
nand U17318 (N_17318,N_10532,N_8381);
nand U17319 (N_17319,N_9187,N_6874);
xnor U17320 (N_17320,N_9327,N_8593);
nand U17321 (N_17321,N_11624,N_10562);
or U17322 (N_17322,N_10393,N_10995);
and U17323 (N_17323,N_9913,N_7956);
nor U17324 (N_17324,N_7483,N_8222);
nor U17325 (N_17325,N_11382,N_12034);
nor U17326 (N_17326,N_12081,N_9401);
xnor U17327 (N_17327,N_6296,N_6362);
nor U17328 (N_17328,N_11492,N_11741);
nand U17329 (N_17329,N_12347,N_8443);
or U17330 (N_17330,N_7513,N_6743);
xnor U17331 (N_17331,N_6936,N_12044);
and U17332 (N_17332,N_7445,N_8003);
nand U17333 (N_17333,N_11636,N_11683);
nand U17334 (N_17334,N_11395,N_8073);
or U17335 (N_17335,N_9237,N_7135);
nor U17336 (N_17336,N_7669,N_11293);
xnor U17337 (N_17337,N_6430,N_7224);
or U17338 (N_17338,N_10940,N_8743);
nand U17339 (N_17339,N_10458,N_9993);
nor U17340 (N_17340,N_9663,N_6633);
nor U17341 (N_17341,N_7179,N_9699);
or U17342 (N_17342,N_8560,N_8090);
nor U17343 (N_17343,N_12472,N_7661);
nor U17344 (N_17344,N_12341,N_12171);
and U17345 (N_17345,N_10195,N_7721);
nand U17346 (N_17346,N_10594,N_8848);
and U17347 (N_17347,N_9054,N_12495);
xnor U17348 (N_17348,N_8202,N_6457);
nor U17349 (N_17349,N_11350,N_10239);
or U17350 (N_17350,N_11460,N_6471);
or U17351 (N_17351,N_11455,N_7115);
nor U17352 (N_17352,N_8705,N_7752);
xor U17353 (N_17353,N_8096,N_9917);
nor U17354 (N_17354,N_11406,N_6827);
or U17355 (N_17355,N_7109,N_10173);
or U17356 (N_17356,N_12015,N_8748);
nand U17357 (N_17357,N_12010,N_9852);
nand U17358 (N_17358,N_11123,N_10016);
xor U17359 (N_17359,N_9418,N_8328);
nand U17360 (N_17360,N_7864,N_10108);
and U17361 (N_17361,N_7315,N_6482);
or U17362 (N_17362,N_9197,N_7873);
xnor U17363 (N_17363,N_6875,N_10154);
nand U17364 (N_17364,N_11050,N_12163);
or U17365 (N_17365,N_10530,N_8427);
nor U17366 (N_17366,N_7149,N_6519);
or U17367 (N_17367,N_10674,N_9856);
or U17368 (N_17368,N_10803,N_6870);
and U17369 (N_17369,N_11687,N_8933);
and U17370 (N_17370,N_8168,N_8807);
nand U17371 (N_17371,N_6283,N_11118);
nand U17372 (N_17372,N_7837,N_8116);
nand U17373 (N_17373,N_8423,N_12030);
and U17374 (N_17374,N_11070,N_9969);
nor U17375 (N_17375,N_11472,N_8178);
nand U17376 (N_17376,N_9468,N_6270);
or U17377 (N_17377,N_7749,N_6761);
and U17378 (N_17378,N_12415,N_10285);
xnor U17379 (N_17379,N_6563,N_9410);
or U17380 (N_17380,N_8439,N_8967);
or U17381 (N_17381,N_7340,N_11054);
xor U17382 (N_17382,N_8674,N_8315);
nand U17383 (N_17383,N_9751,N_8853);
xor U17384 (N_17384,N_10350,N_8137);
or U17385 (N_17385,N_10902,N_12282);
nand U17386 (N_17386,N_11876,N_7444);
nor U17387 (N_17387,N_6879,N_7275);
xnor U17388 (N_17388,N_8167,N_8189);
nor U17389 (N_17389,N_11352,N_10082);
and U17390 (N_17390,N_10629,N_11793);
nand U17391 (N_17391,N_11645,N_9481);
nand U17392 (N_17392,N_6665,N_9923);
nor U17393 (N_17393,N_9185,N_6478);
xnor U17394 (N_17394,N_8479,N_6275);
nor U17395 (N_17395,N_12196,N_12199);
and U17396 (N_17396,N_7716,N_11495);
nor U17397 (N_17397,N_10836,N_6272);
nor U17398 (N_17398,N_9092,N_9854);
nand U17399 (N_17399,N_10046,N_7602);
and U17400 (N_17400,N_6514,N_10156);
nand U17401 (N_17401,N_7273,N_11071);
and U17402 (N_17402,N_8375,N_10388);
and U17403 (N_17403,N_11785,N_9326);
xor U17404 (N_17404,N_6831,N_10118);
and U17405 (N_17405,N_11213,N_10556);
or U17406 (N_17406,N_6586,N_11218);
and U17407 (N_17407,N_11325,N_10812);
and U17408 (N_17408,N_12353,N_8582);
xnor U17409 (N_17409,N_11480,N_7681);
or U17410 (N_17410,N_11874,N_10767);
and U17411 (N_17411,N_7789,N_10201);
nor U17412 (N_17412,N_6808,N_10356);
or U17413 (N_17413,N_8938,N_7783);
and U17414 (N_17414,N_7257,N_9212);
nand U17415 (N_17415,N_8576,N_10663);
nand U17416 (N_17416,N_9132,N_9428);
nand U17417 (N_17417,N_6678,N_6646);
and U17418 (N_17418,N_9972,N_7896);
nor U17419 (N_17419,N_10381,N_7521);
nand U17420 (N_17420,N_10748,N_8172);
nand U17421 (N_17421,N_12362,N_9416);
nand U17422 (N_17422,N_7103,N_10662);
and U17423 (N_17423,N_8406,N_8687);
nand U17424 (N_17424,N_11073,N_8143);
and U17425 (N_17425,N_6962,N_10047);
xor U17426 (N_17426,N_11338,N_7466);
or U17427 (N_17427,N_7003,N_6492);
nand U17428 (N_17428,N_8706,N_9312);
nor U17429 (N_17429,N_7513,N_9938);
nand U17430 (N_17430,N_8174,N_8553);
or U17431 (N_17431,N_9894,N_8623);
or U17432 (N_17432,N_8121,N_8223);
and U17433 (N_17433,N_12322,N_7509);
nand U17434 (N_17434,N_11362,N_8062);
and U17435 (N_17435,N_6753,N_8985);
and U17436 (N_17436,N_12461,N_11767);
nand U17437 (N_17437,N_10829,N_7441);
nor U17438 (N_17438,N_6608,N_9265);
nor U17439 (N_17439,N_10560,N_9452);
xor U17440 (N_17440,N_8909,N_6480);
nand U17441 (N_17441,N_11296,N_8168);
and U17442 (N_17442,N_11571,N_11429);
xnor U17443 (N_17443,N_9060,N_10949);
or U17444 (N_17444,N_7190,N_11383);
nand U17445 (N_17445,N_9725,N_6303);
and U17446 (N_17446,N_12329,N_8937);
or U17447 (N_17447,N_6552,N_6446);
xnor U17448 (N_17448,N_11802,N_9140);
nand U17449 (N_17449,N_10934,N_12265);
nor U17450 (N_17450,N_6394,N_6293);
or U17451 (N_17451,N_11588,N_11993);
nor U17452 (N_17452,N_7741,N_10787);
nand U17453 (N_17453,N_8149,N_7577);
xor U17454 (N_17454,N_11577,N_9763);
nand U17455 (N_17455,N_9048,N_11490);
xor U17456 (N_17456,N_10848,N_8920);
nand U17457 (N_17457,N_12471,N_12414);
or U17458 (N_17458,N_11997,N_11183);
or U17459 (N_17459,N_7129,N_11213);
xnor U17460 (N_17460,N_12120,N_12059);
and U17461 (N_17461,N_12049,N_11632);
and U17462 (N_17462,N_11225,N_8573);
xnor U17463 (N_17463,N_9408,N_9452);
nand U17464 (N_17464,N_11199,N_11581);
or U17465 (N_17465,N_9112,N_8291);
nand U17466 (N_17466,N_8766,N_9463);
nor U17467 (N_17467,N_8930,N_8256);
or U17468 (N_17468,N_12342,N_12154);
or U17469 (N_17469,N_8446,N_10581);
nand U17470 (N_17470,N_7592,N_9735);
and U17471 (N_17471,N_6926,N_7605);
or U17472 (N_17472,N_8551,N_8054);
xor U17473 (N_17473,N_10769,N_9723);
nor U17474 (N_17474,N_9566,N_10096);
and U17475 (N_17475,N_10747,N_8781);
nand U17476 (N_17476,N_10147,N_8888);
or U17477 (N_17477,N_12319,N_7173);
nor U17478 (N_17478,N_6577,N_8538);
xnor U17479 (N_17479,N_6695,N_7086);
nor U17480 (N_17480,N_6326,N_7932);
xor U17481 (N_17481,N_8878,N_9246);
nor U17482 (N_17482,N_11547,N_8248);
and U17483 (N_17483,N_12322,N_10642);
or U17484 (N_17484,N_7649,N_8463);
nor U17485 (N_17485,N_8206,N_10703);
xor U17486 (N_17486,N_11060,N_6608);
and U17487 (N_17487,N_9522,N_12256);
or U17488 (N_17488,N_10493,N_11114);
nand U17489 (N_17489,N_10702,N_11299);
nor U17490 (N_17490,N_9934,N_12243);
nand U17491 (N_17491,N_6911,N_12005);
nor U17492 (N_17492,N_11327,N_10794);
nor U17493 (N_17493,N_9032,N_11699);
nor U17494 (N_17494,N_8928,N_7946);
or U17495 (N_17495,N_7763,N_7245);
nor U17496 (N_17496,N_7067,N_8268);
nor U17497 (N_17497,N_11704,N_11553);
or U17498 (N_17498,N_10708,N_7054);
or U17499 (N_17499,N_11844,N_12217);
xnor U17500 (N_17500,N_10332,N_10259);
and U17501 (N_17501,N_10397,N_9451);
and U17502 (N_17502,N_10987,N_9563);
nor U17503 (N_17503,N_10390,N_9914);
xor U17504 (N_17504,N_6610,N_8147);
or U17505 (N_17505,N_10196,N_9395);
or U17506 (N_17506,N_6333,N_10068);
xnor U17507 (N_17507,N_11115,N_9707);
or U17508 (N_17508,N_9144,N_11100);
nand U17509 (N_17509,N_7743,N_7548);
nand U17510 (N_17510,N_11056,N_12029);
or U17511 (N_17511,N_9678,N_11643);
nand U17512 (N_17512,N_7912,N_9485);
nor U17513 (N_17513,N_6791,N_7962);
nor U17514 (N_17514,N_11373,N_7465);
or U17515 (N_17515,N_8441,N_11366);
and U17516 (N_17516,N_6691,N_9701);
and U17517 (N_17517,N_6914,N_9503);
or U17518 (N_17518,N_10870,N_11057);
xor U17519 (N_17519,N_12366,N_8404);
nand U17520 (N_17520,N_9225,N_7885);
nor U17521 (N_17521,N_12093,N_12279);
or U17522 (N_17522,N_10525,N_9646);
and U17523 (N_17523,N_9248,N_11906);
nand U17524 (N_17524,N_8364,N_9642);
xor U17525 (N_17525,N_10863,N_9118);
and U17526 (N_17526,N_8140,N_10584);
nor U17527 (N_17527,N_11444,N_11462);
xnor U17528 (N_17528,N_6961,N_11487);
nand U17529 (N_17529,N_10540,N_7772);
nor U17530 (N_17530,N_10886,N_10955);
nand U17531 (N_17531,N_6905,N_10048);
and U17532 (N_17532,N_10139,N_10878);
nor U17533 (N_17533,N_9621,N_10079);
nor U17534 (N_17534,N_10575,N_7969);
and U17535 (N_17535,N_11315,N_9252);
or U17536 (N_17536,N_6456,N_10612);
xor U17537 (N_17537,N_10026,N_11373);
xnor U17538 (N_17538,N_7094,N_11278);
or U17539 (N_17539,N_10090,N_8805);
nor U17540 (N_17540,N_11589,N_10557);
nor U17541 (N_17541,N_6935,N_12165);
and U17542 (N_17542,N_6376,N_9105);
nand U17543 (N_17543,N_6530,N_10972);
and U17544 (N_17544,N_9340,N_9497);
xor U17545 (N_17545,N_7264,N_7262);
xor U17546 (N_17546,N_6489,N_12416);
xnor U17547 (N_17547,N_6450,N_9449);
xnor U17548 (N_17548,N_7535,N_8835);
xnor U17549 (N_17549,N_10304,N_7308);
nor U17550 (N_17550,N_10270,N_8001);
and U17551 (N_17551,N_7410,N_6673);
nor U17552 (N_17552,N_10029,N_7913);
and U17553 (N_17553,N_12025,N_10610);
and U17554 (N_17554,N_7814,N_7647);
and U17555 (N_17555,N_9837,N_9078);
and U17556 (N_17556,N_10673,N_11291);
and U17557 (N_17557,N_9800,N_9667);
nor U17558 (N_17558,N_6474,N_6371);
and U17559 (N_17559,N_7420,N_9864);
or U17560 (N_17560,N_8149,N_9987);
or U17561 (N_17561,N_8712,N_11990);
nor U17562 (N_17562,N_10719,N_7925);
nand U17563 (N_17563,N_7755,N_6423);
and U17564 (N_17564,N_9156,N_8617);
nor U17565 (N_17565,N_9348,N_6437);
nand U17566 (N_17566,N_10289,N_10255);
and U17567 (N_17567,N_8476,N_8019);
nor U17568 (N_17568,N_6894,N_6873);
nor U17569 (N_17569,N_8806,N_9851);
xnor U17570 (N_17570,N_11113,N_7962);
xor U17571 (N_17571,N_11881,N_8983);
or U17572 (N_17572,N_11832,N_7715);
nor U17573 (N_17573,N_8229,N_7986);
nand U17574 (N_17574,N_10189,N_7263);
or U17575 (N_17575,N_10277,N_9285);
xor U17576 (N_17576,N_11268,N_7415);
nand U17577 (N_17577,N_11371,N_12340);
or U17578 (N_17578,N_10925,N_12020);
nor U17579 (N_17579,N_12001,N_6607);
nand U17580 (N_17580,N_11965,N_12086);
xnor U17581 (N_17581,N_10841,N_12432);
nand U17582 (N_17582,N_12030,N_11080);
or U17583 (N_17583,N_10051,N_11128);
nand U17584 (N_17584,N_10313,N_7235);
nor U17585 (N_17585,N_6417,N_11672);
nor U17586 (N_17586,N_9754,N_11772);
nand U17587 (N_17587,N_8562,N_8542);
xnor U17588 (N_17588,N_7976,N_10526);
nor U17589 (N_17589,N_8909,N_11143);
nor U17590 (N_17590,N_10254,N_7883);
nor U17591 (N_17591,N_6976,N_11671);
or U17592 (N_17592,N_6535,N_9365);
nand U17593 (N_17593,N_9479,N_9993);
nor U17594 (N_17594,N_8369,N_6387);
nor U17595 (N_17595,N_6793,N_6920);
or U17596 (N_17596,N_11658,N_9415);
nor U17597 (N_17597,N_7252,N_7622);
nand U17598 (N_17598,N_11831,N_10157);
nor U17599 (N_17599,N_9376,N_7219);
or U17600 (N_17600,N_8786,N_9767);
nand U17601 (N_17601,N_7134,N_9334);
or U17602 (N_17602,N_8052,N_11776);
or U17603 (N_17603,N_10558,N_10673);
xor U17604 (N_17604,N_8029,N_9828);
nor U17605 (N_17605,N_7560,N_7055);
nor U17606 (N_17606,N_7264,N_7156);
xor U17607 (N_17607,N_9172,N_8843);
xnor U17608 (N_17608,N_11210,N_7631);
nor U17609 (N_17609,N_11616,N_12131);
xor U17610 (N_17610,N_8505,N_7450);
and U17611 (N_17611,N_9586,N_8178);
nand U17612 (N_17612,N_9078,N_6295);
xnor U17613 (N_17613,N_11467,N_12098);
and U17614 (N_17614,N_12285,N_11863);
nand U17615 (N_17615,N_8178,N_12486);
and U17616 (N_17616,N_10843,N_6726);
nor U17617 (N_17617,N_6383,N_12138);
nand U17618 (N_17618,N_10484,N_7611);
xor U17619 (N_17619,N_11608,N_10742);
or U17620 (N_17620,N_6960,N_9945);
xor U17621 (N_17621,N_11097,N_8865);
nand U17622 (N_17622,N_11675,N_9267);
and U17623 (N_17623,N_9112,N_10972);
xor U17624 (N_17624,N_6974,N_10043);
nor U17625 (N_17625,N_8413,N_11445);
or U17626 (N_17626,N_10840,N_12333);
nor U17627 (N_17627,N_8494,N_8300);
xnor U17628 (N_17628,N_7219,N_8092);
or U17629 (N_17629,N_9404,N_7850);
xnor U17630 (N_17630,N_10329,N_11039);
nor U17631 (N_17631,N_9749,N_9127);
nor U17632 (N_17632,N_9784,N_7054);
nand U17633 (N_17633,N_8609,N_9890);
xnor U17634 (N_17634,N_10734,N_6563);
nand U17635 (N_17635,N_9736,N_7250);
xnor U17636 (N_17636,N_9582,N_9298);
nand U17637 (N_17637,N_7703,N_11378);
nor U17638 (N_17638,N_9955,N_9549);
xnor U17639 (N_17639,N_7254,N_7838);
xnor U17640 (N_17640,N_6252,N_10065);
nand U17641 (N_17641,N_6639,N_10700);
nor U17642 (N_17642,N_6766,N_11918);
nand U17643 (N_17643,N_6776,N_7175);
xor U17644 (N_17644,N_9811,N_10205);
nand U17645 (N_17645,N_12090,N_10300);
and U17646 (N_17646,N_8328,N_10723);
nor U17647 (N_17647,N_9927,N_8793);
and U17648 (N_17648,N_9238,N_8670);
nor U17649 (N_17649,N_6606,N_9800);
nor U17650 (N_17650,N_9681,N_6841);
and U17651 (N_17651,N_11323,N_7939);
and U17652 (N_17652,N_9845,N_7292);
xnor U17653 (N_17653,N_10958,N_8901);
xor U17654 (N_17654,N_11188,N_11491);
nand U17655 (N_17655,N_6405,N_9582);
or U17656 (N_17656,N_9083,N_8203);
and U17657 (N_17657,N_7727,N_10123);
nor U17658 (N_17658,N_7113,N_8001);
and U17659 (N_17659,N_12358,N_8172);
xnor U17660 (N_17660,N_8322,N_6756);
xor U17661 (N_17661,N_10509,N_9805);
or U17662 (N_17662,N_11944,N_7189);
xor U17663 (N_17663,N_7133,N_9632);
and U17664 (N_17664,N_12331,N_12316);
nand U17665 (N_17665,N_10595,N_6968);
xor U17666 (N_17666,N_10509,N_6845);
nor U17667 (N_17667,N_8833,N_6748);
nor U17668 (N_17668,N_8769,N_11787);
and U17669 (N_17669,N_7141,N_7465);
xor U17670 (N_17670,N_9548,N_6692);
nor U17671 (N_17671,N_8861,N_12456);
xor U17672 (N_17672,N_6474,N_9635);
nand U17673 (N_17673,N_8912,N_10697);
or U17674 (N_17674,N_8108,N_9526);
nand U17675 (N_17675,N_6784,N_8814);
and U17676 (N_17676,N_6501,N_12410);
or U17677 (N_17677,N_12402,N_11261);
or U17678 (N_17678,N_11772,N_9934);
nor U17679 (N_17679,N_11192,N_7637);
nor U17680 (N_17680,N_9709,N_7587);
and U17681 (N_17681,N_6629,N_11122);
or U17682 (N_17682,N_8305,N_8741);
xnor U17683 (N_17683,N_6381,N_11313);
or U17684 (N_17684,N_12165,N_12134);
and U17685 (N_17685,N_7352,N_8256);
xor U17686 (N_17686,N_10960,N_7444);
nand U17687 (N_17687,N_8008,N_10391);
xor U17688 (N_17688,N_9631,N_8253);
nor U17689 (N_17689,N_10418,N_9305);
xnor U17690 (N_17690,N_9108,N_11190);
nand U17691 (N_17691,N_8410,N_7454);
and U17692 (N_17692,N_9355,N_8526);
nor U17693 (N_17693,N_9392,N_9185);
xor U17694 (N_17694,N_7784,N_6485);
xnor U17695 (N_17695,N_11137,N_7150);
or U17696 (N_17696,N_10186,N_12350);
xnor U17697 (N_17697,N_9636,N_11197);
nor U17698 (N_17698,N_9884,N_8864);
and U17699 (N_17699,N_10281,N_6431);
and U17700 (N_17700,N_10843,N_11380);
or U17701 (N_17701,N_11448,N_8082);
or U17702 (N_17702,N_10208,N_6361);
or U17703 (N_17703,N_9972,N_9897);
nand U17704 (N_17704,N_6272,N_11018);
or U17705 (N_17705,N_6879,N_8031);
nand U17706 (N_17706,N_6693,N_11325);
or U17707 (N_17707,N_9354,N_6401);
and U17708 (N_17708,N_11702,N_12298);
and U17709 (N_17709,N_10092,N_10209);
and U17710 (N_17710,N_8857,N_11507);
nand U17711 (N_17711,N_11218,N_8826);
or U17712 (N_17712,N_11294,N_11817);
nor U17713 (N_17713,N_12376,N_9615);
nand U17714 (N_17714,N_12048,N_8597);
xor U17715 (N_17715,N_8517,N_10457);
nor U17716 (N_17716,N_9392,N_7192);
xor U17717 (N_17717,N_12149,N_11035);
nand U17718 (N_17718,N_10843,N_6817);
xor U17719 (N_17719,N_11718,N_9230);
and U17720 (N_17720,N_12181,N_6283);
nand U17721 (N_17721,N_6737,N_9027);
and U17722 (N_17722,N_6553,N_10413);
nor U17723 (N_17723,N_8782,N_6912);
xnor U17724 (N_17724,N_9937,N_11268);
nor U17725 (N_17725,N_8372,N_9159);
nor U17726 (N_17726,N_8304,N_10701);
and U17727 (N_17727,N_8723,N_10172);
xor U17728 (N_17728,N_6568,N_7966);
and U17729 (N_17729,N_9439,N_8611);
and U17730 (N_17730,N_9986,N_10534);
and U17731 (N_17731,N_8413,N_8996);
or U17732 (N_17732,N_9867,N_11170);
and U17733 (N_17733,N_9108,N_7672);
or U17734 (N_17734,N_9820,N_10820);
xnor U17735 (N_17735,N_10356,N_11021);
and U17736 (N_17736,N_8870,N_11491);
xnor U17737 (N_17737,N_6416,N_7421);
nor U17738 (N_17738,N_7114,N_10915);
nand U17739 (N_17739,N_9758,N_7634);
and U17740 (N_17740,N_8409,N_8452);
nand U17741 (N_17741,N_6537,N_12043);
or U17742 (N_17742,N_7114,N_8389);
nand U17743 (N_17743,N_7442,N_7143);
and U17744 (N_17744,N_8121,N_6967);
nand U17745 (N_17745,N_6335,N_10104);
or U17746 (N_17746,N_10249,N_9724);
nor U17747 (N_17747,N_11995,N_12385);
and U17748 (N_17748,N_8224,N_9805);
and U17749 (N_17749,N_8101,N_8758);
or U17750 (N_17750,N_7297,N_8073);
or U17751 (N_17751,N_7363,N_8764);
nand U17752 (N_17752,N_6636,N_8784);
nand U17753 (N_17753,N_8394,N_8041);
and U17754 (N_17754,N_9460,N_6361);
xor U17755 (N_17755,N_12029,N_10595);
or U17756 (N_17756,N_9318,N_9750);
or U17757 (N_17757,N_8639,N_9999);
nor U17758 (N_17758,N_8911,N_9358);
and U17759 (N_17759,N_9224,N_10831);
xnor U17760 (N_17760,N_8879,N_11839);
nand U17761 (N_17761,N_11896,N_6651);
xor U17762 (N_17762,N_10131,N_9928);
nand U17763 (N_17763,N_9272,N_6358);
nor U17764 (N_17764,N_11412,N_12150);
nor U17765 (N_17765,N_10098,N_10693);
xor U17766 (N_17766,N_8108,N_7105);
xor U17767 (N_17767,N_8337,N_7421);
and U17768 (N_17768,N_6640,N_9064);
or U17769 (N_17769,N_8675,N_10326);
xnor U17770 (N_17770,N_8956,N_9295);
nor U17771 (N_17771,N_9586,N_9770);
or U17772 (N_17772,N_7904,N_11836);
xor U17773 (N_17773,N_7408,N_10630);
nand U17774 (N_17774,N_8831,N_8029);
xor U17775 (N_17775,N_6901,N_11142);
xor U17776 (N_17776,N_9087,N_7003);
nor U17777 (N_17777,N_6858,N_11286);
nand U17778 (N_17778,N_12091,N_6529);
nor U17779 (N_17779,N_11383,N_8848);
and U17780 (N_17780,N_10897,N_11937);
xnor U17781 (N_17781,N_9823,N_8347);
nor U17782 (N_17782,N_6771,N_11574);
nor U17783 (N_17783,N_11279,N_6689);
nor U17784 (N_17784,N_7465,N_6607);
xor U17785 (N_17785,N_8207,N_9783);
and U17786 (N_17786,N_10432,N_7241);
nand U17787 (N_17787,N_10271,N_9349);
nor U17788 (N_17788,N_8396,N_12074);
and U17789 (N_17789,N_10443,N_10757);
xor U17790 (N_17790,N_11150,N_7601);
xnor U17791 (N_17791,N_8985,N_7848);
xnor U17792 (N_17792,N_6621,N_7732);
nor U17793 (N_17793,N_8799,N_9784);
nor U17794 (N_17794,N_10048,N_11254);
or U17795 (N_17795,N_12213,N_11849);
nor U17796 (N_17796,N_11254,N_9734);
xnor U17797 (N_17797,N_11699,N_10590);
nand U17798 (N_17798,N_12490,N_11206);
and U17799 (N_17799,N_9908,N_11121);
nor U17800 (N_17800,N_8021,N_10166);
xor U17801 (N_17801,N_8887,N_7691);
and U17802 (N_17802,N_7140,N_10560);
nor U17803 (N_17803,N_8874,N_11172);
and U17804 (N_17804,N_7079,N_9856);
nand U17805 (N_17805,N_9290,N_11478);
xnor U17806 (N_17806,N_11703,N_8055);
and U17807 (N_17807,N_7523,N_7982);
or U17808 (N_17808,N_11648,N_6691);
and U17809 (N_17809,N_10610,N_11241);
nand U17810 (N_17810,N_11108,N_8503);
or U17811 (N_17811,N_6376,N_9846);
nor U17812 (N_17812,N_11591,N_10703);
or U17813 (N_17813,N_10618,N_6610);
and U17814 (N_17814,N_7687,N_8975);
and U17815 (N_17815,N_8912,N_10575);
nor U17816 (N_17816,N_8290,N_10935);
nor U17817 (N_17817,N_9990,N_8068);
or U17818 (N_17818,N_9495,N_6454);
nor U17819 (N_17819,N_9058,N_9096);
nand U17820 (N_17820,N_7940,N_10748);
and U17821 (N_17821,N_8225,N_11010);
nor U17822 (N_17822,N_10211,N_7766);
nand U17823 (N_17823,N_12241,N_9743);
nor U17824 (N_17824,N_8672,N_8053);
nor U17825 (N_17825,N_11452,N_9181);
xor U17826 (N_17826,N_10319,N_6956);
xnor U17827 (N_17827,N_6439,N_6386);
nand U17828 (N_17828,N_10530,N_11185);
xnor U17829 (N_17829,N_8695,N_7486);
nand U17830 (N_17830,N_9241,N_6940);
nor U17831 (N_17831,N_11114,N_11111);
nand U17832 (N_17832,N_9295,N_11373);
nor U17833 (N_17833,N_11597,N_6520);
or U17834 (N_17834,N_11449,N_10454);
and U17835 (N_17835,N_9247,N_10525);
and U17836 (N_17836,N_10855,N_8401);
or U17837 (N_17837,N_11719,N_10490);
nand U17838 (N_17838,N_10028,N_12126);
nand U17839 (N_17839,N_11099,N_6486);
or U17840 (N_17840,N_7679,N_8496);
nand U17841 (N_17841,N_8453,N_10518);
and U17842 (N_17842,N_8614,N_11935);
nor U17843 (N_17843,N_6706,N_10897);
xor U17844 (N_17844,N_11410,N_7998);
nor U17845 (N_17845,N_6996,N_8540);
nand U17846 (N_17846,N_9859,N_9785);
xor U17847 (N_17847,N_6653,N_10367);
nor U17848 (N_17848,N_11421,N_11371);
and U17849 (N_17849,N_7569,N_7536);
nand U17850 (N_17850,N_7286,N_9872);
nand U17851 (N_17851,N_7144,N_10884);
nor U17852 (N_17852,N_9290,N_8156);
xnor U17853 (N_17853,N_6645,N_11481);
nand U17854 (N_17854,N_8109,N_6592);
nor U17855 (N_17855,N_9120,N_10637);
and U17856 (N_17856,N_11355,N_7384);
nand U17857 (N_17857,N_9519,N_11080);
or U17858 (N_17858,N_8383,N_6339);
xor U17859 (N_17859,N_6437,N_12096);
and U17860 (N_17860,N_8003,N_6783);
and U17861 (N_17861,N_7279,N_11321);
xor U17862 (N_17862,N_11586,N_11566);
and U17863 (N_17863,N_8344,N_8236);
nand U17864 (N_17864,N_9896,N_8496);
xor U17865 (N_17865,N_9697,N_8110);
nand U17866 (N_17866,N_9988,N_10004);
or U17867 (N_17867,N_8940,N_10378);
nor U17868 (N_17868,N_6651,N_7071);
xor U17869 (N_17869,N_7722,N_8984);
or U17870 (N_17870,N_10576,N_8675);
or U17871 (N_17871,N_8753,N_11732);
xnor U17872 (N_17872,N_7420,N_8421);
xnor U17873 (N_17873,N_11051,N_11088);
and U17874 (N_17874,N_6554,N_11264);
and U17875 (N_17875,N_6595,N_7460);
or U17876 (N_17876,N_9431,N_11380);
and U17877 (N_17877,N_6822,N_6753);
and U17878 (N_17878,N_9901,N_8818);
and U17879 (N_17879,N_10896,N_6627);
xnor U17880 (N_17880,N_10838,N_11043);
or U17881 (N_17881,N_9058,N_6260);
nor U17882 (N_17882,N_6912,N_6315);
and U17883 (N_17883,N_8647,N_12311);
nand U17884 (N_17884,N_6614,N_8524);
and U17885 (N_17885,N_7087,N_9865);
or U17886 (N_17886,N_11310,N_10216);
or U17887 (N_17887,N_8380,N_10091);
or U17888 (N_17888,N_10352,N_7736);
xnor U17889 (N_17889,N_9270,N_8655);
nand U17890 (N_17890,N_9120,N_9134);
nand U17891 (N_17891,N_9057,N_9294);
nor U17892 (N_17892,N_8116,N_8982);
xor U17893 (N_17893,N_12038,N_6586);
and U17894 (N_17894,N_12158,N_6387);
and U17895 (N_17895,N_7971,N_8014);
nand U17896 (N_17896,N_9114,N_11900);
or U17897 (N_17897,N_9644,N_9110);
xnor U17898 (N_17898,N_11544,N_10282);
or U17899 (N_17899,N_8611,N_11467);
and U17900 (N_17900,N_6510,N_11813);
nand U17901 (N_17901,N_8319,N_11985);
nor U17902 (N_17902,N_7949,N_8116);
and U17903 (N_17903,N_7610,N_7676);
nand U17904 (N_17904,N_8365,N_10051);
or U17905 (N_17905,N_7182,N_6478);
nand U17906 (N_17906,N_6844,N_9756);
xnor U17907 (N_17907,N_11294,N_10866);
nor U17908 (N_17908,N_10248,N_11670);
xor U17909 (N_17909,N_12211,N_11800);
nor U17910 (N_17910,N_11170,N_11450);
or U17911 (N_17911,N_10765,N_8866);
nor U17912 (N_17912,N_9050,N_6944);
and U17913 (N_17913,N_11195,N_6517);
nand U17914 (N_17914,N_11462,N_9430);
xor U17915 (N_17915,N_8341,N_6915);
and U17916 (N_17916,N_7806,N_6568);
nand U17917 (N_17917,N_10575,N_8314);
nand U17918 (N_17918,N_11980,N_12274);
nand U17919 (N_17919,N_6777,N_6943);
nand U17920 (N_17920,N_6807,N_6588);
nor U17921 (N_17921,N_9968,N_11598);
nor U17922 (N_17922,N_11759,N_12293);
and U17923 (N_17923,N_10833,N_8951);
xor U17924 (N_17924,N_12082,N_9953);
and U17925 (N_17925,N_8980,N_6865);
or U17926 (N_17926,N_12300,N_11295);
xnor U17927 (N_17927,N_11825,N_8605);
xor U17928 (N_17928,N_12283,N_9731);
xor U17929 (N_17929,N_11310,N_11883);
and U17930 (N_17930,N_8483,N_9716);
xor U17931 (N_17931,N_8964,N_9794);
nand U17932 (N_17932,N_6273,N_6905);
nand U17933 (N_17933,N_6636,N_9154);
xnor U17934 (N_17934,N_6522,N_12136);
or U17935 (N_17935,N_12328,N_7066);
nor U17936 (N_17936,N_7221,N_6315);
nand U17937 (N_17937,N_10821,N_11163);
or U17938 (N_17938,N_12102,N_10244);
nor U17939 (N_17939,N_7320,N_10530);
and U17940 (N_17940,N_8345,N_9058);
xnor U17941 (N_17941,N_8536,N_8426);
nand U17942 (N_17942,N_9468,N_7965);
and U17943 (N_17943,N_10298,N_7373);
nor U17944 (N_17944,N_12453,N_8565);
xor U17945 (N_17945,N_10125,N_6325);
nor U17946 (N_17946,N_11110,N_10766);
and U17947 (N_17947,N_9228,N_10732);
xor U17948 (N_17948,N_11167,N_10639);
and U17949 (N_17949,N_7700,N_10041);
and U17950 (N_17950,N_9385,N_6451);
and U17951 (N_17951,N_7444,N_8595);
xor U17952 (N_17952,N_9442,N_8350);
nand U17953 (N_17953,N_12400,N_11930);
and U17954 (N_17954,N_11577,N_8614);
or U17955 (N_17955,N_9708,N_6628);
or U17956 (N_17956,N_10541,N_8227);
nor U17957 (N_17957,N_12344,N_10095);
nand U17958 (N_17958,N_12011,N_6742);
nand U17959 (N_17959,N_12099,N_6471);
xor U17960 (N_17960,N_8004,N_9630);
and U17961 (N_17961,N_10970,N_11504);
or U17962 (N_17962,N_10733,N_9734);
xor U17963 (N_17963,N_9724,N_11215);
nand U17964 (N_17964,N_6587,N_7167);
xor U17965 (N_17965,N_8244,N_10604);
or U17966 (N_17966,N_11208,N_7518);
xnor U17967 (N_17967,N_11589,N_12032);
or U17968 (N_17968,N_8088,N_11893);
nand U17969 (N_17969,N_9157,N_8937);
xor U17970 (N_17970,N_6981,N_10819);
nor U17971 (N_17971,N_8869,N_9445);
nand U17972 (N_17972,N_11451,N_12233);
and U17973 (N_17973,N_10753,N_9261);
nor U17974 (N_17974,N_9878,N_6526);
nand U17975 (N_17975,N_8186,N_7579);
or U17976 (N_17976,N_7867,N_11346);
or U17977 (N_17977,N_8796,N_8534);
and U17978 (N_17978,N_8620,N_10237);
or U17979 (N_17979,N_9399,N_9434);
nor U17980 (N_17980,N_6977,N_11898);
and U17981 (N_17981,N_12151,N_9081);
or U17982 (N_17982,N_11820,N_7174);
xor U17983 (N_17983,N_7205,N_6780);
and U17984 (N_17984,N_6264,N_10368);
or U17985 (N_17985,N_9495,N_12235);
and U17986 (N_17986,N_9385,N_11315);
and U17987 (N_17987,N_6536,N_6922);
or U17988 (N_17988,N_7086,N_11877);
nor U17989 (N_17989,N_11724,N_12295);
nor U17990 (N_17990,N_11122,N_9687);
xnor U17991 (N_17991,N_7318,N_12435);
nor U17992 (N_17992,N_9520,N_10554);
xor U17993 (N_17993,N_10794,N_11604);
and U17994 (N_17994,N_11036,N_11916);
and U17995 (N_17995,N_11599,N_10929);
nor U17996 (N_17996,N_6277,N_11495);
nand U17997 (N_17997,N_6904,N_6698);
nand U17998 (N_17998,N_12289,N_9902);
nand U17999 (N_17999,N_8695,N_6860);
and U18000 (N_18000,N_7839,N_8729);
or U18001 (N_18001,N_10957,N_10260);
nand U18002 (N_18002,N_7005,N_10178);
nand U18003 (N_18003,N_6728,N_12429);
or U18004 (N_18004,N_6436,N_11533);
and U18005 (N_18005,N_8576,N_11478);
nand U18006 (N_18006,N_10609,N_8231);
nand U18007 (N_18007,N_10869,N_8614);
and U18008 (N_18008,N_9773,N_10454);
nor U18009 (N_18009,N_6325,N_8875);
or U18010 (N_18010,N_11106,N_9182);
or U18011 (N_18011,N_9191,N_8160);
or U18012 (N_18012,N_9694,N_6295);
or U18013 (N_18013,N_7936,N_11090);
and U18014 (N_18014,N_9375,N_7538);
xor U18015 (N_18015,N_11742,N_12079);
xor U18016 (N_18016,N_7502,N_8054);
nand U18017 (N_18017,N_12318,N_11654);
nand U18018 (N_18018,N_8861,N_8577);
nand U18019 (N_18019,N_6641,N_12255);
or U18020 (N_18020,N_9759,N_7286);
or U18021 (N_18021,N_9671,N_7994);
or U18022 (N_18022,N_7528,N_7384);
or U18023 (N_18023,N_10860,N_12191);
or U18024 (N_18024,N_11140,N_12379);
or U18025 (N_18025,N_6879,N_7662);
nor U18026 (N_18026,N_7195,N_10674);
nand U18027 (N_18027,N_7450,N_7773);
or U18028 (N_18028,N_7788,N_10276);
and U18029 (N_18029,N_11388,N_9474);
nor U18030 (N_18030,N_6491,N_8129);
nor U18031 (N_18031,N_6764,N_8773);
xor U18032 (N_18032,N_9872,N_8275);
nand U18033 (N_18033,N_8793,N_10201);
nand U18034 (N_18034,N_11485,N_11231);
and U18035 (N_18035,N_11781,N_10693);
and U18036 (N_18036,N_9153,N_10055);
or U18037 (N_18037,N_7369,N_10468);
or U18038 (N_18038,N_6482,N_7233);
nand U18039 (N_18039,N_8297,N_8200);
xnor U18040 (N_18040,N_9589,N_7812);
nor U18041 (N_18041,N_12229,N_7891);
and U18042 (N_18042,N_11019,N_10264);
or U18043 (N_18043,N_7442,N_8734);
nand U18044 (N_18044,N_7022,N_7532);
xor U18045 (N_18045,N_7715,N_6845);
nand U18046 (N_18046,N_7955,N_8833);
nor U18047 (N_18047,N_7997,N_9165);
and U18048 (N_18048,N_10470,N_8980);
nor U18049 (N_18049,N_8986,N_6478);
nor U18050 (N_18050,N_8463,N_11759);
and U18051 (N_18051,N_11332,N_11986);
xnor U18052 (N_18052,N_11953,N_8557);
and U18053 (N_18053,N_10504,N_6636);
nor U18054 (N_18054,N_8092,N_7228);
xor U18055 (N_18055,N_7035,N_10867);
nand U18056 (N_18056,N_10664,N_6798);
or U18057 (N_18057,N_9014,N_7225);
nand U18058 (N_18058,N_8089,N_8732);
nand U18059 (N_18059,N_12343,N_10698);
and U18060 (N_18060,N_10157,N_8137);
nor U18061 (N_18061,N_12084,N_8920);
xnor U18062 (N_18062,N_11395,N_9387);
nand U18063 (N_18063,N_6593,N_7394);
nand U18064 (N_18064,N_7169,N_6715);
nor U18065 (N_18065,N_10685,N_6412);
xor U18066 (N_18066,N_11024,N_8206);
and U18067 (N_18067,N_10673,N_6431);
nand U18068 (N_18068,N_7586,N_9203);
xor U18069 (N_18069,N_8439,N_10974);
xnor U18070 (N_18070,N_12172,N_9531);
or U18071 (N_18071,N_8332,N_8487);
xnor U18072 (N_18072,N_7903,N_8412);
xor U18073 (N_18073,N_12041,N_11589);
or U18074 (N_18074,N_7631,N_11902);
nor U18075 (N_18075,N_6921,N_7265);
or U18076 (N_18076,N_8760,N_9777);
or U18077 (N_18077,N_6565,N_6838);
or U18078 (N_18078,N_8261,N_7463);
xor U18079 (N_18079,N_6628,N_10143);
nand U18080 (N_18080,N_6695,N_12221);
and U18081 (N_18081,N_10738,N_11777);
xnor U18082 (N_18082,N_6651,N_7376);
nand U18083 (N_18083,N_6299,N_10444);
or U18084 (N_18084,N_7021,N_10254);
nor U18085 (N_18085,N_11258,N_11194);
and U18086 (N_18086,N_6277,N_7693);
nor U18087 (N_18087,N_9328,N_9968);
xor U18088 (N_18088,N_10188,N_9904);
nand U18089 (N_18089,N_10966,N_6907);
xor U18090 (N_18090,N_10683,N_7906);
or U18091 (N_18091,N_8055,N_8625);
or U18092 (N_18092,N_10824,N_10042);
nand U18093 (N_18093,N_11164,N_10875);
xnor U18094 (N_18094,N_12227,N_7352);
and U18095 (N_18095,N_10194,N_7660);
nor U18096 (N_18096,N_10497,N_12473);
nor U18097 (N_18097,N_8610,N_6957);
xor U18098 (N_18098,N_11343,N_7001);
nor U18099 (N_18099,N_11594,N_10837);
nand U18100 (N_18100,N_10579,N_7894);
or U18101 (N_18101,N_11474,N_9867);
or U18102 (N_18102,N_9468,N_6859);
and U18103 (N_18103,N_7035,N_7523);
nor U18104 (N_18104,N_7960,N_7822);
nor U18105 (N_18105,N_10681,N_7025);
and U18106 (N_18106,N_11214,N_9019);
nor U18107 (N_18107,N_8453,N_10666);
nand U18108 (N_18108,N_6324,N_10642);
and U18109 (N_18109,N_11075,N_7547);
or U18110 (N_18110,N_7424,N_7091);
and U18111 (N_18111,N_11045,N_8316);
nor U18112 (N_18112,N_9558,N_12457);
or U18113 (N_18113,N_7096,N_7763);
xor U18114 (N_18114,N_8008,N_9688);
nand U18115 (N_18115,N_12499,N_11573);
or U18116 (N_18116,N_11796,N_9034);
nor U18117 (N_18117,N_7374,N_11814);
nor U18118 (N_18118,N_10098,N_9597);
and U18119 (N_18119,N_8661,N_6657);
xnor U18120 (N_18120,N_12428,N_11646);
nand U18121 (N_18121,N_9121,N_6689);
or U18122 (N_18122,N_7128,N_6996);
and U18123 (N_18123,N_11933,N_7784);
nor U18124 (N_18124,N_11437,N_9693);
nand U18125 (N_18125,N_12115,N_10007);
or U18126 (N_18126,N_7209,N_9791);
nor U18127 (N_18127,N_9739,N_12118);
and U18128 (N_18128,N_11554,N_9486);
or U18129 (N_18129,N_8802,N_8440);
or U18130 (N_18130,N_12079,N_10886);
or U18131 (N_18131,N_9717,N_6627);
and U18132 (N_18132,N_9560,N_11174);
or U18133 (N_18133,N_11367,N_6885);
and U18134 (N_18134,N_10889,N_6260);
nor U18135 (N_18135,N_6295,N_11314);
xnor U18136 (N_18136,N_10893,N_8879);
nor U18137 (N_18137,N_9190,N_11666);
nand U18138 (N_18138,N_6993,N_8615);
nand U18139 (N_18139,N_12402,N_9909);
and U18140 (N_18140,N_11645,N_6484);
nand U18141 (N_18141,N_7446,N_11802);
and U18142 (N_18142,N_8651,N_8056);
xnor U18143 (N_18143,N_8447,N_7692);
and U18144 (N_18144,N_9310,N_12127);
or U18145 (N_18145,N_9393,N_9771);
and U18146 (N_18146,N_7744,N_6998);
and U18147 (N_18147,N_10315,N_9007);
nand U18148 (N_18148,N_10726,N_8968);
and U18149 (N_18149,N_8226,N_10291);
nand U18150 (N_18150,N_8343,N_9585);
xor U18151 (N_18151,N_9416,N_7471);
nor U18152 (N_18152,N_9556,N_11416);
or U18153 (N_18153,N_8756,N_7544);
xor U18154 (N_18154,N_10104,N_9239);
and U18155 (N_18155,N_7594,N_8328);
or U18156 (N_18156,N_11068,N_10314);
and U18157 (N_18157,N_6296,N_8919);
xnor U18158 (N_18158,N_7238,N_8512);
or U18159 (N_18159,N_8024,N_8936);
nand U18160 (N_18160,N_10598,N_7619);
or U18161 (N_18161,N_11354,N_10187);
nand U18162 (N_18162,N_7332,N_11565);
nor U18163 (N_18163,N_8409,N_12202);
and U18164 (N_18164,N_9414,N_11443);
and U18165 (N_18165,N_8698,N_9404);
and U18166 (N_18166,N_8694,N_11332);
xnor U18167 (N_18167,N_11176,N_7299);
and U18168 (N_18168,N_10828,N_6709);
nand U18169 (N_18169,N_10160,N_6456);
and U18170 (N_18170,N_10735,N_6755);
xnor U18171 (N_18171,N_9596,N_10759);
and U18172 (N_18172,N_7857,N_10040);
nor U18173 (N_18173,N_6386,N_10640);
xor U18174 (N_18174,N_6934,N_9912);
and U18175 (N_18175,N_10362,N_8723);
nor U18176 (N_18176,N_10236,N_10157);
nand U18177 (N_18177,N_7629,N_12480);
xnor U18178 (N_18178,N_10744,N_6587);
xnor U18179 (N_18179,N_7976,N_9197);
xnor U18180 (N_18180,N_8360,N_7198);
or U18181 (N_18181,N_10993,N_11512);
and U18182 (N_18182,N_9704,N_11233);
or U18183 (N_18183,N_11007,N_6869);
nor U18184 (N_18184,N_12386,N_8409);
xor U18185 (N_18185,N_7968,N_10404);
xor U18186 (N_18186,N_9586,N_11021);
xnor U18187 (N_18187,N_8502,N_6871);
or U18188 (N_18188,N_11426,N_8017);
xor U18189 (N_18189,N_9079,N_12112);
nand U18190 (N_18190,N_9599,N_7619);
nor U18191 (N_18191,N_9854,N_11113);
xnor U18192 (N_18192,N_8232,N_6955);
or U18193 (N_18193,N_10932,N_7747);
xor U18194 (N_18194,N_8727,N_9836);
xnor U18195 (N_18195,N_6598,N_11648);
nand U18196 (N_18196,N_9361,N_8811);
nor U18197 (N_18197,N_10011,N_7621);
nor U18198 (N_18198,N_12285,N_6701);
xnor U18199 (N_18199,N_12111,N_12131);
xnor U18200 (N_18200,N_11910,N_7088);
and U18201 (N_18201,N_8350,N_12124);
xor U18202 (N_18202,N_7970,N_9082);
nand U18203 (N_18203,N_6990,N_12454);
and U18204 (N_18204,N_12213,N_9921);
and U18205 (N_18205,N_7056,N_7660);
nor U18206 (N_18206,N_9664,N_11080);
xnor U18207 (N_18207,N_7732,N_10766);
xnor U18208 (N_18208,N_11341,N_7624);
xnor U18209 (N_18209,N_12016,N_7447);
or U18210 (N_18210,N_6850,N_10233);
or U18211 (N_18211,N_8403,N_6644);
nand U18212 (N_18212,N_10759,N_12263);
or U18213 (N_18213,N_9513,N_9634);
and U18214 (N_18214,N_7404,N_7919);
and U18215 (N_18215,N_10383,N_8866);
xnor U18216 (N_18216,N_6962,N_9127);
nor U18217 (N_18217,N_12235,N_11216);
and U18218 (N_18218,N_10708,N_11020);
xnor U18219 (N_18219,N_8243,N_10197);
xor U18220 (N_18220,N_10541,N_10445);
nor U18221 (N_18221,N_8212,N_9146);
or U18222 (N_18222,N_9060,N_7716);
or U18223 (N_18223,N_8137,N_10652);
xor U18224 (N_18224,N_9602,N_6864);
xor U18225 (N_18225,N_9245,N_8226);
nor U18226 (N_18226,N_8591,N_11451);
xnor U18227 (N_18227,N_10045,N_9649);
or U18228 (N_18228,N_8867,N_10969);
nand U18229 (N_18229,N_11988,N_7610);
xor U18230 (N_18230,N_11019,N_7188);
and U18231 (N_18231,N_8824,N_10655);
xor U18232 (N_18232,N_10143,N_8494);
xor U18233 (N_18233,N_12451,N_9090);
nand U18234 (N_18234,N_6548,N_6483);
nor U18235 (N_18235,N_12077,N_10752);
nor U18236 (N_18236,N_10656,N_11172);
nor U18237 (N_18237,N_7925,N_8295);
or U18238 (N_18238,N_9908,N_6381);
nand U18239 (N_18239,N_8068,N_10597);
xnor U18240 (N_18240,N_9446,N_12243);
and U18241 (N_18241,N_11425,N_11464);
xnor U18242 (N_18242,N_9750,N_11560);
nor U18243 (N_18243,N_6547,N_6715);
or U18244 (N_18244,N_8945,N_10738);
nand U18245 (N_18245,N_11927,N_7028);
nor U18246 (N_18246,N_6538,N_11043);
xor U18247 (N_18247,N_6742,N_10897);
and U18248 (N_18248,N_9937,N_7984);
or U18249 (N_18249,N_9515,N_7719);
and U18250 (N_18250,N_6949,N_8619);
nor U18251 (N_18251,N_6535,N_11135);
or U18252 (N_18252,N_11426,N_11616);
nand U18253 (N_18253,N_10667,N_8623);
or U18254 (N_18254,N_6268,N_9283);
nand U18255 (N_18255,N_11640,N_6706);
or U18256 (N_18256,N_7651,N_7891);
nor U18257 (N_18257,N_10978,N_8907);
xnor U18258 (N_18258,N_11084,N_8488);
or U18259 (N_18259,N_7192,N_9614);
nand U18260 (N_18260,N_7707,N_8948);
nand U18261 (N_18261,N_9301,N_7525);
xnor U18262 (N_18262,N_9384,N_11287);
nand U18263 (N_18263,N_7236,N_6255);
and U18264 (N_18264,N_9991,N_8713);
nor U18265 (N_18265,N_10125,N_7257);
and U18266 (N_18266,N_7705,N_7156);
or U18267 (N_18267,N_8940,N_12020);
nor U18268 (N_18268,N_12340,N_9749);
nand U18269 (N_18269,N_9126,N_9446);
nand U18270 (N_18270,N_11440,N_11483);
or U18271 (N_18271,N_8664,N_8128);
nor U18272 (N_18272,N_8772,N_7977);
or U18273 (N_18273,N_12212,N_6954);
xnor U18274 (N_18274,N_10936,N_10886);
nand U18275 (N_18275,N_9427,N_10075);
nor U18276 (N_18276,N_10517,N_9958);
nor U18277 (N_18277,N_7385,N_6941);
or U18278 (N_18278,N_9224,N_8910);
and U18279 (N_18279,N_8477,N_11690);
nand U18280 (N_18280,N_12353,N_9794);
nand U18281 (N_18281,N_6383,N_6998);
nand U18282 (N_18282,N_11154,N_7336);
nor U18283 (N_18283,N_12411,N_10888);
nor U18284 (N_18284,N_7066,N_8324);
nor U18285 (N_18285,N_8787,N_12049);
nand U18286 (N_18286,N_10841,N_9895);
nor U18287 (N_18287,N_6800,N_7539);
nor U18288 (N_18288,N_12302,N_10627);
xor U18289 (N_18289,N_7378,N_10314);
or U18290 (N_18290,N_8582,N_8143);
nand U18291 (N_18291,N_7874,N_6716);
xnor U18292 (N_18292,N_10250,N_9249);
nor U18293 (N_18293,N_9361,N_8997);
xor U18294 (N_18294,N_10033,N_8584);
xnor U18295 (N_18295,N_11543,N_7810);
nor U18296 (N_18296,N_11363,N_10467);
xnor U18297 (N_18297,N_11760,N_10432);
nand U18298 (N_18298,N_10221,N_9459);
and U18299 (N_18299,N_9048,N_7722);
and U18300 (N_18300,N_7985,N_6542);
or U18301 (N_18301,N_7007,N_9113);
xnor U18302 (N_18302,N_8294,N_11480);
xor U18303 (N_18303,N_8680,N_7443);
or U18304 (N_18304,N_11822,N_9086);
xor U18305 (N_18305,N_9580,N_6595);
or U18306 (N_18306,N_8461,N_9215);
nor U18307 (N_18307,N_12120,N_8930);
or U18308 (N_18308,N_9975,N_9695);
or U18309 (N_18309,N_6407,N_8743);
xor U18310 (N_18310,N_8705,N_10855);
or U18311 (N_18311,N_12437,N_11527);
nor U18312 (N_18312,N_11814,N_6534);
or U18313 (N_18313,N_9493,N_11119);
xor U18314 (N_18314,N_10500,N_10435);
or U18315 (N_18315,N_9842,N_10665);
nand U18316 (N_18316,N_11102,N_9996);
nor U18317 (N_18317,N_6655,N_7282);
or U18318 (N_18318,N_11972,N_11517);
nor U18319 (N_18319,N_8768,N_7954);
nor U18320 (N_18320,N_6963,N_10348);
or U18321 (N_18321,N_7555,N_8728);
or U18322 (N_18322,N_7034,N_11616);
nor U18323 (N_18323,N_8615,N_8264);
xnor U18324 (N_18324,N_8261,N_7381);
and U18325 (N_18325,N_6345,N_11601);
or U18326 (N_18326,N_11762,N_12022);
and U18327 (N_18327,N_12011,N_10924);
nor U18328 (N_18328,N_9534,N_8128);
nor U18329 (N_18329,N_9720,N_10569);
xor U18330 (N_18330,N_11616,N_7181);
and U18331 (N_18331,N_11471,N_8685);
xor U18332 (N_18332,N_11594,N_8387);
nand U18333 (N_18333,N_10976,N_8934);
nor U18334 (N_18334,N_8996,N_8264);
and U18335 (N_18335,N_11510,N_8562);
nand U18336 (N_18336,N_10709,N_6441);
or U18337 (N_18337,N_7893,N_12208);
or U18338 (N_18338,N_6557,N_9776);
or U18339 (N_18339,N_11387,N_6590);
nor U18340 (N_18340,N_11662,N_8550);
and U18341 (N_18341,N_10227,N_9358);
and U18342 (N_18342,N_8057,N_11913);
nand U18343 (N_18343,N_10288,N_6461);
nor U18344 (N_18344,N_9288,N_9354);
and U18345 (N_18345,N_9565,N_11546);
and U18346 (N_18346,N_11502,N_9181);
nand U18347 (N_18347,N_7802,N_6819);
xnor U18348 (N_18348,N_7246,N_6748);
or U18349 (N_18349,N_12493,N_9434);
nand U18350 (N_18350,N_8167,N_7831);
nor U18351 (N_18351,N_8622,N_8807);
nand U18352 (N_18352,N_8029,N_8142);
nor U18353 (N_18353,N_6495,N_6493);
nand U18354 (N_18354,N_7627,N_9503);
nor U18355 (N_18355,N_12474,N_8414);
or U18356 (N_18356,N_8518,N_12449);
nand U18357 (N_18357,N_10209,N_8672);
or U18358 (N_18358,N_6548,N_12258);
and U18359 (N_18359,N_8743,N_7932);
nand U18360 (N_18360,N_9206,N_10837);
nand U18361 (N_18361,N_9701,N_10061);
or U18362 (N_18362,N_6664,N_8344);
and U18363 (N_18363,N_9775,N_7637);
nor U18364 (N_18364,N_9926,N_12414);
xnor U18365 (N_18365,N_9814,N_7041);
xor U18366 (N_18366,N_9166,N_11803);
and U18367 (N_18367,N_7235,N_7066);
or U18368 (N_18368,N_9733,N_7846);
xnor U18369 (N_18369,N_9601,N_8075);
nor U18370 (N_18370,N_11574,N_7373);
or U18371 (N_18371,N_6534,N_8563);
and U18372 (N_18372,N_12155,N_7683);
and U18373 (N_18373,N_9862,N_11247);
and U18374 (N_18374,N_7878,N_10048);
and U18375 (N_18375,N_10697,N_11304);
xnor U18376 (N_18376,N_8098,N_10563);
nor U18377 (N_18377,N_11748,N_9603);
xor U18378 (N_18378,N_8889,N_9262);
nor U18379 (N_18379,N_12013,N_7039);
nor U18380 (N_18380,N_10389,N_6736);
or U18381 (N_18381,N_6415,N_7079);
nor U18382 (N_18382,N_9660,N_6651);
nand U18383 (N_18383,N_8969,N_8008);
or U18384 (N_18384,N_8859,N_10329);
nor U18385 (N_18385,N_8489,N_11645);
xnor U18386 (N_18386,N_9290,N_12356);
or U18387 (N_18387,N_8630,N_7749);
xnor U18388 (N_18388,N_8927,N_9934);
nand U18389 (N_18389,N_9384,N_9868);
nand U18390 (N_18390,N_6709,N_9973);
nor U18391 (N_18391,N_6639,N_6663);
nand U18392 (N_18392,N_10025,N_7488);
xor U18393 (N_18393,N_6498,N_8173);
and U18394 (N_18394,N_12279,N_6602);
nand U18395 (N_18395,N_7971,N_7461);
nand U18396 (N_18396,N_8621,N_10894);
and U18397 (N_18397,N_7588,N_9615);
nor U18398 (N_18398,N_6606,N_6548);
xor U18399 (N_18399,N_6921,N_8590);
or U18400 (N_18400,N_9163,N_9774);
and U18401 (N_18401,N_12357,N_7275);
xnor U18402 (N_18402,N_10299,N_6484);
and U18403 (N_18403,N_9212,N_10891);
nor U18404 (N_18404,N_10629,N_8298);
and U18405 (N_18405,N_11439,N_9549);
nor U18406 (N_18406,N_11399,N_9990);
nand U18407 (N_18407,N_8315,N_12049);
nor U18408 (N_18408,N_6837,N_12482);
xnor U18409 (N_18409,N_9804,N_11815);
nand U18410 (N_18410,N_9864,N_9524);
and U18411 (N_18411,N_7113,N_12342);
and U18412 (N_18412,N_10225,N_12194);
nor U18413 (N_18413,N_12422,N_11291);
or U18414 (N_18414,N_10145,N_9137);
nand U18415 (N_18415,N_6531,N_6792);
nand U18416 (N_18416,N_12073,N_10314);
nor U18417 (N_18417,N_11659,N_9339);
nand U18418 (N_18418,N_10473,N_10274);
xor U18419 (N_18419,N_8326,N_9670);
and U18420 (N_18420,N_7491,N_10391);
nor U18421 (N_18421,N_8977,N_11301);
and U18422 (N_18422,N_12416,N_11634);
nor U18423 (N_18423,N_10690,N_12073);
nand U18424 (N_18424,N_8467,N_6374);
xor U18425 (N_18425,N_9844,N_9286);
xor U18426 (N_18426,N_6949,N_9673);
nand U18427 (N_18427,N_10729,N_8932);
xnor U18428 (N_18428,N_12461,N_9383);
nor U18429 (N_18429,N_7250,N_7328);
and U18430 (N_18430,N_8888,N_12023);
nor U18431 (N_18431,N_8142,N_8538);
or U18432 (N_18432,N_10655,N_11209);
xnor U18433 (N_18433,N_10863,N_9753);
and U18434 (N_18434,N_8107,N_12309);
nor U18435 (N_18435,N_7315,N_8346);
nand U18436 (N_18436,N_11963,N_10355);
or U18437 (N_18437,N_8845,N_9617);
and U18438 (N_18438,N_9433,N_12481);
or U18439 (N_18439,N_6947,N_8676);
and U18440 (N_18440,N_12095,N_9933);
nand U18441 (N_18441,N_7220,N_7152);
nor U18442 (N_18442,N_12082,N_10067);
or U18443 (N_18443,N_10468,N_12107);
and U18444 (N_18444,N_11989,N_10347);
xnor U18445 (N_18445,N_11051,N_9373);
xor U18446 (N_18446,N_8443,N_11001);
nor U18447 (N_18447,N_9452,N_7148);
and U18448 (N_18448,N_11756,N_7495);
and U18449 (N_18449,N_11061,N_8907);
nand U18450 (N_18450,N_10411,N_11419);
nor U18451 (N_18451,N_6469,N_9245);
xor U18452 (N_18452,N_7754,N_11567);
or U18453 (N_18453,N_9654,N_9531);
or U18454 (N_18454,N_9418,N_9747);
xor U18455 (N_18455,N_8687,N_11489);
and U18456 (N_18456,N_8494,N_7683);
and U18457 (N_18457,N_9251,N_10949);
or U18458 (N_18458,N_11245,N_9195);
nor U18459 (N_18459,N_10256,N_10563);
nor U18460 (N_18460,N_11642,N_7593);
or U18461 (N_18461,N_7338,N_8098);
nand U18462 (N_18462,N_11253,N_10989);
and U18463 (N_18463,N_12468,N_11848);
or U18464 (N_18464,N_9236,N_9096);
nor U18465 (N_18465,N_10303,N_10149);
xor U18466 (N_18466,N_9464,N_8971);
or U18467 (N_18467,N_10330,N_12486);
nor U18468 (N_18468,N_8448,N_10128);
and U18469 (N_18469,N_9669,N_9182);
and U18470 (N_18470,N_9317,N_8781);
nor U18471 (N_18471,N_11393,N_9318);
and U18472 (N_18472,N_7424,N_6397);
and U18473 (N_18473,N_11006,N_10004);
nand U18474 (N_18474,N_9921,N_6668);
nor U18475 (N_18475,N_7815,N_8185);
nor U18476 (N_18476,N_12338,N_7777);
xor U18477 (N_18477,N_9194,N_12407);
nand U18478 (N_18478,N_10221,N_9534);
and U18479 (N_18479,N_6322,N_11079);
nor U18480 (N_18480,N_11631,N_6423);
xnor U18481 (N_18481,N_11378,N_8996);
or U18482 (N_18482,N_7619,N_7042);
and U18483 (N_18483,N_8892,N_6478);
and U18484 (N_18484,N_10059,N_7757);
nand U18485 (N_18485,N_8680,N_8467);
or U18486 (N_18486,N_9737,N_6349);
or U18487 (N_18487,N_7485,N_7569);
nor U18488 (N_18488,N_8961,N_6485);
or U18489 (N_18489,N_11898,N_9751);
nand U18490 (N_18490,N_8089,N_6940);
xnor U18491 (N_18491,N_6322,N_11953);
or U18492 (N_18492,N_6422,N_8311);
xor U18493 (N_18493,N_7994,N_8394);
nand U18494 (N_18494,N_9246,N_6757);
and U18495 (N_18495,N_9702,N_9675);
or U18496 (N_18496,N_11436,N_9503);
and U18497 (N_18497,N_9712,N_11984);
nand U18498 (N_18498,N_9739,N_9965);
and U18499 (N_18499,N_6666,N_9172);
nand U18500 (N_18500,N_12203,N_7289);
and U18501 (N_18501,N_8919,N_7327);
nor U18502 (N_18502,N_8239,N_11853);
or U18503 (N_18503,N_10120,N_9274);
nand U18504 (N_18504,N_12279,N_12397);
xor U18505 (N_18505,N_10440,N_10399);
and U18506 (N_18506,N_12132,N_6544);
nor U18507 (N_18507,N_7800,N_11111);
nand U18508 (N_18508,N_10718,N_9584);
nor U18509 (N_18509,N_7928,N_6530);
nor U18510 (N_18510,N_6787,N_8113);
or U18511 (N_18511,N_9402,N_8114);
xnor U18512 (N_18512,N_9287,N_7506);
nor U18513 (N_18513,N_12391,N_10335);
nor U18514 (N_18514,N_12402,N_10256);
nand U18515 (N_18515,N_12350,N_10545);
nand U18516 (N_18516,N_9777,N_7504);
and U18517 (N_18517,N_10068,N_6271);
and U18518 (N_18518,N_11374,N_8384);
nand U18519 (N_18519,N_7522,N_8445);
xor U18520 (N_18520,N_10822,N_8150);
and U18521 (N_18521,N_6333,N_8949);
nor U18522 (N_18522,N_6367,N_6401);
nor U18523 (N_18523,N_11803,N_10938);
xor U18524 (N_18524,N_8907,N_7891);
or U18525 (N_18525,N_8069,N_9116);
and U18526 (N_18526,N_10191,N_6465);
nand U18527 (N_18527,N_10212,N_12281);
nand U18528 (N_18528,N_10456,N_12042);
or U18529 (N_18529,N_9825,N_9587);
xor U18530 (N_18530,N_7188,N_8277);
and U18531 (N_18531,N_8326,N_10507);
nor U18532 (N_18532,N_7250,N_7628);
or U18533 (N_18533,N_9738,N_6803);
and U18534 (N_18534,N_11734,N_10464);
nand U18535 (N_18535,N_11752,N_9898);
nand U18536 (N_18536,N_6386,N_10988);
or U18537 (N_18537,N_7229,N_7265);
and U18538 (N_18538,N_8472,N_10343);
xnor U18539 (N_18539,N_8258,N_12365);
nor U18540 (N_18540,N_10214,N_7053);
or U18541 (N_18541,N_6573,N_7261);
and U18542 (N_18542,N_9100,N_7010);
nand U18543 (N_18543,N_6479,N_10387);
or U18544 (N_18544,N_6385,N_8283);
nand U18545 (N_18545,N_8535,N_12288);
and U18546 (N_18546,N_9230,N_12000);
xnor U18547 (N_18547,N_6775,N_10746);
and U18548 (N_18548,N_6447,N_12333);
nor U18549 (N_18549,N_6939,N_11736);
and U18550 (N_18550,N_10237,N_6942);
xnor U18551 (N_18551,N_11700,N_7707);
nand U18552 (N_18552,N_9760,N_8970);
nor U18553 (N_18553,N_7323,N_8379);
nor U18554 (N_18554,N_9831,N_7135);
nand U18555 (N_18555,N_9544,N_8668);
xnor U18556 (N_18556,N_12481,N_11096);
or U18557 (N_18557,N_8769,N_11396);
xor U18558 (N_18558,N_11440,N_9743);
and U18559 (N_18559,N_6753,N_11657);
xnor U18560 (N_18560,N_11891,N_9458);
nand U18561 (N_18561,N_9715,N_11330);
or U18562 (N_18562,N_10717,N_6766);
xnor U18563 (N_18563,N_12179,N_10956);
xnor U18564 (N_18564,N_7126,N_7236);
nor U18565 (N_18565,N_7879,N_11766);
or U18566 (N_18566,N_12398,N_8462);
and U18567 (N_18567,N_7618,N_6329);
or U18568 (N_18568,N_6465,N_9868);
xor U18569 (N_18569,N_10917,N_7044);
nand U18570 (N_18570,N_6474,N_7744);
nor U18571 (N_18571,N_7197,N_12325);
and U18572 (N_18572,N_11644,N_10873);
and U18573 (N_18573,N_9269,N_9588);
or U18574 (N_18574,N_6799,N_10034);
nor U18575 (N_18575,N_8658,N_11980);
or U18576 (N_18576,N_10080,N_8898);
xnor U18577 (N_18577,N_9716,N_8173);
nand U18578 (N_18578,N_8953,N_11448);
or U18579 (N_18579,N_6695,N_7133);
xnor U18580 (N_18580,N_9260,N_9672);
and U18581 (N_18581,N_9167,N_11901);
xnor U18582 (N_18582,N_11924,N_9600);
nor U18583 (N_18583,N_12274,N_12353);
or U18584 (N_18584,N_8723,N_11489);
nor U18585 (N_18585,N_10120,N_7552);
or U18586 (N_18586,N_7522,N_7516);
nand U18587 (N_18587,N_10409,N_10936);
nor U18588 (N_18588,N_8604,N_7608);
nor U18589 (N_18589,N_8136,N_11572);
nand U18590 (N_18590,N_11580,N_7953);
xor U18591 (N_18591,N_11184,N_10667);
xor U18592 (N_18592,N_8928,N_10526);
nand U18593 (N_18593,N_8613,N_11190);
or U18594 (N_18594,N_9076,N_7235);
nor U18595 (N_18595,N_10401,N_11403);
nor U18596 (N_18596,N_6634,N_9560);
nand U18597 (N_18597,N_8599,N_10744);
nor U18598 (N_18598,N_9611,N_10512);
and U18599 (N_18599,N_7348,N_8697);
nand U18600 (N_18600,N_11610,N_9478);
xor U18601 (N_18601,N_11148,N_6265);
or U18602 (N_18602,N_10317,N_10291);
xor U18603 (N_18603,N_7543,N_8048);
nand U18604 (N_18604,N_12217,N_12165);
xnor U18605 (N_18605,N_7579,N_11440);
nor U18606 (N_18606,N_9557,N_10034);
or U18607 (N_18607,N_8624,N_9233);
or U18608 (N_18608,N_12495,N_8277);
and U18609 (N_18609,N_9778,N_12316);
xnor U18610 (N_18610,N_11838,N_10816);
and U18611 (N_18611,N_7820,N_12348);
nor U18612 (N_18612,N_10390,N_10236);
and U18613 (N_18613,N_6818,N_7676);
or U18614 (N_18614,N_6533,N_11591);
or U18615 (N_18615,N_8101,N_11302);
xor U18616 (N_18616,N_7398,N_11929);
or U18617 (N_18617,N_11258,N_8236);
nand U18618 (N_18618,N_10971,N_9046);
nor U18619 (N_18619,N_10170,N_9014);
or U18620 (N_18620,N_8247,N_8413);
nand U18621 (N_18621,N_8506,N_8718);
xnor U18622 (N_18622,N_8838,N_7940);
nand U18623 (N_18623,N_12262,N_6574);
or U18624 (N_18624,N_11332,N_7164);
or U18625 (N_18625,N_10628,N_10936);
nand U18626 (N_18626,N_7374,N_8027);
or U18627 (N_18627,N_11451,N_6663);
nor U18628 (N_18628,N_12117,N_7959);
or U18629 (N_18629,N_10204,N_12215);
nor U18630 (N_18630,N_8161,N_12408);
nand U18631 (N_18631,N_11281,N_10963);
nand U18632 (N_18632,N_8838,N_6439);
nand U18633 (N_18633,N_9374,N_8055);
nor U18634 (N_18634,N_8806,N_10016);
xor U18635 (N_18635,N_9661,N_8119);
nand U18636 (N_18636,N_7157,N_8862);
or U18637 (N_18637,N_8144,N_7627);
xnor U18638 (N_18638,N_11171,N_10941);
nor U18639 (N_18639,N_11464,N_11707);
nand U18640 (N_18640,N_8724,N_6551);
nor U18641 (N_18641,N_9456,N_6721);
nand U18642 (N_18642,N_8926,N_6758);
or U18643 (N_18643,N_9038,N_10588);
and U18644 (N_18644,N_10505,N_7084);
or U18645 (N_18645,N_10593,N_11401);
nand U18646 (N_18646,N_7874,N_11849);
and U18647 (N_18647,N_11421,N_7997);
or U18648 (N_18648,N_6275,N_10648);
or U18649 (N_18649,N_6645,N_10942);
or U18650 (N_18650,N_8647,N_11480);
and U18651 (N_18651,N_10021,N_6791);
and U18652 (N_18652,N_9412,N_9732);
nand U18653 (N_18653,N_11643,N_7083);
xnor U18654 (N_18654,N_11892,N_8998);
or U18655 (N_18655,N_7297,N_11888);
and U18656 (N_18656,N_12318,N_11384);
nand U18657 (N_18657,N_8965,N_10148);
xnor U18658 (N_18658,N_6688,N_8148);
nand U18659 (N_18659,N_8596,N_6530);
and U18660 (N_18660,N_11209,N_8847);
or U18661 (N_18661,N_11535,N_10730);
and U18662 (N_18662,N_8781,N_6509);
xor U18663 (N_18663,N_7671,N_8826);
nor U18664 (N_18664,N_8919,N_8756);
nand U18665 (N_18665,N_12013,N_10105);
nand U18666 (N_18666,N_9701,N_10358);
or U18667 (N_18667,N_10072,N_10365);
nor U18668 (N_18668,N_12230,N_10571);
or U18669 (N_18669,N_9293,N_7843);
nand U18670 (N_18670,N_10501,N_10624);
nand U18671 (N_18671,N_10534,N_11599);
and U18672 (N_18672,N_9887,N_11363);
and U18673 (N_18673,N_12056,N_11410);
and U18674 (N_18674,N_9242,N_6651);
or U18675 (N_18675,N_6681,N_7503);
or U18676 (N_18676,N_6922,N_11359);
nor U18677 (N_18677,N_7872,N_11339);
and U18678 (N_18678,N_10505,N_11762);
xnor U18679 (N_18679,N_6596,N_10702);
nand U18680 (N_18680,N_11554,N_9727);
and U18681 (N_18681,N_8197,N_10670);
nor U18682 (N_18682,N_12281,N_11388);
nand U18683 (N_18683,N_7184,N_7954);
nand U18684 (N_18684,N_9350,N_11167);
nor U18685 (N_18685,N_10372,N_8243);
or U18686 (N_18686,N_9678,N_10183);
nand U18687 (N_18687,N_7176,N_6984);
and U18688 (N_18688,N_7169,N_12449);
nand U18689 (N_18689,N_9264,N_8716);
xnor U18690 (N_18690,N_12033,N_8926);
xor U18691 (N_18691,N_8895,N_10126);
xor U18692 (N_18692,N_10613,N_8269);
or U18693 (N_18693,N_11940,N_8955);
or U18694 (N_18694,N_9309,N_10355);
nor U18695 (N_18695,N_11071,N_10804);
xor U18696 (N_18696,N_7438,N_9075);
and U18697 (N_18697,N_10134,N_10715);
nor U18698 (N_18698,N_8092,N_10436);
nand U18699 (N_18699,N_9556,N_12437);
or U18700 (N_18700,N_7875,N_10403);
and U18701 (N_18701,N_6572,N_11091);
nor U18702 (N_18702,N_8204,N_8402);
nand U18703 (N_18703,N_8473,N_8304);
nand U18704 (N_18704,N_6752,N_8941);
xor U18705 (N_18705,N_11489,N_9933);
nor U18706 (N_18706,N_12184,N_12010);
or U18707 (N_18707,N_8482,N_9508);
nand U18708 (N_18708,N_9026,N_6847);
nor U18709 (N_18709,N_9398,N_10592);
and U18710 (N_18710,N_8536,N_12443);
nor U18711 (N_18711,N_11565,N_8978);
nand U18712 (N_18712,N_8026,N_8507);
xnor U18713 (N_18713,N_9934,N_6348);
nand U18714 (N_18714,N_11466,N_8516);
and U18715 (N_18715,N_8658,N_6818);
nand U18716 (N_18716,N_8778,N_8757);
or U18717 (N_18717,N_11985,N_6704);
or U18718 (N_18718,N_11632,N_11723);
nand U18719 (N_18719,N_7469,N_8185);
xnor U18720 (N_18720,N_8383,N_8403);
nand U18721 (N_18721,N_8477,N_10779);
nand U18722 (N_18722,N_6564,N_7194);
and U18723 (N_18723,N_7688,N_8099);
nand U18724 (N_18724,N_9239,N_11107);
nand U18725 (N_18725,N_11323,N_12068);
nor U18726 (N_18726,N_6922,N_12269);
nand U18727 (N_18727,N_11116,N_11259);
and U18728 (N_18728,N_8371,N_9987);
and U18729 (N_18729,N_9004,N_12207);
and U18730 (N_18730,N_7834,N_7201);
xor U18731 (N_18731,N_8149,N_7879);
xnor U18732 (N_18732,N_12486,N_7209);
nor U18733 (N_18733,N_10635,N_11802);
and U18734 (N_18734,N_8693,N_12025);
xnor U18735 (N_18735,N_9285,N_6356);
and U18736 (N_18736,N_9735,N_11538);
nand U18737 (N_18737,N_11799,N_12182);
and U18738 (N_18738,N_9127,N_10802);
nand U18739 (N_18739,N_9693,N_7904);
xnor U18740 (N_18740,N_9144,N_12223);
and U18741 (N_18741,N_10845,N_10383);
or U18742 (N_18742,N_12263,N_10171);
xnor U18743 (N_18743,N_11445,N_7096);
xnor U18744 (N_18744,N_6802,N_11676);
and U18745 (N_18745,N_8889,N_11819);
nand U18746 (N_18746,N_9274,N_11818);
nor U18747 (N_18747,N_7813,N_10313);
nor U18748 (N_18748,N_12084,N_6276);
nand U18749 (N_18749,N_10978,N_9355);
nor U18750 (N_18750,N_14573,N_18333);
nor U18751 (N_18751,N_12848,N_16480);
and U18752 (N_18752,N_13902,N_15736);
or U18753 (N_18753,N_17208,N_14563);
nor U18754 (N_18754,N_16551,N_13868);
nor U18755 (N_18755,N_13110,N_17973);
nand U18756 (N_18756,N_18012,N_13936);
or U18757 (N_18757,N_15889,N_15454);
and U18758 (N_18758,N_14999,N_13627);
nor U18759 (N_18759,N_15174,N_16673);
xnor U18760 (N_18760,N_13032,N_13462);
xnor U18761 (N_18761,N_17367,N_17840);
nand U18762 (N_18762,N_17866,N_15432);
and U18763 (N_18763,N_13607,N_12938);
nand U18764 (N_18764,N_17528,N_13702);
or U18765 (N_18765,N_14387,N_18003);
or U18766 (N_18766,N_16460,N_12648);
nand U18767 (N_18767,N_15412,N_13280);
xor U18768 (N_18768,N_16027,N_15834);
nor U18769 (N_18769,N_16071,N_18555);
or U18770 (N_18770,N_13974,N_18182);
or U18771 (N_18771,N_16465,N_14018);
nand U18772 (N_18772,N_13017,N_18444);
xnor U18773 (N_18773,N_16309,N_18603);
xor U18774 (N_18774,N_16607,N_17689);
xnor U18775 (N_18775,N_15384,N_14155);
nor U18776 (N_18776,N_14161,N_12637);
xor U18777 (N_18777,N_14086,N_13578);
nor U18778 (N_18778,N_15789,N_13687);
xor U18779 (N_18779,N_17307,N_12829);
nand U18780 (N_18780,N_16381,N_16036);
nand U18781 (N_18781,N_14858,N_16701);
or U18782 (N_18782,N_14898,N_14566);
nand U18783 (N_18783,N_17662,N_18184);
xnor U18784 (N_18784,N_15397,N_18623);
nor U18785 (N_18785,N_18339,N_17606);
or U18786 (N_18786,N_13231,N_15415);
or U18787 (N_18787,N_14063,N_14290);
nor U18788 (N_18788,N_14066,N_13637);
xor U18789 (N_18789,N_14552,N_13805);
and U18790 (N_18790,N_15781,N_14405);
xnor U18791 (N_18791,N_12901,N_14150);
nor U18792 (N_18792,N_13363,N_16155);
nand U18793 (N_18793,N_18485,N_14512);
xnor U18794 (N_18794,N_17856,N_16292);
xor U18795 (N_18795,N_13256,N_17389);
nor U18796 (N_18796,N_13931,N_12913);
nand U18797 (N_18797,N_17813,N_12633);
and U18798 (N_18798,N_16569,N_17760);
and U18799 (N_18799,N_17570,N_18427);
and U18800 (N_18800,N_16703,N_18353);
nor U18801 (N_18801,N_14019,N_13755);
nand U18802 (N_18802,N_17568,N_17068);
xor U18803 (N_18803,N_16386,N_15147);
nor U18804 (N_18804,N_12917,N_15217);
or U18805 (N_18805,N_15619,N_12777);
nand U18806 (N_18806,N_17905,N_13618);
nand U18807 (N_18807,N_17296,N_14836);
nor U18808 (N_18808,N_13246,N_16019);
xor U18809 (N_18809,N_14281,N_17516);
nor U18810 (N_18810,N_15051,N_14546);
or U18811 (N_18811,N_14036,N_16267);
xnor U18812 (N_18812,N_13003,N_12998);
nor U18813 (N_18813,N_13398,N_17818);
nor U18814 (N_18814,N_14435,N_17586);
nand U18815 (N_18815,N_14831,N_14645);
xnor U18816 (N_18816,N_13348,N_16960);
xor U18817 (N_18817,N_13123,N_14864);
and U18818 (N_18818,N_16759,N_18356);
nand U18819 (N_18819,N_14445,N_17217);
and U18820 (N_18820,N_17725,N_12719);
nor U18821 (N_18821,N_12755,N_17401);
nor U18822 (N_18822,N_14096,N_17327);
or U18823 (N_18823,N_18556,N_16878);
nand U18824 (N_18824,N_14970,N_16170);
xnor U18825 (N_18825,N_13365,N_14215);
and U18826 (N_18826,N_14583,N_15104);
or U18827 (N_18827,N_17158,N_18710);
or U18828 (N_18828,N_12978,N_16418);
nand U18829 (N_18829,N_15727,N_16814);
nand U18830 (N_18830,N_14298,N_17742);
nor U18831 (N_18831,N_17466,N_15742);
nor U18832 (N_18832,N_15021,N_12532);
and U18833 (N_18833,N_16275,N_15509);
or U18834 (N_18834,N_14111,N_16316);
or U18835 (N_18835,N_15676,N_17686);
or U18836 (N_18836,N_16877,N_17620);
xnor U18837 (N_18837,N_17272,N_13274);
xor U18838 (N_18838,N_14752,N_16149);
and U18839 (N_18839,N_13303,N_13068);
or U18840 (N_18840,N_14853,N_13729);
or U18841 (N_18841,N_13076,N_14536);
and U18842 (N_18842,N_18404,N_12773);
nand U18843 (N_18843,N_14146,N_14109);
and U18844 (N_18844,N_17242,N_14771);
or U18845 (N_18845,N_13440,N_13160);
xor U18846 (N_18846,N_16707,N_14487);
nor U18847 (N_18847,N_13233,N_16307);
or U18848 (N_18848,N_16457,N_13675);
nand U18849 (N_18849,N_16471,N_14083);
nand U18850 (N_18850,N_16745,N_16976);
xor U18851 (N_18851,N_17752,N_17429);
and U18852 (N_18852,N_15242,N_13523);
or U18853 (N_18853,N_16810,N_18539);
and U18854 (N_18854,N_18601,N_13167);
or U18855 (N_18855,N_16073,N_14924);
or U18856 (N_18856,N_16839,N_14555);
nor U18857 (N_18857,N_15106,N_16962);
and U18858 (N_18858,N_16014,N_13946);
and U18859 (N_18859,N_16215,N_12501);
nand U18860 (N_18860,N_18092,N_15478);
or U18861 (N_18861,N_18121,N_17954);
and U18862 (N_18862,N_13991,N_13640);
xor U18863 (N_18863,N_15142,N_13836);
and U18864 (N_18864,N_17665,N_14088);
and U18865 (N_18865,N_15132,N_14455);
and U18866 (N_18866,N_17558,N_15643);
nand U18867 (N_18867,N_14067,N_16604);
nand U18868 (N_18868,N_12572,N_18533);
or U18869 (N_18869,N_12749,N_17613);
and U18870 (N_18870,N_14055,N_14769);
nand U18871 (N_18871,N_17065,N_15350);
xnor U18872 (N_18872,N_12709,N_13494);
nor U18873 (N_18873,N_13404,N_17540);
nand U18874 (N_18874,N_12950,N_13043);
or U18875 (N_18875,N_12527,N_15292);
and U18876 (N_18876,N_15624,N_14490);
nor U18877 (N_18877,N_14903,N_13548);
nand U18878 (N_18878,N_14556,N_17678);
xor U18879 (N_18879,N_12604,N_15832);
and U18880 (N_18880,N_15044,N_17399);
nand U18881 (N_18881,N_13381,N_16077);
xnor U18882 (N_18882,N_12645,N_14190);
nor U18883 (N_18883,N_16299,N_16761);
nand U18884 (N_18884,N_18015,N_15651);
and U18885 (N_18885,N_17358,N_12934);
nand U18886 (N_18886,N_17845,N_16521);
and U18887 (N_18887,N_12561,N_13859);
nor U18888 (N_18888,N_15960,N_14333);
and U18889 (N_18889,N_12549,N_13757);
or U18890 (N_18890,N_17029,N_15869);
nor U18891 (N_18891,N_14976,N_15112);
xnor U18892 (N_18892,N_15237,N_18391);
and U18893 (N_18893,N_17857,N_14632);
nand U18894 (N_18894,N_18004,N_17290);
and U18895 (N_18895,N_17907,N_14906);
xnor U18896 (N_18896,N_16995,N_13832);
nand U18897 (N_18897,N_15860,N_15436);
xor U18898 (N_18898,N_16766,N_18265);
and U18899 (N_18899,N_12518,N_16776);
nor U18900 (N_18900,N_14242,N_17473);
nor U18901 (N_18901,N_18298,N_18136);
xnor U18902 (N_18902,N_14131,N_12568);
nor U18903 (N_18903,N_18660,N_16515);
xor U18904 (N_18904,N_12614,N_15442);
nor U18905 (N_18905,N_16988,N_17387);
nand U18906 (N_18906,N_18511,N_13589);
nor U18907 (N_18907,N_15260,N_13271);
nand U18908 (N_18908,N_16007,N_16142);
nand U18909 (N_18909,N_16946,N_13482);
xor U18910 (N_18910,N_13185,N_18357);
xor U18911 (N_18911,N_18156,N_17163);
nor U18912 (N_18912,N_18747,N_15492);
and U18913 (N_18913,N_13150,N_17007);
nor U18914 (N_18914,N_13019,N_13709);
nor U18915 (N_18915,N_13808,N_12703);
or U18916 (N_18916,N_18477,N_15066);
xor U18917 (N_18917,N_12753,N_15737);
xor U18918 (N_18918,N_13152,N_13560);
and U18919 (N_18919,N_18396,N_12790);
nand U18920 (N_18920,N_13787,N_14670);
or U18921 (N_18921,N_15055,N_16039);
or U18922 (N_18922,N_17582,N_18654);
nand U18923 (N_18923,N_17045,N_13154);
or U18924 (N_18924,N_17566,N_14317);
xor U18925 (N_18925,N_17616,N_17462);
nand U18926 (N_18926,N_17599,N_12575);
and U18927 (N_18927,N_15456,N_17572);
nand U18928 (N_18928,N_17345,N_15855);
and U18929 (N_18929,N_16531,N_18175);
nand U18930 (N_18930,N_15351,N_12973);
nand U18931 (N_18931,N_13432,N_12655);
nor U18932 (N_18932,N_13529,N_18048);
or U18933 (N_18933,N_14646,N_13876);
and U18934 (N_18934,N_15808,N_16028);
nor U18935 (N_18935,N_16102,N_14309);
and U18936 (N_18936,N_17079,N_16268);
xor U18937 (N_18937,N_16391,N_18108);
and U18938 (N_18938,N_13530,N_12706);
nand U18939 (N_18939,N_12885,N_18042);
nor U18940 (N_18940,N_17712,N_18640);
xor U18941 (N_18941,N_14344,N_12944);
nor U18942 (N_18942,N_15959,N_16091);
nor U18943 (N_18943,N_18388,N_16291);
xnor U18944 (N_18944,N_17412,N_16940);
nor U18945 (N_18945,N_15891,N_16263);
xor U18946 (N_18946,N_14894,N_15874);
nor U18947 (N_18947,N_16025,N_15410);
nor U18948 (N_18948,N_15884,N_16499);
nor U18949 (N_18949,N_14790,N_15375);
nand U18950 (N_18950,N_14950,N_14787);
nor U18951 (N_18951,N_13905,N_17977);
xor U18952 (N_18952,N_15148,N_13087);
or U18953 (N_18953,N_12810,N_15581);
or U18954 (N_18954,N_12914,N_14829);
nor U18955 (N_18955,N_13665,N_17078);
or U18956 (N_18956,N_16419,N_18240);
and U18957 (N_18957,N_14712,N_16433);
and U18958 (N_18958,N_14102,N_14401);
or U18959 (N_18959,N_14496,N_18010);
nor U18960 (N_18960,N_15815,N_13466);
and U18961 (N_18961,N_12607,N_16449);
xor U18962 (N_18962,N_13028,N_14998);
and U18963 (N_18963,N_13985,N_17097);
nor U18964 (N_18964,N_14620,N_18118);
xnor U18965 (N_18965,N_14765,N_12688);
nand U18966 (N_18966,N_15023,N_13416);
nor U18967 (N_18967,N_16070,N_18348);
xor U18968 (N_18968,N_17346,N_12821);
and U18969 (N_18969,N_14157,N_13006);
or U18970 (N_18970,N_12783,N_13568);
nor U18971 (N_18971,N_15034,N_18064);
nand U18972 (N_18972,N_14029,N_18061);
nand U18973 (N_18973,N_17793,N_13429);
xor U18974 (N_18974,N_12720,N_16793);
or U18975 (N_18975,N_12727,N_17869);
nor U18976 (N_18976,N_13691,N_13206);
and U18977 (N_18977,N_16675,N_15419);
nor U18978 (N_18978,N_17251,N_16167);
xor U18979 (N_18979,N_13312,N_14817);
and U18980 (N_18980,N_17289,N_15248);
xnor U18981 (N_18981,N_18343,N_12931);
xor U18982 (N_18982,N_18503,N_16127);
xor U18983 (N_18983,N_13008,N_17597);
xnor U18984 (N_18984,N_17180,N_17142);
nor U18985 (N_18985,N_14417,N_12666);
or U18986 (N_18986,N_14235,N_13543);
nor U18987 (N_18987,N_17416,N_15940);
nor U18988 (N_18988,N_15963,N_15511);
nor U18989 (N_18989,N_15853,N_13368);
xor U18990 (N_18990,N_17318,N_17930);
nand U18991 (N_18991,N_12778,N_15517);
nor U18992 (N_18992,N_16430,N_13712);
nand U18993 (N_18993,N_15786,N_15173);
nand U18994 (N_18994,N_15449,N_13510);
or U18995 (N_18995,N_13767,N_18689);
xnor U18996 (N_18996,N_18544,N_12511);
and U18997 (N_18997,N_13881,N_13141);
or U18998 (N_18998,N_15917,N_17967);
and U18999 (N_18999,N_16594,N_18472);
xor U19000 (N_19000,N_16377,N_12864);
or U19001 (N_19001,N_12605,N_18505);
nor U19002 (N_19002,N_15747,N_18664);
and U19003 (N_19003,N_17109,N_12805);
or U19004 (N_19004,N_14814,N_18593);
or U19005 (N_19005,N_15216,N_13388);
xnor U19006 (N_19006,N_15675,N_17567);
and U19007 (N_19007,N_15659,N_13502);
and U19008 (N_19008,N_16547,N_15776);
xor U19009 (N_19009,N_16722,N_16854);
xor U19010 (N_19010,N_17831,N_16772);
or U19011 (N_19011,N_13288,N_17441);
and U19012 (N_19012,N_18540,N_16815);
nand U19013 (N_19013,N_18200,N_14747);
and U19014 (N_19014,N_15613,N_14100);
nor U19015 (N_19015,N_14574,N_18095);
xnor U19016 (N_19016,N_17361,N_16914);
nand U19017 (N_19017,N_16646,N_15686);
and U19018 (N_19018,N_18154,N_15083);
or U19019 (N_19019,N_12508,N_14915);
nor U19020 (N_19020,N_17673,N_16930);
nand U19021 (N_19021,N_13158,N_15561);
or U19022 (N_19022,N_15238,N_15356);
nor U19023 (N_19023,N_13234,N_17483);
and U19024 (N_19024,N_12756,N_16535);
or U19025 (N_19025,N_16483,N_17971);
nand U19026 (N_19026,N_17319,N_12760);
nand U19027 (N_19027,N_13020,N_17283);
xnor U19028 (N_19028,N_16000,N_17796);
xnor U19029 (N_19029,N_13596,N_13677);
nand U19030 (N_19030,N_17199,N_14068);
and U19031 (N_19031,N_14314,N_16736);
xnor U19032 (N_19032,N_13603,N_12853);
xor U19033 (N_19033,N_15510,N_15980);
or U19034 (N_19034,N_14900,N_16851);
xor U19035 (N_19035,N_13034,N_16875);
nand U19036 (N_19036,N_14039,N_16978);
and U19037 (N_19037,N_18523,N_17975);
xnor U19038 (N_19038,N_14085,N_17108);
and U19039 (N_19039,N_18681,N_15470);
or U19040 (N_19040,N_14721,N_18104);
or U19041 (N_19041,N_17415,N_13272);
nor U19042 (N_19042,N_12945,N_12522);
xor U19043 (N_19043,N_17747,N_17000);
or U19044 (N_19044,N_15443,N_14638);
nand U19045 (N_19045,N_18569,N_14237);
nor U19046 (N_19046,N_16208,N_12926);
nand U19047 (N_19047,N_18002,N_13733);
nor U19048 (N_19048,N_18329,N_14193);
and U19049 (N_19049,N_18150,N_15647);
xnor U19050 (N_19050,N_13937,N_15197);
nor U19051 (N_19051,N_17919,N_15764);
xnor U19052 (N_19052,N_18177,N_15153);
and U19053 (N_19053,N_18336,N_15434);
or U19054 (N_19054,N_12535,N_14826);
or U19055 (N_19055,N_16660,N_17368);
nor U19056 (N_19056,N_14069,N_16894);
and U19057 (N_19057,N_13290,N_13044);
xnor U19058 (N_19058,N_12764,N_18442);
or U19059 (N_19059,N_17477,N_17838);
xor U19060 (N_19060,N_13790,N_17578);
xnor U19061 (N_19061,N_17195,N_17829);
nand U19062 (N_19062,N_15017,N_14322);
or U19063 (N_19063,N_16692,N_16934);
nand U19064 (N_19064,N_12576,N_13670);
nor U19065 (N_19065,N_15710,N_14557);
and U19066 (N_19066,N_14611,N_13894);
nor U19067 (N_19067,N_17705,N_17316);
xnor U19068 (N_19068,N_12658,N_13754);
and U19069 (N_19069,N_14470,N_17154);
or U19070 (N_19070,N_18631,N_12712);
nand U19071 (N_19071,N_13250,N_15746);
nand U19072 (N_19072,N_16454,N_14040);
nor U19073 (N_19073,N_18123,N_14818);
or U19074 (N_19074,N_15810,N_15204);
nor U19075 (N_19075,N_14373,N_12767);
or U19076 (N_19076,N_14975,N_14788);
and U19077 (N_19077,N_12502,N_15482);
nor U19078 (N_19078,N_17178,N_12837);
or U19079 (N_19079,N_15868,N_13077);
nor U19080 (N_19080,N_13349,N_14246);
and U19081 (N_19081,N_17347,N_13335);
or U19082 (N_19082,N_17691,N_17336);
and U19083 (N_19083,N_16281,N_16591);
and U19084 (N_19084,N_16785,N_14627);
nand U19085 (N_19085,N_15211,N_13553);
or U19086 (N_19086,N_13503,N_15690);
nor U19087 (N_19087,N_14545,N_14933);
xor U19088 (N_19088,N_16201,N_16754);
and U19089 (N_19089,N_17538,N_15928);
nor U19090 (N_19090,N_14473,N_17481);
nor U19091 (N_19091,N_16219,N_12687);
and U19092 (N_19092,N_17589,N_13140);
nor U19093 (N_19093,N_13258,N_17333);
nor U19094 (N_19094,N_12863,N_12628);
nand U19095 (N_19095,N_14971,N_16026);
xor U19096 (N_19096,N_15180,N_18594);
and U19097 (N_19097,N_13046,N_13093);
nor U19098 (N_19098,N_14597,N_14770);
and U19099 (N_19099,N_14296,N_14554);
and U19100 (N_19100,N_16796,N_15851);
nor U19101 (N_19101,N_17323,N_18328);
nand U19102 (N_19102,N_14139,N_17921);
nor U19103 (N_19103,N_18113,N_16194);
xnor U19104 (N_19104,N_14089,N_16993);
nand U19105 (N_19105,N_13969,N_14682);
xor U19106 (N_19106,N_13444,N_15528);
nand U19107 (N_19107,N_17815,N_15641);
or U19108 (N_19108,N_13725,N_14201);
and U19109 (N_19109,N_13375,N_13809);
or U19110 (N_19110,N_16214,N_13180);
nand U19111 (N_19111,N_15072,N_15912);
and U19112 (N_19112,N_15774,N_18625);
nor U19113 (N_19113,N_18629,N_18393);
nand U19114 (N_19114,N_14378,N_12584);
nor U19115 (N_19115,N_16432,N_18360);
or U19116 (N_19116,N_13564,N_13500);
nand U19117 (N_19117,N_16054,N_15618);
and U19118 (N_19118,N_18284,N_16605);
nor U19119 (N_19119,N_17439,N_15223);
xnor U19120 (N_19120,N_16526,N_17709);
nand U19121 (N_19121,N_17842,N_13883);
nand U19122 (N_19122,N_17761,N_13983);
or U19123 (N_19123,N_17913,N_18155);
nand U19124 (N_19124,N_18675,N_18739);
nor U19125 (N_19125,N_16616,N_15151);
nor U19126 (N_19126,N_14865,N_13166);
xnor U19127 (N_19127,N_16059,N_15467);
or U19128 (N_19128,N_16326,N_15526);
nor U19129 (N_19129,N_14078,N_17833);
xnor U19130 (N_19130,N_13331,N_13639);
nor U19131 (N_19131,N_16100,N_16052);
nor U19132 (N_19132,N_14577,N_13920);
or U19133 (N_19133,N_17153,N_16423);
nor U19134 (N_19134,N_13645,N_17398);
nor U19135 (N_19135,N_18202,N_15672);
xor U19136 (N_19136,N_12947,N_18036);
nand U19137 (N_19137,N_13595,N_15970);
nor U19138 (N_19138,N_14647,N_14600);
and U19139 (N_19139,N_15228,N_14699);
and U19140 (N_19140,N_18137,N_15777);
nand U19141 (N_19141,N_16146,N_15485);
xnor U19142 (N_19142,N_14247,N_17190);
nor U19143 (N_19143,N_17623,N_14441);
and U19144 (N_19144,N_14024,N_18024);
or U19145 (N_19145,N_17261,N_18163);
nand U19146 (N_19146,N_18488,N_16779);
xor U19147 (N_19147,N_14483,N_13664);
xor U19148 (N_19148,N_14974,N_15469);
and U19149 (N_19149,N_15344,N_17775);
nor U19150 (N_19150,N_12716,N_16564);
nor U19151 (N_19151,N_18060,N_16705);
nor U19152 (N_19152,N_15497,N_18090);
nand U19153 (N_19153,N_14634,N_14336);
and U19154 (N_19154,N_16933,N_18377);
and U19155 (N_19155,N_15337,N_14076);
or U19156 (N_19156,N_13407,N_13731);
xnor U19157 (N_19157,N_16967,N_12663);
or U19158 (N_19158,N_15840,N_15165);
and U19159 (N_19159,N_13828,N_14951);
or U19160 (N_19160,N_15437,N_14527);
nand U19161 (N_19161,N_13105,N_12977);
nand U19162 (N_19162,N_16310,N_18234);
or U19163 (N_19163,N_13764,N_16786);
or U19164 (N_19164,N_18126,N_16241);
and U19165 (N_19165,N_16929,N_13644);
nand U19166 (N_19166,N_13345,N_14821);
or U19167 (N_19167,N_18642,N_16282);
nor U19168 (N_19168,N_15172,N_13656);
and U19169 (N_19169,N_15817,N_16013);
xor U19170 (N_19170,N_17010,N_15711);
and U19171 (N_19171,N_16046,N_13916);
nor U19172 (N_19172,N_18268,N_13509);
nor U19173 (N_19173,N_12940,N_17819);
nor U19174 (N_19174,N_13861,N_13948);
and U19175 (N_19175,N_12570,N_17286);
or U19176 (N_19176,N_14371,N_12526);
or U19177 (N_19177,N_12963,N_13489);
nand U19178 (N_19178,N_12758,N_18553);
xnor U19179 (N_19179,N_13322,N_14839);
or U19180 (N_19180,N_13377,N_13875);
nand U19181 (N_19181,N_13865,N_18078);
xnor U19182 (N_19182,N_15290,N_13172);
xor U19183 (N_19183,N_17989,N_18471);
xor U19184 (N_19184,N_15265,N_15504);
or U19185 (N_19185,N_18321,N_13278);
and U19186 (N_19186,N_14129,N_14118);
xnor U19187 (N_19187,N_16697,N_16235);
nor U19188 (N_19188,N_15957,N_15753);
and U19189 (N_19189,N_17210,N_16597);
nand U19190 (N_19190,N_14538,N_18466);
xnor U19191 (N_19191,N_12521,N_17661);
and U19192 (N_19192,N_18194,N_16205);
or U19193 (N_19193,N_15552,N_13067);
and U19194 (N_19194,N_17472,N_16417);
xnor U19195 (N_19195,N_18606,N_18608);
nand U19196 (N_19196,N_13971,N_13934);
or U19197 (N_19197,N_15187,N_13901);
or U19198 (N_19198,N_14683,N_16051);
xnor U19199 (N_19199,N_15288,N_12620);
nand U19200 (N_19200,N_18167,N_18363);
and U19201 (N_19201,N_18026,N_17018);
or U19202 (N_19202,N_13437,N_18584);
or U19203 (N_19203,N_18487,N_18431);
nand U19204 (N_19204,N_18041,N_15661);
xor U19205 (N_19205,N_14197,N_13434);
xor U19206 (N_19206,N_17248,N_17896);
or U19207 (N_19207,N_13210,N_17063);
nor U19208 (N_19208,N_14204,N_14535);
and U19209 (N_19209,N_16202,N_17402);
and U19210 (N_19210,N_14674,N_15982);
xor U19211 (N_19211,N_15885,N_18248);
nand U19212 (N_19212,N_16809,N_15751);
xnor U19213 (N_19213,N_14677,N_18361);
or U19214 (N_19214,N_13385,N_17161);
or U19215 (N_19215,N_13561,N_14165);
nand U19216 (N_19216,N_16191,N_15579);
and U19217 (N_19217,N_16668,N_13460);
nand U19218 (N_19218,N_15625,N_18469);
and U19219 (N_19219,N_14996,N_13780);
nor U19220 (N_19220,N_15766,N_15176);
or U19221 (N_19221,N_15068,N_12603);
nand U19222 (N_19222,N_18717,N_17436);
nor U19223 (N_19223,N_17554,N_12902);
nand U19224 (N_19224,N_13449,N_13856);
nand U19225 (N_19225,N_16846,N_15287);
or U19226 (N_19226,N_14792,N_16643);
xor U19227 (N_19227,N_18645,N_15493);
or U19228 (N_19228,N_18562,N_17820);
nor U19229 (N_19229,N_18693,N_14003);
nor U19230 (N_19230,N_13533,N_17293);
or U19231 (N_19231,N_13557,N_17996);
nand U19232 (N_19232,N_14099,N_17646);
nor U19233 (N_19233,N_13458,N_18616);
nand U19234 (N_19234,N_14307,N_14700);
nand U19235 (N_19235,N_13559,N_16904);
nand U19236 (N_19236,N_13831,N_18346);
nand U19237 (N_19237,N_17580,N_17379);
nand U19238 (N_19238,N_15206,N_12644);
xor U19239 (N_19239,N_18062,N_13359);
or U19240 (N_19240,N_12673,N_16818);
xnor U19241 (N_19241,N_16990,N_16251);
and U19242 (N_19242,N_18205,N_14572);
nand U19243 (N_19243,N_18014,N_16247);
and U19244 (N_19244,N_18083,N_13211);
nand U19245 (N_19245,N_16507,N_15405);
nand U19246 (N_19246,N_18340,N_14326);
nor U19247 (N_19247,N_15864,N_17268);
or U19248 (N_19248,N_18044,N_13427);
xnor U19249 (N_19249,N_12957,N_13378);
xnor U19250 (N_19250,N_14101,N_14891);
nand U19251 (N_19251,N_12730,N_15146);
nand U19252 (N_19252,N_15945,N_13759);
and U19253 (N_19253,N_12506,N_13193);
xor U19254 (N_19254,N_12548,N_14219);
or U19255 (N_19255,N_16139,N_17933);
nand U19256 (N_19256,N_15650,N_17166);
nor U19257 (N_19257,N_15518,N_15052);
nor U19258 (N_19258,N_17987,N_14457);
nor U19259 (N_19259,N_12700,N_18033);
nand U19260 (N_19260,N_15585,N_16476);
xor U19261 (N_19261,N_17049,N_13218);
or U19262 (N_19262,N_16264,N_17810);
nand U19263 (N_19263,N_16301,N_13111);
or U19264 (N_19264,N_16966,N_12779);
or U19265 (N_19265,N_14436,N_15326);
nand U19266 (N_19266,N_17407,N_17156);
xnor U19267 (N_19267,N_14211,N_15196);
xnor U19268 (N_19268,N_16314,N_14114);
nand U19269 (N_19269,N_14113,N_14888);
or U19270 (N_19270,N_15723,N_15700);
nor U19271 (N_19271,N_17998,N_16548);
nand U19272 (N_19272,N_14684,N_15253);
or U19273 (N_19273,N_12524,N_14753);
and U19274 (N_19274,N_16141,N_12830);
nor U19275 (N_19275,N_15016,N_14628);
xor U19276 (N_19276,N_13129,N_14442);
nand U19277 (N_19277,N_18047,N_14272);
xor U19278 (N_19278,N_17509,N_13041);
or U19279 (N_19279,N_15591,N_16985);
and U19280 (N_19280,N_15322,N_13997);
or U19281 (N_19281,N_16509,N_12857);
or U19282 (N_19282,N_15681,N_15534);
nand U19283 (N_19283,N_16229,N_15439);
nor U19284 (N_19284,N_16343,N_17099);
or U19285 (N_19285,N_15429,N_15827);
and U19286 (N_19286,N_12785,N_18144);
nor U19287 (N_19287,N_15924,N_12724);
or U19288 (N_19288,N_16355,N_13619);
xnor U19289 (N_19289,N_17601,N_15163);
nand U19290 (N_19290,N_17549,N_15655);
nor U19291 (N_19291,N_16357,N_15936);
nor U19292 (N_19292,N_16725,N_15157);
and U19293 (N_19293,N_17562,N_15065);
nand U19294 (N_19294,N_13127,N_18162);
and U19295 (N_19295,N_17759,N_17330);
and U19296 (N_19296,N_13480,N_18452);
xnor U19297 (N_19297,N_17891,N_13397);
nor U19298 (N_19298,N_18592,N_13804);
or U19299 (N_19299,N_14561,N_14617);
nand U19300 (N_19300,N_12916,N_14758);
nand U19301 (N_19301,N_17836,N_16633);
nor U19302 (N_19302,N_15767,N_13491);
and U19303 (N_19303,N_16541,N_14213);
nor U19304 (N_19304,N_15367,N_13414);
xnor U19305 (N_19305,N_14087,N_15822);
nor U19306 (N_19306,N_13657,N_14012);
and U19307 (N_19307,N_12677,N_18085);
or U19308 (N_19308,N_16171,N_16869);
xor U19309 (N_19309,N_14008,N_16936);
or U19310 (N_19310,N_16132,N_12560);
or U19311 (N_19311,N_15161,N_17808);
nand U19312 (N_19312,N_16627,N_12592);
and U19313 (N_19313,N_16802,N_18542);
and U19314 (N_19314,N_17434,N_12831);
nor U19315 (N_19315,N_14722,N_16169);
nand U19316 (N_19316,N_14376,N_16126);
nor U19317 (N_19317,N_18525,N_15348);
nor U19318 (N_19318,N_15839,N_18327);
and U19319 (N_19319,N_17356,N_16719);
nand U19320 (N_19320,N_18632,N_15126);
and U19321 (N_19321,N_13148,N_15630);
nand U19322 (N_19322,N_16678,N_15110);
nor U19323 (N_19323,N_17826,N_13925);
and U19324 (N_19324,N_14230,N_15922);
nor U19325 (N_19325,N_12748,N_16378);
xor U19326 (N_19326,N_14565,N_12500);
nand U19327 (N_19327,N_13768,N_13356);
or U19328 (N_19328,N_15154,N_17993);
xnor U19329 (N_19329,N_15593,N_12669);
nand U19330 (N_19330,N_12589,N_17638);
nand U19331 (N_19331,N_17343,N_15053);
xor U19332 (N_19332,N_16233,N_14729);
or U19333 (N_19333,N_16213,N_17209);
xor U19334 (N_19334,N_13389,N_13992);
or U19335 (N_19335,N_17730,N_17104);
nand U19336 (N_19336,N_18129,N_13009);
nor U19337 (N_19337,N_13518,N_14443);
nor U19338 (N_19338,N_13949,N_12960);
nand U19339 (N_19339,N_17488,N_13428);
nand U19340 (N_19340,N_12976,N_17040);
nand U19341 (N_19341,N_16489,N_14337);
or U19342 (N_19342,N_12598,N_13487);
xor U19343 (N_19343,N_16808,N_15530);
and U19344 (N_19344,N_14588,N_16506);
nor U19345 (N_19345,N_15732,N_18534);
and U19346 (N_19346,N_13134,N_18159);
and U19347 (N_19347,N_17497,N_14453);
nand U19348 (N_19348,N_12995,N_14319);
nor U19349 (N_19349,N_15213,N_14093);
or U19350 (N_19350,N_15575,N_18424);
xnor U19351 (N_19351,N_17344,N_15328);
nor U19352 (N_19352,N_16917,N_18076);
or U19353 (N_19353,N_14988,N_17325);
xnor U19354 (N_19354,N_16832,N_16274);
xor U19355 (N_19355,N_16952,N_18125);
nor U19356 (N_19356,N_13243,N_12555);
nor U19357 (N_19357,N_15977,N_12841);
and U19358 (N_19358,N_17768,N_14756);
nand U19359 (N_19359,N_17183,N_17541);
and U19360 (N_19360,N_17478,N_12824);
nor U19361 (N_19361,N_17608,N_17467);
and U19362 (N_19362,N_18410,N_17471);
nand U19363 (N_19363,N_15658,N_16156);
nand U19364 (N_19364,N_17984,N_14515);
nor U19365 (N_19365,N_17258,N_18103);
and U19366 (N_19366,N_14200,N_13994);
xnor U19367 (N_19367,N_18242,N_16987);
or U19368 (N_19368,N_14509,N_18618);
or U19369 (N_19369,N_18220,N_13203);
xor U19370 (N_19370,N_18145,N_17100);
xor U19371 (N_19371,N_13522,N_12908);
nand U19372 (N_19372,N_15633,N_13366);
or U19373 (N_19373,N_15387,N_12836);
nand U19374 (N_19374,N_12606,N_12967);
nor U19375 (N_19375,N_17906,N_16397);
nand U19376 (N_19376,N_14418,N_13155);
or U19377 (N_19377,N_12519,N_13684);
nor U19378 (N_19378,N_17703,N_17278);
or U19379 (N_19379,N_15010,N_17892);
nor U19380 (N_19380,N_16599,N_18493);
and U19381 (N_19381,N_18124,N_16426);
and U19382 (N_19382,N_15438,N_17435);
or U19383 (N_19383,N_17870,N_13168);
nand U19384 (N_19384,N_17405,N_15878);
and U19385 (N_19385,N_18414,N_17236);
nor U19386 (N_19386,N_13403,N_15958);
nand U19387 (N_19387,N_15702,N_12751);
and U19388 (N_19388,N_14059,N_13514);
xnor U19389 (N_19389,N_17124,N_14952);
nand U19390 (N_19390,N_14399,N_13751);
or U19391 (N_19391,N_15644,N_15677);
nand U19392 (N_19392,N_16520,N_13197);
nor U19393 (N_19393,N_15787,N_12698);
or U19394 (N_19394,N_12578,N_18079);
nand U19395 (N_19395,N_12966,N_13800);
and U19396 (N_19396,N_16573,N_13903);
nand U19397 (N_19397,N_18588,N_15671);
nand U19398 (N_19398,N_17410,N_15089);
xnor U19399 (N_19399,N_15533,N_16017);
nand U19400 (N_19400,N_12795,N_17423);
nor U19401 (N_19401,N_17788,N_13837);
or U19402 (N_19402,N_15105,N_13913);
xor U19403 (N_19403,N_18699,N_17548);
nand U19404 (N_19404,N_18001,N_15584);
nand U19405 (N_19405,N_13058,N_15252);
nand U19406 (N_19406,N_16035,N_16020);
or U19407 (N_19407,N_12580,N_14140);
nor U19408 (N_19408,N_18180,N_14172);
nand U19409 (N_19409,N_14269,N_18418);
nand U19410 (N_19410,N_15941,N_14031);
nand U19411 (N_19411,N_15961,N_12746);
nor U19412 (N_19412,N_16311,N_16368);
nand U19413 (N_19413,N_16473,N_15560);
xnor U19414 (N_19414,N_13478,N_15369);
nor U19415 (N_19415,N_14195,N_15863);
nor U19416 (N_19416,N_14255,N_13834);
nor U19417 (N_19417,N_18250,N_12503);
or U19418 (N_19418,N_12641,N_17197);
xnor U19419 (N_19419,N_17521,N_15920);
or U19420 (N_19420,N_15218,N_15050);
xor U19421 (N_19421,N_17298,N_18138);
or U19422 (N_19422,N_14595,N_18696);
nor U19423 (N_19423,N_14440,N_17002);
xnor U19424 (N_19424,N_18748,N_15303);
nor U19425 (N_19425,N_15531,N_14760);
and U19426 (N_19426,N_17802,N_16047);
nand U19427 (N_19427,N_16884,N_15955);
nand U19428 (N_19428,N_12611,N_14972);
nor U19429 (N_19429,N_14812,N_16239);
xnor U19430 (N_19430,N_13952,N_13841);
nand U19431 (N_19431,N_14559,N_15305);
or U19432 (N_19432,N_16886,N_18222);
xnor U19433 (N_19433,N_18119,N_17406);
xnor U19434 (N_19434,N_17602,N_16651);
and U19435 (N_19435,N_17171,N_17688);
nor U19436 (N_19436,N_14631,N_13606);
or U19437 (N_19437,N_15362,N_15116);
nor U19438 (N_19438,N_16655,N_12667);
nand U19439 (N_19439,N_15683,N_16286);
and U19440 (N_19440,N_18521,N_14902);
xor U19441 (N_19441,N_18350,N_18102);
xnor U19442 (N_19442,N_17865,N_15850);
nand U19443 (N_19443,N_13626,N_14208);
or U19444 (N_19444,N_12714,N_12674);
or U19445 (N_19445,N_14978,N_16408);
nand U19446 (N_19446,N_18671,N_15911);
and U19447 (N_19447,N_18619,N_14926);
nand U19448 (N_19448,N_17349,N_13165);
or U19449 (N_19449,N_16819,N_17924);
xnor U19450 (N_19450,N_16777,N_14351);
and U19451 (N_19451,N_14295,N_15857);
or U19452 (N_19452,N_12949,N_16477);
nand U19453 (N_19453,N_13912,N_15606);
nand U19454 (N_19454,N_15247,N_12569);
xor U19455 (N_19455,N_12981,N_14433);
nor U19456 (N_19456,N_16897,N_15335);
xor U19457 (N_19457,N_16530,N_17706);
nor U19458 (N_19458,N_13526,N_14449);
and U19459 (N_19459,N_17927,N_14353);
or U19460 (N_19460,N_14862,N_17304);
xnor U19461 (N_19461,N_18437,N_17041);
xnor U19462 (N_19462,N_14801,N_16532);
and U19463 (N_19463,N_13964,N_13026);
nor U19464 (N_19464,N_16768,N_17702);
or U19465 (N_19465,N_18100,N_13783);
nand U19466 (N_19466,N_17234,N_15212);
or U19467 (N_19467,N_17576,N_15663);
nor U19468 (N_19468,N_13412,N_18577);
nor U19469 (N_19469,N_14830,N_17020);
or U19470 (N_19470,N_14503,N_15615);
and U19471 (N_19471,N_12504,N_15507);
xnor U19472 (N_19472,N_15061,N_14080);
and U19473 (N_19473,N_13297,N_15640);
and U19474 (N_19474,N_18419,N_14908);
and U19475 (N_19475,N_18198,N_12786);
nor U19476 (N_19476,N_16037,N_16781);
or U19477 (N_19477,N_16319,N_17594);
nor U19478 (N_19478,N_17750,N_14277);
nor U19479 (N_19479,N_15487,N_12646);
nor U19480 (N_19480,N_17556,N_13748);
nand U19481 (N_19481,N_15200,N_13820);
nand U19482 (N_19482,N_16401,N_13852);
or U19483 (N_19483,N_14724,N_13138);
or U19484 (N_19484,N_17110,N_13737);
nor U19485 (N_19485,N_17338,N_14469);
nand U19486 (N_19486,N_15080,N_13315);
or U19487 (N_19487,N_16040,N_15379);
xnor U19488 (N_19488,N_12794,N_13396);
xnor U19489 (N_19489,N_14304,N_14773);
xnor U19490 (N_19490,N_16182,N_17492);
or U19491 (N_19491,N_16690,N_16587);
and U19492 (N_19492,N_13289,N_14875);
xor U19493 (N_19493,N_13900,N_15688);
xnor U19494 (N_19494,N_18708,N_14510);
or U19495 (N_19495,N_13690,N_18066);
or U19496 (N_19496,N_16947,N_12650);
xnor U19497 (N_19497,N_13962,N_14198);
xor U19498 (N_19498,N_13007,N_15741);
and U19499 (N_19499,N_15214,N_18494);
xnor U19500 (N_19500,N_13650,N_17611);
xnor U19501 (N_19501,N_14142,N_13079);
nor U19502 (N_19502,N_13293,N_18382);
xor U19503 (N_19503,N_15926,N_18527);
xnor U19504 (N_19504,N_17968,N_18308);
xor U19505 (N_19505,N_13666,N_14285);
xor U19506 (N_19506,N_15611,N_16780);
and U19507 (N_19507,N_17944,N_13499);
xnor U19508 (N_19508,N_13305,N_14034);
and U19509 (N_19509,N_13450,N_13268);
or U19510 (N_19510,N_17463,N_15258);
nand U19511 (N_19511,N_18302,N_15547);
nand U19512 (N_19512,N_16550,N_18115);
nand U19513 (N_19513,N_12930,N_14491);
nor U19514 (N_19514,N_15143,N_15758);
xor U19515 (N_19515,N_14364,N_17230);
nor U19516 (N_19516,N_15183,N_18636);
xnor U19517 (N_19517,N_18405,N_12685);
or U19518 (N_19518,N_16536,N_12818);
or U19519 (N_19519,N_12820,N_18131);
and U19520 (N_19520,N_15739,N_13588);
or U19521 (N_19521,N_15012,N_14594);
nand U19522 (N_19522,N_17920,N_15998);
or U19523 (N_19523,N_14495,N_16434);
xor U19524 (N_19524,N_17592,N_15149);
and U19525 (N_19525,N_12918,N_13697);
or U19526 (N_19526,N_15555,N_14254);
or U19527 (N_19527,N_15833,N_17284);
and U19528 (N_19528,N_15967,N_15568);
and U19529 (N_19529,N_16921,N_16023);
and U19530 (N_19530,N_16164,N_14979);
and U19531 (N_19531,N_16840,N_14250);
and U19532 (N_19532,N_16345,N_13581);
nand U19533 (N_19533,N_17957,N_15024);
xnor U19534 (N_19534,N_16954,N_16999);
nor U19535 (N_19535,N_15468,N_16848);
nand U19536 (N_19536,N_13633,N_16979);
or U19537 (N_19537,N_13039,N_16880);
nand U19538 (N_19538,N_16254,N_12733);
or U19539 (N_19539,N_14709,N_17884);
nand U19540 (N_19540,N_15128,N_13535);
and U19541 (N_19541,N_17422,N_14644);
or U19542 (N_19542,N_17828,N_18415);
nor U19543 (N_19543,N_14262,N_14049);
and U19544 (N_19544,N_17245,N_13151);
nor U19545 (N_19545,N_15599,N_14354);
and U19546 (N_19546,N_15162,N_13786);
nand U19547 (N_19547,N_13542,N_13951);
nor U19548 (N_19548,N_14061,N_15471);
and U19549 (N_19549,N_13097,N_18249);
nand U19550 (N_19550,N_13889,N_14824);
nor U19551 (N_19551,N_12541,N_17247);
nand U19552 (N_19552,N_13975,N_18400);
nand U19553 (N_19553,N_18282,N_14664);
xor U19554 (N_19554,N_16740,N_16795);
and U19555 (N_19555,N_16682,N_18397);
nor U19556 (N_19556,N_13658,N_15339);
nand U19557 (N_19557,N_14993,N_15652);
or U19558 (N_19558,N_14320,N_17118);
nor U19559 (N_19559,N_15795,N_14786);
or U19560 (N_19560,N_13393,N_12659);
xnor U19561 (N_19561,N_14504,N_18208);
nor U19562 (N_19562,N_15124,N_17939);
or U19563 (N_19563,N_12649,N_13692);
nand U19564 (N_19564,N_14789,N_15986);
nand U19565 (N_19565,N_13267,N_16487);
or U19566 (N_19566,N_13850,N_16297);
xor U19567 (N_19567,N_17774,N_13255);
nand U19568 (N_19568,N_16441,N_18725);
and U19569 (N_19569,N_16277,N_18035);
nor U19570 (N_19570,N_14370,N_17265);
or U19571 (N_19571,N_17164,N_16135);
nor U19572 (N_19572,N_18399,N_18670);
nor U19573 (N_19573,N_14928,N_14465);
nor U19574 (N_19574,N_13205,N_18007);
and U19575 (N_19575,N_16029,N_16295);
or U19576 (N_19576,N_16159,N_13734);
xor U19577 (N_19577,N_13463,N_16352);
nor U19578 (N_19578,N_14589,N_12618);
nor U19579 (N_19579,N_16172,N_14261);
xnor U19580 (N_19580,N_13707,N_16446);
nand U19581 (N_19581,N_16206,N_17859);
nand U19582 (N_19582,N_17042,N_14446);
nor U19583 (N_19583,N_16083,N_14959);
xnor U19584 (N_19584,N_17495,N_12736);
xnor U19585 (N_19585,N_13663,N_16683);
and U19586 (N_19586,N_13344,N_15067);
nand U19587 (N_19587,N_17779,N_13064);
nor U19588 (N_19588,N_16056,N_16098);
and U19589 (N_19589,N_14576,N_15329);
and U19590 (N_19590,N_14313,N_14476);
or U19591 (N_19591,N_16691,N_14984);
and U19592 (N_19592,N_15257,N_14339);
or U19593 (N_19593,N_17873,N_17354);
nor U19594 (N_19594,N_16911,N_15709);
nand U19595 (N_19595,N_17753,N_13227);
and U19596 (N_19596,N_15537,N_17843);
nor U19597 (N_19597,N_15805,N_15102);
and U19598 (N_19598,N_15730,N_13372);
nand U19599 (N_19599,N_12889,N_17326);
xor U19600 (N_19600,N_12574,N_16050);
or U19601 (N_19601,N_17176,N_15978);
and U19602 (N_19602,N_17952,N_12806);
xor U19603 (N_19603,N_18668,N_17916);
or U19604 (N_19604,N_18254,N_15610);
nand U19605 (N_19605,N_12525,N_13321);
nand U19606 (N_19606,N_15500,N_18698);
and U19607 (N_19607,N_16015,N_15453);
and U19608 (N_19608,N_13010,N_16058);
or U19609 (N_19609,N_12701,N_14909);
xor U19610 (N_19610,N_17882,N_16906);
nor U19611 (N_19611,N_16905,N_13750);
xnor U19612 (N_19612,N_13281,N_17449);
nand U19613 (N_19613,N_12621,N_18433);
nand U19614 (N_19614,N_14458,N_18063);
nor U19615 (N_19615,N_14209,N_18347);
or U19616 (N_19616,N_14777,N_16289);
nand U19617 (N_19617,N_14966,N_18206);
nand U19618 (N_19618,N_13456,N_14685);
or U19619 (N_19619,N_17340,N_17806);
and U19620 (N_19620,N_17848,N_15607);
or U19621 (N_19621,N_17931,N_14745);
nor U19622 (N_19622,N_16396,N_18341);
xor U19623 (N_19623,N_15099,N_17525);
and U19624 (N_19624,N_13549,N_14517);
and U19625 (N_19625,N_15261,N_13694);
or U19626 (N_19626,N_16393,N_17915);
and U19627 (N_19627,N_12690,N_13213);
and U19628 (N_19628,N_17360,N_13066);
nor U19629 (N_19629,N_16173,N_13212);
nor U19630 (N_19630,N_13332,N_15342);
or U19631 (N_19631,N_17559,N_18238);
xnor U19632 (N_19632,N_14394,N_15060);
or U19633 (N_19633,N_15229,N_17684);
nor U19634 (N_19634,N_16045,N_15284);
xnor U19635 (N_19635,N_13291,N_14842);
nand U19636 (N_19636,N_17696,N_18617);
or U19637 (N_19637,N_15596,N_18295);
nand U19638 (N_19638,N_14282,N_17461);
or U19639 (N_19639,N_14424,N_17524);
and U19640 (N_19640,N_12850,N_14893);
xnor U19641 (N_19641,N_17846,N_15081);
or U19642 (N_19642,N_17642,N_17951);
or U19643 (N_19643,N_17082,N_15355);
and U19644 (N_19644,N_12543,N_13373);
xor U19645 (N_19645,N_15030,N_14006);
and U19646 (N_19646,N_18589,N_14478);
or U19647 (N_19647,N_17519,N_16180);
and U19648 (N_19648,N_15310,N_14920);
xor U19649 (N_19649,N_14944,N_13204);
xor U19650 (N_19650,N_16792,N_16941);
xnor U19651 (N_19651,N_14977,N_13228);
xnor U19652 (N_19652,N_13661,N_13114);
or U19653 (N_19653,N_13538,N_12647);
and U19654 (N_19654,N_18648,N_13042);
nand U19655 (N_19655,N_13260,N_16945);
and U19656 (N_19656,N_14762,N_15423);
or U19657 (N_19657,N_15020,N_16699);
and U19658 (N_19658,N_17312,N_18372);
or U19659 (N_19659,N_12662,N_17083);
or U19660 (N_19660,N_13337,N_17036);
nand U19661 (N_19661,N_16708,N_16068);
xnor U19662 (N_19662,N_14223,N_15797);
nor U19663 (N_19663,N_13735,N_13993);
or U19664 (N_19664,N_16816,N_14562);
nand U19665 (N_19665,N_15400,N_17275);
and U19666 (N_19666,N_15201,N_17844);
or U19667 (N_19667,N_14860,N_13002);
and U19668 (N_19668,N_17685,N_16844);
or U19669 (N_19669,N_17054,N_12968);
nor U19670 (N_19670,N_17372,N_15378);
or U19671 (N_19671,N_18247,N_13672);
and U19672 (N_19672,N_16244,N_18098);
xor U19673 (N_19673,N_17381,N_16637);
xnor U19674 (N_19674,N_14592,N_14229);
or U19675 (N_19675,N_13961,N_17339);
xnor U19676 (N_19676,N_14749,N_13179);
nand U19677 (N_19677,N_13200,N_17129);
and U19678 (N_19678,N_15324,N_14757);
and U19679 (N_19679,N_15301,N_17946);
nor U19680 (N_19680,N_13988,N_13652);
and U19681 (N_19681,N_16369,N_15232);
xnor U19682 (N_19682,N_16950,N_17385);
nor U19683 (N_19683,N_16992,N_16016);
xor U19684 (N_19684,N_15386,N_13801);
and U19685 (N_19685,N_12520,N_12577);
nor U19686 (N_19686,N_13842,N_14022);
nand U19687 (N_19687,N_13726,N_15090);
and U19688 (N_19688,N_16470,N_12660);
and U19689 (N_19689,N_15494,N_15441);
nor U19690 (N_19690,N_13353,N_15202);
nor U19691 (N_19691,N_12552,N_18701);
or U19692 (N_19692,N_13909,N_17334);
nor U19693 (N_19693,N_16727,N_14057);
nand U19694 (N_19694,N_16729,N_14822);
or U19695 (N_19695,N_14716,N_12729);
and U19696 (N_19696,N_17229,N_17862);
xor U19697 (N_19697,N_16866,N_16074);
nand U19698 (N_19698,N_14431,N_16367);
nor U19699 (N_19699,N_18236,N_17149);
nor U19700 (N_19700,N_15341,N_18380);
nand U19701 (N_19701,N_14454,N_13081);
nor U19702 (N_19702,N_14382,N_13120);
nand U19703 (N_19703,N_12567,N_14938);
nand U19704 (N_19704,N_12816,N_14098);
nand U19705 (N_19705,N_13890,N_14260);
xor U19706 (N_19706,N_14501,N_16842);
nor U19707 (N_19707,N_16221,N_12610);
nor U19708 (N_19708,N_18174,N_17598);
xor U19709 (N_19709,N_16502,N_12894);
nor U19710 (N_19710,N_18287,N_14932);
nand U19711 (N_19711,N_15150,N_17762);
nor U19712 (N_19712,N_15476,N_17943);
or U19713 (N_19713,N_13035,N_14081);
or U19714 (N_19714,N_13173,N_14618);
xor U19715 (N_19715,N_18223,N_18020);
nand U19716 (N_19716,N_18203,N_14768);
or U19717 (N_19717,N_14990,N_18227);
and U19718 (N_19718,N_14419,N_14911);
xor U19719 (N_19719,N_13198,N_18724);
nand U19720 (N_19720,N_16714,N_13911);
or U19721 (N_19721,N_17085,N_18262);
nor U19722 (N_19722,N_13144,N_16245);
or U19723 (N_19723,N_13343,N_13515);
and U19724 (N_19724,N_14017,N_14225);
or U19725 (N_19725,N_17934,N_13631);
nor U19726 (N_19726,N_17593,N_17331);
nor U19727 (N_19727,N_13338,N_16813);
or U19728 (N_19728,N_16977,N_16413);
or U19729 (N_19729,N_16863,N_16728);
nand U19730 (N_19730,N_14251,N_13318);
or U19731 (N_19731,N_13550,N_13923);
nor U19732 (N_19732,N_14112,N_15459);
nor U19733 (N_19733,N_17061,N_15120);
nand U19734 (N_19734,N_15082,N_17746);
or U19735 (N_19735,N_15848,N_12952);
xnor U19736 (N_19736,N_15871,N_18732);
nand U19737 (N_19737,N_13399,N_13217);
xor U19738 (N_19738,N_14332,N_18492);
nor U19739 (N_19739,N_17803,N_16385);
nand U19740 (N_19740,N_13872,N_18510);
xor U19741 (N_19741,N_15984,N_13888);
or U19742 (N_19742,N_14464,N_16871);
or U19743 (N_19743,N_13854,N_13771);
and U19744 (N_19744,N_17841,N_17297);
or U19745 (N_19745,N_16634,N_17370);
nand U19746 (N_19746,N_16304,N_12691);
and U19747 (N_19747,N_15841,N_14661);
nor U19748 (N_19748,N_14502,N_18673);
and U19749 (N_19749,N_15852,N_13636);
xnor U19750 (N_19750,N_15396,N_15921);
or U19751 (N_19751,N_14186,N_16374);
xor U19752 (N_19752,N_16494,N_14635);
nand U19753 (N_19753,N_13417,N_18316);
xor U19754 (N_19754,N_17694,N_18622);
and U19755 (N_19755,N_18147,N_14460);
or U19756 (N_19756,N_13452,N_16204);
nand U19757 (N_19757,N_17494,N_15293);
xnor U19758 (N_19758,N_16888,N_17172);
nand U19759 (N_19759,N_12735,N_18195);
or U19760 (N_19760,N_17088,N_16002);
nor U19761 (N_19761,N_16998,N_13350);
nand U19762 (N_19762,N_18470,N_14740);
nor U19763 (N_19763,N_13178,N_16410);
or U19764 (N_19764,N_14127,N_15152);
or U19765 (N_19765,N_16332,N_16008);
and U19766 (N_19766,N_13791,N_17015);
nand U19767 (N_19767,N_14153,N_17748);
xor U19768 (N_19768,N_15664,N_15349);
and U19769 (N_19769,N_14945,N_16234);
and U19770 (N_19770,N_17737,N_13237);
and U19771 (N_19771,N_14511,N_17948);
and U19772 (N_19772,N_14624,N_15452);
or U19773 (N_19773,N_14256,N_14953);
nor U19774 (N_19774,N_12900,N_17321);
and U19775 (N_19775,N_16971,N_18549);
nor U19776 (N_19776,N_17650,N_17132);
xnor U19777 (N_19777,N_15073,N_15800);
xor U19778 (N_19778,N_16174,N_15569);
and U19779 (N_19779,N_16111,N_16305);
and U19780 (N_19780,N_18463,N_16915);
xnor U19781 (N_19781,N_13843,N_17899);
or U19782 (N_19782,N_13918,N_12832);
nand U19783 (N_19783,N_13325,N_15856);
nor U19784 (N_19784,N_15273,N_14406);
or U19785 (N_19785,N_15207,N_16949);
nand U19786 (N_19786,N_14855,N_14714);
or U19787 (N_19787,N_18054,N_16064);
or U19788 (N_19788,N_16125,N_16496);
xor U19789 (N_19789,N_12681,N_17735);
and U19790 (N_19790,N_16876,N_16442);
nor U19791 (N_19791,N_17139,N_15274);
nand U19792 (N_19792,N_12992,N_17395);
and U19793 (N_19793,N_18317,N_12815);
nand U19794 (N_19794,N_17249,N_12925);
and U19795 (N_19795,N_14516,N_16123);
or U19796 (N_19796,N_14693,N_12856);
nand U19797 (N_19797,N_16666,N_16031);
nand U19798 (N_19798,N_16072,N_14701);
xor U19799 (N_19799,N_15352,N_17584);
and U19800 (N_19800,N_18557,N_15905);
and U19801 (N_19801,N_13669,N_12759);
nand U19802 (N_19802,N_18570,N_14227);
or U19803 (N_19803,N_15309,N_15170);
and U19804 (N_19804,N_12640,N_14580);
xor U19805 (N_19805,N_17274,N_13853);
nor U19806 (N_19806,N_15424,N_18273);
and U19807 (N_19807,N_16746,N_17306);
nand U19808 (N_19808,N_13811,N_17628);
or U19809 (N_19809,N_18721,N_18439);
nor U19810 (N_19810,N_14408,N_12780);
or U19811 (N_19811,N_14539,N_17804);
or U19812 (N_19812,N_17404,N_14041);
or U19813 (N_19813,N_16412,N_17231);
nor U19814 (N_19814,N_18685,N_15880);
xnor U19815 (N_19815,N_16831,N_16350);
nand U19816 (N_19816,N_17937,N_12822);
and U19817 (N_19817,N_14607,N_12534);
nor U19818 (N_19818,N_18046,N_17600);
and U19819 (N_19819,N_14717,N_17024);
nor U19820 (N_19820,N_13304,N_14447);
xor U19821 (N_19821,N_18120,N_14599);
or U19822 (N_19822,N_13784,N_14610);
nand U19823 (N_19823,N_18716,N_14438);
xnor U19824 (N_19824,N_14188,N_15179);
xor U19825 (N_19825,N_15323,N_16336);
xor U19826 (N_19826,N_13147,N_14547);
nor U19827 (N_19827,N_13616,N_16662);
xor U19828 (N_19828,N_18583,N_13294);
xor U19829 (N_19829,N_16733,N_15343);
or U19830 (N_19830,N_16448,N_16237);
nor U19831 (N_19831,N_16317,N_14011);
nor U19832 (N_19832,N_13188,N_16331);
nand U19833 (N_19833,N_12807,N_15557);
xor U19834 (N_19834,N_14169,N_14253);
nor U19835 (N_19835,N_12897,N_18678);
xor U19836 (N_19836,N_18421,N_17914);
xor U19837 (N_19837,N_17571,N_18094);
and U19838 (N_19838,N_15743,N_15881);
nor U19839 (N_19839,N_12796,N_16519);
or U19840 (N_19840,N_17309,N_14955);
xnor U19841 (N_19841,N_17724,N_12915);
nand U19842 (N_19842,N_18323,N_17496);
nor U19843 (N_19843,N_15813,N_16003);
nor U19844 (N_19844,N_16136,N_16259);
nand U19845 (N_19845,N_18722,N_16955);
nor U19846 (N_19846,N_16379,N_17003);
and U19847 (N_19847,N_18425,N_17469);
nor U19848 (N_19848,N_16112,N_14004);
nor U19849 (N_19849,N_13857,N_16409);
nand U19850 (N_19850,N_13600,N_12997);
nor U19851 (N_19851,N_13738,N_15108);
nand U19852 (N_19852,N_14715,N_15422);
or U19853 (N_19853,N_18445,N_15353);
nand U19854 (N_19854,N_13638,N_17969);
xnor U19855 (N_19855,N_14793,N_12629);
and U19856 (N_19856,N_15895,N_13895);
xor U19857 (N_19857,N_17305,N_14236);
and U19858 (N_19858,N_13109,N_14744);
and U19859 (N_19859,N_12948,N_13686);
nor U19860 (N_19860,N_18186,N_14639);
or U19861 (N_19861,N_14050,N_17064);
or U19862 (N_19862,N_12664,N_14300);
or U19863 (N_19863,N_14838,N_18398);
or U19864 (N_19864,N_18345,N_16735);
xnor U19865 (N_19865,N_13944,N_13070);
nor U19866 (N_19866,N_15125,N_18344);
nor U19867 (N_19867,N_15902,N_13766);
and U19868 (N_19868,N_13714,N_15306);
nor U19869 (N_19869,N_15347,N_17133);
xnor U19870 (N_19870,N_13376,N_15263);
nand U19871 (N_19871,N_13630,N_16384);
nor U19872 (N_19872,N_18135,N_17978);
xnor U19873 (N_19873,N_14205,N_16865);
nor U19874 (N_19874,N_14949,N_14907);
nand U19875 (N_19875,N_16817,N_12718);
nor U19876 (N_19876,N_15477,N_17636);
nor U19877 (N_19877,N_13252,N_13769);
nand U19878 (N_19878,N_13601,N_14210);
or U19879 (N_19879,N_15657,N_16524);
nand U19880 (N_19880,N_17113,N_16983);
or U19881 (N_19881,N_15109,N_18166);
nor U19882 (N_19882,N_16712,N_14124);
xor U19883 (N_19883,N_13891,N_18590);
nand U19884 (N_19884,N_18239,N_14804);
nor U19885 (N_19885,N_18016,N_15275);
nor U19886 (N_19886,N_14147,N_18504);
nor U19887 (N_19887,N_16133,N_13706);
nand U19888 (N_19888,N_16501,N_14871);
nand U19889 (N_19889,N_13016,N_12825);
nor U19890 (N_19890,N_16445,N_15551);
or U19891 (N_19891,N_12962,N_17380);
or U19892 (N_19892,N_14160,N_16404);
or U19893 (N_19893,N_14358,N_17464);
nor U19894 (N_19894,N_17604,N_15931);
nand U19895 (N_19895,N_17823,N_15484);
xnor U19896 (N_19896,N_12529,N_12986);
or U19897 (N_19897,N_18311,N_14750);
and U19898 (N_19898,N_16570,N_14016);
or U19899 (N_19899,N_17877,N_14841);
nand U19900 (N_19900,N_14613,N_18086);
nor U19901 (N_19901,N_18358,N_12596);
and U19902 (N_19902,N_13037,N_13336);
nand U19903 (N_19903,N_15704,N_17476);
nor U19904 (N_19904,N_15175,N_12819);
xnor U19905 (N_19905,N_17560,N_18365);
xnor U19906 (N_19906,N_14301,N_13390);
nand U19907 (N_19907,N_13386,N_18005);
nor U19908 (N_19908,N_12979,N_15177);
nor U19909 (N_19909,N_12732,N_14654);
nor U19910 (N_19910,N_15968,N_14244);
nor U19911 (N_19911,N_18420,N_14847);
or U19912 (N_19912,N_14802,N_12717);
xnor U19913 (N_19913,N_14245,N_18301);
xnor U19914 (N_19914,N_15278,N_15135);
and U19915 (N_19915,N_12686,N_14481);
nand U19916 (N_19916,N_16694,N_14958);
or U19917 (N_19917,N_15914,N_16324);
nor U19918 (N_19918,N_13324,N_18597);
nor U19919 (N_19919,N_15948,N_17655);
or U19920 (N_19920,N_15873,N_18628);
xor U19921 (N_19921,N_14143,N_14779);
and U19922 (N_19922,N_14104,N_12597);
nand U19923 (N_19923,N_17076,N_15101);
nor U19924 (N_19924,N_16088,N_14107);
nor U19925 (N_19925,N_17159,N_13585);
and U19926 (N_19926,N_14946,N_16217);
and U19927 (N_19927,N_14303,N_17514);
xor U19928 (N_19928,N_13469,N_12707);
nor U19929 (N_19929,N_15033,N_16402);
nor U19930 (N_19930,N_15417,N_15270);
nand U19931 (N_19931,N_17500,N_13908);
and U19932 (N_19932,N_16283,N_17281);
or U19933 (N_19933,N_12769,N_13794);
and U19934 (N_19934,N_12788,N_12936);
or U19935 (N_19935,N_14386,N_16901);
nand U19936 (N_19936,N_17861,N_13011);
or U19937 (N_19937,N_18538,N_12866);
nand U19938 (N_19938,N_16879,N_18275);
nor U19939 (N_19939,N_15406,N_18190);
xor U19940 (N_19940,N_17935,N_17659);
nand U19941 (N_19941,N_17365,N_15549);
or U19942 (N_19942,N_16422,N_16760);
nand U19943 (N_19943,N_14015,N_17991);
nand U19944 (N_19944,N_12776,N_18148);
or U19945 (N_19945,N_16344,N_13728);
nand U19946 (N_19946,N_12941,N_17790);
or U19947 (N_19947,N_14404,N_18475);
nor U19948 (N_19948,N_15844,N_16452);
nand U19949 (N_19949,N_17456,N_15798);
xor U19950 (N_19950,N_13261,N_15285);
nand U19951 (N_19951,N_15992,N_15972);
and U19952 (N_19952,N_16415,N_12711);
and U19953 (N_19953,N_15985,N_18403);
xnor U19954 (N_19954,N_13824,N_16734);
xnor U19955 (N_19955,N_15192,N_15697);
or U19956 (N_19956,N_14043,N_12639);
nand U19957 (N_19957,N_16340,N_13696);
or U19958 (N_19958,N_17201,N_12838);
nor U19959 (N_19959,N_18719,N_13742);
or U19960 (N_19960,N_17134,N_18213);
xnor U19961 (N_19961,N_14324,N_15876);
and U19962 (N_19962,N_15508,N_18669);
nand U19963 (N_19963,N_14761,N_12539);
nor U19964 (N_19964,N_15567,N_15897);
and U19965 (N_19965,N_16236,N_13744);
and U19966 (N_19966,N_14718,N_15842);
nor U19967 (N_19967,N_17639,N_12766);
and U19968 (N_19968,N_15336,N_16556);
and U19969 (N_19969,N_13527,N_15818);
or U19970 (N_19970,N_18401,N_13159);
xor U19971 (N_19971,N_15357,N_12619);
and U19972 (N_19972,N_13713,N_16624);
nand U19973 (N_19973,N_17660,N_13308);
or U19974 (N_19974,N_17403,N_12624);
xnor U19975 (N_19975,N_18253,N_13194);
or U19976 (N_19976,N_16260,N_17522);
xor U19977 (N_19977,N_18656,N_16788);
and U19978 (N_19978,N_14189,N_16970);
and U19979 (N_19979,N_15843,N_16669);
and U19980 (N_19980,N_18178,N_17743);
and U19981 (N_19981,N_16461,N_15949);
xnor U19982 (N_19982,N_13525,N_16137);
nor U19983 (N_19983,N_18021,N_12919);
and U19984 (N_19984,N_15892,N_14119);
or U19985 (N_19985,N_13528,N_12715);
nor U19986 (N_19986,N_17239,N_15966);
nand U19987 (N_19987,N_15382,N_18551);
and U19988 (N_19988,N_15632,N_17677);
nor U19989 (N_19989,N_13674,N_18117);
and U19990 (N_19990,N_12865,N_17501);
or U19991 (N_19991,N_14852,N_15361);
nand U19992 (N_19992,N_16103,N_12679);
or U19993 (N_19993,N_18743,N_17983);
nand U19994 (N_19994,N_13545,N_12955);
nand U19995 (N_19995,N_15115,N_15407);
xor U19996 (N_19996,N_15295,N_16211);
xnor U19997 (N_19997,N_13431,N_18070);
nor U19998 (N_19998,N_13520,N_15828);
or U19999 (N_19999,N_16892,N_18199);
and U20000 (N_20000,N_14922,N_16252);
or U20001 (N_20001,N_16085,N_18607);
xor U20002 (N_20002,N_13459,N_13101);
xnor U20003 (N_20003,N_14667,N_15245);
and U20004 (N_20004,N_14070,N_18498);
or U20005 (N_20005,N_13423,N_14411);
xnor U20006 (N_20006,N_15501,N_14434);
and U20007 (N_20007,N_16942,N_13699);
or U20008 (N_20008,N_13209,N_15806);
xor U20009 (N_20009,N_17027,N_16145);
nand U20010 (N_20010,N_13307,N_13507);
or U20011 (N_20011,N_15934,N_12689);
xnor U20012 (N_20012,N_14028,N_14321);
xor U20013 (N_20013,N_14166,N_13383);
xnor U20014 (N_20014,N_14763,N_16636);
xnor U20015 (N_20015,N_16881,N_15093);
nand U20016 (N_20016,N_17502,N_16713);
or U20017 (N_20017,N_12988,N_14231);
nand U20018 (N_20018,N_13556,N_17974);
nand U20019 (N_20019,N_14352,N_14274);
nor U20020 (N_20020,N_15235,N_15014);
and U20021 (N_20021,N_14365,N_16216);
or U20022 (N_20022,N_15621,N_13415);
xnor U20023 (N_20023,N_15144,N_14936);
nand U20024 (N_20024,N_18737,N_15374);
and U20025 (N_20025,N_18720,N_16629);
or U20026 (N_20026,N_16925,N_16063);
or U20027 (N_20027,N_17618,N_13446);
nand U20028 (N_20028,N_15904,N_16723);
or U20029 (N_20029,N_12565,N_13497);
and U20030 (N_20030,N_17985,N_13761);
and U20031 (N_20031,N_14741,N_18043);
nand U20032 (N_20032,N_12694,N_14947);
xor U20033 (N_20033,N_14492,N_15100);
and U20034 (N_20034,N_18099,N_16500);
xnor U20035 (N_20035,N_16642,N_13182);
nand U20036 (N_20036,N_12752,N_13505);
or U20037 (N_20037,N_17999,N_13777);
nor U20038 (N_20038,N_16545,N_13330);
or U20039 (N_20039,N_16273,N_18128);
nor U20040 (N_20040,N_17189,N_15589);
nor U20041 (N_20041,N_15587,N_15879);
or U20042 (N_20042,N_14751,N_14123);
xnor U20043 (N_20043,N_18259,N_18417);
or U20044 (N_20044,N_13191,N_18441);
xnor U20045 (N_20045,N_12933,N_12920);
and U20046 (N_20046,N_13451,N_17925);
xnor U20047 (N_20047,N_14316,N_14605);
or U20048 (N_20048,N_18332,N_17026);
or U20049 (N_20049,N_14957,N_18655);
nor U20050 (N_20050,N_15861,N_16687);
or U20051 (N_20051,N_17990,N_14474);
nand U20052 (N_20052,N_16554,N_12804);
nor U20053 (N_20053,N_13807,N_13286);
and U20054 (N_20054,N_17211,N_14233);
and U20055 (N_20055,N_16986,N_17112);
and U20056 (N_20056,N_12887,N_14273);
nand U20057 (N_20057,N_14158,N_18714);
xor U20058 (N_20058,N_17713,N_15791);
or U20059 (N_20059,N_14593,N_16338);
nand U20060 (N_20060,N_14662,N_16158);
nand U20061 (N_20061,N_13851,N_17267);
nand U20062 (N_20062,N_15465,N_13096);
nor U20063 (N_20063,N_18225,N_16152);
nand U20064 (N_20064,N_14868,N_12741);
xnor U20065 (N_20065,N_12871,N_12798);
nand U20066 (N_20066,N_14669,N_13183);
xor U20067 (N_20067,N_16222,N_16143);
nand U20068 (N_20068,N_12595,N_15648);
or U20069 (N_20069,N_12892,N_17256);
nand U20070 (N_20070,N_16571,N_16370);
nand U20071 (N_20071,N_17077,N_13945);
xor U20072 (N_20072,N_15035,N_13333);
nor U20073 (N_20073,N_16889,N_18153);
or U20074 (N_20074,N_13320,N_14389);
or U20075 (N_20075,N_13470,N_12942);
nor U20076 (N_20076,N_15793,N_17440);
xnor U20077 (N_20077,N_17126,N_16852);
or U20078 (N_20078,N_15616,N_16117);
nor U20079 (N_20079,N_14451,N_14910);
nor U20080 (N_20080,N_16742,N_15762);
and U20081 (N_20081,N_12904,N_13225);
and U20082 (N_20082,N_18285,N_16553);
or U20083 (N_20083,N_17056,N_13275);
or U20084 (N_20084,N_13774,N_13421);
or U20085 (N_20085,N_13919,N_14400);
xnor U20086 (N_20086,N_13104,N_17188);
nor U20087 (N_20087,N_16188,N_13544);
nand U20088 (N_20088,N_14363,N_14294);
nand U20089 (N_20089,N_14331,N_15858);
or U20090 (N_20090,N_14267,N_13795);
nor U20091 (N_20091,N_14171,N_15825);
xor U20092 (N_20092,N_18368,N_13958);
xor U20093 (N_20093,N_18637,N_14866);
nand U20094 (N_20094,N_18134,N_13715);
or U20095 (N_20095,N_13537,N_17972);
and U20096 (N_20096,N_16957,N_16598);
nand U20097 (N_20097,N_13448,N_17885);
xnor U20098 (N_20098,N_17314,N_18495);
nand U20099 (N_20099,N_13219,N_16890);
nor U20100 (N_20100,N_15037,N_16481);
or U20101 (N_20101,N_13387,N_13782);
xor U20102 (N_20102,N_14774,N_17317);
nand U20103 (N_20103,N_18624,N_15370);
nand U20104 (N_20104,N_13967,N_17411);
and U20105 (N_20105,N_16271,N_13239);
nor U20106 (N_20106,N_18734,N_17783);
nor U20107 (N_20107,N_15312,N_15331);
nand U20108 (N_20108,N_14663,N_17072);
and U20109 (N_20109,N_17936,N_12993);
xor U20110 (N_20110,N_13517,N_13778);
xnor U20111 (N_20111,N_15117,N_15794);
or U20112 (N_20112,N_16615,N_15479);
xnor U20113 (N_20113,N_14738,N_15268);
and U20114 (N_20114,N_16383,N_13604);
or U20115 (N_20115,N_16226,N_12747);
nand U20116 (N_20116,N_14187,N_16179);
nor U20117 (N_20117,N_13171,N_18315);
nand U20118 (N_20118,N_15320,N_15638);
or U20119 (N_20119,N_14571,N_15317);
xnor U20120 (N_20120,N_13996,N_18713);
nor U20121 (N_20121,N_14062,N_17772);
or U20122 (N_20122,N_15395,N_16783);
or U20123 (N_20123,N_18013,N_15346);
and U20124 (N_20124,N_15199,N_14791);
and U20125 (N_20125,N_18212,N_12878);
nor U20126 (N_20126,N_16318,N_15077);
and U20127 (N_20127,N_14587,N_15656);
nor U20128 (N_20128,N_17550,N_15227);
nor U20129 (N_20129,N_18558,N_17651);
or U20130 (N_20130,N_18728,N_12811);
nor U20131 (N_20131,N_15474,N_14448);
and U20132 (N_20132,N_13524,N_13086);
xnor U20133 (N_20133,N_15472,N_13426);
and U20134 (N_20134,N_14925,N_13641);
nand U20135 (N_20135,N_17254,N_17216);
or U20136 (N_20136,N_17292,N_17227);
or U20137 (N_20137,N_13128,N_14217);
or U20138 (N_20138,N_15203,N_12772);
and U20139 (N_20139,N_18690,N_14180);
nand U20140 (N_20140,N_13004,N_14499);
or U20141 (N_20141,N_18364,N_16631);
and U20142 (N_20142,N_15191,N_18006);
nand U20143 (N_20143,N_17852,N_16716);
and U20144 (N_20144,N_18680,N_18572);
and U20145 (N_20145,N_16706,N_16874);
and U20146 (N_20146,N_16680,N_17021);
and U20147 (N_20147,N_18072,N_15502);
xor U20148 (N_20148,N_15188,N_18501);
nand U20149 (N_20149,N_12675,N_14398);
nand U20150 (N_20150,N_15605,N_16943);
nor U20151 (N_20151,N_18052,N_16837);
and U20152 (N_20152,N_14901,N_15694);
or U20153 (N_20153,N_13075,N_17479);
nand U20154 (N_20154,N_16018,N_14657);
and U20155 (N_20155,N_12757,N_17711);
or U20156 (N_20156,N_15716,N_15259);
and U20157 (N_20157,N_18201,N_15906);
nand U20158 (N_20158,N_13576,N_16860);
and U20159 (N_20159,N_15721,N_13763);
xnor U20160 (N_20160,N_17263,N_17055);
nor U20161 (N_20161,N_14541,N_18032);
nor U20162 (N_20162,N_17313,N_18359);
nand U20163 (N_20163,N_12668,N_13513);
xor U20164 (N_20164,N_13132,N_12563);
and U20165 (N_20165,N_15527,N_16975);
nand U20166 (N_20166,N_17537,N_16349);
nor U20167 (N_20167,N_14695,N_16207);
or U20168 (N_20168,N_17723,N_17903);
and U20169 (N_20169,N_13965,N_16150);
and U20170 (N_20170,N_13329,N_14347);
xor U20171 (N_20171,N_16300,N_12728);
and U20172 (N_20172,N_18210,N_15660);
xnor U20173 (N_20173,N_18313,N_17131);
xnor U20174 (N_20174,N_15458,N_16099);
nor U20175 (N_20175,N_13409,N_12761);
xor U20176 (N_20176,N_12763,N_13115);
nand U20177 (N_20177,N_17854,N_12765);
and U20178 (N_20178,N_14623,N_15266);
or U20179 (N_20179,N_16909,N_16038);
or U20180 (N_20180,N_15189,N_14239);
xor U20181 (N_20181,N_16144,N_17252);
nor U20182 (N_20182,N_17739,N_16497);
nor U20183 (N_20183,N_14995,N_15130);
and U20184 (N_20184,N_18686,N_14450);
and U20185 (N_20185,N_13342,N_18009);
or U20186 (N_20186,N_17527,N_14343);
xnor U20187 (N_20187,N_18548,N_13927);
or U20188 (N_20188,N_12533,N_13620);
and U20189 (N_20189,N_13306,N_17335);
and U20190 (N_20190,N_17610,N_14159);
or U20191 (N_20191,N_13346,N_14179);
xnor U20192 (N_20192,N_13938,N_18019);
nor U20193 (N_20193,N_18244,N_16192);
xnor U20194 (N_20194,N_16258,N_14609);
nor U20195 (N_20195,N_17741,N_16843);
nand U20196 (N_20196,N_17075,N_12600);
or U20197 (N_20197,N_17332,N_17970);
nor U20198 (N_20198,N_13186,N_16870);
or U20199 (N_20199,N_18658,N_12553);
or U20200 (N_20200,N_12781,N_16453);
xor U20201 (N_20201,N_13632,N_17825);
or U20202 (N_20202,N_15953,N_18303);
or U20203 (N_20203,N_14014,N_13052);
or U20204 (N_20204,N_13295,N_18307);
or U20205 (N_20205,N_13819,N_18172);
nand U20206 (N_20206,N_13827,N_18443);
nor U20207 (N_20207,N_16927,N_12726);
nor U20208 (N_20208,N_16315,N_17797);
xnor U20209 (N_20209,N_17530,N_18612);
nor U20210 (N_20210,N_17929,N_13998);
or U20211 (N_20211,N_14380,N_17719);
and U20212 (N_20212,N_13065,N_16320);
nor U20213 (N_20213,N_18370,N_15475);
nand U20214 (N_20214,N_17080,N_13721);
and U20215 (N_20215,N_12984,N_18192);
xnor U20216 (N_20216,N_15987,N_13877);
nor U20217 (N_20217,N_18049,N_17627);
nor U20218 (N_20218,N_15780,N_17364);
nor U20219 (N_20219,N_13467,N_18025);
nor U20220 (N_20220,N_12970,N_12803);
xor U20221 (N_20221,N_18641,N_17784);
xnor U20222 (N_20222,N_17270,N_17187);
xor U20223 (N_20223,N_17715,N_18352);
xor U20224 (N_20224,N_15594,N_17637);
or U20225 (N_20225,N_15164,N_16677);
and U20226 (N_20226,N_13957,N_12855);
nor U20227 (N_20227,N_14156,N_18065);
nor U20228 (N_20228,N_18657,N_14377);
and U20229 (N_20229,N_18055,N_12974);
or U20230 (N_20230,N_14630,N_14854);
xor U20231 (N_20231,N_15027,N_17887);
xor U20232 (N_20232,N_16824,N_14930);
and U20233 (N_20233,N_14982,N_17114);
or U20234 (N_20234,N_13862,N_17679);
and U20235 (N_20235,N_17563,N_15496);
and U20236 (N_20236,N_17733,N_14177);
xor U20237 (N_20237,N_18304,N_16200);
nor U20238 (N_20238,N_18067,N_14912);
or U20239 (N_20239,N_17428,N_17801);
or U20240 (N_20240,N_17031,N_15129);
or U20241 (N_20241,N_17663,N_15463);
xnor U20242 (N_20242,N_18478,N_13892);
nand U20243 (N_20243,N_15181,N_18575);
and U20244 (N_20244,N_12996,N_14228);
nor U20245 (N_20245,N_14601,N_14426);
or U20246 (N_20246,N_15799,N_14720);
nor U20247 (N_20247,N_16762,N_14278);
nor U20248 (N_20248,N_13986,N_15215);
xnor U20249 (N_20249,N_15057,N_14488);
or U20250 (N_20250,N_13718,N_15890);
and U20251 (N_20251,N_16069,N_12813);
or U20252 (N_20252,N_15829,N_15956);
and U20253 (N_20253,N_15414,N_14330);
nand U20254 (N_20254,N_16512,N_13394);
xnor U20255 (N_20255,N_13049,N_15289);
nor U20256 (N_20256,N_12672,N_13490);
nor U20257 (N_20257,N_16757,N_17816);
nor U20258 (N_20258,N_12678,N_16833);
nand U20259 (N_20259,N_15499,N_18000);
nand U20260 (N_20260,N_14518,N_12899);
nand U20261 (N_20261,N_12903,N_16626);
or U20262 (N_20262,N_18122,N_16951);
xnor U20263 (N_20263,N_16186,N_14659);
or U20264 (N_20264,N_13340,N_12632);
nor U20265 (N_20265,N_14279,N_14297);
and U20266 (N_20266,N_13797,N_13863);
and U20267 (N_20267,N_14191,N_14856);
xnor U20268 (N_20268,N_17033,N_14766);
and U20269 (N_20269,N_14369,N_13847);
nand U20270 (N_20270,N_14596,N_16294);
and U20271 (N_20271,N_18429,N_12961);
and U20272 (N_20272,N_13869,N_13929);
nand U20273 (N_20273,N_13540,N_15695);
xnor U20274 (N_20274,N_16057,N_12906);
or U20275 (N_20275,N_18059,N_18369);
or U20276 (N_20276,N_14884,N_15205);
and U20277 (N_20277,N_18233,N_13723);
xor U20278 (N_20278,N_16523,N_15241);
nor U20279 (N_20279,N_12867,N_15918);
xnor U20280 (N_20280,N_16611,N_17890);
xor U20281 (N_20281,N_18745,N_12879);
or U20282 (N_20282,N_16885,N_14591);
and U20283 (N_20283,N_18214,N_15246);
nor U20284 (N_20284,N_18187,N_17396);
nor U20285 (N_20285,N_14819,N_15572);
and U20286 (N_20286,N_15448,N_16084);
xor U20287 (N_20287,N_13474,N_14084);
nand U20288 (N_20288,N_17744,N_15131);
and U20289 (N_20289,N_17253,N_14748);
nor U20290 (N_20290,N_14444,N_16484);
and U20291 (N_20291,N_17675,N_15883);
or U20292 (N_20292,N_18270,N_15965);
or U20293 (N_20293,N_15279,N_13038);
nand U20294 (N_20294,N_14340,N_15107);
xnor U20295 (N_20295,N_17965,N_17850);
nand U20296 (N_20296,N_13195,N_17510);
or U20297 (N_20297,N_17053,N_18252);
nand U20298 (N_20298,N_12657,N_13098);
or U20299 (N_20299,N_17807,N_13495);
xnor U20300 (N_20300,N_13682,N_15264);
or U20301 (N_20301,N_15029,N_16296);
nor U20302 (N_20302,N_15334,N_14885);
nand U20303 (N_20303,N_12652,N_15026);
xnor U20304 (N_20304,N_17266,N_17329);
and U20305 (N_20305,N_17491,N_14550);
and U20306 (N_20306,N_15666,N_16429);
and U20307 (N_20307,N_14851,N_17722);
xor U20308 (N_20308,N_14268,N_14284);
nand U20309 (N_20309,N_17221,N_17821);
or U20310 (N_20310,N_15390,N_14616);
nand U20311 (N_20311,N_18529,N_16747);
xor U20312 (N_20312,N_12953,N_15291);
and U20313 (N_20313,N_13612,N_14425);
or U20314 (N_20314,N_13955,N_15733);
or U20315 (N_20315,N_12874,N_13082);
or U20316 (N_20316,N_14937,N_13818);
nand U20317 (N_20317,N_12869,N_16093);
xnor U20318 (N_20318,N_18744,N_13433);
nor U20319 (N_20319,N_16830,N_13789);
nor U20320 (N_20320,N_18337,N_14679);
or U20321 (N_20321,N_12743,N_13848);
xnor U20322 (N_20322,N_15158,N_17362);
xnor U20323 (N_20323,N_16269,N_18438);
nor U20324 (N_20324,N_16075,N_18105);
and U20325 (N_20325,N_18216,N_15769);
and U20326 (N_20326,N_16238,N_13442);
and U20327 (N_20327,N_18140,N_16053);
nand U20328 (N_20328,N_17127,N_12847);
or U20329 (N_20329,N_15543,N_18596);
or U20330 (N_20330,N_14184,N_14338);
xor U20331 (N_20331,N_13124,N_14175);
xnor U20332 (N_20332,N_16323,N_16737);
nor U20333 (N_20333,N_14782,N_14857);
or U20334 (N_20334,N_13249,N_17941);
xor U20335 (N_20335,N_15715,N_18586);
nor U20336 (N_20336,N_13796,N_13094);
and U20337 (N_20337,N_16938,N_17392);
or U20338 (N_20338,N_16522,N_17067);
or U20339 (N_20339,N_16730,N_12710);
and U20340 (N_20340,N_15975,N_15631);
nor U20341 (N_20341,N_17791,N_13089);
xor U20342 (N_20342,N_16922,N_14035);
and U20343 (N_20343,N_14614,N_16109);
nor U20344 (N_20344,N_13659,N_16437);
nand U20345 (N_20345,N_18277,N_17136);
xnor U20346 (N_20346,N_18499,N_17117);
xor U20347 (N_20347,N_13655,N_14833);
or U20348 (N_20348,N_12812,N_15812);
nand U20349 (N_20349,N_13788,N_14275);
xor U20350 (N_20350,N_15725,N_13263);
or U20351 (N_20351,N_13411,N_17658);
or U20352 (N_20352,N_18435,N_17125);
xnor U20353 (N_20353,N_16618,N_17257);
xnor U20354 (N_20354,N_15846,N_18450);
and U20355 (N_20355,N_16565,N_14410);
nand U20356 (N_20356,N_16407,N_16775);
xor U20357 (N_20357,N_18028,N_18107);
nand U20358 (N_20358,N_15069,N_12884);
and U20359 (N_20359,N_13565,N_16751);
or U20360 (N_20360,N_16649,N_13156);
xor U20361 (N_20361,N_16140,N_15898);
nor U20362 (N_20362,N_18546,N_18740);
nor U20363 (N_20363,N_17950,N_15491);
and U20364 (N_20364,N_16110,N_16469);
and U20365 (N_20365,N_13806,N_12676);
or U20366 (N_20366,N_15078,N_18742);
nand U20367 (N_20367,N_13592,N_18383);
nand U20368 (N_20368,N_16546,N_15754);
and U20369 (N_20369,N_15313,N_14374);
and U20370 (N_20370,N_16769,N_17106);
or U20371 (N_20371,N_16495,N_13400);
and U20372 (N_20372,N_14869,N_14723);
nand U20373 (N_20373,N_14734,N_16231);
xor U20374 (N_20374,N_14162,N_18428);
nand U20375 (N_20375,N_13380,N_17520);
nand U20376 (N_20376,N_18573,N_14005);
xor U20377 (N_20377,N_18068,N_13208);
and U20378 (N_20378,N_13615,N_17119);
nand U20379 (N_20379,N_17107,N_18554);
or U20380 (N_20380,N_12852,N_13475);
and U20381 (N_20381,N_18300,N_13355);
or U20382 (N_20382,N_13622,N_13504);
and U20383 (N_20383,N_16185,N_17490);
nor U20384 (N_20384,N_15582,N_12951);
nor U20385 (N_20385,N_17727,N_16585);
and U20386 (N_20386,N_14521,N_12537);
nor U20387 (N_20387,N_12546,N_17992);
or U20388 (N_20388,N_13483,N_12731);
nand U20389 (N_20389,N_17376,N_14312);
nor U20390 (N_20390,N_17493,N_16165);
and U20391 (N_20391,N_13454,N_12802);
nor U20392 (N_20392,N_17059,N_16087);
and U20393 (N_20393,N_17596,N_13732);
or U20394 (N_20394,N_18649,N_15969);
and U20395 (N_20395,N_13575,N_17764);
nor U20396 (N_20396,N_14327,N_15979);
xor U20397 (N_20397,N_14544,N_13688);
and U20398 (N_20398,N_12594,N_18491);
and U20399 (N_20399,N_16012,N_17667);
and U20400 (N_20400,N_13084,N_12797);
xnor U20401 (N_20401,N_14466,N_13050);
nor U20402 (N_20402,N_18738,N_14144);
nand U20403 (N_20403,N_18169,N_16763);
or U20404 (N_20404,N_12507,N_14007);
nand U20405 (N_20405,N_14514,N_17102);
xnor U20406 (N_20406,N_13300,N_15464);
nor U20407 (N_20407,N_15950,N_16908);
and U20408 (N_20408,N_14676,N_14381);
nor U20409 (N_20409,N_14042,N_14379);
or U20410 (N_20410,N_16290,N_17453);
nand U20411 (N_20411,N_15009,N_17529);
xnor U20412 (N_20412,N_15368,N_17868);
and U20413 (N_20413,N_16076,N_17081);
and U20414 (N_20414,N_12682,N_14133);
xor U20415 (N_20415,N_16328,N_12858);
and U20416 (N_20416,N_17940,N_15802);
and U20417 (N_20417,N_15031,N_16346);
nor U20418 (N_20418,N_16095,N_15925);
and U20419 (N_20419,N_14811,N_17359);
and U20420 (N_20420,N_18468,N_15849);
nor U20421 (N_20421,N_14482,N_14680);
nand U20422 (N_20422,N_15765,N_15629);
nand U20423 (N_20423,N_14305,N_13189);
or U20424 (N_20424,N_13551,N_17300);
xnor U20425 (N_20425,N_13296,N_16567);
nand U20426 (N_20426,N_13170,N_17487);
xnor U20427 (N_20427,N_15678,N_15234);
or U20428 (N_20428,N_12893,N_13700);
nor U20429 (N_20429,N_13668,N_18093);
nand U20430 (N_20430,N_16468,N_16405);
or U20431 (N_20431,N_12754,N_14137);
or U20432 (N_20432,N_12770,N_13662);
xnor U20433 (N_20433,N_16262,N_14283);
nor U20434 (N_20434,N_12593,N_18269);
or U20435 (N_20435,N_13317,N_15811);
nor U20436 (N_20436,N_18390,N_18330);
xnor U20437 (N_20437,N_17146,N_13283);
xnor U20438 (N_20438,N_13242,N_18384);
xnor U20439 (N_20439,N_17191,N_15804);
nand U20440 (N_20440,N_13717,N_18568);
or U20441 (N_20441,N_18263,N_15867);
nor U20442 (N_20442,N_15156,N_16770);
and U20443 (N_20443,N_17632,N_15254);
and U20444 (N_20444,N_15990,N_16303);
or U20445 (N_20445,N_17447,N_16749);
or U20446 (N_20446,N_17262,N_14987);
nor U20447 (N_20447,N_15269,N_13085);
and U20448 (N_20448,N_14525,N_16555);
nand U20449 (N_20449,N_13685,N_14678);
nor U20450 (N_20450,N_17669,N_18663);
or U20451 (N_20451,N_17681,N_13438);
or U20452 (N_20452,N_17508,N_17587);
xor U20453 (N_20453,N_13762,N_17485);
nor U20454 (N_20454,N_15058,N_13367);
nand U20455 (N_20455,N_18646,N_14000);
nand U20456 (N_20456,N_14052,N_14784);
and U20457 (N_20457,N_17982,N_14755);
and U20458 (N_20458,N_17864,N_18209);
or U20459 (N_20459,N_16375,N_16543);
or U20460 (N_20460,N_16190,N_12623);
or U20461 (N_20461,N_18215,N_12975);
nor U20462 (N_20462,N_15952,N_12708);
nor U20463 (N_20463,N_15038,N_15086);
nor U20464 (N_20464,N_13033,N_17091);
xnor U20465 (N_20465,N_18692,N_15935);
and U20466 (N_20466,N_16431,N_15583);
nor U20467 (N_20467,N_18731,N_16005);
or U20468 (N_20468,N_18661,N_18051);
or U20469 (N_20469,N_16339,N_17830);
and U20470 (N_20470,N_13845,N_15622);
nand U20471 (N_20471,N_15302,N_12742);
nand U20472 (N_20472,N_15639,N_18158);
or U20473 (N_20473,N_13112,N_13119);
and U20474 (N_20474,N_18040,N_13716);
and U20475 (N_20475,N_15141,N_15943);
xor U20476 (N_20476,N_15063,N_16359);
xnor U20477 (N_20477,N_17302,N_14543);
and U20478 (N_20478,N_15160,N_13339);
nor U20479 (N_20479,N_12704,N_17046);
or U20480 (N_20480,N_13539,N_14619);
or U20481 (N_20481,N_12775,N_17303);
nand U20482 (N_20482,N_15558,N_17763);
nor U20483 (N_20483,N_17511,N_12929);
xnor U20484 (N_20484,N_15801,N_14531);
or U20485 (N_20485,N_14560,N_17475);
and U20486 (N_20486,N_18718,N_13708);
and U20487 (N_20487,N_14629,N_17895);
nand U20488 (N_20488,N_15689,N_15870);
xor U20489 (N_20489,N_17445,N_13816);
nor U20490 (N_20490,N_12886,N_16333);
nand U20491 (N_20491,N_16122,N_17945);
nor U20492 (N_20492,N_17740,N_15079);
nor U20493 (N_20493,N_13855,N_15835);
xnor U20494 (N_20494,N_17038,N_14065);
and U20495 (N_20495,N_16043,N_14271);
xnor U20496 (N_20496,N_13298,N_18385);
nand U20497 (N_20497,N_16648,N_13651);
and U20498 (N_20498,N_16049,N_15041);
and U20499 (N_20499,N_18702,N_16010);
or U20500 (N_20500,N_14985,N_13248);
nor U20501 (N_20501,N_17052,N_14151);
nand U20502 (N_20502,N_13262,N_18486);
xor U20503 (N_20503,N_13519,N_15535);
nand U20504 (N_20504,N_16187,N_17355);
nor U20505 (N_20505,N_14222,N_18392);
xor U20506 (N_20506,N_15137,N_16577);
nor U20507 (N_20507,N_16841,N_12705);
nor U20508 (N_20508,N_17351,N_15425);
nor U20509 (N_20509,N_18031,N_17151);
or U20510 (N_20510,N_16820,N_13871);
or U20511 (N_20511,N_16748,N_15745);
or U20512 (N_20512,N_13598,N_13610);
and U20513 (N_20513,N_16861,N_16354);
and U20514 (N_20514,N_16935,N_14221);
or U20515 (N_20515,N_15719,N_14553);
nand U20516 (N_20516,N_16443,N_18559);
or U20517 (N_20517,N_16129,N_14524);
nor U20518 (N_20518,N_14781,N_17452);
nand U20519 (N_20519,N_13316,N_14575);
and U20520 (N_20520,N_12636,N_14529);
nor U20521 (N_20521,N_17244,N_15546);
nor U20522 (N_20522,N_18532,N_14785);
nand U20523 (N_20523,N_13201,N_14918);
xor U20524 (N_20524,N_13812,N_13932);
or U20525 (N_20525,N_17674,N_13436);
nor U20526 (N_20526,N_16836,N_15821);
nor U20527 (N_20527,N_15773,N_14798);
and U20528 (N_20528,N_15532,N_13508);
and U20529 (N_20529,N_18566,N_16278);
nand U20530 (N_20530,N_18474,N_16560);
and U20531 (N_20531,N_14293,N_16576);
nand U20532 (N_20532,N_15523,N_17963);
or U20533 (N_20533,N_16670,N_14033);
nand U20534 (N_20534,N_13864,N_16322);
nand U20535 (N_20535,N_13770,N_14637);
nand U20536 (N_20536,N_16826,N_12616);
xor U20537 (N_20537,N_15047,N_13027);
and U20538 (N_20538,N_16450,N_17111);
xor U20539 (N_20539,N_15524,N_14608);
xor U20540 (N_20540,N_15408,N_17630);
and U20541 (N_20541,N_14415,N_16388);
nand U20542 (N_20542,N_14214,N_12843);
and U20543 (N_20543,N_12643,N_13711);
nand U20544 (N_20544,N_16744,N_16887);
nor U20545 (N_20545,N_12513,N_15545);
xnor U20546 (N_20546,N_13145,N_14702);
xor U20547 (N_20547,N_14913,N_15838);
xor U20548 (N_20548,N_17374,N_15084);
nand U20549 (N_20549,N_18729,N_14881);
and U20550 (N_20550,N_16572,N_14241);
nor U20551 (N_20551,N_15391,N_13379);
xor U20552 (N_20552,N_16893,N_17718);
and U20553 (N_20553,N_13506,N_12782);
nor U20554 (N_20554,N_14666,N_16685);
nor U20555 (N_20555,N_17876,N_16078);
and U20556 (N_20556,N_15680,N_15032);
and U20557 (N_20557,N_15896,N_12626);
or U20558 (N_20558,N_13703,N_15734);
and U20559 (N_20559,N_16664,N_18651);
or U20560 (N_20560,N_18650,N_12905);
or U20561 (N_20561,N_12923,N_15991);
nand U20562 (N_20562,N_12544,N_17755);
or U20563 (N_20563,N_14196,N_13369);
or U20564 (N_20564,N_14579,N_14276);
or U20565 (N_20565,N_18141,N_18476);
xnor U20566 (N_20566,N_16021,N_16364);
or U20567 (N_20567,N_18536,N_14390);
nand U20568 (N_20568,N_15782,N_18412);
or U20569 (N_20569,N_17671,N_17458);
nor U20570 (N_20570,N_17656,N_13678);
and U20571 (N_20571,N_18230,N_15062);
and U20572 (N_20572,N_18426,N_15759);
nor U20573 (N_20573,N_18513,N_13012);
nor U20574 (N_20574,N_12564,N_16883);
or U20575 (N_20575,N_17507,N_14522);
nor U20576 (N_20576,N_15836,N_17147);
xor U20577 (N_20577,N_15865,N_15428);
or U20578 (N_20578,N_14961,N_16086);
xnor U20579 (N_20579,N_16867,N_14797);
nor U20580 (N_20580,N_12635,N_14633);
or U20581 (N_20581,N_17165,N_15380);
or U20582 (N_20582,N_17644,N_16394);
nor U20583 (N_20583,N_16628,N_18674);
and U20584 (N_20584,N_15480,N_12622);
and U20585 (N_20585,N_14202,N_16134);
and U20586 (N_20586,N_15947,N_16944);
nand U20587 (N_20587,N_15665,N_15590);
and U20588 (N_20588,N_17575,N_18621);
and U20589 (N_20589,N_13024,N_12566);
nor U20590 (N_20590,N_15364,N_13244);
and U20591 (N_20591,N_13435,N_17786);
nor U20592 (N_20592,N_12985,N_16847);
nor U20593 (N_20593,N_15048,N_17798);
nand U20594 (N_20594,N_12551,N_16601);
nand U20595 (N_20595,N_15381,N_18310);
and U20596 (N_20596,N_13301,N_18164);
and U20597 (N_20597,N_18168,N_15937);
or U20598 (N_20598,N_13629,N_15240);
xor U20599 (N_20599,N_17767,N_16153);
or U20600 (N_20600,N_17011,N_15286);
or U20601 (N_20601,N_15194,N_17811);
or U20602 (N_20602,N_14569,N_18272);
nand U20603 (N_20603,N_13384,N_16981);
xor U20604 (N_20604,N_18027,N_13468);
xor U20605 (N_20605,N_16891,N_18142);
xor U20606 (N_20606,N_16392,N_17881);
xor U20607 (N_20607,N_18707,N_14621);
nand U20608 (N_20608,N_13781,N_13873);
and U20609 (N_20609,N_17030,N_16853);
xnor U20610 (N_20610,N_13840,N_16223);
and U20611 (N_20611,N_15418,N_16838);
nor U20612 (N_20612,N_14116,N_15332);
or U20613 (N_20613,N_15565,N_14461);
nand U20614 (N_20614,N_16302,N_14874);
and U20615 (N_20615,N_16048,N_17444);
or U20616 (N_20616,N_17738,N_17771);
nor U20617 (N_20617,N_16424,N_14335);
nor U20618 (N_20618,N_14350,N_18387);
xnor U20619 (N_20619,N_16365,N_17377);
nor U20620 (N_20620,N_14897,N_14372);
nor U20621 (N_20621,N_12898,N_14308);
and U20622 (N_20622,N_14934,N_14073);
and U20623 (N_20623,N_16490,N_13571);
nand U20624 (N_20624,N_14671,N_17012);
or U20625 (N_20625,N_17420,N_18058);
nor U20626 (N_20626,N_16505,N_13587);
nor U20627 (N_20627,N_16387,N_15015);
or U20628 (N_20628,N_13092,N_15402);
and U20629 (N_20629,N_15628,N_16160);
or U20630 (N_20630,N_17765,N_17781);
and U20631 (N_20631,N_15809,N_14128);
xnor U20632 (N_20632,N_14030,N_14257);
and U20633 (N_20633,N_17555,N_15506);
or U20634 (N_20634,N_17736,N_14542);
and U20635 (N_20635,N_15505,N_16121);
nor U20636 (N_20636,N_18524,N_18627);
and U20637 (N_20637,N_13319,N_17693);
and U20638 (N_20638,N_15831,N_15542);
and U20639 (N_20639,N_16062,N_13279);
or U20640 (N_20640,N_18071,N_17382);
nand U20641 (N_20641,N_15901,N_17337);
and U20642 (N_20642,N_18602,N_18088);
and U20643 (N_20643,N_15450,N_16420);
nor U20644 (N_20644,N_17605,N_13760);
nor U20645 (N_20645,N_13995,N_13254);
xnor U20646 (N_20646,N_15556,N_18229);
xnor U20647 (N_20647,N_17196,N_13361);
nor U20648 (N_20648,N_14023,N_17641);
nor U20649 (N_20649,N_14540,N_12982);
nand U20650 (N_20650,N_17287,N_17773);
and U20651 (N_20651,N_18582,N_13683);
nor U20652 (N_20652,N_17947,N_17409);
nor U20653 (N_20653,N_15691,N_16080);
nor U20654 (N_20654,N_15006,N_17878);
nor U20655 (N_20655,N_13341,N_14598);
nand U20656 (N_20656,N_18197,N_15319);
xor U20657 (N_20657,N_14806,N_18688);
xor U20658 (N_20658,N_18289,N_12737);
or U20659 (N_20659,N_15318,N_13536);
or U20660 (N_20660,N_16667,N_12509);
xor U20661 (N_20661,N_18258,N_14058);
nor U20662 (N_20662,N_17315,N_16240);
xnor U20663 (N_20663,N_14519,N_18545);
nand U20664 (N_20664,N_17959,N_15738);
nor U20665 (N_20665,N_14656,N_12699);
and U20666 (N_20666,N_18267,N_14286);
nand U20667 (N_20667,N_16356,N_16411);
nand U20668 (N_20668,N_15913,N_16928);
nor U20669 (N_20669,N_14706,N_14887);
or U20670 (N_20670,N_14234,N_15929);
or U20671 (N_20671,N_15573,N_15763);
or U20672 (N_20672,N_18672,N_13643);
nor U20673 (N_20673,N_14238,N_17591);
nand U20674 (N_20674,N_12571,N_16916);
nand U20675 (N_20675,N_14216,N_15515);
nand U20676 (N_20676,N_14074,N_18091);
and U20677 (N_20677,N_13798,N_15536);
nor U20678 (N_20678,N_14427,N_15435);
and U20679 (N_20679,N_18069,N_13161);
nand U20680 (N_20680,N_13000,N_16285);
xnor U20681 (N_20681,N_16903,N_13935);
or U20682 (N_20682,N_15713,N_12696);
and U20683 (N_20683,N_17486,N_17025);
xor U20684 (N_20684,N_15907,N_13302);
xnor U20685 (N_20685,N_17680,N_14148);
nand U20686 (N_20686,N_15667,N_18512);
nor U20687 (N_20687,N_15298,N_15756);
nor U20688 (N_20688,N_17039,N_13772);
and U20689 (N_20689,N_13473,N_14361);
nor U20690 (N_20690,N_14366,N_13040);
xnor U20691 (N_20691,N_16414,N_15074);
xor U20692 (N_20692,N_17446,N_14174);
xor U20693 (N_20693,N_18309,N_13184);
nor U20694 (N_20694,N_14134,N_17795);
nor U20695 (N_20695,N_18232,N_14432);
and U20696 (N_20696,N_14152,N_14795);
or U20697 (N_20697,N_17942,N_16731);
nand U20698 (N_20698,N_13963,N_15092);
nor U20699 (N_20699,N_16586,N_13045);
nor U20700 (N_20700,N_15946,N_12799);
and U20701 (N_20701,N_15692,N_14796);
and U20702 (N_20702,N_14306,N_14688);
or U20703 (N_20703,N_15521,N_13933);
and U20704 (N_20704,N_18116,N_14692);
or U20705 (N_20705,N_14578,N_18157);
nand U20706 (N_20706,N_14590,N_18600);
xor U20707 (N_20707,N_16189,N_17757);
nor U20708 (N_20708,N_13199,N_15140);
nor U20709 (N_20709,N_16872,N_13485);
nand U20710 (N_20710,N_13970,N_17645);
and U20711 (N_20711,N_15294,N_17962);
nand U20712 (N_20712,N_18188,N_12695);
or U20713 (N_20713,N_14520,N_17995);
and U20714 (N_20714,N_18073,N_17310);
xnor U20715 (N_20715,N_17167,N_16488);
xor U20716 (N_20716,N_13314,N_18522);
nand U20717 (N_20717,N_15095,N_15096);
or U20718 (N_20718,N_13106,N_18687);
xor U20719 (N_20719,N_16097,N_17366);
nand U20720 (N_20720,N_13689,N_17832);
nor U20721 (N_20721,N_18082,N_14713);
or U20722 (N_20722,N_15251,N_17205);
xnor U20723 (N_20723,N_17143,N_14258);
and U20724 (N_20724,N_18726,N_18354);
nor U20725 (N_20725,N_13915,N_13126);
nor U20726 (N_20726,N_15447,N_17005);
or U20727 (N_20727,N_13867,N_17430);
and U20728 (N_20728,N_18050,N_15007);
and U20729 (N_20729,N_15540,N_14564);
nand U20730 (N_20730,N_13613,N_13486);
nor U20731 (N_20731,N_15954,N_17837);
and U20732 (N_20732,N_18053,N_13015);
or U20733 (N_20733,N_14969,N_13023);
or U20734 (N_20734,N_14681,N_15859);
and U20735 (N_20735,N_13591,N_14266);
nand U20736 (N_20736,N_17988,N_18440);
nor U20737 (N_20737,N_15684,N_17682);
or U20738 (N_20738,N_14660,N_14288);
xnor U20739 (N_20739,N_17574,N_13990);
or U20740 (N_20740,N_13401,N_14880);
nor U20741 (N_20741,N_14001,N_18286);
and U20742 (N_20742,N_14173,N_18251);
or U20743 (N_20743,N_16242,N_15909);
xor U20744 (N_20744,N_17480,N_17383);
or U20745 (N_20745,N_16513,N_16362);
or U20746 (N_20746,N_17961,N_16119);
xnor U20747 (N_20747,N_16676,N_16493);
or U20748 (N_20748,N_18256,N_18217);
xor U20749 (N_20749,N_18749,N_17770);
or U20750 (N_20750,N_16248,N_12875);
nor U20751 (N_20751,N_17577,N_17276);
xor U20752 (N_20752,N_13870,N_13897);
and U20753 (N_20753,N_15894,N_18030);
or U20754 (N_20754,N_17901,N_15190);
nor U20755 (N_20755,N_14507,N_14106);
nand U20756 (N_20756,N_16044,N_18386);
and U20757 (N_20757,N_17499,N_12670);
or U20758 (N_20758,N_13352,N_17955);
or U20759 (N_20759,N_16518,N_15466);
nor U20760 (N_20760,N_18023,N_15772);
nor U20761 (N_20761,N_13131,N_14497);
nor U20762 (N_20762,N_13157,N_17617);
xor U20763 (N_20763,N_14045,N_17893);
nor U20764 (N_20764,N_13584,N_12630);
nand U20765 (N_20765,N_13583,N_14077);
or U20766 (N_20766,N_12581,N_14047);
and U20767 (N_20767,N_16342,N_18257);
nand U20768 (N_20768,N_18355,N_13921);
or U20769 (N_20769,N_14484,N_14532);
nor U20770 (N_20770,N_13552,N_17016);
nor U20771 (N_20771,N_17624,N_17532);
nand U20772 (N_20772,N_16463,N_15888);
or U20773 (N_20773,N_17573,N_14725);
nor U20774 (N_20774,N_16800,N_16774);
xor U20775 (N_20775,N_14356,N_16918);
and U20776 (N_20776,N_16595,N_14581);
and U20777 (N_20777,N_18179,N_13125);
nand U20778 (N_20778,N_15903,N_14675);
nand U20779 (N_20779,N_14325,N_14360);
or U20780 (N_20780,N_15816,N_13364);
or U20781 (N_20781,N_12591,N_18367);
nor U20782 (N_20782,N_15138,N_15091);
or U20783 (N_20783,N_14090,N_12808);
nor U20784 (N_20784,N_13941,N_14883);
nor U20785 (N_20785,N_13439,N_18695);
nand U20786 (N_20786,N_13597,N_16451);
nand U20787 (N_20787,N_16581,N_16958);
and U20788 (N_20788,N_14815,N_13190);
nand U20789 (N_20789,N_13136,N_16166);
xnor U20790 (N_20790,N_17400,N_17653);
and U20791 (N_20791,N_16218,N_14329);
and U20792 (N_20792,N_13730,N_18183);
and U20793 (N_20793,N_15003,N_16348);
and U20794 (N_20794,N_15674,N_15059);
xor U20795 (N_20795,N_18727,N_14697);
nand U20796 (N_20796,N_15330,N_15602);
and U20797 (N_20797,N_14703,N_17853);
or U20798 (N_20798,N_15385,N_16209);
and U20799 (N_20799,N_15770,N_14707);
nor U20800 (N_20800,N_13984,N_13910);
nand U20801 (N_20801,N_12994,N_15788);
or U20802 (N_20802,N_15750,N_17228);
or U20803 (N_20803,N_17649,N_13135);
nor U20804 (N_20804,N_14010,N_14192);
or U20805 (N_20805,N_17535,N_15139);
xor U20806 (N_20806,N_15951,N_17912);
nor U20807 (N_20807,N_18411,N_17433);
nor U20808 (N_20808,N_15118,N_17203);
or U20809 (N_20809,N_13447,N_13357);
or U20810 (N_20810,N_14963,N_15735);
and U20811 (N_20811,N_16514,N_13162);
or U20812 (N_20812,N_17092,N_13327);
xnor U20813 (N_20813,N_15722,N_13879);
xnor U20814 (N_20814,N_18547,N_17341);
nor U20815 (N_20815,N_13558,N_12959);
or U20816 (N_20816,N_14846,N_13259);
nor U20817 (N_20817,N_16504,N_12762);
or U20818 (N_20818,N_12846,N_15595);
or U20819 (N_20819,N_13177,N_13270);
or U20820 (N_20820,N_17710,N_14462);
or U20821 (N_20821,N_17908,N_18730);
or U20822 (N_20822,N_16804,N_15043);
xor U20823 (N_20823,N_15701,N_13532);
and U20824 (N_20824,N_12851,N_14075);
nor U20825 (N_20825,N_17048,N_14095);
and U20826 (N_20826,N_13061,N_14413);
and U20827 (N_20827,N_14940,N_16902);
nand U20828 (N_20828,N_15820,N_18271);
or U20829 (N_20829,N_13776,N_14407);
xor U20830 (N_20830,N_15119,N_14776);
or U20831 (N_20831,N_16400,N_13241);
xnor U20832 (N_20832,N_16638,N_18574);
and U20833 (N_20833,N_15757,N_15785);
nand U20834 (N_20834,N_12721,N_12638);
xor U20835 (N_20835,N_12540,N_15620);
or U20836 (N_20836,N_12531,N_17028);
nand U20837 (N_20837,N_16659,N_16371);
nand U20838 (N_20838,N_15862,N_18507);
xor U20839 (N_20839,N_17421,N_16540);
xor U20840 (N_20840,N_15707,N_13698);
or U20841 (N_20841,N_17271,N_13563);
nand U20842 (N_20842,N_15726,N_16782);
and U20843 (N_20843,N_12823,N_13785);
or U20844 (N_20844,N_15267,N_13722);
nand U20845 (N_20845,N_17546,N_15195);
and U20846 (N_20846,N_17966,N_17093);
or U20847 (N_20847,N_17544,N_16444);
nand U20848 (N_20848,N_17116,N_17235);
nor U20849 (N_20849,N_15366,N_17223);
and U20850 (N_20850,N_14468,N_17141);
nand U20851 (N_20851,N_13817,N_16900);
or U20852 (N_20852,N_15307,N_17515);
xor U20853 (N_20853,N_16724,N_16665);
or U20854 (N_20854,N_18139,N_17687);
and U20855 (N_20855,N_15601,N_13593);
and U20856 (N_20856,N_13939,N_14505);
nand U20857 (N_20857,N_16617,N_18515);
and U20858 (N_20858,N_18684,N_17621);
nor U20859 (N_20859,N_15637,N_16306);
xor U20860 (N_20860,N_14494,N_17672);
or U20861 (N_20861,N_12734,N_13846);
or U20862 (N_20862,N_16406,N_18149);
nand U20863 (N_20863,N_16580,N_16382);
nand U20864 (N_20864,N_13405,N_13031);
nand U20865 (N_20865,N_18736,N_18526);
xor U20866 (N_20866,N_17035,N_14428);
nand U20867 (N_20867,N_18576,N_13904);
nor U20868 (N_20868,N_13207,N_18430);
nor U20869 (N_20869,N_17273,N_16372);
nand U20870 (N_20870,N_17526,N_13103);
nor U20871 (N_20871,N_16582,N_16592);
nand U20872 (N_20872,N_13455,N_14658);
or U20873 (N_20873,N_17910,N_17328);
xor U20874 (N_20874,N_15995,N_12828);
or U20875 (N_20875,N_13676,N_16330);
nor U20876 (N_20876,N_17792,N_17777);
nand U20877 (N_20877,N_15824,N_13402);
and U20878 (N_20878,N_18226,N_17551);
xor U20879 (N_20879,N_16764,N_17393);
nand U20880 (N_20880,N_15592,N_14044);
xor U20881 (N_20881,N_15280,N_17260);
nor U20882 (N_20882,N_13196,N_14226);
nand U20883 (N_20883,N_16794,N_12888);
and U20884 (N_20884,N_17531,N_18111);
and U20885 (N_20885,N_14348,N_14122);
and U20886 (N_20886,N_13572,N_14954);
nand U20887 (N_20887,N_18320,N_17348);
nor U20888 (N_20888,N_18039,N_16065);
or U20889 (N_20889,N_13062,N_14437);
xor U20890 (N_20890,N_15321,N_17363);
or U20891 (N_20891,N_17698,N_17352);
nor U20892 (N_20892,N_18171,N_17633);
xnor U20893 (N_20893,N_15042,N_16695);
xnor U20894 (N_20894,N_13979,N_15703);
or U20895 (N_20895,N_17150,N_12615);
nand U20896 (N_20896,N_18255,N_17849);
xor U20897 (N_20897,N_15354,N_17174);
xnor U20898 (N_20898,N_17193,N_13671);
or U20899 (N_20899,N_18458,N_16224);
nor U20900 (N_20900,N_13752,N_18598);
nor U20901 (N_20901,N_17583,N_15389);
nand U20902 (N_20902,N_12683,N_17614);
xnor U20903 (N_20903,N_12793,N_15636);
nor U20904 (N_20904,N_15923,N_12653);
xnor U20905 (N_20905,N_14694,N_15973);
and U20906 (N_20906,N_16681,N_14456);
nor U20907 (N_20907,N_15045,N_13673);
or U20908 (N_20908,N_18081,N_16161);
or U20909 (N_20909,N_18299,N_16996);
nand U20910 (N_20910,N_17384,N_15698);
and U20911 (N_20911,N_17123,N_18110);
xor U20912 (N_20912,N_18457,N_17565);
xor U20913 (N_20913,N_15514,N_17050);
nor U20914 (N_20914,N_17949,N_17503);
or U20915 (N_20915,N_17647,N_13498);
xnor U20916 (N_20916,N_13424,N_15224);
xor U20917 (N_20917,N_14218,N_17581);
xor U20918 (N_20918,N_18482,N_12692);
xnor U20919 (N_20919,N_14696,N_15416);
and U20920 (N_20920,N_14138,N_17697);
nor U20921 (N_20921,N_16525,N_17301);
and U20922 (N_20922,N_16756,N_17220);
nor U20923 (N_20923,N_17069,N_15409);
xor U20924 (N_20924,N_18326,N_13821);
and U20925 (N_20925,N_15209,N_18266);
xor U20926 (N_20926,N_13878,N_16351);
and U20927 (N_20927,N_17886,N_18697);
nand U20928 (N_20928,N_13222,N_15586);
xnor U20929 (N_20929,N_12725,N_13223);
nand U20930 (N_20930,N_14009,N_18700);
xor U20931 (N_20931,N_16721,N_14727);
and U20932 (N_20932,N_14873,N_14805);
and U20933 (N_20933,N_12515,N_13358);
xnor U20934 (N_20934,N_15900,N_13839);
nand U20935 (N_20935,N_16196,N_15221);
or U20936 (N_20936,N_14287,N_18112);
and U20937 (N_20937,N_17222,N_16686);
and U20938 (N_20938,N_13413,N_15277);
nand U20939 (N_20939,N_16510,N_13617);
xor U20940 (N_20940,N_12656,N_15282);
nand U20941 (N_20941,N_15169,N_13947);
or U20942 (N_20942,N_18379,N_17695);
nor U20943 (N_20943,N_14834,N_16022);
and U20944 (N_20944,N_14323,N_16089);
and U20945 (N_20945,N_16503,N_17734);
and U20946 (N_20946,N_14941,N_16390);
or U20947 (N_20947,N_14021,N_17545);
and U20948 (N_20948,N_14167,N_14168);
nand U20949 (N_20949,N_15404,N_13220);
or U20950 (N_20950,N_18712,N_15577);
nor U20951 (N_20951,N_12693,N_13579);
xnor U20952 (N_20952,N_16195,N_18045);
nand U20953 (N_20953,N_16717,N_13978);
nor U20954 (N_20954,N_15462,N_12792);
xor U20955 (N_20955,N_12956,N_15446);
and U20956 (N_20956,N_15988,N_15635);
and U20957 (N_20957,N_12980,N_12873);
nand U20958 (N_20958,N_17218,N_15748);
xnor U20959 (N_20959,N_16811,N_15372);
and U20960 (N_20960,N_16491,N_16630);
nor U20961 (N_20961,N_13814,N_18319);
xnor U20962 (N_20962,N_16373,N_15490);
nand U20963 (N_20963,N_13310,N_14879);
or U20964 (N_20964,N_14199,N_12860);
nand U20965 (N_20965,N_13608,N_12588);
and U20966 (N_20966,N_14206,N_16511);
and U20967 (N_20967,N_15999,N_12827);
and U20968 (N_20968,N_16989,N_14927);
nor U20969 (N_20969,N_13088,N_14778);
or U20970 (N_20970,N_16475,N_14835);
nor U20971 (N_20971,N_17152,N_13646);
or U20972 (N_20972,N_18500,N_13492);
nand U20973 (N_20973,N_16959,N_16184);
and U20974 (N_20974,N_17371,N_15837);
nand U20975 (N_20975,N_13163,N_15563);
and U20976 (N_20976,N_15186,N_14731);
nor U20977 (N_20977,N_17250,N_12983);
or U20978 (N_20978,N_18243,N_16835);
nor U20979 (N_20979,N_13240,N_13311);
or U20980 (N_20980,N_17243,N_14551);
and U20981 (N_20981,N_14048,N_18314);
or U20982 (N_20982,N_15103,N_17839);
xor U20983 (N_20983,N_13107,N_15529);
or U20984 (N_20984,N_17506,N_14710);
nor U20985 (N_20985,N_12771,N_14612);
xnor U20986 (N_20986,N_15779,N_14800);
nor U20987 (N_20987,N_14643,N_13232);
nand U20988 (N_20988,N_13605,N_14249);
nor U20989 (N_20989,N_16528,N_15377);
and U20990 (N_20990,N_17206,N_18461);
or U20991 (N_20991,N_13501,N_15673);
nor U20992 (N_20992,N_18746,N_17219);
or U20993 (N_20993,N_13739,N_17484);
nand U20994 (N_20994,N_12958,N_16750);
nand U20995 (N_20995,N_13741,N_16436);
and U20996 (N_20996,N_16656,N_12601);
nand U20997 (N_20997,N_17980,N_16395);
nor U20998 (N_20998,N_16284,N_16438);
or U20999 (N_20999,N_14421,N_14291);
and U21000 (N_21000,N_15714,N_17858);
nand U21001 (N_21001,N_15994,N_16738);
nand U21002 (N_21002,N_17022,N_16791);
or U21003 (N_21003,N_14668,N_14092);
and U21004 (N_21004,N_16131,N_16178);
xor U21005 (N_21005,N_17860,N_12661);
and U21006 (N_21006,N_14149,N_14082);
nor U21007 (N_21007,N_14832,N_15685);
nand U21008 (N_21008,N_13371,N_13117);
xnor U21009 (N_21009,N_16249,N_18096);
and U21010 (N_21010,N_17094,N_13968);
xnor U21011 (N_21011,N_14844,N_12627);
and U21012 (N_21012,N_18278,N_18288);
xor U21013 (N_21013,N_18581,N_16253);
xor U21014 (N_21014,N_13512,N_18408);
xor U21015 (N_21015,N_15612,N_17523);
nand U21016 (N_21016,N_12987,N_15122);
xnor U21017 (N_21017,N_12921,N_15171);
or U21018 (N_21018,N_17782,N_15997);
nand U21019 (N_21019,N_17918,N_14807);
nand U21020 (N_21020,N_15075,N_14981);
and U21021 (N_21021,N_18683,N_14506);
nor U21022 (N_21022,N_13621,N_15036);
or U21023 (N_21023,N_16589,N_13108);
nor U21024 (N_21024,N_17238,N_12972);
xnor U21025 (N_21025,N_14650,N_18643);
or U21026 (N_21026,N_12891,N_18132);
nor U21027 (N_21027,N_15564,N_12826);
nand U21028 (N_21028,N_17994,N_16280);
nor U21029 (N_21029,N_16991,N_15706);
or U21030 (N_21030,N_16641,N_17122);
xnor U21031 (N_21031,N_16439,N_15440);
and U21032 (N_21032,N_15603,N_17664);
nor U21033 (N_21033,N_16913,N_12579);
and U21034 (N_21034,N_12844,N_15887);
nand U21035 (N_21035,N_13710,N_13813);
xor U21036 (N_21036,N_12791,N_15028);
xor U21037 (N_21037,N_16363,N_16720);
nor U21038 (N_21038,N_16255,N_15916);
nand U21039 (N_21039,N_13914,N_16827);
nand U21040 (N_21040,N_13799,N_18204);
and U21041 (N_21041,N_18561,N_17958);
xnor U21042 (N_21042,N_18371,N_15076);
nand U21043 (N_21043,N_14973,N_18580);
nor U21044 (N_21044,N_12587,N_14479);
nor U21045 (N_21045,N_13430,N_15250);
and U21046 (N_21046,N_13959,N_18456);
nor U21047 (N_21047,N_13309,N_15744);
or U21048 (N_21048,N_17778,N_14176);
nand U21049 (N_21049,N_15872,N_13580);
nor U21050 (N_21050,N_16176,N_16061);
nor U21051 (N_21051,N_14585,N_14935);
nand U21052 (N_21052,N_15155,N_17098);
or U21053 (N_21053,N_17034,N_13137);
and U21054 (N_21054,N_14905,N_17539);
and U21055 (N_21055,N_13360,N_18297);
or U21056 (N_21056,N_17442,N_17202);
nor U21057 (N_21057,N_18514,N_13773);
xnor U21058 (N_21058,N_17871,N_13477);
nor U21059 (N_21059,N_17751,N_15046);
or U21060 (N_21060,N_13461,N_13693);
or U21061 (N_21061,N_16261,N_18665);
nand U21062 (N_21062,N_13554,N_16661);
nor U21063 (N_21063,N_14754,N_13849);
nand U21064 (N_21064,N_16674,N_17157);
or U21065 (N_21065,N_14794,N_16534);
and U21066 (N_21066,N_17789,N_13511);
nor U21067 (N_21067,N_16257,N_15696);
or U21068 (N_21068,N_12880,N_15168);
nand U21069 (N_21069,N_18591,N_16212);
nand U21070 (N_21070,N_17809,N_18694);
or U21071 (N_21071,N_14739,N_15019);
nor U21072 (N_21072,N_13073,N_17726);
and U21073 (N_21073,N_16163,N_16644);
xor U21074 (N_21074,N_16658,N_15566);
nor U21075 (N_21075,N_13273,N_16055);
or U21076 (N_21076,N_13815,N_14876);
and U21077 (N_21077,N_17291,N_13036);
xnor U21078 (N_21078,N_12538,N_15544);
and U21079 (N_21079,N_13264,N_17776);
or U21080 (N_21080,N_12609,N_13153);
xor U21081 (N_21081,N_17704,N_14060);
nor U21082 (N_21082,N_13102,N_13235);
nand U21083 (N_21083,N_13100,N_18709);
or U21084 (N_21084,N_14711,N_14733);
nand U21085 (N_21085,N_17749,N_12523);
nor U21086 (N_21086,N_16243,N_18207);
or U21087 (N_21087,N_15399,N_16266);
or U21088 (N_21088,N_18389,N_18170);
and U21089 (N_21089,N_14395,N_13420);
or U21090 (N_21090,N_13642,N_16778);
xor U21091 (N_21091,N_15718,N_14046);
or U21092 (N_21092,N_16568,N_14170);
nor U21093 (N_21093,N_18448,N_17902);
and U21094 (N_21094,N_18378,N_15373);
xnor U21095 (N_21095,N_12922,N_17375);
nor U21096 (N_21096,N_14328,N_13457);
or U21097 (N_21097,N_14849,N_17607);
nor U21098 (N_21098,N_18609,N_17213);
and U21099 (N_21099,N_18682,N_15600);
and U21100 (N_21100,N_14889,N_15522);
or U21101 (N_21101,N_18706,N_15316);
and U21102 (N_21102,N_18018,N_15236);
nor U21103 (N_21103,N_13030,N_16898);
nand U21104 (N_21104,N_16177,N_14477);
xor U21105 (N_21105,N_16456,N_13582);
nor U21106 (N_21106,N_13516,N_16758);
nor U21107 (N_21107,N_18447,N_15444);
and U21108 (N_21108,N_16230,N_17232);
nand U21109 (N_21109,N_15609,N_16559);
or U21110 (N_21110,N_15383,N_18029);
or U21111 (N_21111,N_17666,N_12586);
nand U21112 (N_21112,N_18634,N_13573);
nand U21113 (N_21113,N_13083,N_13347);
or U21114 (N_21114,N_15008,N_17212);
or U21115 (N_21115,N_18599,N_15388);
nor U21116 (N_21116,N_18160,N_17240);
nand U21117 (N_21117,N_13960,N_17169);
and U21118 (N_21118,N_13029,N_17451);
nor U21119 (N_21119,N_14375,N_13091);
and U21120 (N_21120,N_13826,N_18528);
nand U21121 (N_21121,N_14914,N_13966);
xnor U21122 (N_21122,N_14641,N_14767);
xnor U21123 (N_21123,N_13276,N_18483);
or U21124 (N_21124,N_16753,N_17834);
xnor U21125 (N_21125,N_18056,N_15304);
nand U21126 (N_21126,N_16353,N_14493);
nor U21127 (N_21127,N_13880,N_15243);
nand U21128 (N_21128,N_15001,N_14837);
nor U21129 (N_21129,N_16082,N_18432);
and U21130 (N_21130,N_15516,N_15783);
nor U21131 (N_21131,N_17579,N_18292);
nor U21132 (N_21132,N_12550,N_17585);
and U21133 (N_21133,N_17282,N_18274);
or U21134 (N_21134,N_16621,N_14726);
nor U21135 (N_21135,N_12642,N_18615);
and U21136 (N_21136,N_17084,N_16321);
and U21137 (N_21137,N_13649,N_15908);
nor U21138 (N_21138,N_12702,N_12602);
and U21139 (N_21139,N_14383,N_17285);
nor U21140 (N_21140,N_16538,N_16004);
nor U21141 (N_21141,N_17800,N_16474);
xor U21142 (N_21142,N_17378,N_16361);
nor U21143 (N_21143,N_14965,N_18479);
nand U21144 (N_21144,N_14558,N_14943);
nor U21145 (N_21145,N_17057,N_17670);
nand U21146 (N_21146,N_18630,N_18571);
or U21147 (N_21147,N_17438,N_15167);
nand U21148 (N_21148,N_16529,N_16516);
and U21149 (N_21149,N_17448,N_17437);
and U21150 (N_21150,N_14248,N_16596);
nor U21151 (N_21151,N_18679,N_14302);
nor U21152 (N_21152,N_18151,N_15847);
and U21153 (N_21153,N_14983,N_16755);
or U21154 (N_21154,N_18011,N_17564);
nor U21155 (N_21155,N_14872,N_13230);
or U21156 (N_21156,N_12896,N_17676);
nand U21157 (N_21157,N_17460,N_16696);
and U21158 (N_21158,N_16982,N_17505);
or U21159 (N_21159,N_12964,N_13882);
nor U21160 (N_21160,N_18087,N_15668);
nor U21161 (N_21161,N_16803,N_14890);
and U21162 (N_21162,N_14690,N_17863);
or U21163 (N_21163,N_14392,N_18647);
and U21164 (N_21164,N_16710,N_16997);
and U21165 (N_21165,N_17629,N_16092);
and U21166 (N_21166,N_14135,N_18161);
xor U21167 (N_21167,N_17626,N_13844);
nor U21168 (N_21168,N_12861,N_16743);
and U21169 (N_21169,N_15784,N_14154);
xor U21170 (N_21170,N_14412,N_17648);
nand U21171 (N_21171,N_16492,N_13078);
or U21172 (N_21172,N_18366,N_14108);
or U21173 (N_21173,N_17668,N_14528);
and U21174 (N_21174,N_17017,N_12876);
nor U21175 (N_21175,N_17872,N_16329);
or U21176 (N_21176,N_16428,N_13071);
nand U21177 (N_21177,N_15430,N_16128);
xnor U21178 (N_21178,N_17894,N_18613);
and U21179 (N_21179,N_13169,N_13287);
xnor U21180 (N_21180,N_13118,N_13569);
and U21181 (N_21181,N_17071,N_17622);
xnor U21182 (N_21182,N_17186,N_17060);
or U21183 (N_21183,N_17019,N_15011);
nor U21184 (N_21184,N_18331,N_17692);
and U21185 (N_21185,N_15513,N_15981);
nand U21186 (N_21186,N_16718,N_14032);
or U21187 (N_21187,N_17552,N_16198);
nor U21188 (N_21188,N_15778,N_14956);
xnor U21189 (N_21189,N_18465,N_17173);
nor U21190 (N_21190,N_14110,N_16825);
or U21191 (N_21191,N_14094,N_13269);
or U21192 (N_21192,N_12862,N_15823);
nor U21193 (N_21193,N_18037,N_18662);
nor U21194 (N_21194,N_15803,N_17255);
nand U21195 (N_21195,N_14056,N_17294);
and U21196 (N_21196,N_13323,N_15571);
nand U21197 (N_21197,N_18381,N_12911);
nor U21198 (N_21198,N_15394,N_17051);
nand U21199 (N_21199,N_13282,N_17720);
nor U21200 (N_21200,N_16147,N_13382);
nand U21201 (N_21201,N_17769,N_17037);
xor U21202 (N_21202,N_12939,N_12684);
nor U21203 (N_21203,N_14136,N_13245);
and U21204 (N_21204,N_15403,N_18283);
or U21205 (N_21205,N_15004,N_12895);
and U21206 (N_21206,N_17997,N_16557);
or U21207 (N_21207,N_16862,N_12784);
and U21208 (N_21208,N_13488,N_16148);
or U21209 (N_21209,N_18453,N_13833);
xor U21210 (N_21210,N_17794,N_18395);
and U21211 (N_21211,N_13095,N_14843);
xnor U21212 (N_21212,N_14848,N_16609);
and U21213 (N_21213,N_18460,N_14665);
and U21214 (N_21214,N_18374,N_17847);
nand U21215 (N_21215,N_15944,N_15281);
nor U21216 (N_21216,N_18281,N_12937);
nand U21217 (N_21217,N_16635,N_16956);
nand U21218 (N_21218,N_16858,N_12840);
and U21219 (N_21219,N_12881,N_13823);
and U21220 (N_21220,N_16060,N_17096);
xnor U21221 (N_21221,N_13758,N_17233);
and U21222 (N_21222,N_15519,N_14280);
nor U21223 (N_21223,N_16467,N_18564);
nor U21224 (N_21224,N_13555,N_18705);
nand U21225 (N_21225,N_17824,N_12910);
xnor U21226 (N_21226,N_16175,N_15642);
xnor U21227 (N_21227,N_17534,N_14992);
and U21228 (N_21228,N_12585,N_16067);
and U21229 (N_21229,N_13858,N_14243);
nor U21230 (N_21230,N_16256,N_15393);
or U21231 (N_21231,N_16104,N_15771);
nand U21232 (N_21232,N_13987,N_14863);
xnor U21233 (N_21233,N_17214,N_15626);
nor U21234 (N_21234,N_17557,N_15145);
and U21235 (N_21235,N_14549,N_12558);
nand U21236 (N_21236,N_16602,N_16948);
nand U21237 (N_21237,N_15729,N_18473);
and U21238 (N_21238,N_16864,N_18567);
and U21239 (N_21239,N_13143,N_18306);
nor U21240 (N_21240,N_16066,N_17900);
xor U21241 (N_21241,N_17086,N_13779);
or U21242 (N_21242,N_13253,N_18667);
nand U21243 (N_21243,N_13628,N_15646);
nor U21244 (N_21244,N_18541,N_15731);
and U21245 (N_21245,N_18193,N_18080);
or U21246 (N_21246,N_13884,N_14877);
xnor U21247 (N_21247,N_14942,N_18034);
nor U21248 (N_21248,N_14264,N_16376);
nand U21249 (N_21249,N_16732,N_16619);
xnor U21250 (N_21250,N_14141,N_13005);
and U21251 (N_21251,N_13896,N_13822);
or U21252 (N_21252,N_17135,N_16542);
and U21253 (N_21253,N_15345,N_13705);
and U21254 (N_21254,N_13534,N_16366);
nor U21255 (N_21255,N_17635,N_14178);
nor U21256 (N_21256,N_16032,N_15002);
and U21257 (N_21257,N_16279,N_13326);
and U21258 (N_21258,N_17498,N_15314);
nand U21259 (N_21259,N_15845,N_17590);
and U21260 (N_21260,N_17058,N_15974);
xor U21261 (N_21261,N_15457,N_16590);
nand U21262 (N_21262,N_16912,N_16105);
and U21263 (N_21263,N_18502,N_13224);
or U21264 (N_21264,N_14500,N_17701);
nand U21265 (N_21265,N_18585,N_18578);
xor U21266 (N_21266,N_15360,N_16709);
and U21267 (N_21267,N_16227,N_13013);
nand U21268 (N_21268,N_14020,N_12713);
xor U21269 (N_21269,N_12613,N_17700);
xor U21270 (N_21270,N_14672,N_12516);
nor U21271 (N_21271,N_13594,N_17089);
or U21272 (N_21272,N_18652,N_14989);
or U21273 (N_21273,N_16118,N_13634);
xnor U21274 (N_21274,N_16472,N_13887);
nand U21275 (N_21275,N_13943,N_13047);
nor U21276 (N_21276,N_12530,N_18109);
or U21277 (N_21277,N_17090,N_18464);
xor U21278 (N_21278,N_15796,N_13602);
nor U21279 (N_21279,N_17489,N_18407);
nor U21280 (N_21280,N_14105,N_14342);
nand U21281 (N_21281,N_16193,N_17721);
nor U21282 (N_21282,N_14939,N_12882);
xnor U21283 (N_21283,N_14357,N_13802);
nor U21284 (N_21284,N_13116,N_13236);
nor U21285 (N_21285,N_13122,N_14359);
or U21286 (N_21286,N_13214,N_14391);
nand U21287 (N_21287,N_13727,N_13391);
nand U21288 (N_21288,N_16963,N_14845);
or U21289 (N_21289,N_12510,N_14452);
nand U21290 (N_21290,N_17835,N_15005);
nor U21291 (N_21291,N_14182,N_14604);
nor U21292 (N_21292,N_12928,N_16482);
xnor U21293 (N_21293,N_18127,N_16834);
or U21294 (N_21294,N_14606,N_14904);
or U21295 (N_21295,N_15662,N_18362);
or U21296 (N_21296,N_18231,N_15296);
xnor U21297 (N_21297,N_17414,N_12787);
nand U21298 (N_21298,N_15226,N_17880);
and U21299 (N_21299,N_18075,N_18626);
nor U21300 (N_21300,N_17320,N_17115);
xor U21301 (N_21301,N_17450,N_15262);
and U21302 (N_21302,N_12849,N_13792);
or U21303 (N_21303,N_14919,N_14986);
xor U21304 (N_21304,N_14053,N_13940);
nand U21305 (N_21305,N_17170,N_14388);
or U21306 (N_21306,N_14533,N_15121);
or U21307 (N_21307,N_13989,N_16250);
or U21308 (N_21308,N_18305,N_18057);
or U21309 (N_21309,N_14730,N_14051);
and U21310 (N_21310,N_12631,N_16462);
or U21311 (N_21311,N_13226,N_14463);
nor U21312 (N_21312,N_13072,N_12722);
xnor U21313 (N_21313,N_14403,N_17923);
nor U21314 (N_21314,N_14472,N_16920);
and U21315 (N_21315,N_14960,N_13803);
nor U21316 (N_21316,N_13886,N_16578);
nor U21317 (N_21317,N_16704,N_16923);
nor U21318 (N_21318,N_17168,N_13257);
nor U21319 (N_21319,N_16287,N_17140);
or U21320 (N_21320,N_16823,N_13973);
xnor U21321 (N_21321,N_14054,N_15488);
and U21322 (N_21322,N_17643,N_12814);
xnor U21323 (N_21323,N_17431,N_18635);
nor U21324 (N_21324,N_15996,N_14704);
nor U21325 (N_21325,N_14368,N_14409);
and U21326 (N_21326,N_14878,N_12817);
nor U21327 (N_21327,N_13647,N_15899);
nand U21328 (N_21328,N_16856,N_14962);
xor U21329 (N_21329,N_13229,N_15455);
and U21330 (N_21330,N_12872,N_13121);
nand U21331 (N_21331,N_14916,N_14439);
xor U21332 (N_21332,N_16974,N_15539);
or U21333 (N_21333,N_14997,N_13874);
and U21334 (N_21334,N_15649,N_18611);
xor U21335 (N_21335,N_14292,N_14346);
nand U21336 (N_21336,N_16549,N_14349);
nor U21337 (N_21337,N_12768,N_12590);
xor U21338 (N_21338,N_15297,N_17911);
or U21339 (N_21339,N_13648,N_16850);
nor U21340 (N_21340,N_16574,N_14899);
nor U21341 (N_21341,N_18176,N_16679);
nand U21342 (N_21342,N_17185,N_13164);
nor U21343 (N_21343,N_17155,N_17465);
or U21344 (N_21344,N_18610,N_17787);
and U21345 (N_21345,N_16220,N_18280);
xnor U21346 (N_21346,N_15111,N_15220);
or U21347 (N_21347,N_17397,N_14810);
nand U21348 (N_21348,N_15933,N_14163);
and U21349 (N_21349,N_15538,N_17964);
nand U21350 (N_21350,N_14414,N_17246);
nor U21351 (N_21351,N_17160,N_16980);
nor U21352 (N_21352,N_18451,N_18490);
or U21353 (N_21353,N_18516,N_18077);
xnor U21354 (N_21354,N_13547,N_18219);
and U21355 (N_21355,N_14991,N_13266);
nor U21356 (N_21356,N_14803,N_15740);
and U21357 (N_21357,N_18537,N_18293);
nand U21358 (N_21358,N_18666,N_13022);
and U21359 (N_21359,N_15830,N_15554);
xnor U21360 (N_21360,N_14212,N_13586);
and U21361 (N_21361,N_18173,N_14097);
or U21362 (N_21362,N_15604,N_15877);
nor U21363 (N_21363,N_17707,N_12835);
nor U21364 (N_21364,N_15598,N_14485);
nor U21365 (N_21365,N_17308,N_12723);
and U21366 (N_21366,N_12744,N_14625);
or U21367 (N_21367,N_16041,N_14642);
and U21368 (N_21368,N_13247,N_16895);
nand U21369 (N_21369,N_13653,N_17619);
or U21370 (N_21370,N_13018,N_18711);
and U21371 (N_21371,N_15064,N_14850);
nor U21372 (N_21372,N_14698,N_14181);
xor U21373 (N_21373,N_14651,N_13930);
xor U21374 (N_21374,N_16614,N_18563);
and U21375 (N_21375,N_16684,N_16689);
xnor U21376 (N_21376,N_12654,N_17812);
and U21377 (N_21377,N_15893,N_17851);
and U21378 (N_21378,N_16246,N_18416);
or U21379 (N_21379,N_16625,N_18550);
nor U21380 (N_21380,N_16347,N_15623);
xor U21381 (N_21381,N_18715,N_16969);
nand U21382 (N_21382,N_17120,N_15550);
nand U21383 (N_21383,N_17855,N_13956);
nor U21384 (N_21384,N_14968,N_13443);
xor U21385 (N_21385,N_17425,N_17279);
or U21386 (N_21386,N_12554,N_16270);
or U21387 (N_21387,N_18677,N_17408);
nor U21388 (N_21388,N_13221,N_16455);
or U21389 (N_21389,N_17342,N_17390);
nand U21390 (N_21390,N_18520,N_15133);
xnor U21391 (N_21391,N_17615,N_13590);
and U21392 (N_21392,N_12612,N_15411);
or U21393 (N_21393,N_17879,N_18413);
nor U21394 (N_21394,N_17427,N_18189);
nand U21395 (N_21395,N_18449,N_13362);
or U21396 (N_21396,N_13740,N_18484);
xnor U21397 (N_21397,N_12932,N_17953);
xor U21398 (N_21398,N_18422,N_15398);
xor U21399 (N_21399,N_16806,N_14203);
xor U21400 (N_21400,N_13743,N_15311);
xor U21401 (N_21401,N_12625,N_14530);
nand U21402 (N_21402,N_14586,N_13453);
and U21403 (N_21403,N_15708,N_18467);
and U21404 (N_21404,N_15712,N_18221);
nand U21405 (N_21405,N_16398,N_13187);
nand U21406 (N_21406,N_18133,N_18260);
nor U21407 (N_21407,N_13667,N_14686);
xor U21408 (N_21408,N_15427,N_14508);
nand U21409 (N_21409,N_13476,N_14103);
nor U21410 (N_21410,N_16486,N_14896);
xor U21411 (N_21411,N_13611,N_18676);
nor U21412 (N_21412,N_12671,N_16479);
and U21413 (N_21413,N_16790,N_14091);
xor U21414 (N_21414,N_14764,N_16784);
xor U21415 (N_21415,N_12514,N_16096);
nor U21416 (N_21416,N_18152,N_17062);
or U21417 (N_21417,N_16447,N_16552);
xor U21418 (N_21418,N_13063,N_17391);
nand U21419 (N_21419,N_13419,N_13635);
nand U21420 (N_21420,N_15184,N_12547);
and U21421 (N_21421,N_18322,N_13701);
and U21422 (N_21422,N_13609,N_16688);
or U21423 (N_21423,N_16584,N_18312);
and U21424 (N_21424,N_16561,N_18480);
and U21425 (N_21425,N_16647,N_15315);
xor U21426 (N_21426,N_18114,N_17424);
nand U21427 (N_21427,N_13749,N_14240);
nand U21428 (N_21428,N_18455,N_17103);
and U21429 (N_21429,N_13113,N_17875);
xnor U21430 (N_21430,N_13928,N_16855);
nand U21431 (N_21431,N_18296,N_14652);
and U21432 (N_21432,N_15094,N_14232);
and U21433 (N_21433,N_16197,N_12599);
nor U21434 (N_21434,N_14828,N_13284);
and U21435 (N_21435,N_17569,N_15679);
xor U21436 (N_21436,N_18604,N_17926);
and U21437 (N_21437,N_14840,N_17225);
or U21438 (N_21438,N_15210,N_14691);
and U21439 (N_21439,N_17008,N_15401);
nor U21440 (N_21440,N_15962,N_15070);
nor U21441 (N_21441,N_18614,N_14072);
nand U21442 (N_21442,N_13285,N_13251);
xor U21443 (N_21443,N_16822,N_15136);
nor U21444 (N_21444,N_18264,N_12739);
and U21445 (N_21445,N_17883,N_16009);
nand U21446 (N_21446,N_16558,N_18587);
nor U21447 (N_21447,N_15483,N_14772);
nor U21448 (N_21448,N_15231,N_17728);
nor U21449 (N_21449,N_18191,N_16789);
xnor U21450 (N_21450,N_16606,N_15166);
or U21451 (N_21451,N_17468,N_18530);
xnor U21452 (N_21452,N_14121,N_17350);
nor U21453 (N_21453,N_15938,N_16812);
nand U21454 (N_21454,N_17917,N_14534);
xor U21455 (N_21455,N_18294,N_16805);
or U21456 (N_21456,N_17432,N_15682);
nor U21457 (N_21457,N_16829,N_15249);
and U21458 (N_21458,N_18261,N_16797);
and U21459 (N_21459,N_14471,N_14037);
and U21460 (N_21460,N_18543,N_14568);
and U21461 (N_21461,N_17162,N_16276);
nor U21462 (N_21462,N_17756,N_14994);
and U21463 (N_21463,N_17237,N_13174);
nand U21464 (N_21464,N_18434,N_15193);
or U21465 (N_21465,N_15127,N_18291);
xor U21466 (N_21466,N_15930,N_16639);
xor U21467 (N_21467,N_15244,N_13577);
nand U21468 (N_21468,N_15882,N_18376);
nor U21469 (N_21469,N_17200,N_17553);
nor U21470 (N_21470,N_16440,N_15230);
xor U21471 (N_21471,N_12651,N_15588);
or U21472 (N_21472,N_17280,N_17394);
nand U21473 (N_21473,N_17976,N_18496);
nor U21474 (N_21474,N_13133,N_17073);
xor U21475 (N_21475,N_13493,N_16225);
nor U21476 (N_21476,N_15614,N_18489);
xor U21477 (N_21477,N_13441,N_17758);
nand U21478 (N_21478,N_13541,N_15525);
and U21479 (N_21479,N_16798,N_18462);
nor U21480 (N_21480,N_14362,N_18620);
nand U21481 (N_21481,N_15693,N_13950);
and U21482 (N_21482,N_18481,N_13566);
or U21483 (N_21483,N_13980,N_18518);
nand U21484 (N_21484,N_18008,N_16767);
nor U21485 (N_21485,N_15627,N_14548);
xor U21486 (N_21486,N_18097,N_18644);
nor U21487 (N_21487,N_14886,N_16113);
or U21488 (N_21488,N_13149,N_18703);
or U21489 (N_21489,N_14224,N_16612);
or U21490 (N_21490,N_16360,N_16030);
nand U21491 (N_21491,N_15670,N_13765);
or U21492 (N_21492,N_15056,N_16498);
xor U21493 (N_21493,N_13479,N_13055);
and U21494 (N_21494,N_15333,N_16857);
nor U21495 (N_21495,N_16845,N_15325);
or U21496 (N_21496,N_17295,N_16849);
xor U21497 (N_21497,N_16698,N_16090);
nor U21498 (N_21498,N_13216,N_17716);
xor U21499 (N_21499,N_13408,N_15085);
or U21500 (N_21500,N_13835,N_17897);
and U21501 (N_21501,N_16183,N_14385);
nor U21502 (N_21502,N_17032,N_16101);
nand U21503 (N_21503,N_12680,N_16527);
or U21504 (N_21504,N_16403,N_14130);
xor U21505 (N_21505,N_15025,N_14480);
nor U21506 (N_21506,N_17418,N_16868);
nor U21507 (N_21507,N_15000,N_15114);
nand U21508 (N_21508,N_17612,N_15276);
nor U21509 (N_21509,N_18373,N_16425);
nor U21510 (N_21510,N_16859,N_15553);
nand U21511 (N_21511,N_15578,N_15473);
and U21512 (N_21512,N_14584,N_12883);
xnor U21513 (N_21513,N_12505,N_18245);
xnor U21514 (N_21514,N_17259,N_15498);
nor U21515 (N_21515,N_14735,N_14870);
xor U21516 (N_21516,N_16313,N_12556);
nand U21517 (N_21517,N_14653,N_15886);
nor U21518 (N_21518,N_13054,N_15562);
xnor U21519 (N_21519,N_18181,N_17023);
xor U21520 (N_21520,N_12542,N_16114);
nor U21521 (N_21521,N_13056,N_14867);
or U21522 (N_21522,N_12634,N_14132);
nor U21523 (N_21523,N_14743,N_12789);
or U21524 (N_21524,N_15363,N_18224);
nand U21525 (N_21525,N_13014,N_14820);
or U21526 (N_21526,N_13090,N_14736);
nand U21527 (N_21527,N_15486,N_15775);
and U21528 (N_21528,N_16033,N_16081);
nor U21529 (N_21529,N_14827,N_14921);
xor U21530 (N_21530,N_16312,N_13893);
nand U21531 (N_21531,N_14183,N_13057);
nand U21532 (N_21532,N_16335,N_16654);
xnor U21533 (N_21533,N_13048,N_17066);
xnor U21534 (N_21534,N_18143,N_12935);
or U21535 (N_21535,N_17095,N_15942);
xor U21536 (N_21536,N_16265,N_15768);
nor U21537 (N_21537,N_14964,N_14079);
or U21538 (N_21538,N_13410,N_15989);
nand U21539 (N_21539,N_13562,N_14334);
nand U21540 (N_21540,N_14931,N_17904);
and U21541 (N_21541,N_16168,N_17634);
nor U21542 (N_21542,N_14422,N_17683);
or U21543 (N_21543,N_18653,N_14655);
nor U21544 (N_21544,N_17130,N_16399);
or U21545 (N_21545,N_13445,N_13756);
and U21546 (N_21546,N_14420,N_13999);
and U21547 (N_21547,N_14002,N_13976);
or U21548 (N_21548,N_14220,N_12750);
and U21549 (N_21549,N_16672,N_13130);
nand U21550 (N_21550,N_14498,N_14809);
xnor U21551 (N_21551,N_15597,N_12877);
nand U21552 (N_21552,N_12617,N_13181);
or U21553 (N_21553,N_17144,N_13484);
nand U21554 (N_21554,N_18228,N_16563);
nand U21555 (N_21555,N_16882,N_18638);
and U21556 (N_21556,N_17175,N_17137);
nor U21557 (N_21557,N_12665,N_16801);
nand U21558 (N_21558,N_17814,N_16932);
or U21559 (N_21559,N_18605,N_15687);
nor U21560 (N_21560,N_18235,N_15866);
and U21561 (N_21561,N_17817,N_18704);
xnor U21562 (N_21562,N_17822,N_15359);
and U21563 (N_21563,N_15790,N_16539);
and U21564 (N_21564,N_13142,N_16640);
xor U21565 (N_21565,N_17001,N_16973);
xor U21566 (N_21566,N_15699,N_13202);
xnor U21567 (N_21567,N_14759,N_17353);
or U21568 (N_21568,N_15451,N_17986);
nor U21569 (N_21569,N_15461,N_16079);
xnor U21570 (N_21570,N_16931,N_17470);
nor U21571 (N_21571,N_12528,N_13695);
nor U21572 (N_21572,N_16517,N_15570);
and U21573 (N_21573,N_12971,N_17101);
and U21574 (N_21574,N_16610,N_15358);
and U21575 (N_21575,N_13907,N_12833);
and U21576 (N_21576,N_15814,N_17654);
nor U21577 (N_21577,N_13354,N_14705);
nand U21578 (N_21578,N_17474,N_17889);
nor U21579 (N_21579,N_15208,N_16327);
nor U21580 (N_21580,N_14318,N_13265);
xor U21581 (N_21581,N_15054,N_16272);
nand U21582 (N_21582,N_18335,N_18735);
or U21583 (N_21583,N_13954,N_14859);
nor U21584 (N_21584,N_16741,N_13418);
nand U21585 (N_21585,N_16919,N_14310);
and U21586 (N_21586,N_18375,N_13746);
and U21587 (N_21587,N_18406,N_15445);
nor U21588 (N_21588,N_17898,N_16726);
nand U21589 (N_21589,N_18659,N_14467);
nor U21590 (N_21590,N_17277,N_16464);
nand U21591 (N_21591,N_18185,N_18318);
and U21592 (N_21592,N_12834,N_17981);
nand U21593 (N_21593,N_14719,N_13406);
and U21594 (N_21594,N_12927,N_18519);
xor U21595 (N_21595,N_15123,N_15919);
or U21596 (N_21596,N_13351,N_14582);
or U21597 (N_21597,N_16293,N_14071);
nor U21598 (N_21598,N_17731,N_14145);
xnor U21599 (N_21599,N_16566,N_14636);
and U21600 (N_21600,N_15971,N_17609);
or U21601 (N_21601,N_14746,N_17207);
or U21602 (N_21602,N_12859,N_15222);
xor U21603 (N_21603,N_15299,N_16380);
xnor U21604 (N_21604,N_15927,N_15939);
or U21605 (N_21605,N_17536,N_15548);
xnor U21606 (N_21606,N_13481,N_17224);
nor U21607 (N_21607,N_16653,N_15654);
nand U21608 (N_21608,N_15018,N_15178);
or U21609 (N_21609,N_13215,N_12943);
nor U21610 (N_21610,N_13704,N_17454);
nand U21611 (N_21611,N_14603,N_18733);
nand U21612 (N_21612,N_17373,N_17513);
nor U21613 (N_21613,N_17074,N_12991);
nor U21614 (N_21614,N_17426,N_18074);
or U21615 (N_21615,N_18324,N_15761);
xor U21616 (N_21616,N_17533,N_17014);
and U21617 (N_21617,N_16416,N_13926);
nand U21618 (N_21618,N_17457,N_16232);
nor U21619 (N_21619,N_16298,N_14194);
xnor U21620 (N_21620,N_14892,N_15826);
and U21621 (N_21621,N_13719,N_17043);
nand U21622 (N_21622,N_13830,N_15340);
nand U21623 (N_21623,N_14622,N_18459);
nor U21624 (N_21624,N_13906,N_15481);
nand U21625 (N_21625,N_16485,N_16334);
nor U21626 (N_21626,N_15724,N_13313);
and U21627 (N_21627,N_17652,N_13810);
xor U21628 (N_21628,N_17179,N_16389);
xor U21629 (N_21629,N_14808,N_13982);
nor U21630 (N_21630,N_14948,N_16533);
nor U21631 (N_21631,N_17766,N_16358);
and U21632 (N_21632,N_13898,N_15088);
and U21633 (N_21633,N_17504,N_15413);
or U21634 (N_21634,N_13001,N_18218);
nor U21635 (N_21635,N_13465,N_16001);
or U21636 (N_21636,N_16671,N_17732);
xnor U21637 (N_21637,N_16042,N_15503);
or U21638 (N_21638,N_14823,N_17241);
nor U21639 (N_21639,N_14265,N_14737);
or U21640 (N_21640,N_12697,N_13981);
or U21641 (N_21641,N_18436,N_16124);
nand U21642 (N_21642,N_18497,N_14259);
or U21643 (N_21643,N_18196,N_16964);
nor U21644 (N_21644,N_14115,N_16034);
and U21645 (N_21645,N_14126,N_14825);
and U21646 (N_21646,N_17269,N_18146);
nor U21647 (N_21647,N_18089,N_13472);
nand U21648 (N_21648,N_15233,N_18246);
xor U21649 (N_21649,N_13724,N_16435);
and U21650 (N_21650,N_14423,N_18517);
nor U21651 (N_21651,N_13829,N_13922);
xnor U21652 (N_21652,N_14513,N_16650);
nand U21653 (N_21653,N_13775,N_12912);
nor U21654 (N_21654,N_15819,N_17204);
nor U21655 (N_21655,N_16508,N_17215);
or U21656 (N_21656,N_12965,N_15460);
xor U21657 (N_21657,N_13885,N_14673);
nor U21658 (N_21658,N_14732,N_12990);
xnor U21659 (N_21659,N_16421,N_15097);
and U21660 (N_21660,N_15040,N_12809);
xor U21661 (N_21661,N_16562,N_13021);
xnor U21662 (N_21662,N_16937,N_16608);
and U21663 (N_21663,N_14355,N_16157);
nand U21664 (N_21664,N_16130,N_13745);
nand U21665 (N_21665,N_13972,N_15617);
or U21666 (N_21666,N_15255,N_14895);
xnor U21667 (N_21667,N_18639,N_13917);
or U21668 (N_21668,N_14164,N_12559);
nor U21669 (N_21669,N_12989,N_16711);
xnor U21670 (N_21670,N_16288,N_14486);
or U21671 (N_21671,N_14816,N_17087);
or U21672 (N_21672,N_16210,N_13334);
xor U21673 (N_21673,N_15559,N_14299);
nand U21674 (N_21674,N_16024,N_14263);
nor U21675 (N_21675,N_16466,N_18351);
nor U21676 (N_21676,N_13069,N_17518);
xor U21677 (N_21677,N_15669,N_17013);
nor U21678 (N_21678,N_14929,N_14026);
and U21679 (N_21679,N_15185,N_15993);
xor U21680 (N_21680,N_16108,N_15039);
nor U21681 (N_21681,N_14475,N_15256);
or U21682 (N_21682,N_16537,N_12745);
nand U21683 (N_21683,N_17956,N_18211);
xnor U21684 (N_21684,N_16154,N_13370);
and U21685 (N_21685,N_16011,N_15327);
nand U21686 (N_21686,N_13614,N_16821);
xnor U21687 (N_21687,N_14489,N_13025);
xnor U21688 (N_21688,N_14397,N_13074);
or U21689 (N_21689,N_18535,N_13374);
or U21690 (N_21690,N_17369,N_13570);
or U21691 (N_21691,N_17145,N_13567);
xnor U21692 (N_21692,N_17324,N_13292);
or U21693 (N_21693,N_13080,N_17745);
nand U21694 (N_21694,N_15915,N_18022);
or U21695 (N_21695,N_18565,N_17388);
or U21696 (N_21696,N_15431,N_18423);
and U21697 (N_21697,N_12512,N_15113);
nor U21698 (N_21698,N_18017,N_17148);
or U21699 (N_21699,N_13747,N_17517);
or U21700 (N_21700,N_14384,N_17543);
nand U21701 (N_21701,N_14125,N_12774);
and U21702 (N_21702,N_15087,N_17413);
xor U21703 (N_21703,N_18402,N_17443);
nand U21704 (N_21704,N_16984,N_14064);
xor U21705 (N_21705,N_15182,N_17482);
or U21706 (N_21706,N_14013,N_16593);
nand U21707 (N_21707,N_17184,N_16715);
and U21708 (N_21708,N_13425,N_17182);
or U21709 (N_21709,N_15983,N_18290);
nand U21710 (N_21710,N_16899,N_16427);
and U21711 (N_21711,N_14967,N_15433);
nand U21712 (N_21712,N_17105,N_12907);
xor U21713 (N_21713,N_16151,N_16116);
nor U21714 (N_21714,N_17827,N_17177);
nor U21715 (N_21715,N_14602,N_13977);
xor U21716 (N_21716,N_15134,N_14813);
and U21717 (N_21717,N_12801,N_16579);
or U21718 (N_21718,N_16739,N_18560);
and U21719 (N_21719,N_14923,N_13753);
nand U21720 (N_21720,N_16622,N_17455);
xnor U21721 (N_21721,N_17419,N_15705);
and U21722 (N_21722,N_15760,N_15728);
nor U21723 (N_21723,N_17909,N_18349);
xor U21724 (N_21724,N_15376,N_18723);
and U21725 (N_21725,N_12924,N_12842);
and U21726 (N_21726,N_18276,N_18595);
xor U21727 (N_21727,N_17928,N_16994);
nor U21728 (N_21728,N_16771,N_13654);
nand U21729 (N_21729,N_15308,N_16575);
nand U21730 (N_21730,N_14689,N_15541);
or U21731 (N_21731,N_14315,N_17874);
or U21732 (N_21732,N_15576,N_17938);
xnor U21733 (N_21733,N_18038,N_15645);
and U21734 (N_21734,N_12999,N_12839);
nor U21735 (N_21735,N_15300,N_17785);
and U21736 (N_21736,N_14345,N_14742);
or U21737 (N_21737,N_17386,N_15653);
nand U21738 (N_21738,N_13392,N_13521);
xor U21739 (N_21739,N_18409,N_17547);
and U21740 (N_21740,N_12800,N_15338);
nand U21741 (N_21741,N_17588,N_12517);
xor U21742 (N_21742,N_16199,N_15910);
or U21743 (N_21743,N_13531,N_18130);
xnor U21744 (N_21744,N_16807,N_16765);
and U21745 (N_21745,N_17264,N_13953);
and U21746 (N_21746,N_13838,N_13599);
nor U21747 (N_21747,N_18531,N_12740);
or U21748 (N_21748,N_14648,N_16613);
and U21749 (N_21749,N_14252,N_15512);
nand U21750 (N_21750,N_14537,N_13660);
and U21751 (N_21751,N_12909,N_15792);
xnor U21752 (N_21752,N_17006,N_13942);
and U21753 (N_21753,N_14402,N_12868);
nor U21754 (N_21754,N_17960,N_18106);
nand U21755 (N_21755,N_13720,N_14799);
nor U21756 (N_21756,N_18279,N_12870);
and U21757 (N_21757,N_18325,N_13053);
and U21758 (N_21758,N_13866,N_17009);
xor U21759 (N_21759,N_16341,N_14728);
nor U21760 (N_21760,N_15807,N_12545);
or U21761 (N_21761,N_15198,N_16308);
and U21762 (N_21762,N_16181,N_14783);
nor U21763 (N_21763,N_17417,N_15520);
nor U21764 (N_21764,N_13277,N_13395);
and U21765 (N_21765,N_17595,N_18741);
nor U21766 (N_21766,N_15574,N_13736);
nand U21767 (N_21767,N_16337,N_13238);
nand U21768 (N_21768,N_16972,N_15717);
xor U21769 (N_21769,N_14270,N_14687);
or U21770 (N_21770,N_16632,N_12536);
or U21771 (N_21771,N_16799,N_13059);
xor U21772 (N_21772,N_12573,N_12583);
nand U21773 (N_21773,N_17128,N_16162);
and U21774 (N_21774,N_12562,N_14396);
and U21775 (N_21775,N_18101,N_16939);
nor U21776 (N_21776,N_17004,N_17322);
and U21777 (N_21777,N_14416,N_16926);
xor U21778 (N_21778,N_15371,N_13860);
or U21779 (N_21779,N_17561,N_12890);
or U21780 (N_21780,N_17979,N_15580);
xnor U21781 (N_21781,N_17542,N_13793);
nor U21782 (N_21782,N_18506,N_15608);
and U21783 (N_21783,N_16203,N_14570);
or U21784 (N_21784,N_17044,N_13574);
nor U21785 (N_21785,N_14120,N_14882);
or U21786 (N_21786,N_16583,N_12954);
and U21787 (N_21787,N_15875,N_18509);
nor U21788 (N_21788,N_18579,N_16094);
nor U21789 (N_21789,N_14567,N_17640);
nor U21790 (N_21790,N_14429,N_16107);
or U21791 (N_21791,N_17888,N_16773);
or U21792 (N_21792,N_17932,N_17459);
nand U21793 (N_21793,N_15426,N_13546);
nand U21794 (N_21794,N_17311,N_13496);
nand U21795 (N_21795,N_13899,N_18338);
xor U21796 (N_21796,N_14626,N_13681);
and U21797 (N_21797,N_15489,N_15049);
nand U21798 (N_21798,N_15365,N_16603);
and U21799 (N_21799,N_13299,N_17922);
nor U21800 (N_21800,N_18165,N_15271);
and U21801 (N_21801,N_13624,N_13175);
or U21802 (N_21802,N_15098,N_15720);
and U21803 (N_21803,N_13051,N_17194);
and U21804 (N_21804,N_15225,N_16478);
or U21805 (N_21805,N_18446,N_13176);
nor U21806 (N_21806,N_15421,N_14117);
or U21807 (N_21807,N_12969,N_17690);
nor U21808 (N_21808,N_15013,N_16896);
and U21809 (N_21809,N_16325,N_15976);
nand U21810 (N_21810,N_17226,N_16663);
xor U21811 (N_21811,N_15749,N_16623);
or U21812 (N_21812,N_14615,N_17198);
xor U21813 (N_21813,N_12582,N_13099);
and U21814 (N_21814,N_17657,N_18241);
nor U21815 (N_21815,N_18552,N_17780);
or U21816 (N_21816,N_16228,N_14775);
nand U21817 (N_21817,N_13192,N_13464);
or U21818 (N_21818,N_15272,N_13680);
or U21819 (N_21819,N_16006,N_16873);
nand U21820 (N_21820,N_17625,N_16120);
nor U21821 (N_21821,N_16657,N_17138);
nor U21822 (N_21822,N_17805,N_13825);
xor U21823 (N_21823,N_14025,N_14523);
and U21824 (N_21824,N_12557,N_15420);
and U21825 (N_21825,N_14027,N_15022);
nor U21826 (N_21826,N_12738,N_14367);
nor U21827 (N_21827,N_15159,N_16544);
or U21828 (N_21828,N_14430,N_16700);
nor U21829 (N_21829,N_16458,N_16924);
xor U21830 (N_21830,N_17288,N_16459);
xor U21831 (N_21831,N_15283,N_18334);
or U21832 (N_21832,N_16910,N_13679);
nor U21833 (N_21833,N_15634,N_14289);
nor U21834 (N_21834,N_15392,N_16752);
nor U21835 (N_21835,N_16953,N_16600);
and U21836 (N_21836,N_14980,N_14861);
nand U21837 (N_21837,N_13625,N_18237);
and U21838 (N_21838,N_17299,N_17717);
xnor U21839 (N_21839,N_13623,N_18691);
nand U21840 (N_21840,N_13422,N_17714);
or U21841 (N_21841,N_14640,N_16645);
and U21842 (N_21842,N_17631,N_17121);
or U21843 (N_21843,N_14185,N_18342);
and U21844 (N_21844,N_16968,N_17799);
or U21845 (N_21845,N_13146,N_14917);
and U21846 (N_21846,N_17754,N_15239);
or U21847 (N_21847,N_17181,N_14649);
or U21848 (N_21848,N_13471,N_16588);
nand U21849 (N_21849,N_18508,N_13924);
and U21850 (N_21850,N_14311,N_14038);
or U21851 (N_21851,N_14393,N_16106);
nand U21852 (N_21852,N_15932,N_18633);
nand U21853 (N_21853,N_18454,N_16828);
nor U21854 (N_21854,N_15854,N_16961);
nor U21855 (N_21855,N_17047,N_15752);
nand U21856 (N_21856,N_16787,N_15755);
or U21857 (N_21857,N_17512,N_16965);
xor U21858 (N_21858,N_17867,N_17729);
nand U21859 (N_21859,N_15219,N_16620);
nor U21860 (N_21860,N_17070,N_17192);
or U21861 (N_21861,N_15964,N_15071);
nor U21862 (N_21862,N_14780,N_12845);
nor U21863 (N_21863,N_17603,N_16115);
or U21864 (N_21864,N_13060,N_14459);
and U21865 (N_21865,N_16702,N_18084);
nand U21866 (N_21866,N_13328,N_14341);
nor U21867 (N_21867,N_18394,N_16907);
nand U21868 (N_21868,N_12854,N_13139);
xor U21869 (N_21869,N_16693,N_17357);
nor U21870 (N_21870,N_14207,N_16652);
or U21871 (N_21871,N_17708,N_14526);
nand U21872 (N_21872,N_15495,N_14708);
nand U21873 (N_21873,N_12608,N_17699);
nand U21874 (N_21874,N_16138,N_12946);
nand U21875 (N_21875,N_18123,N_14489);
or U21876 (N_21876,N_16463,N_15819);
or U21877 (N_21877,N_14470,N_14832);
or U21878 (N_21878,N_13985,N_18646);
or U21879 (N_21879,N_14844,N_17956);
nor U21880 (N_21880,N_13909,N_13313);
or U21881 (N_21881,N_13309,N_15623);
and U21882 (N_21882,N_15228,N_17873);
nand U21883 (N_21883,N_18667,N_13442);
nor U21884 (N_21884,N_17639,N_16876);
xor U21885 (N_21885,N_17877,N_14479);
nand U21886 (N_21886,N_12660,N_14243);
nand U21887 (N_21887,N_16795,N_13240);
or U21888 (N_21888,N_18309,N_18523);
nor U21889 (N_21889,N_14488,N_16222);
xnor U21890 (N_21890,N_16448,N_18276);
or U21891 (N_21891,N_16958,N_13471);
nor U21892 (N_21892,N_16367,N_16294);
and U21893 (N_21893,N_18166,N_15863);
nor U21894 (N_21894,N_15294,N_14680);
nor U21895 (N_21895,N_13200,N_17375);
and U21896 (N_21896,N_18108,N_12793);
xnor U21897 (N_21897,N_14227,N_18067);
and U21898 (N_21898,N_18626,N_14819);
or U21899 (N_21899,N_17773,N_18240);
nand U21900 (N_21900,N_17472,N_15400);
and U21901 (N_21901,N_16818,N_15762);
xnor U21902 (N_21902,N_16430,N_13266);
or U21903 (N_21903,N_16207,N_18051);
nand U21904 (N_21904,N_14878,N_16983);
and U21905 (N_21905,N_13685,N_13728);
xnor U21906 (N_21906,N_13963,N_18728);
and U21907 (N_21907,N_17127,N_12612);
or U21908 (N_21908,N_13791,N_18359);
or U21909 (N_21909,N_14416,N_15499);
and U21910 (N_21910,N_15125,N_15257);
or U21911 (N_21911,N_17969,N_12772);
and U21912 (N_21912,N_12751,N_15177);
xor U21913 (N_21913,N_15152,N_14051);
or U21914 (N_21914,N_16248,N_13845);
nor U21915 (N_21915,N_13595,N_15394);
xnor U21916 (N_21916,N_17023,N_18030);
xnor U21917 (N_21917,N_16816,N_16073);
and U21918 (N_21918,N_15956,N_16446);
xor U21919 (N_21919,N_15040,N_13780);
nand U21920 (N_21920,N_18129,N_12580);
and U21921 (N_21921,N_13021,N_15512);
or U21922 (N_21922,N_16990,N_18241);
nor U21923 (N_21923,N_16135,N_12758);
and U21924 (N_21924,N_15543,N_13053);
and U21925 (N_21925,N_17505,N_17439);
nor U21926 (N_21926,N_17619,N_13340);
and U21927 (N_21927,N_13958,N_17362);
and U21928 (N_21928,N_18316,N_15391);
nand U21929 (N_21929,N_16883,N_14130);
or U21930 (N_21930,N_14545,N_15210);
or U21931 (N_21931,N_18251,N_17913);
or U21932 (N_21932,N_16351,N_15880);
xnor U21933 (N_21933,N_18531,N_12814);
and U21934 (N_21934,N_16565,N_16992);
nor U21935 (N_21935,N_16259,N_18181);
nor U21936 (N_21936,N_16529,N_14917);
and U21937 (N_21937,N_13551,N_13261);
nor U21938 (N_21938,N_13062,N_18185);
xnor U21939 (N_21939,N_18083,N_12744);
xor U21940 (N_21940,N_12738,N_16787);
xnor U21941 (N_21941,N_17842,N_17675);
xor U21942 (N_21942,N_12857,N_15654);
or U21943 (N_21943,N_13050,N_13476);
xor U21944 (N_21944,N_17283,N_16664);
nor U21945 (N_21945,N_12747,N_13095);
or U21946 (N_21946,N_16583,N_18480);
and U21947 (N_21947,N_16245,N_14827);
or U21948 (N_21948,N_16270,N_18573);
and U21949 (N_21949,N_15199,N_15026);
nor U21950 (N_21950,N_16131,N_15639);
nor U21951 (N_21951,N_14589,N_15164);
or U21952 (N_21952,N_15797,N_18147);
nand U21953 (N_21953,N_13868,N_13405);
nor U21954 (N_21954,N_13713,N_17655);
or U21955 (N_21955,N_16033,N_18099);
xor U21956 (N_21956,N_12851,N_16648);
and U21957 (N_21957,N_17574,N_14192);
or U21958 (N_21958,N_16684,N_12938);
or U21959 (N_21959,N_14834,N_17550);
nor U21960 (N_21960,N_16921,N_14058);
nand U21961 (N_21961,N_18158,N_18268);
nand U21962 (N_21962,N_18047,N_13993);
xor U21963 (N_21963,N_17073,N_14996);
nand U21964 (N_21964,N_17326,N_14387);
or U21965 (N_21965,N_16588,N_18157);
nand U21966 (N_21966,N_15714,N_16533);
nor U21967 (N_21967,N_18202,N_18710);
or U21968 (N_21968,N_14844,N_14021);
or U21969 (N_21969,N_17115,N_17551);
or U21970 (N_21970,N_16273,N_18319);
xor U21971 (N_21971,N_13103,N_17750);
and U21972 (N_21972,N_18229,N_16996);
and U21973 (N_21973,N_15493,N_14328);
xnor U21974 (N_21974,N_16219,N_13742);
nor U21975 (N_21975,N_14827,N_15134);
and U21976 (N_21976,N_16047,N_17177);
nor U21977 (N_21977,N_16040,N_15827);
or U21978 (N_21978,N_16415,N_13060);
or U21979 (N_21979,N_18367,N_18701);
nor U21980 (N_21980,N_13545,N_14854);
or U21981 (N_21981,N_14638,N_13426);
and U21982 (N_21982,N_15389,N_14605);
xnor U21983 (N_21983,N_15438,N_16454);
or U21984 (N_21984,N_15820,N_16612);
and U21985 (N_21985,N_16503,N_14664);
and U21986 (N_21986,N_15363,N_12764);
xor U21987 (N_21987,N_14233,N_17734);
nor U21988 (N_21988,N_12568,N_15752);
and U21989 (N_21989,N_15722,N_16919);
xnor U21990 (N_21990,N_16852,N_14166);
nor U21991 (N_21991,N_15536,N_17999);
xnor U21992 (N_21992,N_15515,N_13820);
nor U21993 (N_21993,N_17560,N_15396);
nand U21994 (N_21994,N_16704,N_16674);
and U21995 (N_21995,N_15315,N_17670);
and U21996 (N_21996,N_16617,N_12844);
and U21997 (N_21997,N_12697,N_14514);
and U21998 (N_21998,N_14885,N_13088);
nor U21999 (N_21999,N_14563,N_14965);
nand U22000 (N_22000,N_18065,N_16974);
and U22001 (N_22001,N_15369,N_13147);
and U22002 (N_22002,N_15218,N_12905);
nand U22003 (N_22003,N_16736,N_17177);
nand U22004 (N_22004,N_16243,N_16370);
nor U22005 (N_22005,N_18560,N_13103);
or U22006 (N_22006,N_14047,N_12575);
nand U22007 (N_22007,N_18685,N_14903);
or U22008 (N_22008,N_17066,N_16442);
nand U22009 (N_22009,N_16302,N_13330);
xor U22010 (N_22010,N_13958,N_17306);
nor U22011 (N_22011,N_17758,N_15604);
nor U22012 (N_22012,N_15061,N_15849);
nand U22013 (N_22013,N_12947,N_15040);
nand U22014 (N_22014,N_16324,N_17253);
and U22015 (N_22015,N_17596,N_17099);
xnor U22016 (N_22016,N_13640,N_13594);
and U22017 (N_22017,N_15089,N_13194);
or U22018 (N_22018,N_18467,N_13504);
nor U22019 (N_22019,N_17713,N_14712);
xor U22020 (N_22020,N_13874,N_13458);
and U22021 (N_22021,N_13273,N_17787);
nand U22022 (N_22022,N_17524,N_17585);
or U22023 (N_22023,N_18188,N_13103);
xnor U22024 (N_22024,N_12772,N_17232);
nand U22025 (N_22025,N_14638,N_14186);
xor U22026 (N_22026,N_14383,N_14096);
and U22027 (N_22027,N_14175,N_15632);
xor U22028 (N_22028,N_14752,N_14284);
nor U22029 (N_22029,N_15925,N_13270);
and U22030 (N_22030,N_13076,N_18038);
xor U22031 (N_22031,N_15847,N_13635);
nor U22032 (N_22032,N_17990,N_17207);
and U22033 (N_22033,N_15559,N_13444);
nand U22034 (N_22034,N_12996,N_16150);
and U22035 (N_22035,N_18634,N_14353);
xnor U22036 (N_22036,N_13863,N_18076);
nor U22037 (N_22037,N_17009,N_17554);
nand U22038 (N_22038,N_12944,N_16017);
nand U22039 (N_22039,N_17581,N_14336);
nor U22040 (N_22040,N_14444,N_14126);
xor U22041 (N_22041,N_14351,N_13895);
xnor U22042 (N_22042,N_13796,N_14275);
xnor U22043 (N_22043,N_15862,N_17638);
xor U22044 (N_22044,N_15896,N_12629);
and U22045 (N_22045,N_16171,N_14289);
nand U22046 (N_22046,N_15485,N_12707);
nor U22047 (N_22047,N_14799,N_18327);
nor U22048 (N_22048,N_15824,N_14524);
or U22049 (N_22049,N_14962,N_16236);
nand U22050 (N_22050,N_16490,N_13238);
nand U22051 (N_22051,N_13927,N_13193);
nand U22052 (N_22052,N_13628,N_17802);
xor U22053 (N_22053,N_16369,N_16598);
nand U22054 (N_22054,N_15904,N_17514);
nand U22055 (N_22055,N_12957,N_14097);
nand U22056 (N_22056,N_17635,N_17444);
nand U22057 (N_22057,N_18229,N_17448);
nand U22058 (N_22058,N_17315,N_17719);
nand U22059 (N_22059,N_15204,N_15382);
xnor U22060 (N_22060,N_13590,N_14800);
or U22061 (N_22061,N_18112,N_18513);
or U22062 (N_22062,N_17393,N_17026);
xor U22063 (N_22063,N_16519,N_13607);
nor U22064 (N_22064,N_18237,N_17996);
or U22065 (N_22065,N_17248,N_15277);
or U22066 (N_22066,N_13672,N_14343);
nand U22067 (N_22067,N_18326,N_18291);
nor U22068 (N_22068,N_13603,N_13487);
xnor U22069 (N_22069,N_13293,N_14028);
nor U22070 (N_22070,N_17449,N_14386);
nand U22071 (N_22071,N_13678,N_16739);
nand U22072 (N_22072,N_16523,N_17494);
xor U22073 (N_22073,N_14530,N_14051);
xnor U22074 (N_22074,N_13748,N_16654);
nand U22075 (N_22075,N_13019,N_12718);
and U22076 (N_22076,N_18637,N_15673);
nor U22077 (N_22077,N_15163,N_18426);
or U22078 (N_22078,N_17744,N_17164);
nand U22079 (N_22079,N_14226,N_13098);
or U22080 (N_22080,N_16800,N_18656);
nand U22081 (N_22081,N_17249,N_14231);
nor U22082 (N_22082,N_18437,N_14477);
or U22083 (N_22083,N_18013,N_15480);
nand U22084 (N_22084,N_18624,N_14612);
and U22085 (N_22085,N_14247,N_18274);
nand U22086 (N_22086,N_18176,N_13428);
nand U22087 (N_22087,N_16339,N_16234);
xor U22088 (N_22088,N_15993,N_16906);
or U22089 (N_22089,N_15343,N_14374);
nand U22090 (N_22090,N_17911,N_12897);
nand U22091 (N_22091,N_17246,N_17942);
nor U22092 (N_22092,N_13295,N_16124);
nand U22093 (N_22093,N_16981,N_13953);
nand U22094 (N_22094,N_17284,N_15587);
xnor U22095 (N_22095,N_17345,N_17681);
and U22096 (N_22096,N_14448,N_15727);
nand U22097 (N_22097,N_14996,N_14282);
and U22098 (N_22098,N_14102,N_15667);
nand U22099 (N_22099,N_17000,N_15629);
nand U22100 (N_22100,N_12801,N_12994);
or U22101 (N_22101,N_18276,N_13590);
and U22102 (N_22102,N_18517,N_16991);
nand U22103 (N_22103,N_16876,N_14878);
nor U22104 (N_22104,N_15114,N_17425);
nor U22105 (N_22105,N_18205,N_14089);
nor U22106 (N_22106,N_14385,N_15774);
xor U22107 (N_22107,N_15910,N_17379);
or U22108 (N_22108,N_15687,N_18029);
nor U22109 (N_22109,N_18420,N_15170);
xor U22110 (N_22110,N_15027,N_16979);
xnor U22111 (N_22111,N_18656,N_16721);
and U22112 (N_22112,N_18481,N_13820);
nor U22113 (N_22113,N_16907,N_15365);
and U22114 (N_22114,N_18250,N_18148);
xnor U22115 (N_22115,N_13775,N_17912);
or U22116 (N_22116,N_14052,N_12928);
nor U22117 (N_22117,N_17522,N_16686);
nor U22118 (N_22118,N_17035,N_15816);
and U22119 (N_22119,N_17559,N_13605);
and U22120 (N_22120,N_15655,N_12643);
xnor U22121 (N_22121,N_16272,N_12816);
xor U22122 (N_22122,N_16138,N_15787);
and U22123 (N_22123,N_16681,N_16633);
xnor U22124 (N_22124,N_12710,N_18380);
or U22125 (N_22125,N_13527,N_13837);
and U22126 (N_22126,N_13436,N_15294);
xor U22127 (N_22127,N_18313,N_13098);
nor U22128 (N_22128,N_13671,N_14087);
and U22129 (N_22129,N_17893,N_16625);
xnor U22130 (N_22130,N_16444,N_18743);
xor U22131 (N_22131,N_17352,N_12982);
nor U22132 (N_22132,N_18328,N_18320);
and U22133 (N_22133,N_17809,N_15713);
and U22134 (N_22134,N_15587,N_13310);
nand U22135 (N_22135,N_17953,N_17790);
nand U22136 (N_22136,N_16123,N_15949);
xnor U22137 (N_22137,N_13890,N_13590);
nand U22138 (N_22138,N_16887,N_18638);
or U22139 (N_22139,N_14161,N_18095);
or U22140 (N_22140,N_17099,N_17359);
or U22141 (N_22141,N_14292,N_18648);
or U22142 (N_22142,N_13838,N_17477);
xnor U22143 (N_22143,N_15985,N_18250);
nand U22144 (N_22144,N_15338,N_14885);
nand U22145 (N_22145,N_18690,N_14123);
or U22146 (N_22146,N_13457,N_15076);
or U22147 (N_22147,N_14282,N_15009);
xnor U22148 (N_22148,N_14582,N_17004);
nor U22149 (N_22149,N_12767,N_15503);
and U22150 (N_22150,N_18028,N_14715);
xnor U22151 (N_22151,N_12961,N_16620);
and U22152 (N_22152,N_15614,N_17471);
xor U22153 (N_22153,N_13014,N_12808);
nor U22154 (N_22154,N_14834,N_14771);
xor U22155 (N_22155,N_15375,N_13870);
or U22156 (N_22156,N_15719,N_18521);
nor U22157 (N_22157,N_15429,N_17500);
or U22158 (N_22158,N_14558,N_15324);
xnor U22159 (N_22159,N_16312,N_12661);
nand U22160 (N_22160,N_13581,N_16730);
nor U22161 (N_22161,N_17822,N_14874);
xor U22162 (N_22162,N_16601,N_14523);
and U22163 (N_22163,N_18543,N_18688);
or U22164 (N_22164,N_16073,N_14248);
and U22165 (N_22165,N_15797,N_13727);
nor U22166 (N_22166,N_18308,N_15236);
nor U22167 (N_22167,N_18022,N_13714);
nand U22168 (N_22168,N_13110,N_14060);
nor U22169 (N_22169,N_12658,N_13845);
and U22170 (N_22170,N_13688,N_16294);
nor U22171 (N_22171,N_12925,N_13504);
nor U22172 (N_22172,N_17866,N_13584);
nand U22173 (N_22173,N_17160,N_16110);
and U22174 (N_22174,N_14330,N_14194);
xnor U22175 (N_22175,N_13903,N_13262);
xor U22176 (N_22176,N_15947,N_18354);
xor U22177 (N_22177,N_15567,N_16051);
nand U22178 (N_22178,N_13453,N_15375);
xnor U22179 (N_22179,N_17426,N_12667);
or U22180 (N_22180,N_17010,N_13981);
nand U22181 (N_22181,N_18393,N_14635);
nand U22182 (N_22182,N_16700,N_12817);
nand U22183 (N_22183,N_16678,N_16116);
nand U22184 (N_22184,N_13860,N_15452);
or U22185 (N_22185,N_13235,N_16123);
nor U22186 (N_22186,N_14636,N_17792);
nor U22187 (N_22187,N_16354,N_17303);
nor U22188 (N_22188,N_16788,N_17692);
nand U22189 (N_22189,N_18546,N_15095);
or U22190 (N_22190,N_18030,N_14626);
xor U22191 (N_22191,N_17898,N_15193);
nand U22192 (N_22192,N_16652,N_13019);
nor U22193 (N_22193,N_16925,N_18007);
nor U22194 (N_22194,N_12775,N_14571);
nand U22195 (N_22195,N_13990,N_15442);
and U22196 (N_22196,N_16999,N_17287);
and U22197 (N_22197,N_17646,N_14667);
or U22198 (N_22198,N_12934,N_18251);
nand U22199 (N_22199,N_18386,N_15971);
nand U22200 (N_22200,N_15546,N_13027);
xor U22201 (N_22201,N_17003,N_15745);
nand U22202 (N_22202,N_15357,N_15588);
nand U22203 (N_22203,N_16381,N_14568);
or U22204 (N_22204,N_16014,N_16336);
xor U22205 (N_22205,N_13586,N_16374);
xnor U22206 (N_22206,N_17185,N_16796);
nand U22207 (N_22207,N_14680,N_15693);
nor U22208 (N_22208,N_12746,N_18519);
and U22209 (N_22209,N_15520,N_14396);
xor U22210 (N_22210,N_14968,N_14977);
or U22211 (N_22211,N_13515,N_15179);
or U22212 (N_22212,N_15717,N_13224);
nor U22213 (N_22213,N_12823,N_16706);
and U22214 (N_22214,N_17035,N_16809);
nor U22215 (N_22215,N_17419,N_16504);
or U22216 (N_22216,N_17491,N_15354);
xor U22217 (N_22217,N_18489,N_15109);
and U22218 (N_22218,N_14703,N_18644);
xor U22219 (N_22219,N_16186,N_14955);
nand U22220 (N_22220,N_17386,N_14484);
nor U22221 (N_22221,N_15844,N_14213);
nand U22222 (N_22222,N_16595,N_13696);
xor U22223 (N_22223,N_14571,N_18710);
nor U22224 (N_22224,N_14063,N_15238);
nor U22225 (N_22225,N_15914,N_16900);
nand U22226 (N_22226,N_15104,N_14420);
nor U22227 (N_22227,N_14111,N_16809);
and U22228 (N_22228,N_14297,N_15587);
or U22229 (N_22229,N_15702,N_16562);
nor U22230 (N_22230,N_16294,N_14282);
or U22231 (N_22231,N_12696,N_17943);
and U22232 (N_22232,N_13248,N_17516);
nand U22233 (N_22233,N_14474,N_15235);
nand U22234 (N_22234,N_14905,N_16645);
xnor U22235 (N_22235,N_14446,N_16582);
or U22236 (N_22236,N_16903,N_13132);
nand U22237 (N_22237,N_14261,N_18274);
nand U22238 (N_22238,N_12526,N_18446);
nand U22239 (N_22239,N_16553,N_15417);
xor U22240 (N_22240,N_14665,N_15456);
or U22241 (N_22241,N_15258,N_17246);
nor U22242 (N_22242,N_13962,N_12816);
and U22243 (N_22243,N_12655,N_15077);
xor U22244 (N_22244,N_14342,N_13763);
and U22245 (N_22245,N_14642,N_18622);
nor U22246 (N_22246,N_18421,N_14599);
and U22247 (N_22247,N_13708,N_14771);
or U22248 (N_22248,N_18730,N_17595);
and U22249 (N_22249,N_14637,N_15160);
xnor U22250 (N_22250,N_17962,N_14802);
xnor U22251 (N_22251,N_13092,N_13999);
xnor U22252 (N_22252,N_15145,N_13665);
xnor U22253 (N_22253,N_15087,N_17054);
nor U22254 (N_22254,N_17547,N_17714);
nand U22255 (N_22255,N_13081,N_16414);
nor U22256 (N_22256,N_13189,N_12639);
xor U22257 (N_22257,N_16045,N_15643);
or U22258 (N_22258,N_15203,N_13089);
and U22259 (N_22259,N_15660,N_12502);
xor U22260 (N_22260,N_14013,N_14136);
nand U22261 (N_22261,N_13492,N_15173);
xnor U22262 (N_22262,N_17495,N_15602);
nor U22263 (N_22263,N_13631,N_13981);
and U22264 (N_22264,N_15113,N_16869);
xor U22265 (N_22265,N_15993,N_14997);
xnor U22266 (N_22266,N_12758,N_16506);
xnor U22267 (N_22267,N_14896,N_18082);
nor U22268 (N_22268,N_15474,N_15102);
xnor U22269 (N_22269,N_15743,N_16171);
xor U22270 (N_22270,N_15284,N_13589);
xnor U22271 (N_22271,N_17719,N_15877);
nand U22272 (N_22272,N_14822,N_14656);
nand U22273 (N_22273,N_15763,N_15686);
and U22274 (N_22274,N_14756,N_16935);
nor U22275 (N_22275,N_14080,N_13341);
or U22276 (N_22276,N_13658,N_16502);
nor U22277 (N_22277,N_17272,N_17893);
nor U22278 (N_22278,N_18447,N_14953);
or U22279 (N_22279,N_16632,N_12689);
nor U22280 (N_22280,N_15641,N_16755);
and U22281 (N_22281,N_15089,N_16899);
nand U22282 (N_22282,N_14545,N_14267);
xnor U22283 (N_22283,N_16033,N_18378);
or U22284 (N_22284,N_14518,N_16780);
xor U22285 (N_22285,N_18304,N_14477);
nor U22286 (N_22286,N_14917,N_17572);
nor U22287 (N_22287,N_13356,N_14828);
nand U22288 (N_22288,N_18311,N_17497);
and U22289 (N_22289,N_16165,N_15207);
nor U22290 (N_22290,N_18172,N_18372);
nor U22291 (N_22291,N_18349,N_14438);
and U22292 (N_22292,N_14949,N_17048);
nor U22293 (N_22293,N_18344,N_17816);
nor U22294 (N_22294,N_13259,N_16705);
nor U22295 (N_22295,N_14596,N_17526);
nand U22296 (N_22296,N_16341,N_18063);
xor U22297 (N_22297,N_18462,N_14930);
xnor U22298 (N_22298,N_13804,N_15684);
and U22299 (N_22299,N_16465,N_15323);
xor U22300 (N_22300,N_15592,N_13139);
nor U22301 (N_22301,N_17467,N_14427);
nand U22302 (N_22302,N_18651,N_16985);
nor U22303 (N_22303,N_18468,N_13796);
and U22304 (N_22304,N_16659,N_12660);
xor U22305 (N_22305,N_14140,N_16772);
xor U22306 (N_22306,N_16131,N_13208);
nand U22307 (N_22307,N_17271,N_13371);
nand U22308 (N_22308,N_16479,N_14405);
xor U22309 (N_22309,N_18302,N_14240);
xnor U22310 (N_22310,N_17284,N_13182);
and U22311 (N_22311,N_13212,N_17970);
or U22312 (N_22312,N_16417,N_18306);
nor U22313 (N_22313,N_12570,N_16581);
and U22314 (N_22314,N_18192,N_15843);
and U22315 (N_22315,N_12754,N_17909);
nand U22316 (N_22316,N_16452,N_13705);
nand U22317 (N_22317,N_13702,N_13998);
nor U22318 (N_22318,N_16290,N_12506);
nor U22319 (N_22319,N_17586,N_13997);
and U22320 (N_22320,N_16709,N_12612);
nor U22321 (N_22321,N_16252,N_15974);
nor U22322 (N_22322,N_13962,N_13512);
xor U22323 (N_22323,N_12777,N_14756);
or U22324 (N_22324,N_13257,N_15781);
nand U22325 (N_22325,N_16488,N_18178);
xor U22326 (N_22326,N_18044,N_13261);
nand U22327 (N_22327,N_16188,N_13640);
xor U22328 (N_22328,N_17714,N_15766);
or U22329 (N_22329,N_16828,N_12938);
and U22330 (N_22330,N_14713,N_14004);
nor U22331 (N_22331,N_12636,N_14625);
nand U22332 (N_22332,N_15524,N_16030);
nor U22333 (N_22333,N_15267,N_18634);
nand U22334 (N_22334,N_13926,N_12791);
or U22335 (N_22335,N_13856,N_17490);
or U22336 (N_22336,N_16357,N_16417);
and U22337 (N_22337,N_17390,N_14143);
and U22338 (N_22338,N_18300,N_15009);
nand U22339 (N_22339,N_17140,N_16241);
or U22340 (N_22340,N_16447,N_12986);
or U22341 (N_22341,N_13505,N_17712);
nor U22342 (N_22342,N_12621,N_17371);
xnor U22343 (N_22343,N_17616,N_18227);
and U22344 (N_22344,N_14861,N_15671);
or U22345 (N_22345,N_14144,N_17563);
xor U22346 (N_22346,N_13437,N_13823);
or U22347 (N_22347,N_18645,N_17073);
nor U22348 (N_22348,N_13911,N_17262);
and U22349 (N_22349,N_16479,N_13241);
and U22350 (N_22350,N_14907,N_16435);
and U22351 (N_22351,N_15334,N_14601);
xor U22352 (N_22352,N_14498,N_17013);
xnor U22353 (N_22353,N_15297,N_15349);
or U22354 (N_22354,N_14607,N_16540);
or U22355 (N_22355,N_18172,N_16158);
and U22356 (N_22356,N_18433,N_18460);
xor U22357 (N_22357,N_17725,N_17290);
xnor U22358 (N_22358,N_15529,N_15975);
xor U22359 (N_22359,N_17858,N_16221);
or U22360 (N_22360,N_17367,N_16910);
xor U22361 (N_22361,N_15232,N_14398);
or U22362 (N_22362,N_17772,N_14026);
xor U22363 (N_22363,N_12816,N_18603);
xnor U22364 (N_22364,N_15020,N_18437);
xor U22365 (N_22365,N_15722,N_15531);
or U22366 (N_22366,N_14000,N_15082);
nor U22367 (N_22367,N_16639,N_12519);
and U22368 (N_22368,N_15731,N_17706);
nand U22369 (N_22369,N_15998,N_16416);
or U22370 (N_22370,N_14270,N_17431);
nand U22371 (N_22371,N_12634,N_13104);
or U22372 (N_22372,N_15818,N_17162);
nand U22373 (N_22373,N_15660,N_16031);
nor U22374 (N_22374,N_17068,N_17952);
nor U22375 (N_22375,N_17742,N_16341);
or U22376 (N_22376,N_14789,N_18212);
xor U22377 (N_22377,N_14596,N_17594);
nand U22378 (N_22378,N_13289,N_12511);
xnor U22379 (N_22379,N_17198,N_15838);
xnor U22380 (N_22380,N_18429,N_17079);
nor U22381 (N_22381,N_17938,N_18731);
nand U22382 (N_22382,N_18385,N_15000);
nor U22383 (N_22383,N_18062,N_13851);
or U22384 (N_22384,N_18286,N_14043);
nand U22385 (N_22385,N_18720,N_17804);
nand U22386 (N_22386,N_14202,N_17113);
and U22387 (N_22387,N_13948,N_17997);
or U22388 (N_22388,N_17805,N_14684);
xor U22389 (N_22389,N_13751,N_15053);
or U22390 (N_22390,N_13177,N_17039);
nor U22391 (N_22391,N_18637,N_17310);
nor U22392 (N_22392,N_12970,N_15389);
nand U22393 (N_22393,N_12650,N_15515);
nor U22394 (N_22394,N_18621,N_15003);
and U22395 (N_22395,N_17814,N_17145);
and U22396 (N_22396,N_14012,N_17918);
or U22397 (N_22397,N_18570,N_15479);
or U22398 (N_22398,N_17689,N_15801);
nor U22399 (N_22399,N_13616,N_18134);
xnor U22400 (N_22400,N_15166,N_18155);
or U22401 (N_22401,N_13369,N_12772);
nand U22402 (N_22402,N_14496,N_18384);
nor U22403 (N_22403,N_13642,N_14398);
xor U22404 (N_22404,N_17550,N_17758);
xnor U22405 (N_22405,N_13484,N_16641);
nor U22406 (N_22406,N_12724,N_14924);
nor U22407 (N_22407,N_13036,N_16679);
and U22408 (N_22408,N_16106,N_16388);
nor U22409 (N_22409,N_17853,N_12795);
xor U22410 (N_22410,N_12783,N_14460);
nor U22411 (N_22411,N_16649,N_18203);
xor U22412 (N_22412,N_13795,N_17271);
xor U22413 (N_22413,N_15821,N_17556);
nor U22414 (N_22414,N_18601,N_14858);
xor U22415 (N_22415,N_16816,N_17001);
xnor U22416 (N_22416,N_17545,N_14272);
xnor U22417 (N_22417,N_12760,N_13191);
nor U22418 (N_22418,N_14795,N_16817);
or U22419 (N_22419,N_17361,N_14447);
xor U22420 (N_22420,N_14216,N_17394);
xor U22421 (N_22421,N_17175,N_13896);
nand U22422 (N_22422,N_12868,N_17768);
and U22423 (N_22423,N_14153,N_12791);
nand U22424 (N_22424,N_13482,N_18735);
xor U22425 (N_22425,N_17967,N_13455);
xor U22426 (N_22426,N_15410,N_15475);
or U22427 (N_22427,N_18322,N_16886);
nor U22428 (N_22428,N_18095,N_16980);
and U22429 (N_22429,N_15813,N_13353);
and U22430 (N_22430,N_15389,N_14464);
and U22431 (N_22431,N_17024,N_13368);
xor U22432 (N_22432,N_14446,N_15296);
nand U22433 (N_22433,N_17476,N_14825);
and U22434 (N_22434,N_15392,N_12585);
nor U22435 (N_22435,N_18242,N_18241);
nor U22436 (N_22436,N_15273,N_18591);
nor U22437 (N_22437,N_18034,N_13951);
nand U22438 (N_22438,N_13371,N_15150);
nor U22439 (N_22439,N_15102,N_17437);
and U22440 (N_22440,N_15181,N_14742);
and U22441 (N_22441,N_13890,N_18098);
or U22442 (N_22442,N_17840,N_16723);
or U22443 (N_22443,N_17773,N_12686);
nor U22444 (N_22444,N_15046,N_15294);
or U22445 (N_22445,N_18481,N_13505);
and U22446 (N_22446,N_16067,N_14313);
or U22447 (N_22447,N_17947,N_17785);
nor U22448 (N_22448,N_17242,N_13900);
xnor U22449 (N_22449,N_15796,N_15610);
and U22450 (N_22450,N_16132,N_17846);
and U22451 (N_22451,N_15201,N_16408);
xor U22452 (N_22452,N_14062,N_13348);
nand U22453 (N_22453,N_12787,N_13171);
nand U22454 (N_22454,N_17491,N_18116);
xor U22455 (N_22455,N_16228,N_18461);
nand U22456 (N_22456,N_17819,N_17504);
nor U22457 (N_22457,N_17709,N_13462);
xor U22458 (N_22458,N_16802,N_17598);
or U22459 (N_22459,N_15483,N_16292);
or U22460 (N_22460,N_14299,N_18061);
or U22461 (N_22461,N_16556,N_15473);
xnor U22462 (N_22462,N_16623,N_18695);
nor U22463 (N_22463,N_13141,N_17144);
xor U22464 (N_22464,N_18508,N_16133);
and U22465 (N_22465,N_18626,N_15820);
nand U22466 (N_22466,N_12703,N_15977);
nor U22467 (N_22467,N_15051,N_14602);
nand U22468 (N_22468,N_13715,N_16429);
nor U22469 (N_22469,N_16712,N_14416);
nor U22470 (N_22470,N_13498,N_12883);
nand U22471 (N_22471,N_17613,N_13411);
or U22472 (N_22472,N_15850,N_17194);
and U22473 (N_22473,N_14083,N_18671);
nand U22474 (N_22474,N_17356,N_13395);
nand U22475 (N_22475,N_14025,N_15336);
nor U22476 (N_22476,N_16866,N_17756);
xor U22477 (N_22477,N_17264,N_14127);
or U22478 (N_22478,N_17952,N_15515);
or U22479 (N_22479,N_13175,N_17672);
nand U22480 (N_22480,N_14754,N_13027);
and U22481 (N_22481,N_17087,N_17197);
nor U22482 (N_22482,N_14252,N_14428);
and U22483 (N_22483,N_15022,N_12609);
and U22484 (N_22484,N_14410,N_16911);
or U22485 (N_22485,N_17287,N_13947);
xnor U22486 (N_22486,N_15287,N_12669);
nand U22487 (N_22487,N_13106,N_16981);
xor U22488 (N_22488,N_13859,N_16701);
xnor U22489 (N_22489,N_16526,N_17177);
nand U22490 (N_22490,N_16890,N_13158);
nand U22491 (N_22491,N_16279,N_13722);
nand U22492 (N_22492,N_16450,N_15622);
nand U22493 (N_22493,N_13392,N_15379);
nor U22494 (N_22494,N_15405,N_15036);
or U22495 (N_22495,N_13074,N_14141);
or U22496 (N_22496,N_16207,N_14211);
nor U22497 (N_22497,N_12569,N_18092);
nor U22498 (N_22498,N_12583,N_13866);
and U22499 (N_22499,N_18371,N_18161);
and U22500 (N_22500,N_17058,N_14952);
xor U22501 (N_22501,N_16784,N_17832);
nand U22502 (N_22502,N_18743,N_15212);
and U22503 (N_22503,N_16358,N_12750);
xor U22504 (N_22504,N_18204,N_16664);
nor U22505 (N_22505,N_14407,N_15634);
xor U22506 (N_22506,N_13307,N_13925);
and U22507 (N_22507,N_13385,N_17766);
xnor U22508 (N_22508,N_13465,N_13379);
and U22509 (N_22509,N_16851,N_15106);
or U22510 (N_22510,N_16405,N_16946);
xor U22511 (N_22511,N_14256,N_18629);
nor U22512 (N_22512,N_13689,N_13680);
or U22513 (N_22513,N_14164,N_17155);
nand U22514 (N_22514,N_13335,N_17943);
xnor U22515 (N_22515,N_17917,N_12742);
and U22516 (N_22516,N_13902,N_15027);
xnor U22517 (N_22517,N_15054,N_15137);
xnor U22518 (N_22518,N_15206,N_18633);
and U22519 (N_22519,N_14550,N_17784);
or U22520 (N_22520,N_13182,N_16006);
nor U22521 (N_22521,N_15578,N_17024);
or U22522 (N_22522,N_15292,N_13637);
nand U22523 (N_22523,N_15008,N_12740);
nor U22524 (N_22524,N_18158,N_17349);
and U22525 (N_22525,N_14596,N_12948);
xor U22526 (N_22526,N_13018,N_17804);
and U22527 (N_22527,N_17560,N_13814);
and U22528 (N_22528,N_18476,N_15803);
or U22529 (N_22529,N_15015,N_13581);
nand U22530 (N_22530,N_17290,N_17229);
and U22531 (N_22531,N_18354,N_17081);
or U22532 (N_22532,N_17671,N_18013);
nor U22533 (N_22533,N_13156,N_12842);
or U22534 (N_22534,N_15103,N_18350);
or U22535 (N_22535,N_12723,N_13816);
nand U22536 (N_22536,N_14549,N_18723);
nor U22537 (N_22537,N_14550,N_13174);
or U22538 (N_22538,N_14980,N_17045);
xor U22539 (N_22539,N_15416,N_14907);
and U22540 (N_22540,N_17210,N_12847);
nand U22541 (N_22541,N_16727,N_17930);
xor U22542 (N_22542,N_16406,N_18583);
nor U22543 (N_22543,N_17124,N_13611);
nor U22544 (N_22544,N_15959,N_14093);
or U22545 (N_22545,N_18021,N_13264);
nand U22546 (N_22546,N_15640,N_18406);
and U22547 (N_22547,N_16160,N_18712);
xnor U22548 (N_22548,N_15581,N_16636);
xor U22549 (N_22549,N_18217,N_13756);
or U22550 (N_22550,N_15467,N_18309);
xnor U22551 (N_22551,N_16844,N_18748);
nand U22552 (N_22552,N_16982,N_15565);
xor U22553 (N_22553,N_12647,N_13107);
and U22554 (N_22554,N_13932,N_17995);
and U22555 (N_22555,N_13913,N_15710);
xnor U22556 (N_22556,N_15710,N_15001);
xnor U22557 (N_22557,N_17927,N_14298);
or U22558 (N_22558,N_14347,N_18156);
or U22559 (N_22559,N_13217,N_13562);
and U22560 (N_22560,N_15048,N_17392);
or U22561 (N_22561,N_12621,N_14244);
xor U22562 (N_22562,N_17741,N_12829);
nand U22563 (N_22563,N_15014,N_17317);
nor U22564 (N_22564,N_18168,N_13591);
and U22565 (N_22565,N_16165,N_13346);
nand U22566 (N_22566,N_16756,N_16250);
or U22567 (N_22567,N_18074,N_13186);
or U22568 (N_22568,N_14428,N_15144);
xor U22569 (N_22569,N_18518,N_14167);
nand U22570 (N_22570,N_12828,N_13573);
nand U22571 (N_22571,N_13072,N_17331);
xnor U22572 (N_22572,N_14101,N_15697);
and U22573 (N_22573,N_14146,N_14314);
or U22574 (N_22574,N_16779,N_16607);
or U22575 (N_22575,N_18076,N_17086);
xnor U22576 (N_22576,N_12970,N_12651);
xor U22577 (N_22577,N_15485,N_14852);
nand U22578 (N_22578,N_13797,N_17700);
nand U22579 (N_22579,N_13315,N_13090);
xnor U22580 (N_22580,N_15434,N_18194);
and U22581 (N_22581,N_14170,N_12965);
and U22582 (N_22582,N_16222,N_12882);
nor U22583 (N_22583,N_18118,N_16927);
or U22584 (N_22584,N_14548,N_14383);
nor U22585 (N_22585,N_17351,N_18526);
and U22586 (N_22586,N_16109,N_14750);
nor U22587 (N_22587,N_17255,N_14226);
nor U22588 (N_22588,N_13666,N_16925);
nor U22589 (N_22589,N_14201,N_13291);
and U22590 (N_22590,N_12526,N_18357);
nand U22591 (N_22591,N_15371,N_13579);
or U22592 (N_22592,N_16723,N_15148);
or U22593 (N_22593,N_15219,N_12749);
xnor U22594 (N_22594,N_14516,N_16130);
xor U22595 (N_22595,N_13826,N_17952);
nand U22596 (N_22596,N_12823,N_12592);
or U22597 (N_22597,N_12756,N_16581);
xor U22598 (N_22598,N_18240,N_16806);
nand U22599 (N_22599,N_13890,N_12939);
or U22600 (N_22600,N_15839,N_17422);
and U22601 (N_22601,N_14810,N_14650);
xor U22602 (N_22602,N_12920,N_13532);
or U22603 (N_22603,N_17380,N_13996);
and U22604 (N_22604,N_15524,N_17170);
nand U22605 (N_22605,N_18194,N_14084);
and U22606 (N_22606,N_15184,N_18277);
or U22607 (N_22607,N_16417,N_13448);
and U22608 (N_22608,N_13310,N_15946);
or U22609 (N_22609,N_16235,N_16830);
and U22610 (N_22610,N_17330,N_15115);
nor U22611 (N_22611,N_13576,N_15134);
xor U22612 (N_22612,N_16755,N_13507);
or U22613 (N_22613,N_12880,N_17235);
or U22614 (N_22614,N_16383,N_15290);
nor U22615 (N_22615,N_13415,N_16191);
nand U22616 (N_22616,N_18411,N_14670);
nor U22617 (N_22617,N_17271,N_13049);
or U22618 (N_22618,N_17064,N_15125);
xor U22619 (N_22619,N_13332,N_16637);
or U22620 (N_22620,N_12738,N_18283);
or U22621 (N_22621,N_17453,N_12832);
nor U22622 (N_22622,N_13400,N_16189);
nand U22623 (N_22623,N_17200,N_18165);
or U22624 (N_22624,N_16170,N_18558);
and U22625 (N_22625,N_15995,N_17509);
and U22626 (N_22626,N_14067,N_15684);
or U22627 (N_22627,N_13505,N_16894);
nand U22628 (N_22628,N_18597,N_13488);
xnor U22629 (N_22629,N_15810,N_17470);
nand U22630 (N_22630,N_18439,N_12563);
nand U22631 (N_22631,N_13375,N_18058);
and U22632 (N_22632,N_15238,N_17123);
or U22633 (N_22633,N_18113,N_17886);
xnor U22634 (N_22634,N_18449,N_18290);
and U22635 (N_22635,N_12622,N_14669);
nor U22636 (N_22636,N_13176,N_14573);
nand U22637 (N_22637,N_15715,N_14789);
or U22638 (N_22638,N_18682,N_16300);
nor U22639 (N_22639,N_16201,N_15047);
or U22640 (N_22640,N_17739,N_18739);
nor U22641 (N_22641,N_13568,N_15468);
nor U22642 (N_22642,N_17214,N_14999);
or U22643 (N_22643,N_13498,N_16480);
nand U22644 (N_22644,N_14792,N_14024);
nor U22645 (N_22645,N_15047,N_18617);
or U22646 (N_22646,N_15645,N_18706);
nand U22647 (N_22647,N_15869,N_12516);
or U22648 (N_22648,N_15775,N_17031);
nor U22649 (N_22649,N_17439,N_13525);
or U22650 (N_22650,N_13259,N_12804);
xor U22651 (N_22651,N_15665,N_13194);
nor U22652 (N_22652,N_17958,N_17561);
nand U22653 (N_22653,N_18729,N_17571);
nand U22654 (N_22654,N_12853,N_18092);
or U22655 (N_22655,N_17028,N_17954);
or U22656 (N_22656,N_13105,N_16408);
or U22657 (N_22657,N_16598,N_16783);
nor U22658 (N_22658,N_14519,N_16254);
and U22659 (N_22659,N_17609,N_18056);
xor U22660 (N_22660,N_16849,N_16731);
nand U22661 (N_22661,N_16719,N_14990);
xor U22662 (N_22662,N_18266,N_14374);
xnor U22663 (N_22663,N_14968,N_15513);
and U22664 (N_22664,N_16906,N_18110);
xor U22665 (N_22665,N_12752,N_15347);
and U22666 (N_22666,N_14009,N_14882);
nand U22667 (N_22667,N_15457,N_14125);
nand U22668 (N_22668,N_14942,N_16364);
nor U22669 (N_22669,N_16652,N_12874);
nor U22670 (N_22670,N_13981,N_16668);
or U22671 (N_22671,N_18450,N_18253);
xnor U22672 (N_22672,N_14779,N_16850);
or U22673 (N_22673,N_14312,N_16001);
xor U22674 (N_22674,N_17149,N_15189);
xor U22675 (N_22675,N_12671,N_15225);
nor U22676 (N_22676,N_16076,N_17174);
or U22677 (N_22677,N_17640,N_15932);
nor U22678 (N_22678,N_18108,N_12781);
nor U22679 (N_22679,N_14452,N_16529);
or U22680 (N_22680,N_13978,N_16072);
nand U22681 (N_22681,N_14649,N_18309);
nand U22682 (N_22682,N_17734,N_15929);
nor U22683 (N_22683,N_18418,N_15169);
or U22684 (N_22684,N_15716,N_18352);
and U22685 (N_22685,N_17964,N_17188);
or U22686 (N_22686,N_17732,N_16438);
nor U22687 (N_22687,N_16295,N_15395);
nor U22688 (N_22688,N_16384,N_16550);
nor U22689 (N_22689,N_14430,N_17835);
or U22690 (N_22690,N_17182,N_15739);
xnor U22691 (N_22691,N_14707,N_18707);
xnor U22692 (N_22692,N_14316,N_13019);
nor U22693 (N_22693,N_16000,N_15241);
xnor U22694 (N_22694,N_17804,N_17469);
and U22695 (N_22695,N_13487,N_14931);
nand U22696 (N_22696,N_14933,N_16307);
and U22697 (N_22697,N_13560,N_12977);
or U22698 (N_22698,N_16507,N_13928);
or U22699 (N_22699,N_14645,N_17350);
xor U22700 (N_22700,N_13060,N_17881);
nor U22701 (N_22701,N_14040,N_15239);
nand U22702 (N_22702,N_16580,N_17516);
or U22703 (N_22703,N_14511,N_17281);
nand U22704 (N_22704,N_17095,N_14194);
or U22705 (N_22705,N_16706,N_17170);
or U22706 (N_22706,N_14778,N_16617);
and U22707 (N_22707,N_16102,N_14482);
nor U22708 (N_22708,N_13451,N_13777);
or U22709 (N_22709,N_17366,N_17406);
nand U22710 (N_22710,N_16384,N_13482);
xor U22711 (N_22711,N_14870,N_15144);
or U22712 (N_22712,N_15804,N_16492);
and U22713 (N_22713,N_15530,N_18398);
nor U22714 (N_22714,N_14777,N_18704);
or U22715 (N_22715,N_16640,N_16303);
nand U22716 (N_22716,N_16058,N_17733);
and U22717 (N_22717,N_17395,N_14740);
nor U22718 (N_22718,N_16129,N_17387);
nor U22719 (N_22719,N_12888,N_12765);
nor U22720 (N_22720,N_14414,N_16279);
xnor U22721 (N_22721,N_18730,N_17275);
or U22722 (N_22722,N_15470,N_18186);
or U22723 (N_22723,N_17672,N_14674);
nor U22724 (N_22724,N_17064,N_16409);
xor U22725 (N_22725,N_13172,N_12783);
xor U22726 (N_22726,N_17455,N_17610);
nor U22727 (N_22727,N_17836,N_14812);
or U22728 (N_22728,N_13883,N_12903);
and U22729 (N_22729,N_14734,N_13241);
xnor U22730 (N_22730,N_16015,N_16883);
and U22731 (N_22731,N_16116,N_12602);
nor U22732 (N_22732,N_15069,N_12737);
nor U22733 (N_22733,N_14465,N_14152);
and U22734 (N_22734,N_14607,N_17753);
and U22735 (N_22735,N_13139,N_13531);
nand U22736 (N_22736,N_14689,N_16271);
nor U22737 (N_22737,N_14290,N_14465);
and U22738 (N_22738,N_15141,N_15261);
or U22739 (N_22739,N_18662,N_12891);
or U22740 (N_22740,N_16137,N_15823);
or U22741 (N_22741,N_14238,N_18611);
and U22742 (N_22742,N_17448,N_18223);
nand U22743 (N_22743,N_15595,N_12706);
nor U22744 (N_22744,N_14996,N_14523);
nand U22745 (N_22745,N_15928,N_15031);
and U22746 (N_22746,N_12974,N_17751);
or U22747 (N_22747,N_17525,N_14375);
xor U22748 (N_22748,N_12573,N_17038);
nand U22749 (N_22749,N_16282,N_16909);
or U22750 (N_22750,N_13368,N_14539);
or U22751 (N_22751,N_15454,N_13679);
xnor U22752 (N_22752,N_14423,N_13366);
nor U22753 (N_22753,N_18653,N_14089);
nand U22754 (N_22754,N_15970,N_18376);
and U22755 (N_22755,N_14496,N_14624);
nand U22756 (N_22756,N_15913,N_12813);
or U22757 (N_22757,N_13955,N_15622);
or U22758 (N_22758,N_15050,N_15826);
or U22759 (N_22759,N_15317,N_12725);
or U22760 (N_22760,N_17742,N_15685);
xnor U22761 (N_22761,N_14827,N_17815);
and U22762 (N_22762,N_16417,N_14982);
or U22763 (N_22763,N_15977,N_13848);
nor U22764 (N_22764,N_13108,N_17921);
or U22765 (N_22765,N_18605,N_14514);
or U22766 (N_22766,N_14473,N_17697);
xor U22767 (N_22767,N_15878,N_15417);
xnor U22768 (N_22768,N_14666,N_17494);
and U22769 (N_22769,N_16180,N_16895);
nand U22770 (N_22770,N_13066,N_14072);
or U22771 (N_22771,N_17925,N_16082);
and U22772 (N_22772,N_17818,N_15100);
or U22773 (N_22773,N_14575,N_16318);
or U22774 (N_22774,N_17524,N_18312);
or U22775 (N_22775,N_14265,N_16172);
xnor U22776 (N_22776,N_17811,N_14375);
nor U22777 (N_22777,N_14816,N_13476);
nor U22778 (N_22778,N_14576,N_14150);
xnor U22779 (N_22779,N_15528,N_14616);
xnor U22780 (N_22780,N_13490,N_17213);
and U22781 (N_22781,N_18111,N_17819);
xor U22782 (N_22782,N_13980,N_13893);
or U22783 (N_22783,N_18108,N_15042);
nand U22784 (N_22784,N_15236,N_15143);
nor U22785 (N_22785,N_13772,N_17165);
or U22786 (N_22786,N_14936,N_15954);
and U22787 (N_22787,N_15787,N_13397);
xor U22788 (N_22788,N_15337,N_14552);
nor U22789 (N_22789,N_18246,N_17916);
nand U22790 (N_22790,N_14407,N_18194);
nor U22791 (N_22791,N_17436,N_14192);
xnor U22792 (N_22792,N_14467,N_18516);
or U22793 (N_22793,N_16670,N_16049);
and U22794 (N_22794,N_16376,N_14133);
nand U22795 (N_22795,N_15266,N_14149);
and U22796 (N_22796,N_18473,N_16343);
xnor U22797 (N_22797,N_17681,N_13419);
or U22798 (N_22798,N_15453,N_14930);
xor U22799 (N_22799,N_18600,N_17500);
nand U22800 (N_22800,N_16458,N_16303);
and U22801 (N_22801,N_13527,N_12921);
nor U22802 (N_22802,N_17356,N_14824);
or U22803 (N_22803,N_18330,N_15754);
xor U22804 (N_22804,N_17837,N_15269);
and U22805 (N_22805,N_13331,N_16729);
and U22806 (N_22806,N_15242,N_17781);
nor U22807 (N_22807,N_13955,N_15159);
and U22808 (N_22808,N_14401,N_17817);
or U22809 (N_22809,N_18161,N_16086);
and U22810 (N_22810,N_17430,N_16609);
or U22811 (N_22811,N_18659,N_18318);
or U22812 (N_22812,N_17395,N_14768);
or U22813 (N_22813,N_15362,N_14666);
or U22814 (N_22814,N_18211,N_14597);
xnor U22815 (N_22815,N_15809,N_15289);
and U22816 (N_22816,N_18420,N_14234);
and U22817 (N_22817,N_13636,N_18720);
or U22818 (N_22818,N_14999,N_14502);
or U22819 (N_22819,N_13547,N_16855);
nand U22820 (N_22820,N_17815,N_16193);
or U22821 (N_22821,N_16996,N_18532);
or U22822 (N_22822,N_14783,N_16192);
and U22823 (N_22823,N_12948,N_16939);
xnor U22824 (N_22824,N_14039,N_12621);
and U22825 (N_22825,N_13286,N_16295);
and U22826 (N_22826,N_17000,N_13532);
xnor U22827 (N_22827,N_18690,N_15689);
and U22828 (N_22828,N_14935,N_14161);
or U22829 (N_22829,N_17319,N_14286);
or U22830 (N_22830,N_17138,N_17283);
xnor U22831 (N_22831,N_14065,N_13902);
nand U22832 (N_22832,N_17059,N_13116);
nor U22833 (N_22833,N_15261,N_12693);
or U22834 (N_22834,N_14326,N_16280);
xor U22835 (N_22835,N_12579,N_14499);
nand U22836 (N_22836,N_18243,N_15291);
or U22837 (N_22837,N_14277,N_16853);
and U22838 (N_22838,N_15563,N_13829);
nor U22839 (N_22839,N_16985,N_18704);
xnor U22840 (N_22840,N_12575,N_17880);
nor U22841 (N_22841,N_17905,N_12827);
xnor U22842 (N_22842,N_14724,N_15036);
nor U22843 (N_22843,N_13980,N_18172);
and U22844 (N_22844,N_13045,N_13867);
nor U22845 (N_22845,N_17985,N_17123);
xor U22846 (N_22846,N_13720,N_13805);
and U22847 (N_22847,N_16974,N_12631);
and U22848 (N_22848,N_16392,N_16171);
or U22849 (N_22849,N_15994,N_13940);
nand U22850 (N_22850,N_16639,N_18453);
or U22851 (N_22851,N_13768,N_12655);
or U22852 (N_22852,N_12721,N_18143);
xor U22853 (N_22853,N_15966,N_15699);
nand U22854 (N_22854,N_17027,N_14303);
nand U22855 (N_22855,N_13086,N_14049);
nand U22856 (N_22856,N_18617,N_12650);
nand U22857 (N_22857,N_17422,N_15772);
or U22858 (N_22858,N_12947,N_16691);
xor U22859 (N_22859,N_17895,N_17940);
and U22860 (N_22860,N_17600,N_18062);
xnor U22861 (N_22861,N_17773,N_17483);
xnor U22862 (N_22862,N_13769,N_15117);
xnor U22863 (N_22863,N_14748,N_18743);
and U22864 (N_22864,N_17407,N_16372);
xnor U22865 (N_22865,N_16078,N_12943);
and U22866 (N_22866,N_17229,N_15323);
nand U22867 (N_22867,N_16939,N_13273);
nand U22868 (N_22868,N_12606,N_14216);
or U22869 (N_22869,N_18464,N_12867);
or U22870 (N_22870,N_12888,N_13187);
and U22871 (N_22871,N_17882,N_14718);
xnor U22872 (N_22872,N_18350,N_15647);
and U22873 (N_22873,N_16570,N_14900);
xor U22874 (N_22874,N_17640,N_13531);
or U22875 (N_22875,N_13077,N_15883);
or U22876 (N_22876,N_14164,N_14744);
and U22877 (N_22877,N_13843,N_13154);
xnor U22878 (N_22878,N_16738,N_12863);
xnor U22879 (N_22879,N_14143,N_16918);
or U22880 (N_22880,N_16655,N_15018);
xnor U22881 (N_22881,N_17068,N_14740);
nor U22882 (N_22882,N_16749,N_16747);
nor U22883 (N_22883,N_17200,N_16023);
nand U22884 (N_22884,N_14776,N_12647);
or U22885 (N_22885,N_17583,N_14070);
or U22886 (N_22886,N_17476,N_13707);
or U22887 (N_22887,N_13028,N_15938);
and U22888 (N_22888,N_15999,N_15916);
or U22889 (N_22889,N_18711,N_18399);
xnor U22890 (N_22890,N_15862,N_15760);
and U22891 (N_22891,N_15098,N_18553);
xnor U22892 (N_22892,N_17597,N_14628);
or U22893 (N_22893,N_16096,N_15796);
or U22894 (N_22894,N_13258,N_12834);
nor U22895 (N_22895,N_17860,N_18237);
nand U22896 (N_22896,N_16842,N_16951);
xor U22897 (N_22897,N_13567,N_14411);
nor U22898 (N_22898,N_14095,N_13923);
nor U22899 (N_22899,N_17110,N_14515);
xnor U22900 (N_22900,N_15497,N_17313);
nor U22901 (N_22901,N_17058,N_14983);
xor U22902 (N_22902,N_16309,N_16845);
nor U22903 (N_22903,N_18137,N_17224);
xor U22904 (N_22904,N_13242,N_14347);
nand U22905 (N_22905,N_14479,N_17511);
and U22906 (N_22906,N_13409,N_13572);
nand U22907 (N_22907,N_13414,N_17447);
and U22908 (N_22908,N_15727,N_18264);
nor U22909 (N_22909,N_18617,N_17973);
and U22910 (N_22910,N_16494,N_13099);
nand U22911 (N_22911,N_14990,N_18710);
and U22912 (N_22912,N_17781,N_15970);
nor U22913 (N_22913,N_18064,N_14702);
xor U22914 (N_22914,N_15738,N_18203);
nor U22915 (N_22915,N_14148,N_17487);
nor U22916 (N_22916,N_15591,N_14605);
nand U22917 (N_22917,N_15828,N_16119);
and U22918 (N_22918,N_16869,N_14674);
nand U22919 (N_22919,N_16079,N_17183);
nor U22920 (N_22920,N_16861,N_14336);
nand U22921 (N_22921,N_18651,N_13681);
and U22922 (N_22922,N_13716,N_14184);
nand U22923 (N_22923,N_15997,N_14928);
and U22924 (N_22924,N_16585,N_12944);
or U22925 (N_22925,N_16078,N_16042);
xnor U22926 (N_22926,N_14618,N_17489);
xnor U22927 (N_22927,N_15760,N_12830);
or U22928 (N_22928,N_13582,N_16217);
nor U22929 (N_22929,N_16636,N_18242);
xnor U22930 (N_22930,N_14162,N_13419);
nand U22931 (N_22931,N_17719,N_17109);
nand U22932 (N_22932,N_18244,N_14504);
nand U22933 (N_22933,N_13409,N_16146);
and U22934 (N_22934,N_18527,N_15660);
nor U22935 (N_22935,N_15256,N_12888);
and U22936 (N_22936,N_18134,N_14207);
and U22937 (N_22937,N_15299,N_16942);
nor U22938 (N_22938,N_15815,N_12718);
nor U22939 (N_22939,N_15395,N_14174);
nand U22940 (N_22940,N_16946,N_12538);
nand U22941 (N_22941,N_17882,N_16778);
xor U22942 (N_22942,N_15470,N_16432);
nor U22943 (N_22943,N_14691,N_17106);
and U22944 (N_22944,N_14096,N_17997);
and U22945 (N_22945,N_15917,N_17595);
nor U22946 (N_22946,N_15007,N_13854);
or U22947 (N_22947,N_18396,N_15808);
and U22948 (N_22948,N_14363,N_17924);
nor U22949 (N_22949,N_14502,N_14225);
nand U22950 (N_22950,N_15841,N_16249);
nor U22951 (N_22951,N_16081,N_13810);
or U22952 (N_22952,N_16508,N_16792);
nand U22953 (N_22953,N_13186,N_15106);
or U22954 (N_22954,N_13678,N_15856);
nor U22955 (N_22955,N_13955,N_15265);
xor U22956 (N_22956,N_16121,N_15181);
nor U22957 (N_22957,N_16112,N_15058);
and U22958 (N_22958,N_13015,N_17618);
nand U22959 (N_22959,N_15096,N_16715);
and U22960 (N_22960,N_13610,N_15844);
or U22961 (N_22961,N_14748,N_17882);
nor U22962 (N_22962,N_13606,N_12975);
nand U22963 (N_22963,N_15583,N_18041);
nor U22964 (N_22964,N_13341,N_14078);
nand U22965 (N_22965,N_17649,N_16498);
and U22966 (N_22966,N_13693,N_14334);
nand U22967 (N_22967,N_17012,N_13053);
xnor U22968 (N_22968,N_16321,N_14681);
nor U22969 (N_22969,N_14417,N_15353);
xor U22970 (N_22970,N_17607,N_14800);
xor U22971 (N_22971,N_16318,N_13758);
and U22972 (N_22972,N_12716,N_14584);
xor U22973 (N_22973,N_14101,N_17732);
and U22974 (N_22974,N_18019,N_16505);
nand U22975 (N_22975,N_14682,N_13405);
or U22976 (N_22976,N_13856,N_14684);
and U22977 (N_22977,N_16585,N_16464);
xor U22978 (N_22978,N_16273,N_18485);
or U22979 (N_22979,N_15096,N_15397);
nand U22980 (N_22980,N_12891,N_17576);
nand U22981 (N_22981,N_17517,N_15210);
xor U22982 (N_22982,N_14091,N_14077);
xor U22983 (N_22983,N_13825,N_13684);
nand U22984 (N_22984,N_16175,N_15084);
xor U22985 (N_22985,N_18748,N_12508);
xor U22986 (N_22986,N_17220,N_13402);
nand U22987 (N_22987,N_15530,N_15925);
nand U22988 (N_22988,N_15554,N_17400);
and U22989 (N_22989,N_13218,N_15005);
nand U22990 (N_22990,N_17277,N_14605);
nor U22991 (N_22991,N_14575,N_13914);
or U22992 (N_22992,N_13498,N_17317);
and U22993 (N_22993,N_17488,N_13797);
and U22994 (N_22994,N_17969,N_17820);
nor U22995 (N_22995,N_15090,N_14310);
and U22996 (N_22996,N_15448,N_16565);
nor U22997 (N_22997,N_13485,N_16628);
and U22998 (N_22998,N_14089,N_17896);
or U22999 (N_22999,N_13803,N_16613);
xnor U23000 (N_23000,N_17433,N_13740);
nor U23001 (N_23001,N_16149,N_16614);
nand U23002 (N_23002,N_14801,N_16029);
nor U23003 (N_23003,N_17072,N_13234);
or U23004 (N_23004,N_14370,N_14857);
and U23005 (N_23005,N_16941,N_17707);
or U23006 (N_23006,N_12827,N_18454);
xnor U23007 (N_23007,N_17354,N_17616);
nor U23008 (N_23008,N_16122,N_15204);
xnor U23009 (N_23009,N_15912,N_14229);
nor U23010 (N_23010,N_16855,N_13446);
xor U23011 (N_23011,N_16781,N_15506);
nor U23012 (N_23012,N_17913,N_13615);
and U23013 (N_23013,N_17595,N_16974);
xor U23014 (N_23014,N_14403,N_18704);
nor U23015 (N_23015,N_16201,N_17550);
nor U23016 (N_23016,N_15826,N_13747);
nor U23017 (N_23017,N_17966,N_16160);
nand U23018 (N_23018,N_16983,N_15808);
and U23019 (N_23019,N_14613,N_16810);
and U23020 (N_23020,N_16691,N_14977);
or U23021 (N_23021,N_18423,N_18572);
and U23022 (N_23022,N_13038,N_12700);
nand U23023 (N_23023,N_18055,N_18157);
and U23024 (N_23024,N_16183,N_14254);
nand U23025 (N_23025,N_17100,N_13711);
nand U23026 (N_23026,N_15199,N_16964);
xnor U23027 (N_23027,N_12743,N_14239);
nor U23028 (N_23028,N_13983,N_14274);
and U23029 (N_23029,N_14953,N_13429);
xor U23030 (N_23030,N_13815,N_15566);
nor U23031 (N_23031,N_13171,N_17756);
or U23032 (N_23032,N_15330,N_18494);
nand U23033 (N_23033,N_14062,N_16533);
nand U23034 (N_23034,N_13389,N_13988);
nand U23035 (N_23035,N_18739,N_17973);
xor U23036 (N_23036,N_13413,N_14565);
xor U23037 (N_23037,N_14329,N_13499);
nor U23038 (N_23038,N_16964,N_12814);
or U23039 (N_23039,N_16021,N_17459);
xnor U23040 (N_23040,N_16393,N_16028);
or U23041 (N_23041,N_15613,N_13201);
xor U23042 (N_23042,N_15621,N_17933);
nor U23043 (N_23043,N_14290,N_17086);
or U23044 (N_23044,N_16255,N_17765);
and U23045 (N_23045,N_18470,N_18159);
nand U23046 (N_23046,N_18498,N_15320);
and U23047 (N_23047,N_14436,N_16628);
and U23048 (N_23048,N_17914,N_14618);
xor U23049 (N_23049,N_13093,N_17390);
and U23050 (N_23050,N_16642,N_14394);
nand U23051 (N_23051,N_16890,N_16161);
or U23052 (N_23052,N_14770,N_17683);
or U23053 (N_23053,N_13606,N_14684);
nand U23054 (N_23054,N_15928,N_18533);
and U23055 (N_23055,N_16358,N_14733);
nand U23056 (N_23056,N_14820,N_16490);
xnor U23057 (N_23057,N_17412,N_14246);
and U23058 (N_23058,N_18142,N_14887);
xnor U23059 (N_23059,N_17638,N_13469);
nand U23060 (N_23060,N_17349,N_15256);
or U23061 (N_23061,N_17859,N_13479);
xnor U23062 (N_23062,N_14771,N_12629);
and U23063 (N_23063,N_17300,N_17971);
and U23064 (N_23064,N_14282,N_13288);
nor U23065 (N_23065,N_15450,N_13077);
nand U23066 (N_23066,N_14011,N_18175);
or U23067 (N_23067,N_16711,N_15463);
nand U23068 (N_23068,N_16562,N_14936);
nor U23069 (N_23069,N_14282,N_14345);
xor U23070 (N_23070,N_17828,N_14741);
xor U23071 (N_23071,N_13651,N_16523);
and U23072 (N_23072,N_16016,N_13649);
nand U23073 (N_23073,N_14253,N_14900);
or U23074 (N_23074,N_18610,N_18578);
nor U23075 (N_23075,N_13845,N_12761);
and U23076 (N_23076,N_14038,N_16396);
nor U23077 (N_23077,N_14223,N_17044);
and U23078 (N_23078,N_15612,N_16200);
and U23079 (N_23079,N_13218,N_15829);
nor U23080 (N_23080,N_14495,N_16628);
xor U23081 (N_23081,N_15767,N_15361);
or U23082 (N_23082,N_17149,N_16070);
xnor U23083 (N_23083,N_12771,N_18232);
nor U23084 (N_23084,N_15491,N_13823);
xnor U23085 (N_23085,N_15662,N_18149);
nor U23086 (N_23086,N_12758,N_18480);
nor U23087 (N_23087,N_18126,N_14648);
nor U23088 (N_23088,N_14770,N_14807);
nor U23089 (N_23089,N_16722,N_14192);
or U23090 (N_23090,N_13493,N_12998);
nand U23091 (N_23091,N_17430,N_16503);
and U23092 (N_23092,N_16479,N_15764);
or U23093 (N_23093,N_12731,N_13823);
nand U23094 (N_23094,N_18252,N_18461);
nor U23095 (N_23095,N_18353,N_16180);
nand U23096 (N_23096,N_16644,N_16903);
and U23097 (N_23097,N_17833,N_18431);
nand U23098 (N_23098,N_18578,N_15029);
nand U23099 (N_23099,N_12662,N_17925);
and U23100 (N_23100,N_14328,N_17135);
xor U23101 (N_23101,N_16751,N_14003);
xnor U23102 (N_23102,N_12682,N_17183);
nand U23103 (N_23103,N_14051,N_18083);
and U23104 (N_23104,N_17776,N_12906);
or U23105 (N_23105,N_13220,N_12538);
or U23106 (N_23106,N_17033,N_16909);
or U23107 (N_23107,N_15296,N_18567);
nor U23108 (N_23108,N_14143,N_15811);
or U23109 (N_23109,N_13643,N_18512);
nor U23110 (N_23110,N_12520,N_15286);
nand U23111 (N_23111,N_12877,N_18212);
or U23112 (N_23112,N_15930,N_18664);
and U23113 (N_23113,N_12693,N_15299);
and U23114 (N_23114,N_17585,N_13480);
nor U23115 (N_23115,N_15064,N_13854);
xnor U23116 (N_23116,N_14979,N_12768);
or U23117 (N_23117,N_12768,N_15139);
xor U23118 (N_23118,N_14251,N_15931);
nor U23119 (N_23119,N_13375,N_12648);
nor U23120 (N_23120,N_14415,N_13561);
nand U23121 (N_23121,N_14838,N_15950);
xnor U23122 (N_23122,N_17879,N_15702);
nor U23123 (N_23123,N_13661,N_16856);
or U23124 (N_23124,N_16673,N_15493);
nor U23125 (N_23125,N_15346,N_14913);
and U23126 (N_23126,N_14467,N_14685);
or U23127 (N_23127,N_14935,N_13215);
or U23128 (N_23128,N_14753,N_12986);
nand U23129 (N_23129,N_15180,N_13922);
nor U23130 (N_23130,N_12514,N_16062);
nor U23131 (N_23131,N_12991,N_17066);
and U23132 (N_23132,N_16851,N_17374);
and U23133 (N_23133,N_13575,N_16534);
nor U23134 (N_23134,N_15515,N_14338);
nor U23135 (N_23135,N_13838,N_18248);
nor U23136 (N_23136,N_13906,N_12755);
and U23137 (N_23137,N_14014,N_13234);
nor U23138 (N_23138,N_18255,N_17676);
xor U23139 (N_23139,N_18512,N_16414);
or U23140 (N_23140,N_17862,N_15904);
or U23141 (N_23141,N_15459,N_14479);
nor U23142 (N_23142,N_15387,N_14341);
nand U23143 (N_23143,N_15332,N_17231);
or U23144 (N_23144,N_15338,N_16999);
nand U23145 (N_23145,N_18164,N_13548);
nand U23146 (N_23146,N_17147,N_13610);
nand U23147 (N_23147,N_15273,N_14887);
or U23148 (N_23148,N_17494,N_14104);
xnor U23149 (N_23149,N_18365,N_14279);
and U23150 (N_23150,N_14966,N_17688);
nand U23151 (N_23151,N_14859,N_16185);
and U23152 (N_23152,N_16770,N_18471);
nor U23153 (N_23153,N_16385,N_18657);
xnor U23154 (N_23154,N_13221,N_13161);
xnor U23155 (N_23155,N_12975,N_14782);
nor U23156 (N_23156,N_17166,N_13378);
xnor U23157 (N_23157,N_18216,N_17945);
nand U23158 (N_23158,N_13732,N_17531);
and U23159 (N_23159,N_15994,N_14131);
nor U23160 (N_23160,N_17900,N_14148);
or U23161 (N_23161,N_16835,N_18562);
nor U23162 (N_23162,N_18428,N_18003);
nand U23163 (N_23163,N_16570,N_16101);
or U23164 (N_23164,N_12731,N_16893);
nor U23165 (N_23165,N_16767,N_14934);
or U23166 (N_23166,N_16306,N_13875);
or U23167 (N_23167,N_14568,N_13986);
nor U23168 (N_23168,N_15616,N_17772);
nand U23169 (N_23169,N_14072,N_13063);
or U23170 (N_23170,N_12521,N_17394);
and U23171 (N_23171,N_17602,N_16529);
or U23172 (N_23172,N_13508,N_13319);
or U23173 (N_23173,N_14740,N_14644);
nor U23174 (N_23174,N_12778,N_13999);
xnor U23175 (N_23175,N_17525,N_12735);
and U23176 (N_23176,N_14239,N_17632);
or U23177 (N_23177,N_17339,N_17472);
or U23178 (N_23178,N_13922,N_16814);
or U23179 (N_23179,N_18639,N_16232);
xnor U23180 (N_23180,N_13272,N_14499);
and U23181 (N_23181,N_14615,N_17888);
or U23182 (N_23182,N_15343,N_14553);
xnor U23183 (N_23183,N_16053,N_12805);
nor U23184 (N_23184,N_16861,N_16592);
nor U23185 (N_23185,N_15503,N_14418);
or U23186 (N_23186,N_13689,N_15931);
xnor U23187 (N_23187,N_17583,N_16269);
or U23188 (N_23188,N_13324,N_16395);
xor U23189 (N_23189,N_16577,N_12961);
or U23190 (N_23190,N_15117,N_13654);
nor U23191 (N_23191,N_17494,N_14680);
or U23192 (N_23192,N_14470,N_15287);
nor U23193 (N_23193,N_18726,N_13855);
nor U23194 (N_23194,N_15322,N_18055);
nor U23195 (N_23195,N_18350,N_13131);
nand U23196 (N_23196,N_17388,N_16610);
and U23197 (N_23197,N_18581,N_16417);
xnor U23198 (N_23198,N_14185,N_13188);
xor U23199 (N_23199,N_16412,N_18239);
xnor U23200 (N_23200,N_15207,N_18239);
nor U23201 (N_23201,N_17877,N_16753);
nand U23202 (N_23202,N_14008,N_14974);
nand U23203 (N_23203,N_16495,N_18396);
nand U23204 (N_23204,N_15235,N_18187);
or U23205 (N_23205,N_13392,N_12968);
or U23206 (N_23206,N_13856,N_13524);
and U23207 (N_23207,N_16073,N_15370);
nor U23208 (N_23208,N_14990,N_13418);
and U23209 (N_23209,N_14342,N_16477);
xor U23210 (N_23210,N_18030,N_16174);
nand U23211 (N_23211,N_18495,N_18225);
and U23212 (N_23212,N_14099,N_18744);
and U23213 (N_23213,N_13648,N_16597);
or U23214 (N_23214,N_15329,N_14739);
xor U23215 (N_23215,N_14055,N_13495);
nor U23216 (N_23216,N_15741,N_15504);
xor U23217 (N_23217,N_16591,N_18655);
nand U23218 (N_23218,N_17423,N_13465);
and U23219 (N_23219,N_15110,N_18325);
or U23220 (N_23220,N_14938,N_18129);
xor U23221 (N_23221,N_17104,N_13511);
and U23222 (N_23222,N_13434,N_13372);
nand U23223 (N_23223,N_17727,N_12762);
xnor U23224 (N_23224,N_16583,N_17789);
nand U23225 (N_23225,N_12712,N_14045);
and U23226 (N_23226,N_12795,N_17834);
nor U23227 (N_23227,N_16750,N_18655);
xnor U23228 (N_23228,N_13089,N_12920);
or U23229 (N_23229,N_16724,N_16651);
and U23230 (N_23230,N_17912,N_16505);
nor U23231 (N_23231,N_17077,N_16634);
xnor U23232 (N_23232,N_14989,N_18591);
nand U23233 (N_23233,N_13585,N_15467);
xor U23234 (N_23234,N_17504,N_15347);
and U23235 (N_23235,N_17804,N_16663);
or U23236 (N_23236,N_13083,N_17397);
and U23237 (N_23237,N_16818,N_13062);
xnor U23238 (N_23238,N_14944,N_15389);
and U23239 (N_23239,N_16561,N_16238);
or U23240 (N_23240,N_13937,N_18457);
or U23241 (N_23241,N_14811,N_15332);
nor U23242 (N_23242,N_16579,N_18183);
nand U23243 (N_23243,N_13183,N_14509);
xnor U23244 (N_23244,N_13530,N_13418);
nor U23245 (N_23245,N_13920,N_15459);
or U23246 (N_23246,N_13705,N_16471);
nand U23247 (N_23247,N_16326,N_12991);
nor U23248 (N_23248,N_12784,N_16375);
nor U23249 (N_23249,N_17411,N_18515);
or U23250 (N_23250,N_12580,N_14815);
or U23251 (N_23251,N_14514,N_18544);
and U23252 (N_23252,N_14209,N_14563);
nor U23253 (N_23253,N_12921,N_14144);
or U23254 (N_23254,N_14128,N_15196);
nor U23255 (N_23255,N_13040,N_12522);
nor U23256 (N_23256,N_15326,N_15351);
and U23257 (N_23257,N_18128,N_12673);
xor U23258 (N_23258,N_16893,N_17901);
or U23259 (N_23259,N_17247,N_18743);
nand U23260 (N_23260,N_14215,N_17956);
or U23261 (N_23261,N_15865,N_12990);
and U23262 (N_23262,N_13420,N_13017);
or U23263 (N_23263,N_13040,N_18471);
and U23264 (N_23264,N_12523,N_15159);
xor U23265 (N_23265,N_16105,N_15983);
nand U23266 (N_23266,N_18364,N_17649);
or U23267 (N_23267,N_13725,N_17036);
nand U23268 (N_23268,N_18237,N_13082);
and U23269 (N_23269,N_14467,N_13214);
xor U23270 (N_23270,N_15034,N_14904);
or U23271 (N_23271,N_15545,N_17443);
xor U23272 (N_23272,N_18205,N_18664);
xor U23273 (N_23273,N_13937,N_13310);
nand U23274 (N_23274,N_14290,N_17836);
xnor U23275 (N_23275,N_16136,N_14179);
nor U23276 (N_23276,N_15179,N_15989);
nand U23277 (N_23277,N_16408,N_17710);
nor U23278 (N_23278,N_14076,N_16880);
nand U23279 (N_23279,N_17598,N_12971);
nand U23280 (N_23280,N_18381,N_14116);
xnor U23281 (N_23281,N_16014,N_18450);
xnor U23282 (N_23282,N_15464,N_17519);
xnor U23283 (N_23283,N_15421,N_18433);
and U23284 (N_23284,N_18563,N_18527);
or U23285 (N_23285,N_18291,N_14720);
or U23286 (N_23286,N_12968,N_15967);
nand U23287 (N_23287,N_17135,N_14532);
and U23288 (N_23288,N_13983,N_16395);
and U23289 (N_23289,N_14674,N_17982);
or U23290 (N_23290,N_14988,N_16880);
and U23291 (N_23291,N_13757,N_14017);
nor U23292 (N_23292,N_17008,N_16166);
xor U23293 (N_23293,N_16046,N_13712);
xor U23294 (N_23294,N_14210,N_17659);
nor U23295 (N_23295,N_16524,N_13090);
or U23296 (N_23296,N_17262,N_14719);
and U23297 (N_23297,N_17813,N_12849);
and U23298 (N_23298,N_13808,N_15502);
and U23299 (N_23299,N_13268,N_17325);
nand U23300 (N_23300,N_17190,N_15049);
nand U23301 (N_23301,N_13273,N_16011);
nor U23302 (N_23302,N_12912,N_14496);
xor U23303 (N_23303,N_13772,N_14374);
xor U23304 (N_23304,N_16687,N_14249);
nand U23305 (N_23305,N_16565,N_15114);
and U23306 (N_23306,N_18199,N_13037);
xnor U23307 (N_23307,N_16340,N_12680);
or U23308 (N_23308,N_17796,N_17473);
nor U23309 (N_23309,N_14100,N_14095);
and U23310 (N_23310,N_17846,N_12775);
nor U23311 (N_23311,N_18432,N_16089);
and U23312 (N_23312,N_18704,N_14118);
or U23313 (N_23313,N_15952,N_12932);
and U23314 (N_23314,N_14477,N_14822);
nand U23315 (N_23315,N_14094,N_16226);
nor U23316 (N_23316,N_13769,N_15149);
or U23317 (N_23317,N_18709,N_16280);
or U23318 (N_23318,N_18347,N_15346);
or U23319 (N_23319,N_13437,N_15976);
xor U23320 (N_23320,N_15586,N_16725);
or U23321 (N_23321,N_15018,N_17579);
xor U23322 (N_23322,N_18709,N_18280);
nand U23323 (N_23323,N_18437,N_18127);
xor U23324 (N_23324,N_18627,N_12566);
nand U23325 (N_23325,N_14197,N_17103);
and U23326 (N_23326,N_16771,N_18673);
or U23327 (N_23327,N_14047,N_18691);
and U23328 (N_23328,N_17963,N_18436);
nand U23329 (N_23329,N_16336,N_15042);
nor U23330 (N_23330,N_12962,N_12584);
xor U23331 (N_23331,N_16951,N_13653);
nor U23332 (N_23332,N_12639,N_16386);
or U23333 (N_23333,N_16036,N_17928);
xnor U23334 (N_23334,N_13593,N_14020);
and U23335 (N_23335,N_13917,N_17381);
and U23336 (N_23336,N_16424,N_13258);
nand U23337 (N_23337,N_15628,N_13014);
or U23338 (N_23338,N_13285,N_15908);
nor U23339 (N_23339,N_17017,N_13702);
and U23340 (N_23340,N_15568,N_14616);
and U23341 (N_23341,N_13015,N_16244);
or U23342 (N_23342,N_16132,N_12772);
xnor U23343 (N_23343,N_13335,N_12990);
nand U23344 (N_23344,N_18418,N_13578);
and U23345 (N_23345,N_17314,N_15560);
xnor U23346 (N_23346,N_13383,N_15091);
nand U23347 (N_23347,N_18500,N_15461);
nor U23348 (N_23348,N_14513,N_16576);
nor U23349 (N_23349,N_13342,N_16614);
nand U23350 (N_23350,N_12758,N_18286);
or U23351 (N_23351,N_17497,N_13173);
xor U23352 (N_23352,N_17360,N_15996);
nor U23353 (N_23353,N_18331,N_15249);
nand U23354 (N_23354,N_16935,N_16129);
nor U23355 (N_23355,N_13451,N_12812);
nand U23356 (N_23356,N_13657,N_18459);
and U23357 (N_23357,N_12848,N_18204);
xnor U23358 (N_23358,N_12822,N_15569);
nand U23359 (N_23359,N_12914,N_16529);
xnor U23360 (N_23360,N_18577,N_14760);
nor U23361 (N_23361,N_14493,N_14369);
xor U23362 (N_23362,N_14884,N_13309);
nand U23363 (N_23363,N_16150,N_14836);
xnor U23364 (N_23364,N_13662,N_15423);
nand U23365 (N_23365,N_12765,N_13294);
nand U23366 (N_23366,N_15907,N_15100);
xor U23367 (N_23367,N_13902,N_16099);
or U23368 (N_23368,N_16097,N_16365);
and U23369 (N_23369,N_13171,N_13362);
xnor U23370 (N_23370,N_18382,N_15818);
nor U23371 (N_23371,N_15596,N_13892);
xnor U23372 (N_23372,N_18598,N_14214);
and U23373 (N_23373,N_13272,N_16235);
and U23374 (N_23374,N_13084,N_16925);
or U23375 (N_23375,N_16015,N_12969);
xor U23376 (N_23376,N_15151,N_18237);
nand U23377 (N_23377,N_13599,N_13349);
or U23378 (N_23378,N_14223,N_18523);
xor U23379 (N_23379,N_16660,N_14384);
xnor U23380 (N_23380,N_14807,N_13895);
nor U23381 (N_23381,N_13737,N_18001);
or U23382 (N_23382,N_18320,N_13539);
nor U23383 (N_23383,N_14717,N_17035);
and U23384 (N_23384,N_13049,N_18150);
or U23385 (N_23385,N_14289,N_17229);
nand U23386 (N_23386,N_15729,N_16419);
xnor U23387 (N_23387,N_12553,N_12861);
or U23388 (N_23388,N_17255,N_12932);
and U23389 (N_23389,N_17742,N_13165);
or U23390 (N_23390,N_18335,N_15029);
or U23391 (N_23391,N_12780,N_12904);
and U23392 (N_23392,N_17819,N_15426);
and U23393 (N_23393,N_14520,N_13033);
nand U23394 (N_23394,N_14083,N_15170);
nand U23395 (N_23395,N_16236,N_16389);
xnor U23396 (N_23396,N_12551,N_15369);
or U23397 (N_23397,N_13756,N_14052);
nand U23398 (N_23398,N_13048,N_16039);
and U23399 (N_23399,N_18224,N_18638);
nor U23400 (N_23400,N_18324,N_18308);
nor U23401 (N_23401,N_17198,N_15181);
nand U23402 (N_23402,N_17163,N_16596);
or U23403 (N_23403,N_14409,N_15277);
nor U23404 (N_23404,N_18727,N_16229);
and U23405 (N_23405,N_16270,N_15100);
xnor U23406 (N_23406,N_17798,N_12660);
nor U23407 (N_23407,N_16470,N_16239);
xnor U23408 (N_23408,N_13204,N_14011);
and U23409 (N_23409,N_13462,N_14817);
xor U23410 (N_23410,N_18633,N_14543);
or U23411 (N_23411,N_15065,N_13486);
nor U23412 (N_23412,N_14371,N_13453);
nor U23413 (N_23413,N_14383,N_13568);
xor U23414 (N_23414,N_18400,N_12791);
and U23415 (N_23415,N_15952,N_14923);
nor U23416 (N_23416,N_17013,N_16770);
and U23417 (N_23417,N_17899,N_12751);
xor U23418 (N_23418,N_18333,N_18308);
and U23419 (N_23419,N_18526,N_12503);
and U23420 (N_23420,N_12758,N_16143);
nand U23421 (N_23421,N_14383,N_15048);
nand U23422 (N_23422,N_18208,N_13057);
nand U23423 (N_23423,N_16716,N_12525);
or U23424 (N_23424,N_18639,N_16216);
or U23425 (N_23425,N_12842,N_12884);
nand U23426 (N_23426,N_17822,N_13226);
nand U23427 (N_23427,N_15175,N_18280);
nand U23428 (N_23428,N_12769,N_17489);
or U23429 (N_23429,N_15357,N_15036);
nor U23430 (N_23430,N_15697,N_17793);
or U23431 (N_23431,N_17791,N_18296);
and U23432 (N_23432,N_17039,N_17256);
nor U23433 (N_23433,N_13578,N_18453);
nor U23434 (N_23434,N_14521,N_13057);
nand U23435 (N_23435,N_18514,N_18268);
or U23436 (N_23436,N_17209,N_12810);
xnor U23437 (N_23437,N_18364,N_17719);
nand U23438 (N_23438,N_16176,N_15110);
xor U23439 (N_23439,N_17395,N_14733);
and U23440 (N_23440,N_16261,N_13893);
nand U23441 (N_23441,N_12539,N_16232);
and U23442 (N_23442,N_15097,N_13427);
xnor U23443 (N_23443,N_16089,N_15837);
and U23444 (N_23444,N_16702,N_18623);
and U23445 (N_23445,N_16039,N_15956);
xnor U23446 (N_23446,N_13104,N_15299);
and U23447 (N_23447,N_18123,N_15053);
nor U23448 (N_23448,N_15512,N_14062);
nand U23449 (N_23449,N_16043,N_18387);
or U23450 (N_23450,N_16034,N_15261);
nor U23451 (N_23451,N_17546,N_16114);
and U23452 (N_23452,N_14290,N_14452);
nand U23453 (N_23453,N_16457,N_14174);
and U23454 (N_23454,N_14322,N_13968);
nand U23455 (N_23455,N_16005,N_13641);
nor U23456 (N_23456,N_15781,N_17168);
xnor U23457 (N_23457,N_15268,N_16878);
nand U23458 (N_23458,N_13579,N_12525);
and U23459 (N_23459,N_13372,N_16263);
and U23460 (N_23460,N_15597,N_16426);
nand U23461 (N_23461,N_18659,N_15742);
nand U23462 (N_23462,N_14867,N_13874);
nand U23463 (N_23463,N_15285,N_17454);
xnor U23464 (N_23464,N_12557,N_14738);
nand U23465 (N_23465,N_16426,N_14649);
and U23466 (N_23466,N_14172,N_13213);
xnor U23467 (N_23467,N_16323,N_15928);
xor U23468 (N_23468,N_14085,N_17322);
and U23469 (N_23469,N_18564,N_15142);
nand U23470 (N_23470,N_13350,N_18447);
or U23471 (N_23471,N_18136,N_13025);
nand U23472 (N_23472,N_16371,N_16886);
and U23473 (N_23473,N_14251,N_12578);
nor U23474 (N_23474,N_14924,N_18135);
xor U23475 (N_23475,N_17618,N_12540);
nor U23476 (N_23476,N_13051,N_13131);
nand U23477 (N_23477,N_13814,N_16341);
nor U23478 (N_23478,N_13858,N_15379);
nor U23479 (N_23479,N_13159,N_15575);
and U23480 (N_23480,N_13778,N_15535);
nor U23481 (N_23481,N_15116,N_15948);
nor U23482 (N_23482,N_14191,N_14912);
nand U23483 (N_23483,N_15790,N_16901);
and U23484 (N_23484,N_18683,N_16491);
xnor U23485 (N_23485,N_13045,N_12545);
nand U23486 (N_23486,N_17950,N_16887);
and U23487 (N_23487,N_15102,N_16404);
xor U23488 (N_23488,N_12583,N_18381);
and U23489 (N_23489,N_18483,N_12636);
nand U23490 (N_23490,N_14478,N_16162);
or U23491 (N_23491,N_15666,N_16306);
and U23492 (N_23492,N_18535,N_14519);
nand U23493 (N_23493,N_14966,N_14766);
and U23494 (N_23494,N_15885,N_13860);
nand U23495 (N_23495,N_16012,N_16009);
and U23496 (N_23496,N_16346,N_13677);
and U23497 (N_23497,N_14596,N_14672);
and U23498 (N_23498,N_18454,N_15213);
nand U23499 (N_23499,N_14195,N_13544);
xor U23500 (N_23500,N_18693,N_16944);
nor U23501 (N_23501,N_13728,N_17228);
nand U23502 (N_23502,N_15135,N_13966);
and U23503 (N_23503,N_15023,N_12892);
and U23504 (N_23504,N_14942,N_15441);
nand U23505 (N_23505,N_16589,N_15417);
and U23506 (N_23506,N_13406,N_14968);
and U23507 (N_23507,N_18582,N_16189);
nor U23508 (N_23508,N_17881,N_17850);
and U23509 (N_23509,N_14513,N_15644);
or U23510 (N_23510,N_17347,N_16446);
nand U23511 (N_23511,N_18391,N_18321);
nor U23512 (N_23512,N_15599,N_18664);
nor U23513 (N_23513,N_12966,N_18038);
xor U23514 (N_23514,N_17264,N_18078);
xnor U23515 (N_23515,N_17096,N_17842);
or U23516 (N_23516,N_12888,N_16500);
nor U23517 (N_23517,N_18013,N_13954);
nand U23518 (N_23518,N_16382,N_17074);
and U23519 (N_23519,N_12723,N_16980);
or U23520 (N_23520,N_12835,N_16716);
nand U23521 (N_23521,N_15238,N_16269);
xnor U23522 (N_23522,N_15205,N_15571);
and U23523 (N_23523,N_16695,N_15115);
nand U23524 (N_23524,N_15083,N_15430);
nor U23525 (N_23525,N_15744,N_14833);
nor U23526 (N_23526,N_16314,N_14166);
and U23527 (N_23527,N_14345,N_13165);
nand U23528 (N_23528,N_16003,N_18218);
nor U23529 (N_23529,N_13421,N_13637);
or U23530 (N_23530,N_12817,N_16390);
and U23531 (N_23531,N_16567,N_16849);
xor U23532 (N_23532,N_14028,N_13530);
nor U23533 (N_23533,N_18499,N_14236);
or U23534 (N_23534,N_17206,N_13178);
and U23535 (N_23535,N_18377,N_13674);
or U23536 (N_23536,N_15970,N_17257);
or U23537 (N_23537,N_18419,N_16801);
nand U23538 (N_23538,N_16741,N_13945);
nor U23539 (N_23539,N_17594,N_18501);
or U23540 (N_23540,N_14327,N_12754);
or U23541 (N_23541,N_12804,N_18108);
or U23542 (N_23542,N_16608,N_14873);
or U23543 (N_23543,N_13451,N_18497);
or U23544 (N_23544,N_13849,N_15780);
or U23545 (N_23545,N_17362,N_18360);
nand U23546 (N_23546,N_14362,N_18632);
nand U23547 (N_23547,N_14480,N_18602);
and U23548 (N_23548,N_18628,N_14013);
nand U23549 (N_23549,N_18316,N_12587);
xnor U23550 (N_23550,N_14368,N_14308);
nand U23551 (N_23551,N_17368,N_14484);
nand U23552 (N_23552,N_13761,N_17382);
and U23553 (N_23553,N_17751,N_13603);
and U23554 (N_23554,N_15905,N_16166);
nor U23555 (N_23555,N_14749,N_16847);
xor U23556 (N_23556,N_17803,N_14753);
xor U23557 (N_23557,N_18123,N_14984);
and U23558 (N_23558,N_12645,N_16288);
nor U23559 (N_23559,N_16008,N_13461);
or U23560 (N_23560,N_12946,N_16294);
nor U23561 (N_23561,N_17422,N_14082);
xnor U23562 (N_23562,N_13100,N_17159);
and U23563 (N_23563,N_18216,N_14702);
or U23564 (N_23564,N_14728,N_16265);
nor U23565 (N_23565,N_18073,N_17458);
or U23566 (N_23566,N_16960,N_14888);
or U23567 (N_23567,N_14245,N_14454);
xnor U23568 (N_23568,N_14124,N_13587);
or U23569 (N_23569,N_14125,N_13414);
or U23570 (N_23570,N_15021,N_12531);
xor U23571 (N_23571,N_14112,N_17546);
or U23572 (N_23572,N_14640,N_14710);
nor U23573 (N_23573,N_15119,N_15099);
and U23574 (N_23574,N_13654,N_16515);
or U23575 (N_23575,N_15516,N_12560);
and U23576 (N_23576,N_18399,N_14180);
nand U23577 (N_23577,N_18328,N_18482);
nand U23578 (N_23578,N_15827,N_15617);
nor U23579 (N_23579,N_14248,N_14041);
and U23580 (N_23580,N_12669,N_13240);
and U23581 (N_23581,N_16300,N_16030);
nand U23582 (N_23582,N_18522,N_14364);
xnor U23583 (N_23583,N_17806,N_13951);
nor U23584 (N_23584,N_15432,N_16375);
nand U23585 (N_23585,N_14872,N_13364);
nand U23586 (N_23586,N_18281,N_17899);
and U23587 (N_23587,N_16103,N_15914);
or U23588 (N_23588,N_17208,N_15333);
or U23589 (N_23589,N_14087,N_12974);
nor U23590 (N_23590,N_18008,N_16826);
nand U23591 (N_23591,N_17981,N_17549);
nand U23592 (N_23592,N_16688,N_18586);
xnor U23593 (N_23593,N_16791,N_16979);
xnor U23594 (N_23594,N_14127,N_16989);
nand U23595 (N_23595,N_18385,N_14916);
xnor U23596 (N_23596,N_16330,N_17294);
nor U23597 (N_23597,N_13340,N_15807);
and U23598 (N_23598,N_15206,N_17314);
nor U23599 (N_23599,N_17229,N_17160);
and U23600 (N_23600,N_15352,N_18654);
nand U23601 (N_23601,N_17085,N_13777);
nand U23602 (N_23602,N_17344,N_14415);
and U23603 (N_23603,N_16295,N_13427);
or U23604 (N_23604,N_16959,N_16059);
and U23605 (N_23605,N_18097,N_17699);
nand U23606 (N_23606,N_12577,N_13950);
and U23607 (N_23607,N_16652,N_12990);
nor U23608 (N_23608,N_18072,N_16136);
xnor U23609 (N_23609,N_13094,N_15063);
nor U23610 (N_23610,N_16593,N_18744);
nor U23611 (N_23611,N_12850,N_15238);
nor U23612 (N_23612,N_17113,N_17130);
nand U23613 (N_23613,N_13230,N_16265);
nand U23614 (N_23614,N_18133,N_13621);
or U23615 (N_23615,N_13526,N_12987);
nand U23616 (N_23616,N_12881,N_15775);
nor U23617 (N_23617,N_16003,N_13317);
and U23618 (N_23618,N_18655,N_18340);
nand U23619 (N_23619,N_14680,N_14825);
nand U23620 (N_23620,N_13126,N_12759);
or U23621 (N_23621,N_18010,N_13520);
xor U23622 (N_23622,N_13399,N_17516);
nor U23623 (N_23623,N_15067,N_15171);
nor U23624 (N_23624,N_12764,N_17145);
or U23625 (N_23625,N_12665,N_17694);
nor U23626 (N_23626,N_17611,N_12645);
and U23627 (N_23627,N_17765,N_17808);
xor U23628 (N_23628,N_16006,N_18439);
xor U23629 (N_23629,N_13673,N_14843);
and U23630 (N_23630,N_17709,N_17252);
nand U23631 (N_23631,N_12536,N_16067);
nor U23632 (N_23632,N_15091,N_15659);
nand U23633 (N_23633,N_17303,N_14332);
and U23634 (N_23634,N_14620,N_18159);
xnor U23635 (N_23635,N_16897,N_18158);
or U23636 (N_23636,N_12682,N_18112);
nor U23637 (N_23637,N_13491,N_18145);
nor U23638 (N_23638,N_17052,N_12904);
and U23639 (N_23639,N_14316,N_18426);
nand U23640 (N_23640,N_13680,N_13533);
nor U23641 (N_23641,N_12654,N_18572);
and U23642 (N_23642,N_15596,N_18206);
or U23643 (N_23643,N_16518,N_13957);
nand U23644 (N_23644,N_14302,N_16653);
and U23645 (N_23645,N_18304,N_18357);
nor U23646 (N_23646,N_17305,N_15191);
nor U23647 (N_23647,N_13011,N_17129);
xnor U23648 (N_23648,N_17608,N_16577);
nand U23649 (N_23649,N_13718,N_16320);
or U23650 (N_23650,N_12991,N_17518);
nor U23651 (N_23651,N_16036,N_15272);
nand U23652 (N_23652,N_17295,N_13433);
nand U23653 (N_23653,N_16653,N_18049);
nand U23654 (N_23654,N_18615,N_15640);
or U23655 (N_23655,N_13654,N_14015);
xnor U23656 (N_23656,N_18085,N_13429);
and U23657 (N_23657,N_16079,N_15482);
nor U23658 (N_23658,N_13925,N_13629);
nor U23659 (N_23659,N_17114,N_12633);
nor U23660 (N_23660,N_12653,N_16539);
xor U23661 (N_23661,N_15598,N_12529);
nand U23662 (N_23662,N_13769,N_14767);
nand U23663 (N_23663,N_13067,N_13275);
xnor U23664 (N_23664,N_16148,N_12808);
xor U23665 (N_23665,N_17019,N_16420);
nand U23666 (N_23666,N_13711,N_16698);
nor U23667 (N_23667,N_15713,N_16864);
nand U23668 (N_23668,N_14355,N_17749);
xor U23669 (N_23669,N_17028,N_13173);
nand U23670 (N_23670,N_13675,N_12843);
nand U23671 (N_23671,N_15042,N_15234);
nor U23672 (N_23672,N_16048,N_13776);
nand U23673 (N_23673,N_12977,N_15077);
and U23674 (N_23674,N_16953,N_18323);
xor U23675 (N_23675,N_17408,N_16943);
nor U23676 (N_23676,N_16506,N_13132);
nand U23677 (N_23677,N_13200,N_15245);
and U23678 (N_23678,N_16742,N_14879);
xor U23679 (N_23679,N_16111,N_16871);
nor U23680 (N_23680,N_18465,N_16930);
xor U23681 (N_23681,N_16321,N_17432);
nor U23682 (N_23682,N_14435,N_16858);
xnor U23683 (N_23683,N_17843,N_17364);
or U23684 (N_23684,N_15378,N_15499);
or U23685 (N_23685,N_14751,N_13721);
and U23686 (N_23686,N_15283,N_18544);
nor U23687 (N_23687,N_13885,N_18237);
and U23688 (N_23688,N_17448,N_16177);
xor U23689 (N_23689,N_15711,N_15951);
nor U23690 (N_23690,N_13833,N_15736);
and U23691 (N_23691,N_17264,N_14121);
nand U23692 (N_23692,N_14781,N_16149);
nand U23693 (N_23693,N_15366,N_18044);
or U23694 (N_23694,N_16315,N_18484);
and U23695 (N_23695,N_16866,N_13824);
nor U23696 (N_23696,N_16155,N_13787);
nor U23697 (N_23697,N_18221,N_12683);
and U23698 (N_23698,N_14791,N_16094);
or U23699 (N_23699,N_16253,N_17251);
xnor U23700 (N_23700,N_16336,N_15998);
nand U23701 (N_23701,N_17292,N_13536);
nand U23702 (N_23702,N_16410,N_16806);
or U23703 (N_23703,N_16617,N_16809);
or U23704 (N_23704,N_14929,N_16046);
and U23705 (N_23705,N_14060,N_16450);
xor U23706 (N_23706,N_15260,N_17843);
xor U23707 (N_23707,N_17254,N_13631);
xor U23708 (N_23708,N_12578,N_18311);
and U23709 (N_23709,N_13274,N_15991);
or U23710 (N_23710,N_13620,N_14826);
xor U23711 (N_23711,N_14951,N_15017);
nand U23712 (N_23712,N_15955,N_15085);
or U23713 (N_23713,N_12919,N_15892);
xor U23714 (N_23714,N_17533,N_13786);
and U23715 (N_23715,N_18415,N_15877);
nor U23716 (N_23716,N_14518,N_12564);
nor U23717 (N_23717,N_18310,N_15868);
xor U23718 (N_23718,N_12890,N_13457);
nand U23719 (N_23719,N_16146,N_12535);
xor U23720 (N_23720,N_15151,N_13538);
xnor U23721 (N_23721,N_17290,N_16846);
nand U23722 (N_23722,N_17583,N_18726);
nor U23723 (N_23723,N_15310,N_12629);
xor U23724 (N_23724,N_15768,N_17131);
and U23725 (N_23725,N_18286,N_16448);
nand U23726 (N_23726,N_15863,N_18722);
nor U23727 (N_23727,N_14552,N_16748);
nand U23728 (N_23728,N_12741,N_13202);
nor U23729 (N_23729,N_12779,N_18039);
and U23730 (N_23730,N_17173,N_15586);
or U23731 (N_23731,N_15226,N_13835);
nand U23732 (N_23732,N_18190,N_13450);
and U23733 (N_23733,N_14591,N_17724);
nand U23734 (N_23734,N_12551,N_17116);
nand U23735 (N_23735,N_13839,N_13675);
or U23736 (N_23736,N_12881,N_18538);
or U23737 (N_23737,N_14962,N_13188);
or U23738 (N_23738,N_12704,N_13134);
nand U23739 (N_23739,N_12788,N_18478);
xor U23740 (N_23740,N_14183,N_17814);
or U23741 (N_23741,N_13546,N_13234);
nor U23742 (N_23742,N_15873,N_13453);
or U23743 (N_23743,N_17917,N_12673);
nand U23744 (N_23744,N_15335,N_18509);
nand U23745 (N_23745,N_12507,N_18410);
and U23746 (N_23746,N_16237,N_18646);
xor U23747 (N_23747,N_18363,N_16182);
and U23748 (N_23748,N_13648,N_14819);
and U23749 (N_23749,N_18106,N_17866);
or U23750 (N_23750,N_14144,N_17030);
and U23751 (N_23751,N_13276,N_17291);
and U23752 (N_23752,N_17531,N_17626);
nor U23753 (N_23753,N_14880,N_17110);
xor U23754 (N_23754,N_17749,N_12709);
nand U23755 (N_23755,N_12886,N_12978);
nand U23756 (N_23756,N_13310,N_12775);
nand U23757 (N_23757,N_16156,N_16889);
nor U23758 (N_23758,N_17973,N_15494);
nand U23759 (N_23759,N_16366,N_17537);
or U23760 (N_23760,N_14509,N_14311);
nand U23761 (N_23761,N_13858,N_18189);
nor U23762 (N_23762,N_15310,N_17474);
and U23763 (N_23763,N_17261,N_13130);
nand U23764 (N_23764,N_16250,N_18611);
and U23765 (N_23765,N_15801,N_15526);
or U23766 (N_23766,N_13756,N_15579);
and U23767 (N_23767,N_12751,N_17141);
xnor U23768 (N_23768,N_17925,N_15837);
nor U23769 (N_23769,N_12640,N_18147);
or U23770 (N_23770,N_15115,N_15520);
nand U23771 (N_23771,N_14134,N_14877);
nor U23772 (N_23772,N_14999,N_17003);
and U23773 (N_23773,N_15709,N_17068);
nor U23774 (N_23774,N_14430,N_14445);
xnor U23775 (N_23775,N_15536,N_16382);
nand U23776 (N_23776,N_14870,N_13840);
nor U23777 (N_23777,N_18265,N_18725);
nor U23778 (N_23778,N_12790,N_14483);
and U23779 (N_23779,N_12714,N_13463);
or U23780 (N_23780,N_14666,N_12548);
or U23781 (N_23781,N_15845,N_17985);
xor U23782 (N_23782,N_18024,N_18395);
nor U23783 (N_23783,N_12671,N_15031);
and U23784 (N_23784,N_18067,N_17566);
and U23785 (N_23785,N_15861,N_13598);
nand U23786 (N_23786,N_16555,N_18134);
xnor U23787 (N_23787,N_15815,N_13328);
nand U23788 (N_23788,N_15633,N_17578);
or U23789 (N_23789,N_17801,N_16437);
nor U23790 (N_23790,N_16578,N_18341);
or U23791 (N_23791,N_18703,N_13444);
nor U23792 (N_23792,N_18333,N_14166);
nor U23793 (N_23793,N_14432,N_13863);
and U23794 (N_23794,N_15929,N_13253);
nor U23795 (N_23795,N_14378,N_17741);
and U23796 (N_23796,N_16779,N_15815);
nor U23797 (N_23797,N_13354,N_12677);
or U23798 (N_23798,N_16601,N_18425);
and U23799 (N_23799,N_13249,N_18107);
or U23800 (N_23800,N_18733,N_13647);
and U23801 (N_23801,N_12930,N_16407);
xnor U23802 (N_23802,N_18169,N_16836);
or U23803 (N_23803,N_16925,N_18656);
nor U23804 (N_23804,N_17399,N_14355);
and U23805 (N_23805,N_16052,N_12881);
xnor U23806 (N_23806,N_13833,N_15384);
and U23807 (N_23807,N_13608,N_16982);
or U23808 (N_23808,N_12524,N_12720);
nand U23809 (N_23809,N_14359,N_14637);
or U23810 (N_23810,N_12685,N_12829);
nor U23811 (N_23811,N_16021,N_15283);
nand U23812 (N_23812,N_14050,N_13372);
nor U23813 (N_23813,N_12580,N_17064);
nand U23814 (N_23814,N_17663,N_18731);
and U23815 (N_23815,N_16346,N_18440);
or U23816 (N_23816,N_17382,N_17682);
nand U23817 (N_23817,N_18689,N_18270);
xnor U23818 (N_23818,N_13876,N_14259);
and U23819 (N_23819,N_16942,N_15674);
and U23820 (N_23820,N_16211,N_14619);
and U23821 (N_23821,N_16264,N_17480);
nor U23822 (N_23822,N_14856,N_14605);
nand U23823 (N_23823,N_17119,N_18584);
xnor U23824 (N_23824,N_13979,N_16151);
nand U23825 (N_23825,N_15704,N_16882);
xnor U23826 (N_23826,N_12709,N_14380);
nor U23827 (N_23827,N_17122,N_18383);
or U23828 (N_23828,N_12823,N_14537);
nand U23829 (N_23829,N_17753,N_17340);
nand U23830 (N_23830,N_14655,N_17455);
xor U23831 (N_23831,N_15122,N_15292);
and U23832 (N_23832,N_14397,N_12698);
nor U23833 (N_23833,N_15919,N_17035);
or U23834 (N_23834,N_17658,N_13788);
nor U23835 (N_23835,N_17373,N_15237);
or U23836 (N_23836,N_15904,N_16036);
nor U23837 (N_23837,N_15968,N_14881);
or U23838 (N_23838,N_12749,N_18622);
and U23839 (N_23839,N_16921,N_14033);
nand U23840 (N_23840,N_16640,N_14330);
or U23841 (N_23841,N_18073,N_12720);
nor U23842 (N_23842,N_18508,N_15527);
and U23843 (N_23843,N_13562,N_16080);
xor U23844 (N_23844,N_12853,N_18169);
xnor U23845 (N_23845,N_14562,N_13013);
or U23846 (N_23846,N_13518,N_16228);
nand U23847 (N_23847,N_15845,N_13258);
nand U23848 (N_23848,N_12909,N_12758);
nand U23849 (N_23849,N_14925,N_18170);
nor U23850 (N_23850,N_15815,N_15361);
nor U23851 (N_23851,N_14374,N_16951);
xnor U23852 (N_23852,N_13762,N_15052);
nor U23853 (N_23853,N_17410,N_14615);
or U23854 (N_23854,N_16880,N_13926);
nor U23855 (N_23855,N_16542,N_18671);
or U23856 (N_23856,N_16399,N_15149);
nor U23857 (N_23857,N_14631,N_15041);
or U23858 (N_23858,N_17823,N_14701);
nor U23859 (N_23859,N_17765,N_13620);
nor U23860 (N_23860,N_14787,N_13679);
nand U23861 (N_23861,N_18071,N_14280);
and U23862 (N_23862,N_16367,N_17452);
nor U23863 (N_23863,N_17465,N_18749);
xnor U23864 (N_23864,N_15419,N_16496);
nor U23865 (N_23865,N_13902,N_15325);
nand U23866 (N_23866,N_14820,N_15860);
nand U23867 (N_23867,N_13654,N_18726);
nor U23868 (N_23868,N_16529,N_12990);
nand U23869 (N_23869,N_18276,N_15039);
nor U23870 (N_23870,N_18514,N_16138);
nor U23871 (N_23871,N_14765,N_16192);
nor U23872 (N_23872,N_17979,N_13325);
nand U23873 (N_23873,N_16960,N_16030);
or U23874 (N_23874,N_13367,N_12815);
and U23875 (N_23875,N_15571,N_15283);
or U23876 (N_23876,N_18540,N_17632);
xor U23877 (N_23877,N_12910,N_13680);
or U23878 (N_23878,N_16729,N_17533);
and U23879 (N_23879,N_17854,N_17235);
nor U23880 (N_23880,N_13385,N_13836);
and U23881 (N_23881,N_14131,N_15098);
or U23882 (N_23882,N_17227,N_17250);
xnor U23883 (N_23883,N_14128,N_14359);
nor U23884 (N_23884,N_17975,N_15193);
nor U23885 (N_23885,N_13207,N_13396);
and U23886 (N_23886,N_17908,N_17614);
xnor U23887 (N_23887,N_16003,N_17363);
nand U23888 (N_23888,N_12546,N_18021);
xnor U23889 (N_23889,N_14963,N_13720);
nand U23890 (N_23890,N_18099,N_14993);
xor U23891 (N_23891,N_17259,N_13408);
nor U23892 (N_23892,N_16821,N_14146);
and U23893 (N_23893,N_14500,N_18425);
or U23894 (N_23894,N_13308,N_12624);
and U23895 (N_23895,N_16077,N_15002);
nor U23896 (N_23896,N_14102,N_16281);
and U23897 (N_23897,N_17980,N_14138);
or U23898 (N_23898,N_16468,N_15542);
and U23899 (N_23899,N_13828,N_17953);
xor U23900 (N_23900,N_16445,N_15948);
or U23901 (N_23901,N_12638,N_18387);
nor U23902 (N_23902,N_14980,N_12808);
nor U23903 (N_23903,N_15248,N_17082);
nand U23904 (N_23904,N_13644,N_14331);
nor U23905 (N_23905,N_13461,N_14742);
xor U23906 (N_23906,N_14963,N_14646);
xor U23907 (N_23907,N_15465,N_16677);
xnor U23908 (N_23908,N_17005,N_16481);
nand U23909 (N_23909,N_14428,N_14948);
nand U23910 (N_23910,N_17830,N_15052);
nor U23911 (N_23911,N_12538,N_14900);
and U23912 (N_23912,N_16335,N_13891);
nand U23913 (N_23913,N_14501,N_15968);
xnor U23914 (N_23914,N_16382,N_16234);
nor U23915 (N_23915,N_15616,N_17269);
and U23916 (N_23916,N_13404,N_15195);
and U23917 (N_23917,N_13079,N_18269);
or U23918 (N_23918,N_13658,N_12611);
xnor U23919 (N_23919,N_13874,N_15664);
and U23920 (N_23920,N_16074,N_18241);
xnor U23921 (N_23921,N_17364,N_12548);
nand U23922 (N_23922,N_15251,N_15698);
nand U23923 (N_23923,N_14341,N_13764);
nor U23924 (N_23924,N_13359,N_15470);
nand U23925 (N_23925,N_16870,N_15214);
nand U23926 (N_23926,N_15120,N_18093);
or U23927 (N_23927,N_16858,N_13760);
or U23928 (N_23928,N_14476,N_17240);
xor U23929 (N_23929,N_13331,N_13525);
nand U23930 (N_23930,N_13317,N_12793);
and U23931 (N_23931,N_17303,N_14113);
nand U23932 (N_23932,N_17234,N_14730);
xor U23933 (N_23933,N_16223,N_14149);
and U23934 (N_23934,N_12984,N_14101);
nor U23935 (N_23935,N_14799,N_14050);
or U23936 (N_23936,N_18360,N_13413);
or U23937 (N_23937,N_16365,N_15907);
or U23938 (N_23938,N_15547,N_13646);
and U23939 (N_23939,N_17760,N_17183);
or U23940 (N_23940,N_17547,N_17790);
and U23941 (N_23941,N_14210,N_16217);
xnor U23942 (N_23942,N_16176,N_15222);
xor U23943 (N_23943,N_17879,N_15590);
and U23944 (N_23944,N_17196,N_14664);
and U23945 (N_23945,N_17922,N_16587);
xnor U23946 (N_23946,N_16417,N_14920);
nor U23947 (N_23947,N_13900,N_13400);
nand U23948 (N_23948,N_14038,N_16679);
nand U23949 (N_23949,N_15240,N_13174);
nor U23950 (N_23950,N_13695,N_12773);
or U23951 (N_23951,N_14257,N_17998);
nand U23952 (N_23952,N_14561,N_18583);
and U23953 (N_23953,N_17049,N_14077);
xor U23954 (N_23954,N_17979,N_16742);
xnor U23955 (N_23955,N_13031,N_18316);
nand U23956 (N_23956,N_16066,N_14363);
or U23957 (N_23957,N_14414,N_13540);
and U23958 (N_23958,N_17989,N_12772);
nor U23959 (N_23959,N_17050,N_17480);
or U23960 (N_23960,N_16297,N_17437);
nand U23961 (N_23961,N_17392,N_17978);
nor U23962 (N_23962,N_17680,N_14138);
nor U23963 (N_23963,N_12651,N_14675);
and U23964 (N_23964,N_14705,N_12625);
nor U23965 (N_23965,N_13020,N_15832);
and U23966 (N_23966,N_14217,N_18236);
nor U23967 (N_23967,N_17164,N_17154);
and U23968 (N_23968,N_13721,N_12984);
or U23969 (N_23969,N_13264,N_13633);
or U23970 (N_23970,N_17123,N_16352);
nand U23971 (N_23971,N_15438,N_13296);
and U23972 (N_23972,N_16240,N_17456);
nand U23973 (N_23973,N_17490,N_17164);
xnor U23974 (N_23974,N_13885,N_17238);
and U23975 (N_23975,N_17275,N_13245);
nand U23976 (N_23976,N_17106,N_15977);
nor U23977 (N_23977,N_17247,N_12861);
and U23978 (N_23978,N_16434,N_18367);
and U23979 (N_23979,N_12627,N_13030);
and U23980 (N_23980,N_18099,N_15018);
nand U23981 (N_23981,N_14198,N_14566);
or U23982 (N_23982,N_14795,N_14604);
nand U23983 (N_23983,N_14294,N_14737);
or U23984 (N_23984,N_14888,N_16442);
nand U23985 (N_23985,N_14171,N_15850);
xnor U23986 (N_23986,N_16364,N_16187);
or U23987 (N_23987,N_15305,N_14616);
or U23988 (N_23988,N_14305,N_16733);
and U23989 (N_23989,N_13459,N_17272);
or U23990 (N_23990,N_16619,N_12982);
nand U23991 (N_23991,N_18094,N_16027);
or U23992 (N_23992,N_13252,N_13754);
nor U23993 (N_23993,N_15842,N_12607);
nor U23994 (N_23994,N_17781,N_15901);
nand U23995 (N_23995,N_16687,N_13565);
nand U23996 (N_23996,N_15563,N_13600);
nand U23997 (N_23997,N_17973,N_16676);
xor U23998 (N_23998,N_14552,N_18274);
xnor U23999 (N_23999,N_16132,N_12808);
xor U24000 (N_24000,N_14277,N_18640);
or U24001 (N_24001,N_15577,N_13039);
nand U24002 (N_24002,N_13585,N_13825);
or U24003 (N_24003,N_15766,N_15786);
xor U24004 (N_24004,N_12669,N_13352);
or U24005 (N_24005,N_13961,N_16232);
xor U24006 (N_24006,N_13643,N_15200);
nor U24007 (N_24007,N_15800,N_15818);
and U24008 (N_24008,N_17344,N_13147);
and U24009 (N_24009,N_15149,N_17005);
xor U24010 (N_24010,N_16385,N_18689);
xor U24011 (N_24011,N_12696,N_15085);
nand U24012 (N_24012,N_13385,N_16165);
or U24013 (N_24013,N_13973,N_15136);
or U24014 (N_24014,N_17734,N_13662);
nand U24015 (N_24015,N_15876,N_13294);
or U24016 (N_24016,N_13933,N_17253);
or U24017 (N_24017,N_17510,N_12621);
xor U24018 (N_24018,N_13547,N_15333);
or U24019 (N_24019,N_14625,N_16604);
or U24020 (N_24020,N_14537,N_14342);
nand U24021 (N_24021,N_16224,N_14706);
nand U24022 (N_24022,N_15143,N_12913);
or U24023 (N_24023,N_15437,N_15135);
nand U24024 (N_24024,N_17000,N_16112);
and U24025 (N_24025,N_15701,N_14453);
nand U24026 (N_24026,N_15427,N_17537);
nand U24027 (N_24027,N_16825,N_15063);
xor U24028 (N_24028,N_16953,N_16299);
or U24029 (N_24029,N_16499,N_17991);
and U24030 (N_24030,N_13258,N_15688);
or U24031 (N_24031,N_14842,N_12621);
xor U24032 (N_24032,N_12727,N_15713);
or U24033 (N_24033,N_14066,N_13924);
xor U24034 (N_24034,N_13755,N_18440);
nor U24035 (N_24035,N_13587,N_15209);
nand U24036 (N_24036,N_14511,N_15187);
or U24037 (N_24037,N_15189,N_17616);
or U24038 (N_24038,N_16622,N_16568);
xor U24039 (N_24039,N_14790,N_12722);
or U24040 (N_24040,N_17724,N_17243);
and U24041 (N_24041,N_18350,N_16141);
xor U24042 (N_24042,N_17384,N_13780);
or U24043 (N_24043,N_14888,N_18109);
or U24044 (N_24044,N_12789,N_18117);
nor U24045 (N_24045,N_18542,N_16792);
or U24046 (N_24046,N_14332,N_17675);
nand U24047 (N_24047,N_13055,N_17822);
nor U24048 (N_24048,N_17642,N_13716);
xor U24049 (N_24049,N_15609,N_13785);
nand U24050 (N_24050,N_14090,N_13106);
nand U24051 (N_24051,N_12504,N_16704);
nor U24052 (N_24052,N_13912,N_13058);
nand U24053 (N_24053,N_13551,N_16514);
xor U24054 (N_24054,N_16126,N_17293);
nand U24055 (N_24055,N_14655,N_14597);
xnor U24056 (N_24056,N_16334,N_14272);
or U24057 (N_24057,N_16012,N_18719);
xor U24058 (N_24058,N_17657,N_16567);
nor U24059 (N_24059,N_13046,N_16198);
nor U24060 (N_24060,N_15099,N_13627);
nand U24061 (N_24061,N_18406,N_14700);
nor U24062 (N_24062,N_13926,N_16810);
or U24063 (N_24063,N_15574,N_16632);
or U24064 (N_24064,N_14173,N_12713);
xor U24065 (N_24065,N_12662,N_17359);
or U24066 (N_24066,N_14146,N_13843);
and U24067 (N_24067,N_14102,N_18537);
nand U24068 (N_24068,N_16638,N_14349);
nor U24069 (N_24069,N_17455,N_13240);
nand U24070 (N_24070,N_18737,N_13740);
nand U24071 (N_24071,N_13468,N_15588);
xnor U24072 (N_24072,N_14467,N_15112);
or U24073 (N_24073,N_15429,N_17165);
and U24074 (N_24074,N_14465,N_17160);
and U24075 (N_24075,N_13969,N_17374);
or U24076 (N_24076,N_15711,N_18263);
and U24077 (N_24077,N_15815,N_14060);
or U24078 (N_24078,N_16502,N_13100);
and U24079 (N_24079,N_14343,N_16397);
nand U24080 (N_24080,N_15596,N_16748);
or U24081 (N_24081,N_16458,N_13178);
nand U24082 (N_24082,N_16216,N_13456);
and U24083 (N_24083,N_12725,N_16413);
or U24084 (N_24084,N_14481,N_15265);
xor U24085 (N_24085,N_15911,N_16114);
xnor U24086 (N_24086,N_17708,N_15463);
xor U24087 (N_24087,N_12602,N_16753);
and U24088 (N_24088,N_18374,N_13270);
xor U24089 (N_24089,N_13367,N_12622);
xor U24090 (N_24090,N_15423,N_15612);
nor U24091 (N_24091,N_17863,N_15241);
xor U24092 (N_24092,N_16198,N_15106);
or U24093 (N_24093,N_16056,N_16568);
nand U24094 (N_24094,N_15316,N_17320);
nand U24095 (N_24095,N_12975,N_16565);
and U24096 (N_24096,N_13559,N_18051);
and U24097 (N_24097,N_17394,N_13025);
xnor U24098 (N_24098,N_13185,N_13138);
and U24099 (N_24099,N_15195,N_14008);
nor U24100 (N_24100,N_17233,N_14087);
nor U24101 (N_24101,N_12622,N_12964);
xnor U24102 (N_24102,N_18590,N_17805);
and U24103 (N_24103,N_16390,N_18066);
or U24104 (N_24104,N_14228,N_15711);
or U24105 (N_24105,N_18453,N_18181);
nand U24106 (N_24106,N_13792,N_16691);
xor U24107 (N_24107,N_16562,N_14157);
and U24108 (N_24108,N_12604,N_14988);
and U24109 (N_24109,N_14989,N_14964);
and U24110 (N_24110,N_18546,N_16831);
nor U24111 (N_24111,N_12912,N_18380);
xor U24112 (N_24112,N_13333,N_18482);
nor U24113 (N_24113,N_15083,N_18174);
xnor U24114 (N_24114,N_16683,N_16756);
xnor U24115 (N_24115,N_16207,N_13197);
xnor U24116 (N_24116,N_16795,N_16233);
nand U24117 (N_24117,N_14067,N_12555);
nor U24118 (N_24118,N_17902,N_13980);
nor U24119 (N_24119,N_17988,N_16145);
xor U24120 (N_24120,N_15382,N_13552);
nand U24121 (N_24121,N_12848,N_15487);
or U24122 (N_24122,N_15161,N_17801);
nor U24123 (N_24123,N_16709,N_17262);
nand U24124 (N_24124,N_14358,N_15182);
and U24125 (N_24125,N_15218,N_16087);
or U24126 (N_24126,N_14352,N_15317);
or U24127 (N_24127,N_13577,N_13210);
nor U24128 (N_24128,N_17099,N_13007);
nand U24129 (N_24129,N_15195,N_15446);
or U24130 (N_24130,N_16546,N_15344);
xnor U24131 (N_24131,N_13833,N_14549);
and U24132 (N_24132,N_18333,N_13351);
or U24133 (N_24133,N_17761,N_15402);
xnor U24134 (N_24134,N_13056,N_17066);
xor U24135 (N_24135,N_14876,N_14081);
or U24136 (N_24136,N_15897,N_14540);
and U24137 (N_24137,N_13704,N_13755);
and U24138 (N_24138,N_15501,N_18610);
xor U24139 (N_24139,N_14861,N_15011);
nand U24140 (N_24140,N_12549,N_17258);
nor U24141 (N_24141,N_16279,N_16886);
xor U24142 (N_24142,N_14369,N_14179);
nand U24143 (N_24143,N_13786,N_16169);
nor U24144 (N_24144,N_13596,N_16150);
xor U24145 (N_24145,N_16692,N_17025);
xnor U24146 (N_24146,N_13809,N_15402);
nor U24147 (N_24147,N_12694,N_14693);
xnor U24148 (N_24148,N_15467,N_16685);
nor U24149 (N_24149,N_16186,N_15588);
nor U24150 (N_24150,N_18511,N_16157);
nor U24151 (N_24151,N_18509,N_18283);
nor U24152 (N_24152,N_16387,N_13611);
nor U24153 (N_24153,N_13709,N_18221);
and U24154 (N_24154,N_12929,N_17528);
or U24155 (N_24155,N_14142,N_18201);
nor U24156 (N_24156,N_13724,N_17681);
or U24157 (N_24157,N_13754,N_16330);
nand U24158 (N_24158,N_17986,N_16029);
nand U24159 (N_24159,N_17894,N_18344);
nor U24160 (N_24160,N_16061,N_17577);
xnor U24161 (N_24161,N_15051,N_17279);
xor U24162 (N_24162,N_17488,N_17578);
and U24163 (N_24163,N_12724,N_18665);
and U24164 (N_24164,N_15106,N_17933);
nand U24165 (N_24165,N_15582,N_16779);
xnor U24166 (N_24166,N_13113,N_17557);
and U24167 (N_24167,N_17226,N_17000);
and U24168 (N_24168,N_16610,N_13320);
or U24169 (N_24169,N_15448,N_18460);
xnor U24170 (N_24170,N_14637,N_16103);
nand U24171 (N_24171,N_15273,N_12513);
nand U24172 (N_24172,N_17319,N_16427);
xnor U24173 (N_24173,N_17439,N_13174);
xor U24174 (N_24174,N_13605,N_15350);
or U24175 (N_24175,N_14659,N_18527);
and U24176 (N_24176,N_14690,N_13058);
and U24177 (N_24177,N_17233,N_13456);
and U24178 (N_24178,N_17721,N_15457);
nor U24179 (N_24179,N_17945,N_18592);
or U24180 (N_24180,N_14666,N_18642);
xnor U24181 (N_24181,N_12879,N_17109);
nand U24182 (N_24182,N_14012,N_17840);
xnor U24183 (N_24183,N_17388,N_18264);
or U24184 (N_24184,N_18140,N_14820);
and U24185 (N_24185,N_14501,N_15166);
or U24186 (N_24186,N_13982,N_13444);
nand U24187 (N_24187,N_16211,N_17142);
xnor U24188 (N_24188,N_17226,N_18463);
or U24189 (N_24189,N_14976,N_18426);
or U24190 (N_24190,N_15760,N_12704);
or U24191 (N_24191,N_17169,N_13552);
or U24192 (N_24192,N_17616,N_12578);
and U24193 (N_24193,N_14296,N_15009);
nor U24194 (N_24194,N_16451,N_16305);
or U24195 (N_24195,N_14273,N_16839);
or U24196 (N_24196,N_14986,N_17385);
nand U24197 (N_24197,N_15514,N_16800);
nor U24198 (N_24198,N_16544,N_15590);
nand U24199 (N_24199,N_18006,N_16830);
nand U24200 (N_24200,N_14461,N_12599);
and U24201 (N_24201,N_18313,N_18095);
xor U24202 (N_24202,N_13305,N_16781);
nor U24203 (N_24203,N_15167,N_15128);
nor U24204 (N_24204,N_16884,N_13045);
xnor U24205 (N_24205,N_18252,N_15983);
or U24206 (N_24206,N_15952,N_16688);
and U24207 (N_24207,N_18720,N_12714);
and U24208 (N_24208,N_14550,N_14043);
or U24209 (N_24209,N_16059,N_14436);
nand U24210 (N_24210,N_18553,N_17780);
nor U24211 (N_24211,N_16895,N_17093);
nor U24212 (N_24212,N_17532,N_17366);
nand U24213 (N_24213,N_14950,N_13674);
or U24214 (N_24214,N_15382,N_14559);
xnor U24215 (N_24215,N_14507,N_13375);
nand U24216 (N_24216,N_16007,N_15073);
nand U24217 (N_24217,N_13495,N_12675);
nand U24218 (N_24218,N_18620,N_16132);
and U24219 (N_24219,N_16189,N_14734);
xor U24220 (N_24220,N_14206,N_14018);
and U24221 (N_24221,N_12632,N_13582);
xnor U24222 (N_24222,N_15472,N_15646);
nand U24223 (N_24223,N_18461,N_14390);
xnor U24224 (N_24224,N_15884,N_18024);
or U24225 (N_24225,N_18294,N_17350);
xor U24226 (N_24226,N_15643,N_18167);
and U24227 (N_24227,N_17241,N_17523);
xnor U24228 (N_24228,N_13950,N_17996);
or U24229 (N_24229,N_16709,N_17585);
nor U24230 (N_24230,N_12796,N_15899);
xnor U24231 (N_24231,N_16510,N_14703);
nor U24232 (N_24232,N_17095,N_15069);
and U24233 (N_24233,N_13894,N_17375);
nand U24234 (N_24234,N_18560,N_18080);
nor U24235 (N_24235,N_18025,N_14917);
nand U24236 (N_24236,N_16231,N_13310);
or U24237 (N_24237,N_18173,N_16912);
or U24238 (N_24238,N_16519,N_17483);
nand U24239 (N_24239,N_13983,N_17914);
and U24240 (N_24240,N_13243,N_17249);
nand U24241 (N_24241,N_15094,N_15649);
or U24242 (N_24242,N_12849,N_18555);
or U24243 (N_24243,N_16313,N_17878);
or U24244 (N_24244,N_13523,N_15614);
nor U24245 (N_24245,N_18407,N_14540);
nand U24246 (N_24246,N_14943,N_17691);
xnor U24247 (N_24247,N_17336,N_17590);
or U24248 (N_24248,N_16332,N_15755);
nand U24249 (N_24249,N_18718,N_13173);
nor U24250 (N_24250,N_15750,N_13931);
or U24251 (N_24251,N_15352,N_16400);
or U24252 (N_24252,N_13977,N_13938);
and U24253 (N_24253,N_14083,N_14817);
nor U24254 (N_24254,N_13353,N_17492);
nand U24255 (N_24255,N_15927,N_14256);
nand U24256 (N_24256,N_14741,N_13937);
or U24257 (N_24257,N_13405,N_12819);
xor U24258 (N_24258,N_14839,N_17808);
nand U24259 (N_24259,N_16521,N_12732);
and U24260 (N_24260,N_17161,N_15859);
nand U24261 (N_24261,N_17965,N_15769);
or U24262 (N_24262,N_18566,N_17521);
or U24263 (N_24263,N_17393,N_14398);
nand U24264 (N_24264,N_13714,N_14132);
and U24265 (N_24265,N_14921,N_13086);
xor U24266 (N_24266,N_15892,N_15319);
and U24267 (N_24267,N_13722,N_14701);
nand U24268 (N_24268,N_13896,N_16307);
and U24269 (N_24269,N_16532,N_12923);
and U24270 (N_24270,N_14855,N_17329);
nand U24271 (N_24271,N_16057,N_12664);
xor U24272 (N_24272,N_17755,N_15378);
nand U24273 (N_24273,N_16178,N_17331);
and U24274 (N_24274,N_14080,N_17283);
or U24275 (N_24275,N_12600,N_15139);
or U24276 (N_24276,N_16815,N_15832);
xnor U24277 (N_24277,N_16566,N_16403);
or U24278 (N_24278,N_14188,N_15202);
nor U24279 (N_24279,N_16600,N_12779);
xor U24280 (N_24280,N_18135,N_13848);
xor U24281 (N_24281,N_12791,N_18498);
or U24282 (N_24282,N_17124,N_18182);
or U24283 (N_24283,N_17028,N_18593);
nor U24284 (N_24284,N_13713,N_18029);
nand U24285 (N_24285,N_17256,N_15888);
or U24286 (N_24286,N_16088,N_15581);
nand U24287 (N_24287,N_16061,N_13310);
nor U24288 (N_24288,N_14742,N_17861);
and U24289 (N_24289,N_16491,N_15416);
or U24290 (N_24290,N_14461,N_13800);
and U24291 (N_24291,N_15799,N_18292);
and U24292 (N_24292,N_14218,N_12637);
nand U24293 (N_24293,N_15469,N_17667);
and U24294 (N_24294,N_15966,N_17487);
and U24295 (N_24295,N_17803,N_17502);
xnor U24296 (N_24296,N_14264,N_15687);
or U24297 (N_24297,N_15074,N_15554);
xor U24298 (N_24298,N_16257,N_18393);
nor U24299 (N_24299,N_13502,N_18611);
nor U24300 (N_24300,N_13157,N_16363);
nand U24301 (N_24301,N_15285,N_17655);
nand U24302 (N_24302,N_16449,N_15593);
nor U24303 (N_24303,N_15881,N_13069);
xnor U24304 (N_24304,N_14812,N_14261);
nand U24305 (N_24305,N_16237,N_15808);
and U24306 (N_24306,N_18010,N_13114);
and U24307 (N_24307,N_17599,N_14929);
nand U24308 (N_24308,N_16751,N_14678);
and U24309 (N_24309,N_13180,N_17102);
xor U24310 (N_24310,N_13126,N_13954);
and U24311 (N_24311,N_16065,N_17522);
nor U24312 (N_24312,N_14649,N_15094);
or U24313 (N_24313,N_16767,N_13616);
xnor U24314 (N_24314,N_16979,N_13526);
nor U24315 (N_24315,N_16521,N_16536);
or U24316 (N_24316,N_14159,N_15075);
or U24317 (N_24317,N_17373,N_15284);
xor U24318 (N_24318,N_17370,N_14832);
or U24319 (N_24319,N_12659,N_14851);
xor U24320 (N_24320,N_17546,N_17676);
xnor U24321 (N_24321,N_17270,N_12905);
or U24322 (N_24322,N_17208,N_13080);
or U24323 (N_24323,N_16288,N_18140);
nand U24324 (N_24324,N_13626,N_13310);
nand U24325 (N_24325,N_14579,N_12612);
nand U24326 (N_24326,N_14416,N_13961);
or U24327 (N_24327,N_13000,N_16427);
xnor U24328 (N_24328,N_15752,N_15161);
or U24329 (N_24329,N_16617,N_14287);
nor U24330 (N_24330,N_16787,N_17341);
and U24331 (N_24331,N_16096,N_15693);
nor U24332 (N_24332,N_13221,N_15222);
xor U24333 (N_24333,N_18305,N_15500);
nand U24334 (N_24334,N_12792,N_14555);
nand U24335 (N_24335,N_13156,N_13336);
xor U24336 (N_24336,N_15627,N_16704);
or U24337 (N_24337,N_16964,N_16025);
nor U24338 (N_24338,N_12706,N_17675);
nand U24339 (N_24339,N_17487,N_14611);
nand U24340 (N_24340,N_16013,N_16422);
and U24341 (N_24341,N_18528,N_18619);
and U24342 (N_24342,N_14698,N_14540);
nand U24343 (N_24343,N_17660,N_13553);
nand U24344 (N_24344,N_14063,N_12940);
or U24345 (N_24345,N_14074,N_12560);
and U24346 (N_24346,N_16036,N_14353);
nand U24347 (N_24347,N_16407,N_18539);
nand U24348 (N_24348,N_15187,N_17873);
nand U24349 (N_24349,N_13859,N_15174);
or U24350 (N_24350,N_14839,N_15737);
xnor U24351 (N_24351,N_17404,N_18606);
nand U24352 (N_24352,N_14758,N_14021);
or U24353 (N_24353,N_13638,N_17799);
or U24354 (N_24354,N_15685,N_17061);
and U24355 (N_24355,N_12590,N_12635);
and U24356 (N_24356,N_13288,N_18264);
xnor U24357 (N_24357,N_14765,N_15900);
xor U24358 (N_24358,N_17705,N_15930);
nand U24359 (N_24359,N_13983,N_15278);
and U24360 (N_24360,N_13620,N_14048);
or U24361 (N_24361,N_17443,N_15432);
and U24362 (N_24362,N_16039,N_12955);
xnor U24363 (N_24363,N_18687,N_14632);
nand U24364 (N_24364,N_15965,N_18298);
or U24365 (N_24365,N_14176,N_15801);
and U24366 (N_24366,N_16645,N_13649);
nand U24367 (N_24367,N_17815,N_12944);
xor U24368 (N_24368,N_15149,N_16511);
nand U24369 (N_24369,N_16730,N_15668);
or U24370 (N_24370,N_12730,N_18474);
xnor U24371 (N_24371,N_12813,N_13290);
and U24372 (N_24372,N_16142,N_18024);
nor U24373 (N_24373,N_17951,N_17064);
or U24374 (N_24374,N_16397,N_16322);
xnor U24375 (N_24375,N_14286,N_13264);
nor U24376 (N_24376,N_14804,N_17293);
nand U24377 (N_24377,N_17163,N_14059);
nand U24378 (N_24378,N_13515,N_17190);
nor U24379 (N_24379,N_15280,N_15673);
and U24380 (N_24380,N_17415,N_16893);
nand U24381 (N_24381,N_15353,N_12957);
or U24382 (N_24382,N_14158,N_13962);
or U24383 (N_24383,N_16732,N_15995);
nand U24384 (N_24384,N_12896,N_12955);
and U24385 (N_24385,N_16295,N_12821);
xnor U24386 (N_24386,N_16896,N_17266);
xor U24387 (N_24387,N_15396,N_17657);
nand U24388 (N_24388,N_16204,N_16031);
nand U24389 (N_24389,N_18594,N_15830);
nor U24390 (N_24390,N_18637,N_18044);
xor U24391 (N_24391,N_13199,N_13950);
xnor U24392 (N_24392,N_12659,N_16161);
nor U24393 (N_24393,N_15624,N_17011);
or U24394 (N_24394,N_13192,N_12756);
or U24395 (N_24395,N_12897,N_14798);
or U24396 (N_24396,N_18582,N_16671);
or U24397 (N_24397,N_17053,N_14707);
xor U24398 (N_24398,N_18175,N_16979);
or U24399 (N_24399,N_14697,N_12659);
nor U24400 (N_24400,N_17221,N_14694);
xor U24401 (N_24401,N_15247,N_15952);
and U24402 (N_24402,N_13826,N_16304);
xor U24403 (N_24403,N_14539,N_17569);
nor U24404 (N_24404,N_12879,N_16683);
nand U24405 (N_24405,N_14259,N_14651);
and U24406 (N_24406,N_13556,N_18027);
and U24407 (N_24407,N_14251,N_16548);
and U24408 (N_24408,N_13828,N_16797);
and U24409 (N_24409,N_18075,N_13076);
and U24410 (N_24410,N_14219,N_13286);
xor U24411 (N_24411,N_13605,N_17766);
xnor U24412 (N_24412,N_13173,N_13661);
nand U24413 (N_24413,N_13615,N_17492);
or U24414 (N_24414,N_13521,N_17472);
nand U24415 (N_24415,N_13743,N_17510);
and U24416 (N_24416,N_12533,N_16587);
nor U24417 (N_24417,N_15425,N_14771);
or U24418 (N_24418,N_14618,N_16873);
nor U24419 (N_24419,N_14079,N_14516);
nor U24420 (N_24420,N_15243,N_13896);
or U24421 (N_24421,N_17774,N_13706);
nor U24422 (N_24422,N_15957,N_17858);
or U24423 (N_24423,N_16807,N_13982);
nand U24424 (N_24424,N_13556,N_12907);
nand U24425 (N_24425,N_12633,N_14239);
nand U24426 (N_24426,N_15339,N_16275);
nand U24427 (N_24427,N_16959,N_17880);
nand U24428 (N_24428,N_18716,N_15007);
xor U24429 (N_24429,N_18471,N_16746);
xor U24430 (N_24430,N_14713,N_13949);
and U24431 (N_24431,N_13579,N_17660);
or U24432 (N_24432,N_15335,N_15342);
and U24433 (N_24433,N_17058,N_18504);
nand U24434 (N_24434,N_15191,N_13220);
xor U24435 (N_24435,N_13230,N_15315);
nand U24436 (N_24436,N_17469,N_14945);
nand U24437 (N_24437,N_16507,N_12907);
and U24438 (N_24438,N_13715,N_16233);
xor U24439 (N_24439,N_18585,N_15417);
or U24440 (N_24440,N_12919,N_13314);
xnor U24441 (N_24441,N_14148,N_18125);
or U24442 (N_24442,N_16989,N_16874);
nand U24443 (N_24443,N_12883,N_13084);
xnor U24444 (N_24444,N_16040,N_15929);
and U24445 (N_24445,N_16999,N_17637);
xor U24446 (N_24446,N_13881,N_13496);
or U24447 (N_24447,N_15628,N_15345);
nand U24448 (N_24448,N_14458,N_15434);
or U24449 (N_24449,N_15522,N_15831);
xor U24450 (N_24450,N_16448,N_17014);
nand U24451 (N_24451,N_12911,N_18534);
nand U24452 (N_24452,N_13399,N_16358);
or U24453 (N_24453,N_17946,N_15140);
nand U24454 (N_24454,N_12812,N_18302);
and U24455 (N_24455,N_13759,N_17835);
xor U24456 (N_24456,N_13605,N_15605);
or U24457 (N_24457,N_14240,N_14298);
or U24458 (N_24458,N_15032,N_15311);
and U24459 (N_24459,N_12732,N_17848);
nor U24460 (N_24460,N_17686,N_18091);
and U24461 (N_24461,N_15691,N_17573);
or U24462 (N_24462,N_17931,N_13102);
and U24463 (N_24463,N_15602,N_16046);
nor U24464 (N_24464,N_12697,N_16947);
nor U24465 (N_24465,N_15276,N_17813);
nor U24466 (N_24466,N_18054,N_17384);
nor U24467 (N_24467,N_17495,N_13858);
xnor U24468 (N_24468,N_17415,N_17119);
xnor U24469 (N_24469,N_16422,N_17642);
nand U24470 (N_24470,N_16252,N_16264);
nand U24471 (N_24471,N_13440,N_15512);
nor U24472 (N_24472,N_12914,N_15272);
and U24473 (N_24473,N_14576,N_13883);
and U24474 (N_24474,N_12519,N_15612);
xor U24475 (N_24475,N_13368,N_15529);
nor U24476 (N_24476,N_18166,N_15047);
nand U24477 (N_24477,N_13734,N_13368);
xnor U24478 (N_24478,N_12632,N_13192);
or U24479 (N_24479,N_12909,N_17906);
xnor U24480 (N_24480,N_13325,N_14334);
or U24481 (N_24481,N_14272,N_13117);
or U24482 (N_24482,N_14198,N_15962);
nor U24483 (N_24483,N_16157,N_13133);
nor U24484 (N_24484,N_18563,N_13410);
nor U24485 (N_24485,N_18309,N_13682);
nand U24486 (N_24486,N_16941,N_17351);
and U24487 (N_24487,N_14861,N_18631);
xnor U24488 (N_24488,N_13895,N_16336);
nand U24489 (N_24489,N_14814,N_18652);
and U24490 (N_24490,N_13324,N_12881);
nor U24491 (N_24491,N_13843,N_16235);
nor U24492 (N_24492,N_15379,N_17146);
nand U24493 (N_24493,N_17985,N_15902);
or U24494 (N_24494,N_13368,N_15376);
nor U24495 (N_24495,N_12937,N_15012);
nor U24496 (N_24496,N_13969,N_15867);
xnor U24497 (N_24497,N_15218,N_16838);
and U24498 (N_24498,N_14513,N_18352);
nor U24499 (N_24499,N_17904,N_17008);
xor U24500 (N_24500,N_16698,N_15730);
or U24501 (N_24501,N_14280,N_14626);
and U24502 (N_24502,N_15584,N_13685);
nor U24503 (N_24503,N_16237,N_18156);
xnor U24504 (N_24504,N_15439,N_18170);
or U24505 (N_24505,N_12607,N_12602);
nor U24506 (N_24506,N_12747,N_15775);
and U24507 (N_24507,N_15055,N_18640);
nand U24508 (N_24508,N_18210,N_17816);
nor U24509 (N_24509,N_17778,N_12643);
nand U24510 (N_24510,N_14181,N_17438);
xor U24511 (N_24511,N_12771,N_16816);
and U24512 (N_24512,N_14285,N_14808);
nor U24513 (N_24513,N_18222,N_13934);
xor U24514 (N_24514,N_16046,N_18292);
and U24515 (N_24515,N_15520,N_17713);
nand U24516 (N_24516,N_12722,N_12777);
or U24517 (N_24517,N_13033,N_16605);
nor U24518 (N_24518,N_14419,N_16179);
or U24519 (N_24519,N_13374,N_13528);
nand U24520 (N_24520,N_17659,N_18403);
and U24521 (N_24521,N_16592,N_16115);
or U24522 (N_24522,N_15886,N_18651);
xor U24523 (N_24523,N_16219,N_13958);
nor U24524 (N_24524,N_16545,N_13992);
or U24525 (N_24525,N_14372,N_16767);
nand U24526 (N_24526,N_16984,N_14927);
or U24527 (N_24527,N_13990,N_17371);
xor U24528 (N_24528,N_17046,N_12715);
or U24529 (N_24529,N_17116,N_14537);
nand U24530 (N_24530,N_13690,N_17109);
xor U24531 (N_24531,N_12575,N_12706);
nor U24532 (N_24532,N_12552,N_16841);
nand U24533 (N_24533,N_14812,N_15676);
and U24534 (N_24534,N_17812,N_14988);
nand U24535 (N_24535,N_16925,N_16739);
nand U24536 (N_24536,N_12587,N_17776);
nor U24537 (N_24537,N_17122,N_14759);
xor U24538 (N_24538,N_15156,N_15669);
or U24539 (N_24539,N_14176,N_15273);
nand U24540 (N_24540,N_17095,N_13154);
or U24541 (N_24541,N_15280,N_12962);
or U24542 (N_24542,N_14919,N_15809);
nand U24543 (N_24543,N_15391,N_14893);
and U24544 (N_24544,N_13006,N_12655);
xor U24545 (N_24545,N_17094,N_16633);
xnor U24546 (N_24546,N_17539,N_17669);
and U24547 (N_24547,N_14724,N_16997);
nand U24548 (N_24548,N_15266,N_15868);
xnor U24549 (N_24549,N_13828,N_17615);
nand U24550 (N_24550,N_17577,N_16894);
xnor U24551 (N_24551,N_12729,N_17750);
nand U24552 (N_24552,N_18741,N_13676);
and U24553 (N_24553,N_13214,N_15708);
nand U24554 (N_24554,N_16362,N_17418);
nand U24555 (N_24555,N_18566,N_16826);
nor U24556 (N_24556,N_14135,N_15051);
xnor U24557 (N_24557,N_12927,N_16518);
or U24558 (N_24558,N_12976,N_14153);
nand U24559 (N_24559,N_16141,N_12904);
or U24560 (N_24560,N_13291,N_15886);
nor U24561 (N_24561,N_16011,N_12896);
nand U24562 (N_24562,N_15370,N_14563);
or U24563 (N_24563,N_17415,N_15190);
xnor U24564 (N_24564,N_17778,N_15749);
nor U24565 (N_24565,N_12718,N_17618);
nor U24566 (N_24566,N_13905,N_15487);
or U24567 (N_24567,N_18669,N_13111);
xor U24568 (N_24568,N_13490,N_14225);
xnor U24569 (N_24569,N_14438,N_14740);
xnor U24570 (N_24570,N_16255,N_16675);
nand U24571 (N_24571,N_13523,N_18441);
nor U24572 (N_24572,N_16122,N_16112);
xnor U24573 (N_24573,N_13440,N_18619);
nand U24574 (N_24574,N_18288,N_18477);
nand U24575 (N_24575,N_17595,N_13955);
or U24576 (N_24576,N_12735,N_13192);
xnor U24577 (N_24577,N_17759,N_16586);
xnor U24578 (N_24578,N_13832,N_17021);
and U24579 (N_24579,N_14155,N_16361);
and U24580 (N_24580,N_15807,N_15594);
nand U24581 (N_24581,N_13899,N_17801);
or U24582 (N_24582,N_15296,N_16847);
or U24583 (N_24583,N_15491,N_17654);
nand U24584 (N_24584,N_17720,N_17000);
xnor U24585 (N_24585,N_16401,N_15786);
and U24586 (N_24586,N_18730,N_13017);
nor U24587 (N_24587,N_15553,N_16978);
xnor U24588 (N_24588,N_17961,N_15644);
nand U24589 (N_24589,N_17412,N_13128);
nor U24590 (N_24590,N_16920,N_15319);
xor U24591 (N_24591,N_18742,N_15872);
or U24592 (N_24592,N_15592,N_15806);
or U24593 (N_24593,N_17973,N_12641);
or U24594 (N_24594,N_17818,N_18640);
or U24595 (N_24595,N_13447,N_17033);
and U24596 (N_24596,N_14743,N_13088);
or U24597 (N_24597,N_18402,N_15478);
and U24598 (N_24598,N_12981,N_12567);
nand U24599 (N_24599,N_16041,N_13914);
or U24600 (N_24600,N_12714,N_14585);
nor U24601 (N_24601,N_15232,N_15473);
nand U24602 (N_24602,N_14099,N_15446);
nor U24603 (N_24603,N_15165,N_14212);
nor U24604 (N_24604,N_18426,N_14640);
nor U24605 (N_24605,N_18169,N_15947);
xor U24606 (N_24606,N_16452,N_16178);
or U24607 (N_24607,N_15791,N_13618);
and U24608 (N_24608,N_13601,N_14257);
nand U24609 (N_24609,N_16804,N_17869);
nand U24610 (N_24610,N_13166,N_17297);
xnor U24611 (N_24611,N_14654,N_16914);
nand U24612 (N_24612,N_15274,N_17923);
nand U24613 (N_24613,N_14313,N_18616);
and U24614 (N_24614,N_14433,N_18321);
or U24615 (N_24615,N_16654,N_18228);
nor U24616 (N_24616,N_16885,N_15424);
or U24617 (N_24617,N_18301,N_18563);
nor U24618 (N_24618,N_15245,N_18310);
and U24619 (N_24619,N_12683,N_13843);
or U24620 (N_24620,N_15571,N_16574);
or U24621 (N_24621,N_16378,N_14897);
and U24622 (N_24622,N_16181,N_16937);
or U24623 (N_24623,N_13656,N_15399);
nand U24624 (N_24624,N_17194,N_13323);
or U24625 (N_24625,N_14464,N_17048);
xnor U24626 (N_24626,N_17827,N_17092);
nand U24627 (N_24627,N_16895,N_16425);
xor U24628 (N_24628,N_15360,N_17743);
nand U24629 (N_24629,N_16549,N_14469);
and U24630 (N_24630,N_17927,N_12630);
nor U24631 (N_24631,N_17952,N_15242);
nor U24632 (N_24632,N_15830,N_14429);
or U24633 (N_24633,N_15983,N_14595);
nor U24634 (N_24634,N_13448,N_16058);
xor U24635 (N_24635,N_15320,N_14995);
and U24636 (N_24636,N_13298,N_13235);
nand U24637 (N_24637,N_12883,N_12532);
nand U24638 (N_24638,N_12521,N_13125);
nand U24639 (N_24639,N_17385,N_18512);
and U24640 (N_24640,N_17786,N_13994);
nand U24641 (N_24641,N_18086,N_12562);
nor U24642 (N_24642,N_12534,N_17504);
nor U24643 (N_24643,N_15774,N_12869);
xnor U24644 (N_24644,N_15286,N_17125);
xnor U24645 (N_24645,N_14114,N_16197);
nor U24646 (N_24646,N_16106,N_18190);
xnor U24647 (N_24647,N_15926,N_14043);
nor U24648 (N_24648,N_15972,N_15019);
xor U24649 (N_24649,N_12670,N_17962);
and U24650 (N_24650,N_18160,N_14958);
and U24651 (N_24651,N_17880,N_15653);
and U24652 (N_24652,N_17858,N_18170);
or U24653 (N_24653,N_14886,N_17234);
and U24654 (N_24654,N_17835,N_15624);
nand U24655 (N_24655,N_17237,N_17399);
nand U24656 (N_24656,N_14877,N_17739);
and U24657 (N_24657,N_14850,N_14042);
xor U24658 (N_24658,N_18745,N_15399);
nor U24659 (N_24659,N_15272,N_16795);
nand U24660 (N_24660,N_16863,N_13229);
xnor U24661 (N_24661,N_16748,N_14189);
nand U24662 (N_24662,N_18193,N_16793);
and U24663 (N_24663,N_12784,N_18703);
nor U24664 (N_24664,N_18369,N_18715);
nor U24665 (N_24665,N_16919,N_16830);
nor U24666 (N_24666,N_18176,N_15038);
nand U24667 (N_24667,N_18118,N_14353);
or U24668 (N_24668,N_13230,N_17067);
or U24669 (N_24669,N_14094,N_16717);
xor U24670 (N_24670,N_15561,N_14136);
and U24671 (N_24671,N_16753,N_17274);
or U24672 (N_24672,N_13527,N_16810);
xor U24673 (N_24673,N_17632,N_17124);
xor U24674 (N_24674,N_16213,N_16469);
and U24675 (N_24675,N_17041,N_14516);
xor U24676 (N_24676,N_15428,N_18703);
and U24677 (N_24677,N_16407,N_13029);
nand U24678 (N_24678,N_18152,N_17621);
nor U24679 (N_24679,N_13652,N_14243);
or U24680 (N_24680,N_17178,N_17961);
xnor U24681 (N_24681,N_18134,N_15994);
and U24682 (N_24682,N_17674,N_15219);
or U24683 (N_24683,N_12952,N_18018);
nor U24684 (N_24684,N_14127,N_16072);
or U24685 (N_24685,N_15300,N_18713);
and U24686 (N_24686,N_14814,N_13676);
nand U24687 (N_24687,N_13427,N_17361);
and U24688 (N_24688,N_16626,N_18718);
or U24689 (N_24689,N_13216,N_14988);
or U24690 (N_24690,N_17980,N_17348);
nand U24691 (N_24691,N_13479,N_17032);
or U24692 (N_24692,N_13910,N_18749);
and U24693 (N_24693,N_15261,N_13952);
nor U24694 (N_24694,N_16617,N_15016);
xor U24695 (N_24695,N_12670,N_16772);
nor U24696 (N_24696,N_13714,N_16229);
xnor U24697 (N_24697,N_17682,N_13255);
or U24698 (N_24698,N_17316,N_16728);
and U24699 (N_24699,N_15007,N_12643);
nor U24700 (N_24700,N_15861,N_15928);
nor U24701 (N_24701,N_18204,N_13284);
nor U24702 (N_24702,N_16611,N_17394);
xnor U24703 (N_24703,N_18391,N_15739);
and U24704 (N_24704,N_16782,N_13573);
or U24705 (N_24705,N_14899,N_16629);
nor U24706 (N_24706,N_17615,N_17844);
xnor U24707 (N_24707,N_14607,N_17825);
or U24708 (N_24708,N_18509,N_13153);
and U24709 (N_24709,N_17313,N_16387);
nand U24710 (N_24710,N_15857,N_16634);
xnor U24711 (N_24711,N_15708,N_16364);
nand U24712 (N_24712,N_14183,N_14617);
nor U24713 (N_24713,N_16972,N_12710);
nor U24714 (N_24714,N_13545,N_17679);
xnor U24715 (N_24715,N_14719,N_14754);
nor U24716 (N_24716,N_14116,N_15917);
nor U24717 (N_24717,N_14069,N_13322);
nand U24718 (N_24718,N_14822,N_16431);
or U24719 (N_24719,N_16819,N_15430);
and U24720 (N_24720,N_13547,N_16955);
and U24721 (N_24721,N_18592,N_16924);
xnor U24722 (N_24722,N_16175,N_14046);
xor U24723 (N_24723,N_13014,N_17639);
or U24724 (N_24724,N_12634,N_16830);
and U24725 (N_24725,N_12719,N_13683);
nand U24726 (N_24726,N_15555,N_13545);
nand U24727 (N_24727,N_18219,N_17709);
or U24728 (N_24728,N_14584,N_18727);
nor U24729 (N_24729,N_16181,N_12722);
nand U24730 (N_24730,N_13122,N_17538);
nand U24731 (N_24731,N_15562,N_15167);
or U24732 (N_24732,N_17902,N_13351);
xor U24733 (N_24733,N_18710,N_15068);
or U24734 (N_24734,N_17425,N_16221);
and U24735 (N_24735,N_15321,N_16493);
or U24736 (N_24736,N_18546,N_13650);
or U24737 (N_24737,N_13050,N_18710);
or U24738 (N_24738,N_15469,N_16019);
nor U24739 (N_24739,N_13946,N_16896);
nand U24740 (N_24740,N_15500,N_17747);
and U24741 (N_24741,N_12572,N_15280);
xnor U24742 (N_24742,N_13755,N_17740);
or U24743 (N_24743,N_17768,N_13618);
nor U24744 (N_24744,N_13386,N_13102);
xnor U24745 (N_24745,N_15111,N_12843);
nand U24746 (N_24746,N_14725,N_13038);
or U24747 (N_24747,N_14557,N_14129);
xor U24748 (N_24748,N_17153,N_16526);
or U24749 (N_24749,N_17696,N_18703);
xor U24750 (N_24750,N_13766,N_14083);
nor U24751 (N_24751,N_14087,N_14343);
xor U24752 (N_24752,N_17201,N_15262);
nand U24753 (N_24753,N_16899,N_15293);
and U24754 (N_24754,N_16010,N_13613);
xnor U24755 (N_24755,N_14752,N_13056);
nor U24756 (N_24756,N_16425,N_18681);
or U24757 (N_24757,N_17707,N_18583);
nor U24758 (N_24758,N_17844,N_13676);
or U24759 (N_24759,N_12808,N_14310);
and U24760 (N_24760,N_16733,N_12947);
nand U24761 (N_24761,N_13732,N_13862);
xor U24762 (N_24762,N_16380,N_18168);
and U24763 (N_24763,N_13100,N_15590);
nand U24764 (N_24764,N_14200,N_14823);
nand U24765 (N_24765,N_17977,N_14721);
nor U24766 (N_24766,N_14520,N_14085);
or U24767 (N_24767,N_16622,N_17861);
nor U24768 (N_24768,N_14752,N_17390);
nor U24769 (N_24769,N_13257,N_16354);
nand U24770 (N_24770,N_15489,N_16102);
nor U24771 (N_24771,N_14116,N_15322);
xor U24772 (N_24772,N_16048,N_16025);
nor U24773 (N_24773,N_18652,N_17681);
xnor U24774 (N_24774,N_13780,N_16125);
or U24775 (N_24775,N_15316,N_18270);
nor U24776 (N_24776,N_13726,N_16538);
and U24777 (N_24777,N_14956,N_15162);
nor U24778 (N_24778,N_17143,N_14699);
or U24779 (N_24779,N_18279,N_17260);
or U24780 (N_24780,N_15156,N_14974);
xnor U24781 (N_24781,N_17024,N_13089);
nand U24782 (N_24782,N_18624,N_18348);
xor U24783 (N_24783,N_14148,N_16749);
and U24784 (N_24784,N_16853,N_14563);
and U24785 (N_24785,N_17052,N_14770);
nand U24786 (N_24786,N_17838,N_14055);
xor U24787 (N_24787,N_14641,N_17924);
or U24788 (N_24788,N_18057,N_18008);
nor U24789 (N_24789,N_16190,N_13432);
nand U24790 (N_24790,N_15581,N_13112);
nand U24791 (N_24791,N_14065,N_17117);
or U24792 (N_24792,N_16025,N_17461);
xor U24793 (N_24793,N_13425,N_14614);
and U24794 (N_24794,N_14859,N_14853);
or U24795 (N_24795,N_17915,N_16575);
nand U24796 (N_24796,N_18346,N_16970);
or U24797 (N_24797,N_18353,N_12981);
nand U24798 (N_24798,N_13030,N_15440);
and U24799 (N_24799,N_15101,N_16659);
or U24800 (N_24800,N_17030,N_14826);
or U24801 (N_24801,N_15216,N_14063);
or U24802 (N_24802,N_17872,N_18413);
nand U24803 (N_24803,N_14315,N_14394);
nand U24804 (N_24804,N_13552,N_16206);
or U24805 (N_24805,N_12710,N_13219);
or U24806 (N_24806,N_15098,N_14909);
or U24807 (N_24807,N_16243,N_14034);
nand U24808 (N_24808,N_13360,N_15351);
and U24809 (N_24809,N_16107,N_16674);
nor U24810 (N_24810,N_14206,N_16249);
nand U24811 (N_24811,N_14789,N_14095);
nor U24812 (N_24812,N_14263,N_17211);
and U24813 (N_24813,N_17574,N_16193);
and U24814 (N_24814,N_12764,N_13541);
nor U24815 (N_24815,N_18432,N_17049);
or U24816 (N_24816,N_13456,N_13104);
or U24817 (N_24817,N_15718,N_16693);
nor U24818 (N_24818,N_18112,N_13298);
and U24819 (N_24819,N_13921,N_13264);
xnor U24820 (N_24820,N_14796,N_17421);
xnor U24821 (N_24821,N_17514,N_15765);
nor U24822 (N_24822,N_16884,N_16913);
and U24823 (N_24823,N_16300,N_12726);
nor U24824 (N_24824,N_16932,N_15461);
or U24825 (N_24825,N_16674,N_18629);
nor U24826 (N_24826,N_18469,N_13206);
and U24827 (N_24827,N_17694,N_16407);
xnor U24828 (N_24828,N_17888,N_18207);
and U24829 (N_24829,N_17677,N_14570);
nor U24830 (N_24830,N_16696,N_13824);
and U24831 (N_24831,N_18541,N_14468);
and U24832 (N_24832,N_15604,N_18236);
nand U24833 (N_24833,N_16413,N_17142);
and U24834 (N_24834,N_17287,N_16343);
nand U24835 (N_24835,N_18736,N_15411);
xor U24836 (N_24836,N_18489,N_14506);
xnor U24837 (N_24837,N_17593,N_15367);
and U24838 (N_24838,N_14442,N_14680);
nand U24839 (N_24839,N_13127,N_17623);
nand U24840 (N_24840,N_16569,N_15107);
xor U24841 (N_24841,N_13798,N_17745);
nand U24842 (N_24842,N_14765,N_14881);
or U24843 (N_24843,N_15293,N_15245);
or U24844 (N_24844,N_14573,N_14585);
nor U24845 (N_24845,N_18488,N_17720);
and U24846 (N_24846,N_16300,N_16050);
or U24847 (N_24847,N_17327,N_14280);
and U24848 (N_24848,N_18069,N_14655);
nand U24849 (N_24849,N_15245,N_18047);
nor U24850 (N_24850,N_14272,N_18635);
and U24851 (N_24851,N_17809,N_14418);
or U24852 (N_24852,N_14185,N_15676);
and U24853 (N_24853,N_15622,N_13865);
or U24854 (N_24854,N_14035,N_16316);
nor U24855 (N_24855,N_17219,N_13614);
nor U24856 (N_24856,N_13192,N_15715);
or U24857 (N_24857,N_12648,N_15243);
xnor U24858 (N_24858,N_17232,N_13364);
nor U24859 (N_24859,N_13089,N_17581);
and U24860 (N_24860,N_12861,N_16574);
xor U24861 (N_24861,N_16419,N_18675);
xnor U24862 (N_24862,N_13185,N_17450);
nor U24863 (N_24863,N_18569,N_13595);
nor U24864 (N_24864,N_18166,N_18211);
nand U24865 (N_24865,N_17585,N_17714);
and U24866 (N_24866,N_17222,N_13303);
nor U24867 (N_24867,N_14620,N_15762);
xnor U24868 (N_24868,N_14964,N_18123);
xnor U24869 (N_24869,N_13160,N_16676);
xor U24870 (N_24870,N_12562,N_13367);
and U24871 (N_24871,N_18724,N_17630);
or U24872 (N_24872,N_16124,N_15229);
nand U24873 (N_24873,N_14153,N_17558);
xnor U24874 (N_24874,N_16226,N_15932);
or U24875 (N_24875,N_16276,N_14597);
nor U24876 (N_24876,N_17312,N_15717);
nand U24877 (N_24877,N_15141,N_12802);
nor U24878 (N_24878,N_14192,N_12871);
nand U24879 (N_24879,N_14933,N_15261);
nor U24880 (N_24880,N_18388,N_15028);
nand U24881 (N_24881,N_14034,N_17902);
nor U24882 (N_24882,N_16142,N_16858);
and U24883 (N_24883,N_14427,N_13271);
and U24884 (N_24884,N_16719,N_16734);
or U24885 (N_24885,N_16774,N_13635);
or U24886 (N_24886,N_13857,N_15381);
nand U24887 (N_24887,N_15655,N_15992);
nand U24888 (N_24888,N_13247,N_16458);
or U24889 (N_24889,N_13099,N_18685);
xor U24890 (N_24890,N_12618,N_14530);
and U24891 (N_24891,N_17816,N_17430);
nand U24892 (N_24892,N_12704,N_16090);
and U24893 (N_24893,N_16772,N_13424);
and U24894 (N_24894,N_13775,N_13566);
nand U24895 (N_24895,N_17777,N_13776);
nor U24896 (N_24896,N_15930,N_17410);
nand U24897 (N_24897,N_13214,N_17607);
nand U24898 (N_24898,N_13179,N_17841);
or U24899 (N_24899,N_13357,N_16632);
xor U24900 (N_24900,N_18402,N_15936);
nor U24901 (N_24901,N_13525,N_16896);
xor U24902 (N_24902,N_13045,N_13003);
or U24903 (N_24903,N_18545,N_13117);
or U24904 (N_24904,N_13397,N_14302);
and U24905 (N_24905,N_13304,N_17353);
or U24906 (N_24906,N_14437,N_13571);
and U24907 (N_24907,N_16225,N_14478);
xnor U24908 (N_24908,N_13182,N_17744);
and U24909 (N_24909,N_13041,N_18337);
nand U24910 (N_24910,N_13862,N_14728);
and U24911 (N_24911,N_13450,N_14461);
nand U24912 (N_24912,N_12544,N_18666);
nand U24913 (N_24913,N_15524,N_17919);
nand U24914 (N_24914,N_15920,N_13574);
xnor U24915 (N_24915,N_15271,N_15913);
or U24916 (N_24916,N_16336,N_15567);
nand U24917 (N_24917,N_12964,N_17164);
or U24918 (N_24918,N_13454,N_15780);
nor U24919 (N_24919,N_17921,N_17140);
or U24920 (N_24920,N_16760,N_18567);
xnor U24921 (N_24921,N_12896,N_12693);
and U24922 (N_24922,N_16950,N_13375);
nor U24923 (N_24923,N_15610,N_18734);
xnor U24924 (N_24924,N_17921,N_12562);
xor U24925 (N_24925,N_15588,N_12792);
and U24926 (N_24926,N_14778,N_18176);
xnor U24927 (N_24927,N_12705,N_13566);
nor U24928 (N_24928,N_17485,N_14537);
nor U24929 (N_24929,N_16660,N_13564);
nand U24930 (N_24930,N_13982,N_15728);
nor U24931 (N_24931,N_17286,N_15270);
or U24932 (N_24932,N_14323,N_14523);
nand U24933 (N_24933,N_16925,N_15243);
and U24934 (N_24934,N_16118,N_18088);
nand U24935 (N_24935,N_12560,N_17141);
nor U24936 (N_24936,N_13863,N_16945);
or U24937 (N_24937,N_14657,N_18552);
nor U24938 (N_24938,N_13703,N_15580);
nor U24939 (N_24939,N_18007,N_17208);
nor U24940 (N_24940,N_18709,N_13250);
or U24941 (N_24941,N_18590,N_12684);
and U24942 (N_24942,N_17029,N_13067);
xnor U24943 (N_24943,N_17134,N_17578);
and U24944 (N_24944,N_13236,N_16530);
or U24945 (N_24945,N_17224,N_16212);
nand U24946 (N_24946,N_18658,N_13221);
nor U24947 (N_24947,N_12604,N_13001);
nor U24948 (N_24948,N_13556,N_16486);
and U24949 (N_24949,N_13409,N_14885);
nand U24950 (N_24950,N_14695,N_12665);
nor U24951 (N_24951,N_18528,N_17464);
or U24952 (N_24952,N_16311,N_14007);
or U24953 (N_24953,N_15178,N_14593);
nand U24954 (N_24954,N_12992,N_16771);
or U24955 (N_24955,N_13197,N_15357);
and U24956 (N_24956,N_17659,N_15324);
xor U24957 (N_24957,N_17970,N_17740);
and U24958 (N_24958,N_16376,N_15671);
nor U24959 (N_24959,N_13334,N_15906);
or U24960 (N_24960,N_17410,N_17045);
and U24961 (N_24961,N_14536,N_12970);
nor U24962 (N_24962,N_17152,N_18022);
nor U24963 (N_24963,N_16795,N_17571);
and U24964 (N_24964,N_12941,N_12581);
and U24965 (N_24965,N_15447,N_15520);
and U24966 (N_24966,N_12998,N_18532);
nand U24967 (N_24967,N_16172,N_13267);
and U24968 (N_24968,N_16561,N_13708);
xor U24969 (N_24969,N_12552,N_18114);
nand U24970 (N_24970,N_14668,N_15922);
or U24971 (N_24971,N_17379,N_13204);
or U24972 (N_24972,N_14336,N_14642);
and U24973 (N_24973,N_16750,N_17891);
nor U24974 (N_24974,N_15841,N_14325);
nor U24975 (N_24975,N_15607,N_16157);
nand U24976 (N_24976,N_14775,N_14316);
or U24977 (N_24977,N_15354,N_15408);
and U24978 (N_24978,N_14934,N_14124);
nand U24979 (N_24979,N_17878,N_16867);
and U24980 (N_24980,N_15448,N_15336);
xnor U24981 (N_24981,N_17771,N_15465);
and U24982 (N_24982,N_13125,N_16353);
or U24983 (N_24983,N_16406,N_12609);
xor U24984 (N_24984,N_15982,N_13446);
or U24985 (N_24985,N_12842,N_15034);
nor U24986 (N_24986,N_14456,N_15707);
and U24987 (N_24987,N_18618,N_15606);
and U24988 (N_24988,N_14516,N_16102);
nand U24989 (N_24989,N_13868,N_14246);
or U24990 (N_24990,N_16386,N_18598);
nor U24991 (N_24991,N_12921,N_15756);
nand U24992 (N_24992,N_17797,N_12738);
and U24993 (N_24993,N_13260,N_15813);
and U24994 (N_24994,N_18354,N_13404);
xor U24995 (N_24995,N_14379,N_14995);
or U24996 (N_24996,N_14004,N_13517);
nor U24997 (N_24997,N_13202,N_12527);
nor U24998 (N_24998,N_18441,N_14386);
and U24999 (N_24999,N_12588,N_15305);
nor UO_0 (O_0,N_20251,N_24348);
nand UO_1 (O_1,N_24240,N_20809);
nand UO_2 (O_2,N_24826,N_24782);
or UO_3 (O_3,N_19286,N_21863);
nand UO_4 (O_4,N_21211,N_20403);
nand UO_5 (O_5,N_22639,N_20061);
xnor UO_6 (O_6,N_20115,N_24101);
nand UO_7 (O_7,N_22042,N_23077);
xor UO_8 (O_8,N_22521,N_22400);
or UO_9 (O_9,N_19832,N_22920);
or UO_10 (O_10,N_24688,N_22231);
and UO_11 (O_11,N_23170,N_21970);
nand UO_12 (O_12,N_24349,N_21719);
nand UO_13 (O_13,N_21157,N_21770);
or UO_14 (O_14,N_22543,N_21916);
and UO_15 (O_15,N_22898,N_23877);
or UO_16 (O_16,N_21800,N_21897);
nor UO_17 (O_17,N_22754,N_18868);
nand UO_18 (O_18,N_19483,N_20461);
xor UO_19 (O_19,N_24104,N_19028);
and UO_20 (O_20,N_23564,N_23349);
nor UO_21 (O_21,N_20959,N_18968);
or UO_22 (O_22,N_21163,N_22383);
and UO_23 (O_23,N_21330,N_23034);
or UO_24 (O_24,N_21316,N_21373);
and UO_25 (O_25,N_23626,N_21969);
and UO_26 (O_26,N_20122,N_23152);
nor UO_27 (O_27,N_21956,N_21248);
or UO_28 (O_28,N_23722,N_24951);
nand UO_29 (O_29,N_24062,N_19271);
or UO_30 (O_30,N_19632,N_21574);
xor UO_31 (O_31,N_19743,N_24004);
and UO_32 (O_32,N_21007,N_22725);
xor UO_33 (O_33,N_24265,N_23359);
or UO_34 (O_34,N_20968,N_23772);
nor UO_35 (O_35,N_20368,N_23389);
or UO_36 (O_36,N_18785,N_22313);
or UO_37 (O_37,N_22593,N_19659);
nand UO_38 (O_38,N_19046,N_20041);
nand UO_39 (O_39,N_24996,N_24135);
nor UO_40 (O_40,N_23577,N_22923);
xnor UO_41 (O_41,N_21277,N_23076);
nor UO_42 (O_42,N_21059,N_24868);
nor UO_43 (O_43,N_24865,N_24791);
nor UO_44 (O_44,N_23930,N_23067);
or UO_45 (O_45,N_21551,N_19032);
nor UO_46 (O_46,N_24120,N_19801);
or UO_47 (O_47,N_23064,N_20993);
nor UO_48 (O_48,N_22538,N_19983);
nand UO_49 (O_49,N_24803,N_21822);
and UO_50 (O_50,N_24140,N_19667);
or UO_51 (O_51,N_20969,N_24846);
xnor UO_52 (O_52,N_23169,N_23512);
and UO_53 (O_53,N_19173,N_22225);
nor UO_54 (O_54,N_19042,N_20415);
xnor UO_55 (O_55,N_20473,N_21544);
xnor UO_56 (O_56,N_21933,N_19330);
xnor UO_57 (O_57,N_19843,N_23892);
nand UO_58 (O_58,N_22372,N_21240);
nor UO_59 (O_59,N_20654,N_23806);
and UO_60 (O_60,N_24965,N_23517);
xnor UO_61 (O_61,N_23847,N_22824);
nor UO_62 (O_62,N_21466,N_21066);
and UO_63 (O_63,N_23675,N_21795);
and UO_64 (O_64,N_20526,N_23246);
xor UO_65 (O_65,N_20818,N_18899);
nor UO_66 (O_66,N_20760,N_24032);
nor UO_67 (O_67,N_23704,N_23238);
nand UO_68 (O_68,N_20377,N_20678);
xor UO_69 (O_69,N_20136,N_20046);
nor UO_70 (O_70,N_22195,N_22286);
and UO_71 (O_71,N_24732,N_22850);
or UO_72 (O_72,N_19343,N_21790);
nor UO_73 (O_73,N_22496,N_20164);
nand UO_74 (O_74,N_18890,N_22476);
xor UO_75 (O_75,N_21412,N_24350);
xor UO_76 (O_76,N_24736,N_20998);
nor UO_77 (O_77,N_19248,N_23501);
and UO_78 (O_78,N_22147,N_21782);
or UO_79 (O_79,N_24531,N_20937);
nand UO_80 (O_80,N_23645,N_22122);
nand UO_81 (O_81,N_20347,N_23908);
and UO_82 (O_82,N_21402,N_20936);
xor UO_83 (O_83,N_24804,N_19337);
xnor UO_84 (O_84,N_24013,N_22838);
or UO_85 (O_85,N_24312,N_21834);
and UO_86 (O_86,N_20383,N_19257);
nor UO_87 (O_87,N_19578,N_19398);
or UO_88 (O_88,N_19334,N_21292);
or UO_89 (O_89,N_24997,N_23778);
nand UO_90 (O_90,N_20074,N_19666);
and UO_91 (O_91,N_20262,N_22897);
xor UO_92 (O_92,N_20168,N_19966);
nor UO_93 (O_93,N_24008,N_22517);
nand UO_94 (O_94,N_23914,N_20180);
or UO_95 (O_95,N_24408,N_22646);
or UO_96 (O_96,N_22422,N_22590);
and UO_97 (O_97,N_22085,N_20325);
nor UO_98 (O_98,N_24392,N_21246);
or UO_99 (O_99,N_20768,N_20844);
nand UO_100 (O_100,N_22057,N_23696);
nor UO_101 (O_101,N_21669,N_22919);
nand UO_102 (O_102,N_19041,N_19723);
nand UO_103 (O_103,N_21003,N_23058);
or UO_104 (O_104,N_21692,N_24538);
nor UO_105 (O_105,N_23159,N_23166);
xnor UO_106 (O_106,N_23252,N_21132);
xnor UO_107 (O_107,N_22698,N_24933);
xor UO_108 (O_108,N_20769,N_23776);
nand UO_109 (O_109,N_24816,N_19044);
or UO_110 (O_110,N_24875,N_24703);
xnor UO_111 (O_111,N_20631,N_19179);
xor UO_112 (O_112,N_19389,N_21938);
nand UO_113 (O_113,N_19288,N_19193);
or UO_114 (O_114,N_19868,N_19366);
or UO_115 (O_115,N_22633,N_20045);
xnor UO_116 (O_116,N_24671,N_23145);
xor UO_117 (O_117,N_23328,N_20832);
or UO_118 (O_118,N_22772,N_21428);
nand UO_119 (O_119,N_20627,N_23727);
nor UO_120 (O_120,N_23198,N_23943);
xnor UO_121 (O_121,N_22140,N_21722);
nor UO_122 (O_122,N_24344,N_24387);
nor UO_123 (O_123,N_23812,N_22311);
or UO_124 (O_124,N_20200,N_24313);
xor UO_125 (O_125,N_22531,N_20542);
xnor UO_126 (O_126,N_19855,N_19228);
and UO_127 (O_127,N_19925,N_20563);
xor UO_128 (O_128,N_22624,N_24748);
nor UO_129 (O_129,N_24234,N_22664);
and UO_130 (O_130,N_23391,N_19072);
nand UO_131 (O_131,N_20591,N_24869);
nor UO_132 (O_132,N_20567,N_20110);
nand UO_133 (O_133,N_20313,N_23054);
and UO_134 (O_134,N_23010,N_23043);
or UO_135 (O_135,N_21924,N_22363);
nand UO_136 (O_136,N_21497,N_24162);
nand UO_137 (O_137,N_22851,N_22800);
nand UO_138 (O_138,N_20362,N_19611);
xor UO_139 (O_139,N_22036,N_23516);
or UO_140 (O_140,N_24841,N_24903);
nor UO_141 (O_141,N_18879,N_20210);
nand UO_142 (O_142,N_20063,N_18829);
nor UO_143 (O_143,N_20559,N_19778);
nand UO_144 (O_144,N_18975,N_24220);
nor UO_145 (O_145,N_21545,N_24278);
and UO_146 (O_146,N_23709,N_18820);
xor UO_147 (O_147,N_24775,N_24051);
or UO_148 (O_148,N_19112,N_24365);
xor UO_149 (O_149,N_22070,N_23523);
nand UO_150 (O_150,N_23381,N_24171);
and UO_151 (O_151,N_20039,N_22779);
and UO_152 (O_152,N_21523,N_23459);
nand UO_153 (O_153,N_24304,N_21032);
nand UO_154 (O_154,N_22325,N_19121);
nor UO_155 (O_155,N_19479,N_23753);
nor UO_156 (O_156,N_24818,N_23940);
nor UO_157 (O_157,N_23640,N_19740);
and UO_158 (O_158,N_23421,N_18994);
nand UO_159 (O_159,N_22098,N_21119);
or UO_160 (O_160,N_21829,N_20469);
and UO_161 (O_161,N_19853,N_22704);
or UO_162 (O_162,N_23606,N_22510);
nand UO_163 (O_163,N_24132,N_22366);
xor UO_164 (O_164,N_24850,N_20203);
nor UO_165 (O_165,N_19134,N_23890);
xnor UO_166 (O_166,N_21632,N_23912);
and UO_167 (O_167,N_19970,N_24363);
nor UO_168 (O_168,N_22882,N_20273);
xor UO_169 (O_169,N_24173,N_22960);
and UO_170 (O_170,N_20482,N_23443);
or UO_171 (O_171,N_24050,N_20698);
and UO_172 (O_172,N_19640,N_23862);
nor UO_173 (O_173,N_24619,N_21210);
and UO_174 (O_174,N_19305,N_24535);
xor UO_175 (O_175,N_24719,N_20390);
xor UO_176 (O_176,N_19293,N_23397);
or UO_177 (O_177,N_23815,N_19512);
nor UO_178 (O_178,N_20558,N_23572);
nor UO_179 (O_179,N_19268,N_19936);
and UO_180 (O_180,N_20763,N_22828);
and UO_181 (O_181,N_21671,N_23872);
nor UO_182 (O_182,N_23673,N_22438);
and UO_183 (O_183,N_23615,N_23655);
and UO_184 (O_184,N_21973,N_19461);
or UO_185 (O_185,N_19695,N_23228);
and UO_186 (O_186,N_22099,N_19652);
nor UO_187 (O_187,N_22217,N_20731);
or UO_188 (O_188,N_21726,N_20225);
xnor UO_189 (O_189,N_19907,N_24972);
and UO_190 (O_190,N_23851,N_21890);
nor UO_191 (O_191,N_19976,N_18812);
and UO_192 (O_192,N_23467,N_21037);
and UO_193 (O_193,N_22843,N_22364);
nor UO_194 (O_194,N_23670,N_23643);
or UO_195 (O_195,N_23573,N_20928);
xor UO_196 (O_196,N_19470,N_21242);
xnor UO_197 (O_197,N_21962,N_24272);
xnor UO_198 (O_198,N_22522,N_18895);
xnor UO_199 (O_199,N_23850,N_22226);
nor UO_200 (O_200,N_21755,N_21873);
nor UO_201 (O_201,N_22058,N_20995);
nor UO_202 (O_202,N_24910,N_20219);
or UO_203 (O_203,N_22738,N_24341);
nor UO_204 (O_204,N_20786,N_20712);
nor UO_205 (O_205,N_18789,N_18932);
and UO_206 (O_206,N_22253,N_23402);
nor UO_207 (O_207,N_24783,N_19076);
nand UO_208 (O_208,N_23023,N_24587);
nor UO_209 (O_209,N_21876,N_20116);
nor UO_210 (O_210,N_19498,N_23868);
or UO_211 (O_211,N_21126,N_19353);
or UO_212 (O_212,N_24604,N_22551);
nand UO_213 (O_213,N_18769,N_24152);
and UO_214 (O_214,N_22464,N_23500);
nor UO_215 (O_215,N_21764,N_23519);
nand UO_216 (O_216,N_20195,N_18861);
xnor UO_217 (O_217,N_22013,N_19050);
xnor UO_218 (O_218,N_19562,N_23481);
and UO_219 (O_219,N_18800,N_24561);
and UO_220 (O_220,N_24212,N_21459);
or UO_221 (O_221,N_24343,N_21255);
and UO_222 (O_222,N_20681,N_19854);
nor UO_223 (O_223,N_18971,N_21352);
or UO_224 (O_224,N_22236,N_24206);
nand UO_225 (O_225,N_23775,N_18772);
and UO_226 (O_226,N_18892,N_24581);
or UO_227 (O_227,N_23158,N_23649);
nand UO_228 (O_228,N_21323,N_19735);
xnor UO_229 (O_229,N_24059,N_19517);
xnor UO_230 (O_230,N_20571,N_19097);
xor UO_231 (O_231,N_19249,N_21057);
nor UO_232 (O_232,N_24863,N_19616);
xnor UO_233 (O_233,N_24342,N_23207);
or UO_234 (O_234,N_23916,N_19945);
nor UO_235 (O_235,N_22813,N_23038);
nor UO_236 (O_236,N_24263,N_20719);
and UO_237 (O_237,N_22459,N_23855);
nor UO_238 (O_238,N_20239,N_20165);
nor UO_239 (O_239,N_18765,N_19670);
or UO_240 (O_240,N_24222,N_22404);
and UO_241 (O_241,N_24683,N_21096);
and UO_242 (O_242,N_24917,N_22494);
or UO_243 (O_243,N_18825,N_19733);
nor UO_244 (O_244,N_19894,N_21704);
and UO_245 (O_245,N_20534,N_21546);
or UO_246 (O_246,N_24280,N_20006);
nor UO_247 (O_247,N_21317,N_24968);
nor UO_248 (O_248,N_22421,N_20687);
nand UO_249 (O_249,N_24261,N_24753);
nor UO_250 (O_250,N_23910,N_23094);
xor UO_251 (O_251,N_21085,N_24115);
and UO_252 (O_252,N_21023,N_23642);
or UO_253 (O_253,N_19837,N_22426);
nor UO_254 (O_254,N_22737,N_21053);
or UO_255 (O_255,N_21682,N_20851);
xor UO_256 (O_256,N_20677,N_23757);
or UO_257 (O_257,N_24293,N_19335);
nor UO_258 (O_258,N_22905,N_23630);
nor UO_259 (O_259,N_18842,N_20169);
and UO_260 (O_260,N_22280,N_22602);
xnor UO_261 (O_261,N_20833,N_22932);
or UO_262 (O_262,N_20946,N_22651);
nor UO_263 (O_263,N_22405,N_21937);
xnor UO_264 (O_264,N_24180,N_21004);
nand UO_265 (O_265,N_20892,N_24471);
xnor UO_266 (O_266,N_23596,N_24837);
nand UO_267 (O_267,N_22869,N_21407);
nor UO_268 (O_268,N_19281,N_18960);
nor UO_269 (O_269,N_21056,N_24891);
xnor UO_270 (O_270,N_24256,N_24749);
nor UO_271 (O_271,N_19057,N_20471);
nand UO_272 (O_272,N_19947,N_24467);
and UO_273 (O_273,N_21074,N_19447);
or UO_274 (O_274,N_21295,N_24176);
nor UO_275 (O_275,N_23959,N_23587);
xor UO_276 (O_276,N_20396,N_20800);
nor UO_277 (O_277,N_19926,N_21678);
nor UO_278 (O_278,N_24824,N_21108);
nand UO_279 (O_279,N_22533,N_21353);
nand UO_280 (O_280,N_21215,N_22973);
and UO_281 (O_281,N_24969,N_23110);
nand UO_282 (O_282,N_19534,N_23999);
or UO_283 (O_283,N_24412,N_22184);
xor UO_284 (O_284,N_24836,N_21364);
or UO_285 (O_285,N_24641,N_21251);
xnor UO_286 (O_286,N_23889,N_22867);
nor UO_287 (O_287,N_22992,N_23030);
nand UO_288 (O_288,N_20323,N_21917);
or UO_289 (O_289,N_24434,N_24254);
nand UO_290 (O_290,N_22860,N_20408);
nand UO_291 (O_291,N_20158,N_22335);
xnor UO_292 (O_292,N_19574,N_19919);
and UO_293 (O_293,N_22655,N_24662);
and UO_294 (O_294,N_22834,N_24497);
and UO_295 (O_295,N_23963,N_22667);
nand UO_296 (O_296,N_21592,N_20400);
or UO_297 (O_297,N_22658,N_23794);
nand UO_298 (O_298,N_21585,N_23611);
and UO_299 (O_299,N_23939,N_21271);
or UO_300 (O_300,N_21149,N_19836);
or UO_301 (O_301,N_22793,N_19705);
xnor UO_302 (O_302,N_20032,N_19588);
xor UO_303 (O_303,N_20431,N_21511);
nand UO_304 (O_304,N_22244,N_23700);
xor UO_305 (O_305,N_24959,N_22520);
nor UO_306 (O_306,N_20353,N_21156);
xnor UO_307 (O_307,N_24664,N_19978);
and UO_308 (O_308,N_24296,N_21014);
or UO_309 (O_309,N_23821,N_22903);
xnor UO_310 (O_310,N_20111,N_23991);
nor UO_311 (O_311,N_22564,N_22954);
and UO_312 (O_312,N_23144,N_24609);
xor UO_313 (O_313,N_20062,N_19886);
nand UO_314 (O_314,N_23653,N_19979);
xor UO_315 (O_315,N_22949,N_20367);
nand UO_316 (O_316,N_23679,N_22018);
or UO_317 (O_317,N_19184,N_20711);
and UO_318 (O_318,N_19438,N_20749);
or UO_319 (O_319,N_24924,N_23786);
and UO_320 (O_320,N_20226,N_23051);
xnor UO_321 (O_321,N_21673,N_21280);
nand UO_322 (O_322,N_20220,N_22312);
and UO_323 (O_323,N_23751,N_19665);
and UO_324 (O_324,N_19055,N_20505);
nand UO_325 (O_325,N_19903,N_23347);
nand UO_326 (O_326,N_22773,N_19982);
nor UO_327 (O_327,N_18889,N_20010);
nand UO_328 (O_328,N_21664,N_23430);
and UO_329 (O_329,N_22321,N_24200);
and UO_330 (O_330,N_24257,N_19972);
nand UO_331 (O_331,N_24201,N_19296);
and UO_332 (O_332,N_20275,N_19715);
xnor UO_333 (O_333,N_24747,N_23027);
or UO_334 (O_334,N_24058,N_21598);
nand UO_335 (O_335,N_20382,N_21676);
xnor UO_336 (O_336,N_19719,N_22755);
nand UO_337 (O_337,N_19848,N_18974);
xnor UO_338 (O_338,N_19027,N_21047);
and UO_339 (O_339,N_23551,N_23084);
and UO_340 (O_340,N_21533,N_19796);
nor UO_341 (O_341,N_19320,N_22911);
xnor UO_342 (O_342,N_19682,N_22615);
and UO_343 (O_343,N_22211,N_18947);
and UO_344 (O_344,N_24729,N_23689);
nand UO_345 (O_345,N_23131,N_22560);
nor UO_346 (O_346,N_21753,N_24511);
nor UO_347 (O_347,N_21324,N_21244);
xnor UO_348 (O_348,N_22833,N_19948);
xor UO_349 (O_349,N_21435,N_18816);
and UO_350 (O_350,N_20495,N_21575);
and UO_351 (O_351,N_20371,N_23104);
or UO_352 (O_352,N_24774,N_24279);
xnor UO_353 (O_353,N_23146,N_22428);
nand UO_354 (O_354,N_24596,N_19358);
nor UO_355 (O_355,N_19630,N_18792);
nand UO_356 (O_356,N_23783,N_22389);
xor UO_357 (O_357,N_21670,N_24992);
nor UO_358 (O_358,N_20043,N_20737);
nand UO_359 (O_359,N_24243,N_20142);
xnor UO_360 (O_360,N_22050,N_23526);
xnor UO_361 (O_361,N_20720,N_23631);
xnor UO_362 (O_362,N_22410,N_22921);
xor UO_363 (O_363,N_24166,N_24372);
or UO_364 (O_364,N_22866,N_24324);
and UO_365 (O_365,N_21254,N_24126);
or UO_366 (O_366,N_24784,N_23913);
xor UO_367 (O_367,N_20821,N_23278);
nand UO_368 (O_368,N_24915,N_18751);
nor UO_369 (O_369,N_22720,N_23856);
and UO_370 (O_370,N_22008,N_22740);
nand UO_371 (O_371,N_22640,N_24527);
nor UO_372 (O_372,N_18802,N_22855);
nor UO_373 (O_373,N_19457,N_21432);
xnor UO_374 (O_374,N_23841,N_20320);
and UO_375 (O_375,N_22500,N_20523);
xor UO_376 (O_376,N_20055,N_23180);
or UO_377 (O_377,N_18884,N_18837);
or UO_378 (O_378,N_24667,N_19986);
xnor UO_379 (O_379,N_23147,N_24438);
xnor UO_380 (O_380,N_24160,N_21525);
nand UO_381 (O_381,N_19045,N_19506);
or UO_382 (O_382,N_24575,N_21162);
or UO_383 (O_383,N_23824,N_24404);
nor UO_384 (O_384,N_22181,N_23834);
and UO_385 (O_385,N_24988,N_21894);
nand UO_386 (O_386,N_20765,N_24090);
xnor UO_387 (O_387,N_24983,N_21573);
xnor UO_388 (O_388,N_20243,N_24643);
nand UO_389 (O_389,N_20375,N_24827);
nand UO_390 (O_390,N_19949,N_19724);
xor UO_391 (O_391,N_23002,N_23548);
and UO_392 (O_392,N_19386,N_21654);
nor UO_393 (O_393,N_22718,N_21448);
and UO_394 (O_394,N_22831,N_21887);
xor UO_395 (O_395,N_19964,N_19149);
or UO_396 (O_396,N_20589,N_21817);
and UO_397 (O_397,N_21780,N_22189);
and UO_398 (O_398,N_22474,N_20676);
or UO_399 (O_399,N_21257,N_24702);
nand UO_400 (O_400,N_19487,N_21434);
and UO_401 (O_401,N_19164,N_22254);
nand UO_402 (O_402,N_20673,N_20775);
nand UO_403 (O_403,N_21796,N_23579);
or UO_404 (O_404,N_20398,N_23965);
nor UO_405 (O_405,N_23306,N_21880);
nor UO_406 (O_406,N_22635,N_19669);
and UO_407 (O_407,N_23819,N_24923);
nand UO_408 (O_408,N_20084,N_21856);
nor UO_409 (O_409,N_20541,N_22574);
or UO_410 (O_410,N_20460,N_22981);
nand UO_411 (O_411,N_20124,N_22536);
nand UO_412 (O_412,N_20171,N_23752);
nor UO_413 (O_413,N_24435,N_19087);
xnor UO_414 (O_414,N_21715,N_20592);
or UO_415 (O_415,N_19107,N_20759);
nor UO_416 (O_416,N_20788,N_22977);
or UO_417 (O_417,N_23632,N_23769);
xor UO_418 (O_418,N_23463,N_23309);
or UO_419 (O_419,N_23787,N_22413);
and UO_420 (O_420,N_24642,N_22934);
or UO_421 (O_421,N_21942,N_20036);
nand UO_422 (O_422,N_20613,N_18927);
or UO_423 (O_423,N_21232,N_23119);
and UO_424 (O_424,N_22270,N_21071);
nand UO_425 (O_425,N_20642,N_22310);
or UO_426 (O_426,N_23881,N_22495);
nand UO_427 (O_427,N_20267,N_21198);
nor UO_428 (O_428,N_19527,N_21449);
nand UO_429 (O_429,N_20117,N_22466);
xnor UO_430 (O_430,N_24249,N_20662);
nand UO_431 (O_431,N_22395,N_20729);
and UO_432 (O_432,N_20475,N_18860);
nor UO_433 (O_433,N_23203,N_24622);
or UO_434 (O_434,N_19959,N_19060);
xor UO_435 (O_435,N_22082,N_22539);
xnor UO_436 (O_436,N_21761,N_22238);
xor UO_437 (O_437,N_20878,N_21841);
nand UO_438 (O_438,N_23070,N_23546);
nand UO_439 (O_439,N_22110,N_22762);
and UO_440 (O_440,N_20830,N_21142);
xor UO_441 (O_441,N_23575,N_19946);
or UO_442 (O_442,N_22991,N_20372);
xor UO_443 (O_443,N_21898,N_22681);
nor UO_444 (O_444,N_18989,N_22654);
xnor UO_445 (O_445,N_19962,N_21044);
and UO_446 (O_446,N_20008,N_18793);
nor UO_447 (O_447,N_19744,N_20284);
nor UO_448 (O_448,N_19409,N_24146);
nor UO_449 (O_449,N_22307,N_21850);
xor UO_450 (O_450,N_22447,N_19700);
or UO_451 (O_451,N_21583,N_22830);
nand UO_452 (O_452,N_23542,N_24405);
nor UO_453 (O_453,N_24213,N_19143);
and UO_454 (O_454,N_22825,N_23961);
xnor UO_455 (O_455,N_19074,N_24246);
nand UO_456 (O_456,N_24698,N_23374);
nand UO_457 (O_457,N_19441,N_24556);
nor UO_458 (O_458,N_20957,N_19381);
and UO_459 (O_459,N_23904,N_22582);
and UO_460 (O_460,N_23461,N_21883);
nand UO_461 (O_461,N_21996,N_24031);
or UO_462 (O_462,N_24123,N_19233);
xor UO_463 (O_463,N_19614,N_20333);
or UO_464 (O_464,N_24084,N_22205);
nor UO_465 (O_465,N_19590,N_20498);
or UO_466 (O_466,N_19392,N_22741);
and UO_467 (O_467,N_19231,N_24223);
nand UO_468 (O_468,N_23441,N_24862);
or UO_469 (O_469,N_22812,N_22396);
nand UO_470 (O_470,N_22805,N_19646);
or UO_471 (O_471,N_21418,N_22048);
and UO_472 (O_472,N_19975,N_18925);
or UO_473 (O_473,N_19295,N_22846);
nor UO_474 (O_474,N_23258,N_20030);
and UO_475 (O_475,N_20297,N_19712);
nor UO_476 (O_476,N_22318,N_21907);
xor UO_477 (O_477,N_22734,N_20773);
nand UO_478 (O_478,N_18963,N_21823);
xnor UO_479 (O_479,N_20746,N_23156);
and UO_480 (O_480,N_22432,N_23452);
and UO_481 (O_481,N_22007,N_23488);
nor UO_482 (O_482,N_19454,N_20813);
nand UO_483 (O_483,N_19219,N_23938);
nand UO_484 (O_484,N_24015,N_20869);
or UO_485 (O_485,N_24794,N_20190);
nand UO_486 (O_486,N_21980,N_21522);
xnor UO_487 (O_487,N_19301,N_22465);
and UO_488 (O_488,N_21339,N_20064);
nand UO_489 (O_489,N_24925,N_20544);
nand UO_490 (O_490,N_20628,N_19473);
and UO_491 (O_491,N_23663,N_24275);
nor UO_492 (O_492,N_19440,N_19887);
or UO_493 (O_493,N_21769,N_19376);
nand UO_494 (O_494,N_19602,N_20489);
nor UO_495 (O_495,N_24501,N_19309);
nor UO_496 (O_496,N_19345,N_23174);
nand UO_497 (O_497,N_24118,N_21010);
nor UO_498 (O_498,N_21661,N_21724);
nand UO_499 (O_499,N_24672,N_20421);
nor UO_500 (O_500,N_21981,N_20067);
xnor UO_501 (O_501,N_19130,N_21848);
nor UO_502 (O_502,N_23229,N_23765);
or UO_503 (O_503,N_24188,N_22198);
or UO_504 (O_504,N_24239,N_23747);
nor UO_505 (O_505,N_19000,N_23243);
nand UO_506 (O_506,N_22671,N_19102);
and UO_507 (O_507,N_19623,N_23957);
xor UO_508 (O_508,N_22179,N_22235);
or UO_509 (O_509,N_18788,N_19279);
and UO_510 (O_510,N_21387,N_19773);
and UO_511 (O_511,N_24982,N_24876);
and UO_512 (O_512,N_21147,N_21901);
xnor UO_513 (O_513,N_24790,N_24006);
nand UO_514 (O_514,N_18770,N_19525);
nor UO_515 (O_515,N_18813,N_22431);
xor UO_516 (O_516,N_20660,N_23405);
nor UO_517 (O_517,N_23401,N_24878);
or UO_518 (O_518,N_23075,N_24495);
and UO_519 (O_519,N_20801,N_21845);
nor UO_520 (O_520,N_19998,N_18779);
and UO_521 (O_521,N_19240,N_19111);
nor UO_522 (O_522,N_20128,N_19493);
nor UO_523 (O_523,N_19198,N_21182);
nand UO_524 (O_524,N_22512,N_20975);
and UO_525 (O_525,N_22794,N_23213);
nor UO_526 (O_526,N_22360,N_22910);
nand UO_527 (O_527,N_22776,N_21570);
xnor UO_528 (O_528,N_20549,N_19742);
and UO_529 (O_529,N_24195,N_22937);
or UO_530 (O_530,N_20641,N_19782);
and UO_531 (O_531,N_21816,N_23383);
xnor UO_532 (O_532,N_22154,N_22202);
nor UO_533 (O_533,N_19663,N_19952);
nor UO_534 (O_534,N_24483,N_18806);
nor UO_535 (O_535,N_24484,N_24442);
and UO_536 (O_536,N_20896,N_23662);
and UO_537 (O_537,N_22054,N_24011);
nor UO_538 (O_538,N_22508,N_23385);
nor UO_539 (O_539,N_24230,N_19621);
and UO_540 (O_540,N_21388,N_24418);
nor UO_541 (O_541,N_19507,N_23333);
nor UO_542 (O_542,N_23226,N_21018);
or UO_543 (O_543,N_23483,N_20253);
or UO_544 (O_544,N_22606,N_23279);
nand UO_545 (O_545,N_24632,N_21098);
xor UO_546 (O_546,N_18952,N_23239);
or UO_547 (O_547,N_20299,N_22103);
nand UO_548 (O_548,N_23493,N_21143);
xor UO_549 (O_549,N_21019,N_20365);
nand UO_550 (O_550,N_23756,N_23011);
xnor UO_551 (O_551,N_19607,N_24251);
xnor UO_552 (O_552,N_23220,N_23249);
or UO_553 (O_553,N_19720,N_22966);
and UO_554 (O_554,N_24266,N_24900);
nand UO_555 (O_555,N_23091,N_22791);
nor UO_556 (O_556,N_20976,N_24161);
nor UO_557 (O_557,N_19989,N_19357);
and UO_558 (O_558,N_20105,N_24454);
xor UO_559 (O_559,N_24231,N_24253);
nor UO_560 (O_560,N_22319,N_23932);
nand UO_561 (O_561,N_20805,N_20380);
and UO_562 (O_562,N_21781,N_21604);
xnor UO_563 (O_563,N_21732,N_22151);
nand UO_564 (O_564,N_24335,N_23789);
and UO_565 (O_565,N_23683,N_22457);
or UO_566 (O_566,N_20071,N_23138);
xnor UO_567 (O_567,N_22798,N_22746);
or UO_568 (O_568,N_20600,N_20296);
nand UO_569 (O_569,N_24157,N_18855);
and UO_570 (O_570,N_24976,N_22358);
or UO_571 (O_571,N_22854,N_21927);
and UO_572 (O_572,N_24192,N_19410);
and UO_573 (O_573,N_21204,N_24071);
xor UO_574 (O_574,N_24494,N_20757);
and UO_575 (O_575,N_18946,N_23434);
nand UO_576 (O_576,N_24806,N_21716);
xnor UO_577 (O_577,N_22818,N_22971);
or UO_578 (O_578,N_21964,N_24446);
nand UO_579 (O_579,N_20364,N_19960);
nand UO_580 (O_580,N_24894,N_19749);
nand UO_581 (O_581,N_20556,N_19603);
nor UO_582 (O_582,N_21252,N_19898);
xor UO_583 (O_583,N_24492,N_18999);
xnor UO_584 (O_584,N_22126,N_18835);
and UO_585 (O_585,N_22545,N_20014);
and UO_586 (O_586,N_22708,N_23942);
xor UO_587 (O_587,N_24842,N_21011);
or UO_588 (O_588,N_24410,N_19559);
xor UO_589 (O_589,N_21843,N_24966);
and UO_590 (O_590,N_20004,N_21442);
xor UO_591 (O_591,N_20433,N_22694);
xnor UO_592 (O_592,N_18876,N_21900);
xnor UO_593 (O_593,N_21736,N_18784);
and UO_594 (O_594,N_23685,N_21329);
nand UO_595 (O_595,N_21611,N_24208);
nor UO_596 (O_596,N_19036,N_19077);
nand UO_597 (O_597,N_20459,N_20503);
xor UO_598 (O_598,N_19849,N_24145);
and UO_599 (O_599,N_22033,N_19197);
nor UO_600 (O_600,N_22162,N_22972);
nand UO_601 (O_601,N_18921,N_19140);
and UO_602 (O_602,N_22853,N_20161);
nor UO_603 (O_603,N_24457,N_21405);
nand UO_604 (O_604,N_24136,N_20250);
nand UO_605 (O_605,N_24439,N_21872);
xnor UO_606 (O_606,N_24477,N_23041);
xor UO_607 (O_607,N_23474,N_19784);
xor UO_608 (O_608,N_23634,N_22367);
and UO_609 (O_609,N_23539,N_21117);
or UO_610 (O_610,N_19344,N_19349);
nor UO_611 (O_611,N_20130,N_20651);
xnor UO_612 (O_612,N_20934,N_22032);
or UO_613 (O_613,N_22343,N_21855);
nor UO_614 (O_614,N_21743,N_20311);
or UO_615 (O_615,N_20564,N_21391);
nor UO_616 (O_616,N_18956,N_24658);
nand UO_617 (O_617,N_24695,N_22993);
nor UO_618 (O_618,N_20401,N_21740);
or UO_619 (O_619,N_20581,N_19557);
and UO_620 (O_620,N_23337,N_20279);
nor UO_621 (O_621,N_22893,N_21717);
xnor UO_622 (O_622,N_23322,N_19867);
or UO_623 (O_623,N_22584,N_19278);
and UO_624 (O_624,N_20939,N_24367);
nor UO_625 (O_625,N_23831,N_21600);
and UO_626 (O_626,N_19653,N_20785);
nor UO_627 (O_627,N_22145,N_21231);
nor UO_628 (O_628,N_23188,N_24360);
and UO_629 (O_629,N_21506,N_23281);
or UO_630 (O_630,N_19236,N_22717);
and UO_631 (O_631,N_20445,N_18823);
and UO_632 (O_632,N_18900,N_24559);
or UO_633 (O_633,N_23607,N_23254);
nor UO_634 (O_634,N_22810,N_24590);
or UO_635 (O_635,N_24020,N_19132);
and UO_636 (O_636,N_21282,N_24310);
or UO_637 (O_637,N_20842,N_22929);
or UO_638 (O_638,N_19808,N_24395);
nand UO_639 (O_639,N_19078,N_24207);
or UO_640 (O_640,N_24684,N_22706);
or UO_641 (O_641,N_22030,N_24326);
nor UO_642 (O_642,N_23729,N_20500);
or UO_643 (O_643,N_22449,N_22331);
and UO_644 (O_644,N_20949,N_20249);
nor UO_645 (O_645,N_21325,N_24444);
and UO_646 (O_646,N_23953,N_19374);
nor UO_647 (O_647,N_21808,N_20327);
xnor UO_648 (O_648,N_22849,N_23045);
nand UO_649 (O_649,N_21778,N_18973);
xor UO_650 (O_650,N_19429,N_19156);
and UO_651 (O_651,N_22439,N_24696);
and UO_652 (O_652,N_24832,N_20834);
nor UO_653 (O_653,N_21516,N_24056);
nor UO_654 (O_654,N_21104,N_20202);
nor UO_655 (O_655,N_24958,N_21043);
and UO_656 (O_656,N_18926,N_22901);
xor UO_657 (O_657,N_21453,N_22233);
or UO_658 (O_658,N_21952,N_21589);
or UO_659 (O_659,N_24985,N_21430);
or UO_660 (O_660,N_20280,N_23005);
xnor UO_661 (O_661,N_22802,N_20861);
xnor UO_662 (O_662,N_20294,N_24537);
nand UO_663 (O_663,N_22997,N_21478);
xnor UO_664 (O_664,N_22316,N_24994);
nor UO_665 (O_665,N_21217,N_23906);
or UO_666 (O_666,N_19110,N_23650);
xor UO_667 (O_667,N_20217,N_20695);
and UO_668 (O_668,N_19194,N_24423);
nand UO_669 (O_669,N_24053,N_22819);
or UO_670 (O_670,N_23694,N_20714);
nand UO_671 (O_671,N_23102,N_22697);
nand UO_672 (O_672,N_23208,N_24077);
xor UO_673 (O_673,N_21343,N_21383);
and UO_674 (O_674,N_20565,N_21291);
nand UO_675 (O_675,N_19499,N_23978);
or UO_676 (O_676,N_19969,N_23718);
nand UO_677 (O_677,N_23455,N_23440);
xnor UO_678 (O_678,N_19505,N_23767);
or UO_679 (O_679,N_19830,N_19647);
nand UO_680 (O_680,N_21509,N_23209);
nand UO_681 (O_681,N_23003,N_20574);
or UO_682 (O_682,N_24174,N_21027);
or UO_683 (O_683,N_23376,N_24989);
xnor UO_684 (O_684,N_24757,N_21771);
nand UO_685 (O_685,N_21318,N_19119);
or UO_686 (O_686,N_21065,N_19478);
nor UO_687 (O_687,N_23412,N_23193);
and UO_688 (O_688,N_21045,N_24845);
xor UO_689 (O_689,N_22446,N_24428);
xor UO_690 (O_690,N_20670,N_24714);
and UO_691 (O_691,N_20187,N_21176);
or UO_692 (O_692,N_19661,N_19468);
nor UO_693 (O_693,N_22159,N_22513);
or UO_694 (O_694,N_18942,N_23267);
xnor UO_695 (O_695,N_20443,N_23227);
xor UO_696 (O_696,N_21200,N_20048);
nand UO_697 (O_697,N_21734,N_20255);
xor UO_698 (O_698,N_24024,N_24124);
and UO_699 (O_699,N_19348,N_20446);
nand UO_700 (O_700,N_21700,N_19234);
nand UO_701 (O_701,N_21479,N_24975);
nand UO_702 (O_702,N_22962,N_24111);
xnor UO_703 (O_703,N_21809,N_23487);
or UO_704 (O_704,N_19626,N_21285);
xnor UO_705 (O_705,N_22770,N_22095);
or UO_706 (O_706,N_23941,N_22857);
or UO_707 (O_707,N_24317,N_23480);
nor UO_708 (O_708,N_23922,N_22306);
or UO_709 (O_709,N_20103,N_20629);
nand UO_710 (O_710,N_23251,N_19354);
nor UO_711 (O_711,N_22344,N_19306);
nor UO_712 (O_712,N_21234,N_23048);
xor UO_713 (O_713,N_20437,N_22340);
nand UO_714 (O_714,N_20507,N_18898);
nor UO_715 (O_715,N_23864,N_19269);
and UO_716 (O_716,N_19788,N_22806);
nor UO_717 (O_717,N_18791,N_19011);
or UO_718 (O_718,N_18951,N_20942);
and UO_719 (O_719,N_22670,N_22037);
nor UO_720 (O_720,N_23554,N_22302);
nor UO_721 (O_721,N_24330,N_23154);
or UO_722 (O_722,N_20625,N_21892);
nand UO_723 (O_723,N_22351,N_21015);
and UO_724 (O_724,N_21739,N_22148);
nor UO_725 (O_725,N_21521,N_20221);
nand UO_726 (O_726,N_23608,N_21861);
and UO_727 (O_727,N_20578,N_22260);
and UO_728 (O_728,N_23420,N_24133);
or UO_729 (O_729,N_22090,N_24070);
nand UO_730 (O_730,N_24598,N_21495);
xnor UO_731 (O_731,N_20439,N_23581);
or UO_732 (O_732,N_19326,N_20470);
xnor UO_733 (O_733,N_21895,N_24733);
or UO_734 (O_734,N_22899,N_20979);
nand UO_735 (O_735,N_19275,N_21360);
or UO_736 (O_736,N_21068,N_20025);
nand UO_737 (O_737,N_21814,N_21139);
and UO_738 (O_738,N_23348,N_19679);
and UO_739 (O_739,N_20127,N_18787);
or UO_740 (O_740,N_22946,N_22884);
nand UO_741 (O_741,N_23414,N_21785);
or UO_742 (O_742,N_19839,N_19681);
nand UO_743 (O_743,N_22769,N_20322);
nor UO_744 (O_744,N_22131,N_20806);
and UO_745 (O_745,N_24797,N_21083);
nand UO_746 (O_746,N_19648,N_23446);
and UO_747 (O_747,N_20965,N_21346);
nand UO_748 (O_748,N_19459,N_22647);
and UO_749 (O_749,N_23971,N_24610);
or UO_750 (O_750,N_24485,N_19062);
nor UO_751 (O_751,N_22519,N_24214);
xor UO_752 (O_752,N_24415,N_19012);
nor UO_753 (O_753,N_18911,N_19997);
and UO_754 (O_754,N_19528,N_19239);
or UO_755 (O_755,N_23636,N_23610);
nor UO_756 (O_756,N_18944,N_20533);
xor UO_757 (O_757,N_23211,N_19363);
xnor UO_758 (O_758,N_23829,N_24088);
nand UO_759 (O_759,N_21501,N_21103);
and UO_760 (O_760,N_21035,N_21982);
nand UO_761 (O_761,N_20990,N_19406);
xnor UO_762 (O_762,N_19526,N_24829);
or UO_763 (O_763,N_24651,N_19421);
nand UO_764 (O_764,N_19596,N_19284);
and UO_765 (O_765,N_20996,N_21136);
nand UO_766 (O_766,N_21185,N_21298);
nor UO_767 (O_767,N_21754,N_19685);
nor UO_768 (O_768,N_19023,N_24669);
nor UO_769 (O_769,N_24922,N_19212);
and UO_770 (O_770,N_20513,N_18894);
or UO_771 (O_771,N_22451,N_23085);
nand UO_772 (O_772,N_24617,N_21804);
nand UO_773 (O_773,N_23123,N_19609);
and UO_774 (O_774,N_18901,N_24639);
xor UO_775 (O_775,N_23289,N_24420);
and UO_776 (O_776,N_19202,N_20597);
or UO_777 (O_777,N_24526,N_19283);
or UO_778 (O_778,N_21050,N_24640);
nor UO_779 (O_779,N_23997,N_24346);
nor UO_780 (O_780,N_20260,N_20741);
or UO_781 (O_781,N_22693,N_19683);
nand UO_782 (O_782,N_23559,N_22322);
and UO_783 (O_783,N_24844,N_19692);
or UO_784 (O_784,N_21899,N_19531);
xor UO_785 (O_785,N_19865,N_22876);
or UO_786 (O_786,N_24034,N_19569);
or UO_787 (O_787,N_24548,N_20209);
nor UO_788 (O_788,N_24828,N_24158);
or UO_789 (O_789,N_20974,N_22006);
nand UO_790 (O_790,N_20412,N_19834);
nor UO_791 (O_791,N_24194,N_22847);
or UO_792 (O_792,N_23918,N_20791);
nand UO_793 (O_793,N_19001,N_24810);
nand UO_794 (O_794,N_23873,N_19797);
xnor UO_795 (O_795,N_24033,N_22332);
nor UO_796 (O_796,N_19444,N_22504);
nand UO_797 (O_797,N_23234,N_21946);
nand UO_798 (O_798,N_20357,N_22692);
or UO_799 (O_799,N_18807,N_23503);
nand UO_800 (O_800,N_24402,N_21607);
xor UO_801 (O_801,N_19445,N_24674);
and UO_802 (O_802,N_24196,N_19956);
or UO_803 (O_803,N_23472,N_19196);
nand UO_804 (O_804,N_19594,N_22592);
xnor UO_805 (O_805,N_21555,N_24184);
and UO_806 (O_806,N_21487,N_20012);
xnor UO_807 (O_807,N_21485,N_23122);
nand UO_808 (O_808,N_24715,N_24129);
or UO_809 (O_809,N_23885,N_22865);
xor UO_810 (O_810,N_23637,N_24938);
xnor UO_811 (O_811,N_22713,N_24193);
or UO_812 (O_812,N_24001,N_20727);
nor UO_813 (O_813,N_20351,N_23688);
or UO_814 (O_814,N_23671,N_24588);
and UO_815 (O_815,N_22493,N_22499);
xnor UO_816 (O_816,N_22611,N_20211);
nand UO_817 (O_817,N_19336,N_19615);
or UO_818 (O_818,N_24455,N_21454);
xor UO_819 (O_819,N_20033,N_20397);
and UO_820 (O_820,N_21207,N_24361);
nor UO_821 (O_821,N_21560,N_24252);
nand UO_822 (O_822,N_22251,N_19108);
nor UO_823 (O_823,N_22080,N_22197);
xnor UO_824 (O_824,N_24496,N_20406);
and UO_825 (O_825,N_20853,N_19270);
nand UO_826 (O_826,N_24401,N_24096);
nor UO_827 (O_827,N_22158,N_19910);
or UO_828 (O_828,N_24909,N_21052);
nand UO_829 (O_829,N_19360,N_23173);
nor UO_830 (O_830,N_20587,N_21385);
nand UO_831 (O_831,N_19644,N_23724);
nor UO_832 (O_832,N_21189,N_22662);
and UO_833 (O_833,N_24765,N_23731);
xor UO_834 (O_834,N_20404,N_21358);
and UO_835 (O_835,N_24597,N_19934);
or UO_836 (O_836,N_20289,N_24366);
nand UO_837 (O_837,N_20783,N_24699);
and UO_838 (O_838,N_20229,N_20888);
nor UO_839 (O_839,N_19482,N_23714);
nand UO_840 (O_840,N_21909,N_19380);
or UO_841 (O_841,N_20693,N_24607);
nor UO_842 (O_842,N_21630,N_19052);
nor UO_843 (O_843,N_19752,N_22067);
nand UO_844 (O_844,N_22996,N_23846);
and UO_845 (O_845,N_18846,N_22809);
and UO_846 (O_846,N_22392,N_23870);
and UO_847 (O_847,N_22956,N_22059);
nor UO_848 (O_848,N_24830,N_21344);
xor UO_849 (O_849,N_22811,N_23707);
or UO_850 (O_850,N_22565,N_21333);
nand UO_851 (O_851,N_19745,N_22758);
nand UO_852 (O_852,N_19922,N_23504);
nor UO_853 (O_853,N_24741,N_23042);
nand UO_854 (O_854,N_22094,N_22454);
and UO_855 (O_855,N_19765,N_22213);
xor UO_856 (O_856,N_24697,N_20989);
xnor UO_857 (O_857,N_23296,N_24143);
nand UO_858 (O_858,N_21167,N_22473);
or UO_859 (O_859,N_23882,N_19464);
nand UO_860 (O_860,N_23149,N_19856);
and UO_861 (O_861,N_19104,N_24165);
and UO_862 (O_862,N_24042,N_22262);
nand UO_863 (O_863,N_24432,N_19382);
nand UO_864 (O_864,N_23962,N_21810);
and UO_865 (O_865,N_19864,N_23869);
and UO_866 (O_866,N_20241,N_23613);
nand UO_867 (O_867,N_20917,N_24450);
nand UO_868 (O_868,N_22927,N_24509);
and UO_869 (O_869,N_24183,N_21179);
or UO_870 (O_870,N_24308,N_24764);
nand UO_871 (O_871,N_22787,N_21547);
nand UO_872 (O_872,N_23400,N_19368);
nand UO_873 (O_873,N_24627,N_20648);
or UO_874 (O_874,N_21482,N_24521);
xor UO_875 (O_875,N_22621,N_22064);
nand UO_876 (O_876,N_23515,N_24175);
nand UO_877 (O_877,N_19546,N_18762);
nand UO_878 (O_878,N_20118,N_23797);
or UO_879 (O_879,N_20906,N_19139);
xnor UO_880 (O_880,N_24399,N_24000);
nand UO_881 (O_881,N_23735,N_22004);
or UO_882 (O_882,N_19157,N_23116);
nor UO_883 (O_883,N_19980,N_23026);
xor UO_884 (O_884,N_21274,N_19963);
and UO_885 (O_885,N_23451,N_19372);
nand UO_886 (O_886,N_20468,N_22628);
nor UO_887 (O_887,N_21008,N_22448);
or UO_888 (O_888,N_22724,N_24487);
or UO_889 (O_889,N_19658,N_18986);
or UO_890 (O_890,N_21542,N_20667);
nor UO_891 (O_891,N_24406,N_20945);
nand UO_892 (O_892,N_22742,N_21513);
and UO_893 (O_893,N_21256,N_18887);
and UO_894 (O_894,N_23183,N_23134);
and UO_895 (O_895,N_23126,N_19034);
nor UO_896 (O_896,N_19384,N_20784);
nand UO_897 (O_897,N_20933,N_20579);
or UO_898 (O_898,N_19302,N_20252);
and UO_899 (O_899,N_20901,N_18983);
nor UO_900 (O_900,N_23106,N_19504);
nand UO_901 (O_901,N_21864,N_19452);
and UO_902 (O_902,N_18933,N_18930);
xnor UO_903 (O_903,N_19746,N_19828);
nand UO_904 (O_904,N_21087,N_20825);
or UO_905 (O_905,N_21309,N_19747);
xnor UO_906 (O_906,N_19629,N_19207);
nor UO_907 (O_907,N_19882,N_19144);
and UO_908 (O_908,N_19480,N_20223);
and UO_909 (O_909,N_18979,N_24649);
nor UO_910 (O_910,N_20155,N_20758);
xor UO_911 (O_911,N_20958,N_24105);
nand UO_912 (O_912,N_23482,N_24153);
and UO_913 (O_913,N_20743,N_20339);
xnor UO_914 (O_914,N_19757,N_22304);
xor UO_915 (O_915,N_24731,N_20972);
xor UO_916 (O_916,N_24390,N_21130);
nand UO_917 (O_917,N_20512,N_19127);
nand UO_918 (O_918,N_19090,N_24241);
and UO_919 (O_919,N_21552,N_24431);
xnor UO_920 (O_920,N_18830,N_18827);
nor UO_921 (O_921,N_20781,N_18948);
and UO_922 (O_922,N_20601,N_20053);
nor UO_923 (O_923,N_23592,N_19957);
or UO_924 (O_924,N_23521,N_19313);
and UO_925 (O_925,N_24935,N_22686);
xnor UO_926 (O_926,N_19988,N_24142);
xor UO_927 (O_927,N_24233,N_24203);
nand UO_928 (O_928,N_20885,N_24680);
nand UO_929 (O_929,N_19518,N_22230);
and UO_930 (O_930,N_19466,N_24443);
xor UO_931 (O_931,N_23568,N_23413);
nor UO_932 (O_932,N_19608,N_23247);
nor UO_933 (O_933,N_23498,N_23556);
and UO_934 (O_934,N_21991,N_24522);
or UO_935 (O_935,N_22382,N_19537);
and UO_936 (O_936,N_18928,N_24650);
xnor UO_937 (O_937,N_22516,N_19754);
or UO_938 (O_938,N_21830,N_19955);
or UO_939 (O_939,N_20370,N_21751);
xor UO_940 (O_940,N_19133,N_23814);
nand UO_941 (O_941,N_23973,N_19200);
nor UO_942 (O_942,N_21984,N_19243);
and UO_943 (O_943,N_23837,N_24998);
nand UO_944 (O_944,N_21802,N_19287);
or UO_945 (O_945,N_21903,N_22357);
and UO_946 (O_946,N_24685,N_24295);
xnor UO_947 (O_947,N_23711,N_20925);
and UO_948 (O_948,N_19731,N_20706);
and UO_949 (O_949,N_20538,N_20194);
xor UO_950 (O_950,N_24594,N_19532);
nor UO_951 (O_951,N_20182,N_21621);
and UO_952 (O_952,N_18866,N_24210);
and UO_953 (O_953,N_21989,N_20496);
and UO_954 (O_954,N_19577,N_19850);
xor UO_955 (O_955,N_24355,N_18918);
and UO_956 (O_956,N_19794,N_23710);
xor UO_957 (O_957,N_23528,N_22294);
and UO_958 (O_958,N_22377,N_19475);
xnor UO_959 (O_959,N_22379,N_22721);
and UO_960 (O_960,N_24321,N_23601);
xor UO_961 (O_961,N_20423,N_23665);
nor UO_962 (O_962,N_21811,N_23895);
nand UO_963 (O_963,N_20887,N_24323);
or UO_964 (O_964,N_23931,N_21446);
or UO_965 (O_965,N_23612,N_22186);
nand UO_966 (O_966,N_24463,N_21386);
xnor UO_967 (O_967,N_19587,N_23715);
nand UO_968 (O_968,N_19160,N_18880);
and UO_969 (O_969,N_22568,N_21092);
and UO_970 (O_970,N_23407,N_18781);
or UO_971 (O_971,N_24602,N_24269);
or UO_972 (O_972,N_20497,N_22214);
nand UO_973 (O_973,N_20035,N_19066);
or UO_974 (O_974,N_19800,N_21742);
or UO_975 (O_975,N_19232,N_24505);
or UO_976 (O_976,N_19054,N_21972);
or UO_977 (O_977,N_22619,N_24948);
or UO_978 (O_978,N_19789,N_20242);
and UO_979 (O_979,N_21997,N_21000);
xnor UO_980 (O_980,N_20665,N_23734);
nand UO_981 (O_981,N_18870,N_21965);
nor UO_982 (O_982,N_19613,N_24393);
xor UO_983 (O_983,N_21539,N_20312);
nor UO_984 (O_984,N_19370,N_22580);
nand UO_985 (O_985,N_24777,N_21151);
or UO_986 (O_986,N_23927,N_23703);
or UO_987 (O_987,N_19009,N_19425);
nand UO_988 (O_988,N_22074,N_19162);
nor UO_989 (O_989,N_19708,N_20944);
xnor UO_990 (O_990,N_19792,N_19610);
nor UO_991 (O_991,N_19123,N_21707);
nand UO_992 (O_992,N_20804,N_23771);
and UO_993 (O_993,N_19687,N_18962);
xnor UO_994 (O_994,N_24690,N_19169);
nor UO_995 (O_995,N_20355,N_20977);
nand UO_996 (O_996,N_22524,N_23712);
or UO_997 (O_997,N_23060,N_23167);
nor UO_998 (O_998,N_21279,N_20490);
xor UO_999 (O_999,N_21727,N_23590);
nor UO_1000 (O_1000,N_21321,N_21155);
or UO_1001 (O_1001,N_24840,N_21912);
xnor UO_1002 (O_1002,N_21465,N_22223);
nor UO_1003 (O_1003,N_21679,N_21284);
nor UO_1004 (O_1004,N_21806,N_23866);
or UO_1005 (O_1005,N_23049,N_22393);
or UO_1006 (O_1006,N_23549,N_24356);
nor UO_1007 (O_1007,N_20524,N_20555);
or UO_1008 (O_1008,N_19893,N_19880);
nor UO_1009 (O_1009,N_24082,N_19142);
and UO_1010 (O_1010,N_21953,N_21548);
and UO_1011 (O_1011,N_19158,N_24595);
nand UO_1012 (O_1012,N_20066,N_21559);
or UO_1013 (O_1013,N_22133,N_18903);
nor UO_1014 (O_1014,N_21079,N_22002);
and UO_1015 (O_1015,N_22100,N_22232);
and UO_1016 (O_1016,N_24623,N_23547);
and UO_1017 (O_1017,N_22591,N_20157);
nor UO_1018 (O_1018,N_20511,N_20040);
and UO_1019 (O_1019,N_23433,N_19932);
and UO_1020 (O_1020,N_21963,N_20616);
or UO_1021 (O_1021,N_19413,N_20683);
nand UO_1022 (O_1022,N_19323,N_19364);
nand UO_1023 (O_1023,N_20517,N_20848);
nor UO_1024 (O_1024,N_21571,N_21974);
and UO_1025 (O_1025,N_20324,N_21350);
xor UO_1026 (O_1026,N_20744,N_23900);
or UO_1027 (O_1027,N_22576,N_22761);
or UO_1028 (O_1028,N_19774,N_22250);
or UO_1029 (O_1029,N_21636,N_18759);
and UO_1030 (O_1030,N_21695,N_21939);
or UO_1031 (O_1031,N_18857,N_19761);
nor UO_1032 (O_1032,N_24798,N_20774);
or UO_1033 (O_1033,N_19699,N_21150);
or UO_1034 (O_1034,N_19450,N_19831);
xnor UO_1035 (O_1035,N_19040,N_23272);
nand UO_1036 (O_1036,N_22514,N_21112);
nor UO_1037 (O_1037,N_20847,N_21472);
nand UO_1038 (O_1038,N_20419,N_21567);
and UO_1039 (O_1039,N_22888,N_20738);
xor UO_1040 (O_1040,N_24569,N_22677);
xnor UO_1041 (O_1041,N_24856,N_19015);
nand UO_1042 (O_1042,N_24912,N_21696);
or UO_1043 (O_1043,N_19147,N_23191);
and UO_1044 (O_1044,N_24920,N_21051);
nand UO_1045 (O_1045,N_20960,N_19793);
nand UO_1046 (O_1046,N_24211,N_22822);
xnor UO_1047 (O_1047,N_23295,N_24267);
or UO_1048 (O_1048,N_19726,N_22823);
or UO_1049 (O_1049,N_18906,N_21263);
nor UO_1050 (O_1050,N_21426,N_24357);
xnor UO_1051 (O_1051,N_21470,N_20492);
xor UO_1052 (O_1052,N_21875,N_24907);
nand UO_1053 (O_1053,N_22430,N_23172);
and UO_1054 (O_1054,N_21886,N_21224);
xor UO_1055 (O_1055,N_19694,N_19914);
nand UO_1056 (O_1056,N_21359,N_20568);
xor UO_1057 (O_1057,N_20904,N_20913);
or UO_1058 (O_1058,N_24665,N_22689);
and UO_1059 (O_1059,N_21416,N_19242);
nor UO_1060 (O_1060,N_19515,N_21517);
and UO_1061 (O_1061,N_20144,N_20655);
nand UO_1062 (O_1062,N_24080,N_23290);
and UO_1063 (O_1063,N_21031,N_21069);
xor UO_1064 (O_1064,N_23223,N_21537);
and UO_1065 (O_1065,N_23915,N_21889);
and UO_1066 (O_1066,N_21138,N_22365);
nand UO_1067 (O_1067,N_24259,N_18976);
and UO_1068 (O_1068,N_20089,N_23358);
xnor UO_1069 (O_1069,N_23986,N_23248);
nand UO_1070 (O_1070,N_19717,N_22117);
xor UO_1071 (O_1071,N_22247,N_24339);
or UO_1072 (O_1072,N_19449,N_21602);
or UO_1073 (O_1073,N_24219,N_22661);
nor UO_1074 (O_1074,N_20909,N_19122);
nor UO_1075 (O_1075,N_20042,N_19318);
nor UO_1076 (O_1076,N_24010,N_24768);
xor UO_1077 (O_1077,N_20611,N_21677);
xnor UO_1078 (O_1078,N_23161,N_24529);
nor UO_1079 (O_1079,N_23854,N_23860);
xor UO_1080 (O_1080,N_22188,N_19861);
nor UO_1081 (O_1081,N_23760,N_20843);
and UO_1082 (O_1082,N_20029,N_21036);
nor UO_1083 (O_1083,N_24608,N_22329);
xnor UO_1084 (O_1084,N_19510,N_19155);
nand UO_1085 (O_1085,N_19430,N_22904);
nor UO_1086 (O_1086,N_20539,N_24297);
nand UO_1087 (O_1087,N_21433,N_20902);
nand UO_1088 (O_1088,N_22450,N_24754);
nand UO_1089 (O_1089,N_24802,N_21569);
nand UO_1090 (O_1090,N_22066,N_23664);
nor UO_1091 (O_1091,N_20447,N_22108);
nor UO_1092 (O_1092,N_24519,N_22716);
xnor UO_1093 (O_1093,N_21975,N_24771);
nand UO_1094 (O_1094,N_20868,N_20520);
nor UO_1095 (O_1095,N_20047,N_19662);
and UO_1096 (O_1096,N_20086,N_23460);
nor UO_1097 (O_1097,N_19812,N_19673);
xor UO_1098 (O_1098,N_22423,N_24852);
or UO_1099 (O_1099,N_20315,N_22894);
or UO_1100 (O_1100,N_19545,N_20483);
xor UO_1101 (O_1101,N_22636,N_19884);
or UO_1102 (O_1102,N_24073,N_21776);
nor UO_1103 (O_1103,N_22829,N_22573);
or UO_1104 (O_1104,N_19993,N_20407);
nor UO_1105 (O_1105,N_19325,N_22887);
nand UO_1106 (O_1106,N_24315,N_20897);
nand UO_1107 (O_1107,N_23363,N_20488);
and UO_1108 (O_1108,N_23344,N_19810);
nor UO_1109 (O_1109,N_21221,N_20288);
or UO_1110 (O_1110,N_23301,N_20213);
or UO_1111 (O_1111,N_24691,N_24636);
nor UO_1112 (O_1112,N_24134,N_23723);
xnor UO_1113 (O_1113,N_20326,N_23589);
nor UO_1114 (O_1114,N_20174,N_22607);
or UO_1115 (O_1115,N_20093,N_19397);
xnor UO_1116 (O_1116,N_23533,N_21638);
nor UO_1117 (O_1117,N_19584,N_23269);
nand UO_1118 (O_1118,N_19356,N_22586);
or UO_1119 (O_1119,N_21060,N_23018);
and UO_1120 (O_1120,N_20941,N_20560);
nand UO_1121 (O_1121,N_20952,N_19418);
or UO_1122 (O_1122,N_20166,N_21915);
nor UO_1123 (O_1123,N_19718,N_21304);
or UO_1124 (O_1124,N_22942,N_24288);
nand UO_1125 (O_1125,N_20898,N_20346);
nor UO_1126 (O_1126,N_21213,N_21577);
nor UO_1127 (O_1127,N_20427,N_23343);
nor UO_1128 (O_1128,N_21705,N_24493);
or UO_1129 (O_1129,N_21738,N_24726);
xnor UO_1130 (O_1130,N_22023,N_21406);
nand UO_1131 (O_1131,N_21413,N_23340);
xor UO_1132 (O_1132,N_21794,N_21694);
nor UO_1133 (O_1133,N_21265,N_22506);
nand UO_1134 (O_1134,N_22975,N_24012);
nand UO_1135 (O_1135,N_19024,N_19561);
nor UO_1136 (O_1136,N_22221,N_19205);
or UO_1137 (O_1137,N_22475,N_23777);
nor UO_1138 (O_1138,N_19347,N_19738);
xnor UO_1139 (O_1139,N_20426,N_18965);
nand UO_1140 (O_1140,N_21746,N_23318);
or UO_1141 (O_1141,N_23950,N_24599);
nand UO_1142 (O_1142,N_24905,N_22001);
nand UO_1143 (O_1143,N_21766,N_20602);
or UO_1144 (O_1144,N_21264,N_20509);
nand UO_1145 (O_1145,N_20465,N_22917);
nand UO_1146 (O_1146,N_18908,N_21911);
nand UO_1147 (O_1147,N_19579,N_19170);
nor UO_1148 (O_1148,N_19190,N_22535);
nand UO_1149 (O_1149,N_23805,N_24547);
xnor UO_1150 (O_1150,N_22061,N_23809);
or UO_1151 (O_1151,N_20132,N_20713);
nand UO_1152 (O_1152,N_24921,N_19038);
or UO_1153 (O_1153,N_19006,N_20875);
xor UO_1154 (O_1154,N_23429,N_20999);
nor UO_1155 (O_1155,N_21578,N_22974);
and UO_1156 (O_1156,N_24014,N_20997);
or UO_1157 (O_1157,N_20204,N_24488);
or UO_1158 (O_1158,N_20964,N_21175);
nand UO_1159 (O_1159,N_21836,N_20234);
nor UO_1160 (O_1160,N_21666,N_20276);
xor UO_1161 (O_1161,N_23639,N_24303);
or UO_1162 (O_1162,N_19021,N_23143);
xnor UO_1163 (O_1163,N_19634,N_24022);
and UO_1164 (O_1164,N_21599,N_21322);
nor UO_1165 (O_1165,N_20890,N_22352);
and UO_1166 (O_1166,N_24716,N_22368);
nand UO_1167 (O_1167,N_19764,N_24892);
nor UO_1168 (O_1168,N_24264,N_19869);
or UO_1169 (O_1169,N_21192,N_21361);
nand UO_1170 (O_1170,N_20178,N_22456);
nand UO_1171 (O_1171,N_24634,N_21649);
nand UO_1172 (O_1172,N_22156,N_20575);
and UO_1173 (O_1173,N_19213,N_23730);
nand UO_1174 (O_1174,N_19083,N_21400);
xor UO_1175 (O_1175,N_24065,N_23062);
xnor UO_1176 (O_1176,N_18782,N_21267);
xnor UO_1177 (O_1177,N_23693,N_21095);
nor UO_1178 (O_1178,N_20149,N_21936);
xor UO_1179 (O_1179,N_19927,N_21749);
nand UO_1180 (O_1180,N_21220,N_21945);
nor UO_1181 (O_1181,N_19385,N_23792);
and UO_1182 (O_1182,N_20109,N_19216);
nand UO_1183 (O_1183,N_24301,N_19702);
and UO_1184 (O_1184,N_21968,N_19224);
nand UO_1185 (O_1185,N_20797,N_21919);
or UO_1186 (O_1186,N_22285,N_21055);
nand UO_1187 (O_1187,N_18917,N_19159);
or UO_1188 (O_1188,N_22760,N_19795);
nand UO_1189 (O_1189,N_19842,N_21576);
and UO_1190 (O_1190,N_18858,N_22327);
nand UO_1191 (O_1191,N_24131,N_23428);
xnor UO_1192 (O_1192,N_20369,N_19636);
nand UO_1193 (O_1193,N_21745,N_23387);
xor UO_1194 (O_1194,N_22218,N_20590);
nor UO_1195 (O_1195,N_23124,N_20966);
and UO_1196 (O_1196,N_24083,N_22104);
or UO_1197 (O_1197,N_23262,N_24117);
nor UO_1198 (O_1198,N_24319,N_20604);
nand UO_1199 (O_1199,N_22191,N_22610);
or UO_1200 (O_1200,N_21683,N_21398);
nor UO_1201 (O_1201,N_19471,N_20302);
xnor UO_1202 (O_1202,N_23286,N_22821);
nor UO_1203 (O_1203,N_23071,N_22778);
xor UO_1204 (O_1204,N_23352,N_21181);
nor UO_1205 (O_1205,N_24993,N_21021);
xor UO_1206 (O_1206,N_19331,N_22134);
xnor UO_1207 (O_1207,N_19266,N_23454);
nand UO_1208 (O_1208,N_20140,N_20092);
nand UO_1209 (O_1209,N_19237,N_19684);
and UO_1210 (O_1210,N_19238,N_24855);
or UO_1211 (O_1211,N_23350,N_20606);
xor UO_1212 (O_1212,N_24991,N_24376);
nor UO_1213 (O_1213,N_19153,N_21779);
nor UO_1214 (O_1214,N_20448,N_21805);
and UO_1215 (O_1215,N_24934,N_24906);
and UO_1216 (O_1216,N_20755,N_23654);
or UO_1217 (O_1217,N_23749,N_20884);
or UO_1218 (O_1218,N_20912,N_20281);
or UO_1219 (O_1219,N_18815,N_22638);
or UO_1220 (O_1220,N_22547,N_24813);
nand UO_1221 (O_1221,N_23886,N_23571);
and UO_1222 (O_1222,N_23758,N_23618);
xor UO_1223 (O_1223,N_22641,N_20356);
xor UO_1224 (O_1224,N_19706,N_24347);
nand UO_1225 (O_1225,N_20119,N_23934);
nand UO_1226 (O_1226,N_20248,N_21870);
and UO_1227 (O_1227,N_23633,N_20129);
nor UO_1228 (O_1228,N_21667,N_23743);
nand UO_1229 (O_1229,N_18888,N_21634);
or UO_1230 (O_1230,N_22241,N_21543);
or UO_1231 (O_1231,N_23424,N_19401);
xnor UO_1232 (O_1232,N_22701,N_24949);
or UO_1233 (O_1233,N_19005,N_23656);
or UO_1234 (O_1234,N_19402,N_23378);
nor UO_1235 (O_1235,N_24728,N_24564);
xor UO_1236 (O_1236,N_23969,N_19262);
nor UO_1237 (O_1237,N_21166,N_22890);
xor UO_1238 (O_1238,N_23366,N_22472);
xnor UO_1239 (O_1239,N_20872,N_24770);
nand UO_1240 (O_1240,N_19218,N_21113);
and UO_1241 (O_1241,N_20464,N_23737);
or UO_1242 (O_1242,N_22913,N_22482);
xor UO_1243 (O_1243,N_24558,N_20702);
nor UO_1244 (O_1244,N_19753,N_20077);
nand UO_1245 (O_1245,N_21768,N_24677);
xor UO_1246 (O_1246,N_23597,N_19020);
xnor UO_1247 (O_1247,N_23708,N_24956);
xor UO_1248 (O_1248,N_22722,N_23520);
and UO_1249 (O_1249,N_18752,N_23408);
nor UO_1250 (O_1250,N_18756,N_19771);
and UO_1251 (O_1251,N_22411,N_23151);
nor UO_1252 (O_1252,N_20955,N_20924);
xor UO_1253 (O_1253,N_22200,N_19897);
nor UO_1254 (O_1254,N_22153,N_21674);
or UO_1255 (O_1255,N_23660,N_23111);
nor UO_1256 (O_1256,N_24359,N_23177);
nand UO_1257 (O_1257,N_23113,N_24898);
xor UO_1258 (O_1258,N_24075,N_23739);
and UO_1259 (O_1259,N_19691,N_19082);
and UO_1260 (O_1260,N_21993,N_24799);
or UO_1261 (O_1261,N_19511,N_22452);
or UO_1262 (O_1262,N_24692,N_20663);
nor UO_1263 (O_1263,N_21283,N_22594);
and UO_1264 (O_1264,N_22959,N_23692);
and UO_1265 (O_1265,N_22407,N_18993);
nor UO_1266 (O_1266,N_19245,N_20143);
xor UO_1267 (O_1267,N_20839,N_22418);
nor UO_1268 (O_1268,N_21687,N_19241);
and UO_1269 (O_1269,N_22281,N_22719);
or UO_1270 (O_1270,N_22276,N_22875);
and UO_1271 (O_1271,N_21328,N_21457);
or UO_1272 (O_1272,N_19378,N_22113);
xor UO_1273 (O_1273,N_23848,N_24338);
or UO_1274 (O_1274,N_23813,N_21114);
and UO_1275 (O_1275,N_24291,N_20392);
and UO_1276 (O_1276,N_22171,N_21659);
and UO_1277 (O_1277,N_20577,N_24932);
and UO_1278 (O_1278,N_22114,N_21853);
nand UO_1279 (O_1279,N_21499,N_22928);
nor UO_1280 (O_1280,N_20414,N_19981);
or UO_1281 (O_1281,N_22361,N_24858);
nor UO_1282 (O_1282,N_23791,N_22799);
and UO_1283 (O_1283,N_20073,N_23935);
and UO_1284 (O_1284,N_20515,N_24416);
and UO_1285 (O_1285,N_23648,N_20987);
xnor UO_1286 (O_1286,N_21538,N_19524);
nor UO_1287 (O_1287,N_21914,N_20268);
nor UO_1288 (O_1288,N_24276,N_20815);
and UO_1289 (O_1289,N_20545,N_21233);
nor UO_1290 (O_1290,N_23726,N_21268);
xor UO_1291 (O_1291,N_20644,N_22425);
nand UO_1292 (O_1292,N_21473,N_19671);
nor UO_1293 (O_1293,N_21763,N_22599);
or UO_1294 (O_1294,N_20599,N_22745);
and UO_1295 (O_1295,N_23431,N_23770);
and UO_1296 (O_1296,N_23668,N_20017);
or UO_1297 (O_1297,N_23686,N_19541);
nand UO_1298 (O_1298,N_19116,N_20207);
nand UO_1299 (O_1299,N_22259,N_19299);
and UO_1300 (O_1300,N_24637,N_22222);
nor UO_1301 (O_1301,N_23365,N_22659);
nor UO_1302 (O_1302,N_21803,N_19277);
nor UO_1303 (O_1303,N_24112,N_19635);
nand UO_1304 (O_1304,N_22041,N_21169);
xor UO_1305 (O_1305,N_23796,N_19124);
and UO_1306 (O_1306,N_24579,N_24273);
xnor UO_1307 (O_1307,N_23852,N_20506);
nor UO_1308 (O_1308,N_22743,N_23534);
xnor UO_1309 (O_1309,N_24616,N_20630);
xnor UO_1310 (O_1310,N_20894,N_24255);
nand UO_1311 (O_1311,N_19815,N_22570);
nand UO_1312 (O_1312,N_22394,N_23259);
nor UO_1313 (O_1313,N_19656,N_19486);
and UO_1314 (O_1314,N_19114,N_24298);
nand UO_1315 (O_1315,N_19564,N_23569);
or UO_1316 (O_1316,N_19167,N_20907);
or UO_1317 (O_1317,N_24644,N_23478);
nor UO_1318 (O_1318,N_19315,N_23136);
nand UO_1319 (O_1319,N_21940,N_22649);
xor UO_1320 (O_1320,N_23346,N_21314);
or UO_1321 (O_1321,N_19093,N_22121);
xnor UO_1322 (O_1322,N_22955,N_20988);
nand UO_1323 (O_1323,N_22963,N_22442);
and UO_1324 (O_1324,N_19026,N_23902);
and UO_1325 (O_1325,N_18780,N_23719);
xor UO_1326 (O_1326,N_24331,N_22518);
nor UO_1327 (O_1327,N_21414,N_20384);
nand UO_1328 (O_1328,N_19954,N_22256);
nand UO_1329 (O_1329,N_23917,N_19521);
or UO_1330 (O_1330,N_22674,N_18808);
and UO_1331 (O_1331,N_19497,N_18847);
xnor UO_1332 (O_1332,N_19600,N_23646);
xor UO_1333 (O_1333,N_21270,N_23447);
nor UO_1334 (O_1334,N_23713,N_23009);
and UO_1335 (O_1335,N_18988,N_20416);
nor UO_1336 (O_1336,N_23845,N_20298);
or UO_1337 (O_1337,N_23832,N_24808);
nor UO_1338 (O_1338,N_20867,N_23016);
or UO_1339 (O_1339,N_23265,N_20836);
and UO_1340 (O_1340,N_22480,N_23120);
nand UO_1341 (O_1341,N_24536,N_19539);
nor UO_1342 (O_1342,N_21401,N_22071);
nand UO_1343 (O_1343,N_19650,N_19477);
nor UO_1344 (O_1344,N_24530,N_24889);
nor UO_1345 (O_1345,N_19455,N_21789);
nor UO_1346 (O_1346,N_24085,N_22086);
xor UO_1347 (O_1347,N_22237,N_22744);
and UO_1348 (O_1348,N_20790,N_22187);
nor UO_1349 (O_1349,N_21756,N_18840);
or UO_1350 (O_1350,N_19890,N_20622);
nand UO_1351 (O_1351,N_22598,N_20125);
and UO_1352 (O_1352,N_21951,N_19829);
nor UO_1353 (O_1353,N_23840,N_20113);
or UO_1354 (O_1354,N_21262,N_24164);
nor UO_1355 (O_1355,N_20236,N_23604);
or UO_1356 (O_1356,N_18773,N_22970);
nor UO_1357 (O_1357,N_19043,N_19944);
or UO_1358 (O_1358,N_20306,N_21422);
and UO_1359 (O_1359,N_23684,N_22292);
or UO_1360 (O_1360,N_24767,N_19737);
and UO_1361 (O_1361,N_20269,N_24378);
xor UO_1362 (O_1362,N_20709,N_22350);
nand UO_1363 (O_1363,N_20232,N_22527);
nor UO_1364 (O_1364,N_23168,N_23677);
xor UO_1365 (O_1365,N_22248,N_22435);
nor UO_1366 (O_1366,N_20728,N_24628);
nor UO_1367 (O_1367,N_23237,N_19080);
nor UO_1368 (O_1368,N_21629,N_21641);
nand UO_1369 (O_1369,N_22353,N_24645);
and UO_1370 (O_1370,N_23224,N_19176);
nor UO_1371 (O_1371,N_21135,N_20814);
and UO_1372 (O_1372,N_19820,N_19453);
nand UO_1373 (O_1373,N_19937,N_22998);
and UO_1374 (O_1374,N_19722,N_23450);
or UO_1375 (O_1375,N_20277,N_19664);
nor UO_1376 (O_1376,N_24606,N_20812);
nor UO_1377 (O_1377,N_19208,N_19365);
nand UO_1378 (O_1378,N_19940,N_19729);
nand UO_1379 (O_1379,N_19051,N_22461);
nor UO_1380 (O_1380,N_24226,N_24633);
xnor UO_1381 (O_1381,N_22642,N_19258);
xor UO_1382 (O_1382,N_21581,N_20658);
and UO_1383 (O_1383,N_19833,N_20981);
or UO_1384 (O_1384,N_21100,N_19099);
and UO_1385 (O_1385,N_24801,N_24413);
and UO_1386 (O_1386,N_20264,N_24648);
nor UO_1387 (O_1387,N_24035,N_24687);
xnor UO_1388 (O_1388,N_18804,N_23307);
nor UO_1389 (O_1389,N_19226,N_21493);
and UO_1390 (O_1390,N_22534,N_21662);
nand UO_1391 (O_1391,N_23392,N_22759);
or UO_1392 (O_1392,N_20360,N_22385);
nand UO_1393 (O_1393,N_22102,N_21362);
nand UO_1394 (O_1394,N_20716,N_24620);
or UO_1395 (O_1395,N_21259,N_20373);
and UO_1396 (O_1396,N_20341,N_20256);
nor UO_1397 (O_1397,N_21235,N_19767);
xor UO_1398 (O_1398,N_22046,N_20290);
and UO_1399 (O_1399,N_21891,N_21315);
or UO_1400 (O_1400,N_22957,N_22947);
or UO_1401 (O_1401,N_24807,N_22771);
xnor UO_1402 (O_1402,N_24941,N_23949);
xnor UO_1403 (O_1403,N_20474,N_19943);
and UO_1404 (O_1404,N_20724,N_24886);
xnor UO_1405 (O_1405,N_23072,N_20206);
xnor UO_1406 (O_1406,N_22453,N_20285);
xor UO_1407 (O_1407,N_20521,N_18959);
nor UO_1408 (O_1408,N_21159,N_18833);
or UO_1409 (O_1409,N_21786,N_23988);
nor UO_1410 (O_1410,N_20021,N_23808);
xnor UO_1411 (O_1411,N_19859,N_18915);
or UO_1412 (O_1412,N_20338,N_22951);
xor UO_1413 (O_1413,N_22408,N_20530);
or UO_1414 (O_1414,N_22715,N_18864);
or UO_1415 (O_1415,N_21206,N_20479);
nand UO_1416 (O_1416,N_23801,N_19628);
nand UO_1417 (O_1417,N_22780,N_21381);
or UO_1418 (O_1418,N_22691,N_22022);
nand UO_1419 (O_1419,N_24822,N_22079);
nor UO_1420 (O_1420,N_22055,N_21410);
nand UO_1421 (O_1421,N_24944,N_19805);
nand UO_1422 (O_1422,N_23763,N_21122);
or UO_1423 (O_1423,N_20699,N_21528);
nand UO_1424 (O_1424,N_23356,N_19612);
and UO_1425 (O_1425,N_23037,N_23199);
nand UO_1426 (O_1426,N_18811,N_21319);
nor UO_1427 (O_1427,N_20994,N_22792);
and UO_1428 (O_1428,N_20798,N_24018);
xor UO_1429 (O_1429,N_21846,N_24103);
and UO_1430 (O_1430,N_20188,N_21177);
xor UO_1431 (O_1431,N_21396,N_22918);
or UO_1432 (O_1432,N_20610,N_21793);
nor UO_1433 (O_1433,N_18984,N_23360);
and UO_1434 (O_1434,N_20391,N_22766);
and UO_1435 (O_1435,N_24584,N_20696);
or UO_1436 (O_1436,N_22797,N_22862);
xnor UO_1437 (O_1437,N_19921,N_24793);
or UO_1438 (O_1438,N_21144,N_20792);
and UO_1439 (O_1439,N_23205,N_19876);
and UO_1440 (O_1440,N_23330,N_19689);
nor UO_1441 (O_1441,N_23417,N_21905);
nor UO_1442 (O_1442,N_20603,N_22939);
nor UO_1443 (O_1443,N_24038,N_23065);
and UO_1444 (O_1444,N_20561,N_20747);
nor UO_1445 (O_1445,N_21985,N_21474);
and UO_1446 (O_1446,N_21902,N_20485);
and UO_1447 (O_1447,N_22478,N_20214);
xor UO_1448 (O_1448,N_22346,N_24953);
xor UO_1449 (O_1449,N_19779,N_22477);
nand UO_1450 (O_1450,N_21195,N_24939);
nor UO_1451 (O_1451,N_20838,N_20880);
or UO_1452 (O_1452,N_23560,N_23853);
xnor UO_1453 (O_1453,N_19739,N_19641);
and UO_1454 (O_1454,N_21272,N_23793);
nor UO_1455 (O_1455,N_24593,N_22362);
xor UO_1456 (O_1456,N_20871,N_20685);
xnor UO_1457 (O_1457,N_24977,N_21851);
nor UO_1458 (O_1458,N_22938,N_22750);
nand UO_1459 (O_1459,N_19680,N_19352);
or UO_1460 (O_1460,N_20293,N_19186);
or UO_1461 (O_1461,N_22460,N_24512);
nor UO_1462 (O_1462,N_24447,N_21978);
nand UO_1463 (O_1463,N_20841,N_24163);
xor UO_1464 (O_1464,N_19209,N_23375);
nand UO_1465 (O_1465,N_22600,N_20926);
and UO_1466 (O_1466,N_20857,N_23768);
nor UO_1467 (O_1467,N_20494,N_21140);
nand UO_1468 (O_1468,N_18776,N_22324);
nor UO_1469 (O_1469,N_21278,N_21947);
xor UO_1470 (O_1470,N_23403,N_22732);
xor UO_1471 (O_1471,N_20449,N_20233);
or UO_1472 (O_1472,N_19686,N_24954);
and UO_1473 (O_1473,N_24469,N_24102);
xnor UO_1474 (O_1474,N_23040,N_24821);
nand UO_1475 (O_1475,N_20862,N_22227);
nor UO_1476 (O_1476,N_23292,N_18848);
xor UO_1477 (O_1477,N_20771,N_21461);
and UO_1478 (O_1478,N_20947,N_21423);
or UO_1479 (O_1479,N_21310,N_23380);
nand UO_1480 (O_1480,N_24867,N_24332);
nand UO_1481 (O_1481,N_23398,N_23305);
nor UO_1482 (O_1482,N_24823,N_19554);
xnor UO_1483 (O_1483,N_20007,N_24930);
nand UO_1484 (O_1484,N_20605,N_22266);
and UO_1485 (O_1485,N_19933,N_23171);
xnor UO_1486 (O_1486,N_24345,N_20102);
or UO_1487 (O_1487,N_24583,N_19791);
nor UO_1488 (O_1488,N_21807,N_24281);
and UO_1489 (O_1489,N_23000,N_18935);
nor UO_1490 (O_1490,N_22485,N_23357);
xor UO_1491 (O_1491,N_19950,N_20441);
nor UO_1492 (O_1492,N_24499,N_18856);
or UO_1493 (O_1493,N_19168,N_19620);
nand UO_1494 (O_1494,N_20554,N_19920);
nor UO_1495 (O_1495,N_19781,N_24904);
nand UO_1496 (O_1496,N_19362,N_18953);
nor UO_1497 (O_1497,N_21530,N_20536);
or UO_1498 (O_1498,N_21586,N_24682);
and UO_1499 (O_1499,N_22369,N_21888);
xor UO_1500 (O_1500,N_21110,N_22614);
xnor UO_1501 (O_1501,N_19874,N_22177);
and UO_1502 (O_1502,N_19928,N_24466);
xnor UO_1503 (O_1503,N_19456,N_24743);
xor UO_1504 (O_1504,N_20309,N_24859);
and UO_1505 (O_1505,N_24528,N_21039);
nand UO_1506 (O_1506,N_22370,N_18786);
xnor UO_1507 (O_1507,N_23078,N_24918);
or UO_1508 (O_1508,N_22458,N_20905);
nor UO_1509 (O_1509,N_20310,N_20522);
and UO_1510 (O_1510,N_23666,N_19312);
xnor UO_1511 (O_1511,N_19489,N_23951);
nand UO_1512 (O_1512,N_20967,N_18869);
nor UO_1513 (O_1513,N_22540,N_22139);
and UO_1514 (O_1514,N_21869,N_23484);
and UO_1515 (O_1515,N_19604,N_21357);
nor UO_1516 (O_1516,N_22788,N_22167);
nor UO_1517 (O_1517,N_24475,N_24661);
nor UO_1518 (O_1518,N_22965,N_20707);
xnor UO_1519 (O_1519,N_24274,N_23701);
xnor UO_1520 (O_1520,N_20751,N_19520);
xor UO_1521 (O_1521,N_23553,N_20886);
xor UO_1522 (O_1522,N_24017,N_23422);
nor UO_1523 (O_1523,N_21437,N_22406);
and UO_1524 (O_1524,N_21367,N_19509);
nor UO_1525 (O_1525,N_23527,N_20532);
nor UO_1526 (O_1526,N_20854,N_21464);
nand UO_1527 (O_1527,N_18875,N_19172);
and UO_1528 (O_1528,N_22429,N_19387);
and UO_1529 (O_1529,N_22401,N_19274);
nand UO_1530 (O_1530,N_24358,N_20088);
nor UO_1531 (O_1531,N_24962,N_22412);
or UO_1532 (O_1532,N_23202,N_19103);
and UO_1533 (O_1533,N_24563,N_23907);
nand UO_1534 (O_1534,N_24952,N_20689);
and UO_1535 (O_1535,N_21411,N_21639);
or UO_1536 (O_1536,N_23130,N_18910);
xnor UO_1537 (O_1537,N_18844,N_23599);
or UO_1538 (O_1538,N_19068,N_23979);
nor UO_1539 (O_1539,N_24019,N_20026);
and UO_1540 (O_1540,N_24655,N_23028);
xor UO_1541 (O_1541,N_23898,N_24557);
xor UO_1542 (O_1542,N_23255,N_21622);
nand UO_1543 (O_1543,N_23562,N_24788);
nor UO_1544 (O_1544,N_22021,N_23361);
and UO_1545 (O_1545,N_19690,N_20980);
nor UO_1546 (O_1546,N_20335,N_19668);
and UO_1547 (O_1547,N_22245,N_23624);
and UO_1548 (O_1548,N_20723,N_23865);
xor UO_1549 (O_1549,N_24151,N_22790);
nand UO_1550 (O_1550,N_24881,N_22985);
nand UO_1551 (O_1551,N_24795,N_19161);
nor UO_1552 (O_1552,N_19071,N_21799);
nand UO_1553 (O_1553,N_22804,N_24462);
nor UO_1554 (O_1554,N_22073,N_20019);
nand UO_1555 (O_1555,N_20091,N_20900);
nand UO_1556 (O_1556,N_22052,N_24379);
nor UO_1557 (O_1557,N_22874,N_20930);
nor UO_1558 (O_1558,N_18850,N_24334);
and UO_1559 (O_1559,N_21397,N_23901);
nor UO_1560 (O_1560,N_24542,N_22291);
or UO_1561 (O_1561,N_19566,N_23705);
and UO_1562 (O_1562,N_22136,N_21160);
nand UO_1563 (O_1563,N_23867,N_21109);
or UO_1564 (O_1564,N_23995,N_24571);
and UO_1565 (O_1565,N_22014,N_18967);
xnor UO_1566 (O_1566,N_23473,N_22665);
xnor UO_1567 (O_1567,N_21590,N_21153);
nand UO_1568 (O_1568,N_24833,N_20247);
or UO_1569 (O_1569,N_20038,N_23095);
nor UO_1570 (O_1570,N_24712,N_21515);
and UO_1571 (O_1571,N_22169,N_22525);
nor UO_1572 (O_1572,N_19551,N_23629);
and UO_1573 (O_1573,N_24629,N_23107);
nor UO_1574 (O_1574,N_20254,N_24036);
nor UO_1575 (O_1575,N_24299,N_20686);
xor UO_1576 (O_1576,N_23894,N_23964);
xnor UO_1577 (O_1577,N_19785,N_20948);
nor UO_1578 (O_1578,N_22712,N_20674);
or UO_1579 (O_1579,N_21184,N_19953);
nor UO_1580 (O_1580,N_24734,N_23810);
nor UO_1581 (O_1581,N_20617,N_22528);
or UO_1582 (O_1582,N_22278,N_20235);
nor UO_1583 (O_1583,N_21273,N_21266);
nand UO_1584 (O_1584,N_20100,N_23967);
or UO_1585 (O_1585,N_22172,N_23952);
and UO_1586 (O_1586,N_24093,N_22557);
or UO_1587 (O_1587,N_21990,N_18798);
nor UO_1588 (O_1588,N_21001,N_20929);
nor UO_1589 (O_1589,N_20734,N_20079);
nor UO_1590 (O_1590,N_21253,N_21549);
nor UO_1591 (O_1591,N_23567,N_19798);
xnor UO_1592 (O_1592,N_24568,N_21896);
or UO_1593 (O_1593,N_20179,N_20739);
xnor UO_1594 (O_1594,N_18849,N_22983);
nand UO_1595 (O_1595,N_22906,N_23843);
and UO_1596 (O_1596,N_22523,N_22130);
xnor UO_1597 (O_1597,N_23453,N_20330);
nor UO_1598 (O_1598,N_19597,N_24860);
and UO_1599 (O_1599,N_22603,N_20222);
nand UO_1600 (O_1600,N_24044,N_22676);
nor UO_1601 (O_1601,N_23557,N_22885);
xor UO_1602 (O_1602,N_22271,N_20361);
xnor UO_1603 (O_1603,N_24961,N_21703);
nor UO_1604 (O_1604,N_22730,N_24217);
and UO_1605 (O_1605,N_20802,N_24198);
or UO_1606 (O_1606,N_19259,N_24353);
nor UO_1607 (O_1607,N_24109,N_23818);
nor UO_1608 (O_1608,N_20082,N_22501);
and UO_1609 (O_1609,N_20218,N_20817);
nor UO_1610 (O_1610,N_19458,N_24543);
nor UO_1611 (O_1611,N_23367,N_23828);
nor UO_1612 (O_1612,N_23750,N_23411);
xnor UO_1613 (O_1613,N_20873,N_23074);
xnor UO_1614 (O_1614,N_22125,N_20895);
nand UO_1615 (O_1615,N_19138,N_22112);
or UO_1616 (O_1616,N_19529,N_21594);
nor UO_1617 (O_1617,N_24879,N_20197);
or UO_1618 (O_1618,N_19974,N_22990);
and UO_1619 (O_1619,N_21212,N_21858);
nand UO_1620 (O_1620,N_20137,N_22563);
or UO_1621 (O_1621,N_20621,N_24424);
and UO_1622 (O_1622,N_20348,N_19073);
nor UO_1623 (O_1623,N_23377,N_22378);
nand UO_1624 (O_1624,N_22444,N_20016);
nand UO_1625 (O_1625,N_20022,N_24725);
and UO_1626 (O_1626,N_22907,N_23619);
xor UO_1627 (O_1627,N_20099,N_21302);
nor UO_1628 (O_1628,N_19437,N_22650);
xnor UO_1629 (O_1629,N_19710,N_20807);
or UO_1630 (O_1630,N_21881,N_21168);
nand UO_1631 (O_1631,N_20766,N_21510);
and UO_1632 (O_1632,N_21374,N_23033);
or UO_1633 (O_1633,N_19126,N_19004);
nor UO_1634 (O_1634,N_19772,N_20499);
nand UO_1635 (O_1635,N_24490,N_24943);
or UO_1636 (O_1636,N_19251,N_24452);
nand UO_1637 (O_1637,N_20638,N_22601);
xor UO_1638 (O_1638,N_22546,N_22338);
xnor UO_1639 (O_1639,N_22434,N_20580);
nor UO_1640 (O_1640,N_19827,N_22980);
nand UO_1641 (O_1641,N_21275,N_21813);
or UO_1642 (O_1642,N_22815,N_24735);
and UO_1643 (O_1643,N_24061,N_19622);
nor UO_1644 (O_1644,N_24340,N_20614);
nor UO_1645 (O_1645,N_22045,N_20451);
or UO_1646 (O_1646,N_21685,N_19115);
nor UO_1647 (O_1647,N_20420,N_24021);
nand UO_1648 (O_1648,N_19840,N_20916);
or UO_1649 (O_1649,N_23063,N_23574);
xnor UO_1650 (O_1650,N_21837,N_19811);
xnor UO_1651 (O_1651,N_22015,N_19333);
nor UO_1652 (O_1652,N_23524,N_23825);
and UO_1653 (O_1653,N_21145,N_24409);
nand UO_1654 (O_1654,N_21532,N_18862);
xor UO_1655 (O_1655,N_22581,N_22468);
or UO_1656 (O_1656,N_19010,N_19298);
or UO_1657 (O_1657,N_24425,N_22185);
and UO_1658 (O_1658,N_21164,N_20864);
nand UO_1659 (O_1659,N_23396,N_19008);
or UO_1660 (O_1660,N_21208,N_23635);
or UO_1661 (O_1661,N_24498,N_20540);
and UO_1662 (O_1662,N_23585,N_21078);
nor UO_1663 (O_1663,N_21625,N_19210);
and UO_1664 (O_1664,N_24181,N_24245);
nor UO_1665 (O_1665,N_22035,N_19342);
nand UO_1666 (O_1666,N_24352,N_22783);
nor UO_1667 (O_1667,N_19697,N_20793);
xnor UO_1668 (O_1668,N_19813,N_19304);
xnor UO_1669 (O_1669,N_24970,N_23192);
xnor UO_1670 (O_1670,N_18934,N_23842);
nand UO_1671 (O_1671,N_21854,N_19300);
xor UO_1672 (O_1672,N_19346,N_19835);
nor UO_1673 (O_1673,N_23004,N_24660);
and UO_1674 (O_1674,N_24453,N_22555);
nor UO_1675 (O_1675,N_24094,N_24316);
nand UO_1676 (O_1676,N_23186,N_22091);
nor UO_1677 (O_1677,N_20585,N_23947);
xnor UO_1678 (O_1678,N_19375,N_22161);
or UO_1679 (O_1679,N_22710,N_23206);
nor UO_1680 (O_1680,N_22010,N_19150);
or UO_1681 (O_1681,N_19338,N_23956);
nand UO_1682 (O_1682,N_23617,N_23966);
xor UO_1683 (O_1683,N_21983,N_20680);
or UO_1684 (O_1684,N_22339,N_24555);
nor UO_1685 (O_1685,N_22440,N_23264);
xor UO_1686 (O_1686,N_22152,N_21480);
or UO_1687 (O_1687,N_19067,N_21038);
xor UO_1688 (O_1688,N_23945,N_22143);
or UO_1689 (O_1689,N_24760,N_20477);
or UO_1690 (O_1690,N_24087,N_24007);
or UO_1691 (O_1691,N_22040,N_23012);
nand UO_1692 (O_1692,N_22699,N_20703);
xor UO_1693 (O_1693,N_24586,N_20889);
and UO_1694 (O_1694,N_21105,N_21269);
and UO_1695 (O_1695,N_23108,N_24473);
nand UO_1696 (O_1696,N_21223,N_24182);
xnor UO_1697 (O_1697,N_22397,N_21757);
or UO_1698 (O_1698,N_21613,N_20978);
nor UO_1699 (O_1699,N_21054,N_19987);
nor UO_1700 (O_1700,N_19016,N_19230);
nor UO_1701 (O_1701,N_20381,N_19601);
xor UO_1702 (O_1702,N_21107,N_21376);
or UO_1703 (O_1703,N_19766,N_23035);
or UO_1704 (O_1704,N_23418,N_22889);
nor UO_1705 (O_1705,N_20444,N_19501);
or UO_1706 (O_1706,N_19631,N_24601);
nand UO_1707 (O_1707,N_20108,N_19377);
xnor UO_1708 (O_1708,N_21815,N_22424);
xor UO_1709 (O_1709,N_20730,N_21371);
xor UO_1710 (O_1710,N_24507,N_23638);
xnor UO_1711 (O_1711,N_21540,N_19931);
and UO_1712 (O_1712,N_22053,N_23233);
and UO_1713 (O_1713,N_19645,N_20291);
xnor UO_1714 (O_1714,N_24611,N_24689);
xnor UO_1715 (O_1715,N_23444,N_19535);
and UO_1716 (O_1716,N_19063,N_22194);
xor UO_1717 (O_1717,N_24693,N_24854);
nand UO_1718 (O_1718,N_24189,N_20535);
or UO_1719 (O_1719,N_23936,N_20828);
nor UO_1720 (O_1720,N_18854,N_22215);
nand UO_1721 (O_1721,N_19227,N_23210);
nand UO_1722 (O_1722,N_24419,N_22863);
nor UO_1723 (O_1723,N_20318,N_20557);
nand UO_1724 (O_1724,N_20316,N_20303);
and UO_1725 (O_1725,N_20409,N_23874);
nor UO_1726 (O_1726,N_23197,N_23029);
xnor UO_1727 (O_1727,N_21186,N_23716);
and UO_1728 (O_1728,N_24787,N_22296);
and UO_1729 (O_1729,N_19178,N_23140);
or UO_1730 (O_1730,N_21313,N_20595);
nand UO_1731 (O_1731,N_23899,N_24652);
and UO_1732 (O_1732,N_23672,N_21998);
nor UO_1733 (O_1733,N_22505,N_19460);
nand UO_1734 (O_1734,N_23257,N_18922);
and UO_1735 (O_1735,N_20705,N_24403);
and UO_1736 (O_1736,N_21111,N_21347);
or UO_1737 (O_1737,N_21425,N_24215);
nand UO_1738 (O_1738,N_19081,N_19513);
or UO_1739 (O_1739,N_21187,N_19414);
and UO_1740 (O_1740,N_18831,N_22277);
or UO_1741 (O_1741,N_24187,N_19552);
and UO_1742 (O_1742,N_19101,N_24106);
and UO_1743 (O_1743,N_21058,N_22781);
nor UO_1744 (O_1744,N_22135,N_19857);
nand UO_1745 (O_1745,N_21380,N_23162);
nand UO_1746 (O_1746,N_19821,N_23059);
xnor UO_1747 (O_1747,N_24108,N_22328);
or UO_1748 (O_1748,N_23068,N_22883);
nand UO_1749 (O_1749,N_22105,N_20457);
nor UO_1750 (O_1750,N_21089,N_21500);
and UO_1751 (O_1751,N_24973,N_24896);
xor UO_1752 (O_1752,N_19292,N_22748);
nand UO_1753 (O_1753,N_18797,N_22463);
nor UO_1754 (O_1754,N_20106,N_24478);
or UO_1755 (O_1755,N_21646,N_18877);
xor UO_1756 (O_1756,N_19814,N_18754);
nand UO_1757 (O_1757,N_19145,N_23300);
xnor UO_1758 (O_1758,N_23774,N_21820);
nor UO_1759 (O_1759,N_21099,N_24238);
nand UO_1760 (O_1760,N_23830,N_21072);
nand UO_1761 (O_1761,N_22933,N_20175);
nor UO_1762 (O_1762,N_24785,N_19415);
nor UO_1763 (O_1763,N_23362,N_24436);
and UO_1764 (O_1764,N_22572,N_21730);
or UO_1765 (O_1765,N_22964,N_19222);
nand UO_1766 (O_1766,N_20721,N_24978);
xor UO_1767 (O_1767,N_19419,N_19713);
nand UO_1768 (O_1768,N_19674,N_21209);
nor UO_1769 (O_1769,N_21593,N_19565);
nand UO_1770 (O_1770,N_20877,N_22634);
or UO_1771 (O_1771,N_19439,N_21584);
and UO_1772 (O_1772,N_22180,N_22387);
nor UO_1773 (O_1773,N_24902,N_21067);
nor UO_1774 (O_1774,N_24675,N_19003);
and UO_1775 (O_1775,N_20794,N_24260);
or UO_1776 (O_1776,N_22308,N_22333);
nor UO_1777 (O_1777,N_19089,N_21958);
or UO_1778 (O_1778,N_22763,N_21857);
and UO_1779 (O_1779,N_19120,N_19220);
nor UO_1780 (O_1780,N_22832,N_23993);
and UO_1781 (O_1781,N_20358,N_20715);
or UO_1782 (O_1782,N_20080,N_22445);
xor UO_1783 (O_1783,N_22583,N_24744);
and UO_1784 (O_1784,N_20139,N_23628);
and UO_1785 (O_1785,N_20725,N_20691);
or UO_1786 (O_1786,N_24792,N_23089);
nor UO_1787 (O_1787,N_20956,N_23372);
or UO_1788 (O_1788,N_20265,N_21097);
nor UO_1789 (O_1789,N_24283,N_19136);
nand UO_1790 (O_1790,N_19267,N_22150);
or UO_1791 (O_1791,N_18937,N_21447);
nor UO_1792 (O_1792,N_20694,N_20619);
and UO_1793 (O_1793,N_22208,N_21688);
nand UO_1794 (O_1794,N_23748,N_21351);
xor UO_1795 (O_1795,N_20938,N_20643);
and UO_1796 (O_1796,N_24592,N_24700);
nand UO_1797 (O_1797,N_22502,N_19583);
nor UO_1798 (O_1798,N_22902,N_24426);
nand UO_1799 (O_1799,N_24381,N_23017);
or UO_1800 (O_1800,N_24489,N_23985);
xnor UO_1801 (O_1801,N_21821,N_21826);
or UO_1802 (O_1802,N_22940,N_21774);
nor UO_1803 (O_1803,N_24396,N_22012);
and UO_1804 (O_1804,N_18972,N_24002);
xor UO_1805 (O_1805,N_24694,N_22678);
or UO_1806 (O_1806,N_23591,N_21012);
nor UO_1807 (O_1807,N_21229,N_20208);
or UO_1808 (O_1808,N_22076,N_22577);
and UO_1809 (O_1809,N_22597,N_22490);
nor UO_1810 (O_1810,N_24306,N_19888);
xor UO_1811 (O_1811,N_20075,N_19844);
or UO_1812 (O_1812,N_19007,N_21372);
xor UO_1813 (O_1813,N_24472,N_23280);
xor UO_1814 (O_1814,N_20359,N_24394);
and UO_1815 (O_1815,N_20859,N_24967);
nor UO_1816 (O_1816,N_19550,N_24817);
or UO_1817 (O_1817,N_20458,N_19496);
and UO_1818 (O_1818,N_19802,N_21609);
or UO_1819 (O_1819,N_24740,N_23274);
nor UO_1820 (O_1820,N_24271,N_23182);
nor UO_1821 (O_1821,N_22944,N_24779);
and UO_1822 (O_1822,N_22511,N_23253);
nor UO_1823 (O_1823,N_23486,N_21238);
and UO_1824 (O_1824,N_19174,N_18841);
and UO_1825 (O_1825,N_20070,N_20701);
nand UO_1826 (O_1826,N_21016,N_19462);
nor UO_1827 (O_1827,N_19094,N_22605);
nor UO_1828 (O_1828,N_24523,N_19606);
or UO_1829 (O_1829,N_21199,N_24474);
nor UO_1830 (O_1830,N_24063,N_21290);
or UO_1831 (O_1831,N_20566,N_22931);
nand UO_1832 (O_1832,N_19763,N_24236);
nor UO_1833 (O_1833,N_18941,N_20151);
xor UO_1834 (O_1834,N_23605,N_19109);
and UO_1835 (O_1835,N_23052,N_24979);
and UO_1836 (O_1836,N_22263,N_23326);
nand UO_1837 (O_1837,N_21293,N_23909);
or UO_1838 (O_1838,N_19860,N_19432);
or UO_1839 (O_1839,N_19678,N_23092);
xor UO_1840 (O_1840,N_24882,N_24227);
nand UO_1841 (O_1841,N_20050,N_24573);
xnor UO_1842 (O_1842,N_21832,N_24772);
or UO_1843 (O_1843,N_22700,N_19889);
or UO_1844 (O_1844,N_19885,N_22128);
or UO_1845 (O_1845,N_20582,N_20027);
nand UO_1846 (O_1846,N_19014,N_23817);
and UO_1847 (O_1847,N_19547,N_20528);
nor UO_1848 (O_1848,N_22627,N_21710);
or UO_1849 (O_1849,N_24517,N_22293);
xnor UO_1850 (O_1850,N_24947,N_21488);
xor UO_1851 (O_1851,N_19592,N_19047);
xor UO_1852 (O_1852,N_19819,N_22529);
nor UO_1853 (O_1853,N_21767,N_21243);
xnor UO_1854 (O_1854,N_21868,N_22119);
nor UO_1855 (O_1855,N_19935,N_22979);
or UO_1856 (O_1856,N_22729,N_22575);
and UO_1857 (O_1857,N_23863,N_19809);
and UO_1858 (O_1858,N_24113,N_21342);
and UO_1859 (O_1859,N_23625,N_21062);
xor UO_1860 (O_1860,N_23294,N_22553);
nor UO_1861 (O_1861,N_24270,N_23250);
xor UO_1862 (O_1862,N_19625,N_22617);
nor UO_1863 (O_1863,N_23449,N_19756);
xor UO_1864 (O_1864,N_22109,N_22796);
or UO_1865 (O_1865,N_19891,N_23790);
nor UO_1866 (O_1866,N_20918,N_21261);
or UO_1867 (O_1867,N_22673,N_23925);
nor UO_1868 (O_1868,N_23802,N_22354);
xnor UO_1869 (O_1869,N_22537,N_22398);
nor UO_1870 (O_1870,N_21824,N_23998);
and UO_1871 (O_1871,N_22315,N_22785);
nor UO_1872 (O_1872,N_22403,N_22087);
nor UO_1873 (O_1873,N_20502,N_21214);
and UO_1874 (O_1874,N_21424,N_23369);
nand UO_1875 (O_1875,N_20516,N_20261);
xnor UO_1876 (O_1876,N_21624,N_24585);
xnor UO_1877 (O_1877,N_22065,N_19494);
and UO_1878 (O_1878,N_20671,N_19540);
or UO_1879 (O_1879,N_20745,N_23053);
nor UO_1880 (O_1880,N_22178,N_20718);
xnor UO_1881 (O_1881,N_20031,N_24159);
nand UO_1882 (O_1882,N_22283,N_24679);
and UO_1883 (O_1883,N_21081,N_24458);
nand UO_1884 (O_1884,N_24095,N_19991);
nor UO_1885 (O_1885,N_23323,N_24742);
xor UO_1886 (O_1886,N_21950,N_19442);
nor UO_1887 (O_1887,N_24307,N_23621);
or UO_1888 (O_1888,N_20329,N_18945);
xor UO_1889 (O_1889,N_21475,N_21859);
and UO_1890 (O_1890,N_24582,N_23319);
nor UO_1891 (O_1891,N_21860,N_19543);
nor UO_1892 (O_1892,N_23221,N_20593);
and UO_1893 (O_1893,N_22486,N_19866);
and UO_1894 (O_1894,N_22267,N_20037);
nor UO_1895 (O_1895,N_21579,N_21468);
nor UO_1896 (O_1896,N_24539,N_22891);
and UO_1897 (O_1897,N_18940,N_21728);
xnor UO_1898 (O_1898,N_23773,N_22176);
xor UO_1899 (O_1899,N_21595,N_22141);
xnor UO_1900 (O_1900,N_20799,N_18995);
and UO_1901 (O_1901,N_19638,N_19654);
xnor UO_1902 (O_1902,N_24229,N_19022);
xnor UO_1903 (O_1903,N_24235,N_24710);
nor UO_1904 (O_1904,N_19899,N_22157);
xnor UO_1905 (O_1905,N_18914,N_24831);
or UO_1906 (O_1906,N_19560,N_23781);
and UO_1907 (O_1907,N_20750,N_23057);
xnor UO_1908 (O_1908,N_20104,N_19253);
and UO_1909 (O_1909,N_24657,N_24074);
and UO_1910 (O_1910,N_24191,N_19019);
nand UO_1911 (O_1911,N_21029,N_23541);
and UO_1912 (O_1912,N_21943,N_23270);
xnor UO_1913 (O_1913,N_24411,N_20635);
or UO_1914 (O_1914,N_24427,N_23505);
and UO_1915 (O_1915,N_19748,N_22726);
xnor UO_1916 (O_1916,N_19995,N_19199);
or UO_1917 (O_1917,N_21514,N_19503);
nor UO_1918 (O_1918,N_23086,N_19059);
nand UO_1919 (O_1919,N_18821,N_19171);
nand UO_1920 (O_1920,N_20009,N_20808);
nor UO_1921 (O_1921,N_18761,N_21601);
nor UO_1922 (O_1922,N_20395,N_21445);
and UO_1923 (O_1923,N_24383,N_19875);
xnor UO_1924 (O_1924,N_24398,N_23160);
nor UO_1925 (O_1925,N_19092,N_21369);
nor UO_1926 (O_1926,N_22390,N_24814);
or UO_1927 (O_1927,N_21788,N_21226);
nand UO_1928 (O_1928,N_18818,N_19105);
and UO_1929 (O_1929,N_22941,N_21772);
nand UO_1930 (O_1930,N_23994,N_22616);
nand UO_1931 (O_1931,N_20131,N_19399);
nand UO_1932 (O_1932,N_23859,N_21657);
xnor UO_1933 (O_1933,N_24139,N_18938);
xor UO_1934 (O_1934,N_22206,N_20931);
and UO_1935 (O_1935,N_20196,N_24216);
nor UO_1936 (O_1936,N_22948,N_22622);
or UO_1937 (O_1937,N_22604,N_20943);
and UO_1938 (O_1938,N_24520,N_19929);
xor UO_1939 (O_1939,N_23021,N_23456);
xnor UO_1940 (O_1940,N_22388,N_23887);
nand UO_1941 (O_1941,N_22039,N_19290);
xnor UO_1942 (O_1942,N_23245,N_20052);
nand UO_1943 (O_1943,N_22589,N_19488);
and UO_1944 (O_1944,N_24888,N_21024);
xor UO_1945 (O_1945,N_20076,N_22666);
nor UO_1946 (O_1946,N_19675,N_22005);
or UO_1947 (O_1947,N_24812,N_20529);
nor UO_1948 (O_1948,N_24225,N_24763);
or UO_1949 (O_1949,N_19148,N_22571);
or UO_1950 (O_1950,N_22000,N_23891);
or UO_1951 (O_1951,N_24508,N_20176);
xnor UO_1952 (O_1952,N_23897,N_21867);
and UO_1953 (O_1953,N_21866,N_21450);
or UO_1954 (O_1954,N_22801,N_18954);
xor UO_1955 (O_1955,N_21879,N_24397);
nor UO_1956 (O_1956,N_20023,N_19404);
and UO_1957 (O_1957,N_20215,N_21133);
nor UO_1958 (O_1958,N_22488,N_22138);
and UO_1959 (O_1959,N_23081,N_21276);
xnor UO_1960 (O_1960,N_24626,N_24502);
or UO_1961 (O_1961,N_21146,N_23079);
or UO_1962 (O_1962,N_21954,N_23190);
nand UO_1963 (O_1963,N_23044,N_18970);
nand UO_1964 (O_1964,N_21752,N_23285);
xnor UO_1965 (O_1965,N_19858,N_22088);
nor UO_1966 (O_1966,N_21652,N_20624);
nor UO_1967 (O_1967,N_19977,N_21365);
nor UO_1968 (O_1968,N_22467,N_20340);
or UO_1969 (O_1969,N_23006,N_20283);
nor UO_1970 (O_1970,N_21419,N_18929);
nor UO_1971 (O_1971,N_18753,N_23225);
or UO_1972 (O_1972,N_21527,N_24525);
nand UO_1973 (O_1973,N_23178,N_24678);
or UO_1974 (O_1974,N_21421,N_21913);
or UO_1975 (O_1975,N_23196,N_23404);
nor UO_1976 (O_1976,N_23883,N_21885);
or UO_1977 (O_1977,N_22376,N_24156);
or UO_1978 (O_1978,N_21961,N_21723);
or UO_1979 (O_1979,N_23437,N_19407);
nand UO_1980 (O_1980,N_24476,N_23287);
nand UO_1981 (O_1981,N_21994,N_18851);
and UO_1982 (O_1982,N_24329,N_21022);
xor UO_1983 (O_1983,N_21340,N_20518);
and UO_1984 (O_1984,N_19033,N_20620);
xnor UO_1985 (O_1985,N_20147,N_22625);
xor UO_1986 (O_1986,N_20551,N_19255);
and UO_1987 (O_1987,N_19187,N_18992);
and UO_1988 (O_1988,N_24250,N_21839);
nor UO_1989 (O_1989,N_19508,N_22092);
and UO_1990 (O_1990,N_21172,N_21645);
or UO_1991 (O_1991,N_22690,N_19688);
and UO_1992 (O_1992,N_20418,N_20550);
xnor UO_1993 (O_1993,N_20879,N_19758);
or UO_1994 (O_1994,N_23410,N_22845);
nor UO_1995 (O_1995,N_21090,N_18828);
or UO_1996 (O_1996,N_18981,N_20708);
and UO_1997 (O_1997,N_23923,N_20399);
or UO_1998 (O_1998,N_22680,N_23468);
nand UO_1999 (O_1999,N_22952,N_22182);
nand UO_2000 (O_2000,N_22337,N_20199);
and UO_2001 (O_2001,N_21865,N_20493);
xnor UO_2002 (O_2002,N_22909,N_19117);
xor UO_2003 (O_2003,N_19422,N_24456);
nor UO_2004 (O_2004,N_22735,N_20647);
and UO_2005 (O_2005,N_22192,N_21088);
nand UO_2006 (O_2006,N_19902,N_21404);
or UO_2007 (O_2007,N_24864,N_19589);
or UO_2008 (O_2008,N_19420,N_20576);
and UO_2009 (O_2009,N_22556,N_23924);
or UO_2010 (O_2010,N_21009,N_20314);
and UO_2011 (O_2011,N_21923,N_20762);
or UO_2012 (O_2012,N_21733,N_23109);
xor UO_2013 (O_2013,N_19491,N_19923);
xor UO_2014 (O_2014,N_21033,N_23495);
xor UO_2015 (O_2015,N_21308,N_22967);
xor UO_2016 (O_2016,N_18873,N_24514);
nor UO_2017 (O_2017,N_22242,N_20754);
xor UO_2018 (O_2018,N_24202,N_19339);
and UO_2019 (O_2019,N_24380,N_21301);
and UO_2020 (O_2020,N_22786,N_24003);
nand UO_2021 (O_2021,N_19192,N_19591);
xor UO_2022 (O_2022,N_24701,N_19750);
nand UO_2023 (O_2023,N_20820,N_20304);
and UO_2024 (O_2024,N_20855,N_20436);
or UO_2025 (O_2025,N_24320,N_21610);
xnor UO_2026 (O_2026,N_21368,N_19581);
nand UO_2027 (O_2027,N_19484,N_19908);
nand UO_2028 (O_2028,N_19755,N_21311);
nor UO_2029 (O_2029,N_19204,N_21783);
nand UO_2030 (O_2030,N_23302,N_23651);
and UO_2031 (O_2031,N_22968,N_19502);
and UO_2032 (O_2032,N_23494,N_24064);
nand UO_2033 (O_2033,N_19707,N_18939);
or UO_2034 (O_2034,N_19909,N_21979);
or UO_2035 (O_2035,N_23780,N_23082);
nor UO_2036 (O_2036,N_22982,N_22567);
xnor UO_2037 (O_2037,N_23502,N_24421);
nand UO_2038 (O_2038,N_24468,N_23200);
and UO_2039 (O_2039,N_23552,N_23816);
or UO_2040 (O_2040,N_19716,N_23946);
nor UO_2041 (O_2041,N_19575,N_23317);
nand UO_2042 (O_2042,N_23609,N_20028);
nand UO_2043 (O_2043,N_23277,N_22075);
xor UO_2044 (O_2044,N_21878,N_19256);
nand UO_2045 (O_2045,N_22936,N_24897);
nand UO_2046 (O_2046,N_23395,N_23100);
nor UO_2047 (O_2047,N_19878,N_19163);
or UO_2048 (O_2048,N_18799,N_24167);
or UO_2049 (O_2049,N_24847,N_21519);
and UO_2050 (O_2050,N_23623,N_20735);
nand UO_2051 (O_2051,N_21064,N_21644);
or UO_2052 (O_2052,N_22608,N_20424);
and UO_2053 (O_2053,N_22687,N_22873);
xnor UO_2054 (O_2054,N_22969,N_24908);
nand UO_2055 (O_2055,N_21417,N_20881);
nand UO_2056 (O_2056,N_19280,N_21505);
nand UO_2057 (O_2057,N_24914,N_22840);
and UO_2058 (O_2058,N_18805,N_22685);
or UO_2059 (O_2059,N_24986,N_21988);
or UO_2060 (O_2060,N_19390,N_19332);
nor UO_2061 (O_2061,N_24751,N_20761);
and UO_2062 (O_2062,N_21225,N_24141);
and UO_2063 (O_2063,N_21297,N_18902);
or UO_2064 (O_2064,N_20609,N_21596);
or UO_2065 (O_2065,N_22416,N_24148);
xnor UO_2066 (O_2066,N_24029,N_23394);
nor UO_2067 (O_2067,N_21237,N_22347);
nor UO_2068 (O_2068,N_19474,N_24704);
nor UO_2069 (O_2069,N_18763,N_19704);
nor UO_2070 (O_2070,N_24128,N_24449);
nor UO_2071 (O_2071,N_20152,N_22375);
nor UO_2072 (O_2072,N_22844,N_22747);
nor UO_2073 (O_2073,N_20650,N_21491);
and UO_2074 (O_2074,N_23236,N_19013);
and UO_2075 (O_2075,N_24567,N_23499);
nor UO_2076 (O_2076,N_23955,N_24838);
nor UO_2077 (O_2077,N_19264,N_23982);
nand UO_2078 (O_2078,N_22672,N_24150);
or UO_2079 (O_2079,N_21518,N_21835);
nand UO_2080 (O_2080,N_22984,N_23185);
xor UO_2081 (O_2081,N_23485,N_20865);
nor UO_2082 (O_2082,N_23384,N_23271);
or UO_2083 (O_2083,N_20123,N_24638);
nor UO_2084 (O_2084,N_22349,N_24284);
nor UO_2085 (O_2085,N_24717,N_21838);
nand UO_2086 (O_2086,N_21556,N_20777);
or UO_2087 (O_2087,N_23921,N_19154);
nor UO_2088 (O_2088,N_22988,N_22290);
or UO_2089 (O_2089,N_21760,N_23933);
and UO_2090 (O_2090,N_23222,N_21458);
xnor UO_2091 (O_2091,N_23115,N_21203);
nand UO_2092 (O_2092,N_22373,N_18809);
nor UO_2093 (O_2093,N_24711,N_21960);
xnor UO_2094 (O_2094,N_21699,N_19585);
or UO_2095 (O_2095,N_19417,N_22471);
or UO_2096 (O_2096,N_24612,N_21345);
nand UO_2097 (O_2097,N_24713,N_22926);
nor UO_2098 (O_2098,N_20823,N_22836);
nor UO_2099 (O_2099,N_23477,N_21370);
nor UO_2100 (O_2100,N_22675,N_23097);
and UO_2101 (O_2101,N_20005,N_20292);
or UO_2102 (O_2102,N_22548,N_19790);
or UO_2103 (O_2103,N_21787,N_18777);
xnor UO_2104 (O_2104,N_18771,N_20552);
or UO_2105 (O_2105,N_21006,N_23219);
nand UO_2106 (O_2106,N_24122,N_24551);
xor UO_2107 (O_2107,N_20072,N_23576);
nand UO_2108 (O_2108,N_24766,N_20596);
nor UO_2109 (O_2109,N_21180,N_24513);
xor UO_2110 (O_2110,N_23320,N_23976);
nor UO_2111 (O_2111,N_24016,N_22239);
xor UO_2112 (O_2112,N_21289,N_19446);
or UO_2113 (O_2113,N_21668,N_24745);
nor UO_2114 (O_2114,N_22314,N_19826);
or UO_2115 (O_2115,N_24209,N_22009);
xor UO_2116 (O_2116,N_23543,N_23313);
nand UO_2117 (O_2117,N_23681,N_19056);
nand UO_2118 (O_2118,N_19289,N_20466);
and UO_2119 (O_2119,N_23419,N_18924);
xnor UO_2120 (O_2120,N_20618,N_22246);
nand UO_2121 (O_2121,N_22289,N_23345);
and UO_2122 (O_2122,N_19721,N_21831);
or UO_2123 (O_2123,N_21852,N_24097);
and UO_2124 (O_2124,N_20690,N_20481);
nor UO_2125 (O_2125,N_22859,N_18949);
nand UO_2126 (O_2126,N_23047,N_22443);
xnor UO_2127 (O_2127,N_24060,N_20295);
nor UO_2128 (O_2128,N_20795,N_19435);
nand UO_2129 (O_2129,N_21338,N_19434);
xnor UO_2130 (O_2130,N_20454,N_23820);
and UO_2131 (O_2131,N_22595,N_19825);
or UO_2132 (O_2132,N_22144,N_24285);
or UO_2133 (O_2133,N_21456,N_19472);
nor UO_2134 (O_2134,N_21744,N_19542);
nand UO_2135 (O_2135,N_23875,N_24147);
xnor UO_2136 (O_2136,N_23545,N_21349);
xor UO_2137 (O_2137,N_21170,N_19002);
nand UO_2138 (O_2138,N_24369,N_21648);
or UO_2139 (O_2139,N_24382,N_20657);
and UO_2140 (O_2140,N_19393,N_19677);
xor UO_2141 (O_2141,N_23937,N_21443);
xor UO_2142 (O_2142,N_22880,N_21312);
and UO_2143 (O_2143,N_20646,N_20319);
nand UO_2144 (O_2144,N_20623,N_20133);
or UO_2145 (O_2145,N_22003,N_21300);
and UO_2146 (O_2146,N_22204,N_21216);
nand UO_2147 (O_2147,N_24092,N_23785);
and UO_2148 (O_2148,N_23050,N_20321);
nor UO_2149 (O_2149,N_24631,N_19058);
nand UO_2150 (O_2150,N_24110,N_23687);
and UO_2151 (O_2151,N_23983,N_18943);
or UO_2152 (O_2152,N_23800,N_24673);
or UO_2153 (O_2153,N_18757,N_21303);
xor UO_2154 (O_2154,N_23342,N_21957);
xnor UO_2155 (O_2155,N_18872,N_18768);
xor UO_2156 (O_2156,N_24154,N_23099);
or UO_2157 (O_2157,N_19135,N_24098);
nor UO_2158 (O_2158,N_19355,N_21245);
nor UO_2159 (O_2159,N_20286,N_21219);
xor UO_2160 (O_2160,N_24460,N_21086);
nor UO_2161 (O_2161,N_19106,N_24046);
xnor UO_2162 (O_2162,N_19141,N_19195);
nor UO_2163 (O_2163,N_18886,N_22752);
xnor UO_2164 (O_2164,N_20159,N_22137);
or UO_2165 (O_2165,N_19851,N_21642);
nand UO_2166 (O_2166,N_19427,N_21643);
nand UO_2167 (O_2167,N_22056,N_21227);
and UO_2168 (O_2168,N_24911,N_22491);
nor UO_2169 (O_2169,N_21741,N_24999);
or UO_2170 (O_2170,N_21118,N_24268);
or UO_2171 (O_2171,N_20675,N_24759);
nand UO_2172 (O_2172,N_23550,N_21558);
or UO_2173 (O_2173,N_21013,N_22097);
nor UO_2174 (O_2174,N_19586,N_21580);
nor UO_2175 (O_2175,N_24244,N_22765);
and UO_2176 (O_2176,N_19383,N_21183);
or UO_2177 (O_2177,N_18907,N_19317);
and UO_2178 (O_2178,N_24391,N_24479);
and UO_2179 (O_2179,N_21154,N_19131);
or UO_2180 (O_2180,N_23745,N_19770);
or UO_2181 (O_2181,N_22224,N_23476);
and UO_2182 (O_2182,N_21335,N_23015);
and UO_2183 (O_2183,N_19129,N_24565);
or UO_2184 (O_2184,N_22118,N_19906);
and UO_2185 (O_2185,N_22764,N_24354);
nand UO_2186 (O_2186,N_22999,N_20191);
or UO_2187 (O_2187,N_21828,N_20911);
or UO_2188 (O_2188,N_24796,N_24149);
nand UO_2189 (O_2189,N_24890,N_19085);
xor UO_2190 (O_2190,N_24076,N_23244);
or UO_2191 (O_2191,N_21819,N_20819);
nor UO_2192 (O_2192,N_20811,N_21698);
nand UO_2193 (O_2193,N_24853,N_20193);
and UO_2194 (O_2194,N_23153,N_21005);
nor UO_2195 (O_2195,N_24960,N_19660);
nor UO_2196 (O_2196,N_23303,N_24666);
and UO_2197 (O_2197,N_19436,N_24576);
nand UO_2198 (O_2198,N_22663,N_22063);
and UO_2199 (O_2199,N_20840,N_19400);
xnor UO_2200 (O_2200,N_19177,N_18852);
or UO_2201 (O_2201,N_23603,N_21750);
or UO_2202 (O_2202,N_18998,N_22334);
nand UO_2203 (O_2203,N_24388,N_22249);
and UO_2204 (O_2204,N_20098,N_20068);
or UO_2205 (O_2205,N_22541,N_20307);
and UO_2206 (O_2206,N_20726,N_24039);
nor UO_2207 (O_2207,N_22252,N_24510);
xor UO_2208 (O_2208,N_22303,N_22483);
nor UO_2209 (O_2209,N_24722,N_23355);
nor UO_2210 (O_2210,N_20612,N_23399);
nor UO_2211 (O_2211,N_19994,N_24981);
and UO_2212 (O_2212,N_24957,N_20059);
nand UO_2213 (O_2213,N_22986,N_19037);
or UO_2214 (O_2214,N_23926,N_24170);
or UO_2215 (O_2215,N_20413,N_18801);
or UO_2216 (O_2216,N_24834,N_23339);
or UO_2217 (O_2217,N_18817,N_20588);
or UO_2218 (O_2218,N_21077,N_22220);
and UO_2219 (O_2219,N_20001,N_23135);
or UO_2220 (O_2220,N_21849,N_23929);
nor UO_2221 (O_2221,N_22879,N_23415);
and UO_2222 (O_2222,N_18966,N_21093);
nand UO_2223 (O_2223,N_19379,N_20684);
nand UO_2224 (O_2224,N_21920,N_23232);
xnor UO_2225 (O_2225,N_20078,N_22987);
or UO_2226 (O_2226,N_20081,N_20932);
xnor UO_2227 (O_2227,N_21287,N_24769);
and UO_2228 (O_2228,N_23165,N_22265);
nand UO_2229 (O_2229,N_21706,N_21489);
xnor UO_2230 (O_2230,N_24486,N_21247);
and UO_2231 (O_2231,N_23658,N_21017);
nand UO_2232 (O_2232,N_23755,N_21341);
nand UO_2233 (O_2233,N_20919,N_20087);
nor UO_2234 (O_2234,N_19185,N_21731);
and UO_2235 (O_2235,N_19879,N_23754);
xnor UO_2236 (O_2236,N_23133,N_24884);
and UO_2237 (O_2237,N_23466,N_22858);
nor UO_2238 (O_2238,N_22751,N_22596);
and UO_2239 (O_2239,N_19282,N_22558);
or UO_2240 (O_2240,N_21080,N_19416);
xnor UO_2241 (O_2241,N_21775,N_22912);
xnor UO_2242 (O_2242,N_20422,N_23336);
nor UO_2243 (O_2243,N_21191,N_21395);
nand UO_2244 (O_2244,N_20717,N_24414);
nor UO_2245 (O_2245,N_23827,N_23321);
nor UO_2246 (O_2246,N_24333,N_19895);
and UO_2247 (O_2247,N_22807,N_19369);
xnor UO_2248 (O_2248,N_23013,N_22029);
xnor UO_2249 (O_2249,N_21460,N_21438);
nand UO_2250 (O_2250,N_22550,N_23861);
nand UO_2251 (O_2251,N_23598,N_19201);
nor UO_2252 (O_2252,N_21025,N_21631);
and UO_2253 (O_2253,N_20920,N_20826);
nor UO_2254 (O_2254,N_22199,N_23101);
or UO_2255 (O_2255,N_19431,N_23435);
xnor UO_2256 (O_2256,N_23586,N_23788);
xor UO_2257 (O_2257,N_24873,N_22257);
xnor UO_2258 (O_2258,N_22711,N_22644);
xnor UO_2259 (O_2259,N_21918,N_20649);
or UO_2260 (O_2260,N_21120,N_21871);
and UO_2261 (O_2261,N_21337,N_24676);
and UO_2262 (O_2262,N_23782,N_20121);
nand UO_2263 (O_2263,N_23764,N_20387);
nand UO_2264 (O_2264,N_23746,N_21390);
or UO_2265 (O_2265,N_20440,N_22656);
or UO_2266 (O_2266,N_24237,N_23826);
xor UO_2267 (O_2267,N_22757,N_24127);
nand UO_2268 (O_2268,N_20594,N_21030);
nor UO_2269 (O_2269,N_21840,N_23118);
and UO_2270 (O_2270,N_23475,N_23128);
nand UO_2271 (O_2271,N_21116,N_21134);
nor UO_2272 (O_2272,N_19311,N_23698);
or UO_2273 (O_2273,N_19732,N_24533);
nor UO_2274 (O_2274,N_18878,N_22374);
or UO_2275 (O_2275,N_20487,N_20430);
nand UO_2276 (O_2276,N_23717,N_22703);
xnor UO_2277 (O_2277,N_23987,N_24422);
nor UO_2278 (O_2278,N_19070,N_20700);
xor UO_2279 (O_2279,N_20501,N_21617);
and UO_2280 (O_2280,N_18955,N_21507);
and UO_2281 (O_2281,N_20301,N_23580);
or UO_2282 (O_2282,N_19523,N_22203);
and UO_2283 (O_2283,N_24659,N_20491);
nand UO_2284 (O_2284,N_21196,N_24870);
or UO_2285 (O_2285,N_19225,N_20940);
xor UO_2286 (O_2286,N_20543,N_18794);
xnor UO_2287 (O_2287,N_20394,N_19643);
nand UO_2288 (O_2288,N_24430,N_21194);
nor UO_2289 (O_2289,N_20858,N_18905);
nor UO_2290 (O_2290,N_19768,N_18996);
nand UO_2291 (O_2291,N_24262,N_18923);
nand UO_2292 (O_2292,N_21076,N_22892);
nand UO_2293 (O_2293,N_22272,N_24186);
xor UO_2294 (O_2294,N_21477,N_20135);
or UO_2295 (O_2295,N_21701,N_20216);
xor UO_2296 (O_2296,N_23536,N_22210);
and UO_2297 (O_2297,N_20227,N_21620);
nand UO_2298 (O_2298,N_21178,N_20198);
xnor UO_2299 (O_2299,N_19883,N_24464);
and UO_2300 (O_2300,N_24506,N_19818);
xor UO_2301 (O_2301,N_22484,N_19246);
nand UO_2302 (O_2302,N_24037,N_23096);
or UO_2303 (O_2303,N_20266,N_22922);
nand UO_2304 (O_2304,N_20908,N_19637);
nor UO_2305 (O_2305,N_21929,N_21531);
and UO_2306 (O_2306,N_18936,N_20467);
or UO_2307 (O_2307,N_23954,N_19316);
nand UO_2308 (O_2308,N_20863,N_23080);
and UO_2309 (O_2309,N_21904,N_19639);
xor UO_2310 (O_2310,N_22827,N_19725);
nor UO_2311 (O_2311,N_24580,N_21392);
xor UO_2312 (O_2312,N_22749,N_20921);
nor UO_2313 (O_2313,N_24185,N_24851);
nor UO_2314 (O_2314,N_19079,N_18874);
or UO_2315 (O_2315,N_21026,N_22629);
and UO_2316 (O_2316,N_23661,N_23311);
and UO_2317 (O_2317,N_22613,N_20405);
nor UO_2318 (O_2318,N_21825,N_24560);
and UO_2319 (O_2319,N_19576,N_18755);
nor UO_2320 (O_2320,N_24811,N_21484);
or UO_2321 (O_2321,N_22026,N_24541);
or UO_2322 (O_2322,N_20389,N_19476);
or UO_2323 (O_2323,N_23112,N_18881);
nor UO_2324 (O_2324,N_20003,N_21034);
nor UO_2325 (O_2325,N_21684,N_23179);
nand UO_2326 (O_2326,N_24574,N_21377);
and UO_2327 (O_2327,N_22630,N_24277);
or UO_2328 (O_2328,N_21202,N_24861);
and UO_2329 (O_2329,N_19211,N_18883);
nand UO_2330 (O_2330,N_22420,N_24532);
nor UO_2331 (O_2331,N_21748,N_24963);
nand UO_2332 (O_2332,N_20722,N_19206);
nor UO_2333 (O_2333,N_19146,N_18859);
or UO_2334 (O_2334,N_19847,N_21042);
and UO_2335 (O_2335,N_20573,N_19599);
and UO_2336 (O_2336,N_23496,N_21992);
xor UO_2337 (O_2337,N_24668,N_21441);
nand UO_2338 (O_2338,N_22212,N_20201);
nor UO_2339 (O_2339,N_19263,N_19341);
or UO_2340 (O_2340,N_21955,N_24232);
and UO_2341 (O_2341,N_21562,N_24825);
xor UO_2342 (O_2342,N_22784,N_19698);
or UO_2343 (O_2343,N_22345,N_24228);
and UO_2344 (O_2344,N_20640,N_22111);
and UO_2345 (O_2345,N_24172,N_22024);
nand UO_2346 (O_2346,N_20752,N_19672);
or UO_2347 (O_2347,N_18920,N_22207);
nor UO_2348 (O_2348,N_19175,N_23448);
nor UO_2349 (O_2349,N_21286,N_23667);
xor UO_2350 (O_2350,N_24880,N_23332);
nand UO_2351 (O_2351,N_22132,N_19942);
nor UO_2352 (O_2352,N_23105,N_23996);
nand UO_2353 (O_2353,N_21429,N_20184);
xnor UO_2354 (O_2354,N_19605,N_21758);
xnor UO_2355 (O_2355,N_23090,N_23093);
and UO_2356 (O_2356,N_22017,N_22415);
xor UO_2357 (O_2357,N_19223,N_22038);
xor UO_2358 (O_2358,N_20710,N_22848);
or UO_2359 (O_2359,N_20411,N_24242);
xnor UO_2360 (O_2360,N_22047,N_18795);
nor UO_2361 (O_2361,N_20682,N_19075);
and UO_2362 (O_2362,N_20167,N_24518);
or UO_2363 (O_2363,N_19061,N_23977);
nand UO_2364 (O_2364,N_20160,N_20185);
nor UO_2365 (O_2365,N_21469,N_20379);
and UO_2366 (O_2366,N_23471,N_20970);
nor UO_2367 (O_2367,N_23061,N_24549);
or UO_2368 (O_2368,N_23215,N_20732);
nand UO_2369 (O_2369,N_19548,N_20402);
xnor UO_2370 (O_2370,N_19762,N_21690);
xnor UO_2371 (O_2371,N_19069,N_23888);
or UO_2372 (O_2372,N_22123,N_22900);
xnor UO_2373 (O_2373,N_18826,N_18764);
nand UO_2374 (O_2374,N_24028,N_20547);
nor UO_2375 (O_2375,N_20154,N_23733);
xor UO_2376 (O_2376,N_23989,N_20632);
nor UO_2377 (O_2377,N_23354,N_19244);
nand UO_2378 (O_2378,N_22561,N_21535);
xnor UO_2379 (O_2379,N_22300,N_23470);
or UO_2380 (O_2380,N_19053,N_20450);
xnor UO_2381 (O_2381,N_20827,N_23822);
or UO_2382 (O_2382,N_21534,N_19618);
nand UO_2383 (O_2383,N_24168,N_20572);
nor UO_2384 (O_2384,N_24750,N_20753);
nand UO_2385 (O_2385,N_20586,N_22837);
nand UO_2386 (O_2386,N_19714,N_19359);
xor UO_2387 (O_2387,N_23595,N_24534);
and UO_2388 (O_2388,N_24116,N_24600);
nand UO_2389 (O_2389,N_21075,N_19327);
nand UO_2390 (O_2390,N_21420,N_20787);
xnor UO_2391 (O_2391,N_24337,N_24086);
and UO_2392 (O_2392,N_19351,N_21647);
nand UO_2393 (O_2393,N_22427,N_19324);
nor UO_2394 (O_2394,N_19490,N_18750);
and UO_2395 (O_2395,N_23652,N_22852);
nor UO_2396 (O_2396,N_22679,N_21615);
nand UO_2397 (O_2397,N_24718,N_24470);
xnor UO_2398 (O_2398,N_21693,N_22733);
or UO_2399 (O_2399,N_23314,N_22626);
nor UO_2400 (O_2400,N_20337,N_20145);
and UO_2401 (O_2401,N_19582,N_23669);
nand UO_2402 (O_2402,N_22930,N_23676);
nand UO_2403 (O_2403,N_18803,N_22317);
nor UO_2404 (O_2404,N_23507,N_21496);
or UO_2405 (O_2405,N_19125,N_22341);
nand UO_2406 (O_2406,N_19152,N_23438);
or UO_2407 (O_2407,N_20615,N_22044);
and UO_2408 (O_2408,N_24081,N_23784);
xor UO_2409 (O_2409,N_19303,N_20780);
nand UO_2410 (O_2410,N_22820,N_24072);
or UO_2411 (O_2411,N_21941,N_24437);
and UO_2412 (O_2412,N_19881,N_21028);
nand UO_2413 (O_2413,N_19514,N_23690);
nand UO_2414 (O_2414,N_22380,N_18950);
nor UO_2415 (O_2415,N_23014,N_20656);
xnor UO_2416 (O_2416,N_22028,N_23195);
nor UO_2417 (O_2417,N_21627,N_21847);
nand UO_2418 (O_2418,N_22391,N_22175);
and UO_2419 (O_2419,N_19916,N_20527);
nand UO_2420 (O_2420,N_24916,N_19367);
or UO_2421 (O_2421,N_21366,N_22323);
and UO_2422 (O_2422,N_22492,N_24927);
nand UO_2423 (O_2423,N_21455,N_20778);
xnor UO_2424 (O_2424,N_24550,N_23759);
or UO_2425 (O_2425,N_23382,N_19961);
nand UO_2426 (O_2426,N_20740,N_24789);
nand UO_2427 (O_2427,N_21218,N_19189);
or UO_2428 (O_2428,N_19276,N_23260);
and UO_2429 (O_2429,N_22668,N_22609);
or UO_2430 (O_2430,N_24553,N_19180);
nor UO_2431 (O_2431,N_22229,N_20328);
nand UO_2432 (O_2432,N_24078,N_19999);
xnor UO_2433 (O_2433,N_23879,N_20153);
or UO_2434 (O_2434,N_19799,N_23948);
nand UO_2435 (O_2435,N_23370,N_23972);
xor UO_2436 (O_2436,N_22160,N_23036);
xnor UO_2437 (O_2437,N_19958,N_19247);
xor UO_2438 (O_2438,N_24670,N_23514);
and UO_2439 (O_2439,N_19741,N_20331);
or UO_2440 (O_2440,N_21049,N_19624);
nand UO_2441 (O_2441,N_19703,N_24995);
nand UO_2442 (O_2442,N_21536,N_24746);
or UO_2443 (O_2443,N_24781,N_22072);
xor UO_2444 (O_2444,N_22164,N_21557);
and UO_2445 (O_2445,N_23458,N_24138);
and UO_2446 (O_2446,N_23570,N_23538);
and UO_2447 (O_2447,N_24926,N_20476);
nor UO_2448 (O_2448,N_20366,N_24503);
or UO_2449 (O_2449,N_22864,N_21874);
nor UO_2450 (O_2450,N_23088,N_23647);
nand UO_2451 (O_2451,N_21651,N_23282);
and UO_2452 (O_2452,N_20107,N_19823);
or UO_2453 (O_2453,N_24819,N_23368);
or UO_2454 (O_2454,N_24155,N_20049);
nand UO_2455 (O_2455,N_23335,N_21471);
and UO_2456 (O_2456,N_22027,N_24048);
and UO_2457 (O_2457,N_24720,N_23584);
and UO_2458 (O_2458,N_23056,N_24929);
nor UO_2459 (O_2459,N_22081,N_23657);
nand UO_2460 (O_2460,N_18897,N_21503);
xor UO_2461 (O_2461,N_20803,N_21382);
or UO_2462 (O_2462,N_20018,N_20954);
nand UO_2463 (O_2463,N_24199,N_20410);
xnor UO_2464 (O_2464,N_23919,N_21128);
nor UO_2465 (O_2465,N_19573,N_22544);
nor UO_2466 (O_2466,N_21165,N_21930);
or UO_2467 (O_2467,N_21002,N_19553);
nand UO_2468 (O_2468,N_24544,N_24190);
or UO_2469 (O_2469,N_18758,N_20097);
or UO_2470 (O_2470,N_23201,N_23725);
xor UO_2471 (O_2471,N_24681,N_21197);
and UO_2472 (O_2472,N_19593,N_24883);
nand UO_2473 (O_2473,N_23457,N_19165);
and UO_2474 (O_2474,N_24739,N_21355);
and UO_2475 (O_2475,N_22142,N_19291);
xnor UO_2476 (O_2476,N_19571,N_24481);
xnor UO_2477 (O_2477,N_24137,N_23031);
nand UO_2478 (O_2478,N_21348,N_21608);
and UO_2479 (O_2479,N_20672,N_22768);
nor UO_2480 (O_2480,N_21299,N_23235);
and UO_2481 (O_2481,N_21332,N_19941);
nand UO_2482 (O_2482,N_21205,N_20230);
or UO_2483 (O_2483,N_24546,N_21250);
xnor UO_2484 (O_2484,N_22842,N_22371);
and UO_2485 (O_2485,N_22409,N_20141);
xor UO_2486 (O_2486,N_23721,N_20991);
nand UO_2487 (O_2487,N_24893,N_21833);
nor UO_2488 (O_2488,N_22707,N_22489);
xnor UO_2489 (O_2489,N_22234,N_21797);
xnor UO_2490 (O_2490,N_24835,N_24305);
nor UO_2491 (O_2491,N_20742,N_19405);
nor UO_2492 (O_2492,N_20472,N_24052);
xor UO_2493 (O_2493,N_19091,N_24121);
and UO_2494 (O_2494,N_23720,N_21563);
nor UO_2495 (O_2495,N_23439,N_19448);
nand UO_2496 (O_2496,N_22299,N_21582);
xnor UO_2497 (O_2497,N_21827,N_20388);
xor UO_2498 (O_2498,N_19985,N_21141);
or UO_2499 (O_2499,N_22554,N_21258);
nand UO_2500 (O_2500,N_23620,N_20051);
xor UO_2501 (O_2501,N_23627,N_19896);
xor UO_2502 (O_2502,N_21623,N_24778);
nand UO_2503 (O_2503,N_23903,N_19915);
or UO_2504 (O_2504,N_20824,N_21152);
nand UO_2505 (O_2505,N_20300,N_24987);
xnor UO_2506 (O_2506,N_19563,N_23137);
xnor UO_2507 (O_2507,N_22714,N_19901);
xnor UO_2508 (O_2508,N_21320,N_22051);
nand UO_2509 (O_2509,N_19530,N_20428);
nor UO_2510 (O_2510,N_24625,N_24737);
xor UO_2511 (O_2511,N_24089,N_18958);
or UO_2512 (O_2512,N_21747,N_21040);
xnor UO_2513 (O_2513,N_21336,N_22258);
nor UO_2514 (O_2514,N_20915,N_19760);
nand UO_2515 (O_2515,N_23273,N_20733);
nand UO_2516 (O_2516,N_20982,N_22441);
nor UO_2517 (O_2517,N_19183,N_21294);
nand UO_2518 (O_2518,N_24364,N_22950);
xnor UO_2519 (O_2519,N_24314,N_21436);
nand UO_2520 (O_2520,N_24815,N_19904);
or UO_2521 (O_2521,N_18916,N_21306);
or UO_2522 (O_2522,N_19361,N_24931);
xor UO_2523 (O_2523,N_19433,N_22243);
and UO_2524 (O_2524,N_20060,N_23779);
nor UO_2525 (O_2525,N_24654,N_24849);
or UO_2526 (O_2526,N_23659,N_22168);
nor UO_2527 (O_2527,N_23583,N_23588);
and UO_2528 (O_2528,N_19396,N_20537);
nor UO_2529 (O_2529,N_19655,N_23522);
or UO_2530 (O_2530,N_23490,N_19816);
xor UO_2531 (O_2531,N_21987,N_20438);
nor UO_2532 (O_2532,N_23761,N_23839);
nand UO_2533 (O_2533,N_20767,N_24723);
nor UO_2534 (O_2534,N_24100,N_22301);
nor UO_2535 (O_2535,N_20378,N_21926);
and UO_2536 (O_2536,N_24248,N_19394);
or UO_2537 (O_2537,N_20425,N_24375);
or UO_2538 (O_2538,N_20429,N_20156);
or UO_2539 (O_2539,N_23464,N_19619);
nor UO_2540 (O_2540,N_21494,N_24144);
xor UO_2541 (O_2541,N_22817,N_24041);
nand UO_2542 (O_2542,N_19463,N_22077);
nand UO_2543 (O_2543,N_19031,N_22631);
nor UO_2544 (O_2544,N_21481,N_21618);
xor UO_2545 (O_2545,N_21249,N_20455);
or UO_2546 (O_2546,N_19469,N_23157);
nor UO_2547 (O_2547,N_20350,N_18913);
xnor UO_2548 (O_2548,N_19049,N_23762);
and UO_2549 (O_2549,N_23479,N_20562);
or UO_2550 (O_2550,N_20927,N_18980);
or UO_2551 (O_2551,N_21729,N_20985);
and UO_2552 (O_2552,N_22149,N_24776);
or UO_2553 (O_2553,N_23622,N_23019);
xnor UO_2554 (O_2554,N_23324,N_24325);
xor UO_2555 (O_2555,N_19029,N_24562);
xor UO_2556 (O_2556,N_24872,N_24540);
xnor UO_2557 (O_2557,N_21327,N_22871);
nor UO_2558 (O_2558,N_20013,N_19992);
or UO_2559 (O_2559,N_20923,N_21689);
nand UO_2560 (O_2560,N_22916,N_22062);
or UO_2561 (O_2561,N_19556,N_22106);
nor UO_2562 (O_2562,N_21483,N_19151);
nand UO_2563 (O_2563,N_20772,N_24577);
nor UO_2564 (O_2564,N_19544,N_21791);
or UO_2565 (O_2565,N_19098,N_22173);
nor UO_2566 (O_2566,N_23511,N_19252);
nor UO_2567 (O_2567,N_21720,N_20764);
or UO_2568 (O_2568,N_23958,N_20054);
nand UO_2569 (O_2569,N_19676,N_24205);
nor UO_2570 (O_2570,N_21572,N_21041);
or UO_2571 (O_2571,N_24974,N_19310);
and UO_2572 (O_2572,N_20146,N_23212);
or UO_2573 (O_2573,N_23316,N_20504);
and UO_2574 (O_2574,N_24738,N_19930);
and UO_2575 (O_2575,N_23836,N_20860);
xnor UO_2576 (O_2576,N_22767,N_20096);
and UO_2577 (O_2577,N_20748,N_24178);
or UO_2578 (O_2578,N_19217,N_22532);
and UO_2579 (O_2579,N_19911,N_19967);
or UO_2580 (O_2580,N_23231,N_19649);
and UO_2581 (O_2581,N_22569,N_20083);
xor UO_2582 (O_2582,N_24311,N_20024);
and UO_2583 (O_2583,N_24292,N_24433);
or UO_2584 (O_2584,N_20212,N_21637);
xnor UO_2585 (O_2585,N_19905,N_22342);
xnor UO_2586 (O_2586,N_24545,N_20274);
or UO_2587 (O_2587,N_21123,N_24857);
or UO_2588 (O_2588,N_19096,N_23293);
or UO_2589 (O_2589,N_19088,N_21932);
and UO_2590 (O_2590,N_23114,N_22115);
xor UO_2591 (O_2591,N_20173,N_20935);
nor UO_2592 (O_2592,N_24990,N_24300);
nand UO_2593 (O_2593,N_20085,N_20278);
and UO_2594 (O_2594,N_19693,N_23884);
nand UO_2595 (O_2595,N_23024,N_21354);
or UO_2596 (O_2596,N_21504,N_22326);
xnor UO_2597 (O_2597,N_20095,N_24043);
and UO_2598 (O_2598,N_19996,N_21241);
nor UO_2599 (O_2599,N_24504,N_20317);
and UO_2600 (O_2600,N_21451,N_20950);
and UO_2601 (O_2601,N_23445,N_21091);
or UO_2602 (O_2602,N_19751,N_20846);
xnor UO_2603 (O_2603,N_19567,N_23641);
nand UO_2604 (O_2604,N_20453,N_23798);
nor UO_2605 (O_2605,N_23069,N_19841);
xor UO_2606 (O_2606,N_20971,N_21526);
nor UO_2607 (O_2607,N_20393,N_23204);
and UO_2608 (O_2608,N_20065,N_21492);
nand UO_2609 (O_2609,N_24663,N_19580);
and UO_2610 (O_2610,N_21356,N_21672);
nand UO_2611 (O_2611,N_21440,N_19426);
and UO_2612 (O_2612,N_19536,N_23256);
nand UO_2613 (O_2613,N_21046,N_20000);
and UO_2614 (O_2614,N_24045,N_24761);
or UO_2615 (O_2615,N_19711,N_23741);
xnor UO_2616 (O_2616,N_21148,N_23298);
nand UO_2617 (O_2617,N_21680,N_22731);
nand UO_2618 (O_2618,N_21363,N_21818);
or UO_2619 (O_2619,N_24758,N_23905);
xnor UO_2620 (O_2620,N_21663,N_24197);
xor UO_2621 (O_2621,N_24287,N_21712);
or UO_2622 (O_2622,N_21934,N_22320);
or UO_2623 (O_2623,N_24069,N_22728);
xor UO_2624 (O_2624,N_24030,N_24656);
xnor UO_2625 (O_2625,N_23974,N_18978);
nand UO_2626 (O_2626,N_22777,N_19411);
and UO_2627 (O_2627,N_24294,N_23329);
nand UO_2628 (O_2628,N_23614,N_23465);
and UO_2629 (O_2629,N_19191,N_20583);
xor UO_2630 (O_2630,N_20058,N_22089);
xor UO_2631 (O_2631,N_21986,N_24964);
and UO_2632 (O_2632,N_24282,N_24023);
and UO_2633 (O_2633,N_20480,N_23007);
nor UO_2634 (O_2634,N_19572,N_22696);
nor UO_2635 (O_2635,N_22637,N_20849);
or UO_2636 (O_2636,N_22877,N_21550);
and UO_2637 (O_2637,N_22881,N_20150);
xnor UO_2638 (O_2638,N_19340,N_20162);
nand UO_2639 (O_2639,N_19322,N_19261);
xor UO_2640 (O_2640,N_22623,N_23593);
and UO_2641 (O_2641,N_20961,N_18987);
xor UO_2642 (O_2642,N_23600,N_21967);
nor UO_2643 (O_2643,N_22305,N_20240);
and UO_2644 (O_2644,N_20668,N_19025);
nand UO_2645 (O_2645,N_24621,N_23371);
nand UO_2646 (O_2646,N_22330,N_24221);
or UO_2647 (O_2647,N_21115,N_23393);
nor UO_2648 (O_2648,N_20688,N_23742);
nand UO_2649 (O_2649,N_22201,N_24707);
nand UO_2650 (O_2650,N_20363,N_19272);
xor UO_2651 (O_2651,N_20094,N_22736);
nand UO_2652 (O_2652,N_24721,N_21452);
or UO_2653 (O_2653,N_19500,N_21691);
nand UO_2654 (O_2654,N_22709,N_19627);
xnor UO_2655 (O_2655,N_22657,N_22669);
nor UO_2656 (O_2656,N_21959,N_20189);
nor UO_2657 (O_2657,N_19780,N_20263);
nand UO_2658 (O_2658,N_19388,N_24624);
or UO_2659 (O_2659,N_23803,N_21230);
xor UO_2660 (O_2660,N_19467,N_24441);
xor UO_2661 (O_2661,N_21129,N_23155);
and UO_2662 (O_2662,N_20336,N_19321);
and UO_2663 (O_2663,N_19803,N_20664);
nor UO_2664 (O_2664,N_23087,N_23039);
nor UO_2665 (O_2665,N_21714,N_20484);
nand UO_2666 (O_2666,N_24025,N_20835);
nand UO_2667 (O_2667,N_24887,N_23876);
xnor UO_2668 (O_2668,N_20112,N_23032);
nand UO_2669 (O_2669,N_18819,N_23838);
nand UO_2670 (O_2670,N_23691,N_18964);
xnor UO_2671 (O_2671,N_24901,N_23187);
nand UO_2672 (O_2672,N_19873,N_19968);
nor UO_2673 (O_2673,N_20893,N_18836);
and UO_2674 (O_2674,N_19408,N_18990);
xnor UO_2675 (O_2675,N_23555,N_20822);
and UO_2676 (O_2676,N_22989,N_21616);
and UO_2677 (O_2677,N_19863,N_24552);
nor UO_2678 (O_2678,N_18839,N_22069);
nand UO_2679 (O_2679,N_20866,N_24899);
and UO_2680 (O_2680,N_24099,N_24871);
and UO_2681 (O_2681,N_20181,N_19783);
nand UO_2682 (O_2682,N_23388,N_22739);
and UO_2683 (O_2683,N_20177,N_23312);
nand UO_2684 (O_2684,N_19350,N_22269);
nor UO_2685 (O_2685,N_24730,N_22660);
or UO_2686 (O_2686,N_23795,N_19558);
or UO_2687 (O_2687,N_20244,N_21697);
and UO_2688 (O_2688,N_19084,N_20962);
or UO_2689 (O_2689,N_19412,N_22287);
xnor UO_2690 (O_2690,N_19769,N_20272);
xor UO_2691 (O_2691,N_23960,N_21686);
and UO_2692 (O_2692,N_24373,N_22417);
xor UO_2693 (O_2693,N_23706,N_19481);
nand UO_2694 (O_2694,N_21512,N_20992);
or UO_2695 (O_2695,N_21721,N_22695);
and UO_2696 (O_2696,N_23594,N_19913);
nand UO_2697 (O_2697,N_22020,N_22507);
and UO_2698 (O_2698,N_23525,N_21296);
and UO_2699 (O_2699,N_24554,N_24055);
or UO_2700 (O_2700,N_20352,N_23046);
nand UO_2701 (O_2701,N_23240,N_19786);
xnor UO_2702 (O_2702,N_20259,N_19182);
nor UO_2703 (O_2703,N_19308,N_23491);
and UO_2704 (O_2704,N_21281,N_24613);
or UO_2705 (O_2705,N_20056,N_23674);
nor UO_2706 (O_2706,N_20903,N_24351);
or UO_2707 (O_2707,N_24618,N_18977);
and UO_2708 (O_2708,N_24773,N_24417);
nor UO_2709 (O_2709,N_22284,N_18931);
and UO_2710 (O_2710,N_23531,N_18919);
nor UO_2711 (O_2711,N_24429,N_21844);
or UO_2712 (O_2712,N_20837,N_19221);
nor UO_2713 (O_2713,N_23425,N_23911);
nor UO_2714 (O_2714,N_22359,N_22034);
xnor UO_2715 (O_2715,N_23276,N_20510);
nand UO_2716 (O_2716,N_23331,N_22386);
nor UO_2717 (O_2717,N_20432,N_22043);
and UO_2718 (O_2718,N_23736,N_23141);
and UO_2719 (O_2719,N_18766,N_23230);
xnor UO_2720 (O_2720,N_22835,N_22240);
nor UO_2721 (O_2721,N_19806,N_21121);
xor UO_2722 (O_2722,N_22497,N_18845);
and UO_2723 (O_2723,N_21801,N_23968);
or UO_2724 (O_2724,N_20514,N_21239);
nand UO_2725 (O_2725,N_20257,N_22031);
nor UO_2726 (O_2726,N_20305,N_22165);
and UO_2727 (O_2727,N_20633,N_23416);
xnor UO_2728 (O_2728,N_19492,N_19113);
or UO_2729 (O_2729,N_19039,N_24708);
or UO_2730 (O_2730,N_23189,N_19265);
xor UO_2731 (O_2731,N_23427,N_22826);
nor UO_2732 (O_2732,N_23489,N_24322);
and UO_2733 (O_2733,N_22756,N_22166);
and UO_2734 (O_2734,N_22174,N_24461);
or UO_2735 (O_2735,N_20953,N_22068);
xor UO_2736 (O_2736,N_20332,N_21675);
or UO_2737 (O_2737,N_21124,N_22298);
nand UO_2738 (O_2738,N_24928,N_23442);
xnor UO_2739 (O_2739,N_20779,N_20282);
nor UO_2740 (O_2740,N_24603,N_22274);
nand UO_2741 (O_2741,N_18824,N_24327);
and UO_2742 (O_2742,N_21061,N_21331);
nor UO_2743 (O_2743,N_23602,N_21591);
and UO_2744 (O_2744,N_21566,N_20736);
nor UO_2745 (O_2745,N_21893,N_20376);
xnor UO_2746 (O_2746,N_20845,N_21375);
xnor UO_2747 (O_2747,N_24451,N_20666);
or UO_2748 (O_2748,N_21541,N_21524);
or UO_2749 (O_2749,N_19215,N_23025);
and UO_2750 (O_2750,N_20639,N_24809);
or UO_2751 (O_2751,N_20531,N_23680);
nand UO_2752 (O_2752,N_23644,N_21842);
and UO_2753 (O_2753,N_24286,N_20986);
or UO_2754 (O_2754,N_20661,N_20183);
and UO_2755 (O_2755,N_21486,N_21995);
or UO_2756 (O_2756,N_20486,N_21713);
and UO_2757 (O_2757,N_21660,N_23184);
and UO_2758 (O_2758,N_19095,N_22255);
xnor UO_2759 (O_2759,N_24091,N_21173);
and UO_2760 (O_2760,N_22856,N_24057);
nor UO_2761 (O_2761,N_21681,N_22016);
nand UO_2762 (O_2762,N_19870,N_24895);
nor UO_2763 (O_2763,N_24459,N_20796);
nor UO_2764 (O_2764,N_21628,N_24370);
nand UO_2765 (O_2765,N_23509,N_23283);
and UO_2766 (O_2766,N_23334,N_20134);
nor UO_2767 (O_2767,N_23055,N_20192);
or UO_2768 (O_2768,N_22683,N_19845);
and UO_2769 (O_2769,N_19759,N_19657);
and UO_2770 (O_2770,N_22803,N_24635);
and UO_2771 (O_2771,N_22096,N_23364);
xor UO_2772 (O_2772,N_21614,N_21931);
xnor UO_2773 (O_2773,N_22925,N_20831);
or UO_2774 (O_2774,N_23341,N_19838);
xor UO_2775 (O_2775,N_21048,N_19776);
or UO_2776 (O_2776,N_19633,N_20570);
xnor UO_2777 (O_2777,N_22585,N_22436);
xor UO_2778 (O_2778,N_22155,N_19900);
nor UO_2779 (O_2779,N_18778,N_22727);
and UO_2780 (O_2780,N_19443,N_22684);
nand UO_2781 (O_2781,N_20385,N_21597);
nand UO_2782 (O_2782,N_21529,N_22839);
or UO_2783 (O_2783,N_18760,N_20334);
nand UO_2784 (O_2784,N_24756,N_24605);
nor UO_2785 (O_2785,N_19254,N_21084);
or UO_2786 (O_2786,N_22652,N_21948);
xor UO_2787 (O_2787,N_21737,N_22559);
nor UO_2788 (O_2788,N_21921,N_22414);
xnor UO_2789 (O_2789,N_21102,N_23518);
nor UO_2790 (O_2790,N_21444,N_24937);
or UO_2791 (O_2791,N_23268,N_22632);
and UO_2792 (O_2792,N_23510,N_20963);
or UO_2793 (O_2793,N_21565,N_22124);
nor UO_2794 (O_2794,N_23844,N_21260);
xor UO_2795 (O_2795,N_19188,N_21463);
or UO_2796 (O_2796,N_24919,N_20891);
and UO_2797 (O_2797,N_24647,N_22976);
or UO_2798 (O_2798,N_21082,N_20519);
and UO_2799 (O_2799,N_21379,N_23537);
nor UO_2800 (O_2800,N_23699,N_22402);
nand UO_2801 (O_2801,N_21633,N_21326);
nand UO_2802 (O_2802,N_23695,N_22060);
and UO_2803 (O_2803,N_23492,N_22526);
xnor UO_2804 (O_2804,N_20462,N_19391);
or UO_2805 (O_2805,N_20342,N_23561);
and UO_2806 (O_2806,N_19328,N_22101);
nor UO_2807 (O_2807,N_20508,N_21378);
and UO_2808 (O_2808,N_24984,N_24877);
nor UO_2809 (O_2809,N_22264,N_21070);
nor UO_2810 (O_2810,N_23497,N_23241);
nor UO_2811 (O_2811,N_21502,N_23928);
or UO_2812 (O_2812,N_18853,N_20548);
nand UO_2813 (O_2813,N_18904,N_23117);
xnor UO_2814 (O_2814,N_20776,N_20186);
nor UO_2815 (O_2815,N_23176,N_21925);
or UO_2816 (O_2816,N_24589,N_20816);
nand UO_2817 (O_2817,N_24762,N_22355);
or UO_2818 (O_2818,N_20850,N_19984);
nand UO_2819 (O_2819,N_23811,N_24950);
xnor UO_2820 (O_2820,N_21393,N_19990);
xor UO_2821 (O_2821,N_23530,N_20899);
or UO_2822 (O_2822,N_23127,N_19728);
and UO_2823 (O_2823,N_18796,N_22562);
and UO_2824 (O_2824,N_22618,N_22868);
xor UO_2825 (O_2825,N_19617,N_22886);
nor UO_2826 (O_2826,N_23833,N_24940);
or UO_2827 (O_2827,N_23310,N_20882);
nand UO_2828 (O_2828,N_19817,N_21603);
nor UO_2829 (O_2829,N_22578,N_21922);
xnor UO_2830 (O_2830,N_22958,N_21394);
nor UO_2831 (O_2831,N_22789,N_24385);
xor UO_2832 (O_2832,N_24630,N_23218);
and UO_2833 (O_2833,N_23266,N_21759);
nand UO_2834 (O_2834,N_21403,N_24570);
or UO_2835 (O_2835,N_20231,N_23944);
xnor UO_2836 (O_2836,N_21635,N_20044);
xnor UO_2837 (O_2837,N_21812,N_23098);
nor UO_2838 (O_2838,N_19736,N_21127);
and UO_2839 (O_2839,N_23506,N_20810);
nand UO_2840 (O_2840,N_19035,N_21193);
and UO_2841 (O_2841,N_23740,N_23981);
or UO_2842 (O_2842,N_19595,N_22498);
and UO_2843 (O_2843,N_22515,N_21020);
nand UO_2844 (O_2844,N_20883,N_22084);
nor UO_2845 (O_2845,N_21125,N_20463);
and UO_2846 (O_2846,N_20224,N_21884);
nand UO_2847 (O_2847,N_21094,N_19403);
nor UO_2848 (O_2848,N_22470,N_21158);
nand UO_2849 (O_2849,N_23513,N_19730);
xnor UO_2850 (O_2850,N_24805,N_19203);
and UO_2851 (O_2851,N_22399,N_22915);
or UO_2852 (O_2852,N_19495,N_22841);
xnor UO_2853 (O_2853,N_20770,N_22549);
xnor UO_2854 (O_2854,N_19651,N_20228);
nor UO_2855 (O_2855,N_23001,N_23129);
or UO_2856 (O_2856,N_23338,N_23132);
or UO_2857 (O_2857,N_21520,N_20020);
xnor UO_2858 (O_2858,N_24500,N_24040);
nor UO_2859 (O_2859,N_21228,N_22705);
nor UO_2860 (O_2860,N_24049,N_22943);
nand UO_2861 (O_2861,N_19017,N_23288);
nor UO_2862 (O_2862,N_19824,N_19048);
xor UO_2863 (O_2863,N_22588,N_24289);
nand UO_2864 (O_2864,N_22479,N_21553);
or UO_2865 (O_2865,N_23291,N_23970);
xnor UO_2866 (O_2866,N_24646,N_20258);
xor UO_2867 (O_2867,N_20607,N_19485);
nor UO_2868 (O_2868,N_20584,N_22462);
and UO_2869 (O_2869,N_23436,N_23327);
nand UO_2870 (O_2870,N_22083,N_19329);
nand UO_2871 (O_2871,N_20002,N_23150);
and UO_2872 (O_2872,N_21399,N_20914);
nand UO_2873 (O_2873,N_19538,N_21655);
and UO_2874 (O_2874,N_22895,N_21773);
xor UO_2875 (O_2875,N_21161,N_19965);
xnor UO_2876 (O_2876,N_24169,N_22896);
or UO_2877 (O_2877,N_19598,N_20271);
or UO_2878 (O_2878,N_21798,N_20456);
nor UO_2879 (O_2879,N_18775,N_19787);
nand UO_2880 (O_2880,N_21709,N_23469);
nor UO_2881 (O_2881,N_19373,N_23121);
nor UO_2882 (O_2882,N_22127,N_21131);
or UO_2883 (O_2883,N_24368,N_19250);
and UO_2884 (O_2884,N_18783,N_19734);
xnor UO_2885 (O_2885,N_22469,N_19100);
or UO_2886 (O_2886,N_19822,N_20246);
xor UO_2887 (O_2887,N_23857,N_24114);
or UO_2888 (O_2888,N_22295,N_20973);
and UO_2889 (O_2889,N_24936,N_22587);
nor UO_2890 (O_2890,N_23242,N_21971);
or UO_2891 (O_2891,N_23896,N_23409);
nand UO_2892 (O_2892,N_24706,N_22107);
nand UO_2893 (O_2893,N_21174,N_24566);
nor UO_2894 (O_2894,N_19951,N_22872);
nor UO_2895 (O_2895,N_18991,N_22336);
and UO_2896 (O_2896,N_21977,N_20114);
xnor UO_2897 (O_2897,N_23175,N_18885);
or UO_2898 (O_2898,N_19777,N_19727);
xnor UO_2899 (O_2899,N_24389,N_22437);
xor UO_2900 (O_2900,N_24290,N_24177);
xor UO_2901 (O_2901,N_21554,N_18891);
nand UO_2902 (O_2902,N_20126,N_19568);
nand UO_2903 (O_2903,N_24362,N_20645);
and UO_2904 (O_2904,N_19804,N_23578);
or UO_2905 (O_2905,N_24820,N_18822);
or UO_2906 (O_2906,N_23682,N_21777);
and UO_2907 (O_2907,N_22279,N_21490);
nand UO_2908 (O_2908,N_18893,N_18843);
or UO_2909 (O_2909,N_20354,N_19064);
or UO_2910 (O_2910,N_20669,N_20163);
nand UO_2911 (O_2911,N_24491,N_21201);
xor UO_2912 (O_2912,N_19533,N_23304);
or UO_2913 (O_2913,N_24407,N_22795);
nand UO_2914 (O_2914,N_23566,N_24614);
and UO_2915 (O_2915,N_19973,N_22011);
nor UO_2916 (O_2916,N_23066,N_23263);
or UO_2917 (O_2917,N_22196,N_21650);
nand UO_2918 (O_2918,N_24839,N_24247);
nand UO_2919 (O_2919,N_22487,N_19917);
and UO_2920 (O_2920,N_19939,N_22455);
or UO_2921 (O_2921,N_22653,N_23744);
nor UO_2922 (O_2922,N_23823,N_22908);
nand UO_2923 (O_2923,N_21906,N_20829);
or UO_2924 (O_2924,N_21063,N_24374);
nor UO_2925 (O_2925,N_21976,N_23880);
and UO_2926 (O_2926,N_21564,N_18871);
nor UO_2927 (O_2927,N_21236,N_24377);
and UO_2928 (O_2928,N_19451,N_21389);
nor UO_2929 (O_2929,N_22163,N_23020);
xor UO_2930 (O_2930,N_21612,N_20922);
nor UO_2931 (O_2931,N_20270,N_19775);
or UO_2932 (O_2932,N_22924,N_21792);
and UO_2933 (O_2933,N_20435,N_21877);
or UO_2934 (O_2934,N_22170,N_19862);
or UO_2935 (O_2935,N_21910,N_20344);
nor UO_2936 (O_2936,N_21334,N_19924);
xor UO_2937 (O_2937,N_23728,N_22530);
nor UO_2938 (O_2938,N_23217,N_19128);
xnor UO_2939 (O_2939,N_23423,N_20874);
and UO_2940 (O_2940,N_23214,N_21561);
nand UO_2941 (O_2941,N_24309,N_23008);
xnor UO_2942 (O_2942,N_19522,N_23835);
or UO_2943 (O_2943,N_19709,N_21702);
and UO_2944 (O_2944,N_20679,N_22093);
nand UO_2945 (O_2945,N_19642,N_20452);
nor UO_2946 (O_2946,N_20343,N_22261);
nand UO_2947 (O_2947,N_21427,N_23315);
nor UO_2948 (O_2948,N_22228,N_23148);
xnor UO_2949 (O_2949,N_21944,N_19549);
xor UO_2950 (O_2950,N_22542,N_22190);
xnor UO_2951 (O_2951,N_20237,N_22503);
xnor UO_2952 (O_2952,N_23508,N_24705);
and UO_2953 (O_2953,N_22961,N_23163);
nor UO_2954 (O_2954,N_19465,N_20417);
nor UO_2955 (O_2955,N_21665,N_23325);
and UO_2956 (O_2956,N_20983,N_22643);
xor UO_2957 (O_2957,N_21966,N_23799);
nor UO_2958 (O_2958,N_20170,N_22978);
xor UO_2959 (O_2959,N_19912,N_21711);
and UO_2960 (O_2960,N_21935,N_20636);
nor UO_2961 (O_2961,N_22419,N_22209);
and UO_2962 (O_2962,N_18832,N_20205);
xnor UO_2963 (O_2963,N_21415,N_20852);
and UO_2964 (O_2964,N_23103,N_24107);
nor UO_2965 (O_2965,N_22953,N_19371);
nand UO_2966 (O_2966,N_18909,N_21588);
or UO_2967 (O_2967,N_24119,N_24027);
and UO_2968 (O_2968,N_24218,N_18961);
nand UO_2969 (O_2969,N_24130,N_20652);
xor UO_2970 (O_2970,N_18810,N_22078);
or UO_2971 (O_2971,N_23984,N_22782);
xor UO_2972 (O_2972,N_24384,N_21498);
and UO_2973 (O_2973,N_24445,N_20034);
nor UO_2974 (O_2974,N_19260,N_19294);
nand UO_2975 (O_2975,N_18957,N_19892);
nand UO_2976 (O_2976,N_19297,N_24980);
or UO_2977 (O_2977,N_24945,N_21568);
nand UO_2978 (O_2978,N_22995,N_24125);
and UO_2979 (O_2979,N_23582,N_21188);
nor UO_2980 (O_2980,N_24258,N_22381);
xnor UO_2981 (O_2981,N_21762,N_22620);
xnor UO_2982 (O_2982,N_21409,N_20634);
nor UO_2983 (O_2983,N_22914,N_24005);
or UO_2984 (O_2984,N_20308,N_22348);
or UO_2985 (O_2985,N_20442,N_20287);
nor UO_2986 (O_2986,N_24067,N_24302);
and UO_2987 (O_2987,N_22433,N_23558);
nand UO_2988 (O_2988,N_23297,N_23406);
xnor UO_2989 (O_2989,N_22994,N_20637);
or UO_2990 (O_2990,N_24026,N_21784);
and UO_2991 (O_2991,N_24480,N_24516);
or UO_2992 (O_2992,N_20984,N_24068);
and UO_2993 (O_2993,N_20856,N_19065);
nor UO_2994 (O_2994,N_19086,N_22216);
nor UO_2995 (O_2995,N_22579,N_24874);
or UO_2996 (O_2996,N_19018,N_22146);
xnor UO_2997 (O_2997,N_24386,N_20608);
or UO_2998 (O_2998,N_21288,N_22183);
nand UO_2999 (O_2999,N_24204,N_21171);
endmodule