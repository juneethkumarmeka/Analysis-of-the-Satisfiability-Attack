module basic_1500_15000_2000_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_367,In_567);
xnor U1 (N_1,In_548,In_60);
xnor U2 (N_2,In_1147,In_971);
or U3 (N_3,In_1129,In_472);
and U4 (N_4,In_1125,In_1341);
xor U5 (N_5,In_1042,In_1300);
or U6 (N_6,In_599,In_258);
nor U7 (N_7,In_494,In_1224);
or U8 (N_8,In_1182,In_1259);
nor U9 (N_9,In_90,In_1239);
nor U10 (N_10,In_732,In_1005);
xnor U11 (N_11,In_293,In_1396);
nand U12 (N_12,In_937,In_38);
nand U13 (N_13,In_825,In_1170);
nor U14 (N_14,In_1433,In_1205);
or U15 (N_15,In_861,In_1212);
or U16 (N_16,In_1377,In_778);
xor U17 (N_17,In_1420,In_102);
or U18 (N_18,In_1149,In_650);
or U19 (N_19,In_451,In_975);
nor U20 (N_20,In_1288,In_1492);
nor U21 (N_21,In_668,In_680);
and U22 (N_22,In_14,In_974);
xnor U23 (N_23,In_1049,In_1380);
or U24 (N_24,In_1160,In_560);
or U25 (N_25,In_233,In_432);
xnor U26 (N_26,In_192,In_268);
xnor U27 (N_27,In_1483,In_710);
or U28 (N_28,In_346,In_588);
or U29 (N_29,In_1017,In_566);
and U30 (N_30,In_312,In_1027);
xnor U31 (N_31,In_523,In_608);
nand U32 (N_32,In_2,In_744);
nor U33 (N_33,In_927,In_340);
xor U34 (N_34,In_594,In_1355);
xnor U35 (N_35,In_966,In_1207);
nor U36 (N_36,In_748,In_525);
nand U37 (N_37,In_474,In_799);
nor U38 (N_38,In_457,In_1326);
xnor U39 (N_39,In_1011,In_1335);
xnor U40 (N_40,In_1385,In_1194);
xnor U41 (N_41,In_168,In_513);
or U42 (N_42,In_465,In_23);
and U43 (N_43,In_953,In_1436);
xnor U44 (N_44,In_1104,In_662);
xnor U45 (N_45,In_185,In_46);
or U46 (N_46,In_73,In_1426);
or U47 (N_47,In_325,In_481);
or U48 (N_48,In_1280,In_1057);
nand U49 (N_49,In_1107,In_1251);
and U50 (N_50,In_806,In_1046);
nor U51 (N_51,In_1367,In_1219);
or U52 (N_52,In_917,In_1020);
and U53 (N_53,In_967,In_453);
xor U54 (N_54,In_1325,In_1139);
nor U55 (N_55,In_1093,In_94);
and U56 (N_56,In_285,In_106);
or U57 (N_57,In_1068,In_1279);
nor U58 (N_58,In_1069,In_323);
or U59 (N_59,In_657,In_78);
and U60 (N_60,In_1465,In_561);
and U61 (N_61,In_960,In_1254);
xor U62 (N_62,In_549,In_786);
nand U63 (N_63,In_190,In_303);
nand U64 (N_64,In_1430,In_291);
or U65 (N_65,In_981,In_213);
and U66 (N_66,In_123,In_243);
or U67 (N_67,In_762,In_843);
nor U68 (N_68,In_1499,In_507);
nand U69 (N_69,In_1284,In_893);
or U70 (N_70,In_909,In_932);
and U71 (N_71,In_961,In_477);
and U72 (N_72,In_512,In_1120);
nand U73 (N_73,In_332,In_829);
and U74 (N_74,In_1371,In_658);
and U75 (N_75,In_505,In_411);
and U76 (N_76,In_814,In_1099);
nor U77 (N_77,In_1271,In_832);
or U78 (N_78,In_812,In_272);
nor U79 (N_79,In_1175,In_121);
nand U80 (N_80,In_93,In_1432);
nor U81 (N_81,In_946,In_375);
xor U82 (N_82,In_1322,In_1001);
nand U83 (N_83,In_441,In_200);
nor U84 (N_84,In_1378,In_1350);
nand U85 (N_85,In_1275,In_1313);
or U86 (N_86,In_1282,In_818);
nor U87 (N_87,In_1413,In_1406);
nand U88 (N_88,In_313,In_467);
nand U89 (N_89,In_621,In_508);
or U90 (N_90,In_1301,In_1272);
xnor U91 (N_91,In_585,In_654);
xnor U92 (N_92,In_924,In_579);
xor U93 (N_93,In_826,In_464);
and U94 (N_94,In_898,In_434);
nand U95 (N_95,In_498,In_553);
and U96 (N_96,In_18,In_1395);
xnor U97 (N_97,In_1181,In_1050);
nor U98 (N_98,In_386,In_1014);
nor U99 (N_99,In_1145,In_835);
nor U100 (N_100,In_807,In_796);
and U101 (N_101,In_338,In_150);
or U102 (N_102,In_667,In_1333);
or U103 (N_103,In_1091,In_840);
and U104 (N_104,In_906,In_554);
nor U105 (N_105,In_99,In_219);
xnor U106 (N_106,In_759,In_701);
and U107 (N_107,In_968,In_1489);
or U108 (N_108,In_1403,In_724);
nand U109 (N_109,In_1415,In_334);
or U110 (N_110,In_1138,In_1257);
or U111 (N_111,In_808,In_872);
nand U112 (N_112,In_188,In_536);
and U113 (N_113,In_161,In_831);
or U114 (N_114,In_1281,In_563);
xnor U115 (N_115,In_930,In_879);
nor U116 (N_116,In_1440,In_717);
nand U117 (N_117,In_1051,In_128);
xor U118 (N_118,In_857,In_177);
and U119 (N_119,In_938,In_805);
nand U120 (N_120,In_1445,In_478);
nand U121 (N_121,In_297,In_230);
xor U122 (N_122,In_506,In_1043);
or U123 (N_123,In_35,In_1374);
nand U124 (N_124,In_1073,In_1060);
xnor U125 (N_125,In_765,In_965);
xor U126 (N_126,In_1185,In_207);
and U127 (N_127,In_844,In_922);
nor U128 (N_128,In_392,In_1189);
xnor U129 (N_129,In_1140,In_302);
xor U130 (N_130,In_499,In_1235);
xor U131 (N_131,In_152,In_570);
nand U132 (N_132,In_604,In_811);
nand U133 (N_133,In_398,In_845);
nand U134 (N_134,In_624,In_286);
nand U135 (N_135,In_1067,In_1278);
or U136 (N_136,In_3,In_56);
nor U137 (N_137,In_1383,In_714);
or U138 (N_138,In_1299,In_289);
or U139 (N_139,In_307,In_1242);
xor U140 (N_140,In_605,In_823);
nand U141 (N_141,In_1118,In_127);
nand U142 (N_142,In_619,In_795);
and U143 (N_143,In_1464,In_26);
and U144 (N_144,In_859,In_4);
and U145 (N_145,In_888,In_694);
and U146 (N_146,In_42,In_851);
nor U147 (N_147,In_1334,In_834);
or U148 (N_148,In_901,In_53);
and U149 (N_149,In_260,In_389);
and U150 (N_150,In_1066,In_1006);
nand U151 (N_151,In_600,In_562);
and U152 (N_152,In_1382,In_1191);
nand U153 (N_153,In_582,In_1110);
or U154 (N_154,In_887,In_734);
xor U155 (N_155,In_1443,In_659);
nand U156 (N_156,In_727,In_993);
nor U157 (N_157,In_458,In_1037);
nand U158 (N_158,In_841,In_992);
or U159 (N_159,In_883,In_1405);
nand U160 (N_160,In_125,In_584);
xor U161 (N_161,In_257,In_96);
nor U162 (N_162,In_1086,In_596);
nor U163 (N_163,In_1096,In_1474);
or U164 (N_164,In_417,In_1030);
and U165 (N_165,In_679,In_1345);
and U166 (N_166,In_141,In_743);
nand U167 (N_167,In_419,In_983);
nand U168 (N_168,In_856,In_139);
and U169 (N_169,In_1400,In_810);
and U170 (N_170,In_269,In_294);
nor U171 (N_171,In_858,In_1173);
or U172 (N_172,In_707,In_1152);
nor U173 (N_173,In_670,In_437);
and U174 (N_174,In_785,In_1021);
or U175 (N_175,In_1485,In_189);
nor U176 (N_176,In_160,In_578);
and U177 (N_177,In_1270,In_897);
or U178 (N_178,In_1477,In_544);
nor U179 (N_179,In_638,In_1058);
or U180 (N_180,In_357,In_178);
nor U181 (N_181,In_1157,In_319);
and U182 (N_182,In_745,In_822);
xor U183 (N_183,In_1018,In_763);
nand U184 (N_184,In_1421,In_1079);
nor U185 (N_185,In_1461,In_698);
or U186 (N_186,In_645,In_74);
nor U187 (N_187,In_98,In_708);
and U188 (N_188,In_49,In_214);
nor U189 (N_189,In_144,In_774);
nand U190 (N_190,In_5,In_25);
and U191 (N_191,In_1055,In_275);
nand U192 (N_192,In_730,In_138);
nand U193 (N_193,In_1358,In_697);
nor U194 (N_194,In_1494,In_251);
nor U195 (N_195,In_852,In_1065);
or U196 (N_196,In_1187,In_1309);
xnor U197 (N_197,In_410,In_800);
or U198 (N_198,In_767,In_1316);
and U199 (N_199,In_663,In_700);
xor U200 (N_200,In_438,In_84);
xnor U201 (N_201,In_997,In_9);
and U202 (N_202,In_1158,In_347);
or U203 (N_203,In_590,In_1431);
nor U204 (N_204,In_1101,In_719);
nor U205 (N_205,In_267,In_404);
xnor U206 (N_206,In_1416,In_991);
or U207 (N_207,In_385,In_12);
and U208 (N_208,In_1386,In_833);
and U209 (N_209,In_327,In_413);
and U210 (N_210,In_401,In_1072);
xor U211 (N_211,In_364,In_1211);
nor U212 (N_212,In_1491,In_1019);
and U213 (N_213,In_839,In_172);
or U214 (N_214,In_746,In_374);
nor U215 (N_215,In_109,In_1487);
nor U216 (N_216,In_119,In_476);
nor U217 (N_217,In_381,In_480);
nor U218 (N_218,In_819,In_140);
nand U219 (N_219,In_244,In_1336);
and U220 (N_220,In_1,In_925);
and U221 (N_221,In_736,In_36);
xor U222 (N_222,In_43,In_784);
nor U223 (N_223,In_950,In_672);
nand U224 (N_224,In_963,In_1230);
and U225 (N_225,In_1444,In_798);
and U226 (N_226,In_706,In_1372);
nand U227 (N_227,In_820,In_195);
and U228 (N_228,In_878,In_299);
and U229 (N_229,In_637,In_830);
or U230 (N_230,In_7,In_1004);
nor U231 (N_231,In_1222,In_627);
or U232 (N_232,In_1090,In_628);
xor U233 (N_233,In_1266,In_1202);
and U234 (N_234,In_910,In_452);
xor U235 (N_235,In_1226,In_328);
nand U236 (N_236,In_283,In_980);
and U237 (N_237,In_962,In_130);
nand U238 (N_238,In_500,In_871);
nor U239 (N_239,In_41,In_905);
xor U240 (N_240,In_341,In_685);
nand U241 (N_241,In_174,In_253);
nand U242 (N_242,In_634,In_552);
xnor U243 (N_243,In_528,In_1470);
xor U244 (N_244,In_58,In_315);
xor U245 (N_245,In_133,In_492);
xor U246 (N_246,In_827,In_1076);
xnor U247 (N_247,In_540,In_1319);
or U248 (N_248,In_288,In_935);
or U249 (N_249,In_179,In_330);
nor U250 (N_250,In_229,In_1250);
and U251 (N_251,In_186,In_39);
or U252 (N_252,In_40,In_1100);
nor U253 (N_253,In_914,In_1340);
or U254 (N_254,In_331,In_1344);
or U255 (N_255,In_169,In_1032);
nor U256 (N_256,In_1171,In_69);
and U257 (N_257,In_1277,In_1010);
and U258 (N_258,In_716,In_202);
and U259 (N_259,In_1089,In_1248);
xor U260 (N_260,In_1388,In_1304);
or U261 (N_261,In_1422,In_1039);
nand U262 (N_262,In_1478,In_71);
or U263 (N_263,In_723,In_815);
and U264 (N_264,In_661,In_921);
or U265 (N_265,In_739,In_171);
xnor U266 (N_266,In_1407,In_1169);
or U267 (N_267,In_148,In_326);
nand U268 (N_268,In_769,In_1390);
nor U269 (N_269,In_1201,In_606);
nor U270 (N_270,In_1126,In_447);
nand U271 (N_271,In_1484,In_320);
xnor U272 (N_272,In_920,In_1490);
or U273 (N_273,In_50,In_222);
and U274 (N_274,In_1119,In_234);
nor U275 (N_275,In_1190,In_20);
xor U276 (N_276,In_1085,In_273);
xor U277 (N_277,In_67,In_300);
and U278 (N_278,In_550,In_82);
nor U279 (N_279,In_713,In_445);
nand U280 (N_280,In_754,In_757);
and U281 (N_281,In_255,In_352);
or U282 (N_282,In_1314,In_31);
nand U283 (N_283,In_95,In_532);
nand U284 (N_284,In_1134,In_866);
or U285 (N_285,In_354,In_240);
or U286 (N_286,In_136,In_1303);
nand U287 (N_287,In_1476,In_1246);
xnor U288 (N_288,In_1293,In_522);
nand U289 (N_289,In_1176,In_1197);
xnor U290 (N_290,In_985,In_1144);
nor U291 (N_291,In_193,In_249);
nor U292 (N_292,In_1151,In_206);
nor U293 (N_293,In_1297,In_919);
nand U294 (N_294,In_166,In_1462);
nor U295 (N_295,In_649,In_1273);
and U296 (N_296,In_1408,In_693);
or U297 (N_297,In_1180,In_583);
xor U298 (N_298,In_753,In_1497);
nor U299 (N_299,In_68,In_59);
or U300 (N_300,In_837,In_978);
or U301 (N_301,In_1368,N_148);
xor U302 (N_302,N_27,In_613);
nand U303 (N_303,In_1285,In_1123);
xor U304 (N_304,In_1296,In_1327);
nor U305 (N_305,In_836,In_855);
xnor U306 (N_306,In_1074,N_183);
nand U307 (N_307,N_12,In_65);
nor U308 (N_308,In_502,N_188);
nor U309 (N_309,In_1238,N_18);
and U310 (N_310,In_482,In_115);
xor U311 (N_311,N_237,N_10);
nand U312 (N_312,N_286,In_1456);
xor U313 (N_313,In_1264,In_651);
and U314 (N_314,In_362,In_609);
nand U315 (N_315,N_245,In_460);
nand U316 (N_316,In_231,In_644);
xor U317 (N_317,N_150,N_99);
nor U318 (N_318,In_55,N_78);
nand U319 (N_319,N_111,N_109);
xnor U320 (N_320,N_163,In_509);
or U321 (N_321,In_54,In_768);
nor U322 (N_322,N_107,In_252);
nor U323 (N_323,In_51,In_117);
or U324 (N_324,N_221,In_394);
and U325 (N_325,In_1379,In_24);
nor U326 (N_326,In_1389,In_564);
xor U327 (N_327,N_66,In_1471);
nor U328 (N_328,In_868,In_1486);
xor U329 (N_329,N_205,In_317);
and U330 (N_330,In_597,N_159);
and U331 (N_331,N_28,In_863);
and U332 (N_332,In_1357,In_225);
nor U333 (N_333,In_199,In_85);
and U334 (N_334,In_1262,In_1381);
nand U335 (N_335,In_239,In_660);
nand U336 (N_336,In_1150,In_1351);
nand U337 (N_337,In_1342,N_24);
xnor U338 (N_338,In_629,In_1214);
and U339 (N_339,In_862,In_940);
xnor U340 (N_340,In_221,In_1061);
and U341 (N_341,In_137,N_142);
nor U342 (N_342,In_626,N_64);
and U343 (N_343,In_789,In_1466);
or U344 (N_344,N_83,N_141);
nand U345 (N_345,In_1056,In_1034);
and U346 (N_346,N_226,In_704);
nor U347 (N_347,In_747,In_1206);
xnor U348 (N_348,N_235,In_1328);
nor U349 (N_349,In_388,In_310);
xor U350 (N_350,N_70,N_283);
and U351 (N_351,In_918,In_37);
xor U352 (N_352,In_1449,N_181);
or U353 (N_353,In_1063,In_1132);
and U354 (N_354,In_1276,In_489);
or U355 (N_355,In_1164,N_57);
xnor U356 (N_356,N_184,In_537);
xor U357 (N_357,N_23,In_265);
and U358 (N_358,In_1412,N_165);
xnor U359 (N_359,In_1343,In_503);
nor U360 (N_360,In_764,In_13);
and U361 (N_361,In_1114,In_790);
and U362 (N_362,In_729,In_1012);
xor U363 (N_363,In_10,N_96);
and U364 (N_364,In_170,In_895);
and U365 (N_365,N_122,In_1044);
or U366 (N_366,In_83,N_198);
or U367 (N_367,In_8,In_1243);
nor U368 (N_368,In_620,In_643);
nand U369 (N_369,In_1221,In_876);
nand U370 (N_370,N_115,In_737);
or U371 (N_371,In_1493,In_281);
xor U372 (N_372,N_192,N_131);
nor U373 (N_373,In_1035,In_865);
or U374 (N_374,N_285,In_414);
and U375 (N_375,N_217,In_271);
xor U376 (N_376,In_1031,N_259);
xor U377 (N_377,In_903,N_50);
xor U378 (N_378,In_783,In_400);
or U379 (N_379,In_816,In_828);
xnor U380 (N_380,In_21,In_690);
and U381 (N_381,In_952,In_1256);
nor U382 (N_382,In_692,In_1215);
and U383 (N_383,In_776,N_292);
or U384 (N_384,In_402,In_1399);
and U385 (N_385,In_781,In_1302);
or U386 (N_386,N_95,In_390);
and U387 (N_387,N_194,In_486);
and U388 (N_388,In_423,In_555);
nand U389 (N_389,In_1016,In_408);
and U390 (N_390,In_777,In_22);
nor U391 (N_391,In_359,In_89);
nand U392 (N_392,In_568,In_351);
nand U393 (N_393,N_31,In_1209);
and U394 (N_394,In_397,In_1041);
nand U395 (N_395,In_1295,In_422);
xor U396 (N_396,In_151,N_21);
nor U397 (N_397,In_237,In_803);
nor U398 (N_398,N_253,In_1071);
nor U399 (N_399,In_1231,In_979);
nor U400 (N_400,In_145,In_490);
nand U401 (N_401,In_173,In_556);
nor U402 (N_402,In_1115,N_121);
or U403 (N_403,In_1424,N_74);
nor U404 (N_404,N_118,In_902);
and U405 (N_405,In_899,In_6);
or U406 (N_406,In_741,In_682);
or U407 (N_407,N_102,In_733);
nor U408 (N_408,In_142,In_569);
xor U409 (N_409,N_3,In_614);
nand U410 (N_410,N_166,In_1143);
nor U411 (N_411,In_132,In_154);
nand U412 (N_412,N_45,In_396);
and U413 (N_413,In_454,In_1495);
or U414 (N_414,In_470,N_8);
xor U415 (N_415,N_42,In_616);
nand U416 (N_416,In_495,In_994);
and U417 (N_417,N_49,N_230);
and U418 (N_418,In_70,In_377);
and U419 (N_419,In_1167,In_873);
nor U420 (N_420,In_62,In_589);
nand U421 (N_421,In_1003,In_1448);
nand U422 (N_422,In_1080,N_263);
or U423 (N_423,N_227,In_1261);
nor U424 (N_424,In_223,In_944);
and U425 (N_425,In_131,In_1346);
nor U426 (N_426,In_107,In_683);
xor U427 (N_427,In_514,In_1227);
xnor U428 (N_428,In_301,N_160);
xnor U429 (N_429,N_179,In_314);
nand U430 (N_430,N_269,In_1359);
nand U431 (N_431,In_247,In_665);
and U432 (N_432,In_676,In_874);
xnor U433 (N_433,In_175,In_456);
nor U434 (N_434,In_538,In_211);
xnor U435 (N_435,In_1233,N_9);
or U436 (N_436,In_949,N_176);
and U437 (N_437,In_382,In_1365);
xnor U438 (N_438,N_252,In_63);
nand U439 (N_439,In_1193,In_1105);
and U440 (N_440,In_1418,In_262);
nor U441 (N_441,In_656,In_787);
xor U442 (N_442,N_215,In_959);
nand U443 (N_443,In_760,In_1216);
and U444 (N_444,In_424,N_151);
nand U445 (N_445,N_88,In_116);
or U446 (N_446,In_504,In_112);
and U447 (N_447,N_129,In_1198);
nor U448 (N_448,In_854,In_546);
nand U449 (N_449,In_571,In_421);
nand U450 (N_450,N_229,In_1229);
xnor U451 (N_451,In_666,In_1232);
xor U452 (N_452,In_19,In_156);
nor U453 (N_453,In_1458,In_821);
and U454 (N_454,In_196,N_287);
or U455 (N_455,N_276,In_487);
or U456 (N_456,In_1361,In_1108);
and U457 (N_457,In_279,In_120);
nor U458 (N_458,In_970,In_740);
nand U459 (N_459,In_720,In_797);
nor U460 (N_460,N_267,In_162);
nor U461 (N_461,In_270,In_804);
xor U462 (N_462,In_973,In_407);
nor U463 (N_463,N_202,In_488);
nor U464 (N_464,In_542,In_471);
or U465 (N_465,In_129,In_122);
and U466 (N_466,In_877,In_1393);
or U467 (N_467,In_587,In_1077);
or U468 (N_468,In_34,In_999);
or U469 (N_469,In_248,In_576);
and U470 (N_470,In_603,In_1059);
or U471 (N_471,In_306,In_1468);
nand U472 (N_472,In_365,In_731);
nand U473 (N_473,In_1124,In_1136);
xor U474 (N_474,In_100,In_435);
or U475 (N_475,In_850,N_145);
nand U476 (N_476,In_1457,In_860);
or U477 (N_477,N_69,In_61);
and U478 (N_478,In_32,In_337);
nor U479 (N_479,In_750,In_368);
or U480 (N_480,In_220,In_1161);
xnor U481 (N_481,In_551,N_193);
xnor U482 (N_482,N_11,In_324);
or U483 (N_483,In_591,In_915);
nand U484 (N_484,N_47,In_515);
nand U485 (N_485,N_182,In_1204);
nor U486 (N_486,In_1064,N_92);
nand U487 (N_487,In_355,In_403);
or U488 (N_488,In_228,N_275);
and U489 (N_489,In_527,In_900);
xor U490 (N_490,In_430,In_485);
xor U491 (N_491,In_1404,In_611);
nor U492 (N_492,In_420,In_383);
nand U493 (N_493,In_1081,In_1172);
or U494 (N_494,In_1447,In_755);
or U495 (N_495,N_25,In_889);
xnor U496 (N_496,In_964,N_297);
xor U497 (N_497,In_573,In_241);
or U498 (N_498,N_146,N_258);
or U499 (N_499,In_517,In_1425);
or U500 (N_500,In_1347,N_132);
nor U501 (N_501,In_146,In_436);
and U502 (N_502,In_1310,N_97);
nor U503 (N_503,In_907,N_56);
or U504 (N_504,N_153,N_257);
and U505 (N_505,N_261,N_250);
nor U506 (N_506,In_203,In_418);
or U507 (N_507,In_1053,N_123);
or U508 (N_508,In_1442,In_1305);
xnor U509 (N_509,In_847,In_216);
xnor U510 (N_510,In_1323,N_41);
nand U511 (N_511,In_602,In_1435);
and U512 (N_512,In_1146,N_4);
and U513 (N_513,In_1363,In_1122);
nand U514 (N_514,N_117,In_1481);
and U515 (N_515,N_295,In_224);
xor U516 (N_516,In_1247,N_67);
nor U517 (N_517,In_44,In_143);
xnor U518 (N_518,In_1103,In_771);
and U519 (N_519,In_48,N_65);
nand U520 (N_520,In_1133,In_75);
or U521 (N_521,In_735,In_473);
nor U522 (N_522,In_469,N_281);
or U523 (N_523,In_1217,In_110);
xnor U524 (N_524,In_809,N_91);
nand U525 (N_525,In_788,In_881);
xnor U526 (N_526,In_882,In_756);
nand U527 (N_527,N_242,In_995);
nor U528 (N_528,N_232,In_1166);
or U529 (N_529,N_265,In_1312);
or U530 (N_530,In_880,In_1223);
nor U531 (N_531,In_531,In_529);
or U532 (N_532,In_632,In_846);
nand U533 (N_533,In_709,In_598);
and U534 (N_534,In_442,N_254);
nor U535 (N_535,In_976,In_1409);
nand U536 (N_536,N_278,N_211);
and U537 (N_537,In_577,In_321);
or U538 (N_538,In_886,In_80);
nand U539 (N_539,In_1135,In_673);
and U540 (N_540,In_1225,In_1070);
nor U541 (N_541,In_1200,In_593);
nand U542 (N_542,In_664,In_1291);
nor U543 (N_543,In_1289,In_344);
or U544 (N_544,In_1163,In_982);
and U545 (N_545,In_678,In_111);
nor U546 (N_546,In_1315,In_1045);
nand U547 (N_547,In_66,N_260);
nor U548 (N_548,In_1318,In_1029);
xor U549 (N_549,N_294,In_449);
and U550 (N_550,In_718,In_444);
and U551 (N_551,In_105,In_1268);
and U552 (N_552,N_234,In_1240);
or U553 (N_553,In_1084,N_1);
and U554 (N_554,N_206,In_1048);
or U555 (N_555,N_108,In_1178);
and U556 (N_556,In_945,In_998);
and U557 (N_557,In_163,In_227);
and U558 (N_558,In_715,In_1094);
nor U559 (N_559,N_246,N_207);
nand U560 (N_560,In_232,N_36);
or U561 (N_561,In_86,In_1088);
nand U562 (N_562,N_55,In_384);
xor U563 (N_563,In_284,In_926);
xor U564 (N_564,In_164,N_251);
or U565 (N_565,In_1128,In_671);
or U566 (N_566,In_391,N_264);
xnor U567 (N_567,In_1002,In_250);
or U568 (N_568,In_580,In_165);
and U569 (N_569,In_1213,In_305);
or U570 (N_570,In_28,In_316);
and U571 (N_571,In_380,In_647);
nor U572 (N_572,N_60,In_1362);
xnor U573 (N_573,In_936,N_175);
nor U574 (N_574,In_943,In_565);
or U575 (N_575,N_214,N_86);
or U576 (N_576,N_93,In_101);
and U577 (N_577,In_235,In_181);
and U578 (N_578,In_575,In_1253);
xnor U579 (N_579,In_183,N_255);
xor U580 (N_580,N_75,N_296);
and U581 (N_581,In_631,N_233);
xnor U582 (N_582,In_1195,N_219);
and U583 (N_583,In_496,In_1402);
and U584 (N_584,N_274,N_19);
nor U585 (N_585,In_853,In_1098);
xnor U586 (N_586,In_1036,N_225);
nand U587 (N_587,N_53,N_29);
nand U588 (N_588,N_52,In_1286);
and U589 (N_589,N_162,In_1475);
nand U590 (N_590,N_244,N_218);
and U591 (N_591,In_824,In_108);
xor U592 (N_592,In_1102,N_22);
nor U593 (N_593,In_440,N_293);
nand U594 (N_594,In_791,N_236);
nand U595 (N_595,In_483,In_295);
or U596 (N_596,N_105,In_817);
xor U597 (N_597,In_1498,In_842);
and U598 (N_598,N_197,In_989);
and U599 (N_599,In_526,In_209);
or U600 (N_600,N_200,N_509);
nor U601 (N_601,In_1454,N_481);
nor U602 (N_602,In_409,N_310);
nor U603 (N_603,In_610,N_85);
or U604 (N_604,In_468,In_1113);
nand U605 (N_605,N_30,N_270);
nand U606 (N_606,N_138,In_705);
xor U607 (N_607,N_135,In_1141);
nor U608 (N_608,In_1130,N_305);
and U609 (N_609,In_124,N_228);
nand U610 (N_610,In_1000,In_612);
or U611 (N_611,In_1075,In_911);
or U612 (N_612,N_389,In_615);
nor U613 (N_613,In_1112,N_539);
or U614 (N_614,N_386,In_1083);
nand U615 (N_615,In_88,In_521);
or U616 (N_616,N_341,In_292);
nor U617 (N_617,N_119,N_548);
nand U618 (N_618,N_478,N_411);
and U619 (N_619,In_545,In_29);
nand U620 (N_620,N_144,N_407);
nor U621 (N_621,N_409,In_1263);
nand U622 (N_622,In_1387,In_557);
or U623 (N_623,In_1427,N_445);
or U624 (N_624,N_337,In_52);
and U625 (N_625,In_1024,In_439);
and U626 (N_626,In_641,In_543);
nor U627 (N_627,N_101,N_14);
and U628 (N_628,N_403,In_1087);
or U629 (N_629,N_32,N_26);
nor U630 (N_630,In_412,N_213);
nand U631 (N_631,N_579,In_1353);
and U632 (N_632,N_515,In_113);
xnor U633 (N_633,In_493,In_1236);
or U634 (N_634,In_928,N_266);
and U635 (N_635,N_262,In_934);
nand U636 (N_636,In_201,In_1463);
nand U637 (N_637,N_447,N_171);
xor U638 (N_638,N_503,N_470);
and U639 (N_639,N_426,N_59);
nor U640 (N_640,In_702,N_453);
nor U641 (N_641,In_1331,In_1429);
nor U642 (N_642,N_597,In_349);
nand U643 (N_643,In_912,In_266);
nand U644 (N_644,In_1111,In_309);
nor U645 (N_645,In_1013,In_406);
nor U646 (N_646,N_492,N_586);
xor U647 (N_647,N_321,N_133);
or U648 (N_648,N_307,N_532);
nor U649 (N_649,In_298,In_558);
or U650 (N_650,In_1184,N_522);
nor U651 (N_651,N_583,N_493);
nand U652 (N_652,N_545,In_1218);
and U653 (N_653,In_376,N_381);
nand U654 (N_654,N_396,In_923);
and U655 (N_655,In_635,N_593);
xor U656 (N_656,N_571,In_1199);
nor U657 (N_657,In_322,In_114);
xnor U658 (N_658,N_575,N_199);
nand U659 (N_659,N_345,In_1153);
nand U660 (N_660,N_560,N_195);
nand U661 (N_661,N_395,N_116);
nand U662 (N_662,In_363,N_35);
xnor U663 (N_663,In_15,In_931);
xor U664 (N_664,In_838,In_1188);
nand U665 (N_665,N_44,N_537);
nor U666 (N_666,In_1148,N_500);
nand U667 (N_667,N_393,In_155);
nand U668 (N_668,N_525,N_98);
nand U669 (N_669,N_486,N_433);
and U670 (N_670,In_218,N_480);
xor U671 (N_671,N_106,N_374);
xnor U672 (N_672,N_168,In_623);
nand U673 (N_673,In_208,N_185);
and U674 (N_674,In_885,N_499);
xor U675 (N_675,N_114,In_446);
or U676 (N_676,N_323,In_586);
or U677 (N_677,N_566,In_497);
nand U678 (N_678,In_263,In_167);
and U679 (N_679,N_348,N_81);
nor U680 (N_680,N_508,In_1437);
and U681 (N_681,In_639,In_311);
or U682 (N_682,In_674,N_573);
xnor U683 (N_683,In_180,N_322);
nor U684 (N_684,N_549,N_340);
and U685 (N_685,N_420,In_1320);
xor U686 (N_686,N_73,In_688);
nor U687 (N_687,N_482,N_63);
nand U688 (N_688,In_135,In_1026);
and U689 (N_689,In_1450,In_534);
or U690 (N_690,N_352,In_1311);
nor U691 (N_691,In_1054,N_580);
xor U692 (N_692,N_558,In_1203);
and U693 (N_693,In_686,In_1453);
nand U694 (N_694,N_581,N_475);
or U695 (N_695,In_703,N_243);
and U696 (N_696,In_956,In_1446);
nor U697 (N_697,In_511,In_711);
xor U698 (N_698,In_1165,N_312);
nor U699 (N_699,In_793,N_189);
nor U700 (N_700,N_495,N_351);
or U701 (N_701,In_933,N_451);
nand U702 (N_702,In_1317,N_15);
or U703 (N_703,N_288,In_1162);
and U704 (N_704,In_547,N_544);
nor U705 (N_705,In_646,N_303);
nor U706 (N_706,N_113,In_1451);
xor U707 (N_707,N_318,In_1252);
and U708 (N_708,N_458,In_516);
xnor U709 (N_709,N_363,N_38);
xor U710 (N_710,In_1127,In_622);
nand U711 (N_711,N_300,In_264);
xor U712 (N_712,In_655,N_256);
xor U713 (N_713,In_280,In_802);
and U714 (N_714,N_510,In_158);
xnor U715 (N_715,N_452,In_126);
nand U716 (N_716,In_1394,N_314);
xnor U717 (N_717,N_58,In_559);
nor U718 (N_718,N_326,In_1419);
or U719 (N_719,N_437,N_404);
or U720 (N_720,In_491,N_405);
xnor U721 (N_721,N_328,In_640);
xnor U722 (N_722,In_1269,N_5);
nor U723 (N_723,N_186,N_526);
xor U724 (N_724,N_342,In_1177);
nor U725 (N_725,In_1348,In_1452);
nor U726 (N_726,In_1109,In_1283);
xor U727 (N_727,In_369,N_304);
and U728 (N_728,In_371,In_1324);
xor U729 (N_729,N_354,In_79);
nor U730 (N_730,N_39,In_1267);
nand U731 (N_731,In_955,In_1234);
xor U732 (N_732,N_334,N_401);
nand U733 (N_733,N_574,In_510);
nor U734 (N_734,In_1439,In_1245);
nor U735 (N_735,N_6,In_1025);
nor U736 (N_736,N_546,N_172);
or U737 (N_737,N_422,N_414);
or U738 (N_738,In_864,In_261);
and U739 (N_739,N_336,N_100);
nor U740 (N_740,In_572,In_318);
nor U741 (N_741,In_366,N_438);
nand U742 (N_742,N_490,N_2);
nand U743 (N_743,N_594,In_433);
or U744 (N_744,In_1354,In_345);
nor U745 (N_745,In_254,In_894);
or U746 (N_746,In_1459,In_157);
and U747 (N_747,N_585,In_1384);
nor U748 (N_748,In_1292,N_358);
nand U749 (N_749,N_568,N_48);
and U750 (N_750,In_890,In_524);
and U751 (N_751,In_1159,N_370);
xnor U752 (N_752,N_333,In_198);
or U753 (N_753,In_1260,N_212);
xnor U754 (N_754,In_1298,In_77);
xnor U755 (N_755,In_533,In_1472);
nand U756 (N_756,In_520,N_362);
or U757 (N_757,In_236,In_372);
and U758 (N_758,N_474,In_996);
and U759 (N_759,N_551,N_46);
and U760 (N_760,In_501,In_722);
and U761 (N_761,N_557,In_197);
or U762 (N_762,N_462,N_541);
xor U763 (N_763,N_208,N_385);
or U764 (N_764,N_191,In_581);
nor U765 (N_765,In_1062,N_316);
xor U766 (N_766,N_538,N_155);
xnor U767 (N_767,In_57,In_426);
xnor U768 (N_768,In_1174,N_491);
or U769 (N_769,N_435,In_1414);
nand U770 (N_770,N_501,In_752);
xnor U771 (N_771,In_356,N_273);
nor U772 (N_772,In_742,N_317);
nor U773 (N_773,N_124,N_507);
xnor U774 (N_774,In_282,In_675);
nor U775 (N_775,In_256,In_1308);
or U776 (N_776,N_238,In_1116);
and U777 (N_777,In_696,In_695);
nand U778 (N_778,In_677,N_485);
nand U779 (N_779,In_1117,In_45);
or U780 (N_780,In_1397,N_268);
and U781 (N_781,In_405,N_520);
or U782 (N_782,In_1469,In_1131);
nor U783 (N_783,N_456,In_801);
nor U784 (N_784,N_13,N_487);
or U785 (N_785,In_187,N_72);
nand U786 (N_786,In_450,N_154);
nand U787 (N_787,In_977,In_617);
and U788 (N_788,In_287,N_391);
xnor U789 (N_789,In_191,N_443);
or U790 (N_790,N_524,N_330);
and U791 (N_791,In_378,N_309);
xor U792 (N_792,In_278,In_1241);
xor U793 (N_793,N_161,In_1040);
or U794 (N_794,In_147,In_1352);
nor U795 (N_795,In_721,N_591);
nor U796 (N_796,N_335,In_689);
nand U797 (N_797,N_346,N_173);
and U798 (N_798,N_552,N_298);
xor U799 (N_799,In_518,In_296);
and U800 (N_800,In_1417,In_1097);
xnor U801 (N_801,N_450,N_494);
nor U802 (N_802,In_758,In_1237);
nand U803 (N_803,N_576,In_726);
or U804 (N_804,N_128,N_563);
nor U805 (N_805,In_97,In_1028);
or U806 (N_806,In_636,N_353);
or U807 (N_807,In_984,N_324);
xnor U808 (N_808,N_247,In_942);
xor U809 (N_809,In_916,N_37);
nor U810 (N_810,N_588,N_361);
nand U811 (N_811,In_1356,In_725);
or U812 (N_812,In_429,N_169);
nor U813 (N_813,N_0,N_7);
nand U814 (N_814,N_139,In_592);
nand U815 (N_815,N_104,In_870);
and U816 (N_816,N_220,N_112);
nand U817 (N_817,In_176,N_177);
and U818 (N_818,In_395,N_505);
nor U819 (N_819,In_159,In_1210);
nor U820 (N_820,In_459,N_431);
and U821 (N_821,N_511,N_444);
xnor U822 (N_822,N_394,N_380);
xor U823 (N_823,N_239,In_1339);
or U824 (N_824,In_595,In_30);
or U825 (N_825,N_424,In_149);
xnor U826 (N_826,N_530,N_89);
nor U827 (N_827,N_347,In_1460);
nand U828 (N_828,N_378,In_913);
nor U829 (N_829,In_350,N_130);
nand U830 (N_830,N_79,N_339);
nor U831 (N_831,N_223,N_306);
nand U832 (N_832,N_134,N_313);
nand U833 (N_833,N_43,N_222);
nand U834 (N_834,In_884,In_1428);
nor U835 (N_835,N_471,In_370);
and U836 (N_836,In_379,In_1369);
nand U837 (N_837,N_277,In_274);
nand U838 (N_838,N_400,In_892);
nand U839 (N_839,In_245,In_217);
xnor U840 (N_840,In_226,In_1337);
nor U841 (N_841,In_343,In_1401);
nor U842 (N_842,In_1082,In_1192);
or U843 (N_843,N_596,In_17);
and U844 (N_844,In_1441,N_311);
and U845 (N_845,In_92,N_373);
nand U846 (N_846,N_127,In_1467);
xor U847 (N_847,In_353,N_77);
xor U848 (N_848,In_182,In_869);
nand U849 (N_849,N_428,N_398);
nand U850 (N_850,In_751,In_779);
nand U851 (N_851,N_87,N_383);
and U852 (N_852,N_94,In_184);
or U853 (N_853,N_62,N_241);
nand U854 (N_854,In_728,N_506);
nand U855 (N_855,In_425,In_652);
or U856 (N_856,N_329,N_371);
or U857 (N_857,In_479,N_402);
and U858 (N_858,N_479,N_467);
nand U859 (N_859,In_780,In_648);
or U860 (N_860,In_304,In_373);
and U861 (N_861,N_368,N_164);
and U862 (N_862,In_770,N_390);
xor U863 (N_863,N_282,In_416);
nand U864 (N_864,In_1373,In_1496);
or U865 (N_865,N_496,N_299);
or U866 (N_866,In_1455,In_1349);
or U867 (N_867,In_1007,N_349);
nor U868 (N_868,In_342,In_1196);
and U869 (N_869,N_136,N_464);
and U870 (N_870,N_441,In_387);
and U871 (N_871,N_249,N_561);
nand U872 (N_872,In_1479,In_1249);
xnor U873 (N_873,N_488,In_1033);
or U874 (N_874,In_1294,N_512);
nor U875 (N_875,N_290,N_430);
or U876 (N_876,In_0,N_289);
or U877 (N_877,N_449,In_1392);
or U878 (N_878,In_1220,N_463);
or U879 (N_879,In_16,N_421);
or U880 (N_880,N_562,N_469);
nor U881 (N_881,In_749,N_210);
xnor U882 (N_882,N_434,In_849);
or U883 (N_883,In_1391,N_158);
and U884 (N_884,In_1410,N_376);
nand U885 (N_885,In_91,In_947);
nand U886 (N_886,N_248,In_431);
nand U887 (N_887,In_393,In_361);
xor U888 (N_888,N_80,N_367);
nor U889 (N_889,N_71,N_514);
nand U890 (N_890,In_1411,N_343);
nand U891 (N_891,In_1438,In_1008);
and U892 (N_892,N_556,In_1009);
nand U893 (N_893,In_957,In_986);
nand U894 (N_894,In_699,In_335);
xnor U895 (N_895,In_988,In_1015);
xor U896 (N_896,N_460,N_149);
or U897 (N_897,N_569,N_448);
and U898 (N_898,N_216,In_1290);
xor U899 (N_899,In_848,In_210);
and U900 (N_900,N_375,N_833);
or U901 (N_901,N_618,In_618);
nand U902 (N_902,In_775,N_869);
nor U903 (N_903,In_951,In_574);
or U904 (N_904,N_54,In_904);
xor U905 (N_905,In_1154,N_635);
xor U906 (N_906,In_1482,N_847);
or U907 (N_907,N_773,N_392);
nand U908 (N_908,In_339,N_748);
nor U909 (N_909,N_723,N_694);
and U910 (N_910,N_827,In_1287);
nor U911 (N_911,N_706,N_365);
nand U912 (N_912,In_519,In_64);
xor U913 (N_913,N_366,N_319);
and U914 (N_914,In_466,N_344);
and U915 (N_915,N_240,N_631);
nor U916 (N_916,In_1360,In_1366);
nand U917 (N_917,N_301,N_846);
and U918 (N_918,N_427,N_663);
nand U919 (N_919,N_820,N_899);
xnor U920 (N_920,N_855,N_497);
xnor U921 (N_921,N_689,In_1023);
xor U922 (N_922,In_462,N_774);
xor U923 (N_923,In_104,In_633);
and U924 (N_924,N_350,N_799);
and U925 (N_925,N_652,N_610);
nand U926 (N_926,In_1274,In_1078);
or U927 (N_927,N_473,N_805);
nand U928 (N_928,N_701,In_103);
xor U929 (N_929,N_616,N_605);
nand U930 (N_930,In_813,In_72);
xnor U931 (N_931,N_372,N_729);
and U932 (N_932,N_856,In_969);
and U933 (N_933,N_800,N_873);
and U934 (N_934,N_388,N_477);
nand U935 (N_935,In_535,N_582);
nor U936 (N_936,N_879,N_611);
and U937 (N_937,N_627,N_513);
nand U938 (N_938,In_448,In_958);
nand U939 (N_939,N_658,N_459);
or U940 (N_940,N_308,N_531);
xnor U941 (N_941,N_685,N_720);
nand U942 (N_942,N_664,N_457);
xor U943 (N_943,N_178,N_466);
and U944 (N_944,N_82,N_291);
xor U945 (N_945,N_656,In_1434);
and U946 (N_946,N_684,N_564);
nor U947 (N_947,N_741,N_204);
and U948 (N_948,N_896,In_1321);
nor U949 (N_949,N_698,N_721);
xor U950 (N_950,N_782,N_699);
xnor U951 (N_951,N_535,N_766);
nor U952 (N_952,N_408,N_521);
xnor U953 (N_953,N_707,N_752);
or U954 (N_954,N_406,N_40);
and U955 (N_955,N_796,N_875);
nand U956 (N_956,In_1375,N_878);
xnor U957 (N_957,N_484,N_604);
or U958 (N_958,N_798,N_767);
xnor U959 (N_959,In_773,N_355);
and U960 (N_960,In_1022,In_939);
and U961 (N_961,In_1038,N_835);
nor U962 (N_962,In_941,N_650);
nor U963 (N_963,In_1423,N_677);
xnor U964 (N_964,N_623,N_751);
or U965 (N_965,N_651,In_990);
nor U966 (N_966,N_825,N_716);
xor U967 (N_967,N_379,N_753);
xor U968 (N_968,In_463,N_636);
or U969 (N_969,N_893,N_808);
or U970 (N_970,In_329,N_356);
or U971 (N_971,N_703,N_612);
nand U972 (N_972,N_889,N_157);
xor U973 (N_973,In_475,N_803);
nor U974 (N_974,N_647,N_862);
nand U975 (N_975,N_834,N_425);
and U976 (N_976,N_125,N_822);
and U977 (N_977,N_877,In_81);
or U978 (N_978,N_678,N_600);
nand U979 (N_979,N_174,N_676);
or U980 (N_980,N_870,N_821);
xor U981 (N_981,In_455,N_857);
nor U982 (N_982,N_897,In_539);
and U983 (N_983,N_813,In_954);
and U984 (N_984,N_811,N_439);
or U985 (N_985,N_771,N_882);
nor U986 (N_986,N_853,N_446);
xor U987 (N_987,N_843,N_34);
or U988 (N_988,In_630,N_554);
and U989 (N_989,N_887,N_332);
nor U990 (N_990,N_683,N_785);
and U991 (N_991,N_674,N_331);
or U992 (N_992,N_746,N_634);
xnor U993 (N_993,N_814,N_690);
and U994 (N_994,N_572,N_655);
and U995 (N_995,N_577,N_754);
and U996 (N_996,N_33,In_277);
xor U997 (N_997,N_787,N_788);
and U998 (N_998,In_1186,In_601);
or U999 (N_999,N_679,N_147);
or U1000 (N_1000,N_881,N_775);
nor U1001 (N_1001,In_333,N_640);
nor U1002 (N_1002,N_776,N_143);
xor U1003 (N_1003,N_763,N_602);
xnor U1004 (N_1004,In_1121,N_772);
or U1005 (N_1005,In_929,N_625);
nor U1006 (N_1006,N_769,In_669);
xnor U1007 (N_1007,N_359,N_761);
and U1008 (N_1008,N_51,N_620);
and U1009 (N_1009,N_688,N_804);
and U1010 (N_1010,N_137,N_708);
xnor U1011 (N_1011,N_653,In_761);
nand U1012 (N_1012,N_760,N_432);
nor U1013 (N_1013,N_152,In_1338);
nand U1014 (N_1014,N_540,N_693);
nor U1015 (N_1015,In_681,In_1244);
nor U1016 (N_1016,N_780,N_675);
nand U1017 (N_1017,In_399,In_194);
and U1018 (N_1018,N_750,In_428);
and U1019 (N_1019,N_884,N_714);
and U1020 (N_1020,N_504,In_1376);
nand U1021 (N_1021,In_987,N_727);
or U1022 (N_1022,In_212,N_712);
nor U1023 (N_1023,N_736,N_461);
xnor U1024 (N_1024,N_858,N_830);
nor U1025 (N_1025,N_744,N_436);
nand U1026 (N_1026,N_883,N_603);
xnor U1027 (N_1027,N_517,N_615);
or U1028 (N_1028,In_1255,In_1370);
or U1029 (N_1029,In_642,In_204);
nand U1030 (N_1030,N_734,In_27);
nand U1031 (N_1031,N_747,N_885);
xnor U1032 (N_1032,N_608,N_280);
xor U1033 (N_1033,N_824,N_691);
xnor U1034 (N_1034,In_76,N_742);
and U1035 (N_1035,N_542,N_76);
or U1036 (N_1036,N_692,N_888);
nand U1037 (N_1037,N_624,In_1095);
or U1038 (N_1038,N_726,N_733);
nand U1039 (N_1039,N_527,In_712);
and U1040 (N_1040,N_868,In_1168);
or U1041 (N_1041,N_735,In_87);
and U1042 (N_1042,In_336,N_302);
or U1043 (N_1043,N_768,In_891);
nor U1044 (N_1044,N_863,N_781);
nor U1045 (N_1045,N_836,N_892);
nand U1046 (N_1046,N_648,N_377);
nand U1047 (N_1047,N_749,N_840);
or U1048 (N_1048,N_702,N_387);
and U1049 (N_1049,In_772,In_1142);
or U1050 (N_1050,N_871,In_1052);
and U1051 (N_1051,N_613,N_646);
nor U1052 (N_1052,N_806,N_369);
and U1053 (N_1053,N_719,N_419);
nor U1054 (N_1054,In_153,N_170);
or U1055 (N_1055,In_1137,In_972);
and U1056 (N_1056,N_666,N_724);
or U1057 (N_1057,N_682,N_167);
nor U1058 (N_1058,In_1208,N_440);
nor U1059 (N_1059,In_259,N_765);
xor U1060 (N_1060,N_864,N_201);
and U1061 (N_1061,N_794,N_412);
xnor U1062 (N_1062,N_725,N_668);
and U1063 (N_1063,N_790,N_659);
xor U1064 (N_1064,In_530,N_534);
and U1065 (N_1065,N_645,N_849);
nor U1066 (N_1066,N_739,N_284);
and U1067 (N_1067,N_609,N_140);
nand U1068 (N_1068,N_687,N_415);
or U1069 (N_1069,N_786,N_764);
or U1070 (N_1070,N_795,In_766);
xor U1071 (N_1071,N_103,N_880);
nand U1072 (N_1072,N_730,N_801);
nor U1073 (N_1073,N_628,In_1092);
xnor U1074 (N_1074,In_792,N_416);
xor U1075 (N_1075,In_684,N_837);
or U1076 (N_1076,N_529,In_427);
xnor U1077 (N_1077,N_472,N_587);
or U1078 (N_1078,N_823,N_812);
nand U1079 (N_1079,In_242,N_632);
or U1080 (N_1080,N_890,N_783);
xor U1081 (N_1081,N_874,In_875);
or U1082 (N_1082,In_1047,N_271);
and U1083 (N_1083,N_279,N_662);
and U1084 (N_1084,N_553,N_657);
and U1085 (N_1085,In_290,N_644);
and U1086 (N_1086,In_1398,In_1332);
nand U1087 (N_1087,N_543,In_360);
and U1088 (N_1088,In_687,N_815);
nand U1089 (N_1089,In_948,N_797);
or U1090 (N_1090,N_671,N_601);
nor U1091 (N_1091,N_757,N_876);
and U1092 (N_1092,N_630,N_789);
and U1093 (N_1093,N_851,In_607);
or U1094 (N_1094,In_238,In_215);
or U1095 (N_1095,In_443,N_642);
and U1096 (N_1096,N_891,N_850);
and U1097 (N_1097,N_429,N_845);
nand U1098 (N_1098,N_793,N_841);
or U1099 (N_1099,N_423,N_397);
nand U1100 (N_1100,N_590,N_203);
nand U1101 (N_1101,In_205,N_697);
or U1102 (N_1102,N_516,N_384);
xor U1103 (N_1103,N_196,N_818);
xnor U1104 (N_1104,N_859,In_118);
and U1105 (N_1105,In_867,N_629);
or U1106 (N_1106,N_364,N_338);
xnor U1107 (N_1107,In_896,In_653);
or U1108 (N_1108,N_740,N_599);
nor U1109 (N_1109,N_672,N_502);
or U1110 (N_1110,In_1228,N_320);
and U1111 (N_1111,N_713,N_842);
nand U1112 (N_1112,N_327,N_465);
nor U1113 (N_1113,In_33,N_898);
nor U1114 (N_1114,N_831,N_738);
nand U1115 (N_1115,In_246,N_872);
or U1116 (N_1116,N_528,N_802);
or U1117 (N_1117,N_643,N_894);
nand U1118 (N_1118,N_584,N_90);
or U1119 (N_1119,N_180,In_1183);
or U1120 (N_1120,In_47,In_738);
nor U1121 (N_1121,N_886,N_709);
xor U1122 (N_1122,N_325,N_498);
nand U1123 (N_1123,In_415,N_110);
xor U1124 (N_1124,N_732,N_695);
nand U1125 (N_1125,N_728,In_1179);
nor U1126 (N_1126,N_861,N_826);
nor U1127 (N_1127,N_156,N_413);
nor U1128 (N_1128,N_641,In_625);
or U1129 (N_1129,N_399,N_829);
nor U1130 (N_1130,N_866,In_11);
nand U1131 (N_1131,N_567,N_606);
or U1132 (N_1132,N_84,N_686);
and U1133 (N_1133,N_410,N_895);
or U1134 (N_1134,N_68,N_854);
nor U1135 (N_1135,N_578,In_134);
or U1136 (N_1136,N_622,N_489);
and U1137 (N_1137,N_209,N_639);
xor U1138 (N_1138,N_120,N_743);
xnor U1139 (N_1139,N_715,In_1329);
nand U1140 (N_1140,In_1155,In_1307);
nand U1141 (N_1141,N_633,N_770);
xnor U1142 (N_1142,N_722,N_570);
xnor U1143 (N_1143,N_654,N_468);
xor U1144 (N_1144,In_794,N_621);
or U1145 (N_1145,N_816,N_17);
nor U1146 (N_1146,N_848,In_358);
and U1147 (N_1147,N_660,N_759);
or U1148 (N_1148,N_619,N_589);
and U1149 (N_1149,N_661,N_681);
nor U1150 (N_1150,N_758,N_16);
xnor U1151 (N_1151,N_61,N_360);
and U1152 (N_1152,N_592,N_126);
xnor U1153 (N_1153,In_1480,N_417);
xnor U1154 (N_1154,N_731,N_231);
nor U1155 (N_1155,N_190,N_673);
and U1156 (N_1156,In_1364,N_224);
and U1157 (N_1157,N_670,In_782);
or U1158 (N_1158,In_1265,N_555);
or U1159 (N_1159,N_844,N_20);
nor U1160 (N_1160,N_476,In_461);
and U1161 (N_1161,In_308,N_819);
and U1162 (N_1162,N_778,N_315);
nor U1163 (N_1163,N_852,N_696);
or U1164 (N_1164,N_810,N_860);
nor U1165 (N_1165,N_536,N_614);
xor U1166 (N_1166,N_777,N_617);
nor U1167 (N_1167,N_382,N_626);
and U1168 (N_1168,N_595,N_547);
and U1169 (N_1169,N_737,N_523);
nor U1170 (N_1170,N_711,N_680);
and U1171 (N_1171,N_550,N_838);
nand U1172 (N_1172,N_607,N_839);
nand U1173 (N_1173,N_700,In_1258);
and U1174 (N_1174,N_442,N_762);
or U1175 (N_1175,In_1473,N_455);
nor U1176 (N_1176,N_272,N_357);
nor U1177 (N_1177,In_1306,N_710);
xor U1178 (N_1178,In_348,N_704);
nand U1179 (N_1179,N_745,N_667);
nor U1180 (N_1180,N_756,N_717);
xor U1181 (N_1181,N_559,N_649);
nand U1182 (N_1182,N_533,In_1488);
or U1183 (N_1183,N_755,N_418);
xor U1184 (N_1184,N_832,In_1106);
xor U1185 (N_1185,N_669,N_187);
and U1186 (N_1186,In_1330,In_541);
nor U1187 (N_1187,N_817,N_779);
and U1188 (N_1188,N_519,N_638);
nand U1189 (N_1189,N_665,N_705);
xnor U1190 (N_1190,N_598,N_718);
or U1191 (N_1191,N_828,N_867);
xor U1192 (N_1192,In_691,N_865);
and U1193 (N_1193,N_807,In_484);
or U1194 (N_1194,N_454,N_792);
nor U1195 (N_1195,N_637,In_276);
xor U1196 (N_1196,N_809,In_908);
nand U1197 (N_1197,N_565,In_1156);
nand U1198 (N_1198,N_784,N_518);
and U1199 (N_1199,N_483,N_791);
nor U1200 (N_1200,N_1177,N_1162);
nor U1201 (N_1201,N_1073,N_1039);
or U1202 (N_1202,N_994,N_929);
nor U1203 (N_1203,N_953,N_905);
xor U1204 (N_1204,N_1129,N_1182);
xnor U1205 (N_1205,N_1130,N_987);
and U1206 (N_1206,N_982,N_937);
nand U1207 (N_1207,N_1197,N_1150);
xnor U1208 (N_1208,N_909,N_1169);
nand U1209 (N_1209,N_1155,N_972);
or U1210 (N_1210,N_1071,N_1018);
or U1211 (N_1211,N_959,N_1136);
xor U1212 (N_1212,N_1013,N_1151);
xnor U1213 (N_1213,N_983,N_1029);
xnor U1214 (N_1214,N_936,N_1153);
nand U1215 (N_1215,N_1126,N_1066);
xor U1216 (N_1216,N_1164,N_1188);
xor U1217 (N_1217,N_1015,N_1068);
nor U1218 (N_1218,N_971,N_1009);
and U1219 (N_1219,N_1053,N_1120);
nand U1220 (N_1220,N_1091,N_1141);
nand U1221 (N_1221,N_927,N_1063);
xor U1222 (N_1222,N_1006,N_949);
and U1223 (N_1223,N_1149,N_1152);
and U1224 (N_1224,N_1156,N_1125);
or U1225 (N_1225,N_1193,N_911);
or U1226 (N_1226,N_914,N_1195);
xnor U1227 (N_1227,N_919,N_1139);
nand U1228 (N_1228,N_989,N_1027);
and U1229 (N_1229,N_1191,N_944);
and U1230 (N_1230,N_1167,N_1166);
nor U1231 (N_1231,N_1049,N_1019);
or U1232 (N_1232,N_915,N_996);
nor U1233 (N_1233,N_1183,N_1023);
and U1234 (N_1234,N_1030,N_1113);
or U1235 (N_1235,N_1056,N_1154);
or U1236 (N_1236,N_1020,N_1144);
nand U1237 (N_1237,N_1135,N_1158);
nand U1238 (N_1238,N_1021,N_1034);
or U1239 (N_1239,N_951,N_907);
or U1240 (N_1240,N_1111,N_1110);
or U1241 (N_1241,N_1100,N_984);
or U1242 (N_1242,N_1025,N_1106);
or U1243 (N_1243,N_1122,N_1143);
or U1244 (N_1244,N_1165,N_903);
nor U1245 (N_1245,N_1184,N_1000);
or U1246 (N_1246,N_956,N_1115);
or U1247 (N_1247,N_1086,N_1033);
or U1248 (N_1248,N_910,N_1124);
nor U1249 (N_1249,N_1088,N_999);
and U1250 (N_1250,N_1112,N_1052);
xnor U1251 (N_1251,N_1105,N_1163);
xnor U1252 (N_1252,N_1060,N_908);
nor U1253 (N_1253,N_928,N_942);
nor U1254 (N_1254,N_1083,N_1186);
nor U1255 (N_1255,N_931,N_993);
nand U1256 (N_1256,N_1131,N_1045);
and U1257 (N_1257,N_1132,N_997);
nand U1258 (N_1258,N_922,N_1035);
xnor U1259 (N_1259,N_1107,N_1148);
nand U1260 (N_1260,N_1160,N_976);
or U1261 (N_1261,N_1116,N_990);
nor U1262 (N_1262,N_961,N_955);
and U1263 (N_1263,N_1007,N_1147);
and U1264 (N_1264,N_945,N_1189);
or U1265 (N_1265,N_1192,N_1161);
xor U1266 (N_1266,N_900,N_1024);
nand U1267 (N_1267,N_1114,N_995);
xnor U1268 (N_1268,N_935,N_1017);
and U1269 (N_1269,N_1048,N_958);
nor U1270 (N_1270,N_1128,N_943);
and U1271 (N_1271,N_998,N_1046);
xnor U1272 (N_1272,N_1079,N_933);
xor U1273 (N_1273,N_1065,N_979);
or U1274 (N_1274,N_902,N_1095);
nand U1275 (N_1275,N_988,N_924);
or U1276 (N_1276,N_1179,N_977);
nor U1277 (N_1277,N_1103,N_1181);
xnor U1278 (N_1278,N_917,N_1174);
xor U1279 (N_1279,N_934,N_1059);
nand U1280 (N_1280,N_1187,N_1199);
nand U1281 (N_1281,N_1085,N_1074);
or U1282 (N_1282,N_1061,N_1051);
nand U1283 (N_1283,N_1118,N_1084);
or U1284 (N_1284,N_975,N_916);
or U1285 (N_1285,N_1028,N_1062);
nor U1286 (N_1286,N_1138,N_967);
or U1287 (N_1287,N_1078,N_1043);
nor U1288 (N_1288,N_1008,N_1022);
nand U1289 (N_1289,N_1031,N_1157);
or U1290 (N_1290,N_1093,N_1026);
or U1291 (N_1291,N_1185,N_1064);
or U1292 (N_1292,N_1011,N_1082);
or U1293 (N_1293,N_1102,N_1170);
and U1294 (N_1294,N_1109,N_938);
xor U1295 (N_1295,N_970,N_1140);
nor U1296 (N_1296,N_1173,N_962);
or U1297 (N_1297,N_913,N_1090);
nand U1298 (N_1298,N_1094,N_1058);
xnor U1299 (N_1299,N_1054,N_1080);
nor U1300 (N_1300,N_1005,N_1010);
xor U1301 (N_1301,N_1198,N_960);
or U1302 (N_1302,N_1196,N_923);
and U1303 (N_1303,N_904,N_1087);
and U1304 (N_1304,N_965,N_991);
and U1305 (N_1305,N_930,N_954);
and U1306 (N_1306,N_992,N_1108);
or U1307 (N_1307,N_939,N_1190);
xor U1308 (N_1308,N_1044,N_1075);
nor U1309 (N_1309,N_1145,N_1146);
nand U1310 (N_1310,N_1003,N_1098);
nor U1311 (N_1311,N_1077,N_946);
nor U1312 (N_1312,N_1004,N_1101);
nor U1313 (N_1313,N_947,N_1014);
nand U1314 (N_1314,N_1172,N_1099);
or U1315 (N_1315,N_1038,N_1089);
and U1316 (N_1316,N_966,N_1121);
xor U1317 (N_1317,N_1097,N_921);
nor U1318 (N_1318,N_1040,N_950);
xor U1319 (N_1319,N_980,N_1036);
nand U1320 (N_1320,N_1134,N_1123);
or U1321 (N_1321,N_974,N_1137);
or U1322 (N_1322,N_948,N_901);
xor U1323 (N_1323,N_986,N_1117);
nor U1324 (N_1324,N_985,N_973);
and U1325 (N_1325,N_1175,N_1055);
nor U1326 (N_1326,N_1032,N_912);
nor U1327 (N_1327,N_957,N_920);
xor U1328 (N_1328,N_1041,N_1133);
xor U1329 (N_1329,N_1127,N_906);
xnor U1330 (N_1330,N_1070,N_978);
xnor U1331 (N_1331,N_969,N_1096);
nand U1332 (N_1332,N_940,N_1076);
and U1333 (N_1333,N_964,N_932);
xnor U1334 (N_1334,N_1180,N_1057);
and U1335 (N_1335,N_1159,N_1072);
or U1336 (N_1336,N_1050,N_1119);
xnor U1337 (N_1337,N_1168,N_1069);
nand U1338 (N_1338,N_981,N_1081);
nand U1339 (N_1339,N_1037,N_1067);
xor U1340 (N_1340,N_963,N_968);
and U1341 (N_1341,N_925,N_1092);
xnor U1342 (N_1342,N_1142,N_1012);
and U1343 (N_1343,N_1104,N_926);
and U1344 (N_1344,N_1001,N_1178);
and U1345 (N_1345,N_952,N_1002);
and U1346 (N_1346,N_941,N_1171);
xnor U1347 (N_1347,N_1016,N_1042);
or U1348 (N_1348,N_1047,N_1194);
xnor U1349 (N_1349,N_1176,N_918);
xor U1350 (N_1350,N_986,N_1199);
nor U1351 (N_1351,N_1031,N_1092);
nand U1352 (N_1352,N_957,N_1092);
nor U1353 (N_1353,N_1119,N_1152);
and U1354 (N_1354,N_1143,N_1145);
and U1355 (N_1355,N_936,N_940);
or U1356 (N_1356,N_1022,N_1127);
nand U1357 (N_1357,N_900,N_902);
and U1358 (N_1358,N_1187,N_944);
nand U1359 (N_1359,N_1043,N_1012);
nand U1360 (N_1360,N_971,N_1110);
nor U1361 (N_1361,N_981,N_1109);
nand U1362 (N_1362,N_1080,N_1172);
nor U1363 (N_1363,N_1033,N_1010);
nor U1364 (N_1364,N_1161,N_998);
or U1365 (N_1365,N_1005,N_938);
nand U1366 (N_1366,N_919,N_1150);
and U1367 (N_1367,N_1101,N_1112);
nor U1368 (N_1368,N_1182,N_1064);
nand U1369 (N_1369,N_1010,N_1064);
nand U1370 (N_1370,N_998,N_957);
xnor U1371 (N_1371,N_1099,N_1104);
xor U1372 (N_1372,N_938,N_995);
and U1373 (N_1373,N_975,N_1000);
xnor U1374 (N_1374,N_1189,N_1078);
nand U1375 (N_1375,N_912,N_905);
nand U1376 (N_1376,N_1067,N_1145);
nand U1377 (N_1377,N_952,N_1077);
and U1378 (N_1378,N_918,N_1080);
xnor U1379 (N_1379,N_1130,N_969);
and U1380 (N_1380,N_1041,N_990);
and U1381 (N_1381,N_962,N_952);
and U1382 (N_1382,N_936,N_1143);
xnor U1383 (N_1383,N_973,N_991);
nor U1384 (N_1384,N_1084,N_905);
or U1385 (N_1385,N_1155,N_1171);
or U1386 (N_1386,N_1060,N_994);
and U1387 (N_1387,N_1038,N_906);
xor U1388 (N_1388,N_1120,N_1198);
xor U1389 (N_1389,N_940,N_1145);
or U1390 (N_1390,N_1082,N_1102);
xor U1391 (N_1391,N_1128,N_1161);
nor U1392 (N_1392,N_1023,N_1055);
nor U1393 (N_1393,N_924,N_1080);
nand U1394 (N_1394,N_950,N_1119);
nor U1395 (N_1395,N_1199,N_911);
nor U1396 (N_1396,N_1021,N_1083);
and U1397 (N_1397,N_1167,N_919);
and U1398 (N_1398,N_1132,N_1188);
nor U1399 (N_1399,N_1072,N_911);
nor U1400 (N_1400,N_1059,N_993);
and U1401 (N_1401,N_973,N_997);
or U1402 (N_1402,N_1079,N_1192);
and U1403 (N_1403,N_1027,N_958);
nor U1404 (N_1404,N_932,N_1057);
or U1405 (N_1405,N_1059,N_995);
xnor U1406 (N_1406,N_1020,N_1087);
and U1407 (N_1407,N_1162,N_1139);
and U1408 (N_1408,N_1016,N_1048);
and U1409 (N_1409,N_932,N_1128);
nand U1410 (N_1410,N_1109,N_1041);
nor U1411 (N_1411,N_1081,N_1057);
xnor U1412 (N_1412,N_1147,N_1010);
nand U1413 (N_1413,N_939,N_1133);
nor U1414 (N_1414,N_1043,N_1087);
nor U1415 (N_1415,N_1169,N_1072);
nand U1416 (N_1416,N_921,N_1094);
nand U1417 (N_1417,N_1105,N_953);
nor U1418 (N_1418,N_1185,N_1055);
nand U1419 (N_1419,N_942,N_1176);
xor U1420 (N_1420,N_1144,N_1065);
nor U1421 (N_1421,N_1052,N_1102);
or U1422 (N_1422,N_1146,N_1037);
or U1423 (N_1423,N_920,N_1146);
xor U1424 (N_1424,N_1129,N_1033);
nand U1425 (N_1425,N_1010,N_1139);
nand U1426 (N_1426,N_1198,N_1071);
xor U1427 (N_1427,N_1026,N_1016);
nand U1428 (N_1428,N_957,N_1002);
or U1429 (N_1429,N_1165,N_927);
nand U1430 (N_1430,N_1156,N_1151);
xor U1431 (N_1431,N_967,N_1051);
xnor U1432 (N_1432,N_1178,N_986);
or U1433 (N_1433,N_989,N_934);
xnor U1434 (N_1434,N_1059,N_1029);
xor U1435 (N_1435,N_1007,N_1173);
and U1436 (N_1436,N_1198,N_963);
nand U1437 (N_1437,N_1184,N_1087);
or U1438 (N_1438,N_980,N_1019);
or U1439 (N_1439,N_992,N_1077);
or U1440 (N_1440,N_1194,N_914);
xnor U1441 (N_1441,N_1077,N_1140);
and U1442 (N_1442,N_1165,N_972);
nand U1443 (N_1443,N_1161,N_1180);
nand U1444 (N_1444,N_1103,N_1164);
and U1445 (N_1445,N_1083,N_1079);
xnor U1446 (N_1446,N_978,N_941);
xnor U1447 (N_1447,N_1052,N_946);
nand U1448 (N_1448,N_1121,N_1116);
and U1449 (N_1449,N_944,N_1164);
xor U1450 (N_1450,N_938,N_969);
nor U1451 (N_1451,N_997,N_1072);
and U1452 (N_1452,N_968,N_1161);
or U1453 (N_1453,N_973,N_953);
or U1454 (N_1454,N_929,N_1160);
xnor U1455 (N_1455,N_902,N_976);
nand U1456 (N_1456,N_1043,N_1161);
and U1457 (N_1457,N_927,N_1152);
xor U1458 (N_1458,N_1192,N_1193);
nor U1459 (N_1459,N_941,N_1105);
and U1460 (N_1460,N_943,N_1065);
or U1461 (N_1461,N_958,N_1102);
nor U1462 (N_1462,N_1176,N_1030);
xnor U1463 (N_1463,N_950,N_1051);
xor U1464 (N_1464,N_1087,N_1159);
or U1465 (N_1465,N_992,N_923);
or U1466 (N_1466,N_1132,N_926);
nor U1467 (N_1467,N_1065,N_1187);
and U1468 (N_1468,N_1192,N_1119);
nor U1469 (N_1469,N_988,N_1164);
or U1470 (N_1470,N_985,N_957);
nor U1471 (N_1471,N_995,N_1019);
and U1472 (N_1472,N_1133,N_908);
nand U1473 (N_1473,N_937,N_1027);
nand U1474 (N_1474,N_1158,N_1016);
or U1475 (N_1475,N_1178,N_1110);
nor U1476 (N_1476,N_1043,N_1154);
xnor U1477 (N_1477,N_962,N_1054);
or U1478 (N_1478,N_920,N_990);
or U1479 (N_1479,N_1110,N_1170);
and U1480 (N_1480,N_1092,N_988);
nand U1481 (N_1481,N_1163,N_1193);
nor U1482 (N_1482,N_1046,N_910);
xor U1483 (N_1483,N_964,N_1078);
nand U1484 (N_1484,N_974,N_993);
xnor U1485 (N_1485,N_1075,N_1143);
or U1486 (N_1486,N_1165,N_950);
nor U1487 (N_1487,N_1025,N_1133);
and U1488 (N_1488,N_1032,N_1193);
xor U1489 (N_1489,N_974,N_1082);
nand U1490 (N_1490,N_1103,N_982);
and U1491 (N_1491,N_977,N_1019);
nand U1492 (N_1492,N_1054,N_1032);
xnor U1493 (N_1493,N_939,N_942);
and U1494 (N_1494,N_1110,N_1188);
xor U1495 (N_1495,N_983,N_1065);
xor U1496 (N_1496,N_1079,N_1159);
or U1497 (N_1497,N_942,N_1023);
or U1498 (N_1498,N_1105,N_1182);
and U1499 (N_1499,N_967,N_1028);
nand U1500 (N_1500,N_1467,N_1284);
xnor U1501 (N_1501,N_1477,N_1327);
nor U1502 (N_1502,N_1275,N_1436);
xor U1503 (N_1503,N_1261,N_1285);
and U1504 (N_1504,N_1482,N_1274);
and U1505 (N_1505,N_1226,N_1282);
nor U1506 (N_1506,N_1295,N_1200);
and U1507 (N_1507,N_1369,N_1379);
nand U1508 (N_1508,N_1344,N_1389);
and U1509 (N_1509,N_1277,N_1471);
and U1510 (N_1510,N_1245,N_1462);
or U1511 (N_1511,N_1264,N_1307);
nor U1512 (N_1512,N_1268,N_1396);
and U1513 (N_1513,N_1425,N_1298);
nand U1514 (N_1514,N_1331,N_1405);
nor U1515 (N_1515,N_1406,N_1221);
or U1516 (N_1516,N_1337,N_1392);
xor U1517 (N_1517,N_1438,N_1452);
or U1518 (N_1518,N_1232,N_1423);
nor U1519 (N_1519,N_1347,N_1278);
or U1520 (N_1520,N_1464,N_1293);
nand U1521 (N_1521,N_1316,N_1237);
nand U1522 (N_1522,N_1215,N_1465);
and U1523 (N_1523,N_1470,N_1361);
xnor U1524 (N_1524,N_1483,N_1400);
or U1525 (N_1525,N_1312,N_1283);
and U1526 (N_1526,N_1244,N_1443);
and U1527 (N_1527,N_1288,N_1435);
nand U1528 (N_1528,N_1484,N_1383);
nand U1529 (N_1529,N_1371,N_1364);
nand U1530 (N_1530,N_1213,N_1382);
xor U1531 (N_1531,N_1322,N_1272);
and U1532 (N_1532,N_1220,N_1301);
nor U1533 (N_1533,N_1370,N_1447);
nor U1534 (N_1534,N_1402,N_1397);
xor U1535 (N_1535,N_1279,N_1358);
xnor U1536 (N_1536,N_1380,N_1309);
xor U1537 (N_1537,N_1247,N_1418);
and U1538 (N_1538,N_1330,N_1365);
xor U1539 (N_1539,N_1416,N_1388);
xnor U1540 (N_1540,N_1256,N_1335);
or U1541 (N_1541,N_1485,N_1209);
nor U1542 (N_1542,N_1205,N_1254);
nor U1543 (N_1543,N_1219,N_1491);
nand U1544 (N_1544,N_1394,N_1325);
xnor U1545 (N_1545,N_1227,N_1472);
nor U1546 (N_1546,N_1310,N_1299);
or U1547 (N_1547,N_1363,N_1454);
nand U1548 (N_1548,N_1478,N_1313);
and U1549 (N_1549,N_1208,N_1355);
nor U1550 (N_1550,N_1240,N_1429);
and U1551 (N_1551,N_1303,N_1334);
and U1552 (N_1552,N_1225,N_1216);
or U1553 (N_1553,N_1426,N_1249);
or U1554 (N_1554,N_1393,N_1321);
and U1555 (N_1555,N_1258,N_1469);
xnor U1556 (N_1556,N_1257,N_1424);
nor U1557 (N_1557,N_1450,N_1252);
nand U1558 (N_1558,N_1409,N_1350);
or U1559 (N_1559,N_1461,N_1353);
xor U1560 (N_1560,N_1296,N_1456);
and U1561 (N_1561,N_1251,N_1372);
nand U1562 (N_1562,N_1306,N_1399);
or U1563 (N_1563,N_1230,N_1294);
nor U1564 (N_1564,N_1381,N_1466);
and U1565 (N_1565,N_1243,N_1385);
or U1566 (N_1566,N_1229,N_1420);
nor U1567 (N_1567,N_1314,N_1352);
nor U1568 (N_1568,N_1440,N_1433);
nor U1569 (N_1569,N_1366,N_1489);
and U1570 (N_1570,N_1342,N_1319);
nand U1571 (N_1571,N_1441,N_1202);
nor U1572 (N_1572,N_1223,N_1480);
or U1573 (N_1573,N_1292,N_1442);
or U1574 (N_1574,N_1375,N_1486);
and U1575 (N_1575,N_1207,N_1459);
or U1576 (N_1576,N_1412,N_1255);
and U1577 (N_1577,N_1235,N_1408);
and U1578 (N_1578,N_1490,N_1473);
or U1579 (N_1579,N_1476,N_1217);
or U1580 (N_1580,N_1339,N_1326);
nor U1581 (N_1581,N_1286,N_1233);
xnor U1582 (N_1582,N_1302,N_1446);
nand U1583 (N_1583,N_1387,N_1297);
or U1584 (N_1584,N_1455,N_1498);
and U1585 (N_1585,N_1211,N_1404);
nand U1586 (N_1586,N_1373,N_1343);
and U1587 (N_1587,N_1432,N_1269);
xnor U1588 (N_1588,N_1413,N_1360);
or U1589 (N_1589,N_1250,N_1497);
and U1590 (N_1590,N_1242,N_1414);
and U1591 (N_1591,N_1246,N_1341);
nor U1592 (N_1592,N_1468,N_1453);
nor U1593 (N_1593,N_1259,N_1417);
or U1594 (N_1594,N_1234,N_1395);
nor U1595 (N_1595,N_1263,N_1231);
nand U1596 (N_1596,N_1496,N_1362);
and U1597 (N_1597,N_1315,N_1304);
nor U1598 (N_1598,N_1391,N_1434);
and U1599 (N_1599,N_1204,N_1449);
or U1600 (N_1600,N_1287,N_1437);
and U1601 (N_1601,N_1356,N_1346);
or U1602 (N_1602,N_1368,N_1333);
xor U1603 (N_1603,N_1323,N_1445);
nand U1604 (N_1604,N_1289,N_1214);
nand U1605 (N_1605,N_1276,N_1410);
and U1606 (N_1606,N_1457,N_1336);
and U1607 (N_1607,N_1415,N_1487);
nor U1608 (N_1608,N_1444,N_1332);
nand U1609 (N_1609,N_1311,N_1357);
nor U1610 (N_1610,N_1262,N_1499);
nor U1611 (N_1611,N_1458,N_1267);
nor U1612 (N_1612,N_1493,N_1475);
xor U1613 (N_1613,N_1460,N_1273);
and U1614 (N_1614,N_1431,N_1206);
nor U1615 (N_1615,N_1300,N_1407);
and U1616 (N_1616,N_1212,N_1280);
nor U1617 (N_1617,N_1374,N_1266);
or U1618 (N_1618,N_1338,N_1348);
xor U1619 (N_1619,N_1210,N_1203);
nand U1620 (N_1620,N_1281,N_1218);
or U1621 (N_1621,N_1419,N_1403);
nor U1622 (N_1622,N_1451,N_1270);
and U1623 (N_1623,N_1238,N_1354);
xor U1624 (N_1624,N_1488,N_1421);
and U1625 (N_1625,N_1305,N_1239);
xnor U1626 (N_1626,N_1378,N_1376);
nor U1627 (N_1627,N_1401,N_1324);
and U1628 (N_1628,N_1236,N_1260);
nand U1629 (N_1629,N_1265,N_1345);
or U1630 (N_1630,N_1377,N_1329);
and U1631 (N_1631,N_1463,N_1328);
nand U1632 (N_1632,N_1411,N_1228);
nor U1633 (N_1633,N_1253,N_1474);
nor U1634 (N_1634,N_1495,N_1479);
nand U1635 (N_1635,N_1290,N_1349);
or U1636 (N_1636,N_1422,N_1430);
or U1637 (N_1637,N_1222,N_1390);
nor U1638 (N_1638,N_1481,N_1492);
xor U1639 (N_1639,N_1317,N_1201);
xnor U1640 (N_1640,N_1398,N_1494);
and U1641 (N_1641,N_1318,N_1448);
or U1642 (N_1642,N_1291,N_1439);
or U1643 (N_1643,N_1308,N_1427);
and U1644 (N_1644,N_1384,N_1351);
or U1645 (N_1645,N_1241,N_1320);
xor U1646 (N_1646,N_1224,N_1386);
xor U1647 (N_1647,N_1340,N_1428);
xnor U1648 (N_1648,N_1359,N_1271);
xor U1649 (N_1649,N_1367,N_1248);
nand U1650 (N_1650,N_1229,N_1350);
nand U1651 (N_1651,N_1215,N_1289);
or U1652 (N_1652,N_1263,N_1407);
and U1653 (N_1653,N_1325,N_1473);
or U1654 (N_1654,N_1366,N_1297);
nand U1655 (N_1655,N_1216,N_1384);
nand U1656 (N_1656,N_1496,N_1493);
xor U1657 (N_1657,N_1372,N_1362);
or U1658 (N_1658,N_1301,N_1414);
nand U1659 (N_1659,N_1328,N_1277);
nand U1660 (N_1660,N_1467,N_1268);
xnor U1661 (N_1661,N_1213,N_1204);
or U1662 (N_1662,N_1448,N_1477);
and U1663 (N_1663,N_1265,N_1423);
nand U1664 (N_1664,N_1272,N_1400);
or U1665 (N_1665,N_1208,N_1286);
and U1666 (N_1666,N_1362,N_1442);
and U1667 (N_1667,N_1341,N_1395);
nand U1668 (N_1668,N_1221,N_1229);
or U1669 (N_1669,N_1292,N_1242);
and U1670 (N_1670,N_1407,N_1365);
nor U1671 (N_1671,N_1309,N_1222);
or U1672 (N_1672,N_1221,N_1306);
and U1673 (N_1673,N_1314,N_1304);
xor U1674 (N_1674,N_1438,N_1325);
nor U1675 (N_1675,N_1346,N_1374);
or U1676 (N_1676,N_1467,N_1346);
xnor U1677 (N_1677,N_1472,N_1265);
and U1678 (N_1678,N_1422,N_1392);
or U1679 (N_1679,N_1229,N_1328);
or U1680 (N_1680,N_1475,N_1265);
xnor U1681 (N_1681,N_1463,N_1223);
xor U1682 (N_1682,N_1241,N_1318);
and U1683 (N_1683,N_1234,N_1439);
nor U1684 (N_1684,N_1340,N_1475);
xnor U1685 (N_1685,N_1259,N_1256);
nand U1686 (N_1686,N_1438,N_1446);
and U1687 (N_1687,N_1335,N_1392);
or U1688 (N_1688,N_1363,N_1362);
nand U1689 (N_1689,N_1349,N_1451);
nand U1690 (N_1690,N_1400,N_1470);
or U1691 (N_1691,N_1329,N_1450);
xor U1692 (N_1692,N_1265,N_1499);
nand U1693 (N_1693,N_1331,N_1336);
or U1694 (N_1694,N_1481,N_1371);
nor U1695 (N_1695,N_1410,N_1491);
and U1696 (N_1696,N_1430,N_1407);
or U1697 (N_1697,N_1431,N_1306);
nand U1698 (N_1698,N_1223,N_1345);
nand U1699 (N_1699,N_1353,N_1413);
xor U1700 (N_1700,N_1387,N_1250);
or U1701 (N_1701,N_1264,N_1362);
and U1702 (N_1702,N_1259,N_1376);
and U1703 (N_1703,N_1372,N_1287);
and U1704 (N_1704,N_1425,N_1352);
nand U1705 (N_1705,N_1447,N_1479);
and U1706 (N_1706,N_1368,N_1405);
nor U1707 (N_1707,N_1407,N_1259);
nor U1708 (N_1708,N_1204,N_1494);
xor U1709 (N_1709,N_1426,N_1494);
or U1710 (N_1710,N_1303,N_1345);
nand U1711 (N_1711,N_1453,N_1275);
nor U1712 (N_1712,N_1222,N_1244);
nor U1713 (N_1713,N_1355,N_1394);
xnor U1714 (N_1714,N_1372,N_1498);
nor U1715 (N_1715,N_1482,N_1475);
and U1716 (N_1716,N_1307,N_1309);
xor U1717 (N_1717,N_1227,N_1417);
and U1718 (N_1718,N_1387,N_1207);
or U1719 (N_1719,N_1414,N_1361);
nand U1720 (N_1720,N_1324,N_1320);
and U1721 (N_1721,N_1411,N_1255);
or U1722 (N_1722,N_1440,N_1389);
nand U1723 (N_1723,N_1309,N_1490);
and U1724 (N_1724,N_1279,N_1270);
xor U1725 (N_1725,N_1361,N_1392);
xnor U1726 (N_1726,N_1492,N_1472);
nor U1727 (N_1727,N_1304,N_1347);
nand U1728 (N_1728,N_1294,N_1345);
and U1729 (N_1729,N_1282,N_1484);
xnor U1730 (N_1730,N_1284,N_1414);
xor U1731 (N_1731,N_1483,N_1335);
and U1732 (N_1732,N_1307,N_1327);
xor U1733 (N_1733,N_1438,N_1265);
and U1734 (N_1734,N_1449,N_1381);
nor U1735 (N_1735,N_1337,N_1438);
xnor U1736 (N_1736,N_1207,N_1347);
nor U1737 (N_1737,N_1467,N_1222);
xnor U1738 (N_1738,N_1382,N_1202);
nor U1739 (N_1739,N_1250,N_1330);
nor U1740 (N_1740,N_1493,N_1208);
nor U1741 (N_1741,N_1272,N_1262);
and U1742 (N_1742,N_1275,N_1288);
nand U1743 (N_1743,N_1472,N_1251);
xor U1744 (N_1744,N_1448,N_1443);
or U1745 (N_1745,N_1315,N_1285);
xnor U1746 (N_1746,N_1290,N_1365);
xor U1747 (N_1747,N_1470,N_1373);
nand U1748 (N_1748,N_1334,N_1418);
nor U1749 (N_1749,N_1482,N_1296);
and U1750 (N_1750,N_1374,N_1249);
nor U1751 (N_1751,N_1453,N_1469);
and U1752 (N_1752,N_1350,N_1407);
xor U1753 (N_1753,N_1432,N_1379);
nor U1754 (N_1754,N_1337,N_1278);
and U1755 (N_1755,N_1236,N_1476);
nor U1756 (N_1756,N_1422,N_1388);
nand U1757 (N_1757,N_1426,N_1321);
nand U1758 (N_1758,N_1497,N_1253);
or U1759 (N_1759,N_1250,N_1417);
nand U1760 (N_1760,N_1421,N_1212);
xnor U1761 (N_1761,N_1327,N_1438);
and U1762 (N_1762,N_1326,N_1467);
xor U1763 (N_1763,N_1421,N_1222);
nor U1764 (N_1764,N_1358,N_1337);
or U1765 (N_1765,N_1405,N_1209);
or U1766 (N_1766,N_1353,N_1277);
nor U1767 (N_1767,N_1260,N_1225);
or U1768 (N_1768,N_1470,N_1469);
or U1769 (N_1769,N_1297,N_1266);
or U1770 (N_1770,N_1451,N_1351);
or U1771 (N_1771,N_1307,N_1249);
and U1772 (N_1772,N_1366,N_1256);
and U1773 (N_1773,N_1486,N_1420);
nand U1774 (N_1774,N_1217,N_1492);
or U1775 (N_1775,N_1403,N_1226);
nor U1776 (N_1776,N_1441,N_1408);
and U1777 (N_1777,N_1496,N_1419);
nor U1778 (N_1778,N_1416,N_1377);
and U1779 (N_1779,N_1397,N_1255);
and U1780 (N_1780,N_1229,N_1306);
and U1781 (N_1781,N_1470,N_1261);
nor U1782 (N_1782,N_1298,N_1331);
or U1783 (N_1783,N_1478,N_1435);
and U1784 (N_1784,N_1461,N_1403);
nand U1785 (N_1785,N_1487,N_1205);
xor U1786 (N_1786,N_1452,N_1275);
nor U1787 (N_1787,N_1318,N_1333);
or U1788 (N_1788,N_1496,N_1241);
nor U1789 (N_1789,N_1272,N_1415);
nor U1790 (N_1790,N_1357,N_1310);
xnor U1791 (N_1791,N_1497,N_1248);
nor U1792 (N_1792,N_1235,N_1203);
nor U1793 (N_1793,N_1322,N_1377);
xnor U1794 (N_1794,N_1443,N_1282);
and U1795 (N_1795,N_1433,N_1390);
and U1796 (N_1796,N_1389,N_1300);
nand U1797 (N_1797,N_1234,N_1240);
and U1798 (N_1798,N_1440,N_1357);
nand U1799 (N_1799,N_1252,N_1423);
nand U1800 (N_1800,N_1574,N_1723);
and U1801 (N_1801,N_1636,N_1730);
and U1802 (N_1802,N_1595,N_1703);
nand U1803 (N_1803,N_1762,N_1539);
nand U1804 (N_1804,N_1711,N_1594);
nand U1805 (N_1805,N_1562,N_1660);
or U1806 (N_1806,N_1760,N_1624);
xnor U1807 (N_1807,N_1599,N_1577);
or U1808 (N_1808,N_1671,N_1546);
or U1809 (N_1809,N_1572,N_1775);
and U1810 (N_1810,N_1503,N_1558);
or U1811 (N_1811,N_1639,N_1754);
nor U1812 (N_1812,N_1677,N_1581);
nor U1813 (N_1813,N_1783,N_1786);
and U1814 (N_1814,N_1515,N_1683);
or U1815 (N_1815,N_1528,N_1547);
nand U1816 (N_1816,N_1543,N_1611);
and U1817 (N_1817,N_1731,N_1779);
or U1818 (N_1818,N_1759,N_1705);
xor U1819 (N_1819,N_1742,N_1701);
and U1820 (N_1820,N_1522,N_1712);
nor U1821 (N_1821,N_1688,N_1536);
nand U1822 (N_1822,N_1798,N_1641);
and U1823 (N_1823,N_1591,N_1554);
and U1824 (N_1824,N_1715,N_1774);
nand U1825 (N_1825,N_1746,N_1598);
xnor U1826 (N_1826,N_1517,N_1541);
or U1827 (N_1827,N_1691,N_1649);
and U1828 (N_1828,N_1771,N_1619);
and U1829 (N_1829,N_1578,N_1732);
or U1830 (N_1830,N_1606,N_1645);
nand U1831 (N_1831,N_1692,N_1585);
xnor U1832 (N_1832,N_1560,N_1769);
nor U1833 (N_1833,N_1670,N_1655);
nor U1834 (N_1834,N_1700,N_1780);
nor U1835 (N_1835,N_1716,N_1678);
and U1836 (N_1836,N_1766,N_1593);
nand U1837 (N_1837,N_1568,N_1650);
nand U1838 (N_1838,N_1714,N_1796);
nand U1839 (N_1839,N_1752,N_1566);
nand U1840 (N_1840,N_1525,N_1708);
nor U1841 (N_1841,N_1697,N_1721);
nor U1842 (N_1842,N_1596,N_1728);
nand U1843 (N_1843,N_1643,N_1529);
or U1844 (N_1844,N_1637,N_1602);
or U1845 (N_1845,N_1533,N_1513);
xnor U1846 (N_1846,N_1563,N_1506);
and U1847 (N_1847,N_1516,N_1761);
nand U1848 (N_1848,N_1662,N_1584);
or U1849 (N_1849,N_1629,N_1787);
and U1850 (N_1850,N_1665,N_1644);
and U1851 (N_1851,N_1537,N_1699);
xnor U1852 (N_1852,N_1524,N_1550);
nor U1853 (N_1853,N_1505,N_1718);
and U1854 (N_1854,N_1763,N_1621);
and U1855 (N_1855,N_1532,N_1792);
xor U1856 (N_1856,N_1635,N_1628);
or U1857 (N_1857,N_1768,N_1674);
nor U1858 (N_1858,N_1667,N_1686);
nand U1859 (N_1859,N_1733,N_1735);
xor U1860 (N_1860,N_1685,N_1738);
and U1861 (N_1861,N_1592,N_1657);
and U1862 (N_1862,N_1672,N_1616);
or U1863 (N_1863,N_1579,N_1608);
and U1864 (N_1864,N_1615,N_1758);
and U1865 (N_1865,N_1648,N_1545);
and U1866 (N_1866,N_1729,N_1724);
xor U1867 (N_1867,N_1765,N_1666);
nor U1868 (N_1868,N_1642,N_1739);
and U1869 (N_1869,N_1510,N_1534);
xnor U1870 (N_1870,N_1673,N_1613);
nor U1871 (N_1871,N_1632,N_1755);
xor U1872 (N_1872,N_1757,N_1795);
nor U1873 (N_1873,N_1720,N_1736);
and U1874 (N_1874,N_1609,N_1552);
and U1875 (N_1875,N_1740,N_1682);
nand U1876 (N_1876,N_1502,N_1640);
nor U1877 (N_1877,N_1693,N_1734);
or U1878 (N_1878,N_1535,N_1527);
nand U1879 (N_1879,N_1791,N_1514);
nand U1880 (N_1880,N_1538,N_1794);
or U1881 (N_1881,N_1777,N_1744);
or U1882 (N_1882,N_1586,N_1601);
nand U1883 (N_1883,N_1590,N_1508);
nand U1884 (N_1884,N_1509,N_1668);
nand U1885 (N_1885,N_1719,N_1631);
nor U1886 (N_1886,N_1564,N_1694);
nor U1887 (N_1887,N_1764,N_1651);
and U1888 (N_1888,N_1698,N_1512);
nor U1889 (N_1889,N_1751,N_1767);
nand U1890 (N_1890,N_1776,N_1680);
and U1891 (N_1891,N_1523,N_1521);
nor U1892 (N_1892,N_1669,N_1797);
xnor U1893 (N_1893,N_1748,N_1570);
or U1894 (N_1894,N_1737,N_1675);
or U1895 (N_1895,N_1588,N_1747);
or U1896 (N_1896,N_1749,N_1582);
nand U1897 (N_1897,N_1542,N_1713);
xnor U1898 (N_1898,N_1696,N_1600);
xnor U1899 (N_1899,N_1501,N_1571);
and U1900 (N_1900,N_1784,N_1702);
or U1901 (N_1901,N_1553,N_1630);
nor U1902 (N_1902,N_1551,N_1663);
or U1903 (N_1903,N_1531,N_1709);
or U1904 (N_1904,N_1626,N_1638);
and U1905 (N_1905,N_1679,N_1530);
and U1906 (N_1906,N_1726,N_1559);
and U1907 (N_1907,N_1567,N_1633);
or U1908 (N_1908,N_1587,N_1565);
and U1909 (N_1909,N_1526,N_1790);
nor U1910 (N_1910,N_1681,N_1722);
nor U1911 (N_1911,N_1604,N_1684);
and U1912 (N_1912,N_1659,N_1576);
nor U1913 (N_1913,N_1653,N_1612);
xor U1914 (N_1914,N_1557,N_1781);
nand U1915 (N_1915,N_1520,N_1540);
xnor U1916 (N_1916,N_1778,N_1770);
nand U1917 (N_1917,N_1610,N_1706);
or U1918 (N_1918,N_1756,N_1556);
xor U1919 (N_1919,N_1773,N_1789);
or U1920 (N_1920,N_1549,N_1504);
and U1921 (N_1921,N_1597,N_1580);
and U1922 (N_1922,N_1573,N_1753);
xor U1923 (N_1923,N_1676,N_1658);
nand U1924 (N_1924,N_1518,N_1717);
and U1925 (N_1925,N_1695,N_1583);
and U1926 (N_1926,N_1605,N_1710);
or U1927 (N_1927,N_1607,N_1743);
nor U1928 (N_1928,N_1647,N_1622);
and U1929 (N_1929,N_1785,N_1569);
nor U1930 (N_1930,N_1656,N_1687);
xnor U1931 (N_1931,N_1548,N_1652);
nand U1932 (N_1932,N_1614,N_1745);
nand U1933 (N_1933,N_1788,N_1623);
or U1934 (N_1934,N_1544,N_1690);
xor U1935 (N_1935,N_1634,N_1689);
nor U1936 (N_1936,N_1575,N_1741);
nand U1937 (N_1937,N_1617,N_1519);
and U1938 (N_1938,N_1727,N_1793);
nor U1939 (N_1939,N_1782,N_1625);
nor U1940 (N_1940,N_1620,N_1555);
nor U1941 (N_1941,N_1589,N_1725);
and U1942 (N_1942,N_1654,N_1511);
nand U1943 (N_1943,N_1646,N_1664);
and U1944 (N_1944,N_1618,N_1627);
nand U1945 (N_1945,N_1500,N_1603);
or U1946 (N_1946,N_1707,N_1750);
nor U1947 (N_1947,N_1507,N_1772);
or U1948 (N_1948,N_1799,N_1661);
or U1949 (N_1949,N_1704,N_1561);
nand U1950 (N_1950,N_1564,N_1717);
and U1951 (N_1951,N_1621,N_1732);
or U1952 (N_1952,N_1730,N_1785);
and U1953 (N_1953,N_1591,N_1792);
and U1954 (N_1954,N_1666,N_1647);
nor U1955 (N_1955,N_1646,N_1704);
nand U1956 (N_1956,N_1585,N_1704);
and U1957 (N_1957,N_1723,N_1753);
xor U1958 (N_1958,N_1594,N_1577);
nand U1959 (N_1959,N_1646,N_1726);
nand U1960 (N_1960,N_1792,N_1649);
xor U1961 (N_1961,N_1778,N_1550);
or U1962 (N_1962,N_1637,N_1798);
or U1963 (N_1963,N_1679,N_1649);
and U1964 (N_1964,N_1506,N_1610);
xnor U1965 (N_1965,N_1619,N_1758);
and U1966 (N_1966,N_1589,N_1719);
nand U1967 (N_1967,N_1587,N_1564);
nand U1968 (N_1968,N_1650,N_1550);
xnor U1969 (N_1969,N_1500,N_1706);
or U1970 (N_1970,N_1783,N_1707);
nor U1971 (N_1971,N_1664,N_1536);
nor U1972 (N_1972,N_1766,N_1571);
nor U1973 (N_1973,N_1532,N_1585);
and U1974 (N_1974,N_1730,N_1589);
nor U1975 (N_1975,N_1571,N_1743);
and U1976 (N_1976,N_1678,N_1567);
or U1977 (N_1977,N_1512,N_1766);
nand U1978 (N_1978,N_1734,N_1727);
xnor U1979 (N_1979,N_1551,N_1662);
nand U1980 (N_1980,N_1562,N_1536);
xor U1981 (N_1981,N_1550,N_1502);
xor U1982 (N_1982,N_1502,N_1617);
nand U1983 (N_1983,N_1712,N_1636);
nor U1984 (N_1984,N_1742,N_1709);
and U1985 (N_1985,N_1685,N_1671);
and U1986 (N_1986,N_1569,N_1707);
xor U1987 (N_1987,N_1543,N_1519);
and U1988 (N_1988,N_1783,N_1527);
and U1989 (N_1989,N_1748,N_1671);
and U1990 (N_1990,N_1764,N_1715);
nand U1991 (N_1991,N_1662,N_1500);
and U1992 (N_1992,N_1518,N_1665);
xor U1993 (N_1993,N_1522,N_1728);
xor U1994 (N_1994,N_1733,N_1720);
nand U1995 (N_1995,N_1543,N_1532);
xnor U1996 (N_1996,N_1788,N_1713);
nor U1997 (N_1997,N_1600,N_1786);
or U1998 (N_1998,N_1532,N_1523);
nand U1999 (N_1999,N_1579,N_1690);
nand U2000 (N_2000,N_1653,N_1697);
xnor U2001 (N_2001,N_1526,N_1632);
nand U2002 (N_2002,N_1741,N_1591);
and U2003 (N_2003,N_1570,N_1560);
xor U2004 (N_2004,N_1590,N_1743);
nor U2005 (N_2005,N_1752,N_1754);
nand U2006 (N_2006,N_1740,N_1725);
and U2007 (N_2007,N_1697,N_1678);
nor U2008 (N_2008,N_1690,N_1556);
xor U2009 (N_2009,N_1640,N_1624);
nor U2010 (N_2010,N_1549,N_1711);
or U2011 (N_2011,N_1763,N_1728);
and U2012 (N_2012,N_1672,N_1766);
xnor U2013 (N_2013,N_1774,N_1504);
nor U2014 (N_2014,N_1680,N_1725);
or U2015 (N_2015,N_1594,N_1784);
or U2016 (N_2016,N_1599,N_1769);
and U2017 (N_2017,N_1555,N_1505);
xnor U2018 (N_2018,N_1560,N_1624);
xnor U2019 (N_2019,N_1625,N_1576);
nand U2020 (N_2020,N_1695,N_1687);
nand U2021 (N_2021,N_1586,N_1535);
nor U2022 (N_2022,N_1696,N_1506);
or U2023 (N_2023,N_1766,N_1768);
or U2024 (N_2024,N_1680,N_1540);
xor U2025 (N_2025,N_1562,N_1620);
and U2026 (N_2026,N_1791,N_1777);
or U2027 (N_2027,N_1507,N_1727);
xor U2028 (N_2028,N_1614,N_1739);
nor U2029 (N_2029,N_1660,N_1549);
and U2030 (N_2030,N_1693,N_1567);
nor U2031 (N_2031,N_1596,N_1532);
and U2032 (N_2032,N_1761,N_1729);
and U2033 (N_2033,N_1744,N_1780);
or U2034 (N_2034,N_1536,N_1574);
nand U2035 (N_2035,N_1538,N_1666);
or U2036 (N_2036,N_1565,N_1526);
xnor U2037 (N_2037,N_1754,N_1610);
and U2038 (N_2038,N_1714,N_1600);
nand U2039 (N_2039,N_1688,N_1624);
xnor U2040 (N_2040,N_1760,N_1745);
or U2041 (N_2041,N_1568,N_1673);
xor U2042 (N_2042,N_1732,N_1553);
or U2043 (N_2043,N_1552,N_1515);
nand U2044 (N_2044,N_1518,N_1792);
and U2045 (N_2045,N_1716,N_1675);
nor U2046 (N_2046,N_1554,N_1710);
or U2047 (N_2047,N_1589,N_1724);
or U2048 (N_2048,N_1777,N_1749);
nor U2049 (N_2049,N_1509,N_1622);
or U2050 (N_2050,N_1510,N_1710);
and U2051 (N_2051,N_1679,N_1687);
xor U2052 (N_2052,N_1726,N_1508);
nor U2053 (N_2053,N_1618,N_1560);
and U2054 (N_2054,N_1726,N_1669);
nor U2055 (N_2055,N_1694,N_1601);
xor U2056 (N_2056,N_1727,N_1685);
or U2057 (N_2057,N_1590,N_1539);
and U2058 (N_2058,N_1593,N_1712);
and U2059 (N_2059,N_1615,N_1745);
or U2060 (N_2060,N_1781,N_1673);
xnor U2061 (N_2061,N_1606,N_1507);
or U2062 (N_2062,N_1546,N_1522);
nor U2063 (N_2063,N_1514,N_1767);
nor U2064 (N_2064,N_1564,N_1586);
or U2065 (N_2065,N_1739,N_1503);
nand U2066 (N_2066,N_1670,N_1746);
nor U2067 (N_2067,N_1678,N_1665);
or U2068 (N_2068,N_1731,N_1646);
or U2069 (N_2069,N_1727,N_1788);
nor U2070 (N_2070,N_1743,N_1788);
xnor U2071 (N_2071,N_1718,N_1612);
and U2072 (N_2072,N_1603,N_1620);
nor U2073 (N_2073,N_1634,N_1714);
xor U2074 (N_2074,N_1500,N_1631);
nor U2075 (N_2075,N_1571,N_1592);
nand U2076 (N_2076,N_1718,N_1620);
or U2077 (N_2077,N_1549,N_1554);
and U2078 (N_2078,N_1660,N_1739);
or U2079 (N_2079,N_1794,N_1685);
nor U2080 (N_2080,N_1713,N_1623);
xor U2081 (N_2081,N_1552,N_1523);
xnor U2082 (N_2082,N_1534,N_1553);
nor U2083 (N_2083,N_1596,N_1754);
or U2084 (N_2084,N_1536,N_1658);
or U2085 (N_2085,N_1646,N_1608);
or U2086 (N_2086,N_1749,N_1790);
and U2087 (N_2087,N_1696,N_1683);
and U2088 (N_2088,N_1553,N_1649);
xnor U2089 (N_2089,N_1775,N_1666);
xnor U2090 (N_2090,N_1623,N_1603);
xor U2091 (N_2091,N_1720,N_1521);
nor U2092 (N_2092,N_1527,N_1653);
nor U2093 (N_2093,N_1662,N_1790);
or U2094 (N_2094,N_1638,N_1598);
nor U2095 (N_2095,N_1685,N_1682);
xnor U2096 (N_2096,N_1676,N_1519);
and U2097 (N_2097,N_1582,N_1617);
xnor U2098 (N_2098,N_1531,N_1559);
and U2099 (N_2099,N_1589,N_1518);
or U2100 (N_2100,N_1850,N_1907);
nor U2101 (N_2101,N_2071,N_2064);
and U2102 (N_2102,N_1948,N_1977);
nand U2103 (N_2103,N_1988,N_1959);
or U2104 (N_2104,N_1963,N_1923);
or U2105 (N_2105,N_2055,N_1950);
xor U2106 (N_2106,N_1897,N_1875);
and U2107 (N_2107,N_1935,N_2043);
or U2108 (N_2108,N_1856,N_1934);
or U2109 (N_2109,N_2081,N_1927);
and U2110 (N_2110,N_1840,N_1857);
xor U2111 (N_2111,N_1849,N_2034);
nor U2112 (N_2112,N_1867,N_1929);
and U2113 (N_2113,N_1917,N_1839);
nor U2114 (N_2114,N_1976,N_1951);
and U2115 (N_2115,N_1933,N_1932);
or U2116 (N_2116,N_1810,N_1825);
xor U2117 (N_2117,N_2046,N_1922);
and U2118 (N_2118,N_1961,N_1985);
and U2119 (N_2119,N_1982,N_2020);
nand U2120 (N_2120,N_1994,N_1800);
xor U2121 (N_2121,N_1868,N_2051);
and U2122 (N_2122,N_2076,N_1989);
nand U2123 (N_2123,N_1892,N_1823);
xor U2124 (N_2124,N_2011,N_1848);
nand U2125 (N_2125,N_1805,N_1811);
xnor U2126 (N_2126,N_2066,N_1979);
nor U2127 (N_2127,N_1945,N_1854);
or U2128 (N_2128,N_1835,N_1949);
xnor U2129 (N_2129,N_2023,N_1987);
nor U2130 (N_2130,N_1874,N_1879);
nor U2131 (N_2131,N_2030,N_1964);
nor U2132 (N_2132,N_1896,N_2008);
nor U2133 (N_2133,N_1953,N_2017);
nand U2134 (N_2134,N_2028,N_1807);
and U2135 (N_2135,N_1816,N_1828);
and U2136 (N_2136,N_2084,N_1906);
and U2137 (N_2137,N_1992,N_1926);
and U2138 (N_2138,N_2009,N_1877);
or U2139 (N_2139,N_1946,N_1954);
or U2140 (N_2140,N_1899,N_2018);
nand U2141 (N_2141,N_2058,N_1995);
and U2142 (N_2142,N_1903,N_1912);
or U2143 (N_2143,N_1930,N_2033);
nand U2144 (N_2144,N_2089,N_1938);
and U2145 (N_2145,N_2073,N_2001);
xor U2146 (N_2146,N_1936,N_1806);
and U2147 (N_2147,N_1916,N_2098);
and U2148 (N_2148,N_2053,N_1966);
or U2149 (N_2149,N_2085,N_1815);
and U2150 (N_2150,N_1830,N_1900);
nor U2151 (N_2151,N_1991,N_2003);
xor U2152 (N_2152,N_1838,N_1984);
nand U2153 (N_2153,N_1824,N_2025);
or U2154 (N_2154,N_1822,N_1801);
or U2155 (N_2155,N_1843,N_1813);
and U2156 (N_2156,N_1844,N_1972);
nor U2157 (N_2157,N_1915,N_1853);
nand U2158 (N_2158,N_1847,N_2036);
nand U2159 (N_2159,N_2068,N_2010);
or U2160 (N_2160,N_1837,N_2060);
nand U2161 (N_2161,N_2056,N_1993);
xnor U2162 (N_2162,N_1817,N_2087);
nand U2163 (N_2163,N_1864,N_1866);
and U2164 (N_2164,N_2093,N_1956);
xnor U2165 (N_2165,N_1971,N_1920);
and U2166 (N_2166,N_2002,N_1908);
nor U2167 (N_2167,N_2040,N_2015);
nor U2168 (N_2168,N_2052,N_1852);
or U2169 (N_2169,N_1981,N_1952);
nand U2170 (N_2170,N_1962,N_1970);
xor U2171 (N_2171,N_1858,N_1834);
and U2172 (N_2172,N_2007,N_1913);
nand U2173 (N_2173,N_2061,N_2075);
nor U2174 (N_2174,N_1990,N_2057);
xor U2175 (N_2175,N_1944,N_1855);
nand U2176 (N_2176,N_1888,N_1905);
xnor U2177 (N_2177,N_1902,N_2039);
and U2178 (N_2178,N_1802,N_1865);
nand U2179 (N_2179,N_1898,N_2095);
and U2180 (N_2180,N_1921,N_1942);
or U2181 (N_2181,N_1960,N_2054);
xor U2182 (N_2182,N_2045,N_2005);
or U2183 (N_2183,N_1873,N_2027);
nor U2184 (N_2184,N_1832,N_1872);
xnor U2185 (N_2185,N_1821,N_2042);
nor U2186 (N_2186,N_1863,N_2035);
nand U2187 (N_2187,N_1885,N_2080);
or U2188 (N_2188,N_1870,N_1860);
nand U2189 (N_2189,N_1886,N_1996);
and U2190 (N_2190,N_2049,N_1943);
or U2191 (N_2191,N_1881,N_2016);
xnor U2192 (N_2192,N_2065,N_1974);
or U2193 (N_2193,N_2078,N_1831);
nand U2194 (N_2194,N_1998,N_2091);
and U2195 (N_2195,N_2026,N_2031);
or U2196 (N_2196,N_2072,N_1827);
nor U2197 (N_2197,N_2069,N_1895);
and U2198 (N_2198,N_2082,N_2022);
nand U2199 (N_2199,N_2047,N_1983);
nand U2200 (N_2200,N_2059,N_1803);
and U2201 (N_2201,N_1947,N_1975);
nor U2202 (N_2202,N_1997,N_1967);
and U2203 (N_2203,N_2032,N_2000);
or U2204 (N_2204,N_2037,N_2024);
nor U2205 (N_2205,N_1909,N_1818);
xnor U2206 (N_2206,N_1887,N_1928);
and U2207 (N_2207,N_2013,N_1883);
nor U2208 (N_2208,N_2086,N_1958);
and U2209 (N_2209,N_1980,N_2079);
xnor U2210 (N_2210,N_1876,N_1869);
xnor U2211 (N_2211,N_2019,N_1999);
xor U2212 (N_2212,N_1812,N_2062);
xor U2213 (N_2213,N_1845,N_1836);
xnor U2214 (N_2214,N_1808,N_2094);
and U2215 (N_2215,N_1878,N_1891);
xnor U2216 (N_2216,N_2074,N_2048);
and U2217 (N_2217,N_1809,N_1969);
xor U2218 (N_2218,N_1973,N_1851);
and U2219 (N_2219,N_2006,N_1965);
xor U2220 (N_2220,N_1919,N_1814);
nand U2221 (N_2221,N_1904,N_1914);
and U2222 (N_2222,N_1986,N_2083);
or U2223 (N_2223,N_1884,N_1901);
and U2224 (N_2224,N_1931,N_1925);
and U2225 (N_2225,N_2004,N_1871);
nor U2226 (N_2226,N_2070,N_1941);
nand U2227 (N_2227,N_1882,N_1889);
or U2228 (N_2228,N_1829,N_2077);
or U2229 (N_2229,N_1937,N_1924);
and U2230 (N_2230,N_2044,N_2029);
nor U2231 (N_2231,N_1804,N_1911);
xnor U2232 (N_2232,N_1862,N_1893);
and U2233 (N_2233,N_2038,N_1918);
xor U2234 (N_2234,N_1978,N_1841);
and U2235 (N_2235,N_1826,N_2092);
and U2236 (N_2236,N_1880,N_2014);
nand U2237 (N_2237,N_2096,N_2097);
nand U2238 (N_2238,N_1910,N_2041);
nor U2239 (N_2239,N_2063,N_1940);
xnor U2240 (N_2240,N_1890,N_2050);
or U2241 (N_2241,N_2021,N_1859);
nor U2242 (N_2242,N_2099,N_2012);
xor U2243 (N_2243,N_1846,N_1955);
nand U2244 (N_2244,N_1957,N_1833);
or U2245 (N_2245,N_1820,N_2090);
or U2246 (N_2246,N_2067,N_1819);
nor U2247 (N_2247,N_1842,N_1861);
and U2248 (N_2248,N_1894,N_2088);
xor U2249 (N_2249,N_1939,N_1968);
nor U2250 (N_2250,N_2042,N_2093);
or U2251 (N_2251,N_1891,N_2007);
and U2252 (N_2252,N_2056,N_1851);
nand U2253 (N_2253,N_1882,N_1906);
nor U2254 (N_2254,N_1874,N_1990);
xnor U2255 (N_2255,N_1801,N_1910);
or U2256 (N_2256,N_1882,N_1981);
or U2257 (N_2257,N_1881,N_1883);
or U2258 (N_2258,N_2044,N_1895);
and U2259 (N_2259,N_2060,N_2093);
nand U2260 (N_2260,N_2039,N_2090);
nor U2261 (N_2261,N_1935,N_1849);
nand U2262 (N_2262,N_2040,N_1988);
and U2263 (N_2263,N_1886,N_2072);
xnor U2264 (N_2264,N_1995,N_1828);
and U2265 (N_2265,N_2007,N_1928);
and U2266 (N_2266,N_1934,N_1857);
nand U2267 (N_2267,N_1824,N_2099);
nor U2268 (N_2268,N_2096,N_2050);
and U2269 (N_2269,N_1825,N_1973);
xor U2270 (N_2270,N_2030,N_2012);
nor U2271 (N_2271,N_1956,N_2045);
xor U2272 (N_2272,N_1986,N_2031);
nor U2273 (N_2273,N_1957,N_1919);
xor U2274 (N_2274,N_1809,N_1935);
nor U2275 (N_2275,N_1956,N_1910);
and U2276 (N_2276,N_1847,N_1903);
xnor U2277 (N_2277,N_1999,N_2020);
and U2278 (N_2278,N_1873,N_2010);
xor U2279 (N_2279,N_1898,N_1834);
or U2280 (N_2280,N_2097,N_1884);
xor U2281 (N_2281,N_1977,N_1816);
or U2282 (N_2282,N_1889,N_1979);
and U2283 (N_2283,N_1843,N_1808);
and U2284 (N_2284,N_1868,N_2078);
nand U2285 (N_2285,N_1845,N_1926);
xnor U2286 (N_2286,N_1979,N_2043);
or U2287 (N_2287,N_1992,N_2000);
and U2288 (N_2288,N_1897,N_2098);
nand U2289 (N_2289,N_1939,N_1962);
and U2290 (N_2290,N_1958,N_2027);
or U2291 (N_2291,N_1945,N_1975);
nand U2292 (N_2292,N_1834,N_1908);
nor U2293 (N_2293,N_2097,N_1942);
nand U2294 (N_2294,N_2094,N_1980);
nor U2295 (N_2295,N_1997,N_1833);
or U2296 (N_2296,N_2095,N_1938);
and U2297 (N_2297,N_1980,N_2077);
nor U2298 (N_2298,N_1952,N_2003);
nor U2299 (N_2299,N_1939,N_1896);
nor U2300 (N_2300,N_2037,N_2098);
or U2301 (N_2301,N_1837,N_2004);
nor U2302 (N_2302,N_1845,N_2068);
or U2303 (N_2303,N_1921,N_2025);
xor U2304 (N_2304,N_2089,N_1801);
and U2305 (N_2305,N_1850,N_1855);
and U2306 (N_2306,N_1903,N_1888);
nor U2307 (N_2307,N_1896,N_1813);
and U2308 (N_2308,N_1810,N_2022);
or U2309 (N_2309,N_1878,N_1896);
nand U2310 (N_2310,N_1852,N_1824);
xor U2311 (N_2311,N_1873,N_1920);
xor U2312 (N_2312,N_1804,N_1943);
nor U2313 (N_2313,N_1960,N_2081);
nand U2314 (N_2314,N_2059,N_1956);
or U2315 (N_2315,N_1911,N_2011);
and U2316 (N_2316,N_1864,N_1842);
nand U2317 (N_2317,N_2092,N_1931);
nand U2318 (N_2318,N_2006,N_1834);
nand U2319 (N_2319,N_1974,N_1954);
nand U2320 (N_2320,N_1905,N_1857);
and U2321 (N_2321,N_2048,N_1966);
or U2322 (N_2322,N_1929,N_1980);
and U2323 (N_2323,N_1868,N_1824);
xor U2324 (N_2324,N_2003,N_2051);
and U2325 (N_2325,N_1929,N_1857);
and U2326 (N_2326,N_1982,N_1999);
and U2327 (N_2327,N_2068,N_2083);
nor U2328 (N_2328,N_1921,N_1805);
or U2329 (N_2329,N_2005,N_1956);
or U2330 (N_2330,N_1989,N_1919);
nor U2331 (N_2331,N_2006,N_2026);
and U2332 (N_2332,N_2019,N_1993);
nand U2333 (N_2333,N_2092,N_1953);
nor U2334 (N_2334,N_1956,N_1930);
xor U2335 (N_2335,N_2035,N_1997);
nand U2336 (N_2336,N_2001,N_1852);
xor U2337 (N_2337,N_1946,N_1890);
and U2338 (N_2338,N_1871,N_1853);
nand U2339 (N_2339,N_1888,N_1836);
or U2340 (N_2340,N_2062,N_1894);
nand U2341 (N_2341,N_1865,N_2054);
and U2342 (N_2342,N_1992,N_2068);
nor U2343 (N_2343,N_1974,N_1969);
nand U2344 (N_2344,N_2072,N_1851);
nor U2345 (N_2345,N_2056,N_1858);
xor U2346 (N_2346,N_1843,N_2068);
nand U2347 (N_2347,N_1959,N_1954);
or U2348 (N_2348,N_1977,N_2052);
nor U2349 (N_2349,N_1980,N_2057);
xor U2350 (N_2350,N_1951,N_2051);
or U2351 (N_2351,N_1876,N_1915);
and U2352 (N_2352,N_1920,N_2022);
nor U2353 (N_2353,N_2064,N_1980);
and U2354 (N_2354,N_1937,N_2073);
xor U2355 (N_2355,N_1941,N_1883);
nand U2356 (N_2356,N_1805,N_1946);
nand U2357 (N_2357,N_2050,N_1916);
or U2358 (N_2358,N_1833,N_1823);
nand U2359 (N_2359,N_2012,N_1869);
nand U2360 (N_2360,N_2061,N_1936);
and U2361 (N_2361,N_1883,N_1918);
nand U2362 (N_2362,N_2083,N_1923);
or U2363 (N_2363,N_1955,N_1808);
nand U2364 (N_2364,N_1874,N_1936);
nor U2365 (N_2365,N_1907,N_1901);
nand U2366 (N_2366,N_2034,N_1804);
nor U2367 (N_2367,N_1956,N_1882);
xnor U2368 (N_2368,N_1978,N_1938);
and U2369 (N_2369,N_1827,N_2029);
xnor U2370 (N_2370,N_2065,N_1935);
or U2371 (N_2371,N_1923,N_2084);
or U2372 (N_2372,N_1927,N_1827);
xor U2373 (N_2373,N_2067,N_1909);
and U2374 (N_2374,N_2011,N_1871);
nand U2375 (N_2375,N_2010,N_2034);
xnor U2376 (N_2376,N_1949,N_2041);
xnor U2377 (N_2377,N_1856,N_2079);
nor U2378 (N_2378,N_1928,N_2063);
nor U2379 (N_2379,N_2038,N_1944);
xor U2380 (N_2380,N_1982,N_2049);
nor U2381 (N_2381,N_1879,N_1817);
nand U2382 (N_2382,N_1848,N_2060);
and U2383 (N_2383,N_1989,N_1850);
nor U2384 (N_2384,N_1885,N_1970);
or U2385 (N_2385,N_2016,N_1938);
nand U2386 (N_2386,N_2095,N_1993);
nand U2387 (N_2387,N_1999,N_2057);
nand U2388 (N_2388,N_1875,N_1830);
and U2389 (N_2389,N_2001,N_2069);
xor U2390 (N_2390,N_2082,N_1900);
or U2391 (N_2391,N_1896,N_1866);
xor U2392 (N_2392,N_1979,N_1990);
or U2393 (N_2393,N_2049,N_2086);
nor U2394 (N_2394,N_1879,N_1951);
xnor U2395 (N_2395,N_2044,N_1861);
and U2396 (N_2396,N_1899,N_1886);
or U2397 (N_2397,N_1857,N_1824);
or U2398 (N_2398,N_2088,N_2071);
nor U2399 (N_2399,N_2053,N_2004);
and U2400 (N_2400,N_2398,N_2311);
nor U2401 (N_2401,N_2274,N_2336);
or U2402 (N_2402,N_2265,N_2345);
or U2403 (N_2403,N_2360,N_2239);
xnor U2404 (N_2404,N_2382,N_2152);
and U2405 (N_2405,N_2300,N_2316);
nand U2406 (N_2406,N_2351,N_2186);
and U2407 (N_2407,N_2275,N_2167);
and U2408 (N_2408,N_2225,N_2228);
xor U2409 (N_2409,N_2195,N_2286);
nand U2410 (N_2410,N_2248,N_2134);
or U2411 (N_2411,N_2372,N_2282);
nand U2412 (N_2412,N_2342,N_2333);
and U2413 (N_2413,N_2242,N_2356);
nand U2414 (N_2414,N_2133,N_2137);
xor U2415 (N_2415,N_2174,N_2249);
nand U2416 (N_2416,N_2214,N_2120);
and U2417 (N_2417,N_2289,N_2107);
xor U2418 (N_2418,N_2347,N_2264);
and U2419 (N_2419,N_2381,N_2121);
and U2420 (N_2420,N_2169,N_2375);
nand U2421 (N_2421,N_2288,N_2324);
and U2422 (N_2422,N_2396,N_2117);
or U2423 (N_2423,N_2157,N_2146);
xor U2424 (N_2424,N_2168,N_2308);
nand U2425 (N_2425,N_2335,N_2176);
nand U2426 (N_2426,N_2127,N_2113);
and U2427 (N_2427,N_2226,N_2106);
nor U2428 (N_2428,N_2302,N_2385);
nand U2429 (N_2429,N_2295,N_2217);
nor U2430 (N_2430,N_2171,N_2343);
nand U2431 (N_2431,N_2143,N_2299);
or U2432 (N_2432,N_2389,N_2251);
and U2433 (N_2433,N_2291,N_2243);
nor U2434 (N_2434,N_2196,N_2184);
and U2435 (N_2435,N_2315,N_2271);
nand U2436 (N_2436,N_2313,N_2164);
nor U2437 (N_2437,N_2180,N_2230);
or U2438 (N_2438,N_2367,N_2317);
xor U2439 (N_2439,N_2262,N_2223);
and U2440 (N_2440,N_2210,N_2260);
xor U2441 (N_2441,N_2147,N_2130);
nor U2442 (N_2442,N_2255,N_2399);
nand U2443 (N_2443,N_2211,N_2344);
xor U2444 (N_2444,N_2256,N_2278);
xnor U2445 (N_2445,N_2319,N_2155);
nand U2446 (N_2446,N_2348,N_2364);
nor U2447 (N_2447,N_2323,N_2153);
and U2448 (N_2448,N_2269,N_2188);
and U2449 (N_2449,N_2126,N_2359);
xor U2450 (N_2450,N_2213,N_2154);
nor U2451 (N_2451,N_2170,N_2349);
and U2452 (N_2452,N_2294,N_2338);
nor U2453 (N_2453,N_2236,N_2104);
nand U2454 (N_2454,N_2166,N_2292);
xnor U2455 (N_2455,N_2247,N_2200);
and U2456 (N_2456,N_2379,N_2108);
nor U2457 (N_2457,N_2114,N_2118);
or U2458 (N_2458,N_2337,N_2257);
and U2459 (N_2459,N_2142,N_2116);
and U2460 (N_2460,N_2103,N_2253);
nand U2461 (N_2461,N_2139,N_2207);
or U2462 (N_2462,N_2370,N_2136);
nand U2463 (N_2463,N_2353,N_2362);
and U2464 (N_2464,N_2327,N_2321);
nand U2465 (N_2465,N_2135,N_2306);
nor U2466 (N_2466,N_2202,N_2125);
xnor U2467 (N_2467,N_2105,N_2165);
xnor U2468 (N_2468,N_2394,N_2340);
nor U2469 (N_2469,N_2241,N_2346);
xnor U2470 (N_2470,N_2175,N_2189);
xnor U2471 (N_2471,N_2235,N_2160);
nand U2472 (N_2472,N_2222,N_2112);
xnor U2473 (N_2473,N_2270,N_2383);
nor U2474 (N_2474,N_2215,N_2150);
nor U2475 (N_2475,N_2301,N_2191);
and U2476 (N_2476,N_2290,N_2173);
xnor U2477 (N_2477,N_2197,N_2285);
and U2478 (N_2478,N_2221,N_2314);
xor U2479 (N_2479,N_2326,N_2244);
and U2480 (N_2480,N_2310,N_2201);
xor U2481 (N_2481,N_2216,N_2102);
nand U2482 (N_2482,N_2149,N_2163);
or U2483 (N_2483,N_2287,N_2199);
nor U2484 (N_2484,N_2339,N_2325);
nor U2485 (N_2485,N_2397,N_2304);
xor U2486 (N_2486,N_2266,N_2296);
nand U2487 (N_2487,N_2374,N_2240);
nand U2488 (N_2488,N_2190,N_2272);
nand U2489 (N_2489,N_2387,N_2281);
and U2490 (N_2490,N_2237,N_2129);
and U2491 (N_2491,N_2259,N_2350);
or U2492 (N_2492,N_2307,N_2238);
or U2493 (N_2493,N_2178,N_2145);
or U2494 (N_2494,N_2205,N_2277);
and U2495 (N_2495,N_2330,N_2318);
nor U2496 (N_2496,N_2123,N_2218);
and U2497 (N_2497,N_2212,N_2231);
and U2498 (N_2498,N_2193,N_2172);
and U2499 (N_2499,N_2355,N_2206);
or U2500 (N_2500,N_2388,N_2198);
nand U2501 (N_2501,N_2320,N_2378);
nor U2502 (N_2502,N_2233,N_2391);
and U2503 (N_2503,N_2151,N_2254);
xor U2504 (N_2504,N_2365,N_2395);
or U2505 (N_2505,N_2352,N_2148);
xnor U2506 (N_2506,N_2312,N_2377);
and U2507 (N_2507,N_2280,N_2267);
nand U2508 (N_2508,N_2332,N_2227);
nor U2509 (N_2509,N_2159,N_2128);
and U2510 (N_2510,N_2361,N_2181);
and U2511 (N_2511,N_2261,N_2357);
nor U2512 (N_2512,N_2279,N_2185);
or U2513 (N_2513,N_2177,N_2204);
nand U2514 (N_2514,N_2182,N_2232);
xnor U2515 (N_2515,N_2124,N_2284);
nand U2516 (N_2516,N_2366,N_2297);
xnor U2517 (N_2517,N_2328,N_2309);
xnor U2518 (N_2518,N_2293,N_2268);
and U2519 (N_2519,N_2109,N_2258);
nand U2520 (N_2520,N_2298,N_2219);
and U2521 (N_2521,N_2331,N_2111);
nand U2522 (N_2522,N_2119,N_2100);
nand U2523 (N_2523,N_2208,N_2192);
or U2524 (N_2524,N_2122,N_2371);
and U2525 (N_2525,N_2250,N_2252);
or U2526 (N_2526,N_2245,N_2334);
or U2527 (N_2527,N_2144,N_2276);
xor U2528 (N_2528,N_2393,N_2132);
nor U2529 (N_2529,N_2329,N_2368);
or U2530 (N_2530,N_2373,N_2194);
and U2531 (N_2531,N_2305,N_2322);
or U2532 (N_2532,N_2283,N_2224);
nor U2533 (N_2533,N_2380,N_2263);
or U2534 (N_2534,N_2161,N_2141);
or U2535 (N_2535,N_2303,N_2110);
nand U2536 (N_2536,N_2138,N_2203);
xor U2537 (N_2537,N_2209,N_2363);
nor U2538 (N_2538,N_2101,N_2131);
nand U2539 (N_2539,N_2390,N_2220);
xnor U2540 (N_2540,N_2140,N_2386);
nand U2541 (N_2541,N_2358,N_2392);
nor U2542 (N_2542,N_2162,N_2384);
nor U2543 (N_2543,N_2179,N_2354);
nor U2544 (N_2544,N_2115,N_2234);
nor U2545 (N_2545,N_2187,N_2376);
nand U2546 (N_2546,N_2246,N_2273);
nand U2547 (N_2547,N_2229,N_2183);
xnor U2548 (N_2548,N_2369,N_2156);
or U2549 (N_2549,N_2158,N_2341);
nor U2550 (N_2550,N_2362,N_2368);
nor U2551 (N_2551,N_2327,N_2263);
xor U2552 (N_2552,N_2207,N_2194);
or U2553 (N_2553,N_2180,N_2194);
and U2554 (N_2554,N_2383,N_2113);
nor U2555 (N_2555,N_2180,N_2357);
or U2556 (N_2556,N_2221,N_2117);
nand U2557 (N_2557,N_2201,N_2261);
or U2558 (N_2558,N_2211,N_2317);
xnor U2559 (N_2559,N_2365,N_2372);
nor U2560 (N_2560,N_2104,N_2207);
or U2561 (N_2561,N_2298,N_2341);
nor U2562 (N_2562,N_2117,N_2337);
nor U2563 (N_2563,N_2289,N_2334);
and U2564 (N_2564,N_2323,N_2197);
xnor U2565 (N_2565,N_2111,N_2310);
xor U2566 (N_2566,N_2181,N_2367);
or U2567 (N_2567,N_2334,N_2342);
nand U2568 (N_2568,N_2266,N_2263);
and U2569 (N_2569,N_2385,N_2346);
nand U2570 (N_2570,N_2271,N_2193);
nand U2571 (N_2571,N_2145,N_2153);
nor U2572 (N_2572,N_2277,N_2229);
or U2573 (N_2573,N_2332,N_2261);
and U2574 (N_2574,N_2148,N_2291);
xnor U2575 (N_2575,N_2304,N_2229);
or U2576 (N_2576,N_2188,N_2391);
nor U2577 (N_2577,N_2372,N_2206);
nor U2578 (N_2578,N_2150,N_2343);
nor U2579 (N_2579,N_2362,N_2162);
xor U2580 (N_2580,N_2208,N_2191);
nand U2581 (N_2581,N_2302,N_2334);
and U2582 (N_2582,N_2113,N_2358);
nand U2583 (N_2583,N_2351,N_2220);
xnor U2584 (N_2584,N_2187,N_2266);
nand U2585 (N_2585,N_2321,N_2212);
or U2586 (N_2586,N_2238,N_2217);
or U2587 (N_2587,N_2382,N_2175);
xnor U2588 (N_2588,N_2171,N_2207);
nor U2589 (N_2589,N_2382,N_2325);
or U2590 (N_2590,N_2360,N_2263);
xnor U2591 (N_2591,N_2239,N_2220);
and U2592 (N_2592,N_2202,N_2339);
xnor U2593 (N_2593,N_2135,N_2286);
or U2594 (N_2594,N_2105,N_2167);
and U2595 (N_2595,N_2350,N_2212);
or U2596 (N_2596,N_2323,N_2149);
nand U2597 (N_2597,N_2347,N_2231);
nand U2598 (N_2598,N_2201,N_2326);
and U2599 (N_2599,N_2190,N_2381);
and U2600 (N_2600,N_2295,N_2361);
and U2601 (N_2601,N_2267,N_2374);
nand U2602 (N_2602,N_2147,N_2348);
xnor U2603 (N_2603,N_2154,N_2171);
nor U2604 (N_2604,N_2211,N_2348);
nor U2605 (N_2605,N_2226,N_2228);
or U2606 (N_2606,N_2182,N_2184);
xor U2607 (N_2607,N_2222,N_2219);
and U2608 (N_2608,N_2319,N_2102);
nand U2609 (N_2609,N_2337,N_2289);
nor U2610 (N_2610,N_2289,N_2276);
and U2611 (N_2611,N_2149,N_2249);
and U2612 (N_2612,N_2327,N_2271);
nand U2613 (N_2613,N_2363,N_2311);
and U2614 (N_2614,N_2228,N_2325);
nand U2615 (N_2615,N_2356,N_2324);
nand U2616 (N_2616,N_2132,N_2196);
nand U2617 (N_2617,N_2275,N_2301);
nand U2618 (N_2618,N_2153,N_2287);
or U2619 (N_2619,N_2342,N_2201);
nor U2620 (N_2620,N_2236,N_2320);
xor U2621 (N_2621,N_2286,N_2261);
or U2622 (N_2622,N_2399,N_2102);
and U2623 (N_2623,N_2104,N_2378);
xnor U2624 (N_2624,N_2349,N_2215);
or U2625 (N_2625,N_2304,N_2211);
nor U2626 (N_2626,N_2321,N_2331);
or U2627 (N_2627,N_2148,N_2271);
and U2628 (N_2628,N_2349,N_2103);
or U2629 (N_2629,N_2122,N_2194);
xor U2630 (N_2630,N_2238,N_2125);
and U2631 (N_2631,N_2183,N_2305);
nand U2632 (N_2632,N_2105,N_2357);
nand U2633 (N_2633,N_2322,N_2202);
xor U2634 (N_2634,N_2272,N_2146);
nand U2635 (N_2635,N_2233,N_2174);
or U2636 (N_2636,N_2195,N_2311);
and U2637 (N_2637,N_2319,N_2212);
and U2638 (N_2638,N_2355,N_2225);
and U2639 (N_2639,N_2394,N_2194);
nand U2640 (N_2640,N_2180,N_2366);
xnor U2641 (N_2641,N_2261,N_2101);
nor U2642 (N_2642,N_2386,N_2118);
nand U2643 (N_2643,N_2181,N_2273);
or U2644 (N_2644,N_2385,N_2322);
and U2645 (N_2645,N_2270,N_2302);
nor U2646 (N_2646,N_2301,N_2382);
xnor U2647 (N_2647,N_2168,N_2249);
nor U2648 (N_2648,N_2373,N_2240);
nand U2649 (N_2649,N_2168,N_2398);
nand U2650 (N_2650,N_2382,N_2186);
nand U2651 (N_2651,N_2155,N_2215);
and U2652 (N_2652,N_2106,N_2213);
nand U2653 (N_2653,N_2139,N_2166);
and U2654 (N_2654,N_2144,N_2200);
xor U2655 (N_2655,N_2324,N_2263);
xnor U2656 (N_2656,N_2209,N_2396);
and U2657 (N_2657,N_2233,N_2266);
nor U2658 (N_2658,N_2231,N_2131);
nand U2659 (N_2659,N_2104,N_2126);
or U2660 (N_2660,N_2364,N_2302);
or U2661 (N_2661,N_2236,N_2291);
and U2662 (N_2662,N_2352,N_2214);
nor U2663 (N_2663,N_2233,N_2115);
or U2664 (N_2664,N_2199,N_2344);
and U2665 (N_2665,N_2201,N_2212);
and U2666 (N_2666,N_2277,N_2394);
or U2667 (N_2667,N_2213,N_2163);
nand U2668 (N_2668,N_2251,N_2156);
nor U2669 (N_2669,N_2173,N_2346);
nand U2670 (N_2670,N_2220,N_2375);
and U2671 (N_2671,N_2373,N_2386);
or U2672 (N_2672,N_2176,N_2175);
nor U2673 (N_2673,N_2165,N_2274);
or U2674 (N_2674,N_2192,N_2325);
xor U2675 (N_2675,N_2284,N_2255);
xor U2676 (N_2676,N_2296,N_2231);
and U2677 (N_2677,N_2119,N_2120);
or U2678 (N_2678,N_2154,N_2236);
xor U2679 (N_2679,N_2165,N_2391);
and U2680 (N_2680,N_2283,N_2245);
nor U2681 (N_2681,N_2290,N_2125);
xnor U2682 (N_2682,N_2271,N_2208);
nor U2683 (N_2683,N_2332,N_2339);
nand U2684 (N_2684,N_2162,N_2297);
or U2685 (N_2685,N_2188,N_2162);
nand U2686 (N_2686,N_2228,N_2391);
nor U2687 (N_2687,N_2342,N_2363);
and U2688 (N_2688,N_2212,N_2119);
or U2689 (N_2689,N_2359,N_2245);
nand U2690 (N_2690,N_2331,N_2288);
and U2691 (N_2691,N_2126,N_2224);
or U2692 (N_2692,N_2185,N_2327);
xnor U2693 (N_2693,N_2330,N_2115);
nor U2694 (N_2694,N_2168,N_2219);
nand U2695 (N_2695,N_2225,N_2265);
or U2696 (N_2696,N_2395,N_2283);
and U2697 (N_2697,N_2111,N_2199);
nor U2698 (N_2698,N_2334,N_2387);
or U2699 (N_2699,N_2147,N_2230);
and U2700 (N_2700,N_2634,N_2469);
nand U2701 (N_2701,N_2637,N_2658);
xnor U2702 (N_2702,N_2597,N_2654);
nand U2703 (N_2703,N_2424,N_2480);
nand U2704 (N_2704,N_2483,N_2601);
and U2705 (N_2705,N_2496,N_2416);
xnor U2706 (N_2706,N_2673,N_2514);
or U2707 (N_2707,N_2632,N_2580);
xor U2708 (N_2708,N_2573,N_2524);
nand U2709 (N_2709,N_2608,N_2593);
or U2710 (N_2710,N_2418,N_2607);
and U2711 (N_2711,N_2436,N_2428);
or U2712 (N_2712,N_2663,N_2513);
nor U2713 (N_2713,N_2525,N_2405);
nand U2714 (N_2714,N_2445,N_2693);
nor U2715 (N_2715,N_2472,N_2556);
or U2716 (N_2716,N_2578,N_2511);
nor U2717 (N_2717,N_2498,N_2434);
xor U2718 (N_2718,N_2686,N_2542);
xnor U2719 (N_2719,N_2596,N_2543);
nor U2720 (N_2720,N_2583,N_2629);
nor U2721 (N_2721,N_2660,N_2651);
and U2722 (N_2722,N_2554,N_2550);
xor U2723 (N_2723,N_2640,N_2467);
nand U2724 (N_2724,N_2653,N_2444);
or U2725 (N_2725,N_2455,N_2615);
or U2726 (N_2726,N_2547,N_2666);
nor U2727 (N_2727,N_2588,N_2476);
or U2728 (N_2728,N_2628,N_2645);
nor U2729 (N_2729,N_2675,N_2491);
nor U2730 (N_2730,N_2574,N_2562);
nand U2731 (N_2731,N_2423,N_2544);
nand U2732 (N_2732,N_2517,N_2681);
and U2733 (N_2733,N_2477,N_2478);
and U2734 (N_2734,N_2523,N_2410);
nand U2735 (N_2735,N_2457,N_2501);
xor U2736 (N_2736,N_2603,N_2443);
nand U2737 (N_2737,N_2420,N_2594);
and U2738 (N_2738,N_2407,N_2479);
nor U2739 (N_2739,N_2426,N_2448);
nand U2740 (N_2740,N_2633,N_2577);
nand U2741 (N_2741,N_2493,N_2571);
and U2742 (N_2742,N_2538,N_2452);
or U2743 (N_2743,N_2635,N_2412);
nand U2744 (N_2744,N_2485,N_2581);
or U2745 (N_2745,N_2529,N_2599);
nor U2746 (N_2746,N_2647,N_2429);
xor U2747 (N_2747,N_2585,N_2546);
nand U2748 (N_2748,N_2572,N_2464);
or U2749 (N_2749,N_2674,N_2606);
nand U2750 (N_2750,N_2459,N_2430);
or U2751 (N_2751,N_2619,N_2497);
or U2752 (N_2752,N_2453,N_2520);
nand U2753 (N_2753,N_2522,N_2516);
nand U2754 (N_2754,N_2694,N_2563);
xor U2755 (N_2755,N_2463,N_2630);
and U2756 (N_2756,N_2460,N_2421);
nand U2757 (N_2757,N_2521,N_2440);
and U2758 (N_2758,N_2609,N_2468);
or U2759 (N_2759,N_2617,N_2564);
nand U2760 (N_2760,N_2613,N_2639);
and U2761 (N_2761,N_2665,N_2605);
and U2762 (N_2762,N_2624,N_2502);
and U2763 (N_2763,N_2671,N_2655);
or U2764 (N_2764,N_2614,N_2489);
and U2765 (N_2765,N_2536,N_2461);
nor U2766 (N_2766,N_2621,N_2403);
or U2767 (N_2767,N_2569,N_2692);
and U2768 (N_2768,N_2549,N_2431);
or U2769 (N_2769,N_2490,N_2600);
nand U2770 (N_2770,N_2670,N_2518);
nand U2771 (N_2771,N_2618,N_2551);
nand U2772 (N_2772,N_2406,N_2508);
nor U2773 (N_2773,N_2512,N_2507);
or U2774 (N_2774,N_2540,N_2537);
and U2775 (N_2775,N_2591,N_2590);
nand U2776 (N_2776,N_2503,N_2611);
and U2777 (N_2777,N_2557,N_2530);
or U2778 (N_2778,N_2539,N_2659);
or U2779 (N_2779,N_2528,N_2450);
or U2780 (N_2780,N_2565,N_2417);
nor U2781 (N_2781,N_2589,N_2495);
and U2782 (N_2782,N_2570,N_2648);
or U2783 (N_2783,N_2641,N_2610);
or U2784 (N_2784,N_2494,N_2533);
or U2785 (N_2785,N_2698,N_2622);
nand U2786 (N_2786,N_2462,N_2553);
or U2787 (N_2787,N_2439,N_2531);
and U2788 (N_2788,N_2561,N_2470);
or U2789 (N_2789,N_2656,N_2587);
nand U2790 (N_2790,N_2555,N_2499);
xnor U2791 (N_2791,N_2643,N_2612);
or U2792 (N_2792,N_2471,N_2438);
nand U2793 (N_2793,N_2620,N_2447);
or U2794 (N_2794,N_2481,N_2402);
or U2795 (N_2795,N_2636,N_2576);
or U2796 (N_2796,N_2638,N_2487);
nand U2797 (N_2797,N_2650,N_2408);
nor U2798 (N_2798,N_2400,N_2696);
nor U2799 (N_2799,N_2482,N_2672);
or U2800 (N_2800,N_2486,N_2466);
nor U2801 (N_2801,N_2646,N_2527);
nor U2802 (N_2802,N_2560,N_2644);
nand U2803 (N_2803,N_2682,N_2678);
and U2804 (N_2804,N_2454,N_2676);
or U2805 (N_2805,N_2515,N_2579);
nand U2806 (N_2806,N_2433,N_2506);
nand U2807 (N_2807,N_2680,N_2432);
and U2808 (N_2808,N_2474,N_2567);
nand U2809 (N_2809,N_2598,N_2584);
and U2810 (N_2810,N_2697,N_2484);
xnor U2811 (N_2811,N_2534,N_2669);
and U2812 (N_2812,N_2409,N_2510);
and U2813 (N_2813,N_2558,N_2566);
or U2814 (N_2814,N_2685,N_2526);
or U2815 (N_2815,N_2575,N_2552);
nor U2816 (N_2816,N_2582,N_2652);
xnor U2817 (N_2817,N_2642,N_2427);
xnor U2818 (N_2818,N_2422,N_2602);
nand U2819 (N_2819,N_2616,N_2662);
or U2820 (N_2820,N_2592,N_2441);
xor U2821 (N_2821,N_2488,N_2519);
nand U2822 (N_2822,N_2411,N_2419);
or U2823 (N_2823,N_2492,N_2689);
and U2824 (N_2824,N_2683,N_2509);
or U2825 (N_2825,N_2437,N_2541);
nand U2826 (N_2826,N_2442,N_2649);
or U2827 (N_2827,N_2456,N_2404);
xnor U2828 (N_2828,N_2623,N_2661);
xor U2829 (N_2829,N_2668,N_2690);
nand U2830 (N_2830,N_2415,N_2500);
nor U2831 (N_2831,N_2449,N_2679);
and U2832 (N_2832,N_2667,N_2446);
xnor U2833 (N_2833,N_2699,N_2532);
xor U2834 (N_2834,N_2631,N_2473);
xor U2835 (N_2835,N_2664,N_2505);
xnor U2836 (N_2836,N_2687,N_2695);
nand U2837 (N_2837,N_2458,N_2451);
or U2838 (N_2838,N_2604,N_2627);
nand U2839 (N_2839,N_2677,N_2568);
nor U2840 (N_2840,N_2535,N_2684);
and U2841 (N_2841,N_2548,N_2413);
nor U2842 (N_2842,N_2559,N_2691);
nor U2843 (N_2843,N_2465,N_2475);
xor U2844 (N_2844,N_2586,N_2657);
xor U2845 (N_2845,N_2425,N_2625);
nor U2846 (N_2846,N_2401,N_2504);
and U2847 (N_2847,N_2414,N_2545);
and U2848 (N_2848,N_2626,N_2435);
xor U2849 (N_2849,N_2688,N_2595);
and U2850 (N_2850,N_2433,N_2497);
and U2851 (N_2851,N_2495,N_2461);
and U2852 (N_2852,N_2499,N_2646);
or U2853 (N_2853,N_2415,N_2627);
or U2854 (N_2854,N_2696,N_2564);
nand U2855 (N_2855,N_2670,N_2520);
or U2856 (N_2856,N_2417,N_2583);
xor U2857 (N_2857,N_2471,N_2589);
nor U2858 (N_2858,N_2416,N_2678);
nand U2859 (N_2859,N_2450,N_2501);
nor U2860 (N_2860,N_2453,N_2588);
xor U2861 (N_2861,N_2411,N_2557);
and U2862 (N_2862,N_2511,N_2449);
or U2863 (N_2863,N_2452,N_2617);
and U2864 (N_2864,N_2667,N_2461);
or U2865 (N_2865,N_2432,N_2627);
or U2866 (N_2866,N_2471,N_2694);
nor U2867 (N_2867,N_2524,N_2644);
and U2868 (N_2868,N_2540,N_2632);
or U2869 (N_2869,N_2615,N_2627);
nand U2870 (N_2870,N_2499,N_2564);
nor U2871 (N_2871,N_2510,N_2491);
nand U2872 (N_2872,N_2656,N_2536);
xor U2873 (N_2873,N_2513,N_2456);
or U2874 (N_2874,N_2453,N_2526);
or U2875 (N_2875,N_2628,N_2545);
xor U2876 (N_2876,N_2628,N_2666);
and U2877 (N_2877,N_2660,N_2588);
or U2878 (N_2878,N_2586,N_2444);
and U2879 (N_2879,N_2575,N_2415);
or U2880 (N_2880,N_2409,N_2474);
nor U2881 (N_2881,N_2665,N_2461);
nand U2882 (N_2882,N_2687,N_2566);
nand U2883 (N_2883,N_2625,N_2416);
nor U2884 (N_2884,N_2534,N_2495);
xnor U2885 (N_2885,N_2669,N_2685);
nand U2886 (N_2886,N_2567,N_2435);
nand U2887 (N_2887,N_2594,N_2652);
or U2888 (N_2888,N_2573,N_2432);
or U2889 (N_2889,N_2427,N_2441);
and U2890 (N_2890,N_2659,N_2651);
xor U2891 (N_2891,N_2493,N_2542);
nor U2892 (N_2892,N_2514,N_2493);
nand U2893 (N_2893,N_2431,N_2464);
xor U2894 (N_2894,N_2413,N_2697);
xnor U2895 (N_2895,N_2528,N_2593);
nor U2896 (N_2896,N_2630,N_2495);
nand U2897 (N_2897,N_2638,N_2465);
and U2898 (N_2898,N_2457,N_2660);
and U2899 (N_2899,N_2661,N_2637);
xnor U2900 (N_2900,N_2652,N_2515);
nor U2901 (N_2901,N_2523,N_2572);
or U2902 (N_2902,N_2624,N_2592);
or U2903 (N_2903,N_2524,N_2686);
nor U2904 (N_2904,N_2644,N_2551);
xor U2905 (N_2905,N_2454,N_2616);
nand U2906 (N_2906,N_2483,N_2429);
nand U2907 (N_2907,N_2406,N_2552);
and U2908 (N_2908,N_2662,N_2551);
xnor U2909 (N_2909,N_2678,N_2535);
or U2910 (N_2910,N_2485,N_2564);
or U2911 (N_2911,N_2606,N_2422);
and U2912 (N_2912,N_2457,N_2619);
xnor U2913 (N_2913,N_2559,N_2516);
nor U2914 (N_2914,N_2550,N_2468);
nand U2915 (N_2915,N_2631,N_2552);
or U2916 (N_2916,N_2696,N_2655);
nand U2917 (N_2917,N_2401,N_2590);
nor U2918 (N_2918,N_2423,N_2458);
and U2919 (N_2919,N_2620,N_2699);
nand U2920 (N_2920,N_2509,N_2437);
or U2921 (N_2921,N_2517,N_2540);
and U2922 (N_2922,N_2438,N_2597);
nor U2923 (N_2923,N_2652,N_2463);
nand U2924 (N_2924,N_2409,N_2438);
or U2925 (N_2925,N_2529,N_2458);
nor U2926 (N_2926,N_2495,N_2691);
nor U2927 (N_2927,N_2414,N_2648);
or U2928 (N_2928,N_2692,N_2698);
xor U2929 (N_2929,N_2527,N_2461);
nor U2930 (N_2930,N_2450,N_2601);
nand U2931 (N_2931,N_2411,N_2660);
nand U2932 (N_2932,N_2599,N_2426);
or U2933 (N_2933,N_2411,N_2628);
nor U2934 (N_2934,N_2414,N_2484);
or U2935 (N_2935,N_2565,N_2453);
nand U2936 (N_2936,N_2493,N_2509);
or U2937 (N_2937,N_2449,N_2654);
xnor U2938 (N_2938,N_2559,N_2477);
xor U2939 (N_2939,N_2427,N_2663);
nor U2940 (N_2940,N_2415,N_2588);
or U2941 (N_2941,N_2407,N_2405);
nor U2942 (N_2942,N_2518,N_2478);
xor U2943 (N_2943,N_2512,N_2462);
nor U2944 (N_2944,N_2432,N_2609);
and U2945 (N_2945,N_2472,N_2447);
or U2946 (N_2946,N_2483,N_2696);
nand U2947 (N_2947,N_2644,N_2542);
and U2948 (N_2948,N_2483,N_2612);
nor U2949 (N_2949,N_2490,N_2511);
xor U2950 (N_2950,N_2602,N_2647);
and U2951 (N_2951,N_2453,N_2425);
nor U2952 (N_2952,N_2584,N_2414);
nor U2953 (N_2953,N_2606,N_2525);
and U2954 (N_2954,N_2476,N_2647);
or U2955 (N_2955,N_2500,N_2600);
and U2956 (N_2956,N_2680,N_2507);
and U2957 (N_2957,N_2523,N_2591);
xnor U2958 (N_2958,N_2408,N_2639);
nand U2959 (N_2959,N_2513,N_2628);
xor U2960 (N_2960,N_2538,N_2508);
xnor U2961 (N_2961,N_2578,N_2572);
and U2962 (N_2962,N_2536,N_2694);
nand U2963 (N_2963,N_2451,N_2486);
nor U2964 (N_2964,N_2542,N_2457);
and U2965 (N_2965,N_2697,N_2565);
xnor U2966 (N_2966,N_2692,N_2497);
and U2967 (N_2967,N_2554,N_2616);
nor U2968 (N_2968,N_2660,N_2550);
xnor U2969 (N_2969,N_2434,N_2590);
or U2970 (N_2970,N_2569,N_2521);
and U2971 (N_2971,N_2516,N_2549);
and U2972 (N_2972,N_2556,N_2483);
and U2973 (N_2973,N_2571,N_2615);
nor U2974 (N_2974,N_2474,N_2443);
nor U2975 (N_2975,N_2442,N_2679);
nor U2976 (N_2976,N_2490,N_2572);
nand U2977 (N_2977,N_2634,N_2541);
and U2978 (N_2978,N_2699,N_2409);
and U2979 (N_2979,N_2578,N_2460);
xor U2980 (N_2980,N_2621,N_2599);
nand U2981 (N_2981,N_2623,N_2469);
or U2982 (N_2982,N_2499,N_2479);
xnor U2983 (N_2983,N_2452,N_2634);
and U2984 (N_2984,N_2508,N_2577);
or U2985 (N_2985,N_2614,N_2643);
and U2986 (N_2986,N_2469,N_2599);
or U2987 (N_2987,N_2503,N_2548);
or U2988 (N_2988,N_2554,N_2484);
or U2989 (N_2989,N_2447,N_2465);
xnor U2990 (N_2990,N_2526,N_2506);
or U2991 (N_2991,N_2536,N_2434);
nand U2992 (N_2992,N_2696,N_2668);
nand U2993 (N_2993,N_2516,N_2677);
xnor U2994 (N_2994,N_2662,N_2428);
nor U2995 (N_2995,N_2467,N_2405);
or U2996 (N_2996,N_2436,N_2419);
xnor U2997 (N_2997,N_2683,N_2644);
nand U2998 (N_2998,N_2614,N_2648);
and U2999 (N_2999,N_2455,N_2494);
or U3000 (N_3000,N_2860,N_2882);
nand U3001 (N_3001,N_2734,N_2879);
nand U3002 (N_3002,N_2975,N_2833);
or U3003 (N_3003,N_2985,N_2876);
and U3004 (N_3004,N_2793,N_2867);
xor U3005 (N_3005,N_2785,N_2900);
xnor U3006 (N_3006,N_2792,N_2957);
or U3007 (N_3007,N_2708,N_2883);
nor U3008 (N_3008,N_2790,N_2930);
or U3009 (N_3009,N_2732,N_2722);
nand U3010 (N_3010,N_2786,N_2920);
nand U3011 (N_3011,N_2953,N_2962);
xor U3012 (N_3012,N_2949,N_2841);
nor U3013 (N_3013,N_2801,N_2795);
nand U3014 (N_3014,N_2807,N_2764);
and U3015 (N_3015,N_2846,N_2817);
and U3016 (N_3016,N_2973,N_2948);
xnor U3017 (N_3017,N_2947,N_2946);
or U3018 (N_3018,N_2791,N_2735);
nor U3019 (N_3019,N_2713,N_2877);
nor U3020 (N_3020,N_2970,N_2972);
or U3021 (N_3021,N_2851,N_2995);
nor U3022 (N_3022,N_2963,N_2733);
nand U3023 (N_3023,N_2884,N_2840);
nor U3024 (N_3024,N_2895,N_2951);
nor U3025 (N_3025,N_2940,N_2777);
and U3026 (N_3026,N_2784,N_2829);
nand U3027 (N_3027,N_2767,N_2835);
nor U3028 (N_3028,N_2982,N_2950);
nand U3029 (N_3029,N_2754,N_2766);
xor U3030 (N_3030,N_2988,N_2744);
nand U3031 (N_3031,N_2944,N_2991);
xnor U3032 (N_3032,N_2816,N_2745);
xnor U3033 (N_3033,N_2709,N_2740);
and U3034 (N_3034,N_2729,N_2704);
or U3035 (N_3035,N_2700,N_2756);
or U3036 (N_3036,N_2936,N_2892);
or U3037 (N_3037,N_2911,N_2986);
nand U3038 (N_3038,N_2978,N_2716);
nand U3039 (N_3039,N_2937,N_2712);
and U3040 (N_3040,N_2894,N_2815);
and U3041 (N_3041,N_2763,N_2871);
xnor U3042 (N_3042,N_2913,N_2703);
or U3043 (N_3043,N_2862,N_2711);
and U3044 (N_3044,N_2872,N_2897);
nor U3045 (N_3045,N_2959,N_2902);
and U3046 (N_3046,N_2954,N_2910);
xnor U3047 (N_3047,N_2917,N_2701);
and U3048 (N_3048,N_2852,N_2811);
nand U3049 (N_3049,N_2746,N_2934);
and U3050 (N_3050,N_2865,N_2819);
xnor U3051 (N_3051,N_2783,N_2706);
or U3052 (N_3052,N_2886,N_2908);
or U3053 (N_3053,N_2771,N_2859);
or U3054 (N_3054,N_2762,N_2845);
xor U3055 (N_3055,N_2922,N_2915);
nor U3056 (N_3056,N_2775,N_2820);
and U3057 (N_3057,N_2893,N_2813);
nor U3058 (N_3058,N_2905,N_2822);
and U3059 (N_3059,N_2823,N_2943);
xor U3060 (N_3060,N_2739,N_2914);
xor U3061 (N_3061,N_2728,N_2945);
and U3062 (N_3062,N_2904,N_2929);
xor U3063 (N_3063,N_2921,N_2768);
xor U3064 (N_3064,N_2864,N_2989);
and U3065 (N_3065,N_2715,N_2899);
or U3066 (N_3066,N_2750,N_2942);
or U3067 (N_3067,N_2818,N_2774);
and U3068 (N_3068,N_2993,N_2858);
nand U3069 (N_3069,N_2848,N_2842);
nor U3070 (N_3070,N_2891,N_2977);
nor U3071 (N_3071,N_2887,N_2778);
or U3072 (N_3072,N_2743,N_2889);
xor U3073 (N_3073,N_2997,N_2724);
or U3074 (N_3074,N_2810,N_2702);
xor U3075 (N_3075,N_2738,N_2799);
or U3076 (N_3076,N_2832,N_2881);
nor U3077 (N_3077,N_2961,N_2866);
and U3078 (N_3078,N_2853,N_2916);
nand U3079 (N_3079,N_2971,N_2798);
nor U3080 (N_3080,N_2759,N_2797);
and U3081 (N_3081,N_2907,N_2751);
or U3082 (N_3082,N_2955,N_2870);
and U3083 (N_3083,N_2834,N_2965);
xnor U3084 (N_3084,N_2938,N_2760);
nor U3085 (N_3085,N_2773,N_2794);
and U3086 (N_3086,N_2981,N_2976);
nor U3087 (N_3087,N_2836,N_2974);
xor U3088 (N_3088,N_2928,N_2726);
nor U3089 (N_3089,N_2721,N_2931);
nor U3090 (N_3090,N_2939,N_2839);
and U3091 (N_3091,N_2847,N_2863);
xnor U3092 (N_3092,N_2748,N_2987);
xor U3093 (N_3093,N_2855,N_2838);
and U3094 (N_3094,N_2901,N_2952);
nand U3095 (N_3095,N_2898,N_2979);
or U3096 (N_3096,N_2873,N_2812);
or U3097 (N_3097,N_2753,N_2933);
nor U3098 (N_3098,N_2776,N_2923);
or U3099 (N_3099,N_2875,N_2806);
and U3100 (N_3100,N_2789,N_2805);
nor U3101 (N_3101,N_2856,N_2723);
nand U3102 (N_3102,N_2837,N_2935);
nand U3103 (N_3103,N_2919,N_2958);
nand U3104 (N_3104,N_2868,N_2737);
nand U3105 (N_3105,N_2966,N_2741);
nor U3106 (N_3106,N_2990,N_2969);
nand U3107 (N_3107,N_2999,N_2808);
nor U3108 (N_3108,N_2828,N_2720);
or U3109 (N_3109,N_2731,N_2827);
nor U3110 (N_3110,N_2826,N_2824);
or U3111 (N_3111,N_2821,N_2850);
nor U3112 (N_3112,N_2781,N_2718);
nor U3113 (N_3113,N_2742,N_2924);
and U3114 (N_3114,N_2968,N_2941);
or U3115 (N_3115,N_2926,N_2869);
nor U3116 (N_3116,N_2725,N_2757);
xor U3117 (N_3117,N_2727,N_2903);
nand U3118 (N_3118,N_2927,N_2730);
xor U3119 (N_3119,N_2996,N_2849);
or U3120 (N_3120,N_2752,N_2747);
nor U3121 (N_3121,N_2854,N_2994);
and U3122 (N_3122,N_2890,N_2814);
nor U3123 (N_3123,N_2984,N_2885);
xor U3124 (N_3124,N_2772,N_2809);
nand U3125 (N_3125,N_2918,N_2831);
nand U3126 (N_3126,N_2705,N_2906);
or U3127 (N_3127,N_2758,N_2909);
or U3128 (N_3128,N_2717,N_2874);
nand U3129 (N_3129,N_2878,N_2857);
and U3130 (N_3130,N_2719,N_2992);
nand U3131 (N_3131,N_2749,N_2779);
nand U3132 (N_3132,N_2761,N_2800);
or U3133 (N_3133,N_2714,N_2964);
nor U3134 (N_3134,N_2925,N_2998);
nor U3135 (N_3135,N_2912,N_2787);
nor U3136 (N_3136,N_2788,N_2825);
or U3137 (N_3137,N_2888,N_2736);
nor U3138 (N_3138,N_2861,N_2803);
and U3139 (N_3139,N_2770,N_2844);
or U3140 (N_3140,N_2880,N_2967);
nor U3141 (N_3141,N_2802,N_2765);
and U3142 (N_3142,N_2796,N_2843);
xnor U3143 (N_3143,N_2896,N_2710);
xnor U3144 (N_3144,N_2804,N_2769);
xor U3145 (N_3145,N_2983,N_2932);
or U3146 (N_3146,N_2780,N_2956);
xnor U3147 (N_3147,N_2830,N_2755);
nor U3148 (N_3148,N_2707,N_2782);
xor U3149 (N_3149,N_2980,N_2960);
xnor U3150 (N_3150,N_2757,N_2924);
xnor U3151 (N_3151,N_2788,N_2706);
nand U3152 (N_3152,N_2853,N_2951);
xor U3153 (N_3153,N_2858,N_2944);
nor U3154 (N_3154,N_2783,N_2945);
or U3155 (N_3155,N_2816,N_2718);
or U3156 (N_3156,N_2848,N_2874);
nand U3157 (N_3157,N_2883,N_2809);
xnor U3158 (N_3158,N_2920,N_2840);
nand U3159 (N_3159,N_2972,N_2959);
nor U3160 (N_3160,N_2965,N_2760);
nand U3161 (N_3161,N_2842,N_2786);
nor U3162 (N_3162,N_2943,N_2850);
nand U3163 (N_3163,N_2932,N_2895);
nand U3164 (N_3164,N_2874,N_2900);
nand U3165 (N_3165,N_2929,N_2896);
or U3166 (N_3166,N_2934,N_2735);
or U3167 (N_3167,N_2731,N_2836);
or U3168 (N_3168,N_2858,N_2719);
and U3169 (N_3169,N_2853,N_2710);
xnor U3170 (N_3170,N_2701,N_2804);
nor U3171 (N_3171,N_2726,N_2790);
nand U3172 (N_3172,N_2763,N_2990);
or U3173 (N_3173,N_2892,N_2977);
and U3174 (N_3174,N_2704,N_2871);
nand U3175 (N_3175,N_2791,N_2886);
and U3176 (N_3176,N_2909,N_2870);
and U3177 (N_3177,N_2941,N_2794);
xnor U3178 (N_3178,N_2887,N_2829);
xor U3179 (N_3179,N_2913,N_2957);
and U3180 (N_3180,N_2875,N_2789);
nor U3181 (N_3181,N_2897,N_2782);
nor U3182 (N_3182,N_2809,N_2846);
nand U3183 (N_3183,N_2719,N_2818);
xor U3184 (N_3184,N_2701,N_2905);
nand U3185 (N_3185,N_2993,N_2981);
nand U3186 (N_3186,N_2825,N_2966);
nand U3187 (N_3187,N_2762,N_2957);
nor U3188 (N_3188,N_2747,N_2955);
and U3189 (N_3189,N_2758,N_2938);
or U3190 (N_3190,N_2717,N_2843);
nor U3191 (N_3191,N_2937,N_2999);
xor U3192 (N_3192,N_2734,N_2725);
nor U3193 (N_3193,N_2760,N_2890);
nand U3194 (N_3194,N_2738,N_2917);
nand U3195 (N_3195,N_2705,N_2785);
nor U3196 (N_3196,N_2979,N_2766);
nor U3197 (N_3197,N_2722,N_2984);
or U3198 (N_3198,N_2927,N_2806);
xor U3199 (N_3199,N_2713,N_2795);
xnor U3200 (N_3200,N_2714,N_2913);
nor U3201 (N_3201,N_2987,N_2965);
nor U3202 (N_3202,N_2979,N_2721);
nand U3203 (N_3203,N_2936,N_2769);
nand U3204 (N_3204,N_2700,N_2988);
xnor U3205 (N_3205,N_2711,N_2874);
nor U3206 (N_3206,N_2798,N_2871);
xnor U3207 (N_3207,N_2780,N_2853);
nor U3208 (N_3208,N_2804,N_2993);
xnor U3209 (N_3209,N_2709,N_2728);
nand U3210 (N_3210,N_2818,N_2732);
or U3211 (N_3211,N_2814,N_2940);
nand U3212 (N_3212,N_2811,N_2982);
xnor U3213 (N_3213,N_2906,N_2841);
nand U3214 (N_3214,N_2941,N_2883);
xor U3215 (N_3215,N_2953,N_2735);
xnor U3216 (N_3216,N_2827,N_2971);
or U3217 (N_3217,N_2829,N_2881);
or U3218 (N_3218,N_2752,N_2978);
or U3219 (N_3219,N_2761,N_2816);
or U3220 (N_3220,N_2792,N_2721);
and U3221 (N_3221,N_2942,N_2789);
or U3222 (N_3222,N_2706,N_2845);
nor U3223 (N_3223,N_2797,N_2957);
xnor U3224 (N_3224,N_2834,N_2739);
xor U3225 (N_3225,N_2724,N_2925);
nand U3226 (N_3226,N_2707,N_2736);
nand U3227 (N_3227,N_2914,N_2830);
nor U3228 (N_3228,N_2930,N_2977);
nor U3229 (N_3229,N_2713,N_2834);
nand U3230 (N_3230,N_2979,N_2946);
xnor U3231 (N_3231,N_2973,N_2788);
xor U3232 (N_3232,N_2829,N_2860);
nor U3233 (N_3233,N_2819,N_2786);
nand U3234 (N_3234,N_2755,N_2715);
or U3235 (N_3235,N_2916,N_2805);
nor U3236 (N_3236,N_2826,N_2724);
xor U3237 (N_3237,N_2777,N_2743);
or U3238 (N_3238,N_2869,N_2773);
or U3239 (N_3239,N_2804,N_2755);
xnor U3240 (N_3240,N_2863,N_2895);
xnor U3241 (N_3241,N_2778,N_2982);
or U3242 (N_3242,N_2950,N_2703);
and U3243 (N_3243,N_2786,N_2764);
nor U3244 (N_3244,N_2926,N_2846);
and U3245 (N_3245,N_2738,N_2767);
xor U3246 (N_3246,N_2809,N_2983);
xnor U3247 (N_3247,N_2793,N_2861);
nor U3248 (N_3248,N_2869,N_2714);
xor U3249 (N_3249,N_2907,N_2845);
nand U3250 (N_3250,N_2907,N_2712);
nor U3251 (N_3251,N_2760,N_2745);
and U3252 (N_3252,N_2939,N_2949);
xnor U3253 (N_3253,N_2783,N_2815);
or U3254 (N_3254,N_2918,N_2750);
or U3255 (N_3255,N_2818,N_2768);
or U3256 (N_3256,N_2780,N_2849);
xor U3257 (N_3257,N_2855,N_2865);
nand U3258 (N_3258,N_2835,N_2884);
nor U3259 (N_3259,N_2979,N_2780);
nor U3260 (N_3260,N_2803,N_2804);
xor U3261 (N_3261,N_2738,N_2873);
nand U3262 (N_3262,N_2974,N_2818);
and U3263 (N_3263,N_2875,N_2886);
xnor U3264 (N_3264,N_2892,N_2705);
and U3265 (N_3265,N_2922,N_2977);
or U3266 (N_3266,N_2856,N_2778);
and U3267 (N_3267,N_2852,N_2966);
and U3268 (N_3268,N_2916,N_2921);
or U3269 (N_3269,N_2881,N_2899);
xnor U3270 (N_3270,N_2865,N_2731);
or U3271 (N_3271,N_2943,N_2919);
or U3272 (N_3272,N_2931,N_2890);
xor U3273 (N_3273,N_2749,N_2819);
and U3274 (N_3274,N_2746,N_2794);
nor U3275 (N_3275,N_2780,N_2957);
nor U3276 (N_3276,N_2878,N_2883);
xnor U3277 (N_3277,N_2844,N_2987);
nor U3278 (N_3278,N_2730,N_2999);
xor U3279 (N_3279,N_2812,N_2726);
nor U3280 (N_3280,N_2965,N_2898);
xor U3281 (N_3281,N_2799,N_2789);
and U3282 (N_3282,N_2876,N_2833);
and U3283 (N_3283,N_2821,N_2749);
nand U3284 (N_3284,N_2707,N_2930);
nor U3285 (N_3285,N_2905,N_2947);
nor U3286 (N_3286,N_2907,N_2777);
and U3287 (N_3287,N_2954,N_2797);
xnor U3288 (N_3288,N_2865,N_2708);
nor U3289 (N_3289,N_2968,N_2853);
nand U3290 (N_3290,N_2865,N_2849);
nor U3291 (N_3291,N_2970,N_2830);
and U3292 (N_3292,N_2819,N_2845);
nor U3293 (N_3293,N_2817,N_2786);
nor U3294 (N_3294,N_2942,N_2759);
xnor U3295 (N_3295,N_2978,N_2938);
nand U3296 (N_3296,N_2794,N_2785);
and U3297 (N_3297,N_2832,N_2962);
nand U3298 (N_3298,N_2799,N_2808);
nand U3299 (N_3299,N_2765,N_2984);
xnor U3300 (N_3300,N_3212,N_3085);
or U3301 (N_3301,N_3299,N_3207);
nand U3302 (N_3302,N_3282,N_3252);
xor U3303 (N_3303,N_3167,N_3258);
nor U3304 (N_3304,N_3016,N_3022);
xnor U3305 (N_3305,N_3275,N_3191);
and U3306 (N_3306,N_3263,N_3053);
nor U3307 (N_3307,N_3195,N_3288);
nor U3308 (N_3308,N_3268,N_3209);
nand U3309 (N_3309,N_3074,N_3141);
or U3310 (N_3310,N_3208,N_3034);
nand U3311 (N_3311,N_3023,N_3246);
xor U3312 (N_3312,N_3111,N_3152);
nand U3313 (N_3313,N_3142,N_3079);
nand U3314 (N_3314,N_3230,N_3006);
nor U3315 (N_3315,N_3243,N_3291);
or U3316 (N_3316,N_3244,N_3251);
nor U3317 (N_3317,N_3180,N_3273);
nand U3318 (N_3318,N_3003,N_3179);
and U3319 (N_3319,N_3203,N_3098);
or U3320 (N_3320,N_3270,N_3158);
or U3321 (N_3321,N_3240,N_3118);
xor U3322 (N_3322,N_3174,N_3049);
and U3323 (N_3323,N_3025,N_3127);
or U3324 (N_3324,N_3095,N_3172);
nor U3325 (N_3325,N_3159,N_3238);
and U3326 (N_3326,N_3151,N_3130);
nor U3327 (N_3327,N_3271,N_3051);
or U3328 (N_3328,N_3120,N_3078);
xnor U3329 (N_3329,N_3285,N_3265);
and U3330 (N_3330,N_3287,N_3083);
xnor U3331 (N_3331,N_3002,N_3257);
or U3332 (N_3332,N_3232,N_3068);
nor U3333 (N_3333,N_3165,N_3280);
nor U3334 (N_3334,N_3055,N_3150);
nand U3335 (N_3335,N_3072,N_3201);
and U3336 (N_3336,N_3221,N_3235);
nand U3337 (N_3337,N_3071,N_3199);
or U3338 (N_3338,N_3057,N_3286);
and U3339 (N_3339,N_3135,N_3060);
nand U3340 (N_3340,N_3297,N_3149);
nor U3341 (N_3341,N_3117,N_3131);
or U3342 (N_3342,N_3121,N_3018);
or U3343 (N_3343,N_3234,N_3133);
nand U3344 (N_3344,N_3260,N_3178);
nor U3345 (N_3345,N_3219,N_3173);
nor U3346 (N_3346,N_3146,N_3043);
or U3347 (N_3347,N_3289,N_3254);
and U3348 (N_3348,N_3137,N_3169);
nand U3349 (N_3349,N_3292,N_3267);
or U3350 (N_3350,N_3013,N_3175);
or U3351 (N_3351,N_3164,N_3107);
xnor U3352 (N_3352,N_3272,N_3102);
xor U3353 (N_3353,N_3211,N_3274);
or U3354 (N_3354,N_3004,N_3226);
or U3355 (N_3355,N_3168,N_3124);
nand U3356 (N_3356,N_3281,N_3128);
nand U3357 (N_3357,N_3197,N_3253);
or U3358 (N_3358,N_3262,N_3024);
nand U3359 (N_3359,N_3157,N_3088);
or U3360 (N_3360,N_3198,N_3048);
and U3361 (N_3361,N_3113,N_3064);
nor U3362 (N_3362,N_3020,N_3224);
nand U3363 (N_3363,N_3105,N_3170);
xor U3364 (N_3364,N_3077,N_3223);
nor U3365 (N_3365,N_3041,N_3112);
nor U3366 (N_3366,N_3183,N_3070);
nor U3367 (N_3367,N_3248,N_3109);
nand U3368 (N_3368,N_3000,N_3063);
nor U3369 (N_3369,N_3233,N_3284);
nor U3370 (N_3370,N_3200,N_3047);
nor U3371 (N_3371,N_3269,N_3089);
xnor U3372 (N_3372,N_3249,N_3161);
xnor U3373 (N_3373,N_3144,N_3242);
nand U3374 (N_3374,N_3210,N_3217);
xor U3375 (N_3375,N_3011,N_3104);
and U3376 (N_3376,N_3277,N_3067);
nand U3377 (N_3377,N_3029,N_3103);
nor U3378 (N_3378,N_3114,N_3080);
and U3379 (N_3379,N_3163,N_3017);
nand U3380 (N_3380,N_3228,N_3215);
xor U3381 (N_3381,N_3247,N_3186);
or U3382 (N_3382,N_3036,N_3096);
nor U3383 (N_3383,N_3044,N_3190);
or U3384 (N_3384,N_3222,N_3184);
nand U3385 (N_3385,N_3194,N_3040);
nand U3386 (N_3386,N_3202,N_3166);
and U3387 (N_3387,N_3073,N_3290);
or U3388 (N_3388,N_3139,N_3028);
nand U3389 (N_3389,N_3143,N_3110);
and U3390 (N_3390,N_3213,N_3276);
nand U3391 (N_3391,N_3205,N_3059);
nand U3392 (N_3392,N_3256,N_3177);
nand U3393 (N_3393,N_3106,N_3065);
and U3394 (N_3394,N_3033,N_3032);
or U3395 (N_3395,N_3255,N_3237);
or U3396 (N_3396,N_3015,N_3192);
xnor U3397 (N_3397,N_3182,N_3241);
or U3398 (N_3398,N_3138,N_3039);
nand U3399 (N_3399,N_3081,N_3134);
nand U3400 (N_3400,N_3097,N_3160);
and U3401 (N_3401,N_3052,N_3091);
and U3402 (N_3402,N_3293,N_3101);
and U3403 (N_3403,N_3162,N_3126);
and U3404 (N_3404,N_3093,N_3136);
xor U3405 (N_3405,N_3094,N_3154);
nand U3406 (N_3406,N_3196,N_3031);
and U3407 (N_3407,N_3058,N_3075);
or U3408 (N_3408,N_3218,N_3122);
nand U3409 (N_3409,N_3129,N_3187);
nor U3410 (N_3410,N_3066,N_3239);
and U3411 (N_3411,N_3021,N_3019);
nor U3412 (N_3412,N_3092,N_3245);
or U3413 (N_3413,N_3185,N_3261);
or U3414 (N_3414,N_3278,N_3115);
and U3415 (N_3415,N_3132,N_3050);
nor U3416 (N_3416,N_3216,N_3119);
or U3417 (N_3417,N_3056,N_3227);
or U3418 (N_3418,N_3038,N_3027);
xnor U3419 (N_3419,N_3054,N_3294);
xor U3420 (N_3420,N_3231,N_3087);
xnor U3421 (N_3421,N_3153,N_3012);
nand U3422 (N_3422,N_3188,N_3014);
xor U3423 (N_3423,N_3259,N_3264);
and U3424 (N_3424,N_3099,N_3108);
nand U3425 (N_3425,N_3229,N_3062);
nor U3426 (N_3426,N_3155,N_3030);
or U3427 (N_3427,N_3147,N_3069);
xor U3428 (N_3428,N_3279,N_3061);
nand U3429 (N_3429,N_3171,N_3225);
nor U3430 (N_3430,N_3042,N_3100);
and U3431 (N_3431,N_3076,N_3045);
nor U3432 (N_3432,N_3035,N_3010);
nor U3433 (N_3433,N_3204,N_3283);
and U3434 (N_3434,N_3026,N_3295);
or U3435 (N_3435,N_3181,N_3266);
and U3436 (N_3436,N_3176,N_3193);
nand U3437 (N_3437,N_3250,N_3236);
and U3438 (N_3438,N_3206,N_3037);
or U3439 (N_3439,N_3220,N_3125);
or U3440 (N_3440,N_3086,N_3116);
nand U3441 (N_3441,N_3145,N_3214);
or U3442 (N_3442,N_3007,N_3296);
or U3443 (N_3443,N_3140,N_3001);
nand U3444 (N_3444,N_3123,N_3090);
xor U3445 (N_3445,N_3156,N_3084);
or U3446 (N_3446,N_3008,N_3082);
nor U3447 (N_3447,N_3005,N_3148);
xnor U3448 (N_3448,N_3189,N_3009);
nor U3449 (N_3449,N_3298,N_3046);
nand U3450 (N_3450,N_3067,N_3180);
xnor U3451 (N_3451,N_3053,N_3000);
or U3452 (N_3452,N_3125,N_3156);
xnor U3453 (N_3453,N_3081,N_3021);
or U3454 (N_3454,N_3254,N_3067);
nand U3455 (N_3455,N_3237,N_3256);
xor U3456 (N_3456,N_3225,N_3213);
nor U3457 (N_3457,N_3007,N_3294);
nand U3458 (N_3458,N_3154,N_3077);
and U3459 (N_3459,N_3130,N_3202);
xor U3460 (N_3460,N_3127,N_3110);
nand U3461 (N_3461,N_3193,N_3282);
xor U3462 (N_3462,N_3262,N_3123);
and U3463 (N_3463,N_3156,N_3291);
and U3464 (N_3464,N_3171,N_3178);
nand U3465 (N_3465,N_3123,N_3140);
xor U3466 (N_3466,N_3042,N_3262);
or U3467 (N_3467,N_3239,N_3143);
nand U3468 (N_3468,N_3291,N_3170);
nand U3469 (N_3469,N_3130,N_3192);
or U3470 (N_3470,N_3034,N_3120);
xnor U3471 (N_3471,N_3177,N_3278);
and U3472 (N_3472,N_3129,N_3101);
nor U3473 (N_3473,N_3064,N_3182);
or U3474 (N_3474,N_3104,N_3242);
or U3475 (N_3475,N_3134,N_3184);
or U3476 (N_3476,N_3051,N_3004);
nor U3477 (N_3477,N_3002,N_3039);
and U3478 (N_3478,N_3114,N_3146);
nor U3479 (N_3479,N_3276,N_3176);
or U3480 (N_3480,N_3178,N_3081);
nand U3481 (N_3481,N_3168,N_3257);
xnor U3482 (N_3482,N_3166,N_3160);
and U3483 (N_3483,N_3260,N_3112);
and U3484 (N_3484,N_3105,N_3262);
or U3485 (N_3485,N_3240,N_3129);
nor U3486 (N_3486,N_3094,N_3117);
xnor U3487 (N_3487,N_3224,N_3145);
or U3488 (N_3488,N_3147,N_3251);
xnor U3489 (N_3489,N_3174,N_3284);
and U3490 (N_3490,N_3141,N_3157);
and U3491 (N_3491,N_3061,N_3068);
nor U3492 (N_3492,N_3107,N_3175);
nand U3493 (N_3493,N_3198,N_3235);
nand U3494 (N_3494,N_3091,N_3291);
or U3495 (N_3495,N_3034,N_3271);
nand U3496 (N_3496,N_3093,N_3144);
or U3497 (N_3497,N_3174,N_3009);
nand U3498 (N_3498,N_3176,N_3192);
and U3499 (N_3499,N_3198,N_3169);
nor U3500 (N_3500,N_3011,N_3090);
or U3501 (N_3501,N_3181,N_3234);
xor U3502 (N_3502,N_3102,N_3191);
nor U3503 (N_3503,N_3219,N_3003);
and U3504 (N_3504,N_3044,N_3008);
or U3505 (N_3505,N_3158,N_3216);
xor U3506 (N_3506,N_3275,N_3168);
nand U3507 (N_3507,N_3189,N_3064);
and U3508 (N_3508,N_3131,N_3263);
xnor U3509 (N_3509,N_3163,N_3261);
nor U3510 (N_3510,N_3175,N_3150);
and U3511 (N_3511,N_3061,N_3218);
nand U3512 (N_3512,N_3285,N_3073);
xor U3513 (N_3513,N_3198,N_3224);
nor U3514 (N_3514,N_3125,N_3149);
xor U3515 (N_3515,N_3117,N_3166);
and U3516 (N_3516,N_3112,N_3120);
and U3517 (N_3517,N_3072,N_3015);
nor U3518 (N_3518,N_3277,N_3072);
nor U3519 (N_3519,N_3151,N_3258);
or U3520 (N_3520,N_3195,N_3008);
nor U3521 (N_3521,N_3210,N_3109);
xor U3522 (N_3522,N_3109,N_3048);
nor U3523 (N_3523,N_3050,N_3019);
xor U3524 (N_3524,N_3143,N_3009);
and U3525 (N_3525,N_3121,N_3138);
xnor U3526 (N_3526,N_3254,N_3064);
nand U3527 (N_3527,N_3174,N_3117);
xor U3528 (N_3528,N_3023,N_3028);
nor U3529 (N_3529,N_3286,N_3021);
or U3530 (N_3530,N_3088,N_3173);
or U3531 (N_3531,N_3196,N_3115);
xor U3532 (N_3532,N_3022,N_3127);
nand U3533 (N_3533,N_3265,N_3294);
or U3534 (N_3534,N_3070,N_3089);
or U3535 (N_3535,N_3206,N_3202);
or U3536 (N_3536,N_3236,N_3247);
xor U3537 (N_3537,N_3076,N_3259);
and U3538 (N_3538,N_3107,N_3296);
xor U3539 (N_3539,N_3295,N_3264);
or U3540 (N_3540,N_3247,N_3172);
xor U3541 (N_3541,N_3120,N_3179);
xor U3542 (N_3542,N_3072,N_3224);
or U3543 (N_3543,N_3255,N_3297);
or U3544 (N_3544,N_3205,N_3133);
xnor U3545 (N_3545,N_3191,N_3013);
and U3546 (N_3546,N_3141,N_3124);
or U3547 (N_3547,N_3147,N_3017);
nor U3548 (N_3548,N_3218,N_3198);
xor U3549 (N_3549,N_3116,N_3163);
nand U3550 (N_3550,N_3029,N_3132);
and U3551 (N_3551,N_3099,N_3276);
xor U3552 (N_3552,N_3260,N_3038);
nand U3553 (N_3553,N_3204,N_3152);
xor U3554 (N_3554,N_3184,N_3294);
and U3555 (N_3555,N_3222,N_3147);
nor U3556 (N_3556,N_3211,N_3245);
xor U3557 (N_3557,N_3268,N_3285);
xor U3558 (N_3558,N_3202,N_3105);
nor U3559 (N_3559,N_3010,N_3095);
nor U3560 (N_3560,N_3163,N_3038);
or U3561 (N_3561,N_3115,N_3111);
or U3562 (N_3562,N_3143,N_3242);
xnor U3563 (N_3563,N_3162,N_3061);
or U3564 (N_3564,N_3279,N_3121);
nor U3565 (N_3565,N_3075,N_3156);
nor U3566 (N_3566,N_3119,N_3221);
nand U3567 (N_3567,N_3283,N_3094);
nor U3568 (N_3568,N_3287,N_3050);
xnor U3569 (N_3569,N_3138,N_3065);
and U3570 (N_3570,N_3284,N_3064);
xnor U3571 (N_3571,N_3001,N_3296);
or U3572 (N_3572,N_3188,N_3251);
nand U3573 (N_3573,N_3294,N_3275);
and U3574 (N_3574,N_3155,N_3181);
and U3575 (N_3575,N_3238,N_3072);
xor U3576 (N_3576,N_3285,N_3237);
nor U3577 (N_3577,N_3121,N_3144);
and U3578 (N_3578,N_3087,N_3240);
nor U3579 (N_3579,N_3245,N_3296);
xnor U3580 (N_3580,N_3227,N_3032);
and U3581 (N_3581,N_3254,N_3131);
nand U3582 (N_3582,N_3293,N_3099);
nor U3583 (N_3583,N_3141,N_3230);
nand U3584 (N_3584,N_3079,N_3122);
nor U3585 (N_3585,N_3209,N_3257);
nand U3586 (N_3586,N_3173,N_3051);
or U3587 (N_3587,N_3239,N_3246);
or U3588 (N_3588,N_3051,N_3255);
nor U3589 (N_3589,N_3062,N_3093);
xnor U3590 (N_3590,N_3203,N_3055);
or U3591 (N_3591,N_3139,N_3062);
xnor U3592 (N_3592,N_3239,N_3033);
xnor U3593 (N_3593,N_3206,N_3262);
nand U3594 (N_3594,N_3120,N_3191);
or U3595 (N_3595,N_3076,N_3122);
or U3596 (N_3596,N_3278,N_3131);
or U3597 (N_3597,N_3193,N_3026);
or U3598 (N_3598,N_3160,N_3128);
and U3599 (N_3599,N_3031,N_3071);
and U3600 (N_3600,N_3444,N_3326);
and U3601 (N_3601,N_3565,N_3506);
and U3602 (N_3602,N_3507,N_3478);
or U3603 (N_3603,N_3396,N_3401);
xor U3604 (N_3604,N_3503,N_3447);
nand U3605 (N_3605,N_3422,N_3328);
and U3606 (N_3606,N_3314,N_3317);
and U3607 (N_3607,N_3388,N_3421);
or U3608 (N_3608,N_3410,N_3467);
nand U3609 (N_3609,N_3369,N_3389);
nor U3610 (N_3610,N_3553,N_3484);
or U3611 (N_3611,N_3549,N_3311);
or U3612 (N_3612,N_3350,N_3360);
nor U3613 (N_3613,N_3436,N_3552);
nand U3614 (N_3614,N_3312,N_3362);
xnor U3615 (N_3615,N_3351,N_3408);
xnor U3616 (N_3616,N_3569,N_3468);
and U3617 (N_3617,N_3572,N_3460);
or U3618 (N_3618,N_3409,N_3536);
or U3619 (N_3619,N_3425,N_3342);
or U3620 (N_3620,N_3516,N_3544);
or U3621 (N_3621,N_3511,N_3358);
nand U3622 (N_3622,N_3472,N_3331);
nor U3623 (N_3623,N_3598,N_3502);
or U3624 (N_3624,N_3435,N_3417);
xnor U3625 (N_3625,N_3533,N_3570);
and U3626 (N_3626,N_3325,N_3528);
nor U3627 (N_3627,N_3470,N_3587);
and U3628 (N_3628,N_3488,N_3466);
xor U3629 (N_3629,N_3461,N_3324);
and U3630 (N_3630,N_3306,N_3599);
nand U3631 (N_3631,N_3344,N_3474);
xnor U3632 (N_3632,N_3464,N_3449);
xor U3633 (N_3633,N_3525,N_3391);
xor U3634 (N_3634,N_3384,N_3547);
nor U3635 (N_3635,N_3302,N_3595);
xnor U3636 (N_3636,N_3578,N_3526);
xnor U3637 (N_3637,N_3404,N_3407);
or U3638 (N_3638,N_3381,N_3583);
or U3639 (N_3639,N_3495,N_3385);
and U3640 (N_3640,N_3482,N_3394);
or U3641 (N_3641,N_3367,N_3393);
and U3642 (N_3642,N_3487,N_3451);
or U3643 (N_3643,N_3305,N_3335);
or U3644 (N_3644,N_3441,N_3543);
xnor U3645 (N_3645,N_3522,N_3383);
or U3646 (N_3646,N_3450,N_3571);
nor U3647 (N_3647,N_3490,N_3392);
nand U3648 (N_3648,N_3555,N_3529);
nor U3649 (N_3649,N_3375,N_3568);
or U3650 (N_3650,N_3471,N_3557);
nand U3651 (N_3651,N_3581,N_3323);
nand U3652 (N_3652,N_3303,N_3534);
or U3653 (N_3653,N_3535,N_3395);
nand U3654 (N_3654,N_3315,N_3349);
or U3655 (N_3655,N_3531,N_3548);
xnor U3656 (N_3656,N_3343,N_3370);
xor U3657 (N_3657,N_3562,N_3517);
or U3658 (N_3658,N_3336,N_3428);
nor U3659 (N_3659,N_3424,N_3532);
or U3660 (N_3660,N_3413,N_3567);
and U3661 (N_3661,N_3469,N_3379);
xnor U3662 (N_3662,N_3513,N_3463);
xnor U3663 (N_3663,N_3418,N_3440);
nand U3664 (N_3664,N_3414,N_3426);
xor U3665 (N_3665,N_3398,N_3310);
xor U3666 (N_3666,N_3540,N_3319);
and U3667 (N_3667,N_3564,N_3432);
or U3668 (N_3668,N_3574,N_3445);
and U3669 (N_3669,N_3438,N_3594);
and U3670 (N_3670,N_3456,N_3596);
or U3671 (N_3671,N_3372,N_3521);
nand U3672 (N_3672,N_3420,N_3437);
nor U3673 (N_3673,N_3406,N_3486);
or U3674 (N_3674,N_3542,N_3419);
nor U3675 (N_3675,N_3476,N_3573);
xor U3676 (N_3676,N_3352,N_3356);
nand U3677 (N_3677,N_3537,N_3416);
and U3678 (N_3678,N_3374,N_3518);
nand U3679 (N_3679,N_3538,N_3320);
xnor U3680 (N_3680,N_3489,N_3546);
or U3681 (N_3681,N_3448,N_3399);
nand U3682 (N_3682,N_3558,N_3376);
nor U3683 (N_3683,N_3505,N_3365);
xor U3684 (N_3684,N_3316,N_3443);
nor U3685 (N_3685,N_3430,N_3459);
nand U3686 (N_3686,N_3566,N_3345);
xnor U3687 (N_3687,N_3353,N_3363);
nor U3688 (N_3688,N_3510,N_3504);
xor U3689 (N_3689,N_3499,N_3329);
xnor U3690 (N_3690,N_3318,N_3390);
and U3691 (N_3691,N_3597,N_3498);
and U3692 (N_3692,N_3588,N_3593);
nand U3693 (N_3693,N_3380,N_3494);
and U3694 (N_3694,N_3592,N_3366);
nand U3695 (N_3695,N_3551,N_3497);
and U3696 (N_3696,N_3584,N_3485);
nor U3697 (N_3697,N_3527,N_3338);
nor U3698 (N_3698,N_3477,N_3307);
or U3699 (N_3699,N_3403,N_3589);
nand U3700 (N_3700,N_3327,N_3541);
nand U3701 (N_3701,N_3411,N_3364);
or U3702 (N_3702,N_3465,N_3462);
nor U3703 (N_3703,N_3493,N_3304);
nor U3704 (N_3704,N_3378,N_3346);
nor U3705 (N_3705,N_3539,N_3330);
or U3706 (N_3706,N_3340,N_3301);
nor U3707 (N_3707,N_3341,N_3322);
nand U3708 (N_3708,N_3415,N_3508);
and U3709 (N_3709,N_3357,N_3579);
nand U3710 (N_3710,N_3429,N_3433);
and U3711 (N_3711,N_3530,N_3405);
and U3712 (N_3712,N_3492,N_3300);
and U3713 (N_3713,N_3586,N_3576);
or U3714 (N_3714,N_3455,N_3397);
and U3715 (N_3715,N_3355,N_3427);
or U3716 (N_3716,N_3509,N_3479);
xor U3717 (N_3717,N_3582,N_3458);
and U3718 (N_3718,N_3373,N_3585);
nand U3719 (N_3719,N_3563,N_3577);
xor U3720 (N_3720,N_3545,N_3519);
and U3721 (N_3721,N_3400,N_3308);
nor U3722 (N_3722,N_3514,N_3361);
nor U3723 (N_3723,N_3480,N_3309);
or U3724 (N_3724,N_3556,N_3491);
or U3725 (N_3725,N_3454,N_3386);
nand U3726 (N_3726,N_3554,N_3368);
and U3727 (N_3727,N_3377,N_3337);
xnor U3728 (N_3728,N_3560,N_3473);
nand U3729 (N_3729,N_3550,N_3431);
and U3730 (N_3730,N_3453,N_3334);
nor U3731 (N_3731,N_3457,N_3439);
or U3732 (N_3732,N_3501,N_3523);
nor U3733 (N_3733,N_3434,N_3496);
nor U3734 (N_3734,N_3483,N_3452);
and U3735 (N_3735,N_3575,N_3348);
or U3736 (N_3736,N_3500,N_3412);
nor U3737 (N_3737,N_3515,N_3332);
xor U3738 (N_3738,N_3481,N_3475);
and U3739 (N_3739,N_3512,N_3354);
nor U3740 (N_3740,N_3339,N_3590);
xnor U3741 (N_3741,N_3561,N_3580);
xor U3742 (N_3742,N_3520,N_3313);
nor U3743 (N_3743,N_3382,N_3359);
and U3744 (N_3744,N_3321,N_3591);
and U3745 (N_3745,N_3371,N_3559);
xnor U3746 (N_3746,N_3446,N_3423);
or U3747 (N_3747,N_3333,N_3402);
xnor U3748 (N_3748,N_3347,N_3524);
nand U3749 (N_3749,N_3387,N_3442);
or U3750 (N_3750,N_3549,N_3402);
nand U3751 (N_3751,N_3420,N_3428);
xnor U3752 (N_3752,N_3533,N_3361);
xnor U3753 (N_3753,N_3553,N_3367);
xor U3754 (N_3754,N_3369,N_3449);
or U3755 (N_3755,N_3597,N_3402);
or U3756 (N_3756,N_3477,N_3599);
or U3757 (N_3757,N_3320,N_3360);
nand U3758 (N_3758,N_3509,N_3335);
xor U3759 (N_3759,N_3579,N_3443);
nand U3760 (N_3760,N_3579,N_3498);
nor U3761 (N_3761,N_3328,N_3511);
nand U3762 (N_3762,N_3494,N_3549);
and U3763 (N_3763,N_3453,N_3428);
nor U3764 (N_3764,N_3410,N_3586);
or U3765 (N_3765,N_3449,N_3580);
xor U3766 (N_3766,N_3383,N_3454);
nor U3767 (N_3767,N_3478,N_3556);
nand U3768 (N_3768,N_3591,N_3583);
or U3769 (N_3769,N_3520,N_3359);
or U3770 (N_3770,N_3380,N_3493);
xor U3771 (N_3771,N_3354,N_3520);
xor U3772 (N_3772,N_3303,N_3500);
or U3773 (N_3773,N_3564,N_3502);
xor U3774 (N_3774,N_3302,N_3357);
or U3775 (N_3775,N_3331,N_3410);
or U3776 (N_3776,N_3384,N_3321);
nor U3777 (N_3777,N_3512,N_3401);
nand U3778 (N_3778,N_3381,N_3516);
or U3779 (N_3779,N_3367,N_3482);
and U3780 (N_3780,N_3583,N_3346);
nand U3781 (N_3781,N_3492,N_3526);
and U3782 (N_3782,N_3371,N_3359);
or U3783 (N_3783,N_3457,N_3511);
or U3784 (N_3784,N_3467,N_3530);
or U3785 (N_3785,N_3380,N_3465);
nand U3786 (N_3786,N_3522,N_3359);
nand U3787 (N_3787,N_3511,N_3518);
or U3788 (N_3788,N_3388,N_3406);
or U3789 (N_3789,N_3382,N_3478);
or U3790 (N_3790,N_3598,N_3583);
xor U3791 (N_3791,N_3571,N_3578);
nand U3792 (N_3792,N_3536,N_3473);
nand U3793 (N_3793,N_3465,N_3556);
and U3794 (N_3794,N_3492,N_3412);
xnor U3795 (N_3795,N_3473,N_3508);
and U3796 (N_3796,N_3521,N_3417);
xnor U3797 (N_3797,N_3549,N_3537);
xor U3798 (N_3798,N_3545,N_3569);
xor U3799 (N_3799,N_3352,N_3591);
nand U3800 (N_3800,N_3403,N_3487);
and U3801 (N_3801,N_3569,N_3306);
and U3802 (N_3802,N_3474,N_3412);
nor U3803 (N_3803,N_3485,N_3333);
or U3804 (N_3804,N_3330,N_3557);
and U3805 (N_3805,N_3494,N_3398);
xor U3806 (N_3806,N_3305,N_3304);
nor U3807 (N_3807,N_3571,N_3381);
nand U3808 (N_3808,N_3582,N_3587);
and U3809 (N_3809,N_3425,N_3304);
nor U3810 (N_3810,N_3317,N_3449);
nand U3811 (N_3811,N_3482,N_3595);
nor U3812 (N_3812,N_3395,N_3430);
or U3813 (N_3813,N_3378,N_3325);
nor U3814 (N_3814,N_3564,N_3314);
nand U3815 (N_3815,N_3430,N_3566);
and U3816 (N_3816,N_3449,N_3508);
and U3817 (N_3817,N_3574,N_3303);
or U3818 (N_3818,N_3443,N_3548);
xor U3819 (N_3819,N_3380,N_3358);
and U3820 (N_3820,N_3386,N_3568);
xor U3821 (N_3821,N_3366,N_3338);
nand U3822 (N_3822,N_3563,N_3382);
xnor U3823 (N_3823,N_3545,N_3541);
nor U3824 (N_3824,N_3413,N_3551);
or U3825 (N_3825,N_3485,N_3549);
xor U3826 (N_3826,N_3342,N_3413);
or U3827 (N_3827,N_3468,N_3442);
or U3828 (N_3828,N_3400,N_3497);
and U3829 (N_3829,N_3480,N_3477);
or U3830 (N_3830,N_3350,N_3323);
and U3831 (N_3831,N_3413,N_3564);
or U3832 (N_3832,N_3390,N_3544);
or U3833 (N_3833,N_3500,N_3316);
xor U3834 (N_3834,N_3566,N_3308);
xnor U3835 (N_3835,N_3416,N_3522);
xor U3836 (N_3836,N_3486,N_3360);
nor U3837 (N_3837,N_3416,N_3376);
xor U3838 (N_3838,N_3547,N_3338);
xnor U3839 (N_3839,N_3563,N_3509);
xor U3840 (N_3840,N_3336,N_3314);
or U3841 (N_3841,N_3506,N_3304);
nand U3842 (N_3842,N_3508,N_3392);
nand U3843 (N_3843,N_3532,N_3536);
and U3844 (N_3844,N_3503,N_3593);
nor U3845 (N_3845,N_3373,N_3511);
nand U3846 (N_3846,N_3470,N_3430);
and U3847 (N_3847,N_3446,N_3301);
nand U3848 (N_3848,N_3566,N_3541);
or U3849 (N_3849,N_3551,N_3357);
xnor U3850 (N_3850,N_3338,N_3568);
xor U3851 (N_3851,N_3515,N_3498);
xor U3852 (N_3852,N_3446,N_3441);
nand U3853 (N_3853,N_3506,N_3495);
or U3854 (N_3854,N_3315,N_3343);
xor U3855 (N_3855,N_3511,N_3587);
nand U3856 (N_3856,N_3357,N_3500);
nor U3857 (N_3857,N_3510,N_3485);
nand U3858 (N_3858,N_3477,N_3466);
nor U3859 (N_3859,N_3438,N_3352);
nor U3860 (N_3860,N_3562,N_3577);
and U3861 (N_3861,N_3590,N_3578);
xor U3862 (N_3862,N_3316,N_3568);
xnor U3863 (N_3863,N_3412,N_3448);
or U3864 (N_3864,N_3309,N_3529);
xor U3865 (N_3865,N_3490,N_3350);
nand U3866 (N_3866,N_3591,N_3598);
xnor U3867 (N_3867,N_3517,N_3418);
and U3868 (N_3868,N_3530,N_3333);
and U3869 (N_3869,N_3529,N_3580);
nand U3870 (N_3870,N_3553,N_3399);
nor U3871 (N_3871,N_3491,N_3555);
nand U3872 (N_3872,N_3552,N_3433);
xor U3873 (N_3873,N_3401,N_3592);
xor U3874 (N_3874,N_3553,N_3543);
xor U3875 (N_3875,N_3571,N_3471);
nand U3876 (N_3876,N_3350,N_3595);
and U3877 (N_3877,N_3571,N_3505);
xnor U3878 (N_3878,N_3310,N_3457);
or U3879 (N_3879,N_3323,N_3481);
nand U3880 (N_3880,N_3378,N_3540);
nand U3881 (N_3881,N_3460,N_3349);
nand U3882 (N_3882,N_3325,N_3453);
nor U3883 (N_3883,N_3338,N_3546);
nand U3884 (N_3884,N_3407,N_3452);
or U3885 (N_3885,N_3358,N_3419);
xnor U3886 (N_3886,N_3340,N_3352);
or U3887 (N_3887,N_3318,N_3330);
xor U3888 (N_3888,N_3349,N_3309);
nand U3889 (N_3889,N_3395,N_3564);
nand U3890 (N_3890,N_3479,N_3460);
nor U3891 (N_3891,N_3447,N_3589);
nand U3892 (N_3892,N_3326,N_3432);
xnor U3893 (N_3893,N_3511,N_3426);
nand U3894 (N_3894,N_3478,N_3449);
nand U3895 (N_3895,N_3546,N_3304);
nor U3896 (N_3896,N_3398,N_3516);
nor U3897 (N_3897,N_3420,N_3378);
and U3898 (N_3898,N_3354,N_3587);
and U3899 (N_3899,N_3306,N_3329);
or U3900 (N_3900,N_3702,N_3775);
nand U3901 (N_3901,N_3660,N_3694);
nand U3902 (N_3902,N_3614,N_3705);
nor U3903 (N_3903,N_3770,N_3707);
and U3904 (N_3904,N_3679,N_3888);
nand U3905 (N_3905,N_3665,N_3642);
nand U3906 (N_3906,N_3738,N_3723);
xor U3907 (N_3907,N_3778,N_3895);
nor U3908 (N_3908,N_3818,N_3821);
nor U3909 (N_3909,N_3631,N_3794);
or U3910 (N_3910,N_3715,N_3805);
or U3911 (N_3911,N_3675,N_3887);
nor U3912 (N_3912,N_3883,N_3875);
and U3913 (N_3913,N_3712,N_3717);
nor U3914 (N_3914,N_3754,N_3662);
nor U3915 (N_3915,N_3654,N_3615);
and U3916 (N_3916,N_3852,N_3840);
and U3917 (N_3917,N_3739,N_3800);
nor U3918 (N_3918,N_3892,N_3830);
nor U3919 (N_3919,N_3721,N_3655);
or U3920 (N_3920,N_3652,N_3713);
xor U3921 (N_3921,N_3701,N_3896);
or U3922 (N_3922,N_3756,N_3666);
nor U3923 (N_3923,N_3815,N_3628);
xnor U3924 (N_3924,N_3647,N_3613);
and U3925 (N_3925,N_3606,N_3877);
and U3926 (N_3926,N_3743,N_3710);
xor U3927 (N_3927,N_3685,N_3769);
or U3928 (N_3928,N_3856,N_3760);
nor U3929 (N_3929,N_3726,N_3643);
nand U3930 (N_3930,N_3878,N_3700);
and U3931 (N_3931,N_3746,N_3893);
xor U3932 (N_3932,N_3785,N_3841);
xnor U3933 (N_3933,N_3882,N_3616);
and U3934 (N_3934,N_3859,N_3696);
or U3935 (N_3935,N_3668,N_3811);
nor U3936 (N_3936,N_3798,N_3605);
nand U3937 (N_3937,N_3608,N_3607);
xor U3938 (N_3938,N_3764,N_3693);
nand U3939 (N_3939,N_3784,N_3687);
nand U3940 (N_3940,N_3629,N_3774);
xor U3941 (N_3941,N_3771,N_3753);
nor U3942 (N_3942,N_3803,N_3781);
nand U3943 (N_3943,N_3640,N_3682);
and U3944 (N_3944,N_3879,N_3653);
xor U3945 (N_3945,N_3870,N_3611);
nand U3946 (N_3946,N_3724,N_3644);
or U3947 (N_3947,N_3829,N_3850);
nand U3948 (N_3948,N_3703,N_3826);
nand U3949 (N_3949,N_3734,N_3704);
nor U3950 (N_3950,N_3833,N_3767);
xnor U3951 (N_3951,N_3796,N_3890);
xor U3952 (N_3952,N_3719,N_3737);
nor U3953 (N_3953,N_3789,N_3792);
and U3954 (N_3954,N_3793,N_3897);
nor U3955 (N_3955,N_3637,N_3661);
and U3956 (N_3956,N_3773,N_3788);
nand U3957 (N_3957,N_3757,N_3880);
xor U3958 (N_3958,N_3858,N_3853);
nand U3959 (N_3959,N_3664,N_3672);
or U3960 (N_3960,N_3849,N_3641);
nor U3961 (N_3961,N_3835,N_3657);
nor U3962 (N_3962,N_3632,N_3745);
xor U3963 (N_3963,N_3824,N_3855);
or U3964 (N_3964,N_3797,N_3677);
or U3965 (N_3965,N_3646,N_3808);
and U3966 (N_3966,N_3630,N_3639);
and U3967 (N_3967,N_3722,N_3862);
and U3968 (N_3968,N_3752,N_3891);
xnor U3969 (N_3969,N_3742,N_3609);
xor U3970 (N_3970,N_3716,N_3843);
or U3971 (N_3971,N_3741,N_3868);
nand U3972 (N_3972,N_3699,N_3678);
nand U3973 (N_3973,N_3758,N_3804);
nand U3974 (N_3974,N_3844,N_3720);
nor U3975 (N_3975,N_3780,N_3633);
and U3976 (N_3976,N_3698,N_3747);
or U3977 (N_3977,N_3648,N_3857);
and U3978 (N_3978,N_3671,N_3799);
and U3979 (N_3979,N_3620,N_3684);
or U3980 (N_3980,N_3600,N_3669);
or U3981 (N_3981,N_3626,N_3842);
nand U3982 (N_3982,N_3776,N_3873);
xnor U3983 (N_3983,N_3761,N_3866);
nand U3984 (N_3984,N_3711,N_3865);
and U3985 (N_3985,N_3663,N_3861);
xnor U3986 (N_3986,N_3819,N_3674);
nor U3987 (N_3987,N_3827,N_3656);
nor U3988 (N_3988,N_3689,N_3832);
nand U3989 (N_3989,N_3708,N_3714);
xor U3990 (N_3990,N_3786,N_3766);
nand U3991 (N_3991,N_3728,N_3874);
nand U3992 (N_3992,N_3807,N_3740);
and U3993 (N_3993,N_3680,N_3831);
xor U3994 (N_3994,N_3650,N_3839);
nand U3995 (N_3995,N_3725,N_3816);
xor U3996 (N_3996,N_3881,N_3871);
or U3997 (N_3997,N_3790,N_3820);
and U3998 (N_3998,N_3709,N_3886);
xor U3999 (N_3999,N_3765,N_3894);
nor U4000 (N_4000,N_3884,N_3795);
and U4001 (N_4001,N_3809,N_3762);
and U4002 (N_4002,N_3869,N_3823);
or U4003 (N_4003,N_3867,N_3670);
and U4004 (N_4004,N_3759,N_3812);
xor U4005 (N_4005,N_3601,N_3864);
and U4006 (N_4006,N_3755,N_3847);
nor U4007 (N_4007,N_3692,N_3688);
nand U4008 (N_4008,N_3610,N_3602);
nor U4009 (N_4009,N_3732,N_3889);
xor U4010 (N_4010,N_3872,N_3791);
nand U4011 (N_4011,N_3623,N_3635);
or U4012 (N_4012,N_3636,N_3730);
xor U4013 (N_4013,N_3681,N_3619);
or U4014 (N_4014,N_3733,N_3736);
nor U4015 (N_4015,N_3727,N_3801);
nand U4016 (N_4016,N_3634,N_3731);
or U4017 (N_4017,N_3898,N_3763);
and U4018 (N_4018,N_3612,N_3863);
and U4019 (N_4019,N_3848,N_3718);
nand U4020 (N_4020,N_3683,N_3779);
xnor U4021 (N_4021,N_3625,N_3846);
nand U4022 (N_4022,N_3802,N_3787);
nor U4023 (N_4023,N_3854,N_3690);
or U4024 (N_4024,N_3749,N_3667);
nand U4025 (N_4025,N_3706,N_3603);
xor U4026 (N_4026,N_3772,N_3618);
or U4027 (N_4027,N_3822,N_3837);
nand U4028 (N_4028,N_3676,N_3828);
nor U4029 (N_4029,N_3695,N_3624);
nand U4030 (N_4030,N_3813,N_3651);
xnor U4031 (N_4031,N_3851,N_3817);
and U4032 (N_4032,N_3777,N_3649);
xnor U4033 (N_4033,N_3691,N_3810);
nor U4034 (N_4034,N_3825,N_3729);
or U4035 (N_4035,N_3885,N_3751);
and U4036 (N_4036,N_3658,N_3735);
and U4037 (N_4037,N_3876,N_3783);
nor U4038 (N_4038,N_3617,N_3899);
nand U4039 (N_4039,N_3806,N_3686);
xnor U4040 (N_4040,N_3627,N_3621);
nand U4041 (N_4041,N_3845,N_3697);
nand U4042 (N_4042,N_3834,N_3638);
and U4043 (N_4043,N_3838,N_3782);
nand U4044 (N_4044,N_3673,N_3750);
and U4045 (N_4045,N_3860,N_3604);
nand U4046 (N_4046,N_3814,N_3748);
nand U4047 (N_4047,N_3659,N_3645);
and U4048 (N_4048,N_3836,N_3744);
nor U4049 (N_4049,N_3768,N_3622);
and U4050 (N_4050,N_3626,N_3735);
nor U4051 (N_4051,N_3796,N_3846);
nand U4052 (N_4052,N_3871,N_3887);
nand U4053 (N_4053,N_3611,N_3660);
nand U4054 (N_4054,N_3667,N_3770);
and U4055 (N_4055,N_3639,N_3789);
and U4056 (N_4056,N_3698,N_3686);
nor U4057 (N_4057,N_3857,N_3618);
and U4058 (N_4058,N_3832,N_3756);
xnor U4059 (N_4059,N_3892,N_3653);
xor U4060 (N_4060,N_3788,N_3754);
xnor U4061 (N_4061,N_3748,N_3783);
nor U4062 (N_4062,N_3858,N_3755);
nand U4063 (N_4063,N_3845,N_3646);
xor U4064 (N_4064,N_3781,N_3811);
nor U4065 (N_4065,N_3818,N_3615);
nand U4066 (N_4066,N_3644,N_3884);
or U4067 (N_4067,N_3880,N_3652);
nand U4068 (N_4068,N_3821,N_3800);
and U4069 (N_4069,N_3608,N_3808);
and U4070 (N_4070,N_3871,N_3742);
nor U4071 (N_4071,N_3696,N_3725);
nor U4072 (N_4072,N_3613,N_3625);
xnor U4073 (N_4073,N_3754,N_3720);
and U4074 (N_4074,N_3720,N_3807);
or U4075 (N_4075,N_3896,N_3772);
nand U4076 (N_4076,N_3812,N_3707);
and U4077 (N_4077,N_3655,N_3734);
and U4078 (N_4078,N_3708,N_3759);
or U4079 (N_4079,N_3730,N_3658);
and U4080 (N_4080,N_3827,N_3849);
nand U4081 (N_4081,N_3803,N_3744);
xor U4082 (N_4082,N_3886,N_3847);
or U4083 (N_4083,N_3645,N_3867);
nor U4084 (N_4084,N_3815,N_3666);
or U4085 (N_4085,N_3693,N_3600);
xor U4086 (N_4086,N_3747,N_3647);
or U4087 (N_4087,N_3676,N_3727);
and U4088 (N_4088,N_3724,N_3680);
nor U4089 (N_4089,N_3838,N_3815);
and U4090 (N_4090,N_3884,N_3745);
nor U4091 (N_4091,N_3662,N_3680);
nand U4092 (N_4092,N_3899,N_3878);
xor U4093 (N_4093,N_3722,N_3718);
nand U4094 (N_4094,N_3724,N_3818);
nor U4095 (N_4095,N_3757,N_3625);
and U4096 (N_4096,N_3731,N_3696);
or U4097 (N_4097,N_3748,N_3674);
xnor U4098 (N_4098,N_3688,N_3648);
or U4099 (N_4099,N_3634,N_3657);
xnor U4100 (N_4100,N_3748,N_3650);
nand U4101 (N_4101,N_3860,N_3827);
nand U4102 (N_4102,N_3856,N_3733);
and U4103 (N_4103,N_3624,N_3711);
or U4104 (N_4104,N_3632,N_3711);
nor U4105 (N_4105,N_3610,N_3772);
xnor U4106 (N_4106,N_3631,N_3613);
xnor U4107 (N_4107,N_3745,N_3654);
and U4108 (N_4108,N_3633,N_3685);
nor U4109 (N_4109,N_3681,N_3816);
and U4110 (N_4110,N_3766,N_3742);
nor U4111 (N_4111,N_3855,N_3602);
nor U4112 (N_4112,N_3607,N_3895);
or U4113 (N_4113,N_3601,N_3879);
and U4114 (N_4114,N_3844,N_3703);
nor U4115 (N_4115,N_3608,N_3774);
and U4116 (N_4116,N_3720,N_3895);
and U4117 (N_4117,N_3892,N_3883);
xnor U4118 (N_4118,N_3861,N_3640);
nor U4119 (N_4119,N_3743,N_3798);
nor U4120 (N_4120,N_3816,N_3741);
nor U4121 (N_4121,N_3732,N_3838);
xor U4122 (N_4122,N_3725,N_3677);
nor U4123 (N_4123,N_3650,N_3838);
nor U4124 (N_4124,N_3693,N_3671);
xnor U4125 (N_4125,N_3625,N_3754);
and U4126 (N_4126,N_3770,N_3825);
xnor U4127 (N_4127,N_3871,N_3608);
nand U4128 (N_4128,N_3691,N_3876);
nand U4129 (N_4129,N_3632,N_3749);
nand U4130 (N_4130,N_3800,N_3883);
or U4131 (N_4131,N_3743,N_3773);
xnor U4132 (N_4132,N_3872,N_3884);
and U4133 (N_4133,N_3600,N_3831);
nor U4134 (N_4134,N_3731,N_3752);
nand U4135 (N_4135,N_3785,N_3683);
xor U4136 (N_4136,N_3822,N_3744);
or U4137 (N_4137,N_3663,N_3753);
xor U4138 (N_4138,N_3660,N_3720);
or U4139 (N_4139,N_3606,N_3867);
nand U4140 (N_4140,N_3603,N_3746);
and U4141 (N_4141,N_3733,N_3775);
nor U4142 (N_4142,N_3731,N_3662);
xor U4143 (N_4143,N_3775,N_3744);
nand U4144 (N_4144,N_3693,N_3822);
or U4145 (N_4145,N_3745,N_3788);
nand U4146 (N_4146,N_3838,N_3787);
or U4147 (N_4147,N_3715,N_3623);
and U4148 (N_4148,N_3658,N_3740);
or U4149 (N_4149,N_3637,N_3627);
or U4150 (N_4150,N_3681,N_3677);
and U4151 (N_4151,N_3688,N_3853);
xor U4152 (N_4152,N_3893,N_3729);
nor U4153 (N_4153,N_3893,N_3694);
nand U4154 (N_4154,N_3630,N_3827);
xnor U4155 (N_4155,N_3704,N_3605);
or U4156 (N_4156,N_3676,N_3848);
nand U4157 (N_4157,N_3635,N_3828);
nand U4158 (N_4158,N_3855,N_3631);
xnor U4159 (N_4159,N_3849,N_3850);
or U4160 (N_4160,N_3744,N_3638);
and U4161 (N_4161,N_3871,N_3664);
and U4162 (N_4162,N_3724,N_3676);
and U4163 (N_4163,N_3866,N_3864);
nor U4164 (N_4164,N_3899,N_3667);
nor U4165 (N_4165,N_3894,N_3617);
nand U4166 (N_4166,N_3655,N_3644);
and U4167 (N_4167,N_3709,N_3762);
nand U4168 (N_4168,N_3668,N_3761);
xor U4169 (N_4169,N_3654,N_3641);
xor U4170 (N_4170,N_3869,N_3822);
nor U4171 (N_4171,N_3884,N_3761);
and U4172 (N_4172,N_3818,N_3880);
and U4173 (N_4173,N_3695,N_3860);
and U4174 (N_4174,N_3734,N_3622);
nor U4175 (N_4175,N_3641,N_3841);
or U4176 (N_4176,N_3687,N_3755);
xor U4177 (N_4177,N_3776,N_3720);
or U4178 (N_4178,N_3650,N_3745);
or U4179 (N_4179,N_3849,N_3874);
nand U4180 (N_4180,N_3794,N_3815);
and U4181 (N_4181,N_3622,N_3824);
or U4182 (N_4182,N_3739,N_3625);
nor U4183 (N_4183,N_3657,N_3856);
or U4184 (N_4184,N_3750,N_3699);
or U4185 (N_4185,N_3636,N_3787);
nor U4186 (N_4186,N_3745,N_3874);
or U4187 (N_4187,N_3873,N_3656);
nor U4188 (N_4188,N_3823,N_3677);
nand U4189 (N_4189,N_3687,N_3872);
nor U4190 (N_4190,N_3755,N_3663);
or U4191 (N_4191,N_3835,N_3776);
xnor U4192 (N_4192,N_3866,N_3882);
nor U4193 (N_4193,N_3629,N_3743);
nand U4194 (N_4194,N_3615,N_3862);
and U4195 (N_4195,N_3674,N_3855);
and U4196 (N_4196,N_3687,N_3899);
xor U4197 (N_4197,N_3661,N_3695);
or U4198 (N_4198,N_3678,N_3603);
xor U4199 (N_4199,N_3804,N_3859);
nor U4200 (N_4200,N_4047,N_4163);
xor U4201 (N_4201,N_3930,N_4030);
nand U4202 (N_4202,N_4197,N_4049);
xnor U4203 (N_4203,N_4169,N_4166);
and U4204 (N_4204,N_4160,N_4167);
nor U4205 (N_4205,N_3991,N_4148);
xor U4206 (N_4206,N_4068,N_3972);
nor U4207 (N_4207,N_4004,N_3966);
xor U4208 (N_4208,N_3922,N_3912);
or U4209 (N_4209,N_3974,N_4103);
and U4210 (N_4210,N_4183,N_4143);
and U4211 (N_4211,N_4076,N_4170);
nor U4212 (N_4212,N_4077,N_3903);
nor U4213 (N_4213,N_3959,N_4108);
nor U4214 (N_4214,N_4084,N_4127);
nand U4215 (N_4215,N_4181,N_3946);
or U4216 (N_4216,N_4125,N_4037);
and U4217 (N_4217,N_4048,N_3996);
and U4218 (N_4218,N_4137,N_4132);
nand U4219 (N_4219,N_3990,N_4119);
nor U4220 (N_4220,N_3962,N_4193);
or U4221 (N_4221,N_3908,N_4098);
or U4222 (N_4222,N_3954,N_4097);
xnor U4223 (N_4223,N_3984,N_3905);
and U4224 (N_4224,N_4029,N_4154);
and U4225 (N_4225,N_3950,N_3965);
and U4226 (N_4226,N_4131,N_4052);
nor U4227 (N_4227,N_4012,N_4088);
or U4228 (N_4228,N_3995,N_4139);
xnor U4229 (N_4229,N_3967,N_4152);
nand U4230 (N_4230,N_4023,N_3944);
xor U4231 (N_4231,N_4051,N_3952);
nand U4232 (N_4232,N_4199,N_3999);
xor U4233 (N_4233,N_3979,N_4019);
xnor U4234 (N_4234,N_3915,N_3963);
nor U4235 (N_4235,N_4039,N_3958);
xnor U4236 (N_4236,N_4159,N_4142);
nor U4237 (N_4237,N_3916,N_4109);
nand U4238 (N_4238,N_3917,N_3970);
xor U4239 (N_4239,N_4136,N_4003);
and U4240 (N_4240,N_3977,N_4190);
and U4241 (N_4241,N_4106,N_3909);
and U4242 (N_4242,N_4145,N_3913);
xor U4243 (N_4243,N_3918,N_4079);
and U4244 (N_4244,N_4028,N_4038);
xnor U4245 (N_4245,N_4020,N_4149);
and U4246 (N_4246,N_4112,N_3982);
or U4247 (N_4247,N_4063,N_4042);
nand U4248 (N_4248,N_3947,N_4044);
nor U4249 (N_4249,N_4101,N_4050);
xor U4250 (N_4250,N_3931,N_4086);
and U4251 (N_4251,N_3961,N_3920);
nor U4252 (N_4252,N_4058,N_4006);
nor U4253 (N_4253,N_4123,N_4041);
and U4254 (N_4254,N_4031,N_3914);
or U4255 (N_4255,N_4156,N_4065);
xnor U4256 (N_4256,N_4091,N_4026);
and U4257 (N_4257,N_4054,N_3902);
nor U4258 (N_4258,N_4069,N_4055);
xor U4259 (N_4259,N_4124,N_4128);
nor U4260 (N_4260,N_4032,N_3956);
or U4261 (N_4261,N_4110,N_4196);
xor U4262 (N_4262,N_4191,N_4107);
nand U4263 (N_4263,N_3937,N_3976);
and U4264 (N_4264,N_4158,N_3978);
and U4265 (N_4265,N_4195,N_4083);
xor U4266 (N_4266,N_4095,N_4016);
nor U4267 (N_4267,N_4045,N_4102);
and U4268 (N_4268,N_3925,N_4105);
or U4269 (N_4269,N_4024,N_4185);
and U4270 (N_4270,N_3904,N_4113);
nand U4271 (N_4271,N_4025,N_4085);
nor U4272 (N_4272,N_4171,N_4104);
and U4273 (N_4273,N_4005,N_3964);
or U4274 (N_4274,N_4057,N_4182);
xnor U4275 (N_4275,N_4146,N_4178);
nand U4276 (N_4276,N_4192,N_3940);
nand U4277 (N_4277,N_3981,N_3945);
or U4278 (N_4278,N_4172,N_4053);
nand U4279 (N_4279,N_3971,N_4072);
xnor U4280 (N_4280,N_4071,N_3910);
xor U4281 (N_4281,N_4002,N_4153);
and U4282 (N_4282,N_4114,N_4180);
and U4283 (N_4283,N_4062,N_3968);
and U4284 (N_4284,N_3985,N_3942);
nor U4285 (N_4285,N_4008,N_3935);
nor U4286 (N_4286,N_4080,N_4033);
xor U4287 (N_4287,N_3919,N_4061);
nand U4288 (N_4288,N_4094,N_4151);
nand U4289 (N_4289,N_4116,N_3938);
xnor U4290 (N_4290,N_3994,N_4040);
or U4291 (N_4291,N_3900,N_3997);
and U4292 (N_4292,N_4147,N_4162);
nand U4293 (N_4293,N_3923,N_4036);
xor U4294 (N_4294,N_4070,N_4100);
nor U4295 (N_4295,N_4168,N_3928);
or U4296 (N_4296,N_3927,N_4133);
nor U4297 (N_4297,N_4081,N_4122);
nor U4298 (N_4298,N_4015,N_4189);
or U4299 (N_4299,N_3973,N_3953);
or U4300 (N_4300,N_3987,N_3948);
nor U4301 (N_4301,N_3941,N_4027);
or U4302 (N_4302,N_3988,N_4001);
nor U4303 (N_4303,N_4165,N_4175);
xnor U4304 (N_4304,N_4198,N_4078);
nand U4305 (N_4305,N_3926,N_4067);
nor U4306 (N_4306,N_4187,N_4134);
nand U4307 (N_4307,N_4075,N_4186);
and U4308 (N_4308,N_4140,N_4173);
nor U4309 (N_4309,N_4060,N_3934);
nor U4310 (N_4310,N_4194,N_4184);
or U4311 (N_4311,N_4056,N_4164);
nand U4312 (N_4312,N_4174,N_4021);
nand U4313 (N_4313,N_3936,N_4007);
xnor U4314 (N_4314,N_4043,N_3955);
nand U4315 (N_4315,N_4161,N_4014);
or U4316 (N_4316,N_4017,N_3993);
and U4317 (N_4317,N_4059,N_3989);
xor U4318 (N_4318,N_3929,N_4188);
and U4319 (N_4319,N_4141,N_4176);
and U4320 (N_4320,N_4000,N_3921);
nand U4321 (N_4321,N_4126,N_4018);
nand U4322 (N_4322,N_3998,N_3980);
and U4323 (N_4323,N_4129,N_3983);
nor U4324 (N_4324,N_4111,N_4120);
nor U4325 (N_4325,N_4022,N_4066);
xnor U4326 (N_4326,N_4144,N_3951);
and U4327 (N_4327,N_3975,N_4118);
and U4328 (N_4328,N_4009,N_3933);
or U4329 (N_4329,N_4099,N_4074);
nand U4330 (N_4330,N_4013,N_4082);
nand U4331 (N_4331,N_3911,N_3969);
nor U4332 (N_4332,N_4093,N_3992);
nand U4333 (N_4333,N_3906,N_4115);
and U4334 (N_4334,N_4096,N_3924);
or U4335 (N_4335,N_4121,N_4035);
and U4336 (N_4336,N_4157,N_3943);
nand U4337 (N_4337,N_4087,N_4135);
nor U4338 (N_4338,N_4034,N_4117);
and U4339 (N_4339,N_3957,N_4010);
and U4340 (N_4340,N_4155,N_4011);
xnor U4341 (N_4341,N_3949,N_4092);
or U4342 (N_4342,N_3939,N_4090);
nor U4343 (N_4343,N_4179,N_3901);
or U4344 (N_4344,N_4130,N_3932);
or U4345 (N_4345,N_4150,N_3960);
nor U4346 (N_4346,N_4177,N_4138);
nor U4347 (N_4347,N_4046,N_3907);
and U4348 (N_4348,N_4089,N_4073);
xor U4349 (N_4349,N_4064,N_3986);
xnor U4350 (N_4350,N_3994,N_4014);
and U4351 (N_4351,N_4075,N_4050);
nand U4352 (N_4352,N_4044,N_4016);
xor U4353 (N_4353,N_4096,N_4036);
or U4354 (N_4354,N_4141,N_3957);
xnor U4355 (N_4355,N_3921,N_4128);
or U4356 (N_4356,N_4116,N_4085);
or U4357 (N_4357,N_4053,N_3953);
and U4358 (N_4358,N_4130,N_4022);
nand U4359 (N_4359,N_4086,N_4115);
nor U4360 (N_4360,N_4073,N_3956);
xnor U4361 (N_4361,N_4125,N_4102);
and U4362 (N_4362,N_3992,N_4199);
nor U4363 (N_4363,N_3968,N_4101);
nand U4364 (N_4364,N_3907,N_3922);
and U4365 (N_4365,N_4003,N_4191);
xor U4366 (N_4366,N_4146,N_4048);
nor U4367 (N_4367,N_4035,N_4011);
xnor U4368 (N_4368,N_4037,N_3985);
xor U4369 (N_4369,N_4125,N_3906);
and U4370 (N_4370,N_4013,N_4048);
xor U4371 (N_4371,N_4087,N_3900);
nand U4372 (N_4372,N_4166,N_4076);
and U4373 (N_4373,N_4109,N_3959);
nand U4374 (N_4374,N_3961,N_4070);
and U4375 (N_4375,N_3994,N_3944);
or U4376 (N_4376,N_3984,N_3957);
nand U4377 (N_4377,N_3985,N_4152);
and U4378 (N_4378,N_3933,N_4195);
or U4379 (N_4379,N_4184,N_4038);
nor U4380 (N_4380,N_4045,N_3911);
xor U4381 (N_4381,N_4175,N_4058);
or U4382 (N_4382,N_4058,N_3948);
xor U4383 (N_4383,N_4118,N_4032);
nand U4384 (N_4384,N_4089,N_4060);
nor U4385 (N_4385,N_4079,N_4049);
or U4386 (N_4386,N_4191,N_4079);
xnor U4387 (N_4387,N_4109,N_4079);
and U4388 (N_4388,N_4052,N_4015);
or U4389 (N_4389,N_4060,N_4007);
or U4390 (N_4390,N_4111,N_4015);
nor U4391 (N_4391,N_4062,N_4042);
nor U4392 (N_4392,N_3995,N_4078);
and U4393 (N_4393,N_4118,N_4145);
nor U4394 (N_4394,N_3974,N_3954);
xnor U4395 (N_4395,N_4044,N_3945);
xor U4396 (N_4396,N_4122,N_4044);
or U4397 (N_4397,N_4098,N_3929);
or U4398 (N_4398,N_3922,N_4005);
xnor U4399 (N_4399,N_3937,N_4007);
and U4400 (N_4400,N_3930,N_3988);
or U4401 (N_4401,N_3981,N_4114);
or U4402 (N_4402,N_4154,N_4071);
nor U4403 (N_4403,N_3973,N_4114);
nand U4404 (N_4404,N_4146,N_4065);
and U4405 (N_4405,N_4178,N_4118);
nor U4406 (N_4406,N_4101,N_4012);
xor U4407 (N_4407,N_4037,N_3920);
nand U4408 (N_4408,N_3918,N_4180);
and U4409 (N_4409,N_3942,N_4020);
or U4410 (N_4410,N_4130,N_3994);
and U4411 (N_4411,N_3914,N_3994);
nand U4412 (N_4412,N_4058,N_4034);
or U4413 (N_4413,N_4047,N_4068);
nor U4414 (N_4414,N_3923,N_4181);
or U4415 (N_4415,N_4018,N_4189);
or U4416 (N_4416,N_4008,N_4119);
nand U4417 (N_4417,N_4005,N_4137);
and U4418 (N_4418,N_4111,N_3921);
or U4419 (N_4419,N_3948,N_4195);
nor U4420 (N_4420,N_3950,N_4069);
nor U4421 (N_4421,N_3916,N_4030);
and U4422 (N_4422,N_3901,N_4193);
or U4423 (N_4423,N_4063,N_3987);
and U4424 (N_4424,N_4073,N_3978);
or U4425 (N_4425,N_3948,N_4125);
and U4426 (N_4426,N_4084,N_4075);
or U4427 (N_4427,N_4043,N_4078);
nor U4428 (N_4428,N_4105,N_4170);
or U4429 (N_4429,N_4164,N_4119);
or U4430 (N_4430,N_4107,N_3976);
nand U4431 (N_4431,N_3935,N_4111);
nand U4432 (N_4432,N_4125,N_4026);
and U4433 (N_4433,N_4116,N_3932);
or U4434 (N_4434,N_4075,N_4029);
xnor U4435 (N_4435,N_4066,N_4165);
nand U4436 (N_4436,N_4091,N_4194);
or U4437 (N_4437,N_4105,N_3953);
or U4438 (N_4438,N_3995,N_3972);
nand U4439 (N_4439,N_4164,N_4136);
xor U4440 (N_4440,N_4118,N_4159);
or U4441 (N_4441,N_3973,N_4110);
nand U4442 (N_4442,N_3903,N_4168);
or U4443 (N_4443,N_3976,N_4052);
nor U4444 (N_4444,N_4103,N_4077);
or U4445 (N_4445,N_3940,N_4059);
nand U4446 (N_4446,N_4044,N_3922);
nor U4447 (N_4447,N_4183,N_4118);
and U4448 (N_4448,N_4199,N_4034);
nor U4449 (N_4449,N_3939,N_3948);
nand U4450 (N_4450,N_3915,N_3990);
xor U4451 (N_4451,N_4137,N_4141);
nor U4452 (N_4452,N_4091,N_3900);
and U4453 (N_4453,N_4017,N_4178);
nor U4454 (N_4454,N_4004,N_4145);
nor U4455 (N_4455,N_4149,N_4173);
nor U4456 (N_4456,N_3955,N_3925);
or U4457 (N_4457,N_4044,N_4132);
and U4458 (N_4458,N_4113,N_4003);
xor U4459 (N_4459,N_4093,N_4132);
xnor U4460 (N_4460,N_4074,N_4141);
nand U4461 (N_4461,N_3946,N_4149);
and U4462 (N_4462,N_4156,N_3940);
or U4463 (N_4463,N_4146,N_4180);
and U4464 (N_4464,N_3989,N_3945);
nor U4465 (N_4465,N_3924,N_4172);
nor U4466 (N_4466,N_3997,N_3980);
nand U4467 (N_4467,N_3974,N_4157);
nand U4468 (N_4468,N_3986,N_4035);
and U4469 (N_4469,N_4143,N_4042);
or U4470 (N_4470,N_4180,N_4064);
nand U4471 (N_4471,N_4071,N_4161);
and U4472 (N_4472,N_4126,N_3924);
and U4473 (N_4473,N_3915,N_4089);
or U4474 (N_4474,N_4013,N_3937);
and U4475 (N_4475,N_4073,N_3996);
nor U4476 (N_4476,N_3988,N_4041);
xnor U4477 (N_4477,N_3962,N_3986);
and U4478 (N_4478,N_4154,N_3915);
nor U4479 (N_4479,N_4149,N_3954);
nand U4480 (N_4480,N_4067,N_4113);
or U4481 (N_4481,N_3948,N_4145);
nand U4482 (N_4482,N_4112,N_4099);
and U4483 (N_4483,N_4011,N_3922);
nand U4484 (N_4484,N_4124,N_4130);
and U4485 (N_4485,N_4032,N_4085);
or U4486 (N_4486,N_3912,N_4070);
or U4487 (N_4487,N_3958,N_4076);
or U4488 (N_4488,N_3958,N_3955);
and U4489 (N_4489,N_4137,N_4098);
and U4490 (N_4490,N_3986,N_4105);
xnor U4491 (N_4491,N_4049,N_4030);
xnor U4492 (N_4492,N_4140,N_4105);
xor U4493 (N_4493,N_4150,N_3974);
or U4494 (N_4494,N_4054,N_4132);
and U4495 (N_4495,N_4029,N_4115);
nor U4496 (N_4496,N_4017,N_3933);
nand U4497 (N_4497,N_4122,N_4040);
and U4498 (N_4498,N_3955,N_3983);
nand U4499 (N_4499,N_4167,N_3939);
nand U4500 (N_4500,N_4488,N_4252);
or U4501 (N_4501,N_4348,N_4400);
or U4502 (N_4502,N_4267,N_4249);
and U4503 (N_4503,N_4402,N_4268);
or U4504 (N_4504,N_4395,N_4464);
xnor U4505 (N_4505,N_4292,N_4226);
nand U4506 (N_4506,N_4460,N_4280);
and U4507 (N_4507,N_4328,N_4288);
nor U4508 (N_4508,N_4212,N_4450);
or U4509 (N_4509,N_4347,N_4355);
xor U4510 (N_4510,N_4318,N_4274);
and U4511 (N_4511,N_4410,N_4223);
nor U4512 (N_4512,N_4350,N_4428);
nor U4513 (N_4513,N_4234,N_4326);
xor U4514 (N_4514,N_4325,N_4433);
and U4515 (N_4515,N_4342,N_4467);
nand U4516 (N_4516,N_4277,N_4356);
and U4517 (N_4517,N_4431,N_4437);
and U4518 (N_4518,N_4389,N_4374);
nor U4519 (N_4519,N_4452,N_4391);
or U4520 (N_4520,N_4465,N_4334);
xor U4521 (N_4521,N_4373,N_4451);
and U4522 (N_4522,N_4415,N_4362);
and U4523 (N_4523,N_4243,N_4446);
or U4524 (N_4524,N_4321,N_4336);
xor U4525 (N_4525,N_4304,N_4473);
or U4526 (N_4526,N_4396,N_4412);
nor U4527 (N_4527,N_4447,N_4386);
and U4528 (N_4528,N_4315,N_4414);
or U4529 (N_4529,N_4419,N_4247);
and U4530 (N_4530,N_4361,N_4345);
xnor U4531 (N_4531,N_4285,N_4340);
xor U4532 (N_4532,N_4331,N_4341);
or U4533 (N_4533,N_4385,N_4310);
xor U4534 (N_4534,N_4372,N_4490);
or U4535 (N_4535,N_4338,N_4475);
nor U4536 (N_4536,N_4478,N_4206);
and U4537 (N_4537,N_4456,N_4227);
nand U4538 (N_4538,N_4327,N_4276);
nor U4539 (N_4539,N_4454,N_4269);
xor U4540 (N_4540,N_4388,N_4298);
or U4541 (N_4541,N_4262,N_4346);
or U4542 (N_4542,N_4289,N_4216);
nor U4543 (N_4543,N_4427,N_4471);
or U4544 (N_4544,N_4332,N_4273);
nand U4545 (N_4545,N_4339,N_4364);
nor U4546 (N_4546,N_4429,N_4330);
xnor U4547 (N_4547,N_4312,N_4403);
nand U4548 (N_4548,N_4219,N_4455);
nor U4549 (N_4549,N_4317,N_4263);
xnor U4550 (N_4550,N_4354,N_4401);
nor U4551 (N_4551,N_4204,N_4259);
nor U4552 (N_4552,N_4472,N_4393);
xor U4553 (N_4553,N_4469,N_4418);
or U4554 (N_4554,N_4254,N_4359);
and U4555 (N_4555,N_4294,N_4441);
or U4556 (N_4556,N_4493,N_4217);
or U4557 (N_4557,N_4489,N_4248);
or U4558 (N_4558,N_4498,N_4443);
and U4559 (N_4559,N_4413,N_4224);
and U4560 (N_4560,N_4290,N_4442);
or U4561 (N_4561,N_4398,N_4215);
or U4562 (N_4562,N_4238,N_4213);
and U4563 (N_4563,N_4314,N_4235);
or U4564 (N_4564,N_4240,N_4320);
and U4565 (N_4565,N_4377,N_4371);
or U4566 (N_4566,N_4491,N_4316);
and U4567 (N_4567,N_4264,N_4409);
or U4568 (N_4568,N_4408,N_4335);
xor U4569 (N_4569,N_4201,N_4494);
or U4570 (N_4570,N_4476,N_4375);
and U4571 (N_4571,N_4369,N_4463);
nand U4572 (N_4572,N_4236,N_4322);
nor U4573 (N_4573,N_4458,N_4305);
nor U4574 (N_4574,N_4420,N_4207);
or U4575 (N_4575,N_4363,N_4422);
nor U4576 (N_4576,N_4244,N_4230);
nor U4577 (N_4577,N_4497,N_4272);
xor U4578 (N_4578,N_4482,N_4457);
nor U4579 (N_4579,N_4205,N_4250);
nand U4580 (N_4580,N_4229,N_4261);
nor U4581 (N_4581,N_4436,N_4383);
nor U4582 (N_4582,N_4480,N_4448);
or U4583 (N_4583,N_4421,N_4483);
or U4584 (N_4584,N_4440,N_4211);
nor U4585 (N_4585,N_4461,N_4425);
and U4586 (N_4586,N_4357,N_4344);
nand U4587 (N_4587,N_4468,N_4487);
and U4588 (N_4588,N_4218,N_4381);
nand U4589 (N_4589,N_4343,N_4202);
xor U4590 (N_4590,N_4390,N_4225);
and U4591 (N_4591,N_4439,N_4253);
nand U4592 (N_4592,N_4423,N_4291);
xnor U4593 (N_4593,N_4438,N_4387);
nand U4594 (N_4594,N_4210,N_4445);
and U4595 (N_4595,N_4470,N_4246);
or U4596 (N_4596,N_4379,N_4220);
xnor U4597 (N_4597,N_4417,N_4311);
xnor U4598 (N_4598,N_4271,N_4462);
xor U4599 (N_4599,N_4430,N_4426);
nand U4600 (N_4600,N_4496,N_4399);
nor U4601 (N_4601,N_4208,N_4239);
nor U4602 (N_4602,N_4392,N_4286);
nor U4603 (N_4603,N_4382,N_4351);
xnor U4604 (N_4604,N_4221,N_4495);
and U4605 (N_4605,N_4499,N_4406);
or U4606 (N_4606,N_4245,N_4319);
nand U4607 (N_4607,N_4293,N_4485);
and U4608 (N_4608,N_4278,N_4233);
nand U4609 (N_4609,N_4241,N_4466);
and U4610 (N_4610,N_4486,N_4411);
and U4611 (N_4611,N_4303,N_4257);
nand U4612 (N_4612,N_4203,N_4358);
and U4613 (N_4613,N_4353,N_4484);
xnor U4614 (N_4614,N_4231,N_4232);
or U4615 (N_4615,N_4477,N_4296);
or U4616 (N_4616,N_4366,N_4394);
nand U4617 (N_4617,N_4444,N_4333);
nand U4618 (N_4618,N_4275,N_4367);
or U4619 (N_4619,N_4214,N_4324);
nor U4620 (N_4620,N_4306,N_4474);
and U4621 (N_4621,N_4256,N_4307);
and U4622 (N_4622,N_4242,N_4313);
nor U4623 (N_4623,N_4279,N_4365);
or U4624 (N_4624,N_4397,N_4360);
or U4625 (N_4625,N_4260,N_4295);
xor U4626 (N_4626,N_4297,N_4323);
nor U4627 (N_4627,N_4282,N_4380);
and U4628 (N_4628,N_4237,N_4434);
and U4629 (N_4629,N_4251,N_4481);
nand U4630 (N_4630,N_4405,N_4301);
xor U4631 (N_4631,N_4281,N_4300);
and U4632 (N_4632,N_4432,N_4222);
xnor U4633 (N_4633,N_4492,N_4200);
nand U4634 (N_4634,N_4479,N_4299);
nand U4635 (N_4635,N_4449,N_4258);
nor U4636 (N_4636,N_4309,N_4287);
nand U4637 (N_4637,N_4416,N_4270);
or U4638 (N_4638,N_4368,N_4255);
or U4639 (N_4639,N_4308,N_4407);
xnor U4640 (N_4640,N_4284,N_4265);
xnor U4641 (N_4641,N_4459,N_4384);
and U4642 (N_4642,N_4370,N_4376);
nor U4643 (N_4643,N_4378,N_4349);
or U4644 (N_4644,N_4404,N_4435);
or U4645 (N_4645,N_4453,N_4266);
and U4646 (N_4646,N_4209,N_4302);
xor U4647 (N_4647,N_4329,N_4283);
or U4648 (N_4648,N_4352,N_4424);
nor U4649 (N_4649,N_4228,N_4337);
and U4650 (N_4650,N_4250,N_4258);
nor U4651 (N_4651,N_4203,N_4299);
nor U4652 (N_4652,N_4422,N_4213);
and U4653 (N_4653,N_4428,N_4255);
and U4654 (N_4654,N_4284,N_4377);
or U4655 (N_4655,N_4316,N_4442);
nor U4656 (N_4656,N_4488,N_4217);
nand U4657 (N_4657,N_4250,N_4448);
nor U4658 (N_4658,N_4416,N_4302);
and U4659 (N_4659,N_4321,N_4281);
nor U4660 (N_4660,N_4404,N_4240);
and U4661 (N_4661,N_4237,N_4396);
nor U4662 (N_4662,N_4299,N_4239);
nor U4663 (N_4663,N_4340,N_4487);
nor U4664 (N_4664,N_4282,N_4275);
nand U4665 (N_4665,N_4467,N_4418);
or U4666 (N_4666,N_4261,N_4313);
xnor U4667 (N_4667,N_4498,N_4321);
or U4668 (N_4668,N_4438,N_4398);
xor U4669 (N_4669,N_4418,N_4465);
or U4670 (N_4670,N_4253,N_4356);
nor U4671 (N_4671,N_4243,N_4313);
xor U4672 (N_4672,N_4410,N_4306);
or U4673 (N_4673,N_4297,N_4320);
xnor U4674 (N_4674,N_4245,N_4382);
and U4675 (N_4675,N_4469,N_4497);
xnor U4676 (N_4676,N_4359,N_4490);
or U4677 (N_4677,N_4446,N_4431);
and U4678 (N_4678,N_4341,N_4450);
nand U4679 (N_4679,N_4494,N_4402);
xor U4680 (N_4680,N_4246,N_4450);
or U4681 (N_4681,N_4444,N_4497);
and U4682 (N_4682,N_4372,N_4352);
and U4683 (N_4683,N_4227,N_4407);
nor U4684 (N_4684,N_4452,N_4411);
or U4685 (N_4685,N_4426,N_4249);
xnor U4686 (N_4686,N_4365,N_4397);
xor U4687 (N_4687,N_4426,N_4402);
or U4688 (N_4688,N_4331,N_4380);
and U4689 (N_4689,N_4267,N_4466);
or U4690 (N_4690,N_4287,N_4337);
xnor U4691 (N_4691,N_4479,N_4324);
and U4692 (N_4692,N_4240,N_4374);
nor U4693 (N_4693,N_4247,N_4444);
nor U4694 (N_4694,N_4455,N_4407);
nor U4695 (N_4695,N_4234,N_4235);
xor U4696 (N_4696,N_4325,N_4250);
nor U4697 (N_4697,N_4412,N_4409);
and U4698 (N_4698,N_4402,N_4260);
xor U4699 (N_4699,N_4337,N_4421);
and U4700 (N_4700,N_4386,N_4389);
nor U4701 (N_4701,N_4493,N_4360);
nor U4702 (N_4702,N_4345,N_4430);
xor U4703 (N_4703,N_4489,N_4236);
and U4704 (N_4704,N_4451,N_4369);
nand U4705 (N_4705,N_4318,N_4443);
xor U4706 (N_4706,N_4465,N_4276);
xor U4707 (N_4707,N_4249,N_4494);
and U4708 (N_4708,N_4401,N_4390);
and U4709 (N_4709,N_4406,N_4417);
and U4710 (N_4710,N_4378,N_4221);
nor U4711 (N_4711,N_4366,N_4405);
and U4712 (N_4712,N_4268,N_4216);
nor U4713 (N_4713,N_4410,N_4219);
nand U4714 (N_4714,N_4245,N_4302);
nor U4715 (N_4715,N_4319,N_4468);
nand U4716 (N_4716,N_4253,N_4321);
xnor U4717 (N_4717,N_4269,N_4215);
or U4718 (N_4718,N_4323,N_4408);
and U4719 (N_4719,N_4413,N_4284);
xnor U4720 (N_4720,N_4367,N_4359);
and U4721 (N_4721,N_4276,N_4352);
nor U4722 (N_4722,N_4236,N_4356);
xor U4723 (N_4723,N_4436,N_4277);
nor U4724 (N_4724,N_4487,N_4314);
and U4725 (N_4725,N_4357,N_4203);
nor U4726 (N_4726,N_4468,N_4403);
or U4727 (N_4727,N_4377,N_4382);
or U4728 (N_4728,N_4238,N_4355);
xnor U4729 (N_4729,N_4487,N_4446);
xnor U4730 (N_4730,N_4313,N_4395);
nand U4731 (N_4731,N_4494,N_4355);
and U4732 (N_4732,N_4410,N_4398);
nand U4733 (N_4733,N_4371,N_4455);
or U4734 (N_4734,N_4302,N_4347);
and U4735 (N_4735,N_4345,N_4357);
and U4736 (N_4736,N_4496,N_4318);
nor U4737 (N_4737,N_4245,N_4293);
nand U4738 (N_4738,N_4417,N_4221);
or U4739 (N_4739,N_4258,N_4432);
or U4740 (N_4740,N_4468,N_4388);
or U4741 (N_4741,N_4222,N_4315);
nand U4742 (N_4742,N_4381,N_4217);
xor U4743 (N_4743,N_4492,N_4305);
or U4744 (N_4744,N_4211,N_4488);
and U4745 (N_4745,N_4431,N_4228);
xnor U4746 (N_4746,N_4434,N_4446);
nor U4747 (N_4747,N_4407,N_4484);
xor U4748 (N_4748,N_4217,N_4462);
or U4749 (N_4749,N_4460,N_4254);
xor U4750 (N_4750,N_4362,N_4454);
or U4751 (N_4751,N_4499,N_4455);
or U4752 (N_4752,N_4204,N_4303);
and U4753 (N_4753,N_4373,N_4496);
nand U4754 (N_4754,N_4227,N_4485);
nand U4755 (N_4755,N_4389,N_4392);
and U4756 (N_4756,N_4233,N_4306);
or U4757 (N_4757,N_4347,N_4211);
or U4758 (N_4758,N_4215,N_4235);
xor U4759 (N_4759,N_4467,N_4464);
or U4760 (N_4760,N_4364,N_4244);
and U4761 (N_4761,N_4213,N_4276);
and U4762 (N_4762,N_4426,N_4480);
or U4763 (N_4763,N_4399,N_4309);
nand U4764 (N_4764,N_4435,N_4375);
or U4765 (N_4765,N_4371,N_4394);
or U4766 (N_4766,N_4369,N_4422);
nor U4767 (N_4767,N_4350,N_4465);
nor U4768 (N_4768,N_4263,N_4416);
xor U4769 (N_4769,N_4335,N_4338);
xor U4770 (N_4770,N_4276,N_4380);
xnor U4771 (N_4771,N_4421,N_4465);
nand U4772 (N_4772,N_4307,N_4412);
nor U4773 (N_4773,N_4279,N_4243);
xnor U4774 (N_4774,N_4446,N_4344);
and U4775 (N_4775,N_4220,N_4418);
nor U4776 (N_4776,N_4461,N_4200);
nor U4777 (N_4777,N_4399,N_4454);
nor U4778 (N_4778,N_4427,N_4417);
or U4779 (N_4779,N_4442,N_4407);
and U4780 (N_4780,N_4326,N_4291);
and U4781 (N_4781,N_4294,N_4330);
or U4782 (N_4782,N_4251,N_4302);
or U4783 (N_4783,N_4346,N_4286);
xnor U4784 (N_4784,N_4451,N_4248);
nor U4785 (N_4785,N_4468,N_4386);
nand U4786 (N_4786,N_4328,N_4332);
xnor U4787 (N_4787,N_4446,N_4290);
or U4788 (N_4788,N_4233,N_4227);
and U4789 (N_4789,N_4393,N_4201);
xnor U4790 (N_4790,N_4289,N_4479);
or U4791 (N_4791,N_4288,N_4397);
nor U4792 (N_4792,N_4258,N_4262);
and U4793 (N_4793,N_4214,N_4348);
and U4794 (N_4794,N_4256,N_4371);
xnor U4795 (N_4795,N_4373,N_4275);
nor U4796 (N_4796,N_4436,N_4343);
nor U4797 (N_4797,N_4394,N_4427);
or U4798 (N_4798,N_4455,N_4250);
and U4799 (N_4799,N_4448,N_4367);
nor U4800 (N_4800,N_4728,N_4638);
or U4801 (N_4801,N_4733,N_4695);
or U4802 (N_4802,N_4657,N_4783);
nor U4803 (N_4803,N_4753,N_4773);
nand U4804 (N_4804,N_4745,N_4519);
and U4805 (N_4805,N_4570,N_4748);
and U4806 (N_4806,N_4505,N_4545);
nor U4807 (N_4807,N_4744,N_4617);
xnor U4808 (N_4808,N_4501,N_4633);
nand U4809 (N_4809,N_4698,N_4788);
and U4810 (N_4810,N_4732,N_4701);
or U4811 (N_4811,N_4680,N_4572);
nor U4812 (N_4812,N_4613,N_4781);
and U4813 (N_4813,N_4604,N_4621);
xor U4814 (N_4814,N_4668,N_4500);
xor U4815 (N_4815,N_4567,N_4595);
nand U4816 (N_4816,N_4530,N_4535);
nand U4817 (N_4817,N_4622,N_4772);
nor U4818 (N_4818,N_4771,N_4768);
nor U4819 (N_4819,N_4533,N_4615);
or U4820 (N_4820,N_4606,N_4715);
and U4821 (N_4821,N_4758,N_4516);
xor U4822 (N_4822,N_4560,N_4511);
xor U4823 (N_4823,N_4710,N_4762);
nand U4824 (N_4824,N_4627,N_4760);
nor U4825 (N_4825,N_4655,N_4569);
nor U4826 (N_4826,N_4591,N_4648);
xnor U4827 (N_4827,N_4706,N_4713);
and U4828 (N_4828,N_4678,N_4704);
nand U4829 (N_4829,N_4580,N_4730);
nor U4830 (N_4830,N_4780,N_4746);
or U4831 (N_4831,N_4709,N_4663);
or U4832 (N_4832,N_4656,N_4540);
and U4833 (N_4833,N_4625,N_4679);
nor U4834 (N_4834,N_4575,N_4508);
xnor U4835 (N_4835,N_4798,N_4776);
xnor U4836 (N_4836,N_4611,N_4666);
nor U4837 (N_4837,N_4667,N_4630);
xnor U4838 (N_4838,N_4714,N_4671);
and U4839 (N_4839,N_4724,N_4660);
or U4840 (N_4840,N_4761,N_4644);
and U4841 (N_4841,N_4693,N_4587);
xnor U4842 (N_4842,N_4538,N_4589);
or U4843 (N_4843,N_4683,N_4782);
xnor U4844 (N_4844,N_4568,N_4509);
xnor U4845 (N_4845,N_4703,N_4662);
and U4846 (N_4846,N_4708,N_4791);
and U4847 (N_4847,N_4549,N_4598);
nand U4848 (N_4848,N_4619,N_4739);
xnor U4849 (N_4849,N_4643,N_4528);
nor U4850 (N_4850,N_4583,N_4723);
or U4851 (N_4851,N_4786,N_4716);
nor U4852 (N_4852,N_4717,N_4565);
nor U4853 (N_4853,N_4557,N_4562);
nand U4854 (N_4854,N_4659,N_4646);
xor U4855 (N_4855,N_4523,N_4690);
nand U4856 (N_4856,N_4614,N_4605);
or U4857 (N_4857,N_4684,N_4754);
and U4858 (N_4858,N_4766,N_4658);
and U4859 (N_4859,N_4521,N_4765);
nor U4860 (N_4860,N_4654,N_4741);
nor U4861 (N_4861,N_4696,N_4672);
and U4862 (N_4862,N_4647,N_4774);
nand U4863 (N_4863,N_4797,N_4669);
xnor U4864 (N_4864,N_4525,N_4594);
and U4865 (N_4865,N_4796,N_4737);
or U4866 (N_4866,N_4522,N_4725);
xnor U4867 (N_4867,N_4576,N_4534);
or U4868 (N_4868,N_4742,N_4585);
nand U4869 (N_4869,N_4721,N_4718);
nand U4870 (N_4870,N_4502,N_4531);
nand U4871 (N_4871,N_4513,N_4541);
xnor U4872 (N_4872,N_4778,N_4543);
or U4873 (N_4873,N_4558,N_4661);
xor U4874 (N_4874,N_4649,N_4665);
and U4875 (N_4875,N_4584,N_4601);
and U4876 (N_4876,N_4740,N_4504);
xnor U4877 (N_4877,N_4600,N_4793);
nor U4878 (N_4878,N_4510,N_4597);
or U4879 (N_4879,N_4574,N_4676);
or U4880 (N_4880,N_4712,N_4539);
and U4881 (N_4881,N_4554,N_4691);
nor U4882 (N_4882,N_4692,N_4707);
xor U4883 (N_4883,N_4563,N_4582);
nand U4884 (N_4884,N_4794,N_4542);
or U4885 (N_4885,N_4596,N_4686);
and U4886 (N_4886,N_4700,N_4790);
and U4887 (N_4887,N_4603,N_4720);
and U4888 (N_4888,N_4518,N_4722);
or U4889 (N_4889,N_4756,N_4694);
nor U4890 (N_4890,N_4705,N_4526);
and U4891 (N_4891,N_4593,N_4673);
xnor U4892 (N_4892,N_4677,N_4553);
or U4893 (N_4893,N_4607,N_4527);
nand U4894 (N_4894,N_4650,N_4629);
nand U4895 (N_4895,N_4685,N_4699);
nor U4896 (N_4896,N_4641,N_4799);
nand U4897 (N_4897,N_4620,N_4515);
and U4898 (N_4898,N_4512,N_4503);
or U4899 (N_4899,N_4750,N_4608);
xor U4900 (N_4900,N_4688,N_4586);
and U4901 (N_4901,N_4626,N_4551);
or U4902 (N_4902,N_4792,N_4616);
nor U4903 (N_4903,N_4759,N_4752);
nor U4904 (N_4904,N_4757,N_4581);
or U4905 (N_4905,N_4738,N_4555);
nand U4906 (N_4906,N_4634,N_4785);
and U4907 (N_4907,N_4651,N_4532);
xnor U4908 (N_4908,N_4653,N_4784);
xor U4909 (N_4909,N_4734,N_4751);
nand U4910 (N_4910,N_4578,N_4770);
xnor U4911 (N_4911,N_4609,N_4681);
or U4912 (N_4912,N_4719,N_4520);
xnor U4913 (N_4913,N_4727,N_4612);
nand U4914 (N_4914,N_4645,N_4763);
nand U4915 (N_4915,N_4624,N_4579);
nand U4916 (N_4916,N_4529,N_4637);
nand U4917 (N_4917,N_4636,N_4640);
and U4918 (N_4918,N_4590,N_4735);
nand U4919 (N_4919,N_4564,N_4670);
or U4920 (N_4920,N_4736,N_4729);
or U4921 (N_4921,N_4552,N_4599);
nor U4922 (N_4922,N_4544,N_4507);
nand U4923 (N_4923,N_4514,N_4743);
nor U4924 (N_4924,N_4546,N_4711);
and U4925 (N_4925,N_4697,N_4755);
nand U4926 (N_4926,N_4749,N_4524);
nand U4927 (N_4927,N_4547,N_4642);
xor U4928 (N_4928,N_4747,N_4639);
or U4929 (N_4929,N_4635,N_4702);
xnor U4930 (N_4930,N_4536,N_4537);
or U4931 (N_4931,N_4610,N_4777);
and U4932 (N_4932,N_4506,N_4588);
nor U4933 (N_4933,N_4618,N_4592);
nand U4934 (N_4934,N_4556,N_4764);
xor U4935 (N_4935,N_4559,N_4652);
and U4936 (N_4936,N_4726,N_4682);
xnor U4937 (N_4937,N_4628,N_4664);
and U4938 (N_4938,N_4689,N_4769);
nand U4939 (N_4939,N_4571,N_4602);
and U4940 (N_4940,N_4731,N_4631);
nor U4941 (N_4941,N_4561,N_4548);
and U4942 (N_4942,N_4550,N_4787);
nand U4943 (N_4943,N_4632,N_4674);
xor U4944 (N_4944,N_4623,N_4566);
or U4945 (N_4945,N_4795,N_4767);
nor U4946 (N_4946,N_4517,N_4687);
xor U4947 (N_4947,N_4779,N_4675);
nor U4948 (N_4948,N_4775,N_4573);
nand U4949 (N_4949,N_4577,N_4789);
or U4950 (N_4950,N_4764,N_4509);
xor U4951 (N_4951,N_4778,N_4656);
and U4952 (N_4952,N_4666,N_4793);
xnor U4953 (N_4953,N_4581,N_4600);
xor U4954 (N_4954,N_4716,N_4617);
xnor U4955 (N_4955,N_4771,N_4717);
xor U4956 (N_4956,N_4509,N_4527);
nor U4957 (N_4957,N_4557,N_4798);
xnor U4958 (N_4958,N_4682,N_4548);
nor U4959 (N_4959,N_4619,N_4541);
and U4960 (N_4960,N_4662,N_4684);
or U4961 (N_4961,N_4734,N_4528);
xor U4962 (N_4962,N_4693,N_4555);
or U4963 (N_4963,N_4773,N_4680);
or U4964 (N_4964,N_4736,N_4731);
xor U4965 (N_4965,N_4520,N_4543);
nand U4966 (N_4966,N_4764,N_4584);
or U4967 (N_4967,N_4730,N_4654);
or U4968 (N_4968,N_4727,N_4557);
nand U4969 (N_4969,N_4574,N_4589);
or U4970 (N_4970,N_4524,N_4710);
nor U4971 (N_4971,N_4614,N_4751);
and U4972 (N_4972,N_4587,N_4782);
and U4973 (N_4973,N_4796,N_4653);
nand U4974 (N_4974,N_4505,N_4748);
or U4975 (N_4975,N_4612,N_4614);
xor U4976 (N_4976,N_4514,N_4753);
xnor U4977 (N_4977,N_4786,N_4703);
or U4978 (N_4978,N_4606,N_4571);
xor U4979 (N_4979,N_4516,N_4765);
or U4980 (N_4980,N_4762,N_4597);
nand U4981 (N_4981,N_4596,N_4529);
nor U4982 (N_4982,N_4632,N_4724);
xnor U4983 (N_4983,N_4703,N_4789);
or U4984 (N_4984,N_4559,N_4757);
and U4985 (N_4985,N_4509,N_4553);
xnor U4986 (N_4986,N_4527,N_4588);
xor U4987 (N_4987,N_4509,N_4656);
xnor U4988 (N_4988,N_4602,N_4613);
and U4989 (N_4989,N_4607,N_4566);
or U4990 (N_4990,N_4656,N_4630);
nand U4991 (N_4991,N_4630,N_4706);
nor U4992 (N_4992,N_4714,N_4692);
or U4993 (N_4993,N_4721,N_4709);
and U4994 (N_4994,N_4709,N_4542);
nand U4995 (N_4995,N_4789,N_4539);
nor U4996 (N_4996,N_4582,N_4579);
or U4997 (N_4997,N_4632,N_4660);
and U4998 (N_4998,N_4508,N_4676);
nand U4999 (N_4999,N_4748,N_4744);
nand U5000 (N_5000,N_4579,N_4679);
and U5001 (N_5001,N_4533,N_4636);
and U5002 (N_5002,N_4546,N_4567);
and U5003 (N_5003,N_4757,N_4793);
nor U5004 (N_5004,N_4731,N_4535);
nand U5005 (N_5005,N_4530,N_4773);
or U5006 (N_5006,N_4586,N_4582);
xor U5007 (N_5007,N_4634,N_4599);
and U5008 (N_5008,N_4769,N_4518);
nand U5009 (N_5009,N_4650,N_4739);
or U5010 (N_5010,N_4713,N_4672);
nand U5011 (N_5011,N_4714,N_4694);
nand U5012 (N_5012,N_4684,N_4582);
or U5013 (N_5013,N_4764,N_4599);
xor U5014 (N_5014,N_4785,N_4674);
xor U5015 (N_5015,N_4714,N_4667);
nand U5016 (N_5016,N_4676,N_4734);
nand U5017 (N_5017,N_4757,N_4739);
nor U5018 (N_5018,N_4574,N_4714);
or U5019 (N_5019,N_4692,N_4501);
xnor U5020 (N_5020,N_4739,N_4657);
xor U5021 (N_5021,N_4545,N_4523);
xnor U5022 (N_5022,N_4675,N_4636);
and U5023 (N_5023,N_4682,N_4689);
xor U5024 (N_5024,N_4668,N_4615);
nor U5025 (N_5025,N_4544,N_4794);
nand U5026 (N_5026,N_4576,N_4742);
or U5027 (N_5027,N_4675,N_4690);
or U5028 (N_5028,N_4592,N_4668);
and U5029 (N_5029,N_4517,N_4612);
nor U5030 (N_5030,N_4532,N_4670);
nor U5031 (N_5031,N_4681,N_4640);
or U5032 (N_5032,N_4529,N_4551);
nor U5033 (N_5033,N_4688,N_4635);
nor U5034 (N_5034,N_4765,N_4566);
nand U5035 (N_5035,N_4704,N_4777);
nor U5036 (N_5036,N_4656,N_4695);
or U5037 (N_5037,N_4507,N_4686);
xnor U5038 (N_5038,N_4518,N_4573);
nand U5039 (N_5039,N_4594,N_4774);
or U5040 (N_5040,N_4526,N_4583);
nand U5041 (N_5041,N_4516,N_4706);
xnor U5042 (N_5042,N_4582,N_4506);
and U5043 (N_5043,N_4774,N_4615);
xnor U5044 (N_5044,N_4554,N_4585);
and U5045 (N_5045,N_4740,N_4712);
nand U5046 (N_5046,N_4785,N_4775);
nor U5047 (N_5047,N_4548,N_4730);
or U5048 (N_5048,N_4502,N_4693);
nor U5049 (N_5049,N_4504,N_4781);
nand U5050 (N_5050,N_4690,N_4620);
xor U5051 (N_5051,N_4694,N_4631);
nor U5052 (N_5052,N_4619,N_4633);
and U5053 (N_5053,N_4723,N_4675);
or U5054 (N_5054,N_4522,N_4574);
nor U5055 (N_5055,N_4500,N_4773);
or U5056 (N_5056,N_4648,N_4642);
and U5057 (N_5057,N_4714,N_4681);
nor U5058 (N_5058,N_4765,N_4610);
and U5059 (N_5059,N_4707,N_4592);
nand U5060 (N_5060,N_4776,N_4762);
nor U5061 (N_5061,N_4525,N_4543);
xnor U5062 (N_5062,N_4791,N_4797);
or U5063 (N_5063,N_4638,N_4586);
nor U5064 (N_5064,N_4672,N_4515);
or U5065 (N_5065,N_4604,N_4656);
nor U5066 (N_5066,N_4777,N_4713);
and U5067 (N_5067,N_4542,N_4658);
nor U5068 (N_5068,N_4588,N_4774);
nand U5069 (N_5069,N_4527,N_4774);
nor U5070 (N_5070,N_4578,N_4653);
and U5071 (N_5071,N_4579,N_4661);
nor U5072 (N_5072,N_4712,N_4721);
nor U5073 (N_5073,N_4744,N_4670);
xnor U5074 (N_5074,N_4508,N_4632);
nand U5075 (N_5075,N_4582,N_4737);
nor U5076 (N_5076,N_4780,N_4596);
or U5077 (N_5077,N_4541,N_4582);
nor U5078 (N_5078,N_4511,N_4519);
nand U5079 (N_5079,N_4546,N_4721);
and U5080 (N_5080,N_4675,N_4583);
or U5081 (N_5081,N_4609,N_4707);
and U5082 (N_5082,N_4610,N_4609);
nor U5083 (N_5083,N_4720,N_4680);
and U5084 (N_5084,N_4631,N_4683);
and U5085 (N_5085,N_4682,N_4515);
nor U5086 (N_5086,N_4739,N_4694);
or U5087 (N_5087,N_4770,N_4782);
or U5088 (N_5088,N_4513,N_4769);
nand U5089 (N_5089,N_4559,N_4552);
and U5090 (N_5090,N_4729,N_4732);
nand U5091 (N_5091,N_4699,N_4545);
and U5092 (N_5092,N_4712,N_4789);
or U5093 (N_5093,N_4792,N_4510);
or U5094 (N_5094,N_4793,N_4585);
and U5095 (N_5095,N_4794,N_4687);
and U5096 (N_5096,N_4682,N_4722);
nand U5097 (N_5097,N_4576,N_4669);
xnor U5098 (N_5098,N_4750,N_4728);
and U5099 (N_5099,N_4561,N_4752);
or U5100 (N_5100,N_5016,N_4926);
and U5101 (N_5101,N_4906,N_4913);
nor U5102 (N_5102,N_4993,N_4944);
or U5103 (N_5103,N_4832,N_4857);
nand U5104 (N_5104,N_4883,N_4835);
or U5105 (N_5105,N_5055,N_5061);
and U5106 (N_5106,N_4921,N_4805);
xnor U5107 (N_5107,N_4964,N_4827);
or U5108 (N_5108,N_4822,N_4897);
and U5109 (N_5109,N_4927,N_5071);
nor U5110 (N_5110,N_4922,N_4890);
xor U5111 (N_5111,N_4963,N_4893);
xnor U5112 (N_5112,N_5081,N_4967);
or U5113 (N_5113,N_5072,N_4882);
nand U5114 (N_5114,N_4844,N_4877);
and U5115 (N_5115,N_5039,N_4974);
or U5116 (N_5116,N_4971,N_4986);
or U5117 (N_5117,N_4925,N_4816);
nor U5118 (N_5118,N_4901,N_5091);
nor U5119 (N_5119,N_4942,N_4969);
or U5120 (N_5120,N_4973,N_4841);
nor U5121 (N_5121,N_5022,N_5013);
nand U5122 (N_5122,N_5053,N_5080);
and U5123 (N_5123,N_5059,N_4938);
or U5124 (N_5124,N_5049,N_5074);
xnor U5125 (N_5125,N_4979,N_5032);
or U5126 (N_5126,N_4946,N_4888);
nand U5127 (N_5127,N_4898,N_5082);
nor U5128 (N_5128,N_5008,N_4982);
nor U5129 (N_5129,N_5078,N_4848);
xnor U5130 (N_5130,N_4998,N_5095);
nor U5131 (N_5131,N_5011,N_5030);
or U5132 (N_5132,N_4891,N_4989);
nor U5133 (N_5133,N_5034,N_5027);
or U5134 (N_5134,N_4930,N_4825);
and U5135 (N_5135,N_5067,N_5040);
xor U5136 (N_5136,N_4955,N_4916);
nor U5137 (N_5137,N_5010,N_4996);
nor U5138 (N_5138,N_5014,N_4934);
xnor U5139 (N_5139,N_5088,N_4854);
nor U5140 (N_5140,N_5000,N_4895);
and U5141 (N_5141,N_5066,N_4821);
xnor U5142 (N_5142,N_4988,N_4904);
nor U5143 (N_5143,N_5018,N_5073);
xor U5144 (N_5144,N_5003,N_4937);
nor U5145 (N_5145,N_5009,N_4800);
xnor U5146 (N_5146,N_5051,N_4894);
nor U5147 (N_5147,N_4912,N_4808);
nor U5148 (N_5148,N_5025,N_4802);
nor U5149 (N_5149,N_5038,N_4867);
or U5150 (N_5150,N_4811,N_4886);
xnor U5151 (N_5151,N_4943,N_5046);
or U5152 (N_5152,N_4876,N_4961);
xor U5153 (N_5153,N_4911,N_4960);
nor U5154 (N_5154,N_4815,N_4990);
and U5155 (N_5155,N_4952,N_5076);
xnor U5156 (N_5156,N_4928,N_4980);
nand U5157 (N_5157,N_4957,N_4917);
or U5158 (N_5158,N_4850,N_4845);
and U5159 (N_5159,N_4806,N_4863);
nor U5160 (N_5160,N_4813,N_5063);
and U5161 (N_5161,N_4887,N_4873);
nor U5162 (N_5162,N_5021,N_4981);
nand U5163 (N_5163,N_5075,N_4884);
nand U5164 (N_5164,N_4933,N_4871);
xor U5165 (N_5165,N_5047,N_4801);
nand U5166 (N_5166,N_4866,N_4999);
and U5167 (N_5167,N_4840,N_4966);
and U5168 (N_5168,N_5097,N_4860);
nand U5169 (N_5169,N_4918,N_5015);
and U5170 (N_5170,N_5065,N_4885);
and U5171 (N_5171,N_4948,N_4910);
nand U5172 (N_5172,N_5086,N_4995);
and U5173 (N_5173,N_5023,N_4945);
nor U5174 (N_5174,N_4941,N_5012);
and U5175 (N_5175,N_5099,N_5057);
or U5176 (N_5176,N_4932,N_5054);
nand U5177 (N_5177,N_4899,N_4983);
nand U5178 (N_5178,N_4819,N_4968);
nor U5179 (N_5179,N_4953,N_5083);
nand U5180 (N_5180,N_5019,N_4869);
and U5181 (N_5181,N_4829,N_5064);
or U5182 (N_5182,N_5045,N_4962);
nor U5183 (N_5183,N_4977,N_4929);
nor U5184 (N_5184,N_4812,N_4949);
nand U5185 (N_5185,N_4820,N_5093);
or U5186 (N_5186,N_4853,N_4889);
xor U5187 (N_5187,N_4839,N_4903);
and U5188 (N_5188,N_5001,N_4924);
xor U5189 (N_5189,N_4862,N_4909);
or U5190 (N_5190,N_4920,N_4900);
and U5191 (N_5191,N_5020,N_5068);
or U5192 (N_5192,N_4807,N_4915);
xor U5193 (N_5193,N_5017,N_5087);
nand U5194 (N_5194,N_5002,N_5050);
nand U5195 (N_5195,N_4809,N_4892);
nor U5196 (N_5196,N_4947,N_4936);
xor U5197 (N_5197,N_5062,N_4849);
and U5198 (N_5198,N_5077,N_4856);
or U5199 (N_5199,N_4939,N_4951);
and U5200 (N_5200,N_4975,N_4965);
xnor U5201 (N_5201,N_4843,N_5029);
or U5202 (N_5202,N_5090,N_4935);
nor U5203 (N_5203,N_4831,N_4830);
or U5204 (N_5204,N_4985,N_4838);
nor U5205 (N_5205,N_5058,N_4878);
nand U5206 (N_5206,N_5079,N_5094);
xor U5207 (N_5207,N_5004,N_4826);
and U5208 (N_5208,N_4880,N_4896);
nand U5209 (N_5209,N_4931,N_4905);
nand U5210 (N_5210,N_4864,N_4833);
nand U5211 (N_5211,N_4956,N_5024);
nand U5212 (N_5212,N_4954,N_5069);
xnor U5213 (N_5213,N_4847,N_5052);
xnor U5214 (N_5214,N_4870,N_4908);
nor U5215 (N_5215,N_4872,N_4976);
nand U5216 (N_5216,N_4834,N_5085);
nor U5217 (N_5217,N_4875,N_5098);
nor U5218 (N_5218,N_4902,N_4987);
or U5219 (N_5219,N_4919,N_4914);
nor U5220 (N_5220,N_4959,N_5092);
nand U5221 (N_5221,N_5033,N_4940);
nor U5222 (N_5222,N_4858,N_4804);
or U5223 (N_5223,N_5036,N_4859);
xor U5224 (N_5224,N_4852,N_4881);
or U5225 (N_5225,N_5044,N_4997);
or U5226 (N_5226,N_5048,N_4851);
and U5227 (N_5227,N_4814,N_4907);
or U5228 (N_5228,N_4950,N_4803);
xnor U5229 (N_5229,N_5089,N_5006);
nand U5230 (N_5230,N_4994,N_5096);
xnor U5231 (N_5231,N_5070,N_5043);
or U5232 (N_5232,N_4874,N_4836);
xor U5233 (N_5233,N_4879,N_4978);
xor U5234 (N_5234,N_4842,N_4817);
and U5235 (N_5235,N_5035,N_5056);
xor U5236 (N_5236,N_4991,N_4984);
or U5237 (N_5237,N_5026,N_4824);
nor U5238 (N_5238,N_4818,N_4992);
and U5239 (N_5239,N_5041,N_4810);
nand U5240 (N_5240,N_4958,N_5042);
nand U5241 (N_5241,N_5005,N_4861);
xnor U5242 (N_5242,N_4837,N_4823);
and U5243 (N_5243,N_5028,N_5037);
and U5244 (N_5244,N_5060,N_4846);
and U5245 (N_5245,N_5007,N_4972);
and U5246 (N_5246,N_5031,N_4855);
nand U5247 (N_5247,N_4865,N_4828);
xnor U5248 (N_5248,N_4923,N_4868);
xor U5249 (N_5249,N_5084,N_4970);
nor U5250 (N_5250,N_4922,N_4942);
xnor U5251 (N_5251,N_4913,N_5094);
and U5252 (N_5252,N_5012,N_5081);
nand U5253 (N_5253,N_4929,N_4890);
xor U5254 (N_5254,N_5002,N_4801);
or U5255 (N_5255,N_4968,N_4942);
nor U5256 (N_5256,N_5012,N_4839);
and U5257 (N_5257,N_4883,N_5006);
or U5258 (N_5258,N_4896,N_4962);
xnor U5259 (N_5259,N_4807,N_5075);
and U5260 (N_5260,N_4922,N_4808);
nand U5261 (N_5261,N_4983,N_4956);
nand U5262 (N_5262,N_4962,N_4918);
nand U5263 (N_5263,N_5000,N_4823);
xnor U5264 (N_5264,N_4922,N_4934);
nor U5265 (N_5265,N_4835,N_5073);
nand U5266 (N_5266,N_5010,N_4959);
and U5267 (N_5267,N_4805,N_5029);
or U5268 (N_5268,N_4824,N_4834);
nand U5269 (N_5269,N_4995,N_4911);
nor U5270 (N_5270,N_4850,N_5021);
or U5271 (N_5271,N_4901,N_5071);
and U5272 (N_5272,N_4962,N_4828);
and U5273 (N_5273,N_4853,N_5060);
nand U5274 (N_5274,N_4967,N_4991);
or U5275 (N_5275,N_4979,N_4980);
nand U5276 (N_5276,N_4843,N_4863);
xor U5277 (N_5277,N_4999,N_4989);
or U5278 (N_5278,N_4968,N_5029);
nor U5279 (N_5279,N_5090,N_4962);
nand U5280 (N_5280,N_4977,N_4923);
and U5281 (N_5281,N_4984,N_5016);
nand U5282 (N_5282,N_4902,N_5029);
and U5283 (N_5283,N_5097,N_4821);
nor U5284 (N_5284,N_4876,N_4868);
and U5285 (N_5285,N_5057,N_5049);
nor U5286 (N_5286,N_5088,N_5020);
xor U5287 (N_5287,N_5093,N_4947);
nor U5288 (N_5288,N_5046,N_5044);
or U5289 (N_5289,N_4819,N_4977);
and U5290 (N_5290,N_5047,N_5094);
nand U5291 (N_5291,N_4939,N_4839);
or U5292 (N_5292,N_4805,N_4971);
or U5293 (N_5293,N_4858,N_5083);
or U5294 (N_5294,N_4870,N_4922);
and U5295 (N_5295,N_4899,N_4994);
and U5296 (N_5296,N_5064,N_4828);
nand U5297 (N_5297,N_4824,N_4813);
nand U5298 (N_5298,N_4936,N_4872);
nor U5299 (N_5299,N_4841,N_4999);
nand U5300 (N_5300,N_4903,N_5036);
or U5301 (N_5301,N_5005,N_4850);
nor U5302 (N_5302,N_5015,N_4811);
and U5303 (N_5303,N_4871,N_4937);
or U5304 (N_5304,N_4902,N_4929);
or U5305 (N_5305,N_5077,N_4874);
nand U5306 (N_5306,N_4958,N_4957);
nand U5307 (N_5307,N_4816,N_4994);
nor U5308 (N_5308,N_4829,N_4893);
xnor U5309 (N_5309,N_5068,N_4963);
nand U5310 (N_5310,N_5022,N_4857);
and U5311 (N_5311,N_5003,N_4850);
or U5312 (N_5312,N_4825,N_4909);
and U5313 (N_5313,N_5056,N_4973);
nor U5314 (N_5314,N_5018,N_5028);
nand U5315 (N_5315,N_4991,N_5034);
or U5316 (N_5316,N_4841,N_5018);
and U5317 (N_5317,N_5069,N_5067);
or U5318 (N_5318,N_4865,N_5061);
and U5319 (N_5319,N_5084,N_4838);
and U5320 (N_5320,N_5078,N_4970);
or U5321 (N_5321,N_5071,N_4995);
nand U5322 (N_5322,N_4837,N_5060);
and U5323 (N_5323,N_5050,N_5061);
nand U5324 (N_5324,N_5067,N_5078);
or U5325 (N_5325,N_4998,N_4910);
nand U5326 (N_5326,N_4926,N_5058);
nor U5327 (N_5327,N_4968,N_5082);
and U5328 (N_5328,N_4985,N_4964);
nand U5329 (N_5329,N_4870,N_5035);
xnor U5330 (N_5330,N_4992,N_5071);
xor U5331 (N_5331,N_4908,N_4848);
nand U5332 (N_5332,N_5013,N_4949);
nor U5333 (N_5333,N_4867,N_4998);
or U5334 (N_5334,N_5032,N_4843);
and U5335 (N_5335,N_4882,N_4844);
nor U5336 (N_5336,N_5021,N_4989);
and U5337 (N_5337,N_5006,N_5001);
and U5338 (N_5338,N_5058,N_4888);
and U5339 (N_5339,N_4815,N_4944);
and U5340 (N_5340,N_4943,N_4821);
or U5341 (N_5341,N_5011,N_4976);
or U5342 (N_5342,N_4920,N_4837);
xor U5343 (N_5343,N_4911,N_4914);
nand U5344 (N_5344,N_5098,N_5009);
or U5345 (N_5345,N_4889,N_4847);
or U5346 (N_5346,N_4949,N_4995);
nor U5347 (N_5347,N_4927,N_5054);
nand U5348 (N_5348,N_4958,N_4885);
and U5349 (N_5349,N_4831,N_5009);
and U5350 (N_5350,N_5003,N_5022);
xnor U5351 (N_5351,N_5074,N_5062);
nand U5352 (N_5352,N_5041,N_5081);
xor U5353 (N_5353,N_4991,N_4985);
xnor U5354 (N_5354,N_4870,N_4996);
xor U5355 (N_5355,N_4800,N_4843);
nand U5356 (N_5356,N_4943,N_4808);
and U5357 (N_5357,N_4880,N_5010);
xor U5358 (N_5358,N_4882,N_4941);
or U5359 (N_5359,N_5011,N_5080);
or U5360 (N_5360,N_4865,N_4891);
and U5361 (N_5361,N_4929,N_4993);
nor U5362 (N_5362,N_4935,N_5057);
nor U5363 (N_5363,N_4956,N_4902);
nor U5364 (N_5364,N_5038,N_5096);
nand U5365 (N_5365,N_5045,N_5021);
or U5366 (N_5366,N_4810,N_4908);
or U5367 (N_5367,N_5042,N_4919);
nand U5368 (N_5368,N_4801,N_4955);
or U5369 (N_5369,N_4844,N_4868);
or U5370 (N_5370,N_4807,N_4948);
or U5371 (N_5371,N_5084,N_5011);
or U5372 (N_5372,N_4832,N_4841);
nor U5373 (N_5373,N_5049,N_4869);
and U5374 (N_5374,N_4872,N_4862);
xnor U5375 (N_5375,N_5032,N_5087);
xnor U5376 (N_5376,N_5006,N_4869);
nand U5377 (N_5377,N_5090,N_4998);
nand U5378 (N_5378,N_4886,N_4908);
or U5379 (N_5379,N_4820,N_4880);
and U5380 (N_5380,N_5084,N_4978);
nand U5381 (N_5381,N_5019,N_4961);
nand U5382 (N_5382,N_5023,N_4897);
or U5383 (N_5383,N_5097,N_4953);
nand U5384 (N_5384,N_4944,N_5002);
xnor U5385 (N_5385,N_5013,N_5049);
nand U5386 (N_5386,N_4925,N_4861);
and U5387 (N_5387,N_4926,N_4817);
nor U5388 (N_5388,N_5037,N_5041);
nor U5389 (N_5389,N_5060,N_4864);
nor U5390 (N_5390,N_4880,N_4838);
nor U5391 (N_5391,N_5058,N_4867);
and U5392 (N_5392,N_4900,N_4999);
nand U5393 (N_5393,N_4968,N_5067);
and U5394 (N_5394,N_4944,N_5057);
nand U5395 (N_5395,N_5021,N_4993);
or U5396 (N_5396,N_4948,N_4979);
nand U5397 (N_5397,N_4997,N_5043);
nand U5398 (N_5398,N_4948,N_5053);
xnor U5399 (N_5399,N_5023,N_4980);
nand U5400 (N_5400,N_5270,N_5357);
xnor U5401 (N_5401,N_5255,N_5201);
nand U5402 (N_5402,N_5240,N_5145);
xor U5403 (N_5403,N_5282,N_5301);
nand U5404 (N_5404,N_5109,N_5204);
nand U5405 (N_5405,N_5162,N_5186);
xnor U5406 (N_5406,N_5373,N_5298);
xnor U5407 (N_5407,N_5238,N_5356);
xnor U5408 (N_5408,N_5292,N_5169);
nand U5409 (N_5409,N_5268,N_5253);
nand U5410 (N_5410,N_5206,N_5300);
nand U5411 (N_5411,N_5329,N_5208);
xor U5412 (N_5412,N_5394,N_5260);
and U5413 (N_5413,N_5189,N_5199);
nor U5414 (N_5414,N_5223,N_5166);
xor U5415 (N_5415,N_5264,N_5303);
nand U5416 (N_5416,N_5227,N_5132);
nand U5417 (N_5417,N_5246,N_5221);
nor U5418 (N_5418,N_5274,N_5150);
and U5419 (N_5419,N_5249,N_5386);
nor U5420 (N_5420,N_5396,N_5348);
nor U5421 (N_5421,N_5231,N_5215);
nor U5422 (N_5422,N_5124,N_5216);
or U5423 (N_5423,N_5328,N_5237);
xor U5424 (N_5424,N_5239,N_5382);
or U5425 (N_5425,N_5290,N_5324);
and U5426 (N_5426,N_5359,N_5118);
xnor U5427 (N_5427,N_5320,N_5135);
nand U5428 (N_5428,N_5257,N_5331);
nor U5429 (N_5429,N_5280,N_5106);
nand U5430 (N_5430,N_5306,N_5397);
or U5431 (N_5431,N_5287,N_5136);
and U5432 (N_5432,N_5165,N_5273);
nor U5433 (N_5433,N_5307,N_5358);
nor U5434 (N_5434,N_5338,N_5281);
nor U5435 (N_5435,N_5304,N_5376);
xor U5436 (N_5436,N_5266,N_5184);
nand U5437 (N_5437,N_5291,N_5177);
xor U5438 (N_5438,N_5374,N_5148);
or U5439 (N_5439,N_5326,N_5387);
and U5440 (N_5440,N_5360,N_5188);
and U5441 (N_5441,N_5213,N_5198);
nor U5442 (N_5442,N_5289,N_5119);
or U5443 (N_5443,N_5335,N_5114);
xor U5444 (N_5444,N_5366,N_5267);
xor U5445 (N_5445,N_5183,N_5134);
nand U5446 (N_5446,N_5353,N_5380);
nor U5447 (N_5447,N_5234,N_5196);
xnor U5448 (N_5448,N_5179,N_5247);
xor U5449 (N_5449,N_5113,N_5158);
xor U5450 (N_5450,N_5277,N_5341);
nor U5451 (N_5451,N_5317,N_5195);
or U5452 (N_5452,N_5236,N_5310);
nand U5453 (N_5453,N_5308,N_5147);
nor U5454 (N_5454,N_5286,N_5296);
and U5455 (N_5455,N_5284,N_5211);
and U5456 (N_5456,N_5214,N_5283);
nor U5457 (N_5457,N_5342,N_5302);
or U5458 (N_5458,N_5173,N_5288);
or U5459 (N_5459,N_5220,N_5226);
or U5460 (N_5460,N_5346,N_5171);
xnor U5461 (N_5461,N_5137,N_5276);
xor U5462 (N_5462,N_5131,N_5154);
nand U5463 (N_5463,N_5365,N_5168);
xnor U5464 (N_5464,N_5368,N_5212);
and U5465 (N_5465,N_5232,N_5285);
or U5466 (N_5466,N_5252,N_5385);
and U5467 (N_5467,N_5130,N_5269);
nand U5468 (N_5468,N_5182,N_5122);
nor U5469 (N_5469,N_5101,N_5295);
and U5470 (N_5470,N_5125,N_5369);
xor U5471 (N_5471,N_5210,N_5332);
or U5472 (N_5472,N_5367,N_5395);
nor U5473 (N_5473,N_5399,N_5325);
nor U5474 (N_5474,N_5319,N_5334);
nor U5475 (N_5475,N_5265,N_5343);
nand U5476 (N_5476,N_5108,N_5248);
nor U5477 (N_5477,N_5129,N_5141);
nor U5478 (N_5478,N_5192,N_5185);
xor U5479 (N_5479,N_5263,N_5259);
and U5480 (N_5480,N_5398,N_5378);
xor U5481 (N_5481,N_5163,N_5327);
nor U5482 (N_5482,N_5350,N_5202);
nor U5483 (N_5483,N_5294,N_5377);
and U5484 (N_5484,N_5293,N_5272);
xor U5485 (N_5485,N_5143,N_5244);
nand U5486 (N_5486,N_5224,N_5250);
nand U5487 (N_5487,N_5381,N_5314);
nand U5488 (N_5488,N_5279,N_5205);
xor U5489 (N_5489,N_5209,N_5391);
and U5490 (N_5490,N_5242,N_5116);
or U5491 (N_5491,N_5389,N_5364);
nand U5492 (N_5492,N_5172,N_5339);
nor U5493 (N_5493,N_5133,N_5336);
or U5494 (N_5494,N_5103,N_5174);
and U5495 (N_5495,N_5383,N_5243);
xnor U5496 (N_5496,N_5340,N_5271);
and U5497 (N_5497,N_5371,N_5180);
nand U5498 (N_5498,N_5161,N_5126);
nor U5499 (N_5499,N_5379,N_5318);
and U5500 (N_5500,N_5225,N_5297);
nand U5501 (N_5501,N_5384,N_5102);
nand U5502 (N_5502,N_5390,N_5194);
and U5503 (N_5503,N_5152,N_5170);
and U5504 (N_5504,N_5363,N_5191);
or U5505 (N_5505,N_5347,N_5393);
or U5506 (N_5506,N_5352,N_5313);
and U5507 (N_5507,N_5207,N_5228);
and U5508 (N_5508,N_5230,N_5120);
and U5509 (N_5509,N_5190,N_5218);
nand U5510 (N_5510,N_5159,N_5123);
or U5511 (N_5511,N_5181,N_5261);
xnor U5512 (N_5512,N_5354,N_5117);
xnor U5513 (N_5513,N_5128,N_5157);
or U5514 (N_5514,N_5309,N_5375);
xnor U5515 (N_5515,N_5256,N_5251);
and U5516 (N_5516,N_5321,N_5355);
nand U5517 (N_5517,N_5362,N_5110);
and U5518 (N_5518,N_5151,N_5388);
nor U5519 (N_5519,N_5254,N_5241);
nand U5520 (N_5520,N_5217,N_5315);
and U5521 (N_5521,N_5258,N_5138);
nor U5522 (N_5522,N_5262,N_5193);
and U5523 (N_5523,N_5229,N_5146);
and U5524 (N_5524,N_5197,N_5345);
and U5525 (N_5525,N_5219,N_5370);
or U5526 (N_5526,N_5153,N_5105);
nand U5527 (N_5527,N_5155,N_5222);
or U5528 (N_5528,N_5149,N_5316);
xnor U5529 (N_5529,N_5176,N_5344);
xnor U5530 (N_5530,N_5361,N_5203);
nor U5531 (N_5531,N_5178,N_5278);
xor U5532 (N_5532,N_5140,N_5323);
or U5533 (N_5533,N_5349,N_5333);
and U5534 (N_5534,N_5233,N_5104);
nor U5535 (N_5535,N_5112,N_5322);
nand U5536 (N_5536,N_5311,N_5121);
nand U5537 (N_5537,N_5330,N_5111);
or U5538 (N_5538,N_5100,N_5312);
nor U5539 (N_5539,N_5144,N_5164);
or U5540 (N_5540,N_5245,N_5160);
or U5541 (N_5541,N_5305,N_5175);
and U5542 (N_5542,N_5127,N_5275);
xnor U5543 (N_5543,N_5392,N_5299);
and U5544 (N_5544,N_5372,N_5351);
or U5545 (N_5545,N_5167,N_5107);
and U5546 (N_5546,N_5337,N_5200);
xnor U5547 (N_5547,N_5142,N_5156);
xor U5548 (N_5548,N_5187,N_5139);
and U5549 (N_5549,N_5235,N_5115);
xor U5550 (N_5550,N_5310,N_5203);
and U5551 (N_5551,N_5132,N_5121);
or U5552 (N_5552,N_5170,N_5293);
nand U5553 (N_5553,N_5150,N_5337);
and U5554 (N_5554,N_5261,N_5121);
nor U5555 (N_5555,N_5276,N_5131);
nand U5556 (N_5556,N_5303,N_5312);
and U5557 (N_5557,N_5151,N_5275);
nand U5558 (N_5558,N_5234,N_5208);
nor U5559 (N_5559,N_5142,N_5194);
or U5560 (N_5560,N_5334,N_5123);
or U5561 (N_5561,N_5347,N_5387);
and U5562 (N_5562,N_5269,N_5235);
nor U5563 (N_5563,N_5150,N_5178);
or U5564 (N_5564,N_5143,N_5182);
and U5565 (N_5565,N_5161,N_5366);
nor U5566 (N_5566,N_5177,N_5126);
nor U5567 (N_5567,N_5390,N_5171);
and U5568 (N_5568,N_5203,N_5204);
and U5569 (N_5569,N_5182,N_5356);
or U5570 (N_5570,N_5274,N_5117);
xor U5571 (N_5571,N_5208,N_5231);
nand U5572 (N_5572,N_5182,N_5325);
or U5573 (N_5573,N_5173,N_5251);
and U5574 (N_5574,N_5266,N_5191);
or U5575 (N_5575,N_5103,N_5117);
or U5576 (N_5576,N_5374,N_5337);
or U5577 (N_5577,N_5311,N_5330);
and U5578 (N_5578,N_5171,N_5242);
xnor U5579 (N_5579,N_5386,N_5255);
xnor U5580 (N_5580,N_5342,N_5114);
nand U5581 (N_5581,N_5141,N_5259);
xnor U5582 (N_5582,N_5228,N_5358);
xnor U5583 (N_5583,N_5164,N_5208);
nand U5584 (N_5584,N_5355,N_5186);
nor U5585 (N_5585,N_5103,N_5356);
or U5586 (N_5586,N_5398,N_5177);
nand U5587 (N_5587,N_5325,N_5176);
xor U5588 (N_5588,N_5341,N_5176);
nor U5589 (N_5589,N_5296,N_5394);
nor U5590 (N_5590,N_5123,N_5307);
or U5591 (N_5591,N_5216,N_5383);
nor U5592 (N_5592,N_5235,N_5295);
or U5593 (N_5593,N_5103,N_5386);
nand U5594 (N_5594,N_5130,N_5247);
nor U5595 (N_5595,N_5178,N_5246);
and U5596 (N_5596,N_5281,N_5271);
or U5597 (N_5597,N_5200,N_5398);
nor U5598 (N_5598,N_5115,N_5285);
nor U5599 (N_5599,N_5359,N_5293);
and U5600 (N_5600,N_5180,N_5390);
xnor U5601 (N_5601,N_5199,N_5168);
nor U5602 (N_5602,N_5317,N_5256);
xor U5603 (N_5603,N_5236,N_5314);
or U5604 (N_5604,N_5108,N_5254);
xor U5605 (N_5605,N_5337,N_5389);
or U5606 (N_5606,N_5189,N_5188);
and U5607 (N_5607,N_5203,N_5112);
nor U5608 (N_5608,N_5361,N_5344);
nor U5609 (N_5609,N_5342,N_5326);
nand U5610 (N_5610,N_5258,N_5117);
nor U5611 (N_5611,N_5209,N_5311);
or U5612 (N_5612,N_5138,N_5211);
and U5613 (N_5613,N_5366,N_5396);
nor U5614 (N_5614,N_5242,N_5358);
nand U5615 (N_5615,N_5324,N_5245);
nand U5616 (N_5616,N_5290,N_5153);
xnor U5617 (N_5617,N_5153,N_5134);
or U5618 (N_5618,N_5127,N_5265);
or U5619 (N_5619,N_5171,N_5342);
nor U5620 (N_5620,N_5332,N_5266);
and U5621 (N_5621,N_5294,N_5207);
or U5622 (N_5622,N_5218,N_5162);
or U5623 (N_5623,N_5328,N_5241);
and U5624 (N_5624,N_5133,N_5265);
and U5625 (N_5625,N_5184,N_5110);
or U5626 (N_5626,N_5214,N_5364);
xnor U5627 (N_5627,N_5138,N_5159);
and U5628 (N_5628,N_5129,N_5307);
nand U5629 (N_5629,N_5265,N_5157);
xor U5630 (N_5630,N_5388,N_5103);
xnor U5631 (N_5631,N_5296,N_5216);
xor U5632 (N_5632,N_5398,N_5347);
xnor U5633 (N_5633,N_5387,N_5339);
xnor U5634 (N_5634,N_5382,N_5326);
xnor U5635 (N_5635,N_5208,N_5374);
and U5636 (N_5636,N_5394,N_5355);
or U5637 (N_5637,N_5150,N_5149);
nand U5638 (N_5638,N_5280,N_5122);
and U5639 (N_5639,N_5206,N_5256);
nand U5640 (N_5640,N_5381,N_5299);
xor U5641 (N_5641,N_5169,N_5321);
nand U5642 (N_5642,N_5195,N_5374);
nor U5643 (N_5643,N_5259,N_5330);
nand U5644 (N_5644,N_5105,N_5392);
nand U5645 (N_5645,N_5117,N_5114);
xor U5646 (N_5646,N_5383,N_5183);
xnor U5647 (N_5647,N_5215,N_5292);
nor U5648 (N_5648,N_5129,N_5246);
and U5649 (N_5649,N_5294,N_5393);
and U5650 (N_5650,N_5267,N_5149);
and U5651 (N_5651,N_5285,N_5348);
and U5652 (N_5652,N_5201,N_5149);
and U5653 (N_5653,N_5325,N_5221);
nor U5654 (N_5654,N_5239,N_5103);
or U5655 (N_5655,N_5199,N_5212);
or U5656 (N_5656,N_5333,N_5238);
or U5657 (N_5657,N_5388,N_5243);
or U5658 (N_5658,N_5375,N_5389);
or U5659 (N_5659,N_5248,N_5376);
xnor U5660 (N_5660,N_5327,N_5310);
nand U5661 (N_5661,N_5342,N_5188);
nand U5662 (N_5662,N_5243,N_5292);
nor U5663 (N_5663,N_5389,N_5299);
or U5664 (N_5664,N_5106,N_5399);
nor U5665 (N_5665,N_5382,N_5399);
xnor U5666 (N_5666,N_5355,N_5172);
or U5667 (N_5667,N_5136,N_5295);
and U5668 (N_5668,N_5326,N_5235);
or U5669 (N_5669,N_5213,N_5215);
and U5670 (N_5670,N_5320,N_5333);
nand U5671 (N_5671,N_5346,N_5365);
nor U5672 (N_5672,N_5152,N_5367);
nand U5673 (N_5673,N_5226,N_5207);
xor U5674 (N_5674,N_5191,N_5375);
nand U5675 (N_5675,N_5239,N_5325);
and U5676 (N_5676,N_5385,N_5382);
xor U5677 (N_5677,N_5392,N_5126);
xor U5678 (N_5678,N_5230,N_5139);
xor U5679 (N_5679,N_5231,N_5124);
nor U5680 (N_5680,N_5312,N_5223);
nand U5681 (N_5681,N_5233,N_5193);
or U5682 (N_5682,N_5327,N_5364);
nand U5683 (N_5683,N_5382,N_5161);
or U5684 (N_5684,N_5285,N_5394);
xnor U5685 (N_5685,N_5290,N_5225);
and U5686 (N_5686,N_5226,N_5187);
nand U5687 (N_5687,N_5170,N_5340);
and U5688 (N_5688,N_5218,N_5254);
nor U5689 (N_5689,N_5378,N_5244);
xor U5690 (N_5690,N_5314,N_5389);
or U5691 (N_5691,N_5115,N_5342);
or U5692 (N_5692,N_5233,N_5137);
nor U5693 (N_5693,N_5294,N_5270);
xnor U5694 (N_5694,N_5209,N_5241);
nand U5695 (N_5695,N_5332,N_5181);
nand U5696 (N_5696,N_5354,N_5277);
nand U5697 (N_5697,N_5214,N_5325);
or U5698 (N_5698,N_5152,N_5309);
nor U5699 (N_5699,N_5349,N_5212);
and U5700 (N_5700,N_5483,N_5489);
and U5701 (N_5701,N_5665,N_5473);
nand U5702 (N_5702,N_5551,N_5550);
xnor U5703 (N_5703,N_5617,N_5457);
xnor U5704 (N_5704,N_5479,N_5581);
or U5705 (N_5705,N_5415,N_5436);
xnor U5706 (N_5706,N_5677,N_5521);
xnor U5707 (N_5707,N_5609,N_5655);
or U5708 (N_5708,N_5538,N_5624);
nand U5709 (N_5709,N_5578,N_5498);
xnor U5710 (N_5710,N_5650,N_5645);
xnor U5711 (N_5711,N_5611,N_5475);
and U5712 (N_5712,N_5603,N_5675);
and U5713 (N_5713,N_5541,N_5607);
nor U5714 (N_5714,N_5422,N_5461);
nor U5715 (N_5715,N_5558,N_5486);
nand U5716 (N_5716,N_5574,N_5403);
xor U5717 (N_5717,N_5420,N_5582);
nor U5718 (N_5718,N_5456,N_5468);
nand U5719 (N_5719,N_5513,N_5608);
and U5720 (N_5720,N_5540,N_5549);
and U5721 (N_5721,N_5564,N_5671);
nand U5722 (N_5722,N_5480,N_5657);
nand U5723 (N_5723,N_5529,N_5565);
xnor U5724 (N_5724,N_5462,N_5628);
or U5725 (N_5725,N_5561,N_5517);
or U5726 (N_5726,N_5571,N_5459);
nand U5727 (N_5727,N_5482,N_5426);
nand U5728 (N_5728,N_5643,N_5566);
nand U5729 (N_5729,N_5694,N_5404);
nor U5730 (N_5730,N_5531,N_5474);
or U5731 (N_5731,N_5471,N_5514);
nor U5732 (N_5732,N_5556,N_5481);
or U5733 (N_5733,N_5451,N_5441);
nand U5734 (N_5734,N_5572,N_5661);
xor U5735 (N_5735,N_5535,N_5458);
and U5736 (N_5736,N_5445,N_5648);
nand U5737 (N_5737,N_5669,N_5635);
xor U5738 (N_5738,N_5476,N_5414);
and U5739 (N_5739,N_5522,N_5450);
or U5740 (N_5740,N_5681,N_5692);
nand U5741 (N_5741,N_5599,N_5424);
xor U5742 (N_5742,N_5478,N_5595);
or U5743 (N_5743,N_5680,N_5602);
or U5744 (N_5744,N_5591,N_5672);
nor U5745 (N_5745,N_5434,N_5567);
xor U5746 (N_5746,N_5697,N_5431);
nor U5747 (N_5747,N_5488,N_5670);
nand U5748 (N_5748,N_5658,N_5428);
nor U5749 (N_5749,N_5539,N_5570);
and U5750 (N_5750,N_5530,N_5637);
nor U5751 (N_5751,N_5412,N_5485);
nand U5752 (N_5752,N_5423,N_5644);
nand U5753 (N_5753,N_5686,N_5501);
and U5754 (N_5754,N_5506,N_5685);
xor U5755 (N_5755,N_5408,N_5532);
nand U5756 (N_5756,N_5469,N_5487);
and U5757 (N_5757,N_5548,N_5504);
nand U5758 (N_5758,N_5432,N_5573);
nor U5759 (N_5759,N_5484,N_5455);
nor U5760 (N_5760,N_5569,N_5555);
or U5761 (N_5761,N_5696,N_5663);
nor U5762 (N_5762,N_5491,N_5633);
nor U5763 (N_5763,N_5614,N_5597);
xnor U5764 (N_5764,N_5543,N_5647);
and U5765 (N_5765,N_5467,N_5401);
or U5766 (N_5766,N_5640,N_5575);
nor U5767 (N_5767,N_5623,N_5557);
or U5768 (N_5768,N_5494,N_5673);
or U5769 (N_5769,N_5547,N_5497);
nand U5770 (N_5770,N_5576,N_5579);
and U5771 (N_5771,N_5492,N_5642);
or U5772 (N_5772,N_5520,N_5620);
and U5773 (N_5773,N_5523,N_5600);
and U5774 (N_5774,N_5413,N_5430);
nor U5775 (N_5775,N_5463,N_5630);
and U5776 (N_5776,N_5664,N_5537);
xnor U5777 (N_5777,N_5683,N_5621);
and U5778 (N_5778,N_5405,N_5691);
nor U5779 (N_5779,N_5676,N_5583);
nor U5780 (N_5780,N_5553,N_5588);
xor U5781 (N_5781,N_5693,N_5418);
xor U5782 (N_5782,N_5448,N_5627);
nand U5783 (N_5783,N_5409,N_5667);
nand U5784 (N_5784,N_5622,N_5507);
nor U5785 (N_5785,N_5668,N_5687);
xor U5786 (N_5786,N_5638,N_5634);
nand U5787 (N_5787,N_5525,N_5610);
nand U5788 (N_5788,N_5496,N_5508);
nor U5789 (N_5789,N_5659,N_5552);
or U5790 (N_5790,N_5601,N_5612);
xnor U5791 (N_5791,N_5560,N_5690);
or U5792 (N_5792,N_5527,N_5562);
nor U5793 (N_5793,N_5400,N_5505);
or U5794 (N_5794,N_5613,N_5653);
nand U5795 (N_5795,N_5503,N_5619);
nor U5796 (N_5796,N_5545,N_5511);
and U5797 (N_5797,N_5587,N_5499);
xnor U5798 (N_5798,N_5534,N_5568);
xnor U5799 (N_5799,N_5449,N_5460);
or U5800 (N_5800,N_5447,N_5416);
nor U5801 (N_5801,N_5452,N_5689);
and U5802 (N_5802,N_5666,N_5586);
nor U5803 (N_5803,N_5407,N_5688);
xnor U5804 (N_5804,N_5429,N_5425);
xnor U5805 (N_5805,N_5698,N_5585);
xor U5806 (N_5806,N_5632,N_5629);
or U5807 (N_5807,N_5606,N_5699);
or U5808 (N_5808,N_5427,N_5631);
xnor U5809 (N_5809,N_5500,N_5626);
or U5810 (N_5810,N_5684,N_5584);
nand U5811 (N_5811,N_5616,N_5440);
nand U5812 (N_5812,N_5442,N_5516);
xor U5813 (N_5813,N_5554,N_5559);
and U5814 (N_5814,N_5411,N_5433);
nor U5815 (N_5815,N_5598,N_5510);
or U5816 (N_5816,N_5519,N_5641);
or U5817 (N_5817,N_5592,N_5596);
and U5818 (N_5818,N_5544,N_5615);
nor U5819 (N_5819,N_5493,N_5604);
or U5820 (N_5820,N_5660,N_5466);
and U5821 (N_5821,N_5649,N_5662);
nor U5822 (N_5822,N_5443,N_5651);
xor U5823 (N_5823,N_5464,N_5472);
and U5824 (N_5824,N_5682,N_5654);
nand U5825 (N_5825,N_5515,N_5590);
nand U5826 (N_5826,N_5402,N_5509);
and U5827 (N_5827,N_5437,N_5536);
or U5828 (N_5828,N_5639,N_5580);
and U5829 (N_5829,N_5546,N_5577);
nor U5830 (N_5830,N_5495,N_5477);
and U5831 (N_5831,N_5421,N_5674);
nand U5832 (N_5832,N_5605,N_5652);
nor U5833 (N_5833,N_5512,N_5524);
nor U5834 (N_5834,N_5453,N_5589);
or U5835 (N_5835,N_5695,N_5625);
nand U5836 (N_5836,N_5594,N_5528);
or U5837 (N_5837,N_5646,N_5470);
nor U5838 (N_5838,N_5618,N_5446);
nor U5839 (N_5839,N_5593,N_5656);
and U5840 (N_5840,N_5410,N_5444);
nor U5841 (N_5841,N_5679,N_5465);
or U5842 (N_5842,N_5526,N_5439);
xnor U5843 (N_5843,N_5417,N_5502);
nand U5844 (N_5844,N_5419,N_5563);
nand U5845 (N_5845,N_5438,N_5636);
nor U5846 (N_5846,N_5533,N_5678);
or U5847 (N_5847,N_5454,N_5490);
or U5848 (N_5848,N_5542,N_5435);
xor U5849 (N_5849,N_5406,N_5518);
and U5850 (N_5850,N_5455,N_5476);
or U5851 (N_5851,N_5624,N_5434);
or U5852 (N_5852,N_5401,N_5457);
and U5853 (N_5853,N_5506,N_5610);
or U5854 (N_5854,N_5420,N_5455);
nor U5855 (N_5855,N_5570,N_5441);
and U5856 (N_5856,N_5621,N_5676);
nor U5857 (N_5857,N_5519,N_5438);
nor U5858 (N_5858,N_5541,N_5676);
or U5859 (N_5859,N_5406,N_5402);
nand U5860 (N_5860,N_5414,N_5443);
xnor U5861 (N_5861,N_5543,N_5510);
nand U5862 (N_5862,N_5503,N_5550);
and U5863 (N_5863,N_5573,N_5551);
or U5864 (N_5864,N_5574,N_5504);
xnor U5865 (N_5865,N_5598,N_5491);
and U5866 (N_5866,N_5447,N_5465);
nor U5867 (N_5867,N_5429,N_5606);
nand U5868 (N_5868,N_5518,N_5657);
xor U5869 (N_5869,N_5481,N_5681);
or U5870 (N_5870,N_5414,N_5450);
or U5871 (N_5871,N_5483,N_5436);
nor U5872 (N_5872,N_5631,N_5586);
and U5873 (N_5873,N_5582,N_5579);
and U5874 (N_5874,N_5456,N_5629);
and U5875 (N_5875,N_5594,N_5468);
xnor U5876 (N_5876,N_5493,N_5650);
and U5877 (N_5877,N_5505,N_5613);
and U5878 (N_5878,N_5485,N_5620);
nor U5879 (N_5879,N_5476,N_5644);
nor U5880 (N_5880,N_5450,N_5451);
or U5881 (N_5881,N_5429,N_5418);
and U5882 (N_5882,N_5479,N_5565);
nor U5883 (N_5883,N_5510,N_5424);
nor U5884 (N_5884,N_5416,N_5470);
xnor U5885 (N_5885,N_5639,N_5557);
nand U5886 (N_5886,N_5606,N_5621);
and U5887 (N_5887,N_5507,N_5659);
xor U5888 (N_5888,N_5459,N_5512);
or U5889 (N_5889,N_5619,N_5568);
nor U5890 (N_5890,N_5529,N_5493);
nand U5891 (N_5891,N_5462,N_5686);
xnor U5892 (N_5892,N_5534,N_5618);
xnor U5893 (N_5893,N_5612,N_5465);
and U5894 (N_5894,N_5648,N_5615);
nand U5895 (N_5895,N_5419,N_5629);
or U5896 (N_5896,N_5573,N_5655);
nand U5897 (N_5897,N_5629,N_5575);
xnor U5898 (N_5898,N_5697,N_5648);
nand U5899 (N_5899,N_5461,N_5681);
or U5900 (N_5900,N_5494,N_5479);
and U5901 (N_5901,N_5475,N_5639);
and U5902 (N_5902,N_5538,N_5466);
and U5903 (N_5903,N_5687,N_5466);
or U5904 (N_5904,N_5541,N_5477);
and U5905 (N_5905,N_5615,N_5601);
and U5906 (N_5906,N_5522,N_5543);
xnor U5907 (N_5907,N_5461,N_5485);
xnor U5908 (N_5908,N_5650,N_5679);
nand U5909 (N_5909,N_5483,N_5611);
nand U5910 (N_5910,N_5678,N_5650);
and U5911 (N_5911,N_5638,N_5580);
nor U5912 (N_5912,N_5436,N_5428);
or U5913 (N_5913,N_5597,N_5626);
nor U5914 (N_5914,N_5640,N_5675);
and U5915 (N_5915,N_5550,N_5612);
nand U5916 (N_5916,N_5523,N_5691);
or U5917 (N_5917,N_5456,N_5571);
and U5918 (N_5918,N_5614,N_5629);
or U5919 (N_5919,N_5422,N_5547);
or U5920 (N_5920,N_5430,N_5581);
or U5921 (N_5921,N_5654,N_5588);
nor U5922 (N_5922,N_5655,N_5459);
nor U5923 (N_5923,N_5538,N_5449);
nor U5924 (N_5924,N_5552,N_5651);
and U5925 (N_5925,N_5671,N_5523);
nor U5926 (N_5926,N_5496,N_5416);
nor U5927 (N_5927,N_5684,N_5400);
nand U5928 (N_5928,N_5482,N_5693);
nor U5929 (N_5929,N_5626,N_5422);
nor U5930 (N_5930,N_5572,N_5692);
nand U5931 (N_5931,N_5448,N_5635);
or U5932 (N_5932,N_5654,N_5487);
xnor U5933 (N_5933,N_5511,N_5578);
or U5934 (N_5934,N_5487,N_5420);
and U5935 (N_5935,N_5501,N_5418);
and U5936 (N_5936,N_5581,N_5405);
or U5937 (N_5937,N_5689,N_5697);
nor U5938 (N_5938,N_5401,N_5476);
and U5939 (N_5939,N_5665,N_5510);
nand U5940 (N_5940,N_5567,N_5517);
nor U5941 (N_5941,N_5548,N_5632);
nand U5942 (N_5942,N_5626,N_5658);
nor U5943 (N_5943,N_5405,N_5516);
nor U5944 (N_5944,N_5437,N_5650);
nand U5945 (N_5945,N_5428,N_5674);
nor U5946 (N_5946,N_5458,N_5489);
or U5947 (N_5947,N_5679,N_5491);
or U5948 (N_5948,N_5589,N_5682);
nor U5949 (N_5949,N_5542,N_5583);
xnor U5950 (N_5950,N_5482,N_5447);
and U5951 (N_5951,N_5552,N_5632);
or U5952 (N_5952,N_5694,N_5498);
nor U5953 (N_5953,N_5579,N_5672);
or U5954 (N_5954,N_5494,N_5502);
or U5955 (N_5955,N_5596,N_5647);
nand U5956 (N_5956,N_5501,N_5576);
and U5957 (N_5957,N_5688,N_5654);
nor U5958 (N_5958,N_5478,N_5599);
nand U5959 (N_5959,N_5665,N_5628);
nand U5960 (N_5960,N_5559,N_5454);
nor U5961 (N_5961,N_5606,N_5590);
xor U5962 (N_5962,N_5492,N_5672);
nand U5963 (N_5963,N_5641,N_5415);
xor U5964 (N_5964,N_5617,N_5577);
xor U5965 (N_5965,N_5572,N_5666);
nand U5966 (N_5966,N_5485,N_5448);
xnor U5967 (N_5967,N_5539,N_5676);
and U5968 (N_5968,N_5696,N_5562);
nand U5969 (N_5969,N_5639,N_5436);
nor U5970 (N_5970,N_5623,N_5529);
or U5971 (N_5971,N_5473,N_5671);
xor U5972 (N_5972,N_5662,N_5457);
or U5973 (N_5973,N_5493,N_5593);
and U5974 (N_5974,N_5532,N_5417);
nor U5975 (N_5975,N_5504,N_5658);
and U5976 (N_5976,N_5466,N_5406);
and U5977 (N_5977,N_5475,N_5668);
and U5978 (N_5978,N_5462,N_5682);
nor U5979 (N_5979,N_5494,N_5528);
nor U5980 (N_5980,N_5532,N_5698);
nand U5981 (N_5981,N_5526,N_5658);
xor U5982 (N_5982,N_5502,N_5675);
nand U5983 (N_5983,N_5455,N_5561);
xor U5984 (N_5984,N_5617,N_5439);
xor U5985 (N_5985,N_5563,N_5509);
and U5986 (N_5986,N_5505,N_5604);
nor U5987 (N_5987,N_5455,N_5419);
nand U5988 (N_5988,N_5626,N_5566);
and U5989 (N_5989,N_5660,N_5548);
nand U5990 (N_5990,N_5460,N_5499);
nor U5991 (N_5991,N_5414,N_5682);
or U5992 (N_5992,N_5526,N_5690);
xnor U5993 (N_5993,N_5621,N_5470);
and U5994 (N_5994,N_5617,N_5495);
nand U5995 (N_5995,N_5598,N_5638);
xor U5996 (N_5996,N_5683,N_5662);
xnor U5997 (N_5997,N_5519,N_5507);
nand U5998 (N_5998,N_5567,N_5688);
xnor U5999 (N_5999,N_5562,N_5541);
or U6000 (N_6000,N_5904,N_5781);
and U6001 (N_6001,N_5818,N_5955);
or U6002 (N_6002,N_5712,N_5953);
and U6003 (N_6003,N_5881,N_5887);
and U6004 (N_6004,N_5724,N_5843);
xnor U6005 (N_6005,N_5876,N_5775);
nor U6006 (N_6006,N_5948,N_5758);
nor U6007 (N_6007,N_5812,N_5871);
and U6008 (N_6008,N_5717,N_5831);
nor U6009 (N_6009,N_5718,N_5845);
xor U6010 (N_6010,N_5857,N_5932);
and U6011 (N_6011,N_5872,N_5906);
nand U6012 (N_6012,N_5924,N_5709);
nor U6013 (N_6013,N_5913,N_5725);
nor U6014 (N_6014,N_5859,N_5752);
xnor U6015 (N_6015,N_5926,N_5982);
nor U6016 (N_6016,N_5707,N_5858);
xnor U6017 (N_6017,N_5706,N_5921);
and U6018 (N_6018,N_5715,N_5779);
or U6019 (N_6019,N_5894,N_5825);
xnor U6020 (N_6020,N_5957,N_5928);
nor U6021 (N_6021,N_5959,N_5844);
xor U6022 (N_6022,N_5973,N_5855);
xnor U6023 (N_6023,N_5999,N_5801);
xor U6024 (N_6024,N_5902,N_5942);
nor U6025 (N_6025,N_5726,N_5816);
and U6026 (N_6026,N_5991,N_5738);
nand U6027 (N_6027,N_5968,N_5927);
and U6028 (N_6028,N_5952,N_5977);
nor U6029 (N_6029,N_5979,N_5755);
xnor U6030 (N_6030,N_5842,N_5728);
nand U6031 (N_6031,N_5852,N_5923);
and U6032 (N_6032,N_5869,N_5838);
and U6033 (N_6033,N_5854,N_5804);
nor U6034 (N_6034,N_5848,N_5920);
or U6035 (N_6035,N_5877,N_5774);
xnor U6036 (N_6036,N_5811,N_5949);
xnor U6037 (N_6037,N_5787,N_5765);
nor U6038 (N_6038,N_5736,N_5886);
xor U6039 (N_6039,N_5783,N_5970);
nand U6040 (N_6040,N_5873,N_5967);
nor U6041 (N_6041,N_5864,N_5908);
and U6042 (N_6042,N_5965,N_5743);
or U6043 (N_6043,N_5986,N_5799);
and U6044 (N_6044,N_5897,N_5998);
nor U6045 (N_6045,N_5786,N_5943);
nand U6046 (N_6046,N_5958,N_5769);
nand U6047 (N_6047,N_5827,N_5883);
nor U6048 (N_6048,N_5807,N_5962);
nor U6049 (N_6049,N_5742,N_5810);
and U6050 (N_6050,N_5768,N_5996);
or U6051 (N_6051,N_5995,N_5780);
and U6052 (N_6052,N_5954,N_5898);
nand U6053 (N_6053,N_5803,N_5767);
nor U6054 (N_6054,N_5721,N_5992);
xnor U6055 (N_6055,N_5914,N_5817);
and U6056 (N_6056,N_5939,N_5740);
nand U6057 (N_6057,N_5701,N_5963);
nand U6058 (N_6058,N_5911,N_5824);
or U6059 (N_6059,N_5798,N_5806);
nand U6060 (N_6060,N_5981,N_5994);
xnor U6061 (N_6061,N_5713,N_5891);
or U6062 (N_6062,N_5744,N_5935);
nand U6063 (N_6063,N_5889,N_5940);
nand U6064 (N_6064,N_5761,N_5711);
and U6065 (N_6065,N_5915,N_5944);
xnor U6066 (N_6066,N_5792,N_5766);
or U6067 (N_6067,N_5989,N_5791);
and U6068 (N_6068,N_5951,N_5899);
or U6069 (N_6069,N_5764,N_5972);
or U6070 (N_6070,N_5978,N_5931);
or U6071 (N_6071,N_5947,N_5748);
xnor U6072 (N_6072,N_5704,N_5751);
or U6073 (N_6073,N_5735,N_5700);
and U6074 (N_6074,N_5909,N_5971);
xor U6075 (N_6075,N_5826,N_5985);
nand U6076 (N_6076,N_5878,N_5760);
or U6077 (N_6077,N_5884,N_5796);
and U6078 (N_6078,N_5793,N_5832);
xor U6079 (N_6079,N_5839,N_5819);
or U6080 (N_6080,N_5846,N_5917);
and U6081 (N_6081,N_5849,N_5934);
xnor U6082 (N_6082,N_5734,N_5987);
xnor U6083 (N_6083,N_5875,N_5770);
xor U6084 (N_6084,N_5893,N_5941);
nor U6085 (N_6085,N_5729,N_5772);
xnor U6086 (N_6086,N_5937,N_5933);
or U6087 (N_6087,N_5813,N_5702);
and U6088 (N_6088,N_5800,N_5809);
xor U6089 (N_6089,N_5722,N_5988);
and U6090 (N_6090,N_5851,N_5983);
nor U6091 (N_6091,N_5901,N_5762);
xor U6092 (N_6092,N_5732,N_5739);
and U6093 (N_6093,N_5910,N_5771);
and U6094 (N_6094,N_5874,N_5961);
and U6095 (N_6095,N_5745,N_5747);
xor U6096 (N_6096,N_5746,N_5716);
xor U6097 (N_6097,N_5710,N_5737);
xor U6098 (N_6098,N_5936,N_5823);
or U6099 (N_6099,N_5756,N_5853);
nand U6100 (N_6100,N_5856,N_5720);
and U6101 (N_6101,N_5863,N_5966);
nor U6102 (N_6102,N_5714,N_5794);
nand U6103 (N_6103,N_5990,N_5784);
nor U6104 (N_6104,N_5805,N_5834);
and U6105 (N_6105,N_5836,N_5922);
or U6106 (N_6106,N_5861,N_5750);
xor U6107 (N_6107,N_5895,N_5703);
nand U6108 (N_6108,N_5778,N_5829);
and U6109 (N_6109,N_5789,N_5929);
nor U6110 (N_6110,N_5782,N_5705);
xnor U6111 (N_6111,N_5993,N_5880);
nand U6112 (N_6112,N_5975,N_5860);
nor U6113 (N_6113,N_5916,N_5754);
nor U6114 (N_6114,N_5974,N_5723);
nor U6115 (N_6115,N_5984,N_5719);
or U6116 (N_6116,N_5892,N_5866);
nor U6117 (N_6117,N_5749,N_5945);
or U6118 (N_6118,N_5969,N_5896);
nand U6119 (N_6119,N_5960,N_5790);
nand U6120 (N_6120,N_5850,N_5814);
and U6121 (N_6121,N_5867,N_5733);
nand U6122 (N_6122,N_5882,N_5862);
nor U6123 (N_6123,N_5925,N_5788);
nand U6124 (N_6124,N_5905,N_5830);
nand U6125 (N_6125,N_5795,N_5776);
or U6126 (N_6126,N_5919,N_5808);
or U6127 (N_6127,N_5900,N_5802);
xor U6128 (N_6128,N_5753,N_5907);
or U6129 (N_6129,N_5757,N_5950);
or U6130 (N_6130,N_5837,N_5980);
nand U6131 (N_6131,N_5833,N_5997);
and U6132 (N_6132,N_5879,N_5903);
nand U6133 (N_6133,N_5938,N_5785);
nor U6134 (N_6134,N_5870,N_5841);
nand U6135 (N_6135,N_5828,N_5868);
or U6136 (N_6136,N_5888,N_5727);
xor U6137 (N_6137,N_5708,N_5763);
and U6138 (N_6138,N_5815,N_5741);
and U6139 (N_6139,N_5912,N_5946);
nand U6140 (N_6140,N_5847,N_5731);
xnor U6141 (N_6141,N_5835,N_5777);
nand U6142 (N_6142,N_5820,N_5976);
or U6143 (N_6143,N_5956,N_5773);
and U6144 (N_6144,N_5840,N_5822);
nor U6145 (N_6145,N_5797,N_5918);
and U6146 (N_6146,N_5964,N_5885);
or U6147 (N_6147,N_5730,N_5759);
xor U6148 (N_6148,N_5890,N_5930);
xnor U6149 (N_6149,N_5865,N_5821);
nor U6150 (N_6150,N_5706,N_5904);
and U6151 (N_6151,N_5997,N_5868);
or U6152 (N_6152,N_5708,N_5867);
nand U6153 (N_6153,N_5916,N_5841);
nor U6154 (N_6154,N_5829,N_5824);
xor U6155 (N_6155,N_5727,N_5879);
xor U6156 (N_6156,N_5806,N_5901);
nand U6157 (N_6157,N_5851,N_5745);
xor U6158 (N_6158,N_5855,N_5831);
or U6159 (N_6159,N_5945,N_5840);
xnor U6160 (N_6160,N_5703,N_5733);
nor U6161 (N_6161,N_5909,N_5891);
and U6162 (N_6162,N_5735,N_5757);
nor U6163 (N_6163,N_5730,N_5807);
and U6164 (N_6164,N_5806,N_5823);
or U6165 (N_6165,N_5862,N_5751);
or U6166 (N_6166,N_5828,N_5937);
nand U6167 (N_6167,N_5957,N_5871);
or U6168 (N_6168,N_5726,N_5813);
nor U6169 (N_6169,N_5965,N_5918);
nand U6170 (N_6170,N_5795,N_5950);
and U6171 (N_6171,N_5856,N_5939);
nor U6172 (N_6172,N_5831,N_5897);
or U6173 (N_6173,N_5717,N_5954);
and U6174 (N_6174,N_5822,N_5984);
and U6175 (N_6175,N_5992,N_5989);
or U6176 (N_6176,N_5939,N_5971);
or U6177 (N_6177,N_5814,N_5704);
nor U6178 (N_6178,N_5897,N_5906);
and U6179 (N_6179,N_5912,N_5847);
and U6180 (N_6180,N_5972,N_5724);
xor U6181 (N_6181,N_5822,N_5974);
nor U6182 (N_6182,N_5720,N_5998);
or U6183 (N_6183,N_5842,N_5705);
xnor U6184 (N_6184,N_5929,N_5752);
and U6185 (N_6185,N_5829,N_5791);
xor U6186 (N_6186,N_5752,N_5772);
and U6187 (N_6187,N_5921,N_5871);
nor U6188 (N_6188,N_5849,N_5930);
and U6189 (N_6189,N_5864,N_5927);
xor U6190 (N_6190,N_5919,N_5918);
nand U6191 (N_6191,N_5961,N_5952);
and U6192 (N_6192,N_5798,N_5886);
nor U6193 (N_6193,N_5753,N_5921);
xor U6194 (N_6194,N_5787,N_5749);
nand U6195 (N_6195,N_5836,N_5919);
nand U6196 (N_6196,N_5753,N_5821);
or U6197 (N_6197,N_5948,N_5710);
nor U6198 (N_6198,N_5891,N_5937);
nand U6199 (N_6199,N_5810,N_5776);
or U6200 (N_6200,N_5716,N_5865);
or U6201 (N_6201,N_5929,N_5796);
and U6202 (N_6202,N_5962,N_5920);
xor U6203 (N_6203,N_5984,N_5909);
and U6204 (N_6204,N_5751,N_5718);
or U6205 (N_6205,N_5872,N_5910);
or U6206 (N_6206,N_5799,N_5957);
and U6207 (N_6207,N_5731,N_5841);
nor U6208 (N_6208,N_5914,N_5925);
nand U6209 (N_6209,N_5808,N_5755);
or U6210 (N_6210,N_5734,N_5823);
or U6211 (N_6211,N_5745,N_5814);
and U6212 (N_6212,N_5998,N_5941);
or U6213 (N_6213,N_5802,N_5906);
nor U6214 (N_6214,N_5873,N_5927);
xnor U6215 (N_6215,N_5738,N_5933);
nor U6216 (N_6216,N_5951,N_5842);
or U6217 (N_6217,N_5717,N_5879);
xor U6218 (N_6218,N_5790,N_5879);
or U6219 (N_6219,N_5958,N_5772);
or U6220 (N_6220,N_5755,N_5740);
nand U6221 (N_6221,N_5982,N_5848);
nand U6222 (N_6222,N_5982,N_5935);
nor U6223 (N_6223,N_5795,N_5839);
nor U6224 (N_6224,N_5748,N_5967);
and U6225 (N_6225,N_5879,N_5827);
and U6226 (N_6226,N_5955,N_5707);
and U6227 (N_6227,N_5773,N_5809);
nor U6228 (N_6228,N_5921,N_5851);
and U6229 (N_6229,N_5758,N_5776);
xnor U6230 (N_6230,N_5854,N_5781);
nand U6231 (N_6231,N_5852,N_5976);
nand U6232 (N_6232,N_5942,N_5858);
nand U6233 (N_6233,N_5859,N_5800);
nand U6234 (N_6234,N_5917,N_5747);
or U6235 (N_6235,N_5945,N_5908);
and U6236 (N_6236,N_5989,N_5823);
nand U6237 (N_6237,N_5953,N_5948);
or U6238 (N_6238,N_5865,N_5802);
xor U6239 (N_6239,N_5703,N_5979);
nor U6240 (N_6240,N_5822,N_5989);
nor U6241 (N_6241,N_5902,N_5927);
xor U6242 (N_6242,N_5714,N_5707);
nand U6243 (N_6243,N_5863,N_5954);
or U6244 (N_6244,N_5838,N_5704);
or U6245 (N_6245,N_5922,N_5990);
or U6246 (N_6246,N_5883,N_5917);
xnor U6247 (N_6247,N_5706,N_5929);
nand U6248 (N_6248,N_5907,N_5947);
or U6249 (N_6249,N_5947,N_5727);
or U6250 (N_6250,N_5927,N_5826);
or U6251 (N_6251,N_5994,N_5805);
xnor U6252 (N_6252,N_5874,N_5740);
and U6253 (N_6253,N_5785,N_5948);
xor U6254 (N_6254,N_5811,N_5816);
nand U6255 (N_6255,N_5771,N_5967);
and U6256 (N_6256,N_5896,N_5845);
nor U6257 (N_6257,N_5796,N_5989);
and U6258 (N_6258,N_5822,N_5711);
xor U6259 (N_6259,N_5848,N_5725);
nand U6260 (N_6260,N_5851,N_5777);
or U6261 (N_6261,N_5866,N_5871);
xor U6262 (N_6262,N_5903,N_5856);
nand U6263 (N_6263,N_5850,N_5951);
nor U6264 (N_6264,N_5802,N_5763);
nand U6265 (N_6265,N_5796,N_5931);
xnor U6266 (N_6266,N_5721,N_5936);
or U6267 (N_6267,N_5777,N_5950);
nor U6268 (N_6268,N_5979,N_5947);
or U6269 (N_6269,N_5737,N_5861);
nor U6270 (N_6270,N_5846,N_5784);
nand U6271 (N_6271,N_5762,N_5718);
nand U6272 (N_6272,N_5958,N_5974);
xor U6273 (N_6273,N_5909,N_5865);
xor U6274 (N_6274,N_5944,N_5907);
xor U6275 (N_6275,N_5938,N_5988);
xnor U6276 (N_6276,N_5775,N_5846);
xnor U6277 (N_6277,N_5915,N_5760);
nand U6278 (N_6278,N_5987,N_5908);
xnor U6279 (N_6279,N_5873,N_5923);
or U6280 (N_6280,N_5906,N_5742);
nor U6281 (N_6281,N_5959,N_5833);
xnor U6282 (N_6282,N_5985,N_5721);
nor U6283 (N_6283,N_5814,N_5758);
or U6284 (N_6284,N_5728,N_5847);
nand U6285 (N_6285,N_5734,N_5875);
or U6286 (N_6286,N_5888,N_5932);
or U6287 (N_6287,N_5768,N_5989);
nor U6288 (N_6288,N_5881,N_5965);
nor U6289 (N_6289,N_5712,N_5860);
nand U6290 (N_6290,N_5757,N_5811);
or U6291 (N_6291,N_5783,N_5797);
and U6292 (N_6292,N_5750,N_5830);
nand U6293 (N_6293,N_5930,N_5945);
nor U6294 (N_6294,N_5945,N_5926);
nand U6295 (N_6295,N_5821,N_5893);
nor U6296 (N_6296,N_5789,N_5942);
xor U6297 (N_6297,N_5908,N_5914);
xnor U6298 (N_6298,N_5927,N_5867);
xor U6299 (N_6299,N_5773,N_5962);
nor U6300 (N_6300,N_6060,N_6279);
and U6301 (N_6301,N_6246,N_6023);
or U6302 (N_6302,N_6163,N_6162);
and U6303 (N_6303,N_6137,N_6084);
nor U6304 (N_6304,N_6250,N_6286);
nand U6305 (N_6305,N_6016,N_6225);
or U6306 (N_6306,N_6236,N_6025);
and U6307 (N_6307,N_6121,N_6287);
and U6308 (N_6308,N_6181,N_6109);
or U6309 (N_6309,N_6035,N_6180);
nor U6310 (N_6310,N_6153,N_6045);
xor U6311 (N_6311,N_6059,N_6291);
or U6312 (N_6312,N_6071,N_6085);
and U6313 (N_6313,N_6299,N_6078);
nor U6314 (N_6314,N_6282,N_6005);
or U6315 (N_6315,N_6002,N_6147);
or U6316 (N_6316,N_6042,N_6126);
or U6317 (N_6317,N_6273,N_6129);
xor U6318 (N_6318,N_6221,N_6292);
nand U6319 (N_6319,N_6019,N_6092);
xnor U6320 (N_6320,N_6211,N_6197);
xor U6321 (N_6321,N_6097,N_6011);
and U6322 (N_6322,N_6034,N_6185);
nand U6323 (N_6323,N_6231,N_6081);
xnor U6324 (N_6324,N_6079,N_6058);
xnor U6325 (N_6325,N_6262,N_6048);
or U6326 (N_6326,N_6252,N_6099);
and U6327 (N_6327,N_6064,N_6201);
or U6328 (N_6328,N_6222,N_6149);
xor U6329 (N_6329,N_6191,N_6183);
and U6330 (N_6330,N_6098,N_6090);
and U6331 (N_6331,N_6242,N_6251);
xor U6332 (N_6332,N_6119,N_6104);
and U6333 (N_6333,N_6170,N_6224);
xnor U6334 (N_6334,N_6103,N_6229);
nand U6335 (N_6335,N_6138,N_6200);
nor U6336 (N_6336,N_6074,N_6232);
or U6337 (N_6337,N_6220,N_6261);
nand U6338 (N_6338,N_6050,N_6125);
and U6339 (N_6339,N_6018,N_6265);
or U6340 (N_6340,N_6174,N_6227);
nand U6341 (N_6341,N_6187,N_6043);
nand U6342 (N_6342,N_6159,N_6274);
or U6343 (N_6343,N_6013,N_6101);
or U6344 (N_6344,N_6055,N_6118);
xor U6345 (N_6345,N_6190,N_6175);
or U6346 (N_6346,N_6038,N_6021);
or U6347 (N_6347,N_6066,N_6110);
nor U6348 (N_6348,N_6116,N_6017);
nand U6349 (N_6349,N_6269,N_6131);
xnor U6350 (N_6350,N_6245,N_6128);
xor U6351 (N_6351,N_6293,N_6241);
and U6352 (N_6352,N_6268,N_6167);
or U6353 (N_6353,N_6207,N_6015);
and U6354 (N_6354,N_6150,N_6049);
and U6355 (N_6355,N_6182,N_6053);
nor U6356 (N_6356,N_6248,N_6196);
and U6357 (N_6357,N_6144,N_6106);
nand U6358 (N_6358,N_6230,N_6156);
nor U6359 (N_6359,N_6117,N_6155);
nand U6360 (N_6360,N_6012,N_6255);
nor U6361 (N_6361,N_6148,N_6193);
and U6362 (N_6362,N_6283,N_6047);
nor U6363 (N_6363,N_6031,N_6171);
nand U6364 (N_6364,N_6056,N_6069);
and U6365 (N_6365,N_6022,N_6195);
xor U6366 (N_6366,N_6254,N_6000);
and U6367 (N_6367,N_6146,N_6247);
or U6368 (N_6368,N_6238,N_6253);
or U6369 (N_6369,N_6178,N_6290);
and U6370 (N_6370,N_6223,N_6205);
nand U6371 (N_6371,N_6094,N_6285);
and U6372 (N_6372,N_6214,N_6107);
and U6373 (N_6373,N_6233,N_6204);
nand U6374 (N_6374,N_6249,N_6213);
xnor U6375 (N_6375,N_6086,N_6028);
or U6376 (N_6376,N_6095,N_6206);
or U6377 (N_6377,N_6296,N_6029);
nor U6378 (N_6378,N_6141,N_6271);
and U6379 (N_6379,N_6258,N_6257);
nand U6380 (N_6380,N_6007,N_6041);
and U6381 (N_6381,N_6052,N_6142);
xnor U6382 (N_6382,N_6105,N_6177);
and U6383 (N_6383,N_6152,N_6073);
nand U6384 (N_6384,N_6004,N_6260);
and U6385 (N_6385,N_6140,N_6063);
nor U6386 (N_6386,N_6014,N_6001);
and U6387 (N_6387,N_6003,N_6054);
nor U6388 (N_6388,N_6199,N_6244);
nor U6389 (N_6389,N_6218,N_6184);
or U6390 (N_6390,N_6009,N_6024);
nand U6391 (N_6391,N_6087,N_6194);
nor U6392 (N_6392,N_6033,N_6186);
nor U6393 (N_6393,N_6068,N_6172);
or U6394 (N_6394,N_6032,N_6091);
nand U6395 (N_6395,N_6270,N_6202);
or U6396 (N_6396,N_6093,N_6100);
xnor U6397 (N_6397,N_6208,N_6114);
or U6398 (N_6398,N_6169,N_6295);
or U6399 (N_6399,N_6123,N_6212);
or U6400 (N_6400,N_6188,N_6217);
nor U6401 (N_6401,N_6006,N_6145);
xnor U6402 (N_6402,N_6240,N_6278);
or U6403 (N_6403,N_6189,N_6272);
nor U6404 (N_6404,N_6158,N_6151);
xor U6405 (N_6405,N_6266,N_6275);
or U6406 (N_6406,N_6256,N_6143);
and U6407 (N_6407,N_6239,N_6083);
nand U6408 (N_6408,N_6192,N_6122);
xor U6409 (N_6409,N_6040,N_6124);
nor U6410 (N_6410,N_6044,N_6164);
nand U6411 (N_6411,N_6027,N_6088);
nand U6412 (N_6412,N_6203,N_6267);
xor U6413 (N_6413,N_6165,N_6120);
nor U6414 (N_6414,N_6263,N_6235);
or U6415 (N_6415,N_6135,N_6133);
nand U6416 (N_6416,N_6030,N_6219);
nor U6417 (N_6417,N_6132,N_6161);
and U6418 (N_6418,N_6288,N_6072);
nor U6419 (N_6419,N_6062,N_6096);
nand U6420 (N_6420,N_6080,N_6008);
or U6421 (N_6421,N_6115,N_6127);
nor U6422 (N_6422,N_6067,N_6168);
nor U6423 (N_6423,N_6198,N_6234);
xor U6424 (N_6424,N_6076,N_6026);
nand U6425 (N_6425,N_6036,N_6130);
or U6426 (N_6426,N_6089,N_6037);
nand U6427 (N_6427,N_6046,N_6276);
nand U6428 (N_6428,N_6077,N_6173);
and U6429 (N_6429,N_6277,N_6134);
nand U6430 (N_6430,N_6082,N_6020);
nor U6431 (N_6431,N_6226,N_6209);
nor U6432 (N_6432,N_6108,N_6113);
and U6433 (N_6433,N_6157,N_6111);
nand U6434 (N_6434,N_6243,N_6264);
nand U6435 (N_6435,N_6228,N_6281);
nor U6436 (N_6436,N_6057,N_6065);
nand U6437 (N_6437,N_6284,N_6179);
nor U6438 (N_6438,N_6039,N_6176);
xnor U6439 (N_6439,N_6294,N_6154);
nand U6440 (N_6440,N_6010,N_6259);
nor U6441 (N_6441,N_6237,N_6075);
nand U6442 (N_6442,N_6061,N_6216);
nand U6443 (N_6443,N_6298,N_6102);
nor U6444 (N_6444,N_6160,N_6280);
nand U6445 (N_6445,N_6210,N_6215);
nor U6446 (N_6446,N_6289,N_6112);
nand U6447 (N_6447,N_6297,N_6136);
nor U6448 (N_6448,N_6051,N_6166);
or U6449 (N_6449,N_6070,N_6139);
or U6450 (N_6450,N_6212,N_6291);
nor U6451 (N_6451,N_6241,N_6025);
and U6452 (N_6452,N_6242,N_6079);
xnor U6453 (N_6453,N_6093,N_6081);
or U6454 (N_6454,N_6187,N_6101);
or U6455 (N_6455,N_6200,N_6088);
nand U6456 (N_6456,N_6291,N_6027);
and U6457 (N_6457,N_6101,N_6070);
or U6458 (N_6458,N_6039,N_6283);
xor U6459 (N_6459,N_6034,N_6179);
or U6460 (N_6460,N_6149,N_6217);
nor U6461 (N_6461,N_6025,N_6129);
xor U6462 (N_6462,N_6175,N_6284);
xnor U6463 (N_6463,N_6096,N_6131);
xor U6464 (N_6464,N_6175,N_6050);
or U6465 (N_6465,N_6052,N_6061);
nand U6466 (N_6466,N_6053,N_6086);
nor U6467 (N_6467,N_6226,N_6229);
nand U6468 (N_6468,N_6117,N_6228);
nor U6469 (N_6469,N_6208,N_6197);
nor U6470 (N_6470,N_6240,N_6177);
nor U6471 (N_6471,N_6155,N_6280);
and U6472 (N_6472,N_6129,N_6123);
xnor U6473 (N_6473,N_6274,N_6298);
nand U6474 (N_6474,N_6215,N_6162);
and U6475 (N_6475,N_6128,N_6253);
nor U6476 (N_6476,N_6224,N_6180);
or U6477 (N_6477,N_6096,N_6161);
and U6478 (N_6478,N_6251,N_6165);
xor U6479 (N_6479,N_6161,N_6140);
or U6480 (N_6480,N_6242,N_6269);
nor U6481 (N_6481,N_6191,N_6228);
and U6482 (N_6482,N_6243,N_6289);
and U6483 (N_6483,N_6001,N_6130);
or U6484 (N_6484,N_6281,N_6138);
or U6485 (N_6485,N_6142,N_6105);
and U6486 (N_6486,N_6122,N_6008);
xor U6487 (N_6487,N_6138,N_6003);
xnor U6488 (N_6488,N_6168,N_6007);
and U6489 (N_6489,N_6144,N_6200);
nand U6490 (N_6490,N_6257,N_6071);
xnor U6491 (N_6491,N_6007,N_6115);
nor U6492 (N_6492,N_6101,N_6150);
xnor U6493 (N_6493,N_6202,N_6104);
and U6494 (N_6494,N_6031,N_6121);
or U6495 (N_6495,N_6052,N_6287);
xor U6496 (N_6496,N_6139,N_6273);
nor U6497 (N_6497,N_6124,N_6194);
nor U6498 (N_6498,N_6164,N_6181);
nor U6499 (N_6499,N_6002,N_6009);
xor U6500 (N_6500,N_6217,N_6079);
and U6501 (N_6501,N_6171,N_6071);
nand U6502 (N_6502,N_6295,N_6222);
or U6503 (N_6503,N_6284,N_6272);
nor U6504 (N_6504,N_6019,N_6115);
nand U6505 (N_6505,N_6235,N_6012);
nor U6506 (N_6506,N_6235,N_6042);
nand U6507 (N_6507,N_6039,N_6207);
and U6508 (N_6508,N_6103,N_6140);
and U6509 (N_6509,N_6038,N_6241);
or U6510 (N_6510,N_6128,N_6110);
xor U6511 (N_6511,N_6277,N_6027);
nor U6512 (N_6512,N_6289,N_6275);
nand U6513 (N_6513,N_6022,N_6274);
nor U6514 (N_6514,N_6267,N_6076);
nor U6515 (N_6515,N_6249,N_6083);
or U6516 (N_6516,N_6180,N_6297);
nor U6517 (N_6517,N_6119,N_6102);
and U6518 (N_6518,N_6142,N_6256);
nand U6519 (N_6519,N_6221,N_6147);
nor U6520 (N_6520,N_6116,N_6069);
or U6521 (N_6521,N_6143,N_6119);
nor U6522 (N_6522,N_6271,N_6101);
nor U6523 (N_6523,N_6094,N_6242);
xnor U6524 (N_6524,N_6027,N_6082);
and U6525 (N_6525,N_6107,N_6166);
nand U6526 (N_6526,N_6186,N_6210);
nand U6527 (N_6527,N_6258,N_6073);
xor U6528 (N_6528,N_6082,N_6077);
nand U6529 (N_6529,N_6115,N_6148);
xor U6530 (N_6530,N_6128,N_6252);
nand U6531 (N_6531,N_6237,N_6070);
nand U6532 (N_6532,N_6111,N_6287);
or U6533 (N_6533,N_6074,N_6209);
or U6534 (N_6534,N_6161,N_6244);
nor U6535 (N_6535,N_6022,N_6014);
nor U6536 (N_6536,N_6131,N_6143);
or U6537 (N_6537,N_6160,N_6250);
nor U6538 (N_6538,N_6172,N_6011);
nand U6539 (N_6539,N_6063,N_6121);
xnor U6540 (N_6540,N_6025,N_6053);
or U6541 (N_6541,N_6111,N_6200);
and U6542 (N_6542,N_6079,N_6039);
nor U6543 (N_6543,N_6081,N_6045);
xnor U6544 (N_6544,N_6230,N_6119);
or U6545 (N_6545,N_6257,N_6206);
nand U6546 (N_6546,N_6068,N_6117);
and U6547 (N_6547,N_6189,N_6062);
nor U6548 (N_6548,N_6003,N_6057);
or U6549 (N_6549,N_6118,N_6250);
and U6550 (N_6550,N_6273,N_6240);
xnor U6551 (N_6551,N_6061,N_6037);
nor U6552 (N_6552,N_6052,N_6228);
xnor U6553 (N_6553,N_6100,N_6086);
or U6554 (N_6554,N_6238,N_6284);
or U6555 (N_6555,N_6096,N_6271);
nand U6556 (N_6556,N_6235,N_6044);
and U6557 (N_6557,N_6264,N_6194);
nand U6558 (N_6558,N_6085,N_6006);
xnor U6559 (N_6559,N_6292,N_6150);
nand U6560 (N_6560,N_6296,N_6120);
and U6561 (N_6561,N_6058,N_6291);
xnor U6562 (N_6562,N_6273,N_6002);
nor U6563 (N_6563,N_6057,N_6043);
or U6564 (N_6564,N_6161,N_6257);
nand U6565 (N_6565,N_6049,N_6011);
nand U6566 (N_6566,N_6136,N_6095);
or U6567 (N_6567,N_6152,N_6238);
and U6568 (N_6568,N_6244,N_6073);
nand U6569 (N_6569,N_6023,N_6226);
and U6570 (N_6570,N_6127,N_6231);
or U6571 (N_6571,N_6106,N_6160);
xnor U6572 (N_6572,N_6204,N_6299);
and U6573 (N_6573,N_6059,N_6047);
xor U6574 (N_6574,N_6145,N_6070);
or U6575 (N_6575,N_6284,N_6170);
or U6576 (N_6576,N_6026,N_6245);
and U6577 (N_6577,N_6286,N_6189);
xor U6578 (N_6578,N_6146,N_6232);
nand U6579 (N_6579,N_6035,N_6002);
nor U6580 (N_6580,N_6114,N_6071);
and U6581 (N_6581,N_6025,N_6251);
nor U6582 (N_6582,N_6159,N_6035);
or U6583 (N_6583,N_6166,N_6159);
and U6584 (N_6584,N_6102,N_6137);
and U6585 (N_6585,N_6026,N_6251);
or U6586 (N_6586,N_6196,N_6238);
xor U6587 (N_6587,N_6178,N_6128);
and U6588 (N_6588,N_6131,N_6024);
and U6589 (N_6589,N_6184,N_6254);
nor U6590 (N_6590,N_6118,N_6117);
and U6591 (N_6591,N_6266,N_6170);
xnor U6592 (N_6592,N_6290,N_6286);
and U6593 (N_6593,N_6164,N_6270);
nand U6594 (N_6594,N_6240,N_6014);
nor U6595 (N_6595,N_6082,N_6210);
nor U6596 (N_6596,N_6111,N_6064);
nor U6597 (N_6597,N_6176,N_6232);
and U6598 (N_6598,N_6085,N_6060);
nand U6599 (N_6599,N_6005,N_6103);
and U6600 (N_6600,N_6540,N_6521);
or U6601 (N_6601,N_6442,N_6548);
or U6602 (N_6602,N_6500,N_6302);
nor U6603 (N_6603,N_6400,N_6370);
nor U6604 (N_6604,N_6588,N_6534);
and U6605 (N_6605,N_6563,N_6492);
and U6606 (N_6606,N_6360,N_6533);
nor U6607 (N_6607,N_6408,N_6300);
xor U6608 (N_6608,N_6590,N_6560);
xor U6609 (N_6609,N_6386,N_6527);
or U6610 (N_6610,N_6425,N_6474);
xnor U6611 (N_6611,N_6456,N_6536);
nor U6612 (N_6612,N_6512,N_6564);
nand U6613 (N_6613,N_6486,N_6438);
nand U6614 (N_6614,N_6448,N_6593);
and U6615 (N_6615,N_6517,N_6362);
and U6616 (N_6616,N_6332,N_6365);
or U6617 (N_6617,N_6543,N_6428);
and U6618 (N_6618,N_6509,N_6364);
nand U6619 (N_6619,N_6567,N_6353);
nor U6620 (N_6620,N_6510,N_6462);
or U6621 (N_6621,N_6508,N_6505);
and U6622 (N_6622,N_6317,N_6447);
nand U6623 (N_6623,N_6496,N_6460);
xor U6624 (N_6624,N_6398,N_6561);
or U6625 (N_6625,N_6596,N_6318);
and U6626 (N_6626,N_6587,N_6552);
nand U6627 (N_6627,N_6379,N_6541);
nand U6628 (N_6628,N_6330,N_6491);
or U6629 (N_6629,N_6396,N_6357);
or U6630 (N_6630,N_6352,N_6413);
nor U6631 (N_6631,N_6566,N_6581);
nor U6632 (N_6632,N_6539,N_6390);
xor U6633 (N_6633,N_6380,N_6483);
nand U6634 (N_6634,N_6369,N_6554);
nand U6635 (N_6635,N_6526,N_6482);
nor U6636 (N_6636,N_6472,N_6407);
and U6637 (N_6637,N_6446,N_6591);
nor U6638 (N_6638,N_6454,N_6328);
and U6639 (N_6639,N_6504,N_6417);
and U6640 (N_6640,N_6549,N_6394);
and U6641 (N_6641,N_6439,N_6444);
xnor U6642 (N_6642,N_6363,N_6316);
or U6643 (N_6643,N_6367,N_6524);
xnor U6644 (N_6644,N_6368,N_6572);
and U6645 (N_6645,N_6599,N_6575);
nand U6646 (N_6646,N_6341,N_6349);
nor U6647 (N_6647,N_6597,N_6348);
xor U6648 (N_6648,N_6434,N_6303);
or U6649 (N_6649,N_6494,N_6433);
nand U6650 (N_6650,N_6470,N_6385);
nand U6651 (N_6651,N_6405,N_6412);
nand U6652 (N_6652,N_6522,N_6319);
and U6653 (N_6653,N_6399,N_6595);
nor U6654 (N_6654,N_6573,N_6419);
nand U6655 (N_6655,N_6322,N_6424);
and U6656 (N_6656,N_6535,N_6347);
nor U6657 (N_6657,N_6545,N_6479);
and U6658 (N_6658,N_6329,N_6406);
xor U6659 (N_6659,N_6311,N_6476);
or U6660 (N_6660,N_6324,N_6471);
nor U6661 (N_6661,N_6475,N_6337);
nand U6662 (N_6662,N_6562,N_6520);
or U6663 (N_6663,N_6464,N_6592);
nand U6664 (N_6664,N_6459,N_6503);
nand U6665 (N_6665,N_6309,N_6409);
or U6666 (N_6666,N_6578,N_6421);
and U6667 (N_6667,N_6410,N_6542);
and U6668 (N_6668,N_6507,N_6391);
and U6669 (N_6669,N_6484,N_6555);
and U6670 (N_6670,N_6559,N_6516);
xor U6671 (N_6671,N_6571,N_6314);
nand U6672 (N_6672,N_6450,N_6418);
xor U6673 (N_6673,N_6529,N_6528);
nand U6674 (N_6674,N_6457,N_6315);
and U6675 (N_6675,N_6377,N_6344);
nor U6676 (N_6676,N_6495,N_6339);
nand U6677 (N_6677,N_6537,N_6493);
or U6678 (N_6678,N_6467,N_6589);
and U6679 (N_6679,N_6307,N_6313);
nor U6680 (N_6680,N_6432,N_6582);
and U6681 (N_6681,N_6401,N_6415);
xor U6682 (N_6682,N_6420,N_6381);
nor U6683 (N_6683,N_6331,N_6308);
xnor U6684 (N_6684,N_6373,N_6389);
nand U6685 (N_6685,N_6498,N_6463);
or U6686 (N_6686,N_6305,N_6392);
nand U6687 (N_6687,N_6465,N_6411);
xnor U6688 (N_6688,N_6336,N_6469);
xnor U6689 (N_6689,N_6550,N_6519);
xnor U6690 (N_6690,N_6372,N_6487);
and U6691 (N_6691,N_6544,N_6530);
nor U6692 (N_6692,N_6441,N_6445);
nor U6693 (N_6693,N_6383,N_6477);
nor U6694 (N_6694,N_6436,N_6455);
nor U6695 (N_6695,N_6565,N_6466);
nand U6696 (N_6696,N_6375,N_6378);
nand U6697 (N_6697,N_6478,N_6402);
nand U6698 (N_6698,N_6449,N_6580);
or U6699 (N_6699,N_6335,N_6320);
nand U6700 (N_6700,N_6574,N_6414);
and U6701 (N_6701,N_6387,N_6452);
and U6702 (N_6702,N_6518,N_6359);
xor U6703 (N_6703,N_6501,N_6423);
xor U6704 (N_6704,N_6356,N_6358);
or U6705 (N_6705,N_6404,N_6310);
or U6706 (N_6706,N_6513,N_6345);
xor U6707 (N_6707,N_6384,N_6440);
nor U6708 (N_6708,N_6426,N_6570);
and U6709 (N_6709,N_6304,N_6583);
or U6710 (N_6710,N_6497,N_6351);
nand U6711 (N_6711,N_6395,N_6422);
nand U6712 (N_6712,N_6325,N_6355);
xnor U6713 (N_6713,N_6350,N_6547);
xnor U6714 (N_6714,N_6342,N_6435);
nor U6715 (N_6715,N_6321,N_6382);
nand U6716 (N_6716,N_6343,N_6557);
nor U6717 (N_6717,N_6584,N_6416);
or U6718 (N_6718,N_6468,N_6511);
or U6719 (N_6719,N_6458,N_6338);
nand U6720 (N_6720,N_6576,N_6346);
nor U6721 (N_6721,N_6393,N_6451);
or U6722 (N_6722,N_6514,N_6481);
and U6723 (N_6723,N_6388,N_6598);
nor U6724 (N_6724,N_6553,N_6532);
nand U6725 (N_6725,N_6354,N_6531);
nor U6726 (N_6726,N_6376,N_6431);
xnor U6727 (N_6727,N_6327,N_6443);
or U6728 (N_6728,N_6579,N_6334);
xnor U6729 (N_6729,N_6594,N_6333);
nor U6730 (N_6730,N_6371,N_6546);
xor U6731 (N_6731,N_6556,N_6374);
xnor U6732 (N_6732,N_6506,N_6585);
nand U6733 (N_6733,N_6502,N_6306);
nand U6734 (N_6734,N_6403,N_6499);
nor U6735 (N_6735,N_6490,N_6301);
and U6736 (N_6736,N_6429,N_6586);
or U6737 (N_6737,N_6453,N_6568);
and U6738 (N_6738,N_6480,N_6323);
nor U6739 (N_6739,N_6427,N_6361);
xor U6740 (N_6740,N_6326,N_6366);
and U6741 (N_6741,N_6485,N_6312);
or U6742 (N_6742,N_6430,N_6569);
nor U6743 (N_6743,N_6340,N_6461);
and U6744 (N_6744,N_6488,N_6437);
and U6745 (N_6745,N_6551,N_6577);
or U6746 (N_6746,N_6523,N_6489);
and U6747 (N_6747,N_6558,N_6515);
nand U6748 (N_6748,N_6473,N_6397);
nor U6749 (N_6749,N_6538,N_6525);
xnor U6750 (N_6750,N_6329,N_6573);
and U6751 (N_6751,N_6357,N_6343);
nand U6752 (N_6752,N_6378,N_6558);
xnor U6753 (N_6753,N_6386,N_6480);
or U6754 (N_6754,N_6521,N_6587);
nor U6755 (N_6755,N_6560,N_6371);
and U6756 (N_6756,N_6422,N_6300);
xnor U6757 (N_6757,N_6518,N_6514);
xor U6758 (N_6758,N_6481,N_6394);
and U6759 (N_6759,N_6408,N_6570);
nand U6760 (N_6760,N_6578,N_6497);
and U6761 (N_6761,N_6423,N_6472);
xor U6762 (N_6762,N_6557,N_6303);
or U6763 (N_6763,N_6360,N_6408);
or U6764 (N_6764,N_6362,N_6533);
nor U6765 (N_6765,N_6438,N_6392);
nand U6766 (N_6766,N_6598,N_6336);
nor U6767 (N_6767,N_6394,N_6405);
nand U6768 (N_6768,N_6488,N_6369);
nor U6769 (N_6769,N_6349,N_6577);
xnor U6770 (N_6770,N_6362,N_6496);
or U6771 (N_6771,N_6494,N_6492);
and U6772 (N_6772,N_6372,N_6547);
and U6773 (N_6773,N_6343,N_6350);
nor U6774 (N_6774,N_6420,N_6581);
and U6775 (N_6775,N_6443,N_6428);
nand U6776 (N_6776,N_6471,N_6498);
nor U6777 (N_6777,N_6366,N_6492);
and U6778 (N_6778,N_6380,N_6401);
nand U6779 (N_6779,N_6506,N_6326);
or U6780 (N_6780,N_6493,N_6519);
xnor U6781 (N_6781,N_6521,N_6353);
or U6782 (N_6782,N_6408,N_6305);
or U6783 (N_6783,N_6406,N_6565);
nor U6784 (N_6784,N_6325,N_6451);
xnor U6785 (N_6785,N_6468,N_6374);
or U6786 (N_6786,N_6475,N_6372);
nor U6787 (N_6787,N_6363,N_6381);
xor U6788 (N_6788,N_6430,N_6347);
nor U6789 (N_6789,N_6457,N_6535);
nand U6790 (N_6790,N_6485,N_6364);
nor U6791 (N_6791,N_6541,N_6317);
nand U6792 (N_6792,N_6587,N_6442);
and U6793 (N_6793,N_6447,N_6356);
nor U6794 (N_6794,N_6324,N_6331);
nor U6795 (N_6795,N_6552,N_6570);
or U6796 (N_6796,N_6433,N_6463);
xnor U6797 (N_6797,N_6585,N_6432);
or U6798 (N_6798,N_6583,N_6474);
and U6799 (N_6799,N_6506,N_6385);
xor U6800 (N_6800,N_6569,N_6453);
nor U6801 (N_6801,N_6490,N_6322);
xor U6802 (N_6802,N_6437,N_6388);
xnor U6803 (N_6803,N_6547,N_6323);
and U6804 (N_6804,N_6595,N_6360);
or U6805 (N_6805,N_6371,N_6331);
nand U6806 (N_6806,N_6392,N_6449);
nand U6807 (N_6807,N_6508,N_6352);
or U6808 (N_6808,N_6511,N_6383);
nor U6809 (N_6809,N_6314,N_6456);
nor U6810 (N_6810,N_6325,N_6477);
nand U6811 (N_6811,N_6487,N_6488);
and U6812 (N_6812,N_6444,N_6351);
or U6813 (N_6813,N_6367,N_6420);
nor U6814 (N_6814,N_6409,N_6440);
or U6815 (N_6815,N_6427,N_6430);
nor U6816 (N_6816,N_6459,N_6517);
and U6817 (N_6817,N_6333,N_6379);
nand U6818 (N_6818,N_6549,N_6466);
nor U6819 (N_6819,N_6591,N_6346);
nor U6820 (N_6820,N_6356,N_6407);
or U6821 (N_6821,N_6331,N_6329);
and U6822 (N_6822,N_6333,N_6363);
nor U6823 (N_6823,N_6342,N_6381);
nand U6824 (N_6824,N_6582,N_6451);
xnor U6825 (N_6825,N_6517,N_6366);
nor U6826 (N_6826,N_6552,N_6538);
xor U6827 (N_6827,N_6334,N_6332);
nor U6828 (N_6828,N_6442,N_6388);
nand U6829 (N_6829,N_6448,N_6470);
and U6830 (N_6830,N_6450,N_6508);
or U6831 (N_6831,N_6387,N_6300);
and U6832 (N_6832,N_6397,N_6351);
nor U6833 (N_6833,N_6480,N_6341);
or U6834 (N_6834,N_6553,N_6442);
and U6835 (N_6835,N_6435,N_6410);
nand U6836 (N_6836,N_6518,N_6453);
xor U6837 (N_6837,N_6382,N_6318);
and U6838 (N_6838,N_6342,N_6405);
or U6839 (N_6839,N_6341,N_6472);
and U6840 (N_6840,N_6370,N_6340);
nor U6841 (N_6841,N_6311,N_6528);
nand U6842 (N_6842,N_6508,N_6317);
and U6843 (N_6843,N_6351,N_6452);
nand U6844 (N_6844,N_6450,N_6583);
and U6845 (N_6845,N_6458,N_6482);
nand U6846 (N_6846,N_6326,N_6361);
or U6847 (N_6847,N_6402,N_6452);
or U6848 (N_6848,N_6495,N_6458);
or U6849 (N_6849,N_6366,N_6393);
and U6850 (N_6850,N_6523,N_6300);
nor U6851 (N_6851,N_6539,N_6371);
xnor U6852 (N_6852,N_6431,N_6455);
and U6853 (N_6853,N_6594,N_6481);
xnor U6854 (N_6854,N_6403,N_6384);
and U6855 (N_6855,N_6403,N_6312);
and U6856 (N_6856,N_6417,N_6515);
nor U6857 (N_6857,N_6332,N_6305);
xnor U6858 (N_6858,N_6325,N_6535);
xor U6859 (N_6859,N_6514,N_6517);
xnor U6860 (N_6860,N_6546,N_6567);
and U6861 (N_6861,N_6503,N_6333);
or U6862 (N_6862,N_6583,N_6501);
or U6863 (N_6863,N_6498,N_6512);
and U6864 (N_6864,N_6523,N_6506);
nor U6865 (N_6865,N_6430,N_6584);
xor U6866 (N_6866,N_6537,N_6402);
and U6867 (N_6867,N_6533,N_6331);
and U6868 (N_6868,N_6406,N_6433);
nand U6869 (N_6869,N_6526,N_6317);
or U6870 (N_6870,N_6328,N_6393);
nand U6871 (N_6871,N_6560,N_6567);
and U6872 (N_6872,N_6434,N_6551);
or U6873 (N_6873,N_6379,N_6522);
and U6874 (N_6874,N_6477,N_6388);
xor U6875 (N_6875,N_6314,N_6378);
nor U6876 (N_6876,N_6490,N_6355);
xor U6877 (N_6877,N_6417,N_6438);
or U6878 (N_6878,N_6581,N_6453);
and U6879 (N_6879,N_6322,N_6370);
nand U6880 (N_6880,N_6422,N_6531);
or U6881 (N_6881,N_6445,N_6474);
nor U6882 (N_6882,N_6300,N_6472);
and U6883 (N_6883,N_6413,N_6363);
xor U6884 (N_6884,N_6516,N_6526);
nor U6885 (N_6885,N_6545,N_6372);
nor U6886 (N_6886,N_6315,N_6553);
xnor U6887 (N_6887,N_6410,N_6402);
nand U6888 (N_6888,N_6515,N_6380);
nor U6889 (N_6889,N_6320,N_6573);
or U6890 (N_6890,N_6386,N_6327);
xnor U6891 (N_6891,N_6366,N_6572);
nor U6892 (N_6892,N_6383,N_6348);
nor U6893 (N_6893,N_6321,N_6433);
nand U6894 (N_6894,N_6404,N_6424);
xor U6895 (N_6895,N_6327,N_6302);
nand U6896 (N_6896,N_6523,N_6483);
or U6897 (N_6897,N_6527,N_6309);
and U6898 (N_6898,N_6424,N_6332);
or U6899 (N_6899,N_6589,N_6355);
xnor U6900 (N_6900,N_6626,N_6852);
xor U6901 (N_6901,N_6841,N_6785);
nand U6902 (N_6902,N_6842,N_6862);
xor U6903 (N_6903,N_6748,N_6839);
or U6904 (N_6904,N_6877,N_6725);
nor U6905 (N_6905,N_6708,N_6791);
nand U6906 (N_6906,N_6605,N_6669);
nor U6907 (N_6907,N_6733,N_6884);
or U6908 (N_6908,N_6888,N_6667);
xnor U6909 (N_6909,N_6711,N_6606);
nor U6910 (N_6910,N_6730,N_6719);
xnor U6911 (N_6911,N_6738,N_6643);
nor U6912 (N_6912,N_6706,N_6808);
or U6913 (N_6913,N_6739,N_6767);
xnor U6914 (N_6914,N_6892,N_6766);
or U6915 (N_6915,N_6826,N_6714);
nor U6916 (N_6916,N_6620,N_6628);
and U6917 (N_6917,N_6624,N_6815);
nor U6918 (N_6918,N_6656,N_6891);
or U6919 (N_6919,N_6604,N_6866);
nor U6920 (N_6920,N_6801,N_6872);
nor U6921 (N_6921,N_6810,N_6698);
or U6922 (N_6922,N_6681,N_6752);
or U6923 (N_6923,N_6790,N_6787);
or U6924 (N_6924,N_6607,N_6797);
or U6925 (N_6925,N_6675,N_6881);
and U6926 (N_6926,N_6761,N_6819);
or U6927 (N_6927,N_6772,N_6799);
or U6928 (N_6928,N_6619,N_6736);
xor U6929 (N_6929,N_6735,N_6649);
nand U6930 (N_6930,N_6788,N_6869);
nand U6931 (N_6931,N_6774,N_6610);
xor U6932 (N_6932,N_6613,N_6696);
and U6933 (N_6933,N_6701,N_6700);
nor U6934 (N_6934,N_6794,N_6609);
nor U6935 (N_6935,N_6679,N_6685);
and U6936 (N_6936,N_6641,N_6899);
or U6937 (N_6937,N_6809,N_6779);
nand U6938 (N_6938,N_6849,N_6726);
xor U6939 (N_6939,N_6776,N_6786);
and U6940 (N_6940,N_6835,N_6837);
nor U6941 (N_6941,N_6759,N_6715);
nand U6942 (N_6942,N_6647,N_6769);
and U6943 (N_6943,N_6644,N_6713);
or U6944 (N_6944,N_6789,N_6847);
nor U6945 (N_6945,N_6630,N_6631);
or U6946 (N_6946,N_6792,N_6823);
or U6947 (N_6947,N_6770,N_6690);
xnor U6948 (N_6948,N_6645,N_6781);
xnor U6949 (N_6949,N_6886,N_6636);
nand U6950 (N_6950,N_6639,N_6804);
or U6951 (N_6951,N_6629,N_6845);
and U6952 (N_6952,N_6699,N_6694);
nor U6953 (N_6953,N_6895,N_6763);
xor U6954 (N_6954,N_6898,N_6820);
nand U6955 (N_6955,N_6734,N_6637);
and U6956 (N_6956,N_6704,N_6832);
xor U6957 (N_6957,N_6775,N_6650);
xor U6958 (N_6958,N_6834,N_6634);
nand U6959 (N_6959,N_6844,N_6831);
or U6960 (N_6960,N_6848,N_6855);
nand U6961 (N_6961,N_6851,N_6879);
and U6962 (N_6962,N_6753,N_6611);
nand U6963 (N_6963,N_6850,N_6732);
nor U6964 (N_6964,N_6646,N_6885);
nand U6965 (N_6965,N_6824,N_6671);
xnor U6966 (N_6966,N_6659,N_6840);
and U6967 (N_6967,N_6635,N_6758);
xnor U6968 (N_6968,N_6668,N_6653);
nand U6969 (N_6969,N_6652,N_6755);
nor U6970 (N_6970,N_6747,N_6800);
or U6971 (N_6971,N_6843,N_6859);
or U6972 (N_6972,N_6727,N_6601);
xnor U6973 (N_6973,N_6897,N_6618);
and U6974 (N_6974,N_6664,N_6817);
and U6975 (N_6975,N_6889,N_6853);
xor U6976 (N_6976,N_6724,N_6720);
or U6977 (N_6977,N_6833,N_6603);
xnor U6978 (N_6978,N_6682,N_6757);
or U6979 (N_6979,N_6751,N_6655);
nor U6980 (N_6980,N_6807,N_6865);
and U6981 (N_6981,N_6705,N_6802);
xnor U6982 (N_6982,N_6709,N_6878);
nand U6983 (N_6983,N_6838,N_6821);
or U6984 (N_6984,N_6689,N_6762);
xor U6985 (N_6985,N_6737,N_6796);
or U6986 (N_6986,N_6661,N_6854);
nand U6987 (N_6987,N_6818,N_6666);
nand U6988 (N_6988,N_6625,N_6693);
nor U6989 (N_6989,N_6870,N_6777);
or U6990 (N_6990,N_6780,N_6614);
xor U6991 (N_6991,N_6612,N_6658);
nor U6992 (N_6992,N_6712,N_6868);
nor U6993 (N_6993,N_6710,N_6765);
and U6994 (N_6994,N_6622,N_6608);
nand U6995 (N_6995,N_6729,N_6723);
xor U6996 (N_6996,N_6662,N_6836);
and U6997 (N_6997,N_6632,N_6616);
nor U6998 (N_6998,N_6672,N_6741);
nand U6999 (N_6999,N_6858,N_6602);
nor U7000 (N_7000,N_6740,N_6684);
xnor U7001 (N_7001,N_6871,N_6697);
or U7002 (N_7002,N_6688,N_6703);
or U7003 (N_7003,N_6722,N_6692);
nand U7004 (N_7004,N_6673,N_6728);
xor U7005 (N_7005,N_6882,N_6812);
nand U7006 (N_7006,N_6875,N_6687);
nand U7007 (N_7007,N_6642,N_6873);
and U7008 (N_7008,N_6717,N_6864);
and U7009 (N_7009,N_6768,N_6860);
xor U7010 (N_7010,N_6887,N_6670);
nor U7011 (N_7011,N_6816,N_6827);
or U7012 (N_7012,N_6657,N_6627);
or U7013 (N_7013,N_6795,N_6750);
and U7014 (N_7014,N_6749,N_6783);
and U7015 (N_7015,N_6707,N_6651);
xor U7016 (N_7016,N_6867,N_6876);
xnor U7017 (N_7017,N_6745,N_6773);
nand U7018 (N_7018,N_6678,N_6640);
nand U7019 (N_7019,N_6756,N_6894);
nand U7020 (N_7020,N_6617,N_6830);
nor U7021 (N_7021,N_6805,N_6822);
or U7022 (N_7022,N_6683,N_6615);
nor U7023 (N_7023,N_6846,N_6742);
and U7024 (N_7024,N_6746,N_6893);
nand U7025 (N_7025,N_6676,N_6803);
or U7026 (N_7026,N_6686,N_6674);
or U7027 (N_7027,N_6764,N_6806);
xor U7028 (N_7028,N_6691,N_6754);
nor U7029 (N_7029,N_6880,N_6828);
or U7030 (N_7030,N_6744,N_6883);
or U7031 (N_7031,N_6731,N_6648);
nand U7032 (N_7032,N_6890,N_6861);
or U7033 (N_7033,N_6813,N_6825);
nand U7034 (N_7034,N_6660,N_6654);
xor U7035 (N_7035,N_6829,N_6623);
or U7036 (N_7036,N_6856,N_6782);
nand U7037 (N_7037,N_6857,N_6874);
nor U7038 (N_7038,N_6896,N_6716);
and U7039 (N_7039,N_6600,N_6784);
and U7040 (N_7040,N_6695,N_6863);
xnor U7041 (N_7041,N_6680,N_6798);
or U7042 (N_7042,N_6760,N_6814);
or U7043 (N_7043,N_6811,N_6771);
nand U7044 (N_7044,N_6721,N_6793);
nor U7045 (N_7045,N_6638,N_6677);
nor U7046 (N_7046,N_6621,N_6718);
or U7047 (N_7047,N_6663,N_6633);
nand U7048 (N_7048,N_6702,N_6665);
nor U7049 (N_7049,N_6778,N_6743);
or U7050 (N_7050,N_6855,N_6772);
xnor U7051 (N_7051,N_6780,N_6838);
or U7052 (N_7052,N_6800,N_6614);
or U7053 (N_7053,N_6832,N_6856);
xnor U7054 (N_7054,N_6896,N_6655);
nor U7055 (N_7055,N_6615,N_6612);
nand U7056 (N_7056,N_6899,N_6658);
xnor U7057 (N_7057,N_6655,N_6891);
nor U7058 (N_7058,N_6749,N_6853);
and U7059 (N_7059,N_6716,N_6869);
and U7060 (N_7060,N_6718,N_6720);
nor U7061 (N_7061,N_6636,N_6723);
nor U7062 (N_7062,N_6651,N_6850);
nor U7063 (N_7063,N_6890,N_6722);
nand U7064 (N_7064,N_6893,N_6881);
and U7065 (N_7065,N_6777,N_6646);
and U7066 (N_7066,N_6674,N_6895);
and U7067 (N_7067,N_6821,N_6846);
or U7068 (N_7068,N_6768,N_6792);
nand U7069 (N_7069,N_6817,N_6873);
nand U7070 (N_7070,N_6617,N_6612);
nand U7071 (N_7071,N_6851,N_6746);
or U7072 (N_7072,N_6645,N_6715);
nor U7073 (N_7073,N_6762,N_6776);
and U7074 (N_7074,N_6600,N_6830);
nor U7075 (N_7075,N_6652,N_6649);
and U7076 (N_7076,N_6805,N_6768);
nand U7077 (N_7077,N_6611,N_6663);
nand U7078 (N_7078,N_6737,N_6668);
xnor U7079 (N_7079,N_6683,N_6890);
nand U7080 (N_7080,N_6602,N_6801);
nand U7081 (N_7081,N_6765,N_6884);
and U7082 (N_7082,N_6896,N_6891);
xnor U7083 (N_7083,N_6763,N_6679);
nand U7084 (N_7084,N_6715,N_6780);
nand U7085 (N_7085,N_6659,N_6730);
or U7086 (N_7086,N_6671,N_6879);
and U7087 (N_7087,N_6636,N_6708);
xnor U7088 (N_7088,N_6741,N_6870);
or U7089 (N_7089,N_6883,N_6775);
or U7090 (N_7090,N_6795,N_6736);
and U7091 (N_7091,N_6713,N_6724);
and U7092 (N_7092,N_6707,N_6899);
xnor U7093 (N_7093,N_6809,N_6849);
xor U7094 (N_7094,N_6607,N_6863);
or U7095 (N_7095,N_6702,N_6618);
xor U7096 (N_7096,N_6884,N_6620);
or U7097 (N_7097,N_6648,N_6723);
and U7098 (N_7098,N_6662,N_6737);
nor U7099 (N_7099,N_6782,N_6867);
nand U7100 (N_7100,N_6775,N_6888);
nand U7101 (N_7101,N_6699,N_6864);
and U7102 (N_7102,N_6864,N_6747);
xor U7103 (N_7103,N_6633,N_6893);
or U7104 (N_7104,N_6616,N_6876);
and U7105 (N_7105,N_6670,N_6683);
nor U7106 (N_7106,N_6713,N_6647);
or U7107 (N_7107,N_6733,N_6720);
or U7108 (N_7108,N_6769,N_6704);
xor U7109 (N_7109,N_6611,N_6778);
xor U7110 (N_7110,N_6676,N_6846);
nand U7111 (N_7111,N_6726,N_6690);
or U7112 (N_7112,N_6607,N_6852);
nor U7113 (N_7113,N_6719,N_6832);
and U7114 (N_7114,N_6724,N_6853);
or U7115 (N_7115,N_6666,N_6798);
nand U7116 (N_7116,N_6673,N_6623);
and U7117 (N_7117,N_6799,N_6770);
xor U7118 (N_7118,N_6696,N_6704);
nor U7119 (N_7119,N_6672,N_6774);
or U7120 (N_7120,N_6678,N_6754);
and U7121 (N_7121,N_6856,N_6665);
nor U7122 (N_7122,N_6625,N_6836);
xnor U7123 (N_7123,N_6750,N_6866);
xor U7124 (N_7124,N_6634,N_6606);
nand U7125 (N_7125,N_6836,N_6892);
and U7126 (N_7126,N_6613,N_6852);
nor U7127 (N_7127,N_6822,N_6688);
and U7128 (N_7128,N_6873,N_6774);
or U7129 (N_7129,N_6666,N_6652);
nor U7130 (N_7130,N_6698,N_6821);
xnor U7131 (N_7131,N_6888,N_6855);
nor U7132 (N_7132,N_6690,N_6858);
and U7133 (N_7133,N_6730,N_6800);
nand U7134 (N_7134,N_6606,N_6625);
and U7135 (N_7135,N_6745,N_6881);
nor U7136 (N_7136,N_6733,N_6844);
xnor U7137 (N_7137,N_6889,N_6754);
or U7138 (N_7138,N_6691,N_6803);
xnor U7139 (N_7139,N_6789,N_6765);
and U7140 (N_7140,N_6812,N_6868);
and U7141 (N_7141,N_6774,N_6712);
and U7142 (N_7142,N_6723,N_6706);
xnor U7143 (N_7143,N_6779,N_6655);
nor U7144 (N_7144,N_6702,N_6663);
and U7145 (N_7145,N_6773,N_6643);
nor U7146 (N_7146,N_6716,N_6677);
nor U7147 (N_7147,N_6620,N_6664);
xor U7148 (N_7148,N_6896,N_6865);
xnor U7149 (N_7149,N_6783,N_6693);
or U7150 (N_7150,N_6752,N_6811);
or U7151 (N_7151,N_6713,N_6726);
or U7152 (N_7152,N_6635,N_6733);
nor U7153 (N_7153,N_6626,N_6683);
nor U7154 (N_7154,N_6668,N_6825);
nor U7155 (N_7155,N_6744,N_6843);
and U7156 (N_7156,N_6701,N_6698);
nor U7157 (N_7157,N_6835,N_6736);
xor U7158 (N_7158,N_6605,N_6673);
nor U7159 (N_7159,N_6680,N_6849);
nor U7160 (N_7160,N_6729,N_6819);
and U7161 (N_7161,N_6730,N_6752);
xnor U7162 (N_7162,N_6716,N_6714);
nand U7163 (N_7163,N_6824,N_6621);
nand U7164 (N_7164,N_6853,N_6818);
xnor U7165 (N_7165,N_6694,N_6603);
nor U7166 (N_7166,N_6680,N_6731);
xnor U7167 (N_7167,N_6756,N_6656);
nor U7168 (N_7168,N_6706,N_6739);
xnor U7169 (N_7169,N_6763,N_6887);
or U7170 (N_7170,N_6763,N_6703);
and U7171 (N_7171,N_6679,N_6804);
xnor U7172 (N_7172,N_6719,N_6852);
and U7173 (N_7173,N_6793,N_6644);
nand U7174 (N_7174,N_6840,N_6764);
and U7175 (N_7175,N_6783,N_6747);
nand U7176 (N_7176,N_6725,N_6678);
nand U7177 (N_7177,N_6736,N_6799);
nand U7178 (N_7178,N_6719,N_6668);
and U7179 (N_7179,N_6858,N_6825);
nand U7180 (N_7180,N_6707,N_6686);
or U7181 (N_7181,N_6651,N_6667);
and U7182 (N_7182,N_6749,N_6734);
and U7183 (N_7183,N_6758,N_6896);
or U7184 (N_7184,N_6782,N_6826);
nor U7185 (N_7185,N_6643,N_6718);
or U7186 (N_7186,N_6676,N_6764);
nand U7187 (N_7187,N_6785,N_6805);
nand U7188 (N_7188,N_6855,N_6655);
or U7189 (N_7189,N_6802,N_6608);
nor U7190 (N_7190,N_6664,N_6777);
or U7191 (N_7191,N_6805,N_6647);
xor U7192 (N_7192,N_6764,N_6703);
nor U7193 (N_7193,N_6624,N_6746);
and U7194 (N_7194,N_6871,N_6628);
nand U7195 (N_7195,N_6781,N_6701);
nand U7196 (N_7196,N_6738,N_6625);
xor U7197 (N_7197,N_6682,N_6691);
nor U7198 (N_7198,N_6640,N_6820);
and U7199 (N_7199,N_6791,N_6726);
and U7200 (N_7200,N_7068,N_7053);
nand U7201 (N_7201,N_6969,N_7149);
or U7202 (N_7202,N_7180,N_7148);
and U7203 (N_7203,N_6970,N_6972);
nor U7204 (N_7204,N_6949,N_7135);
and U7205 (N_7205,N_7170,N_7097);
nor U7206 (N_7206,N_7036,N_7160);
nand U7207 (N_7207,N_6911,N_7134);
nor U7208 (N_7208,N_7037,N_7194);
nand U7209 (N_7209,N_7051,N_7031);
nor U7210 (N_7210,N_6989,N_7086);
nand U7211 (N_7211,N_7140,N_6954);
nand U7212 (N_7212,N_7063,N_7105);
xor U7213 (N_7213,N_7023,N_6927);
xor U7214 (N_7214,N_7141,N_7038);
or U7215 (N_7215,N_6980,N_7079);
and U7216 (N_7216,N_7174,N_6978);
and U7217 (N_7217,N_7022,N_7106);
and U7218 (N_7218,N_7027,N_6918);
and U7219 (N_7219,N_6925,N_6942);
xor U7220 (N_7220,N_6923,N_6904);
or U7221 (N_7221,N_7030,N_7172);
or U7222 (N_7222,N_6937,N_7083);
nand U7223 (N_7223,N_7102,N_7146);
or U7224 (N_7224,N_7156,N_7044);
xnor U7225 (N_7225,N_6930,N_6938);
or U7226 (N_7226,N_6908,N_6910);
or U7227 (N_7227,N_7039,N_7055);
and U7228 (N_7228,N_7158,N_7162);
nor U7229 (N_7229,N_6964,N_7154);
and U7230 (N_7230,N_6992,N_7188);
nor U7231 (N_7231,N_6907,N_6955);
xnor U7232 (N_7232,N_6962,N_7192);
xor U7233 (N_7233,N_7076,N_7074);
and U7234 (N_7234,N_7057,N_6924);
xor U7235 (N_7235,N_7157,N_6916);
or U7236 (N_7236,N_6965,N_6966);
nor U7237 (N_7237,N_6919,N_7080);
xnor U7238 (N_7238,N_7011,N_7019);
nand U7239 (N_7239,N_6906,N_7016);
and U7240 (N_7240,N_7077,N_7175);
nor U7241 (N_7241,N_7088,N_7100);
xnor U7242 (N_7242,N_6984,N_7071);
nor U7243 (N_7243,N_7065,N_6905);
nor U7244 (N_7244,N_7118,N_7090);
and U7245 (N_7245,N_7082,N_7042);
and U7246 (N_7246,N_7033,N_7126);
nand U7247 (N_7247,N_6976,N_6933);
xor U7248 (N_7248,N_7072,N_6913);
or U7249 (N_7249,N_7147,N_6993);
nor U7250 (N_7250,N_7161,N_7073);
xnor U7251 (N_7251,N_7142,N_6994);
or U7252 (N_7252,N_7195,N_7110);
and U7253 (N_7253,N_7052,N_7166);
nand U7254 (N_7254,N_6929,N_7003);
nor U7255 (N_7255,N_7153,N_7178);
nor U7256 (N_7256,N_7167,N_7010);
xor U7257 (N_7257,N_7165,N_7133);
or U7258 (N_7258,N_6983,N_6956);
nand U7259 (N_7259,N_7060,N_7089);
xnor U7260 (N_7260,N_7176,N_7115);
and U7261 (N_7261,N_7096,N_7177);
or U7262 (N_7262,N_7066,N_6947);
nand U7263 (N_7263,N_6932,N_7091);
and U7264 (N_7264,N_6999,N_7171);
nand U7265 (N_7265,N_7017,N_6997);
nand U7266 (N_7266,N_6940,N_6982);
nand U7267 (N_7267,N_7056,N_7186);
xor U7268 (N_7268,N_7007,N_7191);
or U7269 (N_7269,N_7163,N_6914);
xnor U7270 (N_7270,N_6939,N_7041);
and U7271 (N_7271,N_6958,N_7045);
xnor U7272 (N_7272,N_7168,N_6936);
or U7273 (N_7273,N_6934,N_7067);
xnor U7274 (N_7274,N_7182,N_7032);
xnor U7275 (N_7275,N_6995,N_7093);
xor U7276 (N_7276,N_6957,N_6901);
and U7277 (N_7277,N_7179,N_7150);
and U7278 (N_7278,N_7005,N_7001);
nand U7279 (N_7279,N_7169,N_6990);
xor U7280 (N_7280,N_7081,N_7139);
nand U7281 (N_7281,N_7025,N_7087);
xor U7282 (N_7282,N_7099,N_7199);
nor U7283 (N_7283,N_7187,N_7014);
nand U7284 (N_7284,N_6960,N_6959);
xor U7285 (N_7285,N_7159,N_7061);
nand U7286 (N_7286,N_7069,N_7152);
xor U7287 (N_7287,N_7018,N_7155);
nor U7288 (N_7288,N_7059,N_7128);
and U7289 (N_7289,N_7123,N_7181);
nor U7290 (N_7290,N_7026,N_7004);
or U7291 (N_7291,N_6988,N_6985);
xor U7292 (N_7292,N_7173,N_7119);
nor U7293 (N_7293,N_7050,N_6967);
and U7294 (N_7294,N_7107,N_6903);
and U7295 (N_7295,N_7129,N_6998);
nand U7296 (N_7296,N_7046,N_7136);
xor U7297 (N_7297,N_6946,N_7108);
or U7298 (N_7298,N_6926,N_7092);
nand U7299 (N_7299,N_6979,N_6975);
or U7300 (N_7300,N_6987,N_7183);
or U7301 (N_7301,N_7125,N_7198);
nor U7302 (N_7302,N_7138,N_7095);
or U7303 (N_7303,N_7084,N_7164);
nand U7304 (N_7304,N_7137,N_6952);
or U7305 (N_7305,N_7151,N_6996);
nor U7306 (N_7306,N_7144,N_6909);
nand U7307 (N_7307,N_7127,N_6920);
nand U7308 (N_7308,N_7013,N_7064);
nor U7309 (N_7309,N_7113,N_7043);
nand U7310 (N_7310,N_7029,N_7070);
xnor U7311 (N_7311,N_7000,N_7028);
nand U7312 (N_7312,N_7075,N_7062);
xor U7313 (N_7313,N_6991,N_7193);
xor U7314 (N_7314,N_7112,N_7190);
nand U7315 (N_7315,N_7103,N_7085);
xnor U7316 (N_7316,N_7098,N_6963);
xor U7317 (N_7317,N_6902,N_7012);
nand U7318 (N_7318,N_7021,N_7124);
or U7319 (N_7319,N_7002,N_7143);
nand U7320 (N_7320,N_7109,N_6948);
nor U7321 (N_7321,N_6951,N_7047);
nor U7322 (N_7322,N_7049,N_7189);
xor U7323 (N_7323,N_7145,N_6928);
or U7324 (N_7324,N_6986,N_7048);
and U7325 (N_7325,N_6977,N_7034);
and U7326 (N_7326,N_6950,N_6968);
nor U7327 (N_7327,N_7078,N_6943);
nor U7328 (N_7328,N_7121,N_7185);
nor U7329 (N_7329,N_7020,N_6941);
nand U7330 (N_7330,N_7122,N_6981);
and U7331 (N_7331,N_6912,N_6921);
and U7332 (N_7332,N_7094,N_6974);
nand U7333 (N_7333,N_6922,N_7008);
xnor U7334 (N_7334,N_7101,N_6931);
nor U7335 (N_7335,N_7009,N_7015);
or U7336 (N_7336,N_7196,N_6900);
or U7337 (N_7337,N_7040,N_7116);
and U7338 (N_7338,N_6917,N_7114);
or U7339 (N_7339,N_7111,N_7130);
nand U7340 (N_7340,N_7006,N_7197);
nand U7341 (N_7341,N_6944,N_6973);
or U7342 (N_7342,N_7131,N_6935);
nand U7343 (N_7343,N_7035,N_6961);
or U7344 (N_7344,N_7058,N_6971);
xnor U7345 (N_7345,N_7184,N_7132);
nand U7346 (N_7346,N_7104,N_6945);
or U7347 (N_7347,N_7117,N_6915);
nor U7348 (N_7348,N_6953,N_7054);
nand U7349 (N_7349,N_7024,N_7120);
xor U7350 (N_7350,N_6906,N_7010);
or U7351 (N_7351,N_7129,N_7156);
and U7352 (N_7352,N_6928,N_7188);
and U7353 (N_7353,N_6902,N_7018);
nor U7354 (N_7354,N_7101,N_6945);
nor U7355 (N_7355,N_6907,N_6983);
xnor U7356 (N_7356,N_6922,N_7089);
or U7357 (N_7357,N_7158,N_7053);
or U7358 (N_7358,N_7187,N_7057);
xnor U7359 (N_7359,N_7197,N_7175);
nand U7360 (N_7360,N_6931,N_7054);
and U7361 (N_7361,N_7199,N_7122);
nor U7362 (N_7362,N_6945,N_7080);
or U7363 (N_7363,N_6935,N_7169);
and U7364 (N_7364,N_7124,N_7080);
and U7365 (N_7365,N_6915,N_6907);
nand U7366 (N_7366,N_7149,N_6922);
nor U7367 (N_7367,N_6930,N_6910);
or U7368 (N_7368,N_6963,N_7103);
xor U7369 (N_7369,N_7058,N_7086);
xnor U7370 (N_7370,N_7027,N_7055);
xor U7371 (N_7371,N_7061,N_7047);
nand U7372 (N_7372,N_7025,N_7070);
and U7373 (N_7373,N_6947,N_7180);
xnor U7374 (N_7374,N_7185,N_6992);
nand U7375 (N_7375,N_7033,N_6959);
nand U7376 (N_7376,N_7061,N_6985);
nor U7377 (N_7377,N_7055,N_7172);
xnor U7378 (N_7378,N_6988,N_7040);
nor U7379 (N_7379,N_7185,N_6990);
or U7380 (N_7380,N_7156,N_7178);
and U7381 (N_7381,N_7127,N_7156);
and U7382 (N_7382,N_6915,N_7061);
or U7383 (N_7383,N_7098,N_6966);
and U7384 (N_7384,N_6904,N_7053);
and U7385 (N_7385,N_7043,N_7039);
nand U7386 (N_7386,N_6920,N_6979);
xor U7387 (N_7387,N_6965,N_7184);
and U7388 (N_7388,N_7139,N_7132);
xnor U7389 (N_7389,N_7076,N_7032);
or U7390 (N_7390,N_7156,N_6992);
xor U7391 (N_7391,N_7094,N_7177);
or U7392 (N_7392,N_7104,N_6954);
nand U7393 (N_7393,N_7060,N_7040);
nor U7394 (N_7394,N_7088,N_6928);
xor U7395 (N_7395,N_6928,N_7031);
or U7396 (N_7396,N_6975,N_7133);
and U7397 (N_7397,N_6948,N_7002);
and U7398 (N_7398,N_7060,N_6949);
nor U7399 (N_7399,N_7048,N_7005);
nand U7400 (N_7400,N_6915,N_7086);
or U7401 (N_7401,N_7129,N_7090);
or U7402 (N_7402,N_7085,N_7006);
nand U7403 (N_7403,N_6972,N_6919);
nand U7404 (N_7404,N_7010,N_7141);
and U7405 (N_7405,N_6977,N_7186);
nor U7406 (N_7406,N_6901,N_7151);
nand U7407 (N_7407,N_6957,N_7188);
or U7408 (N_7408,N_6957,N_7142);
and U7409 (N_7409,N_7156,N_6943);
and U7410 (N_7410,N_7110,N_7060);
or U7411 (N_7411,N_6944,N_7028);
nor U7412 (N_7412,N_6967,N_7162);
nor U7413 (N_7413,N_6953,N_7032);
or U7414 (N_7414,N_7166,N_6952);
or U7415 (N_7415,N_7124,N_6999);
nor U7416 (N_7416,N_6951,N_7153);
xor U7417 (N_7417,N_6929,N_6957);
xnor U7418 (N_7418,N_6934,N_7192);
or U7419 (N_7419,N_7042,N_7025);
xnor U7420 (N_7420,N_6997,N_7152);
nand U7421 (N_7421,N_6935,N_7158);
nand U7422 (N_7422,N_7007,N_6998);
and U7423 (N_7423,N_7025,N_7037);
nor U7424 (N_7424,N_6908,N_7127);
or U7425 (N_7425,N_6949,N_7178);
nand U7426 (N_7426,N_7168,N_7022);
xor U7427 (N_7427,N_7141,N_7114);
and U7428 (N_7428,N_6927,N_6969);
nor U7429 (N_7429,N_7060,N_7022);
xnor U7430 (N_7430,N_6933,N_7097);
or U7431 (N_7431,N_7137,N_6917);
and U7432 (N_7432,N_7106,N_6918);
and U7433 (N_7433,N_6926,N_7014);
and U7434 (N_7434,N_6958,N_6975);
or U7435 (N_7435,N_6973,N_7165);
nand U7436 (N_7436,N_7037,N_7000);
or U7437 (N_7437,N_6900,N_7127);
nand U7438 (N_7438,N_7189,N_6934);
and U7439 (N_7439,N_7022,N_6980);
xnor U7440 (N_7440,N_6941,N_6967);
or U7441 (N_7441,N_7151,N_6953);
nand U7442 (N_7442,N_7139,N_6974);
nor U7443 (N_7443,N_6984,N_6926);
nand U7444 (N_7444,N_6972,N_7092);
or U7445 (N_7445,N_7055,N_6915);
and U7446 (N_7446,N_7103,N_6975);
xor U7447 (N_7447,N_7132,N_6989);
nor U7448 (N_7448,N_7145,N_7063);
and U7449 (N_7449,N_7176,N_6934);
xor U7450 (N_7450,N_6923,N_6919);
and U7451 (N_7451,N_7036,N_7112);
and U7452 (N_7452,N_7175,N_6919);
nand U7453 (N_7453,N_7033,N_7176);
or U7454 (N_7454,N_7032,N_6975);
and U7455 (N_7455,N_6914,N_7034);
and U7456 (N_7456,N_6938,N_6910);
xor U7457 (N_7457,N_7009,N_6946);
and U7458 (N_7458,N_6982,N_6911);
nand U7459 (N_7459,N_6940,N_7027);
and U7460 (N_7460,N_6950,N_7035);
xor U7461 (N_7461,N_7128,N_7055);
and U7462 (N_7462,N_6975,N_7099);
and U7463 (N_7463,N_6937,N_7176);
nand U7464 (N_7464,N_7135,N_7078);
and U7465 (N_7465,N_7139,N_7197);
and U7466 (N_7466,N_7041,N_7075);
nand U7467 (N_7467,N_7078,N_7044);
nor U7468 (N_7468,N_7177,N_7164);
xnor U7469 (N_7469,N_7056,N_7033);
or U7470 (N_7470,N_7000,N_6954);
and U7471 (N_7471,N_7132,N_6970);
nor U7472 (N_7472,N_7139,N_7185);
or U7473 (N_7473,N_7165,N_7054);
xnor U7474 (N_7474,N_7071,N_6989);
and U7475 (N_7475,N_6997,N_6949);
xor U7476 (N_7476,N_7163,N_7074);
nor U7477 (N_7477,N_7042,N_6927);
nor U7478 (N_7478,N_7138,N_7106);
or U7479 (N_7479,N_7085,N_6909);
and U7480 (N_7480,N_7197,N_6902);
or U7481 (N_7481,N_7147,N_7083);
or U7482 (N_7482,N_7134,N_6998);
and U7483 (N_7483,N_7072,N_7021);
xnor U7484 (N_7484,N_7177,N_7097);
xor U7485 (N_7485,N_7143,N_7152);
and U7486 (N_7486,N_7035,N_7130);
xnor U7487 (N_7487,N_7077,N_6949);
nand U7488 (N_7488,N_7190,N_7131);
or U7489 (N_7489,N_7037,N_6944);
and U7490 (N_7490,N_6945,N_7021);
nor U7491 (N_7491,N_6968,N_7181);
nor U7492 (N_7492,N_7133,N_7071);
and U7493 (N_7493,N_6962,N_7043);
and U7494 (N_7494,N_6907,N_6950);
nor U7495 (N_7495,N_6920,N_7116);
xnor U7496 (N_7496,N_7196,N_6906);
and U7497 (N_7497,N_7119,N_6913);
nor U7498 (N_7498,N_7111,N_7067);
xnor U7499 (N_7499,N_6964,N_6933);
nand U7500 (N_7500,N_7385,N_7452);
nor U7501 (N_7501,N_7498,N_7282);
xor U7502 (N_7502,N_7399,N_7367);
nor U7503 (N_7503,N_7233,N_7309);
nor U7504 (N_7504,N_7403,N_7204);
and U7505 (N_7505,N_7372,N_7435);
xor U7506 (N_7506,N_7359,N_7247);
or U7507 (N_7507,N_7412,N_7261);
nor U7508 (N_7508,N_7393,N_7405);
and U7509 (N_7509,N_7292,N_7356);
xnor U7510 (N_7510,N_7303,N_7260);
nand U7511 (N_7511,N_7248,N_7293);
xor U7512 (N_7512,N_7246,N_7387);
and U7513 (N_7513,N_7271,N_7486);
nand U7514 (N_7514,N_7209,N_7379);
or U7515 (N_7515,N_7341,N_7213);
xor U7516 (N_7516,N_7388,N_7242);
nand U7517 (N_7517,N_7304,N_7258);
xnor U7518 (N_7518,N_7429,N_7227);
or U7519 (N_7519,N_7278,N_7232);
nand U7520 (N_7520,N_7342,N_7376);
nor U7521 (N_7521,N_7462,N_7308);
nand U7522 (N_7522,N_7479,N_7208);
nand U7523 (N_7523,N_7382,N_7280);
nand U7524 (N_7524,N_7275,N_7263);
nor U7525 (N_7525,N_7229,N_7255);
nor U7526 (N_7526,N_7228,N_7315);
xor U7527 (N_7527,N_7432,N_7250);
xnor U7528 (N_7528,N_7323,N_7215);
or U7529 (N_7529,N_7224,N_7243);
and U7530 (N_7530,N_7384,N_7348);
nand U7531 (N_7531,N_7488,N_7443);
nand U7532 (N_7532,N_7391,N_7414);
nor U7533 (N_7533,N_7428,N_7395);
and U7534 (N_7534,N_7463,N_7400);
nand U7535 (N_7535,N_7310,N_7381);
nand U7536 (N_7536,N_7217,N_7201);
and U7537 (N_7537,N_7499,N_7410);
nor U7538 (N_7538,N_7324,N_7357);
nor U7539 (N_7539,N_7354,N_7449);
nand U7540 (N_7540,N_7219,N_7313);
nor U7541 (N_7541,N_7458,N_7472);
xnor U7542 (N_7542,N_7314,N_7344);
and U7543 (N_7543,N_7411,N_7477);
nor U7544 (N_7544,N_7312,N_7370);
xor U7545 (N_7545,N_7316,N_7267);
nor U7546 (N_7546,N_7439,N_7471);
and U7547 (N_7547,N_7497,N_7407);
nor U7548 (N_7548,N_7426,N_7490);
nor U7549 (N_7549,N_7301,N_7257);
nor U7550 (N_7550,N_7205,N_7493);
nand U7551 (N_7551,N_7392,N_7339);
or U7552 (N_7552,N_7496,N_7427);
or U7553 (N_7553,N_7328,N_7203);
or U7554 (N_7554,N_7413,N_7396);
and U7555 (N_7555,N_7470,N_7419);
or U7556 (N_7556,N_7474,N_7320);
nor U7557 (N_7557,N_7216,N_7454);
and U7558 (N_7558,N_7417,N_7211);
nand U7559 (N_7559,N_7305,N_7333);
nand U7560 (N_7560,N_7234,N_7398);
and U7561 (N_7561,N_7409,N_7290);
xnor U7562 (N_7562,N_7330,N_7221);
or U7563 (N_7563,N_7289,N_7346);
or U7564 (N_7564,N_7279,N_7369);
or U7565 (N_7565,N_7338,N_7481);
nor U7566 (N_7566,N_7425,N_7416);
nand U7567 (N_7567,N_7302,N_7438);
nand U7568 (N_7568,N_7321,N_7251);
xnor U7569 (N_7569,N_7277,N_7451);
nor U7570 (N_7570,N_7422,N_7483);
or U7571 (N_7571,N_7453,N_7467);
or U7572 (N_7572,N_7448,N_7230);
xnor U7573 (N_7573,N_7495,N_7404);
and U7574 (N_7574,N_7352,N_7468);
nand U7575 (N_7575,N_7340,N_7286);
nand U7576 (N_7576,N_7469,N_7420);
or U7577 (N_7577,N_7358,N_7202);
or U7578 (N_7578,N_7431,N_7223);
and U7579 (N_7579,N_7457,N_7252);
nor U7580 (N_7580,N_7424,N_7386);
or U7581 (N_7581,N_7371,N_7368);
and U7582 (N_7582,N_7222,N_7225);
nor U7583 (N_7583,N_7478,N_7249);
xnor U7584 (N_7584,N_7241,N_7446);
and U7585 (N_7585,N_7297,N_7437);
nor U7586 (N_7586,N_7430,N_7406);
nand U7587 (N_7587,N_7461,N_7281);
and U7588 (N_7588,N_7360,N_7335);
nand U7589 (N_7589,N_7492,N_7377);
nor U7590 (N_7590,N_7415,N_7363);
nand U7591 (N_7591,N_7487,N_7390);
nand U7592 (N_7592,N_7237,N_7466);
xor U7593 (N_7593,N_7259,N_7361);
or U7594 (N_7594,N_7480,N_7264);
nand U7595 (N_7595,N_7475,N_7245);
xnor U7596 (N_7596,N_7295,N_7383);
nand U7597 (N_7597,N_7300,N_7317);
and U7598 (N_7598,N_7418,N_7307);
or U7599 (N_7599,N_7421,N_7455);
and U7600 (N_7600,N_7345,N_7273);
or U7601 (N_7601,N_7401,N_7433);
or U7602 (N_7602,N_7254,N_7253);
nand U7603 (N_7603,N_7287,N_7465);
nand U7604 (N_7604,N_7374,N_7394);
or U7605 (N_7605,N_7336,N_7351);
nand U7606 (N_7606,N_7366,N_7235);
or U7607 (N_7607,N_7276,N_7423);
nand U7608 (N_7608,N_7268,N_7375);
nand U7609 (N_7609,N_7355,N_7491);
or U7610 (N_7610,N_7265,N_7460);
nand U7611 (N_7611,N_7206,N_7402);
xor U7612 (N_7612,N_7484,N_7212);
nand U7613 (N_7613,N_7231,N_7343);
nand U7614 (N_7614,N_7482,N_7331);
or U7615 (N_7615,N_7362,N_7378);
nand U7616 (N_7616,N_7238,N_7288);
nand U7617 (N_7617,N_7236,N_7311);
and U7618 (N_7618,N_7347,N_7269);
xnor U7619 (N_7619,N_7456,N_7485);
and U7620 (N_7620,N_7389,N_7318);
xor U7621 (N_7621,N_7239,N_7207);
xnor U7622 (N_7622,N_7329,N_7332);
nand U7623 (N_7623,N_7337,N_7244);
and U7624 (N_7624,N_7306,N_7436);
nor U7625 (N_7625,N_7272,N_7353);
nor U7626 (N_7626,N_7325,N_7322);
nand U7627 (N_7627,N_7464,N_7440);
or U7628 (N_7628,N_7326,N_7334);
xor U7629 (N_7629,N_7220,N_7291);
xnor U7630 (N_7630,N_7283,N_7296);
nand U7631 (N_7631,N_7489,N_7365);
nor U7632 (N_7632,N_7285,N_7270);
nand U7633 (N_7633,N_7445,N_7459);
or U7634 (N_7634,N_7350,N_7218);
or U7635 (N_7635,N_7444,N_7397);
nand U7636 (N_7636,N_7319,N_7298);
xnor U7637 (N_7637,N_7256,N_7210);
xnor U7638 (N_7638,N_7274,N_7373);
xnor U7639 (N_7639,N_7380,N_7284);
or U7640 (N_7640,N_7441,N_7266);
nor U7641 (N_7641,N_7262,N_7299);
nor U7642 (N_7642,N_7226,N_7214);
nand U7643 (N_7643,N_7327,N_7434);
and U7644 (N_7644,N_7408,N_7447);
nand U7645 (N_7645,N_7476,N_7200);
and U7646 (N_7646,N_7240,N_7473);
nand U7647 (N_7647,N_7364,N_7442);
or U7648 (N_7648,N_7294,N_7450);
xor U7649 (N_7649,N_7349,N_7494);
nand U7650 (N_7650,N_7415,N_7237);
xnor U7651 (N_7651,N_7392,N_7234);
nand U7652 (N_7652,N_7480,N_7481);
nand U7653 (N_7653,N_7329,N_7337);
and U7654 (N_7654,N_7244,N_7431);
xor U7655 (N_7655,N_7461,N_7389);
and U7656 (N_7656,N_7357,N_7430);
xor U7657 (N_7657,N_7470,N_7218);
or U7658 (N_7658,N_7278,N_7214);
or U7659 (N_7659,N_7273,N_7331);
nor U7660 (N_7660,N_7235,N_7280);
or U7661 (N_7661,N_7274,N_7299);
nor U7662 (N_7662,N_7290,N_7336);
nor U7663 (N_7663,N_7471,N_7344);
nor U7664 (N_7664,N_7307,N_7421);
xor U7665 (N_7665,N_7202,N_7279);
or U7666 (N_7666,N_7414,N_7313);
nand U7667 (N_7667,N_7202,N_7241);
nor U7668 (N_7668,N_7486,N_7497);
or U7669 (N_7669,N_7230,N_7323);
nand U7670 (N_7670,N_7470,N_7480);
and U7671 (N_7671,N_7219,N_7214);
nand U7672 (N_7672,N_7448,N_7466);
and U7673 (N_7673,N_7216,N_7462);
and U7674 (N_7674,N_7363,N_7469);
xnor U7675 (N_7675,N_7476,N_7498);
xnor U7676 (N_7676,N_7208,N_7304);
nor U7677 (N_7677,N_7261,N_7490);
nor U7678 (N_7678,N_7468,N_7213);
nor U7679 (N_7679,N_7487,N_7350);
nand U7680 (N_7680,N_7447,N_7487);
xnor U7681 (N_7681,N_7219,N_7258);
or U7682 (N_7682,N_7230,N_7499);
xor U7683 (N_7683,N_7240,N_7234);
or U7684 (N_7684,N_7327,N_7487);
nand U7685 (N_7685,N_7276,N_7320);
nand U7686 (N_7686,N_7218,N_7221);
and U7687 (N_7687,N_7269,N_7222);
nand U7688 (N_7688,N_7367,N_7499);
and U7689 (N_7689,N_7391,N_7261);
nor U7690 (N_7690,N_7267,N_7424);
and U7691 (N_7691,N_7370,N_7403);
or U7692 (N_7692,N_7357,N_7244);
nor U7693 (N_7693,N_7445,N_7477);
and U7694 (N_7694,N_7454,N_7386);
or U7695 (N_7695,N_7249,N_7447);
nand U7696 (N_7696,N_7462,N_7445);
xnor U7697 (N_7697,N_7434,N_7491);
or U7698 (N_7698,N_7242,N_7489);
nand U7699 (N_7699,N_7249,N_7387);
xnor U7700 (N_7700,N_7360,N_7430);
xnor U7701 (N_7701,N_7272,N_7270);
and U7702 (N_7702,N_7380,N_7365);
and U7703 (N_7703,N_7324,N_7331);
and U7704 (N_7704,N_7252,N_7366);
xor U7705 (N_7705,N_7378,N_7202);
and U7706 (N_7706,N_7276,N_7427);
and U7707 (N_7707,N_7212,N_7431);
xor U7708 (N_7708,N_7307,N_7274);
nor U7709 (N_7709,N_7249,N_7400);
nor U7710 (N_7710,N_7269,N_7390);
nor U7711 (N_7711,N_7329,N_7250);
nand U7712 (N_7712,N_7326,N_7442);
nor U7713 (N_7713,N_7432,N_7456);
nor U7714 (N_7714,N_7459,N_7420);
nand U7715 (N_7715,N_7270,N_7409);
or U7716 (N_7716,N_7433,N_7388);
nor U7717 (N_7717,N_7460,N_7497);
xnor U7718 (N_7718,N_7445,N_7437);
nor U7719 (N_7719,N_7361,N_7275);
nor U7720 (N_7720,N_7449,N_7316);
or U7721 (N_7721,N_7445,N_7417);
nand U7722 (N_7722,N_7456,N_7448);
nor U7723 (N_7723,N_7371,N_7333);
xor U7724 (N_7724,N_7311,N_7459);
and U7725 (N_7725,N_7470,N_7479);
nor U7726 (N_7726,N_7299,N_7297);
or U7727 (N_7727,N_7486,N_7218);
or U7728 (N_7728,N_7418,N_7251);
and U7729 (N_7729,N_7329,N_7301);
or U7730 (N_7730,N_7422,N_7320);
nor U7731 (N_7731,N_7252,N_7410);
and U7732 (N_7732,N_7495,N_7212);
nand U7733 (N_7733,N_7348,N_7402);
xor U7734 (N_7734,N_7488,N_7242);
nand U7735 (N_7735,N_7488,N_7317);
xnor U7736 (N_7736,N_7378,N_7449);
nor U7737 (N_7737,N_7467,N_7320);
nand U7738 (N_7738,N_7356,N_7303);
xor U7739 (N_7739,N_7324,N_7280);
xor U7740 (N_7740,N_7489,N_7297);
nor U7741 (N_7741,N_7442,N_7356);
xnor U7742 (N_7742,N_7485,N_7438);
and U7743 (N_7743,N_7472,N_7429);
xor U7744 (N_7744,N_7454,N_7272);
and U7745 (N_7745,N_7465,N_7301);
nor U7746 (N_7746,N_7466,N_7461);
and U7747 (N_7747,N_7496,N_7300);
nand U7748 (N_7748,N_7399,N_7334);
or U7749 (N_7749,N_7353,N_7380);
and U7750 (N_7750,N_7381,N_7405);
and U7751 (N_7751,N_7447,N_7290);
and U7752 (N_7752,N_7464,N_7271);
xnor U7753 (N_7753,N_7286,N_7230);
xor U7754 (N_7754,N_7478,N_7340);
or U7755 (N_7755,N_7295,N_7234);
and U7756 (N_7756,N_7281,N_7227);
xor U7757 (N_7757,N_7458,N_7213);
nand U7758 (N_7758,N_7441,N_7275);
and U7759 (N_7759,N_7468,N_7462);
nor U7760 (N_7760,N_7233,N_7356);
nand U7761 (N_7761,N_7380,N_7350);
xnor U7762 (N_7762,N_7362,N_7223);
or U7763 (N_7763,N_7408,N_7237);
nand U7764 (N_7764,N_7394,N_7200);
or U7765 (N_7765,N_7318,N_7472);
and U7766 (N_7766,N_7471,N_7470);
nor U7767 (N_7767,N_7470,N_7288);
nor U7768 (N_7768,N_7222,N_7230);
nor U7769 (N_7769,N_7374,N_7377);
or U7770 (N_7770,N_7323,N_7363);
nor U7771 (N_7771,N_7467,N_7389);
and U7772 (N_7772,N_7340,N_7273);
and U7773 (N_7773,N_7454,N_7298);
or U7774 (N_7774,N_7388,N_7321);
or U7775 (N_7775,N_7291,N_7446);
or U7776 (N_7776,N_7494,N_7266);
nand U7777 (N_7777,N_7460,N_7310);
xor U7778 (N_7778,N_7284,N_7461);
xor U7779 (N_7779,N_7225,N_7273);
or U7780 (N_7780,N_7499,N_7419);
and U7781 (N_7781,N_7252,N_7413);
xnor U7782 (N_7782,N_7444,N_7357);
and U7783 (N_7783,N_7333,N_7328);
or U7784 (N_7784,N_7301,N_7455);
or U7785 (N_7785,N_7327,N_7400);
or U7786 (N_7786,N_7245,N_7338);
nor U7787 (N_7787,N_7371,N_7389);
xnor U7788 (N_7788,N_7446,N_7317);
or U7789 (N_7789,N_7358,N_7224);
nand U7790 (N_7790,N_7325,N_7288);
nor U7791 (N_7791,N_7484,N_7398);
nand U7792 (N_7792,N_7375,N_7371);
nor U7793 (N_7793,N_7361,N_7377);
xor U7794 (N_7794,N_7458,N_7371);
nor U7795 (N_7795,N_7243,N_7366);
nand U7796 (N_7796,N_7376,N_7477);
nand U7797 (N_7797,N_7451,N_7363);
nor U7798 (N_7798,N_7239,N_7257);
nand U7799 (N_7799,N_7429,N_7399);
nand U7800 (N_7800,N_7724,N_7608);
or U7801 (N_7801,N_7697,N_7506);
nand U7802 (N_7802,N_7541,N_7763);
or U7803 (N_7803,N_7731,N_7781);
nor U7804 (N_7804,N_7571,N_7574);
nand U7805 (N_7805,N_7644,N_7727);
xor U7806 (N_7806,N_7767,N_7569);
xor U7807 (N_7807,N_7699,N_7589);
or U7808 (N_7808,N_7621,N_7796);
and U7809 (N_7809,N_7746,N_7726);
nor U7810 (N_7810,N_7598,N_7749);
nand U7811 (N_7811,N_7691,N_7704);
or U7812 (N_7812,N_7680,N_7786);
nand U7813 (N_7813,N_7531,N_7539);
xnor U7814 (N_7814,N_7661,N_7538);
nor U7815 (N_7815,N_7532,N_7640);
nor U7816 (N_7816,N_7755,N_7504);
or U7817 (N_7817,N_7734,N_7747);
and U7818 (N_7818,N_7718,N_7534);
nand U7819 (N_7819,N_7735,N_7638);
or U7820 (N_7820,N_7525,N_7785);
nor U7821 (N_7821,N_7620,N_7535);
nor U7822 (N_7822,N_7779,N_7543);
and U7823 (N_7823,N_7723,N_7716);
or U7824 (N_7824,N_7593,N_7740);
nand U7825 (N_7825,N_7629,N_7766);
xnor U7826 (N_7826,N_7519,N_7505);
and U7827 (N_7827,N_7641,N_7592);
nand U7828 (N_7828,N_7752,N_7520);
and U7829 (N_7829,N_7654,N_7701);
xor U7830 (N_7830,N_7725,N_7707);
and U7831 (N_7831,N_7764,N_7584);
nor U7832 (N_7832,N_7544,N_7582);
and U7833 (N_7833,N_7774,N_7559);
nor U7834 (N_7834,N_7526,N_7667);
nor U7835 (N_7835,N_7579,N_7791);
xnor U7836 (N_7836,N_7750,N_7770);
xnor U7837 (N_7837,N_7635,N_7596);
xor U7838 (N_7838,N_7687,N_7696);
nor U7839 (N_7839,N_7702,N_7551);
nand U7840 (N_7840,N_7662,N_7633);
and U7841 (N_7841,N_7632,N_7511);
or U7842 (N_7842,N_7686,N_7617);
or U7843 (N_7843,N_7510,N_7722);
nand U7844 (N_7844,N_7650,N_7657);
or U7845 (N_7845,N_7646,N_7760);
xor U7846 (N_7846,N_7611,N_7560);
nor U7847 (N_7847,N_7728,N_7683);
and U7848 (N_7848,N_7768,N_7736);
xor U7849 (N_7849,N_7500,N_7578);
and U7850 (N_7850,N_7795,N_7773);
and U7851 (N_7851,N_7645,N_7743);
nor U7852 (N_7852,N_7706,N_7518);
and U7853 (N_7853,N_7676,N_7503);
nand U7854 (N_7854,N_7690,N_7637);
and U7855 (N_7855,N_7587,N_7549);
or U7856 (N_7856,N_7567,N_7663);
nor U7857 (N_7857,N_7782,N_7751);
nor U7858 (N_7858,N_7554,N_7776);
nor U7859 (N_7859,N_7517,N_7649);
nand U7860 (N_7860,N_7692,N_7636);
or U7861 (N_7861,N_7721,N_7792);
or U7862 (N_7862,N_7788,N_7533);
or U7863 (N_7863,N_7612,N_7597);
and U7864 (N_7864,N_7527,N_7542);
and U7865 (N_7865,N_7540,N_7547);
and U7866 (N_7866,N_7700,N_7684);
or U7867 (N_7867,N_7741,N_7643);
nand U7868 (N_7868,N_7798,N_7745);
or U7869 (N_7869,N_7614,N_7713);
or U7870 (N_7870,N_7647,N_7717);
or U7871 (N_7871,N_7670,N_7607);
xor U7872 (N_7872,N_7602,N_7610);
nor U7873 (N_7873,N_7674,N_7682);
and U7874 (N_7874,N_7628,N_7545);
and U7875 (N_7875,N_7631,N_7573);
nor U7876 (N_7876,N_7627,N_7673);
nor U7877 (N_7877,N_7757,N_7732);
or U7878 (N_7878,N_7705,N_7591);
xor U7879 (N_7879,N_7733,N_7660);
or U7880 (N_7880,N_7585,N_7685);
nor U7881 (N_7881,N_7677,N_7659);
and U7882 (N_7882,N_7555,N_7710);
nand U7883 (N_7883,N_7615,N_7797);
or U7884 (N_7884,N_7548,N_7738);
or U7885 (N_7885,N_7783,N_7678);
xor U7886 (N_7886,N_7619,N_7552);
or U7887 (N_7887,N_7759,N_7772);
xor U7888 (N_7888,N_7566,N_7557);
xnor U7889 (N_7889,N_7675,N_7648);
and U7890 (N_7890,N_7758,N_7515);
xnor U7891 (N_7891,N_7606,N_7575);
nor U7892 (N_7892,N_7521,N_7565);
and U7893 (N_7893,N_7765,N_7501);
xnor U7894 (N_7894,N_7625,N_7689);
xor U7895 (N_7895,N_7600,N_7586);
and U7896 (N_7896,N_7693,N_7708);
nor U7897 (N_7897,N_7715,N_7784);
xor U7898 (N_7898,N_7714,N_7712);
and U7899 (N_7899,N_7528,N_7570);
xnor U7900 (N_7900,N_7630,N_7568);
nand U7901 (N_7901,N_7739,N_7616);
nor U7902 (N_7902,N_7594,N_7588);
nor U7903 (N_7903,N_7626,N_7577);
nand U7904 (N_7904,N_7651,N_7729);
nor U7905 (N_7905,N_7516,N_7550);
and U7906 (N_7906,N_7623,N_7698);
nand U7907 (N_7907,N_7581,N_7679);
or U7908 (N_7908,N_7666,N_7719);
nand U7909 (N_7909,N_7558,N_7695);
and U7910 (N_7910,N_7789,N_7546);
nand U7911 (N_7911,N_7709,N_7595);
and U7912 (N_7912,N_7703,N_7642);
and U7913 (N_7913,N_7769,N_7790);
or U7914 (N_7914,N_7523,N_7730);
or U7915 (N_7915,N_7634,N_7754);
nand U7916 (N_7916,N_7618,N_7771);
or U7917 (N_7917,N_7508,N_7605);
nand U7918 (N_7918,N_7553,N_7622);
and U7919 (N_7919,N_7561,N_7688);
nor U7920 (N_7920,N_7780,N_7529);
nor U7921 (N_7921,N_7778,N_7590);
nor U7922 (N_7922,N_7530,N_7507);
nor U7923 (N_7923,N_7799,N_7664);
nand U7924 (N_7924,N_7793,N_7777);
or U7925 (N_7925,N_7775,N_7536);
xnor U7926 (N_7926,N_7580,N_7624);
and U7927 (N_7927,N_7502,N_7744);
xor U7928 (N_7928,N_7753,N_7668);
and U7929 (N_7929,N_7655,N_7562);
and U7930 (N_7930,N_7669,N_7572);
or U7931 (N_7931,N_7694,N_7576);
or U7932 (N_7932,N_7509,N_7671);
and U7933 (N_7933,N_7514,N_7564);
and U7934 (N_7934,N_7583,N_7563);
or U7935 (N_7935,N_7787,N_7513);
or U7936 (N_7936,N_7656,N_7599);
nor U7937 (N_7937,N_7653,N_7537);
nand U7938 (N_7938,N_7512,N_7756);
and U7939 (N_7939,N_7681,N_7711);
nor U7940 (N_7940,N_7603,N_7762);
xnor U7941 (N_7941,N_7737,N_7761);
and U7942 (N_7942,N_7524,N_7609);
or U7943 (N_7943,N_7639,N_7652);
nor U7944 (N_7944,N_7604,N_7601);
nand U7945 (N_7945,N_7794,N_7748);
nor U7946 (N_7946,N_7613,N_7742);
or U7947 (N_7947,N_7556,N_7522);
nor U7948 (N_7948,N_7720,N_7665);
xor U7949 (N_7949,N_7672,N_7658);
nor U7950 (N_7950,N_7618,N_7796);
xnor U7951 (N_7951,N_7682,N_7646);
nor U7952 (N_7952,N_7774,N_7701);
nand U7953 (N_7953,N_7723,N_7609);
or U7954 (N_7954,N_7664,N_7618);
xnor U7955 (N_7955,N_7672,N_7629);
xor U7956 (N_7956,N_7590,N_7541);
xnor U7957 (N_7957,N_7575,N_7795);
xor U7958 (N_7958,N_7653,N_7766);
xnor U7959 (N_7959,N_7582,N_7691);
xnor U7960 (N_7960,N_7530,N_7501);
nor U7961 (N_7961,N_7520,N_7522);
and U7962 (N_7962,N_7535,N_7504);
or U7963 (N_7963,N_7742,N_7691);
nor U7964 (N_7964,N_7757,N_7585);
nor U7965 (N_7965,N_7723,N_7517);
nand U7966 (N_7966,N_7624,N_7710);
and U7967 (N_7967,N_7611,N_7720);
nand U7968 (N_7968,N_7646,N_7797);
nor U7969 (N_7969,N_7717,N_7733);
and U7970 (N_7970,N_7662,N_7565);
and U7971 (N_7971,N_7789,N_7513);
nor U7972 (N_7972,N_7690,N_7684);
or U7973 (N_7973,N_7655,N_7502);
and U7974 (N_7974,N_7531,N_7790);
or U7975 (N_7975,N_7517,N_7562);
and U7976 (N_7976,N_7742,N_7640);
or U7977 (N_7977,N_7698,N_7502);
or U7978 (N_7978,N_7640,N_7527);
nand U7979 (N_7979,N_7737,N_7609);
or U7980 (N_7980,N_7561,N_7659);
xor U7981 (N_7981,N_7666,N_7650);
nor U7982 (N_7982,N_7777,N_7553);
or U7983 (N_7983,N_7640,N_7660);
or U7984 (N_7984,N_7734,N_7798);
nand U7985 (N_7985,N_7544,N_7539);
nor U7986 (N_7986,N_7776,N_7788);
and U7987 (N_7987,N_7670,N_7775);
xnor U7988 (N_7988,N_7669,N_7710);
nand U7989 (N_7989,N_7661,N_7754);
nor U7990 (N_7990,N_7502,N_7636);
xor U7991 (N_7991,N_7651,N_7657);
and U7992 (N_7992,N_7764,N_7691);
nor U7993 (N_7993,N_7723,N_7632);
or U7994 (N_7994,N_7538,N_7534);
nand U7995 (N_7995,N_7753,N_7784);
nand U7996 (N_7996,N_7511,N_7758);
or U7997 (N_7997,N_7623,N_7743);
and U7998 (N_7998,N_7644,N_7728);
nor U7999 (N_7999,N_7539,N_7575);
or U8000 (N_8000,N_7714,N_7655);
or U8001 (N_8001,N_7739,N_7655);
xnor U8002 (N_8002,N_7743,N_7721);
or U8003 (N_8003,N_7672,N_7602);
nand U8004 (N_8004,N_7522,N_7575);
xnor U8005 (N_8005,N_7535,N_7753);
nor U8006 (N_8006,N_7566,N_7787);
and U8007 (N_8007,N_7608,N_7690);
and U8008 (N_8008,N_7613,N_7714);
nor U8009 (N_8009,N_7684,N_7744);
nor U8010 (N_8010,N_7657,N_7627);
nand U8011 (N_8011,N_7726,N_7652);
or U8012 (N_8012,N_7534,N_7643);
xnor U8013 (N_8013,N_7649,N_7784);
xor U8014 (N_8014,N_7705,N_7725);
nor U8015 (N_8015,N_7522,N_7581);
or U8016 (N_8016,N_7579,N_7575);
nor U8017 (N_8017,N_7759,N_7619);
nand U8018 (N_8018,N_7685,N_7594);
nor U8019 (N_8019,N_7745,N_7629);
xnor U8020 (N_8020,N_7602,N_7759);
or U8021 (N_8021,N_7567,N_7745);
nand U8022 (N_8022,N_7724,N_7761);
nand U8023 (N_8023,N_7601,N_7631);
or U8024 (N_8024,N_7771,N_7536);
nand U8025 (N_8025,N_7543,N_7654);
nor U8026 (N_8026,N_7761,N_7623);
and U8027 (N_8027,N_7564,N_7646);
and U8028 (N_8028,N_7778,N_7653);
xor U8029 (N_8029,N_7540,N_7672);
and U8030 (N_8030,N_7761,N_7591);
nand U8031 (N_8031,N_7690,N_7596);
xor U8032 (N_8032,N_7560,N_7512);
nor U8033 (N_8033,N_7655,N_7684);
nand U8034 (N_8034,N_7618,N_7638);
and U8035 (N_8035,N_7690,N_7751);
or U8036 (N_8036,N_7642,N_7620);
nor U8037 (N_8037,N_7629,N_7786);
nor U8038 (N_8038,N_7688,N_7697);
and U8039 (N_8039,N_7685,N_7709);
and U8040 (N_8040,N_7662,N_7670);
nand U8041 (N_8041,N_7771,N_7676);
nand U8042 (N_8042,N_7655,N_7772);
xor U8043 (N_8043,N_7781,N_7766);
nand U8044 (N_8044,N_7676,N_7511);
and U8045 (N_8045,N_7682,N_7729);
xnor U8046 (N_8046,N_7527,N_7758);
xnor U8047 (N_8047,N_7706,N_7669);
xor U8048 (N_8048,N_7655,N_7710);
and U8049 (N_8049,N_7772,N_7515);
or U8050 (N_8050,N_7629,N_7769);
and U8051 (N_8051,N_7701,N_7742);
or U8052 (N_8052,N_7602,N_7795);
nor U8053 (N_8053,N_7799,N_7695);
and U8054 (N_8054,N_7770,N_7714);
nor U8055 (N_8055,N_7518,N_7612);
nand U8056 (N_8056,N_7728,N_7731);
nand U8057 (N_8057,N_7796,N_7572);
nor U8058 (N_8058,N_7574,N_7588);
nor U8059 (N_8059,N_7634,N_7741);
nand U8060 (N_8060,N_7682,N_7696);
xnor U8061 (N_8061,N_7780,N_7732);
nor U8062 (N_8062,N_7593,N_7687);
nor U8063 (N_8063,N_7517,N_7634);
or U8064 (N_8064,N_7529,N_7525);
xnor U8065 (N_8065,N_7644,N_7523);
xnor U8066 (N_8066,N_7529,N_7794);
xnor U8067 (N_8067,N_7670,N_7754);
nand U8068 (N_8068,N_7692,N_7657);
and U8069 (N_8069,N_7702,N_7518);
nand U8070 (N_8070,N_7634,N_7559);
xor U8071 (N_8071,N_7776,N_7500);
and U8072 (N_8072,N_7731,N_7606);
nor U8073 (N_8073,N_7795,N_7637);
nand U8074 (N_8074,N_7701,N_7578);
nor U8075 (N_8075,N_7735,N_7730);
xor U8076 (N_8076,N_7649,N_7548);
and U8077 (N_8077,N_7770,N_7514);
and U8078 (N_8078,N_7532,N_7577);
or U8079 (N_8079,N_7656,N_7562);
nor U8080 (N_8080,N_7791,N_7784);
or U8081 (N_8081,N_7595,N_7682);
nor U8082 (N_8082,N_7648,N_7720);
nand U8083 (N_8083,N_7534,N_7563);
or U8084 (N_8084,N_7554,N_7725);
or U8085 (N_8085,N_7585,N_7560);
or U8086 (N_8086,N_7778,N_7697);
nand U8087 (N_8087,N_7731,N_7533);
and U8088 (N_8088,N_7556,N_7683);
and U8089 (N_8089,N_7770,N_7684);
xnor U8090 (N_8090,N_7599,N_7622);
or U8091 (N_8091,N_7650,N_7622);
xor U8092 (N_8092,N_7748,N_7738);
xor U8093 (N_8093,N_7780,N_7654);
nor U8094 (N_8094,N_7574,N_7619);
xor U8095 (N_8095,N_7673,N_7621);
xor U8096 (N_8096,N_7653,N_7546);
or U8097 (N_8097,N_7661,N_7718);
xnor U8098 (N_8098,N_7609,N_7707);
or U8099 (N_8099,N_7677,N_7772);
xor U8100 (N_8100,N_7944,N_8011);
xnor U8101 (N_8101,N_7870,N_7837);
or U8102 (N_8102,N_8072,N_8018);
or U8103 (N_8103,N_7881,N_7806);
nor U8104 (N_8104,N_8049,N_7987);
or U8105 (N_8105,N_8090,N_8084);
and U8106 (N_8106,N_8075,N_7822);
xnor U8107 (N_8107,N_7985,N_7810);
nand U8108 (N_8108,N_8060,N_8007);
nand U8109 (N_8109,N_7873,N_7983);
and U8110 (N_8110,N_7920,N_8005);
nand U8111 (N_8111,N_7808,N_7882);
xor U8112 (N_8112,N_7835,N_7804);
or U8113 (N_8113,N_7984,N_7903);
nand U8114 (N_8114,N_7824,N_7884);
xor U8115 (N_8115,N_8097,N_8088);
or U8116 (N_8116,N_8062,N_8071);
nor U8117 (N_8117,N_7931,N_7957);
xnor U8118 (N_8118,N_8030,N_7900);
or U8119 (N_8119,N_8006,N_7805);
xnor U8120 (N_8120,N_8087,N_7886);
nor U8121 (N_8121,N_7830,N_7889);
or U8122 (N_8122,N_7864,N_7818);
or U8123 (N_8123,N_7821,N_7820);
and U8124 (N_8124,N_7828,N_7840);
nand U8125 (N_8125,N_7885,N_8079);
nor U8126 (N_8126,N_7998,N_7912);
xnor U8127 (N_8127,N_7874,N_7976);
and U8128 (N_8128,N_8068,N_8048);
nor U8129 (N_8129,N_8050,N_7981);
nor U8130 (N_8130,N_7858,N_7809);
and U8131 (N_8131,N_8013,N_7817);
nor U8132 (N_8132,N_7993,N_8025);
nor U8133 (N_8133,N_8059,N_7893);
xnor U8134 (N_8134,N_7803,N_7914);
or U8135 (N_8135,N_7844,N_8029);
or U8136 (N_8136,N_7896,N_7802);
nand U8137 (N_8137,N_7898,N_7813);
or U8138 (N_8138,N_8083,N_7954);
nand U8139 (N_8139,N_7868,N_7877);
and U8140 (N_8140,N_7919,N_7849);
xor U8141 (N_8141,N_7847,N_7964);
or U8142 (N_8142,N_7816,N_7909);
or U8143 (N_8143,N_7955,N_7815);
and U8144 (N_8144,N_8016,N_7872);
and U8145 (N_8145,N_7915,N_7906);
nand U8146 (N_8146,N_8010,N_8000);
xor U8147 (N_8147,N_7926,N_7904);
xor U8148 (N_8148,N_7880,N_8033);
xnor U8149 (N_8149,N_7899,N_7859);
or U8150 (N_8150,N_7979,N_7967);
or U8151 (N_8151,N_7950,N_7867);
xor U8152 (N_8152,N_7838,N_8093);
nand U8153 (N_8153,N_7812,N_7856);
xnor U8154 (N_8154,N_8077,N_7945);
xor U8155 (N_8155,N_8015,N_8023);
nand U8156 (N_8156,N_8086,N_7959);
nand U8157 (N_8157,N_8076,N_8008);
and U8158 (N_8158,N_8066,N_7933);
nor U8159 (N_8159,N_7999,N_7911);
nor U8160 (N_8160,N_7897,N_7973);
xor U8161 (N_8161,N_8094,N_7848);
nor U8162 (N_8162,N_7961,N_7947);
xor U8163 (N_8163,N_7829,N_7879);
or U8164 (N_8164,N_7811,N_7845);
nand U8165 (N_8165,N_8026,N_8067);
nand U8166 (N_8166,N_8024,N_7928);
xor U8167 (N_8167,N_7892,N_7935);
or U8168 (N_8168,N_8092,N_8099);
and U8169 (N_8169,N_7850,N_7832);
nand U8170 (N_8170,N_7901,N_8064);
nor U8171 (N_8171,N_7855,N_7865);
nor U8172 (N_8172,N_7997,N_7823);
nor U8173 (N_8173,N_8080,N_7841);
nor U8174 (N_8174,N_7801,N_7907);
nand U8175 (N_8175,N_8085,N_7969);
or U8176 (N_8176,N_8037,N_7982);
xnor U8177 (N_8177,N_7871,N_7991);
nor U8178 (N_8178,N_7827,N_8057);
nor U8179 (N_8179,N_7965,N_7962);
xor U8180 (N_8180,N_7902,N_7953);
and U8181 (N_8181,N_7875,N_8019);
nand U8182 (N_8182,N_7905,N_7938);
nor U8183 (N_8183,N_7932,N_7857);
nor U8184 (N_8184,N_7994,N_7937);
and U8185 (N_8185,N_8002,N_7990);
xor U8186 (N_8186,N_7941,N_8082);
or U8187 (N_8187,N_8096,N_7916);
or U8188 (N_8188,N_8044,N_8004);
nand U8189 (N_8189,N_7940,N_7925);
or U8190 (N_8190,N_8021,N_7952);
and U8191 (N_8191,N_7913,N_7934);
nand U8192 (N_8192,N_7972,N_8058);
nor U8193 (N_8193,N_8031,N_7946);
xor U8194 (N_8194,N_7929,N_7863);
nor U8195 (N_8195,N_8054,N_8028);
nor U8196 (N_8196,N_7943,N_7986);
and U8197 (N_8197,N_7807,N_8051);
nand U8198 (N_8198,N_7956,N_7923);
xnor U8199 (N_8199,N_7927,N_7974);
or U8200 (N_8200,N_7989,N_7843);
xnor U8201 (N_8201,N_8039,N_7842);
xnor U8202 (N_8202,N_8065,N_8061);
and U8203 (N_8203,N_7891,N_7861);
xnor U8204 (N_8204,N_7951,N_8052);
nand U8205 (N_8205,N_7853,N_8022);
or U8206 (N_8206,N_7918,N_7939);
xnor U8207 (N_8207,N_7826,N_7825);
or U8208 (N_8208,N_7958,N_8035);
nor U8209 (N_8209,N_7917,N_7833);
nand U8210 (N_8210,N_7978,N_7948);
and U8211 (N_8211,N_8041,N_8003);
and U8212 (N_8212,N_8070,N_7834);
and U8213 (N_8213,N_7860,N_7971);
and U8214 (N_8214,N_8042,N_8098);
or U8215 (N_8215,N_7890,N_7852);
xnor U8216 (N_8216,N_7895,N_7992);
xnor U8217 (N_8217,N_7908,N_7921);
xnor U8218 (N_8218,N_8009,N_8014);
and U8219 (N_8219,N_8038,N_7894);
nand U8220 (N_8220,N_8040,N_7876);
nor U8221 (N_8221,N_7862,N_7866);
or U8222 (N_8222,N_7995,N_7966);
xnor U8223 (N_8223,N_8012,N_8081);
nor U8224 (N_8224,N_7960,N_8046);
nand U8225 (N_8225,N_8047,N_7888);
nor U8226 (N_8226,N_7977,N_8074);
and U8227 (N_8227,N_8095,N_7836);
nor U8228 (N_8228,N_8034,N_7883);
nor U8229 (N_8229,N_7851,N_8073);
nor U8230 (N_8230,N_7839,N_8045);
and U8231 (N_8231,N_7819,N_8091);
nand U8232 (N_8232,N_7968,N_7846);
nand U8233 (N_8233,N_8032,N_8053);
and U8234 (N_8234,N_7996,N_7910);
xnor U8235 (N_8235,N_8017,N_7970);
xor U8236 (N_8236,N_7800,N_7924);
nand U8237 (N_8237,N_8063,N_8055);
and U8238 (N_8238,N_7869,N_8078);
nand U8239 (N_8239,N_8027,N_7949);
or U8240 (N_8240,N_8001,N_7936);
or U8241 (N_8241,N_7942,N_8020);
or U8242 (N_8242,N_7988,N_8056);
nand U8243 (N_8243,N_7930,N_8036);
nor U8244 (N_8244,N_7922,N_8069);
xnor U8245 (N_8245,N_7963,N_7814);
xnor U8246 (N_8246,N_8089,N_8043);
xnor U8247 (N_8247,N_7854,N_7831);
and U8248 (N_8248,N_7887,N_7980);
nor U8249 (N_8249,N_7878,N_7975);
and U8250 (N_8250,N_7841,N_7824);
nand U8251 (N_8251,N_7864,N_7953);
xnor U8252 (N_8252,N_7862,N_7953);
and U8253 (N_8253,N_7913,N_7986);
nand U8254 (N_8254,N_7870,N_8017);
nor U8255 (N_8255,N_8016,N_8008);
or U8256 (N_8256,N_7850,N_7962);
nor U8257 (N_8257,N_7948,N_8043);
xnor U8258 (N_8258,N_7954,N_7807);
and U8259 (N_8259,N_8081,N_7934);
xnor U8260 (N_8260,N_7868,N_7857);
nand U8261 (N_8261,N_7912,N_8004);
xor U8262 (N_8262,N_7838,N_7832);
and U8263 (N_8263,N_7858,N_7963);
nor U8264 (N_8264,N_7935,N_7833);
or U8265 (N_8265,N_7878,N_8047);
nand U8266 (N_8266,N_8063,N_7895);
or U8267 (N_8267,N_7949,N_7846);
nor U8268 (N_8268,N_8036,N_7972);
nand U8269 (N_8269,N_7852,N_7807);
nor U8270 (N_8270,N_7909,N_7925);
nor U8271 (N_8271,N_8019,N_7833);
nor U8272 (N_8272,N_7901,N_7868);
nor U8273 (N_8273,N_7954,N_7829);
nand U8274 (N_8274,N_8089,N_7845);
and U8275 (N_8275,N_8050,N_7890);
and U8276 (N_8276,N_8045,N_8076);
nand U8277 (N_8277,N_7803,N_7804);
or U8278 (N_8278,N_7934,N_7852);
and U8279 (N_8279,N_7969,N_8092);
or U8280 (N_8280,N_7828,N_8096);
nand U8281 (N_8281,N_7832,N_8049);
or U8282 (N_8282,N_7925,N_7891);
or U8283 (N_8283,N_7810,N_7835);
nand U8284 (N_8284,N_7934,N_7896);
or U8285 (N_8285,N_8023,N_7989);
and U8286 (N_8286,N_7894,N_8099);
or U8287 (N_8287,N_7961,N_7817);
and U8288 (N_8288,N_8045,N_7807);
nor U8289 (N_8289,N_7922,N_8048);
xor U8290 (N_8290,N_7951,N_8039);
nand U8291 (N_8291,N_7996,N_8030);
and U8292 (N_8292,N_7932,N_8033);
or U8293 (N_8293,N_7844,N_7907);
xnor U8294 (N_8294,N_7947,N_8079);
nand U8295 (N_8295,N_7890,N_7923);
and U8296 (N_8296,N_7817,N_7996);
xnor U8297 (N_8297,N_8003,N_8077);
or U8298 (N_8298,N_7917,N_7895);
or U8299 (N_8299,N_7904,N_8045);
or U8300 (N_8300,N_7825,N_8080);
or U8301 (N_8301,N_7828,N_7802);
nand U8302 (N_8302,N_7871,N_7878);
or U8303 (N_8303,N_8017,N_8043);
and U8304 (N_8304,N_8059,N_7805);
nor U8305 (N_8305,N_7962,N_8065);
or U8306 (N_8306,N_7912,N_7890);
nor U8307 (N_8307,N_7849,N_7974);
nor U8308 (N_8308,N_7881,N_7927);
xor U8309 (N_8309,N_8001,N_8056);
nor U8310 (N_8310,N_8083,N_8032);
or U8311 (N_8311,N_7810,N_8010);
nand U8312 (N_8312,N_7978,N_8022);
nand U8313 (N_8313,N_8063,N_7879);
nor U8314 (N_8314,N_7894,N_7943);
or U8315 (N_8315,N_8028,N_7918);
and U8316 (N_8316,N_7921,N_7984);
or U8317 (N_8317,N_7968,N_7808);
xor U8318 (N_8318,N_7817,N_7946);
or U8319 (N_8319,N_7826,N_8025);
or U8320 (N_8320,N_7913,N_7961);
and U8321 (N_8321,N_8013,N_7800);
or U8322 (N_8322,N_7854,N_8062);
nor U8323 (N_8323,N_7914,N_7965);
nor U8324 (N_8324,N_8097,N_8094);
nor U8325 (N_8325,N_8022,N_8037);
xor U8326 (N_8326,N_7890,N_7946);
nor U8327 (N_8327,N_7850,N_8086);
nor U8328 (N_8328,N_7932,N_7920);
nor U8329 (N_8329,N_8044,N_8026);
nand U8330 (N_8330,N_7817,N_8068);
xor U8331 (N_8331,N_7923,N_7876);
xnor U8332 (N_8332,N_7801,N_7832);
and U8333 (N_8333,N_7823,N_7841);
xor U8334 (N_8334,N_7995,N_8022);
or U8335 (N_8335,N_7830,N_7871);
xor U8336 (N_8336,N_7922,N_7976);
and U8337 (N_8337,N_7938,N_8025);
nand U8338 (N_8338,N_7917,N_8024);
nand U8339 (N_8339,N_7907,N_8040);
or U8340 (N_8340,N_8033,N_8022);
xnor U8341 (N_8341,N_7902,N_7912);
and U8342 (N_8342,N_7809,N_7965);
and U8343 (N_8343,N_8094,N_7925);
or U8344 (N_8344,N_7811,N_7945);
or U8345 (N_8345,N_8087,N_7973);
and U8346 (N_8346,N_7986,N_7857);
and U8347 (N_8347,N_7899,N_7969);
nor U8348 (N_8348,N_7896,N_8093);
or U8349 (N_8349,N_8000,N_7992);
or U8350 (N_8350,N_7982,N_7852);
xnor U8351 (N_8351,N_8002,N_8027);
xor U8352 (N_8352,N_7972,N_8025);
nor U8353 (N_8353,N_7869,N_7917);
xnor U8354 (N_8354,N_7991,N_7866);
xor U8355 (N_8355,N_7816,N_7967);
or U8356 (N_8356,N_7917,N_8085);
or U8357 (N_8357,N_8023,N_7834);
or U8358 (N_8358,N_7874,N_7912);
nor U8359 (N_8359,N_7941,N_7949);
nand U8360 (N_8360,N_7830,N_7821);
or U8361 (N_8361,N_7888,N_7991);
nor U8362 (N_8362,N_7862,N_7979);
or U8363 (N_8363,N_8084,N_7845);
or U8364 (N_8364,N_8095,N_7923);
nand U8365 (N_8365,N_7836,N_7986);
and U8366 (N_8366,N_8020,N_7932);
or U8367 (N_8367,N_7851,N_7846);
xnor U8368 (N_8368,N_7805,N_7994);
nor U8369 (N_8369,N_7809,N_7866);
and U8370 (N_8370,N_8006,N_8054);
nand U8371 (N_8371,N_7920,N_7853);
and U8372 (N_8372,N_7948,N_8029);
nand U8373 (N_8373,N_7860,N_7924);
nand U8374 (N_8374,N_7953,N_7997);
nor U8375 (N_8375,N_7914,N_7931);
nor U8376 (N_8376,N_7851,N_7861);
xor U8377 (N_8377,N_7900,N_7911);
or U8378 (N_8378,N_7877,N_8084);
nand U8379 (N_8379,N_8072,N_7912);
and U8380 (N_8380,N_7902,N_7994);
xnor U8381 (N_8381,N_7986,N_7997);
xnor U8382 (N_8382,N_7886,N_7850);
nor U8383 (N_8383,N_8052,N_7901);
or U8384 (N_8384,N_8061,N_8027);
xnor U8385 (N_8385,N_7825,N_7809);
and U8386 (N_8386,N_7963,N_8090);
nand U8387 (N_8387,N_7969,N_8075);
or U8388 (N_8388,N_7954,N_7865);
xnor U8389 (N_8389,N_7803,N_7902);
xor U8390 (N_8390,N_7985,N_8061);
xnor U8391 (N_8391,N_8016,N_7853);
or U8392 (N_8392,N_7991,N_8088);
or U8393 (N_8393,N_7988,N_7841);
nand U8394 (N_8394,N_7811,N_7881);
and U8395 (N_8395,N_8079,N_8050);
and U8396 (N_8396,N_7867,N_8074);
and U8397 (N_8397,N_8027,N_8080);
nand U8398 (N_8398,N_7814,N_7813);
nand U8399 (N_8399,N_8086,N_8055);
xor U8400 (N_8400,N_8309,N_8239);
nand U8401 (N_8401,N_8285,N_8263);
nand U8402 (N_8402,N_8382,N_8190);
nor U8403 (N_8403,N_8158,N_8219);
xor U8404 (N_8404,N_8213,N_8262);
xnor U8405 (N_8405,N_8305,N_8299);
nor U8406 (N_8406,N_8124,N_8232);
nand U8407 (N_8407,N_8274,N_8137);
nor U8408 (N_8408,N_8173,N_8356);
xnor U8409 (N_8409,N_8115,N_8107);
nor U8410 (N_8410,N_8128,N_8399);
or U8411 (N_8411,N_8187,N_8183);
or U8412 (N_8412,N_8130,N_8393);
nor U8413 (N_8413,N_8249,N_8243);
or U8414 (N_8414,N_8209,N_8182);
and U8415 (N_8415,N_8138,N_8149);
nor U8416 (N_8416,N_8254,N_8376);
nand U8417 (N_8417,N_8160,N_8385);
nor U8418 (N_8418,N_8155,N_8349);
xor U8419 (N_8419,N_8324,N_8195);
nand U8420 (N_8420,N_8114,N_8224);
nand U8421 (N_8421,N_8169,N_8250);
nand U8422 (N_8422,N_8180,N_8353);
and U8423 (N_8423,N_8153,N_8246);
nor U8424 (N_8424,N_8216,N_8211);
nand U8425 (N_8425,N_8364,N_8105);
or U8426 (N_8426,N_8301,N_8384);
and U8427 (N_8427,N_8116,N_8127);
xor U8428 (N_8428,N_8375,N_8390);
or U8429 (N_8429,N_8231,N_8192);
nand U8430 (N_8430,N_8238,N_8135);
and U8431 (N_8431,N_8302,N_8331);
and U8432 (N_8432,N_8295,N_8369);
xor U8433 (N_8433,N_8165,N_8259);
nand U8434 (N_8434,N_8111,N_8251);
and U8435 (N_8435,N_8199,N_8379);
or U8436 (N_8436,N_8320,N_8206);
or U8437 (N_8437,N_8342,N_8288);
nand U8438 (N_8438,N_8335,N_8276);
and U8439 (N_8439,N_8119,N_8215);
xor U8440 (N_8440,N_8314,N_8362);
xnor U8441 (N_8441,N_8102,N_8151);
and U8442 (N_8442,N_8359,N_8355);
and U8443 (N_8443,N_8277,N_8374);
xnor U8444 (N_8444,N_8291,N_8395);
or U8445 (N_8445,N_8245,N_8172);
nand U8446 (N_8446,N_8132,N_8330);
or U8447 (N_8447,N_8336,N_8147);
and U8448 (N_8448,N_8131,N_8354);
or U8449 (N_8449,N_8212,N_8150);
or U8450 (N_8450,N_8252,N_8159);
nor U8451 (N_8451,N_8337,N_8312);
and U8452 (N_8452,N_8348,N_8284);
and U8453 (N_8453,N_8134,N_8176);
nor U8454 (N_8454,N_8358,N_8207);
nand U8455 (N_8455,N_8329,N_8113);
nand U8456 (N_8456,N_8126,N_8256);
and U8457 (N_8457,N_8104,N_8185);
or U8458 (N_8458,N_8201,N_8241);
or U8459 (N_8459,N_8363,N_8394);
nor U8460 (N_8460,N_8319,N_8117);
xnor U8461 (N_8461,N_8257,N_8196);
nor U8462 (N_8462,N_8283,N_8178);
and U8463 (N_8463,N_8272,N_8136);
or U8464 (N_8464,N_8214,N_8332);
xnor U8465 (N_8465,N_8168,N_8267);
nor U8466 (N_8466,N_8208,N_8123);
nand U8467 (N_8467,N_8248,N_8120);
nor U8468 (N_8468,N_8181,N_8139);
or U8469 (N_8469,N_8204,N_8109);
nor U8470 (N_8470,N_8265,N_8308);
and U8471 (N_8471,N_8161,N_8121);
nor U8472 (N_8472,N_8280,N_8273);
xor U8473 (N_8473,N_8298,N_8372);
nor U8474 (N_8474,N_8247,N_8327);
or U8475 (N_8475,N_8236,N_8202);
and U8476 (N_8476,N_8322,N_8148);
nor U8477 (N_8477,N_8380,N_8118);
nor U8478 (N_8478,N_8240,N_8106);
and U8479 (N_8479,N_8189,N_8221);
and U8480 (N_8480,N_8296,N_8396);
nand U8481 (N_8481,N_8141,N_8333);
nand U8482 (N_8482,N_8170,N_8205);
or U8483 (N_8483,N_8290,N_8347);
xnor U8484 (N_8484,N_8163,N_8318);
or U8485 (N_8485,N_8268,N_8100);
nand U8486 (N_8486,N_8389,N_8122);
nand U8487 (N_8487,N_8264,N_8146);
and U8488 (N_8488,N_8388,N_8334);
nand U8489 (N_8489,N_8310,N_8186);
xor U8490 (N_8490,N_8378,N_8269);
nor U8491 (N_8491,N_8386,N_8317);
nor U8492 (N_8492,N_8152,N_8357);
xor U8493 (N_8493,N_8345,N_8222);
nor U8494 (N_8494,N_8144,N_8179);
nor U8495 (N_8495,N_8328,N_8242);
nand U8496 (N_8496,N_8392,N_8343);
or U8497 (N_8497,N_8368,N_8171);
and U8498 (N_8498,N_8286,N_8223);
and U8499 (N_8499,N_8381,N_8191);
or U8500 (N_8500,N_8233,N_8391);
and U8501 (N_8501,N_8217,N_8321);
xnor U8502 (N_8502,N_8129,N_8143);
and U8503 (N_8503,N_8300,N_8346);
and U8504 (N_8504,N_8145,N_8307);
and U8505 (N_8505,N_8140,N_8387);
and U8506 (N_8506,N_8255,N_8377);
nand U8507 (N_8507,N_8383,N_8325);
nor U8508 (N_8508,N_8156,N_8167);
and U8509 (N_8509,N_8157,N_8184);
nor U8510 (N_8510,N_8175,N_8101);
and U8511 (N_8511,N_8271,N_8174);
or U8512 (N_8512,N_8360,N_8287);
nor U8513 (N_8513,N_8194,N_8133);
nor U8514 (N_8514,N_8293,N_8266);
and U8515 (N_8515,N_8125,N_8193);
xnor U8516 (N_8516,N_8398,N_8260);
nor U8517 (N_8517,N_8397,N_8370);
or U8518 (N_8518,N_8311,N_8229);
nand U8519 (N_8519,N_8218,N_8371);
or U8520 (N_8520,N_8292,N_8281);
and U8521 (N_8521,N_8315,N_8112);
nand U8522 (N_8522,N_8198,N_8282);
nand U8523 (N_8523,N_8365,N_8244);
nor U8524 (N_8524,N_8313,N_8297);
or U8525 (N_8525,N_8338,N_8270);
and U8526 (N_8526,N_8234,N_8154);
nand U8527 (N_8527,N_8225,N_8279);
xnor U8528 (N_8528,N_8230,N_8188);
xor U8529 (N_8529,N_8237,N_8366);
nor U8530 (N_8530,N_8367,N_8323);
nor U8531 (N_8531,N_8350,N_8352);
xnor U8532 (N_8532,N_8197,N_8316);
nor U8533 (N_8533,N_8226,N_8164);
and U8534 (N_8534,N_8304,N_8294);
nor U8535 (N_8535,N_8108,N_8228);
xor U8536 (N_8536,N_8339,N_8289);
nor U8537 (N_8537,N_8162,N_8340);
nor U8538 (N_8538,N_8142,N_8275);
nor U8539 (N_8539,N_8103,N_8373);
or U8540 (N_8540,N_8258,N_8166);
nor U8541 (N_8541,N_8351,N_8344);
xor U8542 (N_8542,N_8227,N_8326);
nor U8543 (N_8543,N_8235,N_8203);
nand U8544 (N_8544,N_8341,N_8253);
nand U8545 (N_8545,N_8210,N_8220);
nor U8546 (N_8546,N_8278,N_8303);
nand U8547 (N_8547,N_8177,N_8261);
nand U8548 (N_8548,N_8306,N_8200);
xnor U8549 (N_8549,N_8361,N_8110);
nand U8550 (N_8550,N_8183,N_8281);
nand U8551 (N_8551,N_8234,N_8111);
xor U8552 (N_8552,N_8241,N_8384);
and U8553 (N_8553,N_8341,N_8205);
xor U8554 (N_8554,N_8233,N_8357);
or U8555 (N_8555,N_8230,N_8379);
xor U8556 (N_8556,N_8294,N_8356);
nand U8557 (N_8557,N_8355,N_8227);
xor U8558 (N_8558,N_8148,N_8214);
or U8559 (N_8559,N_8207,N_8242);
nor U8560 (N_8560,N_8355,N_8387);
or U8561 (N_8561,N_8187,N_8303);
or U8562 (N_8562,N_8274,N_8324);
and U8563 (N_8563,N_8143,N_8398);
or U8564 (N_8564,N_8311,N_8312);
and U8565 (N_8565,N_8326,N_8235);
or U8566 (N_8566,N_8380,N_8333);
and U8567 (N_8567,N_8161,N_8318);
xnor U8568 (N_8568,N_8140,N_8337);
and U8569 (N_8569,N_8300,N_8116);
and U8570 (N_8570,N_8182,N_8233);
nand U8571 (N_8571,N_8153,N_8282);
nor U8572 (N_8572,N_8228,N_8250);
nand U8573 (N_8573,N_8260,N_8105);
nor U8574 (N_8574,N_8225,N_8121);
nor U8575 (N_8575,N_8190,N_8257);
xor U8576 (N_8576,N_8386,N_8342);
xor U8577 (N_8577,N_8156,N_8187);
and U8578 (N_8578,N_8287,N_8168);
xor U8579 (N_8579,N_8235,N_8337);
and U8580 (N_8580,N_8269,N_8188);
and U8581 (N_8581,N_8275,N_8239);
xnor U8582 (N_8582,N_8348,N_8299);
xor U8583 (N_8583,N_8152,N_8265);
nand U8584 (N_8584,N_8199,N_8351);
or U8585 (N_8585,N_8229,N_8216);
or U8586 (N_8586,N_8172,N_8273);
nor U8587 (N_8587,N_8385,N_8278);
and U8588 (N_8588,N_8306,N_8271);
nand U8589 (N_8589,N_8347,N_8214);
or U8590 (N_8590,N_8204,N_8115);
xor U8591 (N_8591,N_8125,N_8247);
nor U8592 (N_8592,N_8176,N_8169);
and U8593 (N_8593,N_8335,N_8386);
and U8594 (N_8594,N_8314,N_8208);
or U8595 (N_8595,N_8202,N_8390);
nor U8596 (N_8596,N_8364,N_8270);
and U8597 (N_8597,N_8394,N_8316);
and U8598 (N_8598,N_8183,N_8128);
nor U8599 (N_8599,N_8137,N_8302);
nand U8600 (N_8600,N_8373,N_8214);
nor U8601 (N_8601,N_8299,N_8111);
xor U8602 (N_8602,N_8198,N_8371);
and U8603 (N_8603,N_8192,N_8311);
or U8604 (N_8604,N_8254,N_8302);
or U8605 (N_8605,N_8321,N_8203);
nor U8606 (N_8606,N_8137,N_8193);
and U8607 (N_8607,N_8186,N_8136);
nor U8608 (N_8608,N_8361,N_8148);
xnor U8609 (N_8609,N_8337,N_8289);
and U8610 (N_8610,N_8388,N_8196);
or U8611 (N_8611,N_8241,N_8221);
xor U8612 (N_8612,N_8234,N_8281);
xor U8613 (N_8613,N_8301,N_8186);
xnor U8614 (N_8614,N_8130,N_8337);
or U8615 (N_8615,N_8175,N_8388);
xor U8616 (N_8616,N_8373,N_8126);
xnor U8617 (N_8617,N_8369,N_8116);
xnor U8618 (N_8618,N_8213,N_8190);
nand U8619 (N_8619,N_8352,N_8314);
and U8620 (N_8620,N_8347,N_8212);
or U8621 (N_8621,N_8367,N_8210);
or U8622 (N_8622,N_8322,N_8138);
xnor U8623 (N_8623,N_8173,N_8153);
xnor U8624 (N_8624,N_8217,N_8361);
xor U8625 (N_8625,N_8399,N_8284);
nor U8626 (N_8626,N_8226,N_8220);
xnor U8627 (N_8627,N_8391,N_8195);
and U8628 (N_8628,N_8350,N_8392);
nand U8629 (N_8629,N_8356,N_8378);
and U8630 (N_8630,N_8186,N_8278);
nand U8631 (N_8631,N_8310,N_8295);
xnor U8632 (N_8632,N_8148,N_8334);
nand U8633 (N_8633,N_8313,N_8364);
or U8634 (N_8634,N_8381,N_8170);
nand U8635 (N_8635,N_8115,N_8232);
xnor U8636 (N_8636,N_8271,N_8260);
and U8637 (N_8637,N_8324,N_8247);
nor U8638 (N_8638,N_8116,N_8303);
nand U8639 (N_8639,N_8268,N_8204);
xnor U8640 (N_8640,N_8269,N_8218);
xnor U8641 (N_8641,N_8228,N_8196);
xor U8642 (N_8642,N_8392,N_8333);
and U8643 (N_8643,N_8120,N_8294);
or U8644 (N_8644,N_8271,N_8340);
nand U8645 (N_8645,N_8207,N_8213);
or U8646 (N_8646,N_8312,N_8350);
nand U8647 (N_8647,N_8323,N_8241);
or U8648 (N_8648,N_8234,N_8187);
or U8649 (N_8649,N_8137,N_8271);
xor U8650 (N_8650,N_8120,N_8136);
and U8651 (N_8651,N_8234,N_8325);
and U8652 (N_8652,N_8118,N_8162);
nand U8653 (N_8653,N_8212,N_8256);
nor U8654 (N_8654,N_8277,N_8380);
xnor U8655 (N_8655,N_8283,N_8107);
nand U8656 (N_8656,N_8126,N_8370);
and U8657 (N_8657,N_8370,N_8161);
xnor U8658 (N_8658,N_8286,N_8179);
nor U8659 (N_8659,N_8182,N_8169);
or U8660 (N_8660,N_8200,N_8242);
nor U8661 (N_8661,N_8376,N_8141);
nand U8662 (N_8662,N_8280,N_8155);
nor U8663 (N_8663,N_8275,N_8247);
nor U8664 (N_8664,N_8130,N_8258);
xnor U8665 (N_8665,N_8241,N_8249);
xor U8666 (N_8666,N_8261,N_8191);
nor U8667 (N_8667,N_8200,N_8175);
and U8668 (N_8668,N_8111,N_8138);
nor U8669 (N_8669,N_8281,N_8195);
and U8670 (N_8670,N_8305,N_8221);
nand U8671 (N_8671,N_8346,N_8268);
or U8672 (N_8672,N_8105,N_8295);
xor U8673 (N_8673,N_8268,N_8202);
or U8674 (N_8674,N_8327,N_8282);
xor U8675 (N_8675,N_8105,N_8285);
or U8676 (N_8676,N_8380,N_8334);
and U8677 (N_8677,N_8205,N_8316);
or U8678 (N_8678,N_8338,N_8128);
nor U8679 (N_8679,N_8275,N_8189);
or U8680 (N_8680,N_8211,N_8150);
nand U8681 (N_8681,N_8290,N_8362);
and U8682 (N_8682,N_8238,N_8242);
and U8683 (N_8683,N_8376,N_8103);
nor U8684 (N_8684,N_8398,N_8106);
xor U8685 (N_8685,N_8291,N_8360);
and U8686 (N_8686,N_8332,N_8102);
nand U8687 (N_8687,N_8341,N_8325);
nor U8688 (N_8688,N_8258,N_8136);
or U8689 (N_8689,N_8314,N_8234);
nor U8690 (N_8690,N_8283,N_8248);
or U8691 (N_8691,N_8338,N_8181);
nand U8692 (N_8692,N_8170,N_8317);
or U8693 (N_8693,N_8395,N_8234);
nor U8694 (N_8694,N_8189,N_8280);
nor U8695 (N_8695,N_8169,N_8312);
nor U8696 (N_8696,N_8184,N_8210);
and U8697 (N_8697,N_8388,N_8351);
and U8698 (N_8698,N_8356,N_8228);
xnor U8699 (N_8699,N_8367,N_8318);
or U8700 (N_8700,N_8538,N_8453);
nand U8701 (N_8701,N_8498,N_8560);
and U8702 (N_8702,N_8524,N_8545);
or U8703 (N_8703,N_8685,N_8463);
and U8704 (N_8704,N_8662,N_8684);
nand U8705 (N_8705,N_8481,N_8629);
or U8706 (N_8706,N_8586,N_8536);
nor U8707 (N_8707,N_8477,N_8413);
xor U8708 (N_8708,N_8680,N_8509);
nor U8709 (N_8709,N_8480,N_8525);
and U8710 (N_8710,N_8559,N_8646);
nor U8711 (N_8711,N_8659,N_8403);
nor U8712 (N_8712,N_8492,N_8683);
nor U8713 (N_8713,N_8572,N_8682);
nand U8714 (N_8714,N_8535,N_8404);
nor U8715 (N_8715,N_8464,N_8618);
nor U8716 (N_8716,N_8690,N_8512);
and U8717 (N_8717,N_8416,N_8454);
or U8718 (N_8718,N_8444,N_8625);
nand U8719 (N_8719,N_8656,N_8518);
xnor U8720 (N_8720,N_8402,N_8531);
or U8721 (N_8721,N_8540,N_8555);
nand U8722 (N_8722,N_8451,N_8654);
or U8723 (N_8723,N_8636,N_8408);
or U8724 (N_8724,N_8634,N_8537);
and U8725 (N_8725,N_8466,N_8697);
nand U8726 (N_8726,N_8585,N_8595);
nor U8727 (N_8727,N_8426,N_8400);
and U8728 (N_8728,N_8615,N_8551);
nor U8729 (N_8729,N_8489,N_8670);
or U8730 (N_8730,N_8457,N_8485);
nand U8731 (N_8731,N_8621,N_8446);
nand U8732 (N_8732,N_8648,N_8599);
or U8733 (N_8733,N_8476,N_8475);
or U8734 (N_8734,N_8434,N_8582);
nor U8735 (N_8735,N_8503,N_8414);
nand U8736 (N_8736,N_8563,N_8669);
xor U8737 (N_8737,N_8554,N_8473);
nand U8738 (N_8738,N_8678,N_8442);
xor U8739 (N_8739,N_8443,N_8433);
nand U8740 (N_8740,N_8578,N_8513);
xnor U8741 (N_8741,N_8439,N_8411);
nor U8742 (N_8742,N_8462,N_8437);
and U8743 (N_8743,N_8514,N_8627);
xnor U8744 (N_8744,N_8677,N_8543);
nand U8745 (N_8745,N_8651,N_8587);
or U8746 (N_8746,N_8626,N_8583);
xor U8747 (N_8747,N_8522,N_8542);
or U8748 (N_8748,N_8461,N_8552);
nor U8749 (N_8749,N_8455,N_8588);
or U8750 (N_8750,N_8440,N_8698);
xor U8751 (N_8751,N_8521,N_8650);
or U8752 (N_8752,N_8569,N_8630);
xor U8753 (N_8753,N_8639,N_8649);
nand U8754 (N_8754,N_8527,N_8609);
nand U8755 (N_8755,N_8628,N_8465);
nand U8756 (N_8756,N_8484,N_8501);
xnor U8757 (N_8757,N_8529,N_8544);
nor U8758 (N_8758,N_8577,N_8691);
xnor U8759 (N_8759,N_8499,N_8622);
xor U8760 (N_8760,N_8600,N_8488);
or U8761 (N_8761,N_8592,N_8547);
nor U8762 (N_8762,N_8570,N_8665);
nor U8763 (N_8763,N_8546,N_8415);
nor U8764 (N_8764,N_8637,N_8574);
and U8765 (N_8765,N_8493,N_8612);
or U8766 (N_8766,N_8458,N_8644);
and U8767 (N_8767,N_8422,N_8590);
nor U8768 (N_8768,N_8419,N_8568);
nand U8769 (N_8769,N_8429,N_8689);
and U8770 (N_8770,N_8505,N_8658);
and U8771 (N_8771,N_8679,N_8591);
nand U8772 (N_8772,N_8675,N_8616);
nor U8773 (N_8773,N_8407,N_8566);
nand U8774 (N_8774,N_8624,N_8441);
or U8775 (N_8775,N_8594,N_8483);
or U8776 (N_8776,N_8655,N_8478);
or U8777 (N_8777,N_8657,N_8681);
nor U8778 (N_8778,N_8479,N_8496);
and U8779 (N_8779,N_8694,N_8645);
nor U8780 (N_8780,N_8515,N_8597);
nand U8781 (N_8781,N_8581,N_8530);
nor U8782 (N_8782,N_8605,N_8652);
nand U8783 (N_8783,N_8550,N_8516);
and U8784 (N_8784,N_8526,N_8553);
and U8785 (N_8785,N_8664,N_8663);
or U8786 (N_8786,N_8528,N_8614);
and U8787 (N_8787,N_8427,N_8459);
nor U8788 (N_8788,N_8425,N_8508);
nor U8789 (N_8789,N_8676,N_8549);
xor U8790 (N_8790,N_8610,N_8580);
and U8791 (N_8791,N_8673,N_8565);
nand U8792 (N_8792,N_8506,N_8640);
or U8793 (N_8793,N_8661,N_8567);
nand U8794 (N_8794,N_8533,N_8438);
nor U8795 (N_8795,N_8623,N_8604);
and U8796 (N_8796,N_8602,N_8532);
nor U8797 (N_8797,N_8510,N_8534);
or U8798 (N_8798,N_8452,N_8500);
nor U8799 (N_8799,N_8695,N_8406);
nor U8800 (N_8800,N_8671,N_8643);
and U8801 (N_8801,N_8424,N_8571);
xnor U8802 (N_8802,N_8539,N_8467);
xnor U8803 (N_8803,N_8519,N_8558);
xor U8804 (N_8804,N_8601,N_8660);
or U8805 (N_8805,N_8672,N_8638);
and U8806 (N_8806,N_8409,N_8504);
or U8807 (N_8807,N_8561,N_8596);
or U8808 (N_8808,N_8472,N_8410);
and U8809 (N_8809,N_8611,N_8431);
or U8810 (N_8810,N_8632,N_8447);
or U8811 (N_8811,N_8573,N_8647);
nor U8812 (N_8812,N_8693,N_8456);
nor U8813 (N_8813,N_8562,N_8448);
nor U8814 (N_8814,N_8607,N_8470);
nand U8815 (N_8815,N_8468,N_8486);
xnor U8816 (N_8816,N_8631,N_8471);
or U8817 (N_8817,N_8418,N_8401);
or U8818 (N_8818,N_8564,N_8502);
and U8819 (N_8819,N_8541,N_8432);
nand U8820 (N_8820,N_8491,N_8507);
nor U8821 (N_8821,N_8603,N_8474);
nand U8822 (N_8822,N_8653,N_8460);
and U8823 (N_8823,N_8633,N_8635);
and U8824 (N_8824,N_8688,N_8405);
xnor U8825 (N_8825,N_8641,N_8613);
nor U8826 (N_8826,N_8469,N_8619);
nand U8827 (N_8827,N_8482,N_8517);
nand U8828 (N_8828,N_8450,N_8696);
xnor U8829 (N_8829,N_8449,N_8548);
xor U8830 (N_8830,N_8589,N_8497);
or U8831 (N_8831,N_8620,N_8692);
or U8832 (N_8832,N_8428,N_8576);
xnor U8833 (N_8833,N_8436,N_8699);
nand U8834 (N_8834,N_8593,N_8511);
nand U8835 (N_8835,N_8494,N_8490);
xor U8836 (N_8836,N_8487,N_8417);
nand U8837 (N_8837,N_8445,N_8421);
nand U8838 (N_8838,N_8520,N_8642);
and U8839 (N_8839,N_8423,N_8523);
nand U8840 (N_8840,N_8608,N_8606);
and U8841 (N_8841,N_8495,N_8556);
and U8842 (N_8842,N_8579,N_8584);
nand U8843 (N_8843,N_8420,N_8430);
nor U8844 (N_8844,N_8674,N_8667);
or U8845 (N_8845,N_8598,N_8686);
or U8846 (N_8846,N_8435,N_8617);
nand U8847 (N_8847,N_8687,N_8668);
and U8848 (N_8848,N_8666,N_8557);
nand U8849 (N_8849,N_8412,N_8575);
nor U8850 (N_8850,N_8510,N_8417);
xnor U8851 (N_8851,N_8487,N_8653);
nor U8852 (N_8852,N_8609,N_8590);
xnor U8853 (N_8853,N_8464,N_8615);
nand U8854 (N_8854,N_8691,N_8563);
and U8855 (N_8855,N_8684,N_8490);
or U8856 (N_8856,N_8515,N_8485);
or U8857 (N_8857,N_8567,N_8656);
xor U8858 (N_8858,N_8679,N_8464);
nor U8859 (N_8859,N_8678,N_8434);
or U8860 (N_8860,N_8551,N_8666);
nand U8861 (N_8861,N_8605,N_8623);
or U8862 (N_8862,N_8468,N_8674);
nand U8863 (N_8863,N_8570,N_8523);
or U8864 (N_8864,N_8466,N_8508);
xor U8865 (N_8865,N_8639,N_8442);
and U8866 (N_8866,N_8633,N_8550);
nand U8867 (N_8867,N_8519,N_8642);
nand U8868 (N_8868,N_8566,N_8670);
nand U8869 (N_8869,N_8635,N_8574);
nand U8870 (N_8870,N_8575,N_8665);
nor U8871 (N_8871,N_8628,N_8621);
nand U8872 (N_8872,N_8574,N_8504);
xnor U8873 (N_8873,N_8582,N_8685);
and U8874 (N_8874,N_8505,N_8563);
xnor U8875 (N_8875,N_8671,N_8667);
or U8876 (N_8876,N_8675,N_8425);
and U8877 (N_8877,N_8521,N_8553);
and U8878 (N_8878,N_8610,N_8607);
nor U8879 (N_8879,N_8442,N_8575);
or U8880 (N_8880,N_8426,N_8689);
xnor U8881 (N_8881,N_8581,N_8562);
or U8882 (N_8882,N_8404,N_8580);
nor U8883 (N_8883,N_8633,N_8517);
and U8884 (N_8884,N_8542,N_8426);
or U8885 (N_8885,N_8657,N_8687);
nor U8886 (N_8886,N_8646,N_8400);
nor U8887 (N_8887,N_8673,N_8511);
or U8888 (N_8888,N_8681,N_8417);
nor U8889 (N_8889,N_8674,N_8519);
and U8890 (N_8890,N_8413,N_8513);
and U8891 (N_8891,N_8492,N_8692);
or U8892 (N_8892,N_8482,N_8586);
nand U8893 (N_8893,N_8636,N_8686);
nor U8894 (N_8894,N_8687,N_8551);
nand U8895 (N_8895,N_8463,N_8494);
nand U8896 (N_8896,N_8459,N_8460);
nor U8897 (N_8897,N_8655,N_8641);
or U8898 (N_8898,N_8631,N_8675);
or U8899 (N_8899,N_8534,N_8446);
and U8900 (N_8900,N_8639,N_8682);
or U8901 (N_8901,N_8663,N_8694);
nor U8902 (N_8902,N_8653,N_8637);
or U8903 (N_8903,N_8447,N_8548);
or U8904 (N_8904,N_8640,N_8624);
nor U8905 (N_8905,N_8509,N_8419);
and U8906 (N_8906,N_8465,N_8582);
xor U8907 (N_8907,N_8544,N_8698);
nor U8908 (N_8908,N_8600,N_8647);
and U8909 (N_8909,N_8424,N_8525);
nand U8910 (N_8910,N_8415,N_8667);
nand U8911 (N_8911,N_8674,N_8434);
nor U8912 (N_8912,N_8517,N_8473);
nor U8913 (N_8913,N_8444,N_8650);
or U8914 (N_8914,N_8417,N_8460);
xor U8915 (N_8915,N_8654,N_8525);
and U8916 (N_8916,N_8453,N_8654);
nand U8917 (N_8917,N_8423,N_8667);
and U8918 (N_8918,N_8425,N_8529);
or U8919 (N_8919,N_8412,N_8646);
and U8920 (N_8920,N_8506,N_8450);
nor U8921 (N_8921,N_8546,N_8447);
nand U8922 (N_8922,N_8677,N_8438);
and U8923 (N_8923,N_8699,N_8693);
xor U8924 (N_8924,N_8452,N_8633);
and U8925 (N_8925,N_8696,N_8589);
nor U8926 (N_8926,N_8440,N_8676);
nand U8927 (N_8927,N_8631,N_8661);
and U8928 (N_8928,N_8513,N_8687);
nand U8929 (N_8929,N_8687,N_8522);
nand U8930 (N_8930,N_8585,N_8651);
nor U8931 (N_8931,N_8562,N_8531);
or U8932 (N_8932,N_8536,N_8462);
and U8933 (N_8933,N_8496,N_8409);
nand U8934 (N_8934,N_8588,N_8526);
xnor U8935 (N_8935,N_8651,N_8411);
xor U8936 (N_8936,N_8439,N_8595);
and U8937 (N_8937,N_8676,N_8592);
nor U8938 (N_8938,N_8665,N_8638);
and U8939 (N_8939,N_8564,N_8568);
nor U8940 (N_8940,N_8530,N_8623);
nand U8941 (N_8941,N_8466,N_8507);
nor U8942 (N_8942,N_8416,N_8677);
and U8943 (N_8943,N_8571,N_8555);
xnor U8944 (N_8944,N_8601,N_8409);
xnor U8945 (N_8945,N_8529,N_8466);
and U8946 (N_8946,N_8408,N_8454);
and U8947 (N_8947,N_8407,N_8571);
and U8948 (N_8948,N_8666,N_8643);
and U8949 (N_8949,N_8482,N_8435);
xnor U8950 (N_8950,N_8487,N_8631);
nand U8951 (N_8951,N_8586,N_8403);
and U8952 (N_8952,N_8614,N_8669);
and U8953 (N_8953,N_8495,N_8493);
nand U8954 (N_8954,N_8615,N_8675);
and U8955 (N_8955,N_8614,N_8695);
or U8956 (N_8956,N_8539,N_8444);
nor U8957 (N_8957,N_8503,N_8516);
nor U8958 (N_8958,N_8542,N_8483);
nand U8959 (N_8959,N_8610,N_8406);
nor U8960 (N_8960,N_8658,N_8656);
nand U8961 (N_8961,N_8454,N_8440);
nand U8962 (N_8962,N_8453,N_8695);
nand U8963 (N_8963,N_8476,N_8570);
or U8964 (N_8964,N_8560,N_8668);
xnor U8965 (N_8965,N_8673,N_8629);
xor U8966 (N_8966,N_8414,N_8537);
nand U8967 (N_8967,N_8601,N_8690);
nand U8968 (N_8968,N_8664,N_8548);
nand U8969 (N_8969,N_8514,N_8476);
xnor U8970 (N_8970,N_8551,N_8409);
nand U8971 (N_8971,N_8633,N_8405);
and U8972 (N_8972,N_8564,N_8406);
xor U8973 (N_8973,N_8638,N_8546);
nand U8974 (N_8974,N_8675,N_8573);
nor U8975 (N_8975,N_8693,N_8484);
or U8976 (N_8976,N_8680,N_8628);
and U8977 (N_8977,N_8666,N_8671);
xor U8978 (N_8978,N_8548,N_8465);
nor U8979 (N_8979,N_8621,N_8409);
nor U8980 (N_8980,N_8549,N_8512);
nor U8981 (N_8981,N_8404,N_8687);
nor U8982 (N_8982,N_8628,N_8440);
xnor U8983 (N_8983,N_8509,N_8614);
nor U8984 (N_8984,N_8645,N_8464);
or U8985 (N_8985,N_8665,N_8407);
nor U8986 (N_8986,N_8437,N_8615);
xnor U8987 (N_8987,N_8541,N_8633);
xnor U8988 (N_8988,N_8588,N_8539);
xnor U8989 (N_8989,N_8536,N_8661);
or U8990 (N_8990,N_8507,N_8533);
nor U8991 (N_8991,N_8698,N_8672);
and U8992 (N_8992,N_8609,N_8520);
and U8993 (N_8993,N_8527,N_8464);
and U8994 (N_8994,N_8525,N_8426);
xnor U8995 (N_8995,N_8585,N_8547);
and U8996 (N_8996,N_8678,N_8436);
nand U8997 (N_8997,N_8600,N_8631);
nand U8998 (N_8998,N_8534,N_8513);
and U8999 (N_8999,N_8691,N_8519);
nand U9000 (N_9000,N_8756,N_8814);
or U9001 (N_9001,N_8985,N_8937);
and U9002 (N_9002,N_8707,N_8702);
and U9003 (N_9003,N_8921,N_8722);
nand U9004 (N_9004,N_8719,N_8824);
or U9005 (N_9005,N_8741,N_8996);
xnor U9006 (N_9006,N_8984,N_8864);
xor U9007 (N_9007,N_8933,N_8713);
xor U9008 (N_9008,N_8777,N_8839);
or U9009 (N_9009,N_8907,N_8795);
nand U9010 (N_9010,N_8914,N_8769);
or U9011 (N_9011,N_8730,N_8997);
xor U9012 (N_9012,N_8855,N_8759);
or U9013 (N_9013,N_8764,N_8863);
or U9014 (N_9014,N_8762,N_8925);
and U9015 (N_9015,N_8960,N_8938);
xor U9016 (N_9016,N_8705,N_8866);
nor U9017 (N_9017,N_8889,N_8879);
nor U9018 (N_9018,N_8877,N_8782);
and U9019 (N_9019,N_8906,N_8919);
and U9020 (N_9020,N_8706,N_8740);
nor U9021 (N_9021,N_8783,N_8942);
xor U9022 (N_9022,N_8733,N_8884);
xnor U9023 (N_9023,N_8840,N_8749);
nor U9024 (N_9024,N_8941,N_8905);
xor U9025 (N_9025,N_8802,N_8860);
or U9026 (N_9026,N_8931,N_8966);
and U9027 (N_9027,N_8867,N_8904);
xor U9028 (N_9028,N_8980,N_8868);
xnor U9029 (N_9029,N_8735,N_8853);
nor U9030 (N_9030,N_8956,N_8793);
xor U9031 (N_9031,N_8844,N_8896);
or U9032 (N_9032,N_8776,N_8858);
or U9033 (N_9033,N_8750,N_8967);
or U9034 (N_9034,N_8862,N_8943);
xnor U9035 (N_9035,N_8700,N_8848);
or U9036 (N_9036,N_8989,N_8959);
or U9037 (N_9037,N_8987,N_8771);
nand U9038 (N_9038,N_8727,N_8948);
and U9039 (N_9039,N_8913,N_8892);
or U9040 (N_9040,N_8986,N_8708);
and U9041 (N_9041,N_8873,N_8786);
nand U9042 (N_9042,N_8851,N_8871);
nand U9043 (N_9043,N_8843,N_8774);
and U9044 (N_9044,N_8798,N_8974);
xor U9045 (N_9045,N_8990,N_8852);
or U9046 (N_9046,N_8975,N_8809);
and U9047 (N_9047,N_8951,N_8703);
or U9048 (N_9048,N_8901,N_8888);
or U9049 (N_9049,N_8940,N_8953);
or U9050 (N_9050,N_8711,N_8801);
xnor U9051 (N_9051,N_8817,N_8826);
or U9052 (N_9052,N_8882,N_8757);
nor U9053 (N_9053,N_8909,N_8857);
xor U9054 (N_9054,N_8712,N_8977);
and U9055 (N_9055,N_8710,N_8731);
nor U9056 (N_9056,N_8910,N_8761);
nor U9057 (N_9057,N_8954,N_8746);
or U9058 (N_9058,N_8739,N_8994);
nor U9059 (N_9059,N_8726,N_8790);
and U9060 (N_9060,N_8936,N_8821);
xnor U9061 (N_9061,N_8923,N_8898);
nor U9062 (N_9062,N_8766,N_8827);
nand U9063 (N_9063,N_8865,N_8934);
xnor U9064 (N_9064,N_8822,N_8932);
and U9065 (N_9065,N_8788,N_8732);
nor U9066 (N_9066,N_8908,N_8971);
nand U9067 (N_9067,N_8963,N_8995);
and U9068 (N_9068,N_8773,N_8818);
nand U9069 (N_9069,N_8811,N_8955);
xor U9070 (N_9070,N_8847,N_8799);
and U9071 (N_9071,N_8869,N_8830);
or U9072 (N_9072,N_8701,N_8982);
and U9073 (N_9073,N_8881,N_8754);
xnor U9074 (N_9074,N_8856,N_8887);
nor U9075 (N_9075,N_8748,N_8874);
and U9076 (N_9076,N_8778,N_8758);
nand U9077 (N_9077,N_8981,N_8861);
nand U9078 (N_9078,N_8895,N_8765);
or U9079 (N_9079,N_8952,N_8823);
or U9080 (N_9080,N_8886,N_8875);
xnor U9081 (N_9081,N_8893,N_8784);
or U9082 (N_9082,N_8890,N_8787);
nand U9083 (N_9083,N_8880,N_8961);
or U9084 (N_9084,N_8983,N_8806);
and U9085 (N_9085,N_8999,N_8792);
nor U9086 (N_9086,N_8973,N_8946);
or U9087 (N_9087,N_8725,N_8714);
nand U9088 (N_9088,N_8870,N_8922);
nor U9089 (N_9089,N_8841,N_8850);
nor U9090 (N_9090,N_8718,N_8900);
xor U9091 (N_9091,N_8742,N_8717);
nor U9092 (N_9092,N_8838,N_8958);
xor U9093 (N_9093,N_8927,N_8849);
xor U9094 (N_9094,N_8704,N_8715);
nor U9095 (N_9095,N_8835,N_8815);
xnor U9096 (N_9096,N_8816,N_8998);
nand U9097 (N_9097,N_8796,N_8926);
or U9098 (N_9098,N_8785,N_8939);
nor U9099 (N_9099,N_8970,N_8709);
and U9100 (N_9100,N_8859,N_8918);
nand U9101 (N_9101,N_8964,N_8755);
xor U9102 (N_9102,N_8779,N_8807);
nand U9103 (N_9103,N_8969,N_8897);
or U9104 (N_9104,N_8916,N_8902);
xor U9105 (N_9105,N_8834,N_8911);
or U9106 (N_9106,N_8930,N_8976);
nor U9107 (N_9107,N_8944,N_8734);
nor U9108 (N_9108,N_8772,N_8720);
nor U9109 (N_9109,N_8716,N_8878);
or U9110 (N_9110,N_8894,N_8723);
nand U9111 (N_9111,N_8804,N_8978);
nor U9112 (N_9112,N_8770,N_8949);
nand U9113 (N_9113,N_8872,N_8775);
nand U9114 (N_9114,N_8794,N_8763);
nor U9115 (N_9115,N_8979,N_8876);
nand U9116 (N_9116,N_8885,N_8812);
nand U9117 (N_9117,N_8992,N_8842);
and U9118 (N_9118,N_8810,N_8950);
xnor U9119 (N_9119,N_8744,N_8831);
nor U9120 (N_9120,N_8800,N_8743);
or U9121 (N_9121,N_8828,N_8920);
nor U9122 (N_9122,N_8760,N_8968);
and U9123 (N_9123,N_8747,N_8833);
nand U9124 (N_9124,N_8945,N_8803);
and U9125 (N_9125,N_8780,N_8768);
and U9126 (N_9126,N_8846,N_8752);
and U9127 (N_9127,N_8819,N_8737);
and U9128 (N_9128,N_8965,N_8808);
nand U9129 (N_9129,N_8825,N_8728);
and U9130 (N_9130,N_8781,N_8854);
nor U9131 (N_9131,N_8729,N_8829);
xor U9132 (N_9132,N_8845,N_8767);
nor U9133 (N_9133,N_8753,N_8797);
nor U9134 (N_9134,N_8837,N_8899);
nand U9135 (N_9135,N_8993,N_8791);
or U9136 (N_9136,N_8836,N_8805);
nor U9137 (N_9137,N_8929,N_8751);
nor U9138 (N_9138,N_8917,N_8988);
nand U9139 (N_9139,N_8745,N_8915);
xnor U9140 (N_9140,N_8738,N_8991);
and U9141 (N_9141,N_8928,N_8820);
xor U9142 (N_9142,N_8962,N_8947);
nand U9143 (N_9143,N_8957,N_8724);
and U9144 (N_9144,N_8721,N_8883);
nand U9145 (N_9145,N_8789,N_8935);
and U9146 (N_9146,N_8924,N_8891);
nand U9147 (N_9147,N_8736,N_8912);
nand U9148 (N_9148,N_8813,N_8972);
nand U9149 (N_9149,N_8903,N_8832);
nand U9150 (N_9150,N_8807,N_8906);
xnor U9151 (N_9151,N_8831,N_8897);
nand U9152 (N_9152,N_8938,N_8911);
nor U9153 (N_9153,N_8835,N_8740);
and U9154 (N_9154,N_8910,N_8925);
xnor U9155 (N_9155,N_8820,N_8969);
nor U9156 (N_9156,N_8750,N_8838);
nand U9157 (N_9157,N_8990,N_8922);
or U9158 (N_9158,N_8729,N_8862);
xnor U9159 (N_9159,N_8913,N_8926);
or U9160 (N_9160,N_8929,N_8794);
and U9161 (N_9161,N_8753,N_8727);
nor U9162 (N_9162,N_8930,N_8888);
nand U9163 (N_9163,N_8733,N_8921);
xor U9164 (N_9164,N_8771,N_8792);
nand U9165 (N_9165,N_8949,N_8903);
nor U9166 (N_9166,N_8756,N_8739);
nor U9167 (N_9167,N_8932,N_8928);
nand U9168 (N_9168,N_8834,N_8746);
nand U9169 (N_9169,N_8703,N_8784);
nor U9170 (N_9170,N_8903,N_8721);
nand U9171 (N_9171,N_8770,N_8991);
nor U9172 (N_9172,N_8912,N_8977);
nand U9173 (N_9173,N_8945,N_8728);
nand U9174 (N_9174,N_8924,N_8878);
nand U9175 (N_9175,N_8998,N_8795);
or U9176 (N_9176,N_8722,N_8781);
xor U9177 (N_9177,N_8998,N_8802);
nor U9178 (N_9178,N_8839,N_8867);
or U9179 (N_9179,N_8978,N_8823);
nor U9180 (N_9180,N_8913,N_8777);
or U9181 (N_9181,N_8736,N_8843);
nor U9182 (N_9182,N_8866,N_8877);
and U9183 (N_9183,N_8766,N_8769);
nor U9184 (N_9184,N_8911,N_8856);
nor U9185 (N_9185,N_8832,N_8711);
or U9186 (N_9186,N_8835,N_8950);
xor U9187 (N_9187,N_8909,N_8707);
nor U9188 (N_9188,N_8934,N_8856);
nand U9189 (N_9189,N_8887,N_8815);
nor U9190 (N_9190,N_8994,N_8774);
and U9191 (N_9191,N_8827,N_8843);
nand U9192 (N_9192,N_8775,N_8902);
nor U9193 (N_9193,N_8805,N_8876);
nand U9194 (N_9194,N_8711,N_8992);
nand U9195 (N_9195,N_8793,N_8851);
or U9196 (N_9196,N_8738,N_8715);
and U9197 (N_9197,N_8878,N_8900);
xor U9198 (N_9198,N_8731,N_8808);
xor U9199 (N_9199,N_8829,N_8818);
xnor U9200 (N_9200,N_8943,N_8876);
nor U9201 (N_9201,N_8758,N_8958);
xnor U9202 (N_9202,N_8998,N_8735);
nor U9203 (N_9203,N_8894,N_8785);
xnor U9204 (N_9204,N_8920,N_8860);
and U9205 (N_9205,N_8945,N_8707);
nand U9206 (N_9206,N_8843,N_8745);
nor U9207 (N_9207,N_8704,N_8709);
nand U9208 (N_9208,N_8725,N_8909);
nand U9209 (N_9209,N_8795,N_8773);
nor U9210 (N_9210,N_8804,N_8730);
nand U9211 (N_9211,N_8914,N_8860);
nor U9212 (N_9212,N_8956,N_8984);
nor U9213 (N_9213,N_8700,N_8837);
xor U9214 (N_9214,N_8967,N_8991);
xor U9215 (N_9215,N_8844,N_8867);
xnor U9216 (N_9216,N_8821,N_8764);
and U9217 (N_9217,N_8749,N_8923);
and U9218 (N_9218,N_8872,N_8954);
nor U9219 (N_9219,N_8795,N_8879);
xnor U9220 (N_9220,N_8818,N_8887);
xor U9221 (N_9221,N_8989,N_8795);
nor U9222 (N_9222,N_8916,N_8705);
nand U9223 (N_9223,N_8987,N_8873);
and U9224 (N_9224,N_8958,N_8711);
nor U9225 (N_9225,N_8728,N_8903);
nor U9226 (N_9226,N_8796,N_8818);
and U9227 (N_9227,N_8911,N_8918);
xnor U9228 (N_9228,N_8870,N_8978);
and U9229 (N_9229,N_8844,N_8753);
nand U9230 (N_9230,N_8828,N_8780);
xor U9231 (N_9231,N_8827,N_8760);
or U9232 (N_9232,N_8730,N_8797);
and U9233 (N_9233,N_8983,N_8846);
and U9234 (N_9234,N_8923,N_8735);
xor U9235 (N_9235,N_8741,N_8705);
xor U9236 (N_9236,N_8902,N_8927);
nand U9237 (N_9237,N_8953,N_8742);
or U9238 (N_9238,N_8950,N_8900);
nand U9239 (N_9239,N_8723,N_8933);
nand U9240 (N_9240,N_8881,N_8720);
or U9241 (N_9241,N_8700,N_8881);
or U9242 (N_9242,N_8932,N_8830);
and U9243 (N_9243,N_8740,N_8794);
xor U9244 (N_9244,N_8723,N_8777);
or U9245 (N_9245,N_8714,N_8785);
xor U9246 (N_9246,N_8701,N_8946);
xor U9247 (N_9247,N_8780,N_8940);
or U9248 (N_9248,N_8809,N_8928);
nand U9249 (N_9249,N_8765,N_8712);
nand U9250 (N_9250,N_8894,N_8771);
nand U9251 (N_9251,N_8782,N_8783);
or U9252 (N_9252,N_8721,N_8717);
or U9253 (N_9253,N_8915,N_8946);
and U9254 (N_9254,N_8785,N_8866);
or U9255 (N_9255,N_8881,N_8843);
nand U9256 (N_9256,N_8852,N_8714);
or U9257 (N_9257,N_8895,N_8826);
and U9258 (N_9258,N_8702,N_8801);
nand U9259 (N_9259,N_8732,N_8949);
and U9260 (N_9260,N_8872,N_8748);
xnor U9261 (N_9261,N_8969,N_8982);
nor U9262 (N_9262,N_8820,N_8918);
nor U9263 (N_9263,N_8785,N_8893);
or U9264 (N_9264,N_8970,N_8956);
xor U9265 (N_9265,N_8716,N_8984);
nor U9266 (N_9266,N_8845,N_8725);
nand U9267 (N_9267,N_8842,N_8886);
or U9268 (N_9268,N_8995,N_8801);
nor U9269 (N_9269,N_8975,N_8777);
nor U9270 (N_9270,N_8915,N_8803);
nand U9271 (N_9271,N_8947,N_8949);
nor U9272 (N_9272,N_8757,N_8772);
nor U9273 (N_9273,N_8961,N_8930);
or U9274 (N_9274,N_8813,N_8965);
and U9275 (N_9275,N_8794,N_8723);
nor U9276 (N_9276,N_8763,N_8987);
nor U9277 (N_9277,N_8956,N_8722);
and U9278 (N_9278,N_8721,N_8980);
and U9279 (N_9279,N_8936,N_8964);
xor U9280 (N_9280,N_8910,N_8952);
and U9281 (N_9281,N_8987,N_8787);
and U9282 (N_9282,N_8841,N_8762);
or U9283 (N_9283,N_8770,N_8906);
xor U9284 (N_9284,N_8949,N_8942);
nand U9285 (N_9285,N_8967,N_8948);
xnor U9286 (N_9286,N_8844,N_8873);
xnor U9287 (N_9287,N_8875,N_8712);
nor U9288 (N_9288,N_8972,N_8998);
nand U9289 (N_9289,N_8801,N_8928);
or U9290 (N_9290,N_8741,N_8907);
or U9291 (N_9291,N_8949,N_8979);
xor U9292 (N_9292,N_8947,N_8964);
and U9293 (N_9293,N_8889,N_8990);
xor U9294 (N_9294,N_8829,N_8722);
xnor U9295 (N_9295,N_8794,N_8811);
nand U9296 (N_9296,N_8747,N_8719);
xnor U9297 (N_9297,N_8888,N_8833);
and U9298 (N_9298,N_8747,N_8993);
and U9299 (N_9299,N_8948,N_8979);
xor U9300 (N_9300,N_9194,N_9085);
nand U9301 (N_9301,N_9004,N_9128);
nand U9302 (N_9302,N_9141,N_9147);
nor U9303 (N_9303,N_9188,N_9240);
nor U9304 (N_9304,N_9017,N_9193);
xnor U9305 (N_9305,N_9047,N_9173);
or U9306 (N_9306,N_9219,N_9299);
or U9307 (N_9307,N_9296,N_9108);
nor U9308 (N_9308,N_9073,N_9131);
or U9309 (N_9309,N_9214,N_9238);
or U9310 (N_9310,N_9142,N_9282);
nor U9311 (N_9311,N_9092,N_9234);
or U9312 (N_9312,N_9197,N_9094);
and U9313 (N_9313,N_9089,N_9156);
and U9314 (N_9314,N_9080,N_9144);
xor U9315 (N_9315,N_9145,N_9038);
or U9316 (N_9316,N_9235,N_9015);
or U9317 (N_9317,N_9054,N_9140);
xnor U9318 (N_9318,N_9000,N_9143);
or U9319 (N_9319,N_9212,N_9175);
nand U9320 (N_9320,N_9063,N_9130);
or U9321 (N_9321,N_9064,N_9254);
and U9322 (N_9322,N_9158,N_9023);
xnor U9323 (N_9323,N_9151,N_9226);
nand U9324 (N_9324,N_9280,N_9098);
nand U9325 (N_9325,N_9074,N_9203);
and U9326 (N_9326,N_9267,N_9069);
nor U9327 (N_9327,N_9225,N_9198);
or U9328 (N_9328,N_9020,N_9184);
nand U9329 (N_9329,N_9215,N_9230);
and U9330 (N_9330,N_9076,N_9115);
or U9331 (N_9331,N_9272,N_9041);
xnor U9332 (N_9332,N_9290,N_9171);
xnor U9333 (N_9333,N_9291,N_9232);
and U9334 (N_9334,N_9211,N_9228);
nor U9335 (N_9335,N_9132,N_9137);
nand U9336 (N_9336,N_9003,N_9260);
and U9337 (N_9337,N_9164,N_9236);
and U9338 (N_9338,N_9192,N_9163);
or U9339 (N_9339,N_9283,N_9152);
and U9340 (N_9340,N_9106,N_9066);
xnor U9341 (N_9341,N_9072,N_9118);
or U9342 (N_9342,N_9046,N_9071);
xnor U9343 (N_9343,N_9249,N_9129);
xor U9344 (N_9344,N_9185,N_9273);
nor U9345 (N_9345,N_9149,N_9195);
nor U9346 (N_9346,N_9032,N_9202);
nand U9347 (N_9347,N_9006,N_9133);
xnor U9348 (N_9348,N_9010,N_9043);
and U9349 (N_9349,N_9199,N_9084);
and U9350 (N_9350,N_9019,N_9035);
or U9351 (N_9351,N_9079,N_9012);
or U9352 (N_9352,N_9157,N_9264);
nand U9353 (N_9353,N_9159,N_9075);
or U9354 (N_9354,N_9101,N_9088);
nor U9355 (N_9355,N_9077,N_9031);
or U9356 (N_9356,N_9105,N_9252);
or U9357 (N_9357,N_9110,N_9218);
nand U9358 (N_9358,N_9247,N_9204);
or U9359 (N_9359,N_9059,N_9102);
xor U9360 (N_9360,N_9227,N_9025);
and U9361 (N_9361,N_9165,N_9169);
or U9362 (N_9362,N_9055,N_9201);
nand U9363 (N_9363,N_9109,N_9001);
or U9364 (N_9364,N_9170,N_9295);
or U9365 (N_9365,N_9275,N_9253);
nor U9366 (N_9366,N_9274,N_9242);
xnor U9367 (N_9367,N_9208,N_9166);
nor U9368 (N_9368,N_9224,N_9136);
xor U9369 (N_9369,N_9103,N_9243);
and U9370 (N_9370,N_9277,N_9021);
xor U9371 (N_9371,N_9002,N_9206);
and U9372 (N_9372,N_9138,N_9297);
nand U9373 (N_9373,N_9286,N_9030);
nor U9374 (N_9374,N_9107,N_9153);
nand U9375 (N_9375,N_9221,N_9263);
nand U9376 (N_9376,N_9210,N_9276);
or U9377 (N_9377,N_9217,N_9248);
xor U9378 (N_9378,N_9083,N_9177);
nor U9379 (N_9379,N_9150,N_9257);
and U9380 (N_9380,N_9237,N_9011);
nor U9381 (N_9381,N_9082,N_9117);
nand U9382 (N_9382,N_9097,N_9048);
and U9383 (N_9383,N_9258,N_9246);
nand U9384 (N_9384,N_9095,N_9284);
nor U9385 (N_9385,N_9124,N_9014);
xor U9386 (N_9386,N_9172,N_9182);
or U9387 (N_9387,N_9294,N_9278);
nand U9388 (N_9388,N_9281,N_9233);
xnor U9389 (N_9389,N_9087,N_9116);
nor U9390 (N_9390,N_9125,N_9259);
nand U9391 (N_9391,N_9051,N_9178);
or U9392 (N_9392,N_9056,N_9018);
nand U9393 (N_9393,N_9007,N_9288);
nand U9394 (N_9394,N_9070,N_9127);
and U9395 (N_9395,N_9262,N_9062);
xnor U9396 (N_9396,N_9268,N_9005);
nand U9397 (N_9397,N_9112,N_9126);
or U9398 (N_9398,N_9207,N_9053);
and U9399 (N_9399,N_9293,N_9200);
or U9400 (N_9400,N_9086,N_9256);
and U9401 (N_9401,N_9216,N_9036);
xnor U9402 (N_9402,N_9270,N_9067);
nor U9403 (N_9403,N_9060,N_9065);
xnor U9404 (N_9404,N_9090,N_9245);
xnor U9405 (N_9405,N_9050,N_9068);
and U9406 (N_9406,N_9190,N_9146);
and U9407 (N_9407,N_9167,N_9155);
nand U9408 (N_9408,N_9261,N_9134);
xor U9409 (N_9409,N_9162,N_9255);
xor U9410 (N_9410,N_9244,N_9148);
or U9411 (N_9411,N_9220,N_9223);
or U9412 (N_9412,N_9093,N_9289);
and U9413 (N_9413,N_9049,N_9028);
and U9414 (N_9414,N_9292,N_9123);
and U9415 (N_9415,N_9026,N_9027);
nand U9416 (N_9416,N_9231,N_9044);
nand U9417 (N_9417,N_9269,N_9100);
nand U9418 (N_9418,N_9013,N_9168);
and U9419 (N_9419,N_9139,N_9121);
nand U9420 (N_9420,N_9285,N_9271);
xnor U9421 (N_9421,N_9196,N_9120);
or U9422 (N_9422,N_9209,N_9008);
nand U9423 (N_9423,N_9187,N_9287);
xnor U9424 (N_9424,N_9229,N_9265);
nand U9425 (N_9425,N_9042,N_9052);
or U9426 (N_9426,N_9266,N_9174);
xnor U9427 (N_9427,N_9298,N_9250);
nor U9428 (N_9428,N_9176,N_9111);
nand U9429 (N_9429,N_9181,N_9114);
and U9430 (N_9430,N_9183,N_9104);
or U9431 (N_9431,N_9039,N_9029);
xnor U9432 (N_9432,N_9091,N_9161);
xnor U9433 (N_9433,N_9096,N_9058);
and U9434 (N_9434,N_9179,N_9024);
nand U9435 (N_9435,N_9022,N_9037);
nand U9436 (N_9436,N_9186,N_9189);
nand U9437 (N_9437,N_9154,N_9222);
xor U9438 (N_9438,N_9061,N_9180);
or U9439 (N_9439,N_9251,N_9034);
and U9440 (N_9440,N_9122,N_9113);
and U9441 (N_9441,N_9040,N_9033);
nand U9442 (N_9442,N_9081,N_9191);
and U9443 (N_9443,N_9241,N_9279);
and U9444 (N_9444,N_9078,N_9205);
nor U9445 (N_9445,N_9099,N_9045);
or U9446 (N_9446,N_9009,N_9135);
xor U9447 (N_9447,N_9213,N_9239);
or U9448 (N_9448,N_9016,N_9160);
or U9449 (N_9449,N_9119,N_9057);
and U9450 (N_9450,N_9010,N_9223);
or U9451 (N_9451,N_9136,N_9109);
xnor U9452 (N_9452,N_9055,N_9085);
or U9453 (N_9453,N_9092,N_9158);
nor U9454 (N_9454,N_9182,N_9135);
or U9455 (N_9455,N_9022,N_9083);
and U9456 (N_9456,N_9147,N_9005);
xnor U9457 (N_9457,N_9275,N_9266);
xnor U9458 (N_9458,N_9146,N_9017);
and U9459 (N_9459,N_9089,N_9169);
and U9460 (N_9460,N_9083,N_9191);
xor U9461 (N_9461,N_9238,N_9049);
nand U9462 (N_9462,N_9169,N_9069);
nand U9463 (N_9463,N_9013,N_9126);
or U9464 (N_9464,N_9112,N_9176);
or U9465 (N_9465,N_9127,N_9129);
or U9466 (N_9466,N_9108,N_9200);
xor U9467 (N_9467,N_9083,N_9125);
or U9468 (N_9468,N_9061,N_9203);
and U9469 (N_9469,N_9133,N_9244);
nand U9470 (N_9470,N_9289,N_9166);
or U9471 (N_9471,N_9259,N_9179);
nand U9472 (N_9472,N_9179,N_9007);
or U9473 (N_9473,N_9085,N_9076);
or U9474 (N_9474,N_9108,N_9078);
and U9475 (N_9475,N_9110,N_9238);
or U9476 (N_9476,N_9181,N_9207);
and U9477 (N_9477,N_9242,N_9032);
nor U9478 (N_9478,N_9241,N_9228);
and U9479 (N_9479,N_9010,N_9231);
xor U9480 (N_9480,N_9124,N_9142);
or U9481 (N_9481,N_9299,N_9076);
nor U9482 (N_9482,N_9089,N_9036);
or U9483 (N_9483,N_9227,N_9096);
xor U9484 (N_9484,N_9018,N_9028);
or U9485 (N_9485,N_9216,N_9194);
and U9486 (N_9486,N_9049,N_9256);
nor U9487 (N_9487,N_9194,N_9142);
and U9488 (N_9488,N_9190,N_9170);
xor U9489 (N_9489,N_9136,N_9118);
or U9490 (N_9490,N_9259,N_9199);
and U9491 (N_9491,N_9188,N_9002);
and U9492 (N_9492,N_9094,N_9116);
nor U9493 (N_9493,N_9023,N_9155);
or U9494 (N_9494,N_9128,N_9295);
nor U9495 (N_9495,N_9079,N_9159);
nor U9496 (N_9496,N_9231,N_9082);
and U9497 (N_9497,N_9158,N_9250);
nor U9498 (N_9498,N_9163,N_9006);
or U9499 (N_9499,N_9167,N_9203);
or U9500 (N_9500,N_9166,N_9113);
nand U9501 (N_9501,N_9007,N_9084);
and U9502 (N_9502,N_9131,N_9041);
nand U9503 (N_9503,N_9196,N_9135);
and U9504 (N_9504,N_9088,N_9272);
or U9505 (N_9505,N_9100,N_9002);
xor U9506 (N_9506,N_9198,N_9152);
and U9507 (N_9507,N_9113,N_9189);
nand U9508 (N_9508,N_9138,N_9274);
or U9509 (N_9509,N_9253,N_9049);
xnor U9510 (N_9510,N_9130,N_9117);
nand U9511 (N_9511,N_9214,N_9257);
xnor U9512 (N_9512,N_9242,N_9200);
nand U9513 (N_9513,N_9271,N_9258);
xor U9514 (N_9514,N_9194,N_9198);
nand U9515 (N_9515,N_9132,N_9243);
nand U9516 (N_9516,N_9022,N_9019);
and U9517 (N_9517,N_9045,N_9030);
and U9518 (N_9518,N_9169,N_9277);
xnor U9519 (N_9519,N_9189,N_9077);
or U9520 (N_9520,N_9007,N_9151);
and U9521 (N_9521,N_9050,N_9171);
xor U9522 (N_9522,N_9074,N_9103);
and U9523 (N_9523,N_9282,N_9166);
nand U9524 (N_9524,N_9059,N_9054);
and U9525 (N_9525,N_9155,N_9213);
and U9526 (N_9526,N_9024,N_9255);
nor U9527 (N_9527,N_9048,N_9245);
xor U9528 (N_9528,N_9091,N_9047);
nand U9529 (N_9529,N_9139,N_9243);
nand U9530 (N_9530,N_9122,N_9224);
xnor U9531 (N_9531,N_9296,N_9175);
or U9532 (N_9532,N_9135,N_9214);
nand U9533 (N_9533,N_9296,N_9176);
xor U9534 (N_9534,N_9203,N_9059);
nor U9535 (N_9535,N_9193,N_9272);
and U9536 (N_9536,N_9008,N_9110);
nand U9537 (N_9537,N_9170,N_9249);
and U9538 (N_9538,N_9058,N_9013);
nand U9539 (N_9539,N_9152,N_9268);
and U9540 (N_9540,N_9032,N_9187);
xor U9541 (N_9541,N_9216,N_9120);
nor U9542 (N_9542,N_9225,N_9029);
nand U9543 (N_9543,N_9187,N_9021);
nand U9544 (N_9544,N_9128,N_9053);
nor U9545 (N_9545,N_9092,N_9298);
nand U9546 (N_9546,N_9024,N_9073);
nand U9547 (N_9547,N_9003,N_9217);
or U9548 (N_9548,N_9071,N_9007);
xnor U9549 (N_9549,N_9086,N_9105);
xor U9550 (N_9550,N_9130,N_9218);
and U9551 (N_9551,N_9234,N_9209);
and U9552 (N_9552,N_9257,N_9068);
xor U9553 (N_9553,N_9062,N_9240);
and U9554 (N_9554,N_9010,N_9274);
or U9555 (N_9555,N_9216,N_9231);
or U9556 (N_9556,N_9007,N_9116);
and U9557 (N_9557,N_9177,N_9065);
or U9558 (N_9558,N_9292,N_9150);
and U9559 (N_9559,N_9161,N_9123);
and U9560 (N_9560,N_9222,N_9283);
nor U9561 (N_9561,N_9129,N_9040);
and U9562 (N_9562,N_9082,N_9053);
or U9563 (N_9563,N_9181,N_9241);
nor U9564 (N_9564,N_9001,N_9162);
nand U9565 (N_9565,N_9194,N_9129);
and U9566 (N_9566,N_9040,N_9255);
nor U9567 (N_9567,N_9155,N_9224);
and U9568 (N_9568,N_9218,N_9281);
nand U9569 (N_9569,N_9261,N_9064);
nor U9570 (N_9570,N_9274,N_9034);
nor U9571 (N_9571,N_9294,N_9286);
or U9572 (N_9572,N_9116,N_9221);
or U9573 (N_9573,N_9122,N_9089);
nand U9574 (N_9574,N_9237,N_9013);
xnor U9575 (N_9575,N_9068,N_9039);
and U9576 (N_9576,N_9058,N_9292);
and U9577 (N_9577,N_9033,N_9036);
or U9578 (N_9578,N_9184,N_9175);
and U9579 (N_9579,N_9006,N_9260);
nor U9580 (N_9580,N_9002,N_9185);
and U9581 (N_9581,N_9210,N_9195);
xnor U9582 (N_9582,N_9182,N_9091);
nor U9583 (N_9583,N_9111,N_9145);
nand U9584 (N_9584,N_9180,N_9256);
nand U9585 (N_9585,N_9054,N_9249);
or U9586 (N_9586,N_9021,N_9276);
nor U9587 (N_9587,N_9075,N_9231);
and U9588 (N_9588,N_9078,N_9059);
or U9589 (N_9589,N_9051,N_9295);
or U9590 (N_9590,N_9169,N_9296);
or U9591 (N_9591,N_9080,N_9187);
xor U9592 (N_9592,N_9159,N_9190);
nand U9593 (N_9593,N_9169,N_9045);
nor U9594 (N_9594,N_9107,N_9005);
or U9595 (N_9595,N_9272,N_9206);
nor U9596 (N_9596,N_9104,N_9253);
xnor U9597 (N_9597,N_9085,N_9183);
nand U9598 (N_9598,N_9139,N_9049);
xor U9599 (N_9599,N_9213,N_9090);
and U9600 (N_9600,N_9514,N_9385);
xor U9601 (N_9601,N_9392,N_9304);
nand U9602 (N_9602,N_9391,N_9316);
nor U9603 (N_9603,N_9563,N_9310);
xnor U9604 (N_9604,N_9510,N_9548);
nand U9605 (N_9605,N_9408,N_9443);
or U9606 (N_9606,N_9457,N_9415);
or U9607 (N_9607,N_9354,N_9303);
nand U9608 (N_9608,N_9453,N_9545);
xor U9609 (N_9609,N_9557,N_9322);
and U9610 (N_9610,N_9465,N_9592);
xor U9611 (N_9611,N_9412,N_9596);
xor U9612 (N_9612,N_9504,N_9447);
xor U9613 (N_9613,N_9530,N_9405);
nor U9614 (N_9614,N_9461,N_9484);
or U9615 (N_9615,N_9474,N_9559);
and U9616 (N_9616,N_9475,N_9355);
or U9617 (N_9617,N_9452,N_9468);
nand U9618 (N_9618,N_9481,N_9439);
nand U9619 (N_9619,N_9360,N_9571);
xor U9620 (N_9620,N_9471,N_9525);
and U9621 (N_9621,N_9353,N_9448);
and U9622 (N_9622,N_9488,N_9327);
and U9623 (N_9623,N_9527,N_9421);
nand U9624 (N_9624,N_9578,N_9324);
nand U9625 (N_9625,N_9537,N_9584);
nand U9626 (N_9626,N_9547,N_9572);
nand U9627 (N_9627,N_9430,N_9441);
nand U9628 (N_9628,N_9554,N_9365);
and U9629 (N_9629,N_9402,N_9494);
and U9630 (N_9630,N_9541,N_9553);
nand U9631 (N_9631,N_9486,N_9312);
nand U9632 (N_9632,N_9544,N_9406);
nor U9633 (N_9633,N_9321,N_9535);
nor U9634 (N_9634,N_9536,N_9518);
nor U9635 (N_9635,N_9577,N_9466);
nand U9636 (N_9636,N_9463,N_9590);
nor U9637 (N_9637,N_9440,N_9368);
nand U9638 (N_9638,N_9561,N_9422);
nand U9639 (N_9639,N_9582,N_9524);
or U9640 (N_9640,N_9509,N_9338);
xor U9641 (N_9641,N_9476,N_9386);
and U9642 (N_9642,N_9387,N_9459);
nor U9643 (N_9643,N_9332,N_9323);
nand U9644 (N_9644,N_9515,N_9352);
or U9645 (N_9645,N_9529,N_9552);
nor U9646 (N_9646,N_9485,N_9589);
nor U9647 (N_9647,N_9328,N_9302);
nor U9648 (N_9648,N_9482,N_9366);
xnor U9649 (N_9649,N_9330,N_9341);
and U9650 (N_9650,N_9395,N_9523);
xnor U9651 (N_9651,N_9378,N_9361);
or U9652 (N_9652,N_9414,N_9339);
or U9653 (N_9653,N_9428,N_9423);
or U9654 (N_9654,N_9320,N_9307);
and U9655 (N_9655,N_9556,N_9505);
nor U9656 (N_9656,N_9470,N_9326);
or U9657 (N_9657,N_9492,N_9427);
or U9658 (N_9658,N_9319,N_9379);
xor U9659 (N_9659,N_9511,N_9512);
and U9660 (N_9660,N_9346,N_9384);
nand U9661 (N_9661,N_9560,N_9513);
xor U9662 (N_9662,N_9424,N_9426);
and U9663 (N_9663,N_9495,N_9570);
and U9664 (N_9664,N_9493,N_9585);
nand U9665 (N_9665,N_9579,N_9367);
or U9666 (N_9666,N_9543,N_9314);
nor U9667 (N_9667,N_9329,N_9315);
nor U9668 (N_9668,N_9532,N_9507);
xor U9669 (N_9669,N_9540,N_9377);
xor U9670 (N_9670,N_9357,N_9300);
xor U9671 (N_9671,N_9490,N_9587);
nand U9672 (N_9672,N_9508,N_9397);
nand U9673 (N_9673,N_9417,N_9568);
xnor U9674 (N_9674,N_9342,N_9398);
or U9675 (N_9675,N_9337,N_9376);
nor U9676 (N_9676,N_9373,N_9340);
or U9677 (N_9677,N_9413,N_9432);
nand U9678 (N_9678,N_9335,N_9308);
xor U9679 (N_9679,N_9473,N_9374);
and U9680 (N_9680,N_9382,N_9363);
or U9681 (N_9681,N_9549,N_9349);
nand U9682 (N_9682,N_9467,N_9567);
or U9683 (N_9683,N_9450,N_9442);
or U9684 (N_9684,N_9517,N_9479);
and U9685 (N_9685,N_9436,N_9400);
xor U9686 (N_9686,N_9528,N_9516);
nand U9687 (N_9687,N_9588,N_9569);
nor U9688 (N_9688,N_9343,N_9317);
nand U9689 (N_9689,N_9599,N_9401);
nand U9690 (N_9690,N_9478,N_9580);
or U9691 (N_9691,N_9591,N_9456);
and U9692 (N_9692,N_9305,N_9416);
or U9693 (N_9693,N_9375,N_9497);
nor U9694 (N_9694,N_9399,N_9464);
nand U9695 (N_9695,N_9520,N_9434);
or U9696 (N_9696,N_9565,N_9451);
and U9697 (N_9697,N_9502,N_9573);
xnor U9698 (N_9698,N_9438,N_9491);
nand U9699 (N_9699,N_9301,N_9348);
nand U9700 (N_9700,N_9372,N_9534);
and U9701 (N_9701,N_9429,N_9546);
nor U9702 (N_9702,N_9433,N_9519);
nor U9703 (N_9703,N_9487,N_9489);
nand U9704 (N_9704,N_9309,N_9364);
xnor U9705 (N_9705,N_9483,N_9562);
nor U9706 (N_9706,N_9501,N_9435);
and U9707 (N_9707,N_9558,N_9446);
nor U9708 (N_9708,N_9358,N_9566);
xor U9709 (N_9709,N_9318,N_9345);
xnor U9710 (N_9710,N_9499,N_9306);
or U9711 (N_9711,N_9586,N_9503);
xor U9712 (N_9712,N_9351,N_9574);
and U9713 (N_9713,N_9369,N_9595);
or U9714 (N_9714,N_9404,N_9418);
nand U9715 (N_9715,N_9425,N_9454);
xor U9716 (N_9716,N_9531,N_9575);
and U9717 (N_9717,N_9445,N_9458);
and U9718 (N_9718,N_9359,N_9347);
and U9719 (N_9719,N_9370,N_9555);
or U9720 (N_9720,N_9410,N_9576);
xor U9721 (N_9721,N_9593,N_9526);
or U9722 (N_9722,N_9444,N_9477);
nand U9723 (N_9723,N_9431,N_9344);
or U9724 (N_9724,N_9362,N_9325);
xor U9725 (N_9725,N_9313,N_9420);
nand U9726 (N_9726,N_9460,N_9469);
or U9727 (N_9727,N_9383,N_9389);
xnor U9728 (N_9728,N_9597,N_9521);
xor U9729 (N_9729,N_9598,N_9350);
xnor U9730 (N_9730,N_9419,N_9380);
or U9731 (N_9731,N_9333,N_9581);
nor U9732 (N_9732,N_9409,N_9496);
nor U9733 (N_9733,N_9390,N_9533);
nand U9734 (N_9734,N_9480,N_9393);
or U9735 (N_9735,N_9381,N_9388);
and U9736 (N_9736,N_9394,N_9462);
and U9737 (N_9737,N_9542,N_9311);
or U9738 (N_9738,N_9583,N_9407);
or U9739 (N_9739,N_9538,N_9396);
xor U9740 (N_9740,N_9336,N_9498);
xor U9741 (N_9741,N_9455,N_9506);
xor U9742 (N_9742,N_9411,N_9449);
nor U9743 (N_9743,N_9564,N_9551);
nand U9744 (N_9744,N_9356,N_9522);
or U9745 (N_9745,N_9437,N_9334);
nor U9746 (N_9746,N_9472,N_9403);
xnor U9747 (N_9747,N_9371,N_9594);
nor U9748 (N_9748,N_9331,N_9550);
nor U9749 (N_9749,N_9500,N_9539);
and U9750 (N_9750,N_9433,N_9476);
nand U9751 (N_9751,N_9434,N_9425);
nor U9752 (N_9752,N_9314,N_9530);
and U9753 (N_9753,N_9304,N_9383);
nand U9754 (N_9754,N_9559,N_9336);
and U9755 (N_9755,N_9483,N_9545);
or U9756 (N_9756,N_9467,N_9400);
and U9757 (N_9757,N_9519,N_9321);
nand U9758 (N_9758,N_9576,N_9474);
xor U9759 (N_9759,N_9535,N_9484);
xor U9760 (N_9760,N_9598,N_9531);
nor U9761 (N_9761,N_9421,N_9561);
or U9762 (N_9762,N_9437,N_9484);
and U9763 (N_9763,N_9412,N_9454);
or U9764 (N_9764,N_9507,N_9387);
and U9765 (N_9765,N_9506,N_9523);
xnor U9766 (N_9766,N_9589,N_9533);
nor U9767 (N_9767,N_9339,N_9323);
or U9768 (N_9768,N_9573,N_9581);
nor U9769 (N_9769,N_9306,N_9517);
nand U9770 (N_9770,N_9414,N_9448);
nor U9771 (N_9771,N_9353,N_9536);
and U9772 (N_9772,N_9405,N_9437);
or U9773 (N_9773,N_9364,N_9315);
nor U9774 (N_9774,N_9463,N_9520);
nand U9775 (N_9775,N_9500,N_9405);
nand U9776 (N_9776,N_9583,N_9448);
xnor U9777 (N_9777,N_9438,N_9414);
or U9778 (N_9778,N_9423,N_9491);
or U9779 (N_9779,N_9455,N_9582);
or U9780 (N_9780,N_9591,N_9491);
and U9781 (N_9781,N_9582,N_9485);
or U9782 (N_9782,N_9469,N_9353);
or U9783 (N_9783,N_9408,N_9588);
xor U9784 (N_9784,N_9478,N_9346);
or U9785 (N_9785,N_9396,N_9489);
nor U9786 (N_9786,N_9455,N_9524);
xor U9787 (N_9787,N_9467,N_9426);
nand U9788 (N_9788,N_9579,N_9362);
or U9789 (N_9789,N_9474,N_9499);
and U9790 (N_9790,N_9346,N_9393);
nand U9791 (N_9791,N_9361,N_9525);
and U9792 (N_9792,N_9541,N_9381);
nor U9793 (N_9793,N_9325,N_9467);
nor U9794 (N_9794,N_9386,N_9504);
nor U9795 (N_9795,N_9339,N_9418);
nor U9796 (N_9796,N_9461,N_9494);
nor U9797 (N_9797,N_9434,N_9543);
nor U9798 (N_9798,N_9527,N_9540);
and U9799 (N_9799,N_9518,N_9593);
xnor U9800 (N_9800,N_9446,N_9414);
and U9801 (N_9801,N_9497,N_9428);
nand U9802 (N_9802,N_9455,N_9471);
and U9803 (N_9803,N_9570,N_9427);
nor U9804 (N_9804,N_9501,N_9528);
or U9805 (N_9805,N_9492,N_9335);
xnor U9806 (N_9806,N_9579,N_9375);
or U9807 (N_9807,N_9504,N_9416);
or U9808 (N_9808,N_9314,N_9488);
nand U9809 (N_9809,N_9569,N_9386);
nand U9810 (N_9810,N_9443,N_9474);
xor U9811 (N_9811,N_9307,N_9315);
or U9812 (N_9812,N_9413,N_9545);
xor U9813 (N_9813,N_9526,N_9388);
xor U9814 (N_9814,N_9586,N_9371);
nand U9815 (N_9815,N_9574,N_9376);
nor U9816 (N_9816,N_9488,N_9593);
nand U9817 (N_9817,N_9342,N_9326);
nor U9818 (N_9818,N_9478,N_9415);
xor U9819 (N_9819,N_9507,N_9530);
nand U9820 (N_9820,N_9319,N_9400);
nand U9821 (N_9821,N_9372,N_9563);
nand U9822 (N_9822,N_9493,N_9548);
or U9823 (N_9823,N_9494,N_9419);
xnor U9824 (N_9824,N_9477,N_9584);
nor U9825 (N_9825,N_9367,N_9532);
nor U9826 (N_9826,N_9509,N_9476);
or U9827 (N_9827,N_9507,N_9554);
and U9828 (N_9828,N_9475,N_9482);
xnor U9829 (N_9829,N_9555,N_9500);
nand U9830 (N_9830,N_9481,N_9572);
xor U9831 (N_9831,N_9427,N_9436);
or U9832 (N_9832,N_9401,N_9349);
and U9833 (N_9833,N_9345,N_9300);
nand U9834 (N_9834,N_9570,N_9598);
xor U9835 (N_9835,N_9413,N_9394);
or U9836 (N_9836,N_9412,N_9451);
nand U9837 (N_9837,N_9511,N_9555);
xor U9838 (N_9838,N_9487,N_9327);
and U9839 (N_9839,N_9436,N_9489);
or U9840 (N_9840,N_9331,N_9407);
and U9841 (N_9841,N_9414,N_9535);
or U9842 (N_9842,N_9589,N_9302);
and U9843 (N_9843,N_9398,N_9547);
and U9844 (N_9844,N_9521,N_9305);
xor U9845 (N_9845,N_9423,N_9529);
nor U9846 (N_9846,N_9536,N_9587);
nor U9847 (N_9847,N_9516,N_9453);
or U9848 (N_9848,N_9544,N_9357);
nand U9849 (N_9849,N_9556,N_9478);
nor U9850 (N_9850,N_9577,N_9450);
or U9851 (N_9851,N_9579,N_9422);
nor U9852 (N_9852,N_9310,N_9337);
or U9853 (N_9853,N_9585,N_9435);
and U9854 (N_9854,N_9599,N_9473);
or U9855 (N_9855,N_9531,N_9317);
nand U9856 (N_9856,N_9354,N_9496);
nand U9857 (N_9857,N_9460,N_9585);
xnor U9858 (N_9858,N_9310,N_9417);
and U9859 (N_9859,N_9456,N_9487);
or U9860 (N_9860,N_9364,N_9496);
nor U9861 (N_9861,N_9475,N_9309);
nand U9862 (N_9862,N_9524,N_9483);
nand U9863 (N_9863,N_9565,N_9401);
nand U9864 (N_9864,N_9457,N_9347);
nand U9865 (N_9865,N_9429,N_9469);
nand U9866 (N_9866,N_9519,N_9431);
and U9867 (N_9867,N_9463,N_9385);
or U9868 (N_9868,N_9510,N_9433);
and U9869 (N_9869,N_9495,N_9445);
nor U9870 (N_9870,N_9383,N_9408);
or U9871 (N_9871,N_9437,N_9326);
and U9872 (N_9872,N_9371,N_9432);
nand U9873 (N_9873,N_9465,N_9568);
and U9874 (N_9874,N_9309,N_9531);
nor U9875 (N_9875,N_9325,N_9373);
nor U9876 (N_9876,N_9498,N_9416);
nand U9877 (N_9877,N_9426,N_9376);
xor U9878 (N_9878,N_9345,N_9535);
or U9879 (N_9879,N_9580,N_9346);
xnor U9880 (N_9880,N_9551,N_9398);
or U9881 (N_9881,N_9528,N_9573);
xor U9882 (N_9882,N_9332,N_9392);
nor U9883 (N_9883,N_9464,N_9523);
and U9884 (N_9884,N_9378,N_9345);
and U9885 (N_9885,N_9364,N_9392);
nand U9886 (N_9886,N_9328,N_9424);
and U9887 (N_9887,N_9379,N_9527);
and U9888 (N_9888,N_9573,N_9454);
or U9889 (N_9889,N_9355,N_9525);
nand U9890 (N_9890,N_9402,N_9319);
nor U9891 (N_9891,N_9572,N_9542);
nor U9892 (N_9892,N_9533,N_9597);
and U9893 (N_9893,N_9326,N_9377);
nor U9894 (N_9894,N_9440,N_9555);
xnor U9895 (N_9895,N_9380,N_9366);
and U9896 (N_9896,N_9538,N_9581);
or U9897 (N_9897,N_9496,N_9590);
xnor U9898 (N_9898,N_9440,N_9356);
nor U9899 (N_9899,N_9328,N_9363);
nand U9900 (N_9900,N_9714,N_9812);
and U9901 (N_9901,N_9640,N_9737);
or U9902 (N_9902,N_9795,N_9825);
nand U9903 (N_9903,N_9843,N_9747);
nand U9904 (N_9904,N_9628,N_9681);
xnor U9905 (N_9905,N_9601,N_9890);
nand U9906 (N_9906,N_9676,N_9644);
nor U9907 (N_9907,N_9767,N_9892);
and U9908 (N_9908,N_9790,N_9648);
nand U9909 (N_9909,N_9606,N_9808);
xor U9910 (N_9910,N_9818,N_9875);
or U9911 (N_9911,N_9746,N_9777);
nand U9912 (N_9912,N_9610,N_9735);
nor U9913 (N_9913,N_9725,N_9871);
and U9914 (N_9914,N_9876,N_9870);
or U9915 (N_9915,N_9752,N_9798);
nand U9916 (N_9916,N_9664,N_9658);
nor U9917 (N_9917,N_9802,N_9809);
nand U9918 (N_9918,N_9683,N_9776);
nand U9919 (N_9919,N_9759,N_9887);
and U9920 (N_9920,N_9667,N_9797);
nor U9921 (N_9921,N_9660,N_9894);
nand U9922 (N_9922,N_9621,N_9671);
and U9923 (N_9923,N_9708,N_9641);
xnor U9924 (N_9924,N_9873,N_9897);
and U9925 (N_9925,N_9693,N_9784);
nand U9926 (N_9926,N_9835,N_9659);
or U9927 (N_9927,N_9764,N_9794);
and U9928 (N_9928,N_9782,N_9884);
nand U9929 (N_9929,N_9856,N_9674);
and U9930 (N_9930,N_9699,N_9789);
nand U9931 (N_9931,N_9896,N_9841);
nand U9932 (N_9932,N_9779,N_9750);
xnor U9933 (N_9933,N_9891,N_9719);
nor U9934 (N_9934,N_9828,N_9619);
or U9935 (N_9935,N_9743,N_9672);
or U9936 (N_9936,N_9801,N_9691);
nand U9937 (N_9937,N_9637,N_9806);
nor U9938 (N_9938,N_9687,N_9861);
nand U9939 (N_9939,N_9663,N_9624);
and U9940 (N_9940,N_9728,N_9744);
nand U9941 (N_9941,N_9718,N_9736);
and U9942 (N_9942,N_9868,N_9854);
nor U9943 (N_9943,N_9689,N_9706);
and U9944 (N_9944,N_9804,N_9785);
and U9945 (N_9945,N_9766,N_9634);
nor U9946 (N_9946,N_9816,N_9688);
nor U9947 (N_9947,N_9635,N_9888);
xnor U9948 (N_9948,N_9652,N_9703);
nor U9949 (N_9949,N_9788,N_9732);
or U9950 (N_9950,N_9778,N_9768);
and U9951 (N_9951,N_9836,N_9690);
or U9952 (N_9952,N_9857,N_9618);
or U9953 (N_9953,N_9839,N_9655);
or U9954 (N_9954,N_9604,N_9696);
nor U9955 (N_9955,N_9882,N_9810);
and U9956 (N_9956,N_9616,N_9864);
and U9957 (N_9957,N_9846,N_9738);
nor U9958 (N_9958,N_9895,N_9883);
nor U9959 (N_9959,N_9880,N_9613);
and U9960 (N_9960,N_9642,N_9682);
nand U9961 (N_9961,N_9726,N_9755);
and U9962 (N_9962,N_9653,N_9731);
and U9963 (N_9963,N_9847,N_9815);
and U9964 (N_9964,N_9614,N_9729);
nor U9965 (N_9965,N_9860,N_9742);
xor U9966 (N_9966,N_9867,N_9826);
nor U9967 (N_9967,N_9851,N_9669);
and U9968 (N_9968,N_9724,N_9677);
xnor U9969 (N_9969,N_9889,N_9739);
nor U9970 (N_9970,N_9684,N_9760);
nand U9971 (N_9971,N_9709,N_9842);
nand U9972 (N_9972,N_9823,N_9863);
nand U9973 (N_9973,N_9771,N_9831);
nor U9974 (N_9974,N_9878,N_9673);
nand U9975 (N_9975,N_9625,N_9770);
xor U9976 (N_9976,N_9898,N_9765);
and U9977 (N_9977,N_9827,N_9602);
nand U9978 (N_9978,N_9694,N_9899);
and U9979 (N_9979,N_9862,N_9881);
and U9980 (N_9980,N_9710,N_9819);
xor U9981 (N_9981,N_9631,N_9603);
nand U9982 (N_9982,N_9865,N_9716);
xnor U9983 (N_9983,N_9748,N_9787);
and U9984 (N_9984,N_9885,N_9645);
xor U9985 (N_9985,N_9668,N_9840);
xor U9986 (N_9986,N_9649,N_9799);
and U9987 (N_9987,N_9791,N_9774);
xnor U9988 (N_9988,N_9639,N_9609);
and U9989 (N_9989,N_9762,N_9707);
or U9990 (N_9990,N_9761,N_9679);
nor U9991 (N_9991,N_9733,N_9830);
xor U9992 (N_9992,N_9866,N_9763);
nor U9993 (N_9993,N_9886,N_9702);
or U9994 (N_9994,N_9833,N_9786);
or U9995 (N_9995,N_9893,N_9852);
nand U9996 (N_9996,N_9656,N_9734);
nor U9997 (N_9997,N_9745,N_9626);
and U9998 (N_9998,N_9607,N_9723);
and U9999 (N_9999,N_9753,N_9695);
nand U10000 (N_10000,N_9838,N_9800);
nor U10001 (N_10001,N_9670,N_9654);
xnor U10002 (N_10002,N_9872,N_9792);
nor U10003 (N_10003,N_9845,N_9803);
nand U10004 (N_10004,N_9629,N_9781);
xnor U10005 (N_10005,N_9713,N_9853);
and U10006 (N_10006,N_9741,N_9675);
and U10007 (N_10007,N_9775,N_9874);
nand U10008 (N_10008,N_9705,N_9615);
or U10009 (N_10009,N_9769,N_9638);
and U10010 (N_10010,N_9751,N_9754);
or U10011 (N_10011,N_9783,N_9643);
nand U10012 (N_10012,N_9849,N_9807);
nand U10013 (N_10013,N_9756,N_9678);
xor U10014 (N_10014,N_9704,N_9855);
and U10015 (N_10015,N_9820,N_9647);
nor U10016 (N_10016,N_9646,N_9686);
and U10017 (N_10017,N_9662,N_9814);
or U10018 (N_10018,N_9692,N_9832);
and U10019 (N_10019,N_9665,N_9834);
nor U10020 (N_10020,N_9793,N_9700);
and U10021 (N_10021,N_9712,N_9869);
nand U10022 (N_10022,N_9605,N_9811);
or U10023 (N_10023,N_9632,N_9617);
or U10024 (N_10024,N_9796,N_9680);
and U10025 (N_10025,N_9630,N_9877);
nor U10026 (N_10026,N_9608,N_9758);
nor U10027 (N_10027,N_9600,N_9721);
xor U10028 (N_10028,N_9685,N_9697);
and U10029 (N_10029,N_9740,N_9717);
xor U10030 (N_10030,N_9715,N_9651);
or U10031 (N_10031,N_9666,N_9701);
nand U10032 (N_10032,N_9879,N_9722);
or U10033 (N_10033,N_9657,N_9773);
nor U10034 (N_10034,N_9620,N_9821);
and U10035 (N_10035,N_9650,N_9859);
nand U10036 (N_10036,N_9749,N_9661);
xor U10037 (N_10037,N_9848,N_9727);
nand U10038 (N_10038,N_9636,N_9720);
nand U10039 (N_10039,N_9623,N_9730);
and U10040 (N_10040,N_9858,N_9612);
nand U10041 (N_10041,N_9780,N_9622);
or U10042 (N_10042,N_9824,N_9829);
xnor U10043 (N_10043,N_9611,N_9627);
or U10044 (N_10044,N_9698,N_9805);
nand U10045 (N_10045,N_9711,N_9813);
or U10046 (N_10046,N_9633,N_9850);
or U10047 (N_10047,N_9757,N_9844);
nand U10048 (N_10048,N_9822,N_9817);
nand U10049 (N_10049,N_9837,N_9772);
xnor U10050 (N_10050,N_9664,N_9766);
or U10051 (N_10051,N_9722,N_9745);
xnor U10052 (N_10052,N_9879,N_9676);
xor U10053 (N_10053,N_9740,N_9685);
xor U10054 (N_10054,N_9644,N_9649);
or U10055 (N_10055,N_9890,N_9876);
and U10056 (N_10056,N_9726,N_9609);
or U10057 (N_10057,N_9641,N_9772);
nor U10058 (N_10058,N_9675,N_9875);
and U10059 (N_10059,N_9664,N_9629);
and U10060 (N_10060,N_9682,N_9895);
xnor U10061 (N_10061,N_9895,N_9824);
or U10062 (N_10062,N_9720,N_9642);
xnor U10063 (N_10063,N_9792,N_9853);
nor U10064 (N_10064,N_9843,N_9632);
or U10065 (N_10065,N_9696,N_9742);
or U10066 (N_10066,N_9823,N_9837);
or U10067 (N_10067,N_9630,N_9881);
and U10068 (N_10068,N_9673,N_9738);
or U10069 (N_10069,N_9780,N_9611);
xor U10070 (N_10070,N_9784,N_9723);
nor U10071 (N_10071,N_9696,N_9844);
nand U10072 (N_10072,N_9735,N_9824);
xnor U10073 (N_10073,N_9640,N_9757);
xnor U10074 (N_10074,N_9889,N_9860);
nor U10075 (N_10075,N_9620,N_9867);
nand U10076 (N_10076,N_9771,N_9858);
nor U10077 (N_10077,N_9791,N_9885);
xor U10078 (N_10078,N_9712,N_9660);
nor U10079 (N_10079,N_9621,N_9741);
and U10080 (N_10080,N_9850,N_9735);
nand U10081 (N_10081,N_9705,N_9617);
nor U10082 (N_10082,N_9896,N_9694);
nand U10083 (N_10083,N_9680,N_9858);
nor U10084 (N_10084,N_9833,N_9868);
or U10085 (N_10085,N_9625,N_9659);
nand U10086 (N_10086,N_9885,N_9733);
nor U10087 (N_10087,N_9706,N_9708);
and U10088 (N_10088,N_9848,N_9887);
nand U10089 (N_10089,N_9654,N_9745);
xor U10090 (N_10090,N_9871,N_9720);
nor U10091 (N_10091,N_9646,N_9645);
or U10092 (N_10092,N_9898,N_9651);
xor U10093 (N_10093,N_9635,N_9624);
xor U10094 (N_10094,N_9627,N_9781);
nor U10095 (N_10095,N_9860,N_9848);
and U10096 (N_10096,N_9782,N_9784);
and U10097 (N_10097,N_9646,N_9680);
and U10098 (N_10098,N_9737,N_9883);
nand U10099 (N_10099,N_9672,N_9884);
and U10100 (N_10100,N_9867,N_9782);
xnor U10101 (N_10101,N_9699,N_9817);
xnor U10102 (N_10102,N_9711,N_9885);
xnor U10103 (N_10103,N_9665,N_9779);
and U10104 (N_10104,N_9729,N_9863);
and U10105 (N_10105,N_9703,N_9694);
xnor U10106 (N_10106,N_9829,N_9731);
nand U10107 (N_10107,N_9793,N_9735);
nand U10108 (N_10108,N_9784,N_9870);
nand U10109 (N_10109,N_9668,N_9706);
and U10110 (N_10110,N_9737,N_9894);
or U10111 (N_10111,N_9863,N_9607);
xor U10112 (N_10112,N_9892,N_9652);
nand U10113 (N_10113,N_9862,N_9833);
nor U10114 (N_10114,N_9867,N_9786);
nor U10115 (N_10115,N_9828,N_9875);
or U10116 (N_10116,N_9654,N_9864);
and U10117 (N_10117,N_9642,N_9691);
xor U10118 (N_10118,N_9732,N_9886);
nor U10119 (N_10119,N_9786,N_9813);
nor U10120 (N_10120,N_9860,N_9809);
or U10121 (N_10121,N_9800,N_9782);
nand U10122 (N_10122,N_9753,N_9616);
nand U10123 (N_10123,N_9888,N_9777);
or U10124 (N_10124,N_9860,N_9792);
nand U10125 (N_10125,N_9623,N_9648);
or U10126 (N_10126,N_9882,N_9802);
nand U10127 (N_10127,N_9777,N_9635);
xnor U10128 (N_10128,N_9740,N_9731);
nor U10129 (N_10129,N_9814,N_9785);
nand U10130 (N_10130,N_9887,N_9869);
xnor U10131 (N_10131,N_9824,N_9683);
xor U10132 (N_10132,N_9761,N_9808);
or U10133 (N_10133,N_9889,N_9817);
nor U10134 (N_10134,N_9671,N_9646);
nor U10135 (N_10135,N_9669,N_9860);
or U10136 (N_10136,N_9619,N_9713);
or U10137 (N_10137,N_9686,N_9639);
or U10138 (N_10138,N_9738,N_9768);
nand U10139 (N_10139,N_9669,N_9786);
xnor U10140 (N_10140,N_9813,N_9721);
xor U10141 (N_10141,N_9819,N_9713);
or U10142 (N_10142,N_9673,N_9841);
and U10143 (N_10143,N_9751,N_9693);
or U10144 (N_10144,N_9660,N_9705);
xor U10145 (N_10145,N_9708,N_9824);
nand U10146 (N_10146,N_9748,N_9819);
nor U10147 (N_10147,N_9701,N_9631);
and U10148 (N_10148,N_9610,N_9817);
xor U10149 (N_10149,N_9698,N_9761);
xnor U10150 (N_10150,N_9766,N_9810);
or U10151 (N_10151,N_9876,N_9821);
or U10152 (N_10152,N_9618,N_9629);
and U10153 (N_10153,N_9855,N_9778);
nand U10154 (N_10154,N_9616,N_9885);
nor U10155 (N_10155,N_9723,N_9793);
xor U10156 (N_10156,N_9655,N_9643);
or U10157 (N_10157,N_9865,N_9860);
nor U10158 (N_10158,N_9726,N_9774);
nand U10159 (N_10159,N_9737,N_9721);
nor U10160 (N_10160,N_9846,N_9783);
xnor U10161 (N_10161,N_9841,N_9729);
xnor U10162 (N_10162,N_9808,N_9723);
or U10163 (N_10163,N_9811,N_9749);
and U10164 (N_10164,N_9833,N_9635);
nand U10165 (N_10165,N_9878,N_9646);
nor U10166 (N_10166,N_9698,N_9709);
xor U10167 (N_10167,N_9640,N_9731);
or U10168 (N_10168,N_9771,N_9843);
and U10169 (N_10169,N_9884,N_9895);
xor U10170 (N_10170,N_9672,N_9608);
nand U10171 (N_10171,N_9899,N_9852);
or U10172 (N_10172,N_9846,N_9744);
or U10173 (N_10173,N_9696,N_9694);
nand U10174 (N_10174,N_9774,N_9636);
nor U10175 (N_10175,N_9737,N_9634);
nor U10176 (N_10176,N_9610,N_9836);
or U10177 (N_10177,N_9756,N_9884);
and U10178 (N_10178,N_9625,N_9824);
nand U10179 (N_10179,N_9806,N_9785);
xnor U10180 (N_10180,N_9833,N_9893);
nor U10181 (N_10181,N_9684,N_9728);
and U10182 (N_10182,N_9810,N_9867);
or U10183 (N_10183,N_9679,N_9772);
xor U10184 (N_10184,N_9605,N_9601);
or U10185 (N_10185,N_9729,N_9776);
and U10186 (N_10186,N_9873,N_9722);
nand U10187 (N_10187,N_9659,N_9710);
nor U10188 (N_10188,N_9634,N_9806);
nor U10189 (N_10189,N_9617,N_9766);
nand U10190 (N_10190,N_9776,N_9845);
xnor U10191 (N_10191,N_9852,N_9641);
nand U10192 (N_10192,N_9642,N_9801);
or U10193 (N_10193,N_9760,N_9846);
nand U10194 (N_10194,N_9780,N_9615);
or U10195 (N_10195,N_9687,N_9849);
nand U10196 (N_10196,N_9679,N_9715);
nor U10197 (N_10197,N_9607,N_9691);
and U10198 (N_10198,N_9649,N_9781);
xor U10199 (N_10199,N_9696,N_9827);
xor U10200 (N_10200,N_10091,N_10001);
xor U10201 (N_10201,N_10012,N_10197);
or U10202 (N_10202,N_10045,N_10006);
xnor U10203 (N_10203,N_9917,N_9951);
and U10204 (N_10204,N_9944,N_10025);
nor U10205 (N_10205,N_10163,N_10073);
or U10206 (N_10206,N_10058,N_10008);
nor U10207 (N_10207,N_9949,N_10120);
nand U10208 (N_10208,N_9931,N_9952);
nor U10209 (N_10209,N_9909,N_9982);
nand U10210 (N_10210,N_9942,N_10139);
xnor U10211 (N_10211,N_10005,N_9995);
and U10212 (N_10212,N_9924,N_9900);
or U10213 (N_10213,N_10019,N_10127);
nor U10214 (N_10214,N_10157,N_10070);
and U10215 (N_10215,N_10093,N_10056);
xor U10216 (N_10216,N_9934,N_10021);
nor U10217 (N_10217,N_10052,N_9910);
and U10218 (N_10218,N_10123,N_9969);
nor U10219 (N_10219,N_10145,N_9946);
xor U10220 (N_10220,N_10102,N_10071);
nand U10221 (N_10221,N_9928,N_10116);
nor U10222 (N_10222,N_10167,N_10015);
xnor U10223 (N_10223,N_10097,N_9906);
or U10224 (N_10224,N_9962,N_10039);
nor U10225 (N_10225,N_10114,N_10151);
or U10226 (N_10226,N_10180,N_10053);
nor U10227 (N_10227,N_10110,N_9943);
nand U10228 (N_10228,N_10168,N_10169);
or U10229 (N_10229,N_9959,N_9978);
nor U10230 (N_10230,N_9976,N_9945);
nand U10231 (N_10231,N_9994,N_10105);
or U10232 (N_10232,N_9972,N_10095);
nor U10233 (N_10233,N_9991,N_9923);
nand U10234 (N_10234,N_9912,N_10074);
xor U10235 (N_10235,N_10107,N_9974);
nor U10236 (N_10236,N_9993,N_9935);
or U10237 (N_10237,N_10164,N_10049);
nor U10238 (N_10238,N_9913,N_9921);
xor U10239 (N_10239,N_9967,N_9905);
nand U10240 (N_10240,N_10031,N_10106);
nand U10241 (N_10241,N_10065,N_9973);
xnor U10242 (N_10242,N_10124,N_10193);
nand U10243 (N_10243,N_10147,N_10111);
or U10244 (N_10244,N_10038,N_10051);
nand U10245 (N_10245,N_9997,N_10148);
nor U10246 (N_10246,N_9960,N_9987);
xor U10247 (N_10247,N_10166,N_10190);
or U10248 (N_10248,N_10143,N_9933);
and U10249 (N_10249,N_10122,N_9941);
nor U10250 (N_10250,N_10017,N_10196);
nor U10251 (N_10251,N_10077,N_10081);
nand U10252 (N_10252,N_10035,N_10119);
and U10253 (N_10253,N_10092,N_9954);
or U10254 (N_10254,N_10027,N_9992);
nand U10255 (N_10255,N_10162,N_9939);
xnor U10256 (N_10256,N_10068,N_10054);
nand U10257 (N_10257,N_10156,N_10032);
and U10258 (N_10258,N_10055,N_10075);
or U10259 (N_10259,N_9957,N_10048);
and U10260 (N_10260,N_9926,N_10087);
or U10261 (N_10261,N_10041,N_9965);
xnor U10262 (N_10262,N_10125,N_10189);
xor U10263 (N_10263,N_10104,N_10140);
nor U10264 (N_10264,N_9985,N_10018);
or U10265 (N_10265,N_10130,N_10069);
and U10266 (N_10266,N_10170,N_10113);
nand U10267 (N_10267,N_9983,N_10150);
xnor U10268 (N_10268,N_10137,N_10061);
or U10269 (N_10269,N_9970,N_10103);
nor U10270 (N_10270,N_9966,N_10072);
or U10271 (N_10271,N_10090,N_9927);
nor U10272 (N_10272,N_10129,N_9968);
xor U10273 (N_10273,N_10101,N_9908);
nor U10274 (N_10274,N_10036,N_9902);
and U10275 (N_10275,N_10179,N_10082);
nor U10276 (N_10276,N_10152,N_10043);
xor U10277 (N_10277,N_10172,N_10154);
nand U10278 (N_10278,N_10040,N_10014);
nor U10279 (N_10279,N_10086,N_10030);
nand U10280 (N_10280,N_9990,N_10044);
or U10281 (N_10281,N_10013,N_10080);
and U10282 (N_10282,N_10046,N_9989);
nand U10283 (N_10283,N_9963,N_10033);
nand U10284 (N_10284,N_10178,N_9940);
or U10285 (N_10285,N_9929,N_10159);
nand U10286 (N_10286,N_9947,N_10171);
and U10287 (N_10287,N_10134,N_10112);
or U10288 (N_10288,N_9977,N_10192);
and U10289 (N_10289,N_10126,N_10182);
nor U10290 (N_10290,N_9937,N_10083);
nor U10291 (N_10291,N_9914,N_10108);
and U10292 (N_10292,N_10181,N_10003);
nor U10293 (N_10293,N_9903,N_10047);
or U10294 (N_10294,N_10175,N_10177);
xnor U10295 (N_10295,N_10089,N_10016);
and U10296 (N_10296,N_9955,N_10009);
and U10297 (N_10297,N_10060,N_9918);
and U10298 (N_10298,N_10026,N_9920);
nor U10299 (N_10299,N_10117,N_9980);
nor U10300 (N_10300,N_10199,N_10155);
nand U10301 (N_10301,N_9936,N_10165);
nor U10302 (N_10302,N_9953,N_9916);
and U10303 (N_10303,N_9938,N_10142);
or U10304 (N_10304,N_9988,N_10098);
or U10305 (N_10305,N_10088,N_10100);
xor U10306 (N_10306,N_10128,N_10188);
xor U10307 (N_10307,N_10131,N_10133);
nor U10308 (N_10308,N_10138,N_10161);
xnor U10309 (N_10309,N_9911,N_10062);
and U10310 (N_10310,N_10174,N_10085);
nor U10311 (N_10311,N_10136,N_10160);
xor U10312 (N_10312,N_10198,N_9958);
or U10313 (N_10313,N_10004,N_9981);
and U10314 (N_10314,N_9979,N_9904);
or U10315 (N_10315,N_10066,N_10132);
or U10316 (N_10316,N_10029,N_10135);
nand U10317 (N_10317,N_9956,N_10076);
and U10318 (N_10318,N_10050,N_9948);
nand U10319 (N_10319,N_9986,N_10141);
nor U10320 (N_10320,N_10010,N_9901);
nor U10321 (N_10321,N_10195,N_9930);
xor U10322 (N_10322,N_10185,N_10024);
or U10323 (N_10323,N_10064,N_9961);
nor U10324 (N_10324,N_10037,N_10118);
nand U10325 (N_10325,N_10191,N_10067);
and U10326 (N_10326,N_9915,N_10022);
and U10327 (N_10327,N_10079,N_9971);
xor U10328 (N_10328,N_10078,N_10096);
nand U10329 (N_10329,N_9964,N_10184);
and U10330 (N_10330,N_10028,N_10187);
xor U10331 (N_10331,N_10042,N_10176);
and U10332 (N_10332,N_9922,N_10057);
or U10333 (N_10333,N_9998,N_10194);
xor U10334 (N_10334,N_10007,N_9950);
and U10335 (N_10335,N_9919,N_10109);
and U10336 (N_10336,N_10153,N_10173);
xnor U10337 (N_10337,N_10186,N_10121);
nor U10338 (N_10338,N_10000,N_10149);
nor U10339 (N_10339,N_9925,N_10099);
and U10340 (N_10340,N_10146,N_10059);
nor U10341 (N_10341,N_9999,N_10144);
and U10342 (N_10342,N_10020,N_10034);
xor U10343 (N_10343,N_9907,N_10183);
nand U10344 (N_10344,N_9984,N_10023);
xor U10345 (N_10345,N_9932,N_10115);
xnor U10346 (N_10346,N_9996,N_10158);
nand U10347 (N_10347,N_10002,N_10094);
nand U10348 (N_10348,N_10063,N_10011);
and U10349 (N_10349,N_9975,N_10084);
nor U10350 (N_10350,N_10049,N_9945);
xor U10351 (N_10351,N_9916,N_10064);
or U10352 (N_10352,N_9952,N_10086);
or U10353 (N_10353,N_10041,N_10157);
and U10354 (N_10354,N_10004,N_10110);
nand U10355 (N_10355,N_9984,N_10096);
xnor U10356 (N_10356,N_9940,N_10042);
and U10357 (N_10357,N_10170,N_10156);
and U10358 (N_10358,N_9993,N_10081);
and U10359 (N_10359,N_10170,N_10153);
or U10360 (N_10360,N_9938,N_9952);
nand U10361 (N_10361,N_10075,N_10193);
nand U10362 (N_10362,N_9911,N_10066);
xor U10363 (N_10363,N_10102,N_10064);
xnor U10364 (N_10364,N_9952,N_10016);
xor U10365 (N_10365,N_10191,N_10062);
nand U10366 (N_10366,N_10074,N_10167);
xor U10367 (N_10367,N_10034,N_10156);
nand U10368 (N_10368,N_10159,N_10119);
nor U10369 (N_10369,N_9972,N_9915);
nand U10370 (N_10370,N_9946,N_9940);
or U10371 (N_10371,N_10154,N_9956);
xor U10372 (N_10372,N_10188,N_10145);
or U10373 (N_10373,N_10156,N_10188);
or U10374 (N_10374,N_10179,N_9966);
or U10375 (N_10375,N_9941,N_10173);
xnor U10376 (N_10376,N_10182,N_10098);
nand U10377 (N_10377,N_10094,N_10131);
and U10378 (N_10378,N_10066,N_10134);
xor U10379 (N_10379,N_10062,N_10196);
and U10380 (N_10380,N_10175,N_10055);
and U10381 (N_10381,N_9957,N_9987);
nand U10382 (N_10382,N_10084,N_9955);
or U10383 (N_10383,N_10109,N_10010);
xnor U10384 (N_10384,N_10119,N_9952);
nor U10385 (N_10385,N_10151,N_10055);
or U10386 (N_10386,N_10129,N_9902);
nor U10387 (N_10387,N_9958,N_10053);
nand U10388 (N_10388,N_10110,N_9988);
xnor U10389 (N_10389,N_10023,N_9975);
or U10390 (N_10390,N_9991,N_9901);
nand U10391 (N_10391,N_10190,N_10015);
nor U10392 (N_10392,N_10071,N_9963);
or U10393 (N_10393,N_9989,N_10141);
nor U10394 (N_10394,N_10170,N_10044);
nand U10395 (N_10395,N_9971,N_9984);
or U10396 (N_10396,N_10144,N_9988);
or U10397 (N_10397,N_10134,N_10118);
nor U10398 (N_10398,N_10007,N_10064);
nand U10399 (N_10399,N_10054,N_9914);
nor U10400 (N_10400,N_10042,N_10128);
xnor U10401 (N_10401,N_10102,N_10138);
or U10402 (N_10402,N_10022,N_10110);
and U10403 (N_10403,N_10034,N_10196);
nand U10404 (N_10404,N_10050,N_9996);
nand U10405 (N_10405,N_9979,N_9917);
nor U10406 (N_10406,N_9905,N_10134);
nand U10407 (N_10407,N_10084,N_9978);
nor U10408 (N_10408,N_10127,N_10186);
nor U10409 (N_10409,N_10193,N_10125);
nand U10410 (N_10410,N_10039,N_9974);
xnor U10411 (N_10411,N_10054,N_10009);
xnor U10412 (N_10412,N_10070,N_10160);
nor U10413 (N_10413,N_9910,N_9911);
nand U10414 (N_10414,N_10069,N_9923);
xor U10415 (N_10415,N_9994,N_10083);
or U10416 (N_10416,N_10012,N_10027);
nor U10417 (N_10417,N_10100,N_10057);
or U10418 (N_10418,N_9978,N_10067);
nand U10419 (N_10419,N_10146,N_10176);
nor U10420 (N_10420,N_9916,N_9906);
nand U10421 (N_10421,N_10045,N_10075);
nor U10422 (N_10422,N_10082,N_9971);
nand U10423 (N_10423,N_9937,N_9935);
or U10424 (N_10424,N_10072,N_9968);
xnor U10425 (N_10425,N_9973,N_9980);
xor U10426 (N_10426,N_10033,N_10037);
or U10427 (N_10427,N_9960,N_10029);
nand U10428 (N_10428,N_10137,N_9901);
or U10429 (N_10429,N_9949,N_9939);
nor U10430 (N_10430,N_9941,N_10046);
and U10431 (N_10431,N_9999,N_10141);
nand U10432 (N_10432,N_10042,N_10131);
nor U10433 (N_10433,N_9980,N_9941);
nand U10434 (N_10434,N_10025,N_10183);
nand U10435 (N_10435,N_10190,N_9964);
or U10436 (N_10436,N_10088,N_10189);
nor U10437 (N_10437,N_10132,N_10045);
xnor U10438 (N_10438,N_10000,N_10088);
nand U10439 (N_10439,N_9957,N_10185);
and U10440 (N_10440,N_9955,N_9957);
xnor U10441 (N_10441,N_9924,N_10083);
and U10442 (N_10442,N_9978,N_10055);
xnor U10443 (N_10443,N_9936,N_10071);
nor U10444 (N_10444,N_10004,N_10192);
and U10445 (N_10445,N_9918,N_10187);
and U10446 (N_10446,N_10061,N_9986);
nand U10447 (N_10447,N_10171,N_10133);
or U10448 (N_10448,N_10114,N_10091);
or U10449 (N_10449,N_10153,N_9950);
xnor U10450 (N_10450,N_9958,N_9956);
nor U10451 (N_10451,N_10192,N_10172);
or U10452 (N_10452,N_10060,N_9941);
xnor U10453 (N_10453,N_9953,N_10005);
nor U10454 (N_10454,N_10077,N_10026);
or U10455 (N_10455,N_10007,N_10144);
xor U10456 (N_10456,N_9980,N_10189);
nor U10457 (N_10457,N_9940,N_9983);
nor U10458 (N_10458,N_9970,N_10075);
or U10459 (N_10459,N_10096,N_10006);
and U10460 (N_10460,N_10123,N_10044);
and U10461 (N_10461,N_9938,N_10130);
nor U10462 (N_10462,N_10106,N_10007);
xnor U10463 (N_10463,N_10072,N_9905);
nand U10464 (N_10464,N_10106,N_10126);
xnor U10465 (N_10465,N_9948,N_10192);
or U10466 (N_10466,N_9916,N_9968);
nand U10467 (N_10467,N_10122,N_9982);
or U10468 (N_10468,N_9946,N_9972);
nor U10469 (N_10469,N_10174,N_9903);
and U10470 (N_10470,N_9966,N_10136);
and U10471 (N_10471,N_9951,N_10116);
or U10472 (N_10472,N_9924,N_10183);
nor U10473 (N_10473,N_9912,N_9944);
nand U10474 (N_10474,N_10182,N_9935);
and U10475 (N_10475,N_9923,N_9997);
and U10476 (N_10476,N_9932,N_9926);
nand U10477 (N_10477,N_9930,N_9982);
or U10478 (N_10478,N_10149,N_10090);
xor U10479 (N_10479,N_10085,N_9981);
nand U10480 (N_10480,N_10142,N_10189);
xnor U10481 (N_10481,N_10126,N_9963);
nor U10482 (N_10482,N_9903,N_10067);
nand U10483 (N_10483,N_10106,N_10122);
nor U10484 (N_10484,N_10027,N_10153);
and U10485 (N_10485,N_9976,N_10120);
nor U10486 (N_10486,N_9919,N_10120);
nor U10487 (N_10487,N_9962,N_9923);
nand U10488 (N_10488,N_9916,N_9948);
xnor U10489 (N_10489,N_9934,N_10106);
nand U10490 (N_10490,N_10068,N_9921);
or U10491 (N_10491,N_10082,N_9953);
xor U10492 (N_10492,N_10035,N_10062);
and U10493 (N_10493,N_10119,N_9917);
nor U10494 (N_10494,N_9903,N_9927);
xor U10495 (N_10495,N_10169,N_10118);
or U10496 (N_10496,N_10156,N_9951);
or U10497 (N_10497,N_9968,N_10059);
nor U10498 (N_10498,N_10005,N_10146);
or U10499 (N_10499,N_9933,N_10150);
or U10500 (N_10500,N_10311,N_10309);
xor U10501 (N_10501,N_10448,N_10455);
xor U10502 (N_10502,N_10253,N_10355);
or U10503 (N_10503,N_10271,N_10431);
xor U10504 (N_10504,N_10449,N_10492);
or U10505 (N_10505,N_10342,N_10478);
xnor U10506 (N_10506,N_10328,N_10351);
or U10507 (N_10507,N_10273,N_10307);
or U10508 (N_10508,N_10376,N_10456);
nor U10509 (N_10509,N_10274,N_10496);
nor U10510 (N_10510,N_10494,N_10319);
xor U10511 (N_10511,N_10247,N_10336);
and U10512 (N_10512,N_10285,N_10383);
nor U10513 (N_10513,N_10231,N_10256);
and U10514 (N_10514,N_10405,N_10220);
nor U10515 (N_10515,N_10244,N_10467);
or U10516 (N_10516,N_10201,N_10210);
xnor U10517 (N_10517,N_10344,N_10400);
nor U10518 (N_10518,N_10228,N_10442);
xor U10519 (N_10519,N_10391,N_10491);
nand U10520 (N_10520,N_10499,N_10402);
or U10521 (N_10521,N_10332,N_10277);
and U10522 (N_10522,N_10464,N_10430);
xor U10523 (N_10523,N_10421,N_10425);
and U10524 (N_10524,N_10289,N_10334);
and U10525 (N_10525,N_10267,N_10323);
and U10526 (N_10526,N_10490,N_10399);
nand U10527 (N_10527,N_10294,N_10313);
nor U10528 (N_10528,N_10322,N_10394);
or U10529 (N_10529,N_10325,N_10475);
or U10530 (N_10530,N_10388,N_10411);
and U10531 (N_10531,N_10296,N_10374);
nand U10532 (N_10532,N_10485,N_10292);
nor U10533 (N_10533,N_10415,N_10324);
and U10534 (N_10534,N_10329,N_10315);
or U10535 (N_10535,N_10233,N_10424);
xor U10536 (N_10536,N_10214,N_10356);
and U10537 (N_10537,N_10377,N_10218);
or U10538 (N_10538,N_10270,N_10412);
xor U10539 (N_10539,N_10216,N_10452);
or U10540 (N_10540,N_10348,N_10436);
or U10541 (N_10541,N_10359,N_10386);
and U10542 (N_10542,N_10206,N_10275);
nor U10543 (N_10543,N_10462,N_10339);
xor U10544 (N_10544,N_10236,N_10444);
nor U10545 (N_10545,N_10282,N_10370);
nand U10546 (N_10546,N_10230,N_10409);
or U10547 (N_10547,N_10246,N_10366);
xnor U10548 (N_10548,N_10487,N_10213);
or U10549 (N_10549,N_10426,N_10476);
or U10550 (N_10550,N_10299,N_10480);
xor U10551 (N_10551,N_10353,N_10447);
or U10552 (N_10552,N_10343,N_10495);
xnor U10553 (N_10553,N_10207,N_10333);
nand U10554 (N_10554,N_10408,N_10357);
or U10555 (N_10555,N_10440,N_10390);
and U10556 (N_10556,N_10465,N_10489);
or U10557 (N_10557,N_10468,N_10382);
or U10558 (N_10558,N_10364,N_10417);
nor U10559 (N_10559,N_10419,N_10251);
xor U10560 (N_10560,N_10439,N_10320);
xnor U10561 (N_10561,N_10349,N_10397);
or U10562 (N_10562,N_10385,N_10212);
nand U10563 (N_10563,N_10293,N_10261);
nand U10564 (N_10564,N_10451,N_10471);
and U10565 (N_10565,N_10279,N_10316);
nand U10566 (N_10566,N_10393,N_10284);
and U10567 (N_10567,N_10254,N_10262);
or U10568 (N_10568,N_10317,N_10243);
or U10569 (N_10569,N_10486,N_10245);
nand U10570 (N_10570,N_10330,N_10407);
or U10571 (N_10571,N_10276,N_10379);
xor U10572 (N_10572,N_10392,N_10454);
xnor U10573 (N_10573,N_10497,N_10290);
nor U10574 (N_10574,N_10410,N_10481);
nand U10575 (N_10575,N_10266,N_10389);
nor U10576 (N_10576,N_10403,N_10484);
nor U10577 (N_10577,N_10314,N_10373);
nand U10578 (N_10578,N_10345,N_10252);
nand U10579 (N_10579,N_10446,N_10380);
and U10580 (N_10580,N_10362,N_10225);
xor U10581 (N_10581,N_10286,N_10422);
or U10582 (N_10582,N_10209,N_10378);
nor U10583 (N_10583,N_10466,N_10205);
xnor U10584 (N_10584,N_10321,N_10308);
or U10585 (N_10585,N_10303,N_10268);
and U10586 (N_10586,N_10420,N_10483);
and U10587 (N_10587,N_10260,N_10239);
nand U10588 (N_10588,N_10472,N_10375);
and U10589 (N_10589,N_10208,N_10288);
and U10590 (N_10590,N_10404,N_10200);
or U10591 (N_10591,N_10429,N_10217);
nor U10592 (N_10592,N_10250,N_10264);
and U10593 (N_10593,N_10300,N_10283);
and U10594 (N_10594,N_10224,N_10482);
and U10595 (N_10595,N_10287,N_10346);
or U10596 (N_10596,N_10443,N_10398);
or U10597 (N_10597,N_10435,N_10418);
nor U10598 (N_10598,N_10368,N_10453);
xor U10599 (N_10599,N_10434,N_10202);
or U10600 (N_10600,N_10406,N_10413);
xor U10601 (N_10601,N_10432,N_10326);
nand U10602 (N_10602,N_10469,N_10416);
or U10603 (N_10603,N_10445,N_10427);
or U10604 (N_10604,N_10441,N_10360);
nand U10605 (N_10605,N_10257,N_10477);
nor U10606 (N_10606,N_10396,N_10304);
xor U10607 (N_10607,N_10338,N_10352);
and U10608 (N_10608,N_10365,N_10211);
nor U10609 (N_10609,N_10450,N_10291);
nor U10610 (N_10610,N_10222,N_10414);
xnor U10611 (N_10611,N_10318,N_10423);
nor U10612 (N_10612,N_10371,N_10235);
nor U10613 (N_10613,N_10226,N_10305);
nor U10614 (N_10614,N_10363,N_10203);
nand U10615 (N_10615,N_10259,N_10306);
nand U10616 (N_10616,N_10258,N_10437);
and U10617 (N_10617,N_10459,N_10301);
nand U10618 (N_10618,N_10479,N_10241);
xor U10619 (N_10619,N_10237,N_10215);
nor U10620 (N_10620,N_10229,N_10238);
or U10621 (N_10621,N_10310,N_10265);
or U10622 (N_10622,N_10221,N_10438);
nand U10623 (N_10623,N_10249,N_10204);
nor U10624 (N_10624,N_10281,N_10369);
nor U10625 (N_10625,N_10234,N_10474);
nand U10626 (N_10626,N_10387,N_10297);
nand U10627 (N_10627,N_10347,N_10428);
nor U10628 (N_10628,N_10401,N_10223);
xor U10629 (N_10629,N_10255,N_10473);
or U10630 (N_10630,N_10498,N_10337);
xor U10631 (N_10631,N_10272,N_10248);
nor U10632 (N_10632,N_10263,N_10470);
or U10633 (N_10633,N_10350,N_10372);
and U10634 (N_10634,N_10327,N_10461);
xnor U10635 (N_10635,N_10463,N_10457);
nor U10636 (N_10636,N_10340,N_10227);
xor U10637 (N_10637,N_10395,N_10295);
or U10638 (N_10638,N_10433,N_10381);
or U10639 (N_10639,N_10240,N_10361);
nand U10640 (N_10640,N_10488,N_10298);
and U10641 (N_10641,N_10242,N_10493);
nor U10642 (N_10642,N_10312,N_10358);
nand U10643 (N_10643,N_10219,N_10460);
and U10644 (N_10644,N_10341,N_10367);
xnor U10645 (N_10645,N_10335,N_10280);
nor U10646 (N_10646,N_10278,N_10302);
nand U10647 (N_10647,N_10384,N_10354);
xor U10648 (N_10648,N_10331,N_10232);
nor U10649 (N_10649,N_10458,N_10269);
xor U10650 (N_10650,N_10276,N_10439);
xor U10651 (N_10651,N_10267,N_10343);
nand U10652 (N_10652,N_10472,N_10254);
nor U10653 (N_10653,N_10377,N_10330);
xnor U10654 (N_10654,N_10225,N_10204);
and U10655 (N_10655,N_10415,N_10207);
and U10656 (N_10656,N_10446,N_10228);
or U10657 (N_10657,N_10271,N_10263);
or U10658 (N_10658,N_10304,N_10488);
nor U10659 (N_10659,N_10455,N_10254);
or U10660 (N_10660,N_10253,N_10444);
or U10661 (N_10661,N_10330,N_10308);
xor U10662 (N_10662,N_10464,N_10221);
xor U10663 (N_10663,N_10268,N_10326);
or U10664 (N_10664,N_10208,N_10235);
or U10665 (N_10665,N_10438,N_10414);
and U10666 (N_10666,N_10316,N_10203);
and U10667 (N_10667,N_10308,N_10215);
xor U10668 (N_10668,N_10317,N_10255);
xor U10669 (N_10669,N_10494,N_10477);
xor U10670 (N_10670,N_10387,N_10494);
xor U10671 (N_10671,N_10486,N_10417);
or U10672 (N_10672,N_10312,N_10369);
or U10673 (N_10673,N_10436,N_10318);
nor U10674 (N_10674,N_10241,N_10288);
and U10675 (N_10675,N_10482,N_10294);
nor U10676 (N_10676,N_10442,N_10475);
or U10677 (N_10677,N_10267,N_10334);
nor U10678 (N_10678,N_10498,N_10365);
nand U10679 (N_10679,N_10288,N_10375);
or U10680 (N_10680,N_10386,N_10478);
xor U10681 (N_10681,N_10264,N_10497);
xnor U10682 (N_10682,N_10232,N_10304);
nor U10683 (N_10683,N_10425,N_10405);
nor U10684 (N_10684,N_10335,N_10370);
and U10685 (N_10685,N_10467,N_10493);
and U10686 (N_10686,N_10275,N_10366);
or U10687 (N_10687,N_10298,N_10409);
nor U10688 (N_10688,N_10213,N_10440);
nor U10689 (N_10689,N_10224,N_10401);
nand U10690 (N_10690,N_10368,N_10261);
or U10691 (N_10691,N_10484,N_10293);
xnor U10692 (N_10692,N_10465,N_10258);
and U10693 (N_10693,N_10406,N_10211);
nor U10694 (N_10694,N_10465,N_10438);
or U10695 (N_10695,N_10388,N_10256);
and U10696 (N_10696,N_10444,N_10458);
xor U10697 (N_10697,N_10262,N_10289);
xnor U10698 (N_10698,N_10491,N_10433);
xnor U10699 (N_10699,N_10371,N_10495);
nand U10700 (N_10700,N_10361,N_10325);
nand U10701 (N_10701,N_10471,N_10291);
xnor U10702 (N_10702,N_10264,N_10427);
nor U10703 (N_10703,N_10467,N_10250);
and U10704 (N_10704,N_10285,N_10432);
or U10705 (N_10705,N_10355,N_10323);
xnor U10706 (N_10706,N_10415,N_10310);
nand U10707 (N_10707,N_10438,N_10394);
xor U10708 (N_10708,N_10292,N_10309);
or U10709 (N_10709,N_10363,N_10213);
nor U10710 (N_10710,N_10247,N_10433);
nand U10711 (N_10711,N_10390,N_10224);
and U10712 (N_10712,N_10267,N_10358);
nand U10713 (N_10713,N_10334,N_10331);
nor U10714 (N_10714,N_10376,N_10291);
and U10715 (N_10715,N_10231,N_10330);
and U10716 (N_10716,N_10468,N_10457);
or U10717 (N_10717,N_10486,N_10243);
and U10718 (N_10718,N_10324,N_10200);
xnor U10719 (N_10719,N_10377,N_10312);
xor U10720 (N_10720,N_10294,N_10353);
and U10721 (N_10721,N_10211,N_10356);
and U10722 (N_10722,N_10263,N_10498);
nor U10723 (N_10723,N_10473,N_10459);
and U10724 (N_10724,N_10387,N_10473);
or U10725 (N_10725,N_10297,N_10351);
nor U10726 (N_10726,N_10416,N_10438);
and U10727 (N_10727,N_10223,N_10422);
nor U10728 (N_10728,N_10450,N_10485);
nand U10729 (N_10729,N_10441,N_10420);
nor U10730 (N_10730,N_10356,N_10245);
nor U10731 (N_10731,N_10312,N_10359);
xor U10732 (N_10732,N_10437,N_10428);
or U10733 (N_10733,N_10273,N_10441);
nor U10734 (N_10734,N_10417,N_10344);
or U10735 (N_10735,N_10302,N_10386);
and U10736 (N_10736,N_10263,N_10245);
and U10737 (N_10737,N_10477,N_10366);
or U10738 (N_10738,N_10416,N_10289);
nor U10739 (N_10739,N_10460,N_10499);
or U10740 (N_10740,N_10218,N_10336);
nand U10741 (N_10741,N_10450,N_10341);
nor U10742 (N_10742,N_10420,N_10279);
or U10743 (N_10743,N_10235,N_10237);
nand U10744 (N_10744,N_10429,N_10301);
and U10745 (N_10745,N_10427,N_10288);
or U10746 (N_10746,N_10377,N_10406);
and U10747 (N_10747,N_10228,N_10351);
and U10748 (N_10748,N_10454,N_10206);
or U10749 (N_10749,N_10305,N_10265);
or U10750 (N_10750,N_10299,N_10377);
xnor U10751 (N_10751,N_10484,N_10318);
xnor U10752 (N_10752,N_10231,N_10324);
nand U10753 (N_10753,N_10405,N_10257);
nor U10754 (N_10754,N_10424,N_10349);
nor U10755 (N_10755,N_10357,N_10272);
nand U10756 (N_10756,N_10358,N_10266);
nand U10757 (N_10757,N_10420,N_10260);
or U10758 (N_10758,N_10489,N_10205);
or U10759 (N_10759,N_10261,N_10403);
nor U10760 (N_10760,N_10413,N_10489);
or U10761 (N_10761,N_10305,N_10423);
or U10762 (N_10762,N_10489,N_10337);
or U10763 (N_10763,N_10401,N_10290);
nand U10764 (N_10764,N_10431,N_10393);
and U10765 (N_10765,N_10345,N_10492);
and U10766 (N_10766,N_10306,N_10239);
xor U10767 (N_10767,N_10421,N_10403);
nand U10768 (N_10768,N_10207,N_10284);
xor U10769 (N_10769,N_10353,N_10367);
or U10770 (N_10770,N_10344,N_10406);
xor U10771 (N_10771,N_10218,N_10493);
nor U10772 (N_10772,N_10329,N_10366);
nand U10773 (N_10773,N_10417,N_10389);
xnor U10774 (N_10774,N_10497,N_10492);
and U10775 (N_10775,N_10278,N_10444);
and U10776 (N_10776,N_10439,N_10286);
nor U10777 (N_10777,N_10211,N_10355);
nor U10778 (N_10778,N_10356,N_10406);
nor U10779 (N_10779,N_10306,N_10491);
nor U10780 (N_10780,N_10451,N_10499);
nand U10781 (N_10781,N_10431,N_10312);
nand U10782 (N_10782,N_10233,N_10282);
nand U10783 (N_10783,N_10245,N_10320);
nand U10784 (N_10784,N_10299,N_10350);
xnor U10785 (N_10785,N_10453,N_10379);
or U10786 (N_10786,N_10201,N_10489);
or U10787 (N_10787,N_10487,N_10463);
xor U10788 (N_10788,N_10374,N_10221);
and U10789 (N_10789,N_10224,N_10245);
nand U10790 (N_10790,N_10432,N_10477);
nand U10791 (N_10791,N_10470,N_10415);
nand U10792 (N_10792,N_10436,N_10371);
xor U10793 (N_10793,N_10476,N_10275);
or U10794 (N_10794,N_10263,N_10401);
xor U10795 (N_10795,N_10305,N_10457);
and U10796 (N_10796,N_10201,N_10374);
or U10797 (N_10797,N_10237,N_10403);
nor U10798 (N_10798,N_10418,N_10457);
xor U10799 (N_10799,N_10396,N_10231);
nor U10800 (N_10800,N_10621,N_10548);
and U10801 (N_10801,N_10601,N_10637);
nor U10802 (N_10802,N_10654,N_10571);
and U10803 (N_10803,N_10522,N_10638);
or U10804 (N_10804,N_10515,N_10795);
nand U10805 (N_10805,N_10725,N_10681);
nand U10806 (N_10806,N_10784,N_10516);
nor U10807 (N_10807,N_10652,N_10689);
or U10808 (N_10808,N_10728,N_10657);
xor U10809 (N_10809,N_10500,N_10574);
nand U10810 (N_10810,N_10760,N_10691);
or U10811 (N_10811,N_10640,N_10544);
or U10812 (N_10812,N_10650,N_10785);
and U10813 (N_10813,N_10552,N_10506);
and U10814 (N_10814,N_10557,N_10736);
nand U10815 (N_10815,N_10538,N_10723);
nand U10816 (N_10816,N_10519,N_10791);
nor U10817 (N_10817,N_10796,N_10595);
and U10818 (N_10818,N_10521,N_10694);
nor U10819 (N_10819,N_10661,N_10525);
xnor U10820 (N_10820,N_10584,N_10512);
xor U10821 (N_10821,N_10622,N_10587);
and U10822 (N_10822,N_10716,N_10503);
xor U10823 (N_10823,N_10658,N_10729);
or U10824 (N_10824,N_10572,N_10630);
and U10825 (N_10825,N_10733,N_10529);
and U10826 (N_10826,N_10629,N_10666);
xor U10827 (N_10827,N_10594,N_10562);
nand U10828 (N_10828,N_10633,N_10531);
and U10829 (N_10829,N_10581,N_10662);
or U10830 (N_10830,N_10502,N_10697);
nand U10831 (N_10831,N_10509,N_10750);
nor U10832 (N_10832,N_10573,N_10575);
nand U10833 (N_10833,N_10664,N_10618);
xor U10834 (N_10834,N_10636,N_10646);
or U10835 (N_10835,N_10576,N_10756);
or U10836 (N_10836,N_10647,N_10682);
xor U10837 (N_10837,N_10550,N_10765);
and U10838 (N_10838,N_10616,N_10530);
or U10839 (N_10839,N_10588,N_10781);
or U10840 (N_10840,N_10627,N_10596);
and U10841 (N_10841,N_10523,N_10724);
xor U10842 (N_10842,N_10642,N_10679);
nor U10843 (N_10843,N_10589,N_10740);
xor U10844 (N_10844,N_10793,N_10649);
or U10845 (N_10845,N_10704,N_10707);
nor U10846 (N_10846,N_10553,N_10685);
or U10847 (N_10847,N_10563,N_10698);
or U10848 (N_10848,N_10566,N_10695);
nand U10849 (N_10849,N_10614,N_10558);
nor U10850 (N_10850,N_10675,N_10769);
xnor U10851 (N_10851,N_10717,N_10686);
and U10852 (N_10852,N_10655,N_10739);
nand U10853 (N_10853,N_10582,N_10699);
or U10854 (N_10854,N_10612,N_10790);
xor U10855 (N_10855,N_10714,N_10780);
nor U10856 (N_10856,N_10549,N_10770);
nand U10857 (N_10857,N_10577,N_10726);
xnor U10858 (N_10858,N_10602,N_10570);
and U10859 (N_10859,N_10789,N_10518);
or U10860 (N_10860,N_10702,N_10579);
or U10861 (N_10861,N_10692,N_10645);
xor U10862 (N_10862,N_10776,N_10671);
and U10863 (N_10863,N_10641,N_10626);
and U10864 (N_10864,N_10540,N_10585);
or U10865 (N_10865,N_10783,N_10779);
or U10866 (N_10866,N_10510,N_10524);
nand U10867 (N_10867,N_10732,N_10606);
nand U10868 (N_10868,N_10758,N_10745);
or U10869 (N_10869,N_10678,N_10720);
nor U10870 (N_10870,N_10635,N_10747);
nand U10871 (N_10871,N_10684,N_10787);
or U10872 (N_10872,N_10709,N_10773);
nor U10873 (N_10873,N_10623,N_10625);
nor U10874 (N_10874,N_10670,N_10619);
or U10875 (N_10875,N_10539,N_10600);
and U10876 (N_10876,N_10751,N_10718);
nor U10877 (N_10877,N_10713,N_10755);
or U10878 (N_10878,N_10797,N_10528);
xor U10879 (N_10879,N_10708,N_10559);
nor U10880 (N_10880,N_10674,N_10555);
nor U10881 (N_10881,N_10593,N_10527);
nand U10882 (N_10882,N_10688,N_10517);
nor U10883 (N_10883,N_10703,N_10772);
nand U10884 (N_10884,N_10603,N_10734);
nand U10885 (N_10885,N_10741,N_10597);
xor U10886 (N_10886,N_10590,N_10667);
xor U10887 (N_10887,N_10651,N_10774);
xor U10888 (N_10888,N_10547,N_10766);
nor U10889 (N_10889,N_10744,N_10764);
and U10890 (N_10890,N_10565,N_10537);
nand U10891 (N_10891,N_10620,N_10763);
nand U10892 (N_10892,N_10505,N_10680);
nor U10893 (N_10893,N_10788,N_10759);
nor U10894 (N_10894,N_10532,N_10543);
nand U10895 (N_10895,N_10604,N_10541);
xor U10896 (N_10896,N_10771,N_10798);
xnor U10897 (N_10897,N_10607,N_10560);
xor U10898 (N_10898,N_10513,N_10556);
nand U10899 (N_10899,N_10737,N_10504);
nor U10900 (N_10900,N_10511,N_10591);
or U10901 (N_10901,N_10592,N_10617);
and U10902 (N_10902,N_10696,N_10632);
nor U10903 (N_10903,N_10712,N_10631);
or U10904 (N_10904,N_10507,N_10615);
or U10905 (N_10905,N_10676,N_10706);
or U10906 (N_10906,N_10551,N_10526);
nor U10907 (N_10907,N_10777,N_10634);
nor U10908 (N_10908,N_10608,N_10659);
nand U10909 (N_10909,N_10710,N_10613);
nand U10910 (N_10910,N_10719,N_10554);
and U10911 (N_10911,N_10711,N_10799);
xor U10912 (N_10912,N_10792,N_10639);
nor U10913 (N_10913,N_10609,N_10730);
nand U10914 (N_10914,N_10648,N_10663);
nand U10915 (N_10915,N_10520,N_10742);
nand U10916 (N_10916,N_10561,N_10669);
and U10917 (N_10917,N_10546,N_10746);
nand U10918 (N_10918,N_10767,N_10731);
or U10919 (N_10919,N_10643,N_10687);
xnor U10920 (N_10920,N_10721,N_10605);
xnor U10921 (N_10921,N_10700,N_10534);
nor U10922 (N_10922,N_10586,N_10752);
xnor U10923 (N_10923,N_10786,N_10690);
xor U10924 (N_10924,N_10535,N_10735);
or U10925 (N_10925,N_10722,N_10610);
or U10926 (N_10926,N_10599,N_10578);
xnor U10927 (N_10927,N_10705,N_10768);
and U10928 (N_10928,N_10761,N_10673);
or U10929 (N_10929,N_10693,N_10564);
nand U10930 (N_10930,N_10598,N_10748);
nand U10931 (N_10931,N_10624,N_10545);
xnor U10932 (N_10932,N_10583,N_10727);
and U10933 (N_10933,N_10775,N_10514);
xor U10934 (N_10934,N_10757,N_10677);
nor U10935 (N_10935,N_10569,N_10715);
nor U10936 (N_10936,N_10611,N_10749);
or U10937 (N_10937,N_10683,N_10660);
nand U10938 (N_10938,N_10762,N_10754);
and U10939 (N_10939,N_10508,N_10536);
or U10940 (N_10940,N_10653,N_10753);
and U10941 (N_10941,N_10533,N_10701);
or U10942 (N_10942,N_10782,N_10668);
xnor U10943 (N_10943,N_10672,N_10628);
or U10944 (N_10944,N_10656,N_10644);
nand U10945 (N_10945,N_10542,N_10580);
xor U10946 (N_10946,N_10665,N_10567);
and U10947 (N_10947,N_10568,N_10738);
xor U10948 (N_10948,N_10501,N_10794);
xnor U10949 (N_10949,N_10778,N_10743);
and U10950 (N_10950,N_10506,N_10707);
xor U10951 (N_10951,N_10631,N_10510);
nor U10952 (N_10952,N_10741,N_10559);
xor U10953 (N_10953,N_10671,N_10684);
or U10954 (N_10954,N_10500,N_10588);
or U10955 (N_10955,N_10769,N_10556);
or U10956 (N_10956,N_10769,N_10750);
xnor U10957 (N_10957,N_10794,N_10642);
xor U10958 (N_10958,N_10718,N_10689);
and U10959 (N_10959,N_10643,N_10508);
nand U10960 (N_10960,N_10613,N_10629);
xnor U10961 (N_10961,N_10644,N_10796);
nand U10962 (N_10962,N_10764,N_10505);
xor U10963 (N_10963,N_10549,N_10656);
nand U10964 (N_10964,N_10753,N_10531);
and U10965 (N_10965,N_10773,N_10772);
nand U10966 (N_10966,N_10718,N_10665);
nor U10967 (N_10967,N_10672,N_10598);
xnor U10968 (N_10968,N_10509,N_10511);
nor U10969 (N_10969,N_10611,N_10646);
and U10970 (N_10970,N_10594,N_10500);
or U10971 (N_10971,N_10726,N_10698);
xnor U10972 (N_10972,N_10523,N_10635);
and U10973 (N_10973,N_10634,N_10627);
and U10974 (N_10974,N_10543,N_10550);
or U10975 (N_10975,N_10630,N_10709);
or U10976 (N_10976,N_10799,N_10698);
or U10977 (N_10977,N_10541,N_10545);
and U10978 (N_10978,N_10546,N_10739);
nand U10979 (N_10979,N_10500,N_10508);
or U10980 (N_10980,N_10605,N_10594);
nor U10981 (N_10981,N_10672,N_10560);
xor U10982 (N_10982,N_10502,N_10594);
and U10983 (N_10983,N_10638,N_10664);
and U10984 (N_10984,N_10593,N_10610);
and U10985 (N_10985,N_10572,N_10784);
and U10986 (N_10986,N_10637,N_10704);
xnor U10987 (N_10987,N_10658,N_10684);
and U10988 (N_10988,N_10550,N_10556);
nor U10989 (N_10989,N_10701,N_10628);
nand U10990 (N_10990,N_10624,N_10651);
nor U10991 (N_10991,N_10532,N_10591);
nor U10992 (N_10992,N_10632,N_10603);
nor U10993 (N_10993,N_10525,N_10752);
nor U10994 (N_10994,N_10718,N_10647);
or U10995 (N_10995,N_10519,N_10547);
or U10996 (N_10996,N_10670,N_10640);
nand U10997 (N_10997,N_10640,N_10556);
xor U10998 (N_10998,N_10659,N_10793);
nor U10999 (N_10999,N_10601,N_10557);
and U11000 (N_11000,N_10798,N_10747);
and U11001 (N_11001,N_10798,N_10727);
nor U11002 (N_11002,N_10547,N_10581);
or U11003 (N_11003,N_10659,N_10663);
nand U11004 (N_11004,N_10728,N_10681);
nand U11005 (N_11005,N_10512,N_10663);
or U11006 (N_11006,N_10776,N_10678);
and U11007 (N_11007,N_10636,N_10691);
nor U11008 (N_11008,N_10631,N_10500);
or U11009 (N_11009,N_10616,N_10589);
or U11010 (N_11010,N_10594,N_10624);
or U11011 (N_11011,N_10649,N_10747);
and U11012 (N_11012,N_10575,N_10695);
nand U11013 (N_11013,N_10626,N_10665);
and U11014 (N_11014,N_10725,N_10746);
and U11015 (N_11015,N_10742,N_10555);
or U11016 (N_11016,N_10732,N_10677);
nor U11017 (N_11017,N_10601,N_10564);
or U11018 (N_11018,N_10612,N_10638);
nor U11019 (N_11019,N_10638,N_10622);
nand U11020 (N_11020,N_10781,N_10742);
xnor U11021 (N_11021,N_10502,N_10793);
and U11022 (N_11022,N_10705,N_10629);
nand U11023 (N_11023,N_10533,N_10730);
xor U11024 (N_11024,N_10645,N_10727);
nand U11025 (N_11025,N_10796,N_10614);
or U11026 (N_11026,N_10777,N_10759);
and U11027 (N_11027,N_10557,N_10695);
xor U11028 (N_11028,N_10692,N_10798);
and U11029 (N_11029,N_10584,N_10529);
and U11030 (N_11030,N_10634,N_10649);
or U11031 (N_11031,N_10668,N_10566);
and U11032 (N_11032,N_10603,N_10570);
or U11033 (N_11033,N_10784,N_10757);
or U11034 (N_11034,N_10697,N_10599);
and U11035 (N_11035,N_10509,N_10667);
or U11036 (N_11036,N_10680,N_10758);
or U11037 (N_11037,N_10696,N_10639);
xnor U11038 (N_11038,N_10565,N_10704);
nand U11039 (N_11039,N_10534,N_10724);
nand U11040 (N_11040,N_10666,N_10619);
or U11041 (N_11041,N_10669,N_10597);
xnor U11042 (N_11042,N_10746,N_10712);
or U11043 (N_11043,N_10503,N_10780);
nand U11044 (N_11044,N_10790,N_10753);
nand U11045 (N_11045,N_10562,N_10593);
nor U11046 (N_11046,N_10507,N_10737);
nand U11047 (N_11047,N_10745,N_10650);
or U11048 (N_11048,N_10655,N_10537);
or U11049 (N_11049,N_10711,N_10559);
or U11050 (N_11050,N_10561,N_10557);
nand U11051 (N_11051,N_10570,N_10521);
and U11052 (N_11052,N_10782,N_10792);
nand U11053 (N_11053,N_10579,N_10522);
or U11054 (N_11054,N_10764,N_10568);
or U11055 (N_11055,N_10607,N_10509);
nand U11056 (N_11056,N_10635,N_10520);
nand U11057 (N_11057,N_10508,N_10781);
and U11058 (N_11058,N_10744,N_10652);
and U11059 (N_11059,N_10669,N_10708);
nand U11060 (N_11060,N_10766,N_10609);
xnor U11061 (N_11061,N_10647,N_10550);
or U11062 (N_11062,N_10551,N_10634);
nand U11063 (N_11063,N_10506,N_10593);
or U11064 (N_11064,N_10584,N_10516);
xor U11065 (N_11065,N_10526,N_10740);
or U11066 (N_11066,N_10627,N_10590);
or U11067 (N_11067,N_10654,N_10694);
xor U11068 (N_11068,N_10749,N_10554);
and U11069 (N_11069,N_10710,N_10605);
xnor U11070 (N_11070,N_10591,N_10670);
nand U11071 (N_11071,N_10597,N_10680);
nor U11072 (N_11072,N_10633,N_10783);
nand U11073 (N_11073,N_10640,N_10720);
and U11074 (N_11074,N_10743,N_10628);
nor U11075 (N_11075,N_10526,N_10506);
xnor U11076 (N_11076,N_10531,N_10738);
or U11077 (N_11077,N_10651,N_10702);
nor U11078 (N_11078,N_10509,N_10644);
or U11079 (N_11079,N_10775,N_10598);
xnor U11080 (N_11080,N_10613,N_10764);
and U11081 (N_11081,N_10559,N_10775);
and U11082 (N_11082,N_10782,N_10582);
or U11083 (N_11083,N_10669,N_10530);
nor U11084 (N_11084,N_10785,N_10762);
nand U11085 (N_11085,N_10750,N_10672);
xor U11086 (N_11086,N_10620,N_10577);
and U11087 (N_11087,N_10667,N_10704);
xor U11088 (N_11088,N_10774,N_10713);
nor U11089 (N_11089,N_10645,N_10584);
nor U11090 (N_11090,N_10556,N_10647);
or U11091 (N_11091,N_10558,N_10635);
nand U11092 (N_11092,N_10503,N_10746);
or U11093 (N_11093,N_10527,N_10628);
xnor U11094 (N_11094,N_10529,N_10588);
nand U11095 (N_11095,N_10771,N_10680);
or U11096 (N_11096,N_10656,N_10602);
nand U11097 (N_11097,N_10513,N_10658);
or U11098 (N_11098,N_10769,N_10799);
or U11099 (N_11099,N_10657,N_10773);
xnor U11100 (N_11100,N_10985,N_10847);
nand U11101 (N_11101,N_10987,N_11034);
or U11102 (N_11102,N_11003,N_11038);
nor U11103 (N_11103,N_11099,N_10826);
or U11104 (N_11104,N_10886,N_10866);
or U11105 (N_11105,N_10849,N_11065);
xor U11106 (N_11106,N_10812,N_11002);
and U11107 (N_11107,N_10843,N_10909);
nor U11108 (N_11108,N_10890,N_11049);
or U11109 (N_11109,N_10803,N_10901);
nand U11110 (N_11110,N_10859,N_11011);
and U11111 (N_11111,N_11053,N_11080);
or U11112 (N_11112,N_10887,N_10807);
nor U11113 (N_11113,N_10913,N_11076);
or U11114 (N_11114,N_11057,N_10802);
or U11115 (N_11115,N_11030,N_10836);
nand U11116 (N_11116,N_10980,N_10894);
xnor U11117 (N_11117,N_10883,N_10858);
nor U11118 (N_11118,N_10846,N_10820);
nor U11119 (N_11119,N_10902,N_10823);
or U11120 (N_11120,N_10956,N_11075);
nor U11121 (N_11121,N_11022,N_10825);
xnor U11122 (N_11122,N_11010,N_10941);
nand U11123 (N_11123,N_10939,N_10917);
nand U11124 (N_11124,N_10915,N_11087);
and U11125 (N_11125,N_10831,N_10994);
and U11126 (N_11126,N_11071,N_11031);
and U11127 (N_11127,N_11061,N_10923);
nor U11128 (N_11128,N_11067,N_11036);
nor U11129 (N_11129,N_10912,N_11016);
nand U11130 (N_11130,N_10801,N_10844);
nand U11131 (N_11131,N_10863,N_11058);
or U11132 (N_11132,N_10851,N_10918);
or U11133 (N_11133,N_11007,N_11042);
and U11134 (N_11134,N_10869,N_11056);
xnor U11135 (N_11135,N_11025,N_10855);
nor U11136 (N_11136,N_10822,N_10862);
nor U11137 (N_11137,N_11023,N_10930);
or U11138 (N_11138,N_11004,N_10906);
nor U11139 (N_11139,N_10943,N_10947);
nand U11140 (N_11140,N_11045,N_10977);
xor U11141 (N_11141,N_10963,N_11079);
or U11142 (N_11142,N_11054,N_10845);
or U11143 (N_11143,N_10903,N_10905);
or U11144 (N_11144,N_10817,N_10870);
and U11145 (N_11145,N_10891,N_10975);
xnor U11146 (N_11146,N_10920,N_10962);
nor U11147 (N_11147,N_10981,N_11090);
nor U11148 (N_11148,N_10974,N_10976);
xor U11149 (N_11149,N_10884,N_11094);
nor U11150 (N_11150,N_10996,N_11040);
nand U11151 (N_11151,N_10937,N_10986);
nor U11152 (N_11152,N_10919,N_10875);
and U11153 (N_11153,N_11033,N_11089);
xor U11154 (N_11154,N_10856,N_10871);
nand U11155 (N_11155,N_10972,N_11077);
xor U11156 (N_11156,N_11006,N_11028);
nand U11157 (N_11157,N_10935,N_10973);
nor U11158 (N_11158,N_11062,N_10879);
nor U11159 (N_11159,N_10910,N_10874);
or U11160 (N_11160,N_10885,N_10997);
or U11161 (N_11161,N_10818,N_11069);
or U11162 (N_11162,N_11017,N_10848);
xnor U11163 (N_11163,N_10804,N_11008);
and U11164 (N_11164,N_10998,N_10928);
nor U11165 (N_11165,N_10931,N_11029);
nand U11166 (N_11166,N_10893,N_10927);
xnor U11167 (N_11167,N_11021,N_10840);
nor U11168 (N_11168,N_11097,N_11005);
xnor U11169 (N_11169,N_10969,N_11085);
or U11170 (N_11170,N_11060,N_10999);
or U11171 (N_11171,N_11088,N_10979);
nand U11172 (N_11172,N_10934,N_11055);
or U11173 (N_11173,N_10809,N_11070);
nand U11174 (N_11174,N_10867,N_10814);
and U11175 (N_11175,N_11092,N_10800);
xor U11176 (N_11176,N_10970,N_11020);
or U11177 (N_11177,N_11019,N_11095);
nor U11178 (N_11178,N_10982,N_10929);
or U11179 (N_11179,N_11084,N_10932);
xnor U11180 (N_11180,N_10868,N_10907);
xnor U11181 (N_11181,N_10916,N_11096);
or U11182 (N_11182,N_10889,N_10936);
or U11183 (N_11183,N_10957,N_11052);
and U11184 (N_11184,N_11059,N_10881);
nand U11185 (N_11185,N_10834,N_11027);
xnor U11186 (N_11186,N_11043,N_10921);
xnor U11187 (N_11187,N_10908,N_10924);
nor U11188 (N_11188,N_11024,N_10984);
nor U11189 (N_11189,N_10964,N_10938);
nor U11190 (N_11190,N_10983,N_11082);
or U11191 (N_11191,N_10830,N_10819);
and U11192 (N_11192,N_10816,N_11039);
and U11193 (N_11193,N_10968,N_10864);
or U11194 (N_11194,N_10925,N_10990);
or U11195 (N_11195,N_10949,N_11001);
xnor U11196 (N_11196,N_10805,N_10954);
or U11197 (N_11197,N_11068,N_11050);
or U11198 (N_11198,N_11009,N_10948);
nand U11199 (N_11199,N_10951,N_10810);
or U11200 (N_11200,N_11051,N_10961);
nand U11201 (N_11201,N_11078,N_10960);
and U11202 (N_11202,N_11093,N_10876);
nand U11203 (N_11203,N_10991,N_11012);
or U11204 (N_11204,N_10878,N_10940);
or U11205 (N_11205,N_10882,N_10971);
and U11206 (N_11206,N_10877,N_10873);
or U11207 (N_11207,N_11037,N_10911);
or U11208 (N_11208,N_10989,N_10950);
nor U11209 (N_11209,N_10904,N_11035);
and U11210 (N_11210,N_11081,N_11083);
xor U11211 (N_11211,N_10857,N_10835);
nand U11212 (N_11212,N_10899,N_10828);
xor U11213 (N_11213,N_10933,N_11018);
or U11214 (N_11214,N_11041,N_10914);
xor U11215 (N_11215,N_10959,N_10992);
nand U11216 (N_11216,N_11074,N_10955);
xor U11217 (N_11217,N_10806,N_10922);
or U11218 (N_11218,N_10898,N_11044);
or U11219 (N_11219,N_10993,N_11091);
xnor U11220 (N_11220,N_10850,N_10861);
and U11221 (N_11221,N_10860,N_10946);
or U11222 (N_11222,N_10839,N_10958);
and U11223 (N_11223,N_10892,N_10945);
nand U11224 (N_11224,N_10833,N_10815);
nand U11225 (N_11225,N_10897,N_11073);
xnor U11226 (N_11226,N_10813,N_11048);
or U11227 (N_11227,N_11015,N_11014);
xnor U11228 (N_11228,N_10824,N_10832);
or U11229 (N_11229,N_10838,N_10988);
nor U11230 (N_11230,N_10821,N_11066);
and U11231 (N_11231,N_10966,N_11072);
and U11232 (N_11232,N_11063,N_10827);
and U11233 (N_11233,N_10829,N_10811);
nand U11234 (N_11234,N_11032,N_10888);
and U11235 (N_11235,N_10926,N_10965);
or U11236 (N_11236,N_11013,N_11098);
nor U11237 (N_11237,N_10896,N_11026);
and U11238 (N_11238,N_10944,N_10900);
and U11239 (N_11239,N_10853,N_10880);
or U11240 (N_11240,N_10952,N_10865);
nor U11241 (N_11241,N_10967,N_10872);
or U11242 (N_11242,N_10852,N_11047);
xnor U11243 (N_11243,N_10854,N_11086);
nor U11244 (N_11244,N_10895,N_11046);
xor U11245 (N_11245,N_10837,N_10808);
and U11246 (N_11246,N_10842,N_10841);
or U11247 (N_11247,N_11000,N_10942);
or U11248 (N_11248,N_10995,N_11064);
nor U11249 (N_11249,N_10978,N_10953);
nand U11250 (N_11250,N_10941,N_11037);
or U11251 (N_11251,N_11098,N_10850);
nor U11252 (N_11252,N_11021,N_10982);
or U11253 (N_11253,N_10848,N_10874);
or U11254 (N_11254,N_11094,N_11042);
nand U11255 (N_11255,N_10925,N_10803);
nor U11256 (N_11256,N_10863,N_11052);
and U11257 (N_11257,N_11070,N_10861);
and U11258 (N_11258,N_10898,N_10825);
and U11259 (N_11259,N_10947,N_11077);
xor U11260 (N_11260,N_11079,N_11069);
xnor U11261 (N_11261,N_11081,N_10888);
or U11262 (N_11262,N_10862,N_10848);
and U11263 (N_11263,N_10834,N_10865);
or U11264 (N_11264,N_11049,N_10826);
xnor U11265 (N_11265,N_10827,N_11099);
or U11266 (N_11266,N_10855,N_11067);
nand U11267 (N_11267,N_10893,N_10841);
nand U11268 (N_11268,N_10936,N_10844);
or U11269 (N_11269,N_10894,N_11072);
nor U11270 (N_11270,N_11031,N_10895);
or U11271 (N_11271,N_10810,N_10870);
or U11272 (N_11272,N_10811,N_11006);
xnor U11273 (N_11273,N_10996,N_10960);
or U11274 (N_11274,N_10806,N_10937);
nand U11275 (N_11275,N_10861,N_10939);
nor U11276 (N_11276,N_10906,N_10875);
nor U11277 (N_11277,N_10842,N_10916);
nor U11278 (N_11278,N_11095,N_11022);
nand U11279 (N_11279,N_11028,N_10971);
and U11280 (N_11280,N_10899,N_10963);
xnor U11281 (N_11281,N_10886,N_10818);
nand U11282 (N_11282,N_11026,N_11056);
nand U11283 (N_11283,N_10812,N_10946);
or U11284 (N_11284,N_11036,N_10950);
or U11285 (N_11285,N_10985,N_10876);
and U11286 (N_11286,N_11047,N_10813);
or U11287 (N_11287,N_10846,N_10875);
nand U11288 (N_11288,N_11012,N_11089);
and U11289 (N_11289,N_11068,N_10911);
nand U11290 (N_11290,N_11017,N_10891);
or U11291 (N_11291,N_10867,N_11011);
or U11292 (N_11292,N_11020,N_11021);
and U11293 (N_11293,N_10985,N_10961);
nor U11294 (N_11294,N_10991,N_10839);
or U11295 (N_11295,N_10823,N_11072);
nor U11296 (N_11296,N_10961,N_10801);
nor U11297 (N_11297,N_11045,N_10820);
and U11298 (N_11298,N_11061,N_10890);
nand U11299 (N_11299,N_10904,N_11044);
nand U11300 (N_11300,N_10897,N_11006);
and U11301 (N_11301,N_10898,N_10945);
and U11302 (N_11302,N_11049,N_10855);
nor U11303 (N_11303,N_10874,N_11046);
xor U11304 (N_11304,N_10969,N_11032);
xor U11305 (N_11305,N_11056,N_10950);
nor U11306 (N_11306,N_10847,N_10909);
nand U11307 (N_11307,N_10820,N_10919);
and U11308 (N_11308,N_10945,N_10988);
xor U11309 (N_11309,N_10823,N_10892);
xnor U11310 (N_11310,N_10942,N_11036);
xor U11311 (N_11311,N_11075,N_10978);
nand U11312 (N_11312,N_10814,N_11035);
and U11313 (N_11313,N_10887,N_11072);
nand U11314 (N_11314,N_10808,N_10924);
and U11315 (N_11315,N_10845,N_10934);
nor U11316 (N_11316,N_11063,N_10877);
xnor U11317 (N_11317,N_11040,N_10902);
or U11318 (N_11318,N_10973,N_10892);
nand U11319 (N_11319,N_10840,N_10880);
and U11320 (N_11320,N_10971,N_11059);
xnor U11321 (N_11321,N_10992,N_11088);
nor U11322 (N_11322,N_10809,N_10936);
xnor U11323 (N_11323,N_11089,N_10878);
or U11324 (N_11324,N_10975,N_10977);
or U11325 (N_11325,N_11060,N_10942);
nand U11326 (N_11326,N_10894,N_11077);
nand U11327 (N_11327,N_10807,N_10814);
and U11328 (N_11328,N_10806,N_11020);
and U11329 (N_11329,N_10837,N_11005);
nand U11330 (N_11330,N_10924,N_11000);
nand U11331 (N_11331,N_10982,N_11062);
xor U11332 (N_11332,N_10977,N_10869);
xnor U11333 (N_11333,N_11093,N_10894);
nand U11334 (N_11334,N_10898,N_10811);
xor U11335 (N_11335,N_10922,N_11074);
or U11336 (N_11336,N_11002,N_10826);
or U11337 (N_11337,N_10923,N_10970);
or U11338 (N_11338,N_11028,N_10999);
or U11339 (N_11339,N_11002,N_11021);
or U11340 (N_11340,N_11060,N_10890);
or U11341 (N_11341,N_10826,N_10956);
and U11342 (N_11342,N_10819,N_11036);
nor U11343 (N_11343,N_10910,N_10922);
nor U11344 (N_11344,N_11088,N_10937);
or U11345 (N_11345,N_11013,N_10959);
nand U11346 (N_11346,N_10987,N_11013);
and U11347 (N_11347,N_10862,N_10829);
and U11348 (N_11348,N_10957,N_10963);
nand U11349 (N_11349,N_10890,N_10914);
nor U11350 (N_11350,N_11029,N_11060);
or U11351 (N_11351,N_10942,N_10862);
nor U11352 (N_11352,N_10948,N_10807);
nand U11353 (N_11353,N_10855,N_10970);
nand U11354 (N_11354,N_10817,N_10931);
nand U11355 (N_11355,N_11087,N_10992);
and U11356 (N_11356,N_11058,N_10958);
nand U11357 (N_11357,N_10833,N_10886);
nor U11358 (N_11358,N_10893,N_10934);
nor U11359 (N_11359,N_11043,N_11092);
xor U11360 (N_11360,N_11038,N_10916);
xnor U11361 (N_11361,N_10969,N_10883);
nand U11362 (N_11362,N_11053,N_10871);
nor U11363 (N_11363,N_10805,N_10913);
or U11364 (N_11364,N_10978,N_10930);
xnor U11365 (N_11365,N_10921,N_10956);
and U11366 (N_11366,N_10974,N_11082);
or U11367 (N_11367,N_10877,N_10860);
or U11368 (N_11368,N_10912,N_11027);
and U11369 (N_11369,N_10861,N_10983);
nor U11370 (N_11370,N_11085,N_10998);
and U11371 (N_11371,N_10840,N_11084);
nand U11372 (N_11372,N_11045,N_11040);
and U11373 (N_11373,N_11050,N_10932);
nand U11374 (N_11374,N_11021,N_10981);
xnor U11375 (N_11375,N_10871,N_11051);
nor U11376 (N_11376,N_11080,N_11067);
nand U11377 (N_11377,N_11025,N_10989);
and U11378 (N_11378,N_10942,N_10822);
and U11379 (N_11379,N_11085,N_10845);
nor U11380 (N_11380,N_10946,N_10884);
and U11381 (N_11381,N_11010,N_10972);
or U11382 (N_11382,N_10863,N_11054);
and U11383 (N_11383,N_10871,N_10890);
or U11384 (N_11384,N_11013,N_10858);
or U11385 (N_11385,N_10885,N_10890);
or U11386 (N_11386,N_11042,N_10818);
or U11387 (N_11387,N_10916,N_11020);
nand U11388 (N_11388,N_10990,N_10981);
and U11389 (N_11389,N_10857,N_10849);
nor U11390 (N_11390,N_11054,N_10960);
nand U11391 (N_11391,N_10824,N_10939);
or U11392 (N_11392,N_11043,N_10962);
nor U11393 (N_11393,N_10886,N_10897);
nand U11394 (N_11394,N_10800,N_10816);
xor U11395 (N_11395,N_10838,N_11059);
xor U11396 (N_11396,N_11065,N_11024);
nand U11397 (N_11397,N_11083,N_10859);
nor U11398 (N_11398,N_10963,N_10873);
nand U11399 (N_11399,N_10917,N_10862);
nand U11400 (N_11400,N_11385,N_11212);
or U11401 (N_11401,N_11139,N_11276);
nor U11402 (N_11402,N_11309,N_11300);
and U11403 (N_11403,N_11354,N_11389);
xor U11404 (N_11404,N_11103,N_11229);
and U11405 (N_11405,N_11270,N_11214);
nand U11406 (N_11406,N_11337,N_11114);
or U11407 (N_11407,N_11192,N_11327);
and U11408 (N_11408,N_11116,N_11169);
nor U11409 (N_11409,N_11363,N_11340);
nor U11410 (N_11410,N_11272,N_11143);
or U11411 (N_11411,N_11162,N_11197);
nand U11412 (N_11412,N_11240,N_11245);
nor U11413 (N_11413,N_11396,N_11350);
xor U11414 (N_11414,N_11282,N_11283);
or U11415 (N_11415,N_11264,N_11379);
nand U11416 (N_11416,N_11230,N_11320);
or U11417 (N_11417,N_11256,N_11382);
nor U11418 (N_11418,N_11135,N_11304);
and U11419 (N_11419,N_11299,N_11279);
nand U11420 (N_11420,N_11165,N_11301);
xor U11421 (N_11421,N_11374,N_11119);
or U11422 (N_11422,N_11338,N_11369);
nor U11423 (N_11423,N_11265,N_11222);
and U11424 (N_11424,N_11336,N_11190);
and U11425 (N_11425,N_11231,N_11296);
nand U11426 (N_11426,N_11130,N_11360);
or U11427 (N_11427,N_11101,N_11129);
nor U11428 (N_11428,N_11237,N_11258);
nor U11429 (N_11429,N_11148,N_11259);
nand U11430 (N_11430,N_11315,N_11203);
xnor U11431 (N_11431,N_11145,N_11206);
and U11432 (N_11432,N_11275,N_11274);
nor U11433 (N_11433,N_11388,N_11316);
nand U11434 (N_11434,N_11381,N_11368);
nand U11435 (N_11435,N_11251,N_11149);
and U11436 (N_11436,N_11371,N_11106);
xor U11437 (N_11437,N_11321,N_11186);
or U11438 (N_11438,N_11118,N_11141);
nor U11439 (N_11439,N_11226,N_11220);
xnor U11440 (N_11440,N_11397,N_11344);
nor U11441 (N_11441,N_11355,N_11158);
and U11442 (N_11442,N_11399,N_11173);
nand U11443 (N_11443,N_11361,N_11117);
xnor U11444 (N_11444,N_11163,N_11370);
nand U11445 (N_11445,N_11104,N_11310);
or U11446 (N_11446,N_11291,N_11280);
nor U11447 (N_11447,N_11202,N_11288);
or U11448 (N_11448,N_11260,N_11257);
or U11449 (N_11449,N_11312,N_11255);
xnor U11450 (N_11450,N_11234,N_11210);
nor U11451 (N_11451,N_11228,N_11306);
or U11452 (N_11452,N_11215,N_11343);
nand U11453 (N_11453,N_11244,N_11286);
and U11454 (N_11454,N_11236,N_11156);
xor U11455 (N_11455,N_11387,N_11233);
xor U11456 (N_11456,N_11136,N_11191);
and U11457 (N_11457,N_11249,N_11178);
nor U11458 (N_11458,N_11390,N_11225);
or U11459 (N_11459,N_11107,N_11252);
xnor U11460 (N_11460,N_11323,N_11184);
or U11461 (N_11461,N_11305,N_11398);
or U11462 (N_11462,N_11317,N_11324);
or U11463 (N_11463,N_11281,N_11357);
and U11464 (N_11464,N_11395,N_11166);
nor U11465 (N_11465,N_11375,N_11298);
and U11466 (N_11466,N_11378,N_11183);
xnor U11467 (N_11467,N_11289,N_11219);
nor U11468 (N_11468,N_11356,N_11137);
and U11469 (N_11469,N_11261,N_11271);
and U11470 (N_11470,N_11247,N_11221);
nand U11471 (N_11471,N_11151,N_11372);
nor U11472 (N_11472,N_11349,N_11268);
nor U11473 (N_11473,N_11285,N_11150);
nand U11474 (N_11474,N_11170,N_11175);
and U11475 (N_11475,N_11174,N_11154);
nor U11476 (N_11476,N_11110,N_11250);
and U11477 (N_11477,N_11189,N_11105);
or U11478 (N_11478,N_11140,N_11125);
xnor U11479 (N_11479,N_11328,N_11193);
nor U11480 (N_11480,N_11159,N_11134);
and U11481 (N_11481,N_11180,N_11242);
and U11482 (N_11482,N_11112,N_11196);
or U11483 (N_11483,N_11109,N_11188);
or U11484 (N_11484,N_11176,N_11339);
nor U11485 (N_11485,N_11126,N_11380);
xor U11486 (N_11486,N_11120,N_11391);
or U11487 (N_11487,N_11314,N_11152);
nand U11488 (N_11488,N_11364,N_11253);
nor U11489 (N_11489,N_11122,N_11108);
and U11490 (N_11490,N_11346,N_11347);
xor U11491 (N_11491,N_11232,N_11142);
and U11492 (N_11492,N_11102,N_11377);
xnor U11493 (N_11493,N_11345,N_11341);
or U11494 (N_11494,N_11333,N_11123);
nor U11495 (N_11495,N_11208,N_11155);
nand U11496 (N_11496,N_11171,N_11386);
and U11497 (N_11497,N_11157,N_11278);
xnor U11498 (N_11498,N_11313,N_11351);
nand U11499 (N_11499,N_11373,N_11352);
xnor U11500 (N_11500,N_11376,N_11273);
nor U11501 (N_11501,N_11307,N_11209);
xnor U11502 (N_11502,N_11133,N_11172);
nand U11503 (N_11503,N_11128,N_11263);
or U11504 (N_11504,N_11358,N_11287);
nand U11505 (N_11505,N_11290,N_11329);
or U11506 (N_11506,N_11204,N_11182);
xor U11507 (N_11507,N_11223,N_11217);
and U11508 (N_11508,N_11200,N_11367);
nand U11509 (N_11509,N_11332,N_11238);
or U11510 (N_11510,N_11383,N_11277);
xor U11511 (N_11511,N_11113,N_11392);
nand U11512 (N_11512,N_11294,N_11394);
and U11513 (N_11513,N_11235,N_11322);
nor U11514 (N_11514,N_11311,N_11303);
or U11515 (N_11515,N_11144,N_11164);
and U11516 (N_11516,N_11132,N_11269);
nor U11517 (N_11517,N_11262,N_11246);
and U11518 (N_11518,N_11218,N_11198);
nand U11519 (N_11519,N_11199,N_11267);
or U11520 (N_11520,N_11297,N_11124);
nand U11521 (N_11521,N_11131,N_11319);
xor U11522 (N_11522,N_11266,N_11342);
and U11523 (N_11523,N_11161,N_11318);
nand U11524 (N_11524,N_11201,N_11177);
nand U11525 (N_11525,N_11362,N_11195);
nand U11526 (N_11526,N_11153,N_11211);
nand U11527 (N_11527,N_11147,N_11254);
or U11528 (N_11528,N_11207,N_11205);
nand U11529 (N_11529,N_11366,N_11216);
xnor U11530 (N_11530,N_11335,N_11168);
nor U11531 (N_11531,N_11146,N_11292);
xor U11532 (N_11532,N_11302,N_11127);
nand U11533 (N_11533,N_11115,N_11179);
xnor U11534 (N_11534,N_11393,N_11160);
and U11535 (N_11535,N_11308,N_11359);
xnor U11536 (N_11536,N_11194,N_11111);
nand U11537 (N_11537,N_11187,N_11243);
and U11538 (N_11538,N_11121,N_11365);
nand U11539 (N_11539,N_11213,N_11284);
and U11540 (N_11540,N_11353,N_11334);
nor U11541 (N_11541,N_11384,N_11331);
or U11542 (N_11542,N_11293,N_11326);
and U11543 (N_11543,N_11185,N_11241);
xor U11544 (N_11544,N_11248,N_11227);
or U11545 (N_11545,N_11100,N_11295);
and U11546 (N_11546,N_11239,N_11167);
nor U11547 (N_11547,N_11138,N_11348);
xnor U11548 (N_11548,N_11224,N_11325);
nand U11549 (N_11549,N_11330,N_11181);
nand U11550 (N_11550,N_11180,N_11183);
and U11551 (N_11551,N_11125,N_11186);
or U11552 (N_11552,N_11394,N_11146);
xnor U11553 (N_11553,N_11168,N_11123);
xor U11554 (N_11554,N_11136,N_11354);
nor U11555 (N_11555,N_11243,N_11108);
nand U11556 (N_11556,N_11202,N_11344);
and U11557 (N_11557,N_11343,N_11197);
or U11558 (N_11558,N_11152,N_11170);
and U11559 (N_11559,N_11140,N_11137);
nand U11560 (N_11560,N_11296,N_11362);
xnor U11561 (N_11561,N_11342,N_11118);
or U11562 (N_11562,N_11123,N_11170);
or U11563 (N_11563,N_11100,N_11258);
nor U11564 (N_11564,N_11382,N_11301);
or U11565 (N_11565,N_11366,N_11205);
nor U11566 (N_11566,N_11373,N_11364);
xor U11567 (N_11567,N_11133,N_11173);
nand U11568 (N_11568,N_11359,N_11149);
nand U11569 (N_11569,N_11346,N_11179);
xor U11570 (N_11570,N_11321,N_11144);
xor U11571 (N_11571,N_11206,N_11106);
nor U11572 (N_11572,N_11380,N_11185);
and U11573 (N_11573,N_11238,N_11218);
nor U11574 (N_11574,N_11356,N_11174);
or U11575 (N_11575,N_11194,N_11388);
nand U11576 (N_11576,N_11152,N_11272);
xor U11577 (N_11577,N_11144,N_11200);
xor U11578 (N_11578,N_11142,N_11136);
nor U11579 (N_11579,N_11296,N_11375);
xor U11580 (N_11580,N_11314,N_11229);
nand U11581 (N_11581,N_11200,N_11227);
xor U11582 (N_11582,N_11277,N_11392);
nor U11583 (N_11583,N_11371,N_11346);
nor U11584 (N_11584,N_11290,N_11213);
nand U11585 (N_11585,N_11111,N_11198);
xor U11586 (N_11586,N_11323,N_11110);
nor U11587 (N_11587,N_11142,N_11351);
nand U11588 (N_11588,N_11390,N_11311);
nor U11589 (N_11589,N_11389,N_11314);
and U11590 (N_11590,N_11294,N_11365);
or U11591 (N_11591,N_11295,N_11385);
xor U11592 (N_11592,N_11379,N_11313);
or U11593 (N_11593,N_11391,N_11108);
xnor U11594 (N_11594,N_11195,N_11222);
nand U11595 (N_11595,N_11386,N_11261);
nor U11596 (N_11596,N_11215,N_11377);
nand U11597 (N_11597,N_11355,N_11352);
xor U11598 (N_11598,N_11268,N_11267);
and U11599 (N_11599,N_11184,N_11299);
xnor U11600 (N_11600,N_11196,N_11116);
nor U11601 (N_11601,N_11210,N_11339);
xnor U11602 (N_11602,N_11267,N_11238);
nand U11603 (N_11603,N_11102,N_11135);
xnor U11604 (N_11604,N_11365,N_11259);
and U11605 (N_11605,N_11239,N_11276);
nand U11606 (N_11606,N_11128,N_11377);
nor U11607 (N_11607,N_11294,N_11198);
and U11608 (N_11608,N_11284,N_11320);
xnor U11609 (N_11609,N_11392,N_11285);
xnor U11610 (N_11610,N_11271,N_11228);
and U11611 (N_11611,N_11348,N_11174);
or U11612 (N_11612,N_11322,N_11177);
nor U11613 (N_11613,N_11167,N_11316);
xor U11614 (N_11614,N_11240,N_11349);
xnor U11615 (N_11615,N_11166,N_11168);
nor U11616 (N_11616,N_11343,N_11334);
or U11617 (N_11617,N_11383,N_11322);
and U11618 (N_11618,N_11316,N_11190);
nand U11619 (N_11619,N_11232,N_11313);
nand U11620 (N_11620,N_11216,N_11190);
or U11621 (N_11621,N_11221,N_11143);
nand U11622 (N_11622,N_11379,N_11211);
and U11623 (N_11623,N_11342,N_11330);
or U11624 (N_11624,N_11140,N_11299);
xnor U11625 (N_11625,N_11132,N_11243);
nor U11626 (N_11626,N_11323,N_11318);
or U11627 (N_11627,N_11337,N_11396);
nand U11628 (N_11628,N_11119,N_11160);
xor U11629 (N_11629,N_11361,N_11152);
nand U11630 (N_11630,N_11187,N_11256);
nor U11631 (N_11631,N_11185,N_11323);
and U11632 (N_11632,N_11260,N_11153);
and U11633 (N_11633,N_11164,N_11382);
xnor U11634 (N_11634,N_11116,N_11334);
and U11635 (N_11635,N_11396,N_11392);
nor U11636 (N_11636,N_11255,N_11358);
and U11637 (N_11637,N_11326,N_11288);
nor U11638 (N_11638,N_11130,N_11270);
xnor U11639 (N_11639,N_11315,N_11340);
and U11640 (N_11640,N_11343,N_11393);
and U11641 (N_11641,N_11219,N_11377);
nand U11642 (N_11642,N_11176,N_11315);
xor U11643 (N_11643,N_11183,N_11104);
or U11644 (N_11644,N_11308,N_11101);
nand U11645 (N_11645,N_11201,N_11391);
or U11646 (N_11646,N_11266,N_11124);
or U11647 (N_11647,N_11245,N_11235);
nor U11648 (N_11648,N_11360,N_11148);
nor U11649 (N_11649,N_11108,N_11156);
xnor U11650 (N_11650,N_11356,N_11321);
xnor U11651 (N_11651,N_11211,N_11185);
nand U11652 (N_11652,N_11390,N_11236);
nor U11653 (N_11653,N_11211,N_11149);
and U11654 (N_11654,N_11156,N_11357);
nand U11655 (N_11655,N_11312,N_11147);
or U11656 (N_11656,N_11216,N_11253);
and U11657 (N_11657,N_11209,N_11103);
and U11658 (N_11658,N_11263,N_11275);
and U11659 (N_11659,N_11385,N_11324);
or U11660 (N_11660,N_11315,N_11361);
xnor U11661 (N_11661,N_11164,N_11188);
xnor U11662 (N_11662,N_11263,N_11152);
or U11663 (N_11663,N_11324,N_11356);
or U11664 (N_11664,N_11356,N_11348);
nand U11665 (N_11665,N_11327,N_11107);
and U11666 (N_11666,N_11256,N_11208);
nand U11667 (N_11667,N_11158,N_11169);
xor U11668 (N_11668,N_11170,N_11336);
and U11669 (N_11669,N_11322,N_11214);
nor U11670 (N_11670,N_11246,N_11243);
xnor U11671 (N_11671,N_11327,N_11309);
xor U11672 (N_11672,N_11215,N_11385);
nand U11673 (N_11673,N_11327,N_11281);
nor U11674 (N_11674,N_11177,N_11293);
xor U11675 (N_11675,N_11228,N_11291);
xor U11676 (N_11676,N_11179,N_11144);
and U11677 (N_11677,N_11301,N_11143);
and U11678 (N_11678,N_11201,N_11381);
nand U11679 (N_11679,N_11179,N_11257);
or U11680 (N_11680,N_11282,N_11114);
nor U11681 (N_11681,N_11106,N_11164);
nor U11682 (N_11682,N_11374,N_11332);
and U11683 (N_11683,N_11381,N_11206);
nor U11684 (N_11684,N_11108,N_11297);
xor U11685 (N_11685,N_11145,N_11241);
xor U11686 (N_11686,N_11208,N_11119);
nor U11687 (N_11687,N_11129,N_11182);
xor U11688 (N_11688,N_11174,N_11229);
nand U11689 (N_11689,N_11119,N_11200);
and U11690 (N_11690,N_11290,N_11159);
nor U11691 (N_11691,N_11241,N_11343);
xnor U11692 (N_11692,N_11189,N_11305);
and U11693 (N_11693,N_11320,N_11181);
xor U11694 (N_11694,N_11369,N_11176);
nand U11695 (N_11695,N_11393,N_11185);
xnor U11696 (N_11696,N_11220,N_11150);
or U11697 (N_11697,N_11341,N_11127);
nand U11698 (N_11698,N_11317,N_11174);
or U11699 (N_11699,N_11350,N_11374);
xor U11700 (N_11700,N_11401,N_11682);
nand U11701 (N_11701,N_11509,N_11523);
nand U11702 (N_11702,N_11551,N_11593);
and U11703 (N_11703,N_11455,N_11627);
or U11704 (N_11704,N_11442,N_11424);
xnor U11705 (N_11705,N_11651,N_11521);
nand U11706 (N_11706,N_11652,N_11426);
or U11707 (N_11707,N_11404,N_11497);
nand U11708 (N_11708,N_11562,N_11587);
xor U11709 (N_11709,N_11400,N_11576);
nor U11710 (N_11710,N_11644,N_11403);
nor U11711 (N_11711,N_11467,N_11500);
nand U11712 (N_11712,N_11417,N_11406);
and U11713 (N_11713,N_11501,N_11461);
xor U11714 (N_11714,N_11561,N_11583);
and U11715 (N_11715,N_11436,N_11591);
xor U11716 (N_11716,N_11451,N_11645);
and U11717 (N_11717,N_11588,N_11445);
xnor U11718 (N_11718,N_11435,N_11526);
or U11719 (N_11719,N_11678,N_11615);
nand U11720 (N_11720,N_11520,N_11639);
or U11721 (N_11721,N_11533,N_11494);
or U11722 (N_11722,N_11680,N_11676);
or U11723 (N_11723,N_11699,N_11558);
and U11724 (N_11724,N_11548,N_11440);
or U11725 (N_11725,N_11664,N_11646);
xnor U11726 (N_11726,N_11454,N_11609);
nor U11727 (N_11727,N_11517,N_11616);
xnor U11728 (N_11728,N_11546,N_11656);
xor U11729 (N_11729,N_11429,N_11675);
nand U11730 (N_11730,N_11490,N_11574);
nor U11731 (N_11731,N_11507,N_11430);
nand U11732 (N_11732,N_11554,N_11688);
and U11733 (N_11733,N_11492,N_11549);
or U11734 (N_11734,N_11513,N_11522);
and U11735 (N_11735,N_11402,N_11582);
and U11736 (N_11736,N_11453,N_11550);
nand U11737 (N_11737,N_11463,N_11600);
nand U11738 (N_11738,N_11575,N_11466);
and U11739 (N_11739,N_11655,N_11422);
xnor U11740 (N_11740,N_11511,N_11635);
or U11741 (N_11741,N_11612,N_11640);
xnor U11742 (N_11742,N_11568,N_11694);
xor U11743 (N_11743,N_11597,N_11495);
nand U11744 (N_11744,N_11510,N_11665);
or U11745 (N_11745,N_11687,N_11689);
and U11746 (N_11746,N_11653,N_11634);
nor U11747 (N_11747,N_11485,N_11584);
and U11748 (N_11748,N_11496,N_11620);
and U11749 (N_11749,N_11677,N_11498);
and U11750 (N_11750,N_11481,N_11666);
xnor U11751 (N_11751,N_11630,N_11633);
nand U11752 (N_11752,N_11450,N_11519);
nand U11753 (N_11753,N_11654,N_11618);
nor U11754 (N_11754,N_11683,N_11409);
nand U11755 (N_11755,N_11447,N_11547);
xnor U11756 (N_11756,N_11539,N_11679);
nor U11757 (N_11757,N_11613,N_11480);
or U11758 (N_11758,N_11668,N_11469);
nand U11759 (N_11759,N_11599,N_11512);
xor U11760 (N_11760,N_11420,N_11484);
nand U11761 (N_11761,N_11464,N_11610);
nor U11762 (N_11762,N_11564,N_11649);
or U11763 (N_11763,N_11488,N_11592);
or U11764 (N_11764,N_11672,N_11542);
and U11765 (N_11765,N_11658,N_11619);
nand U11766 (N_11766,N_11433,N_11541);
xor U11767 (N_11767,N_11692,N_11617);
xor U11768 (N_11768,N_11604,N_11695);
nor U11769 (N_11769,N_11431,N_11499);
nor U11770 (N_11770,N_11537,N_11421);
or U11771 (N_11771,N_11659,N_11457);
and U11772 (N_11772,N_11531,N_11608);
xor U11773 (N_11773,N_11543,N_11468);
nor U11774 (N_11774,N_11681,N_11662);
xor U11775 (N_11775,N_11477,N_11598);
xnor U11776 (N_11776,N_11514,N_11470);
or U11777 (N_11777,N_11698,N_11524);
or U11778 (N_11778,N_11686,N_11660);
xnor U11779 (N_11779,N_11544,N_11534);
and U11780 (N_11780,N_11573,N_11516);
and U11781 (N_11781,N_11552,N_11505);
or U11782 (N_11782,N_11563,N_11540);
xnor U11783 (N_11783,N_11647,N_11491);
xnor U11784 (N_11784,N_11443,N_11478);
nor U11785 (N_11785,N_11611,N_11473);
nor U11786 (N_11786,N_11460,N_11412);
nor U11787 (N_11787,N_11536,N_11590);
and U11788 (N_11788,N_11601,N_11690);
nor U11789 (N_11789,N_11503,N_11415);
and U11790 (N_11790,N_11545,N_11585);
nor U11791 (N_11791,N_11570,N_11502);
nor U11792 (N_11792,N_11626,N_11529);
nor U11793 (N_11793,N_11553,N_11663);
or U11794 (N_11794,N_11518,N_11595);
and U11795 (N_11795,N_11638,N_11527);
nand U11796 (N_11796,N_11643,N_11418);
or U11797 (N_11797,N_11530,N_11571);
nand U11798 (N_11798,N_11438,N_11579);
and U11799 (N_11799,N_11648,N_11423);
or U11800 (N_11800,N_11458,N_11504);
nor U11801 (N_11801,N_11528,N_11525);
xnor U11802 (N_11802,N_11456,N_11407);
xor U11803 (N_11803,N_11603,N_11661);
nor U11804 (N_11804,N_11486,N_11493);
xnor U11805 (N_11805,N_11432,N_11624);
or U11806 (N_11806,N_11674,N_11459);
nor U11807 (N_11807,N_11566,N_11425);
xor U11808 (N_11808,N_11569,N_11594);
nand U11809 (N_11809,N_11567,N_11691);
and U11810 (N_11810,N_11475,N_11572);
xor U11811 (N_11811,N_11629,N_11589);
nor U11812 (N_11812,N_11555,N_11637);
nand U11813 (N_11813,N_11535,N_11628);
or U11814 (N_11814,N_11483,N_11405);
xor U11815 (N_11815,N_11515,N_11441);
nor U11816 (N_11816,N_11556,N_11625);
xnor U11817 (N_11817,N_11419,N_11565);
or U11818 (N_11818,N_11413,N_11557);
and U11819 (N_11819,N_11614,N_11606);
or U11820 (N_11820,N_11623,N_11506);
nand U11821 (N_11821,N_11410,N_11578);
and U11822 (N_11822,N_11482,N_11685);
nor U11823 (N_11823,N_11434,N_11437);
nand U11824 (N_11824,N_11581,N_11471);
xor U11825 (N_11825,N_11487,N_11673);
nand U11826 (N_11826,N_11650,N_11642);
nor U11827 (N_11827,N_11577,N_11586);
nand U11828 (N_11828,N_11621,N_11411);
nor U11829 (N_11829,N_11559,N_11632);
nand U11830 (N_11830,N_11414,N_11508);
or U11831 (N_11831,N_11636,N_11605);
or U11832 (N_11832,N_11560,N_11452);
nor U11833 (N_11833,N_11479,N_11472);
or U11834 (N_11834,N_11427,N_11641);
nand U11835 (N_11835,N_11596,N_11631);
nor U11836 (N_11836,N_11657,N_11671);
nor U11837 (N_11837,N_11670,N_11439);
xor U11838 (N_11838,N_11476,N_11622);
and U11839 (N_11839,N_11474,N_11449);
nor U11840 (N_11840,N_11462,N_11684);
or U11841 (N_11841,N_11697,N_11428);
or U11842 (N_11842,N_11580,N_11602);
xnor U11843 (N_11843,N_11444,N_11448);
nand U11844 (N_11844,N_11408,N_11667);
nand U11845 (N_11845,N_11696,N_11669);
nor U11846 (N_11846,N_11693,N_11538);
nor U11847 (N_11847,N_11465,N_11446);
nor U11848 (N_11848,N_11607,N_11532);
and U11849 (N_11849,N_11416,N_11489);
nand U11850 (N_11850,N_11649,N_11646);
or U11851 (N_11851,N_11633,N_11574);
xor U11852 (N_11852,N_11664,N_11569);
nor U11853 (N_11853,N_11517,N_11519);
nor U11854 (N_11854,N_11643,N_11686);
xnor U11855 (N_11855,N_11531,N_11650);
nor U11856 (N_11856,N_11694,N_11534);
nand U11857 (N_11857,N_11646,N_11639);
xnor U11858 (N_11858,N_11593,N_11666);
or U11859 (N_11859,N_11475,N_11409);
and U11860 (N_11860,N_11544,N_11686);
nand U11861 (N_11861,N_11643,N_11441);
nor U11862 (N_11862,N_11622,N_11449);
nand U11863 (N_11863,N_11627,N_11573);
and U11864 (N_11864,N_11584,N_11445);
or U11865 (N_11865,N_11557,N_11456);
and U11866 (N_11866,N_11653,N_11453);
xor U11867 (N_11867,N_11657,N_11652);
or U11868 (N_11868,N_11416,N_11618);
nand U11869 (N_11869,N_11554,N_11414);
nor U11870 (N_11870,N_11420,N_11421);
nand U11871 (N_11871,N_11426,N_11406);
nor U11872 (N_11872,N_11674,N_11424);
nand U11873 (N_11873,N_11618,N_11436);
nand U11874 (N_11874,N_11610,N_11408);
nor U11875 (N_11875,N_11548,N_11612);
or U11876 (N_11876,N_11582,N_11574);
xor U11877 (N_11877,N_11525,N_11459);
and U11878 (N_11878,N_11668,N_11663);
or U11879 (N_11879,N_11468,N_11631);
or U11880 (N_11880,N_11486,N_11690);
nand U11881 (N_11881,N_11590,N_11414);
or U11882 (N_11882,N_11508,N_11691);
or U11883 (N_11883,N_11480,N_11550);
and U11884 (N_11884,N_11553,N_11614);
xor U11885 (N_11885,N_11534,N_11439);
nand U11886 (N_11886,N_11442,N_11507);
and U11887 (N_11887,N_11515,N_11424);
and U11888 (N_11888,N_11670,N_11471);
nand U11889 (N_11889,N_11539,N_11557);
or U11890 (N_11890,N_11571,N_11549);
and U11891 (N_11891,N_11629,N_11530);
nand U11892 (N_11892,N_11574,N_11571);
xnor U11893 (N_11893,N_11465,N_11597);
and U11894 (N_11894,N_11695,N_11518);
xnor U11895 (N_11895,N_11625,N_11428);
xnor U11896 (N_11896,N_11661,N_11663);
or U11897 (N_11897,N_11431,N_11639);
nor U11898 (N_11898,N_11662,N_11590);
nand U11899 (N_11899,N_11539,N_11410);
and U11900 (N_11900,N_11586,N_11662);
xnor U11901 (N_11901,N_11639,N_11567);
or U11902 (N_11902,N_11561,N_11578);
and U11903 (N_11903,N_11428,N_11403);
xnor U11904 (N_11904,N_11451,N_11663);
nor U11905 (N_11905,N_11657,N_11459);
xor U11906 (N_11906,N_11642,N_11474);
and U11907 (N_11907,N_11540,N_11458);
or U11908 (N_11908,N_11487,N_11611);
nand U11909 (N_11909,N_11499,N_11632);
xnor U11910 (N_11910,N_11576,N_11552);
nand U11911 (N_11911,N_11499,N_11601);
nand U11912 (N_11912,N_11564,N_11422);
xnor U11913 (N_11913,N_11571,N_11638);
or U11914 (N_11914,N_11607,N_11628);
nor U11915 (N_11915,N_11481,N_11418);
nand U11916 (N_11916,N_11652,N_11553);
nand U11917 (N_11917,N_11403,N_11660);
xor U11918 (N_11918,N_11694,N_11645);
and U11919 (N_11919,N_11458,N_11454);
xnor U11920 (N_11920,N_11436,N_11515);
nand U11921 (N_11921,N_11676,N_11555);
and U11922 (N_11922,N_11558,N_11503);
xnor U11923 (N_11923,N_11563,N_11448);
or U11924 (N_11924,N_11593,N_11686);
xor U11925 (N_11925,N_11583,N_11440);
or U11926 (N_11926,N_11592,N_11536);
xnor U11927 (N_11927,N_11424,N_11465);
nand U11928 (N_11928,N_11564,N_11405);
or U11929 (N_11929,N_11533,N_11629);
and U11930 (N_11930,N_11403,N_11418);
nor U11931 (N_11931,N_11455,N_11413);
xor U11932 (N_11932,N_11436,N_11433);
and U11933 (N_11933,N_11508,N_11479);
nor U11934 (N_11934,N_11514,N_11683);
nor U11935 (N_11935,N_11568,N_11675);
and U11936 (N_11936,N_11645,N_11462);
nand U11937 (N_11937,N_11480,N_11582);
nand U11938 (N_11938,N_11691,N_11541);
nand U11939 (N_11939,N_11501,N_11583);
nand U11940 (N_11940,N_11680,N_11479);
nand U11941 (N_11941,N_11641,N_11441);
xor U11942 (N_11942,N_11612,N_11470);
and U11943 (N_11943,N_11619,N_11474);
and U11944 (N_11944,N_11425,N_11421);
nand U11945 (N_11945,N_11424,N_11625);
and U11946 (N_11946,N_11694,N_11536);
or U11947 (N_11947,N_11497,N_11583);
nor U11948 (N_11948,N_11680,N_11458);
nor U11949 (N_11949,N_11681,N_11618);
or U11950 (N_11950,N_11460,N_11653);
nand U11951 (N_11951,N_11581,N_11461);
nor U11952 (N_11952,N_11619,N_11516);
or U11953 (N_11953,N_11653,N_11651);
or U11954 (N_11954,N_11530,N_11513);
nor U11955 (N_11955,N_11432,N_11420);
nor U11956 (N_11956,N_11522,N_11439);
and U11957 (N_11957,N_11643,N_11499);
xor U11958 (N_11958,N_11429,N_11478);
nand U11959 (N_11959,N_11524,N_11455);
nor U11960 (N_11960,N_11403,N_11408);
or U11961 (N_11961,N_11573,N_11519);
nor U11962 (N_11962,N_11676,N_11610);
xnor U11963 (N_11963,N_11455,N_11656);
nor U11964 (N_11964,N_11572,N_11441);
or U11965 (N_11965,N_11497,N_11664);
and U11966 (N_11966,N_11605,N_11633);
xnor U11967 (N_11967,N_11582,N_11444);
nand U11968 (N_11968,N_11472,N_11432);
xnor U11969 (N_11969,N_11662,N_11424);
xnor U11970 (N_11970,N_11498,N_11633);
nor U11971 (N_11971,N_11473,N_11591);
or U11972 (N_11972,N_11452,N_11617);
xnor U11973 (N_11973,N_11665,N_11421);
xnor U11974 (N_11974,N_11605,N_11486);
and U11975 (N_11975,N_11534,N_11489);
xor U11976 (N_11976,N_11514,N_11532);
nor U11977 (N_11977,N_11516,N_11488);
xor U11978 (N_11978,N_11413,N_11486);
nor U11979 (N_11979,N_11403,N_11662);
nand U11980 (N_11980,N_11441,N_11402);
and U11981 (N_11981,N_11563,N_11566);
nand U11982 (N_11982,N_11511,N_11692);
nand U11983 (N_11983,N_11413,N_11506);
nand U11984 (N_11984,N_11615,N_11630);
and U11985 (N_11985,N_11507,N_11683);
nand U11986 (N_11986,N_11425,N_11616);
xor U11987 (N_11987,N_11650,N_11670);
and U11988 (N_11988,N_11585,N_11531);
or U11989 (N_11989,N_11527,N_11561);
and U11990 (N_11990,N_11658,N_11645);
or U11991 (N_11991,N_11448,N_11630);
or U11992 (N_11992,N_11483,N_11605);
and U11993 (N_11993,N_11519,N_11515);
or U11994 (N_11994,N_11674,N_11613);
or U11995 (N_11995,N_11583,N_11494);
nand U11996 (N_11996,N_11404,N_11462);
or U11997 (N_11997,N_11536,N_11422);
xor U11998 (N_11998,N_11488,N_11405);
nor U11999 (N_11999,N_11596,N_11578);
or U12000 (N_12000,N_11945,N_11883);
nand U12001 (N_12001,N_11745,N_11862);
xor U12002 (N_12002,N_11722,N_11987);
xor U12003 (N_12003,N_11938,N_11819);
xor U12004 (N_12004,N_11820,N_11931);
and U12005 (N_12005,N_11858,N_11876);
or U12006 (N_12006,N_11951,N_11997);
nand U12007 (N_12007,N_11981,N_11793);
nand U12008 (N_12008,N_11720,N_11779);
nand U12009 (N_12009,N_11724,N_11914);
or U12010 (N_12010,N_11888,N_11837);
and U12011 (N_12011,N_11977,N_11864);
or U12012 (N_12012,N_11832,N_11901);
nor U12013 (N_12013,N_11831,N_11767);
and U12014 (N_12014,N_11940,N_11775);
xnor U12015 (N_12015,N_11821,N_11899);
or U12016 (N_12016,N_11814,N_11882);
xnor U12017 (N_12017,N_11941,N_11895);
nor U12018 (N_12018,N_11869,N_11952);
or U12019 (N_12019,N_11826,N_11985);
nor U12020 (N_12020,N_11906,N_11969);
xnor U12021 (N_12021,N_11743,N_11840);
nand U12022 (N_12022,N_11933,N_11991);
or U12023 (N_12023,N_11885,N_11828);
or U12024 (N_12024,N_11884,N_11732);
xor U12025 (N_12025,N_11872,N_11972);
or U12026 (N_12026,N_11966,N_11741);
and U12027 (N_12027,N_11849,N_11769);
nor U12028 (N_12028,N_11776,N_11935);
and U12029 (N_12029,N_11746,N_11948);
or U12030 (N_12030,N_11911,N_11829);
xnor U12031 (N_12031,N_11833,N_11996);
xor U12032 (N_12032,N_11890,N_11807);
nand U12033 (N_12033,N_11727,N_11801);
xnor U12034 (N_12034,N_11762,N_11866);
xnor U12035 (N_12035,N_11980,N_11960);
or U12036 (N_12036,N_11763,N_11770);
nor U12037 (N_12037,N_11706,N_11708);
nand U12038 (N_12038,N_11915,N_11792);
or U12039 (N_12039,N_11744,N_11822);
and U12040 (N_12040,N_11738,N_11843);
and U12041 (N_12041,N_11873,N_11971);
and U12042 (N_12042,N_11936,N_11982);
or U12043 (N_12043,N_11797,N_11900);
xnor U12044 (N_12044,N_11714,N_11859);
nor U12045 (N_12045,N_11925,N_11943);
xor U12046 (N_12046,N_11845,N_11910);
xnor U12047 (N_12047,N_11789,N_11749);
xor U12048 (N_12048,N_11932,N_11913);
and U12049 (N_12049,N_11944,N_11755);
and U12050 (N_12050,N_11817,N_11717);
or U12051 (N_12051,N_11973,N_11855);
nor U12052 (N_12052,N_11927,N_11711);
or U12053 (N_12053,N_11761,N_11897);
nand U12054 (N_12054,N_11988,N_11947);
and U12055 (N_12055,N_11902,N_11918);
xnor U12056 (N_12056,N_11752,N_11841);
or U12057 (N_12057,N_11986,N_11715);
or U12058 (N_12058,N_11788,N_11889);
and U12059 (N_12059,N_11928,N_11796);
nor U12060 (N_12060,N_11959,N_11846);
and U12061 (N_12061,N_11879,N_11750);
and U12062 (N_12062,N_11787,N_11860);
nor U12063 (N_12063,N_11999,N_11754);
or U12064 (N_12064,N_11892,N_11772);
or U12065 (N_12065,N_11707,N_11856);
nand U12066 (N_12066,N_11835,N_11937);
nand U12067 (N_12067,N_11810,N_11736);
nand U12068 (N_12068,N_11823,N_11783);
nor U12069 (N_12069,N_11909,N_11734);
nor U12070 (N_12070,N_11838,N_11989);
nand U12071 (N_12071,N_11993,N_11992);
or U12072 (N_12072,N_11848,N_11771);
xor U12073 (N_12073,N_11861,N_11851);
xor U12074 (N_12074,N_11842,N_11868);
xor U12075 (N_12075,N_11963,N_11757);
nor U12076 (N_12076,N_11917,N_11766);
xor U12077 (N_12077,N_11733,N_11854);
nand U12078 (N_12078,N_11791,N_11967);
and U12079 (N_12079,N_11781,N_11800);
xnor U12080 (N_12080,N_11984,N_11764);
nor U12081 (N_12081,N_11923,N_11773);
or U12082 (N_12082,N_11922,N_11924);
or U12083 (N_12083,N_11825,N_11799);
and U12084 (N_12084,N_11974,N_11718);
or U12085 (N_12085,N_11812,N_11780);
xnor U12086 (N_12086,N_11953,N_11893);
nand U12087 (N_12087,N_11768,N_11785);
or U12088 (N_12088,N_11920,N_11836);
xor U12089 (N_12089,N_11808,N_11905);
or U12090 (N_12090,N_11921,N_11970);
and U12091 (N_12091,N_11705,N_11976);
and U12092 (N_12092,N_11908,N_11839);
and U12093 (N_12093,N_11904,N_11703);
xor U12094 (N_12094,N_11875,N_11994);
nor U12095 (N_12095,N_11930,N_11874);
or U12096 (N_12096,N_11894,N_11815);
nand U12097 (N_12097,N_11853,N_11739);
or U12098 (N_12098,N_11730,N_11760);
and U12099 (N_12099,N_11979,N_11995);
xor U12100 (N_12100,N_11811,N_11954);
and U12101 (N_12101,N_11751,N_11735);
or U12102 (N_12102,N_11975,N_11809);
nor U12103 (N_12103,N_11737,N_11742);
or U12104 (N_12104,N_11778,N_11844);
or U12105 (N_12105,N_11896,N_11723);
xnor U12106 (N_12106,N_11962,N_11891);
or U12107 (N_12107,N_11813,N_11958);
or U12108 (N_12108,N_11965,N_11867);
and U12109 (N_12109,N_11804,N_11961);
xnor U12110 (N_12110,N_11827,N_11955);
nor U12111 (N_12111,N_11926,N_11794);
nand U12112 (N_12112,N_11716,N_11700);
nor U12113 (N_12113,N_11847,N_11704);
or U12114 (N_12114,N_11950,N_11878);
nor U12115 (N_12115,N_11729,N_11712);
or U12116 (N_12116,N_11824,N_11949);
xor U12117 (N_12117,N_11850,N_11834);
or U12118 (N_12118,N_11725,N_11790);
and U12119 (N_12119,N_11774,N_11957);
nand U12120 (N_12120,N_11784,N_11710);
nand U12121 (N_12121,N_11721,N_11740);
and U12122 (N_12122,N_11726,N_11934);
nand U12123 (N_12123,N_11956,N_11765);
nand U12124 (N_12124,N_11857,N_11898);
nor U12125 (N_12125,N_11805,N_11758);
nand U12126 (N_12126,N_11916,N_11887);
xnor U12127 (N_12127,N_11871,N_11702);
and U12128 (N_12128,N_11912,N_11777);
nand U12129 (N_12129,N_11803,N_11990);
nor U12130 (N_12130,N_11753,N_11863);
nand U12131 (N_12131,N_11795,N_11818);
and U12132 (N_12132,N_11719,N_11852);
xnor U12133 (N_12133,N_11759,N_11903);
nor U12134 (N_12134,N_11946,N_11939);
or U12135 (N_12135,N_11802,N_11983);
nand U12136 (N_12136,N_11756,N_11806);
or U12137 (N_12137,N_11798,N_11728);
xnor U12138 (N_12138,N_11877,N_11998);
or U12139 (N_12139,N_11709,N_11881);
nand U12140 (N_12140,N_11816,N_11919);
nor U12141 (N_12141,N_11942,N_11701);
or U12142 (N_12142,N_11731,N_11748);
nand U12143 (N_12143,N_11968,N_11830);
xor U12144 (N_12144,N_11880,N_11978);
nor U12145 (N_12145,N_11907,N_11786);
nor U12146 (N_12146,N_11782,N_11870);
nand U12147 (N_12147,N_11865,N_11929);
and U12148 (N_12148,N_11713,N_11747);
and U12149 (N_12149,N_11886,N_11964);
xor U12150 (N_12150,N_11977,N_11948);
or U12151 (N_12151,N_11979,N_11773);
nand U12152 (N_12152,N_11931,N_11964);
or U12153 (N_12153,N_11951,N_11982);
or U12154 (N_12154,N_11850,N_11965);
nand U12155 (N_12155,N_11713,N_11890);
xor U12156 (N_12156,N_11941,N_11750);
or U12157 (N_12157,N_11922,N_11874);
and U12158 (N_12158,N_11991,N_11967);
xnor U12159 (N_12159,N_11901,N_11821);
nand U12160 (N_12160,N_11995,N_11849);
or U12161 (N_12161,N_11821,N_11936);
or U12162 (N_12162,N_11915,N_11745);
nor U12163 (N_12163,N_11888,N_11776);
nor U12164 (N_12164,N_11932,N_11756);
nand U12165 (N_12165,N_11977,N_11978);
nand U12166 (N_12166,N_11875,N_11822);
nand U12167 (N_12167,N_11720,N_11863);
or U12168 (N_12168,N_11969,N_11865);
nand U12169 (N_12169,N_11966,N_11855);
nor U12170 (N_12170,N_11884,N_11735);
xnor U12171 (N_12171,N_11952,N_11859);
nand U12172 (N_12172,N_11914,N_11881);
or U12173 (N_12173,N_11751,N_11775);
nor U12174 (N_12174,N_11844,N_11773);
and U12175 (N_12175,N_11844,N_11922);
nor U12176 (N_12176,N_11752,N_11774);
nand U12177 (N_12177,N_11965,N_11702);
nand U12178 (N_12178,N_11767,N_11922);
and U12179 (N_12179,N_11737,N_11927);
and U12180 (N_12180,N_11765,N_11826);
or U12181 (N_12181,N_11825,N_11934);
nand U12182 (N_12182,N_11912,N_11891);
nand U12183 (N_12183,N_11944,N_11989);
or U12184 (N_12184,N_11701,N_11845);
nand U12185 (N_12185,N_11983,N_11885);
nand U12186 (N_12186,N_11981,N_11926);
nor U12187 (N_12187,N_11836,N_11717);
xnor U12188 (N_12188,N_11930,N_11975);
and U12189 (N_12189,N_11858,N_11815);
and U12190 (N_12190,N_11747,N_11841);
and U12191 (N_12191,N_11898,N_11721);
or U12192 (N_12192,N_11957,N_11820);
nand U12193 (N_12193,N_11709,N_11815);
nand U12194 (N_12194,N_11989,N_11815);
nor U12195 (N_12195,N_11844,N_11785);
or U12196 (N_12196,N_11772,N_11828);
and U12197 (N_12197,N_11876,N_11845);
nand U12198 (N_12198,N_11923,N_11714);
nor U12199 (N_12199,N_11862,N_11844);
or U12200 (N_12200,N_11929,N_11986);
nand U12201 (N_12201,N_11875,N_11800);
nand U12202 (N_12202,N_11938,N_11809);
nand U12203 (N_12203,N_11895,N_11776);
or U12204 (N_12204,N_11998,N_11762);
xor U12205 (N_12205,N_11952,N_11877);
nor U12206 (N_12206,N_11866,N_11725);
and U12207 (N_12207,N_11712,N_11885);
and U12208 (N_12208,N_11885,N_11812);
and U12209 (N_12209,N_11816,N_11829);
xor U12210 (N_12210,N_11932,N_11766);
xor U12211 (N_12211,N_11711,N_11729);
nand U12212 (N_12212,N_11899,N_11943);
nand U12213 (N_12213,N_11952,N_11825);
or U12214 (N_12214,N_11973,N_11919);
nand U12215 (N_12215,N_11923,N_11835);
xnor U12216 (N_12216,N_11992,N_11738);
xor U12217 (N_12217,N_11784,N_11803);
and U12218 (N_12218,N_11784,N_11976);
or U12219 (N_12219,N_11846,N_11770);
or U12220 (N_12220,N_11851,N_11707);
nor U12221 (N_12221,N_11967,N_11731);
and U12222 (N_12222,N_11742,N_11703);
nand U12223 (N_12223,N_11701,N_11824);
nand U12224 (N_12224,N_11824,N_11997);
or U12225 (N_12225,N_11709,N_11789);
nand U12226 (N_12226,N_11988,N_11819);
nor U12227 (N_12227,N_11719,N_11963);
and U12228 (N_12228,N_11889,N_11909);
nand U12229 (N_12229,N_11743,N_11957);
nand U12230 (N_12230,N_11858,N_11828);
or U12231 (N_12231,N_11721,N_11763);
nor U12232 (N_12232,N_11958,N_11899);
or U12233 (N_12233,N_11983,N_11954);
nand U12234 (N_12234,N_11804,N_11939);
nand U12235 (N_12235,N_11912,N_11991);
and U12236 (N_12236,N_11830,N_11871);
nor U12237 (N_12237,N_11928,N_11789);
nor U12238 (N_12238,N_11757,N_11889);
nor U12239 (N_12239,N_11925,N_11703);
and U12240 (N_12240,N_11996,N_11923);
nor U12241 (N_12241,N_11987,N_11703);
and U12242 (N_12242,N_11940,N_11746);
and U12243 (N_12243,N_11863,N_11758);
xor U12244 (N_12244,N_11766,N_11974);
or U12245 (N_12245,N_11789,N_11712);
xnor U12246 (N_12246,N_11808,N_11801);
nand U12247 (N_12247,N_11885,N_11818);
nand U12248 (N_12248,N_11943,N_11906);
xnor U12249 (N_12249,N_11990,N_11907);
nor U12250 (N_12250,N_11774,N_11827);
or U12251 (N_12251,N_11866,N_11911);
nand U12252 (N_12252,N_11783,N_11857);
and U12253 (N_12253,N_11870,N_11727);
or U12254 (N_12254,N_11822,N_11748);
and U12255 (N_12255,N_11778,N_11878);
nor U12256 (N_12256,N_11738,N_11785);
or U12257 (N_12257,N_11807,N_11898);
nor U12258 (N_12258,N_11824,N_11753);
xnor U12259 (N_12259,N_11753,N_11942);
xnor U12260 (N_12260,N_11701,N_11856);
or U12261 (N_12261,N_11798,N_11883);
or U12262 (N_12262,N_11969,N_11778);
nand U12263 (N_12263,N_11883,N_11956);
xnor U12264 (N_12264,N_11774,N_11780);
or U12265 (N_12265,N_11935,N_11925);
xor U12266 (N_12266,N_11747,N_11905);
nor U12267 (N_12267,N_11998,N_11966);
nand U12268 (N_12268,N_11983,N_11982);
and U12269 (N_12269,N_11843,N_11896);
or U12270 (N_12270,N_11924,N_11966);
nand U12271 (N_12271,N_11952,N_11741);
or U12272 (N_12272,N_11816,N_11968);
nor U12273 (N_12273,N_11795,N_11865);
xnor U12274 (N_12274,N_11780,N_11719);
or U12275 (N_12275,N_11899,N_11963);
and U12276 (N_12276,N_11777,N_11867);
and U12277 (N_12277,N_11890,N_11707);
xnor U12278 (N_12278,N_11808,N_11814);
or U12279 (N_12279,N_11917,N_11738);
nand U12280 (N_12280,N_11710,N_11865);
xor U12281 (N_12281,N_11951,N_11748);
nand U12282 (N_12282,N_11863,N_11915);
nor U12283 (N_12283,N_11912,N_11735);
and U12284 (N_12284,N_11939,N_11809);
and U12285 (N_12285,N_11937,N_11760);
xnor U12286 (N_12286,N_11713,N_11802);
or U12287 (N_12287,N_11893,N_11909);
and U12288 (N_12288,N_11708,N_11915);
or U12289 (N_12289,N_11714,N_11961);
xor U12290 (N_12290,N_11788,N_11904);
xor U12291 (N_12291,N_11754,N_11895);
and U12292 (N_12292,N_11926,N_11934);
or U12293 (N_12293,N_11846,N_11710);
nor U12294 (N_12294,N_11789,N_11924);
nand U12295 (N_12295,N_11753,N_11850);
and U12296 (N_12296,N_11825,N_11985);
or U12297 (N_12297,N_11722,N_11849);
or U12298 (N_12298,N_11918,N_11709);
or U12299 (N_12299,N_11788,N_11983);
xor U12300 (N_12300,N_12204,N_12220);
and U12301 (N_12301,N_12136,N_12199);
xor U12302 (N_12302,N_12277,N_12066);
or U12303 (N_12303,N_12171,N_12144);
nand U12304 (N_12304,N_12002,N_12242);
or U12305 (N_12305,N_12124,N_12182);
and U12306 (N_12306,N_12018,N_12109);
and U12307 (N_12307,N_12013,N_12234);
nor U12308 (N_12308,N_12223,N_12202);
xor U12309 (N_12309,N_12232,N_12226);
nand U12310 (N_12310,N_12095,N_12032);
xnor U12311 (N_12311,N_12150,N_12246);
nor U12312 (N_12312,N_12010,N_12167);
nor U12313 (N_12313,N_12163,N_12101);
nor U12314 (N_12314,N_12156,N_12184);
nand U12315 (N_12315,N_12086,N_12021);
nor U12316 (N_12316,N_12281,N_12123);
and U12317 (N_12317,N_12026,N_12174);
and U12318 (N_12318,N_12057,N_12161);
nand U12319 (N_12319,N_12071,N_12213);
xor U12320 (N_12320,N_12117,N_12279);
and U12321 (N_12321,N_12225,N_12203);
and U12322 (N_12322,N_12272,N_12231);
or U12323 (N_12323,N_12168,N_12129);
or U12324 (N_12324,N_12290,N_12227);
or U12325 (N_12325,N_12073,N_12005);
nor U12326 (N_12326,N_12075,N_12282);
nand U12327 (N_12327,N_12244,N_12169);
nor U12328 (N_12328,N_12023,N_12230);
and U12329 (N_12329,N_12015,N_12056);
nor U12330 (N_12330,N_12110,N_12119);
or U12331 (N_12331,N_12084,N_12143);
nor U12332 (N_12332,N_12134,N_12068);
or U12333 (N_12333,N_12130,N_12160);
nand U12334 (N_12334,N_12042,N_12116);
nand U12335 (N_12335,N_12122,N_12141);
and U12336 (N_12336,N_12022,N_12082);
nor U12337 (N_12337,N_12051,N_12081);
or U12338 (N_12338,N_12236,N_12256);
or U12339 (N_12339,N_12025,N_12205);
nand U12340 (N_12340,N_12218,N_12271);
xor U12341 (N_12341,N_12197,N_12054);
nand U12342 (N_12342,N_12003,N_12243);
or U12343 (N_12343,N_12036,N_12200);
nor U12344 (N_12344,N_12299,N_12052);
and U12345 (N_12345,N_12240,N_12046);
and U12346 (N_12346,N_12099,N_12206);
xnor U12347 (N_12347,N_12148,N_12019);
xor U12348 (N_12348,N_12270,N_12153);
or U12349 (N_12349,N_12298,N_12191);
xor U12350 (N_12350,N_12280,N_12139);
nand U12351 (N_12351,N_12102,N_12009);
nor U12352 (N_12352,N_12105,N_12255);
and U12353 (N_12353,N_12014,N_12106);
or U12354 (N_12354,N_12112,N_12078);
nor U12355 (N_12355,N_12267,N_12048);
xor U12356 (N_12356,N_12120,N_12088);
nand U12357 (N_12357,N_12083,N_12107);
nand U12358 (N_12358,N_12050,N_12257);
nand U12359 (N_12359,N_12175,N_12104);
nand U12360 (N_12360,N_12121,N_12170);
nand U12361 (N_12361,N_12211,N_12189);
nand U12362 (N_12362,N_12193,N_12135);
xnor U12363 (N_12363,N_12162,N_12024);
nand U12364 (N_12364,N_12152,N_12038);
nor U12365 (N_12365,N_12288,N_12297);
xor U12366 (N_12366,N_12286,N_12233);
xor U12367 (N_12367,N_12201,N_12064);
nand U12368 (N_12368,N_12004,N_12185);
nor U12369 (N_12369,N_12035,N_12049);
and U12370 (N_12370,N_12254,N_12079);
nor U12371 (N_12371,N_12179,N_12149);
or U12372 (N_12372,N_12069,N_12118);
xor U12373 (N_12373,N_12262,N_12284);
or U12374 (N_12374,N_12132,N_12289);
xnor U12375 (N_12375,N_12138,N_12017);
nor U12376 (N_12376,N_12198,N_12154);
or U12377 (N_12377,N_12195,N_12011);
nor U12378 (N_12378,N_12251,N_12166);
nor U12379 (N_12379,N_12228,N_12151);
and U12380 (N_12380,N_12261,N_12158);
xnor U12381 (N_12381,N_12089,N_12007);
xor U12382 (N_12382,N_12207,N_12000);
nor U12383 (N_12383,N_12239,N_12173);
and U12384 (N_12384,N_12012,N_12027);
or U12385 (N_12385,N_12028,N_12097);
nand U12386 (N_12386,N_12178,N_12180);
xnor U12387 (N_12387,N_12133,N_12275);
nand U12388 (N_12388,N_12142,N_12033);
nand U12389 (N_12389,N_12128,N_12287);
nor U12390 (N_12390,N_12253,N_12060);
and U12391 (N_12391,N_12031,N_12269);
or U12392 (N_12392,N_12145,N_12008);
and U12393 (N_12393,N_12181,N_12126);
and U12394 (N_12394,N_12065,N_12268);
and U12395 (N_12395,N_12020,N_12029);
xnor U12396 (N_12396,N_12194,N_12094);
and U12397 (N_12397,N_12186,N_12229);
xor U12398 (N_12398,N_12278,N_12072);
nand U12399 (N_12399,N_12146,N_12045);
xnor U12400 (N_12400,N_12214,N_12210);
xnor U12401 (N_12401,N_12062,N_12115);
nor U12402 (N_12402,N_12067,N_12157);
and U12403 (N_12403,N_12040,N_12291);
and U12404 (N_12404,N_12030,N_12241);
and U12405 (N_12405,N_12209,N_12237);
and U12406 (N_12406,N_12285,N_12016);
and U12407 (N_12407,N_12219,N_12187);
nand U12408 (N_12408,N_12212,N_12165);
xnor U12409 (N_12409,N_12238,N_12006);
xor U12410 (N_12410,N_12070,N_12252);
or U12411 (N_12411,N_12147,N_12001);
nand U12412 (N_12412,N_12063,N_12125);
nor U12413 (N_12413,N_12058,N_12039);
nand U12414 (N_12414,N_12164,N_12235);
xor U12415 (N_12415,N_12249,N_12108);
or U12416 (N_12416,N_12091,N_12183);
or U12417 (N_12417,N_12208,N_12041);
and U12418 (N_12418,N_12127,N_12215);
and U12419 (N_12419,N_12096,N_12293);
nand U12420 (N_12420,N_12224,N_12276);
and U12421 (N_12421,N_12188,N_12295);
nand U12422 (N_12422,N_12172,N_12103);
or U12423 (N_12423,N_12217,N_12100);
nor U12424 (N_12424,N_12114,N_12034);
xor U12425 (N_12425,N_12259,N_12221);
or U12426 (N_12426,N_12131,N_12159);
xnor U12427 (N_12427,N_12077,N_12292);
or U12428 (N_12428,N_12093,N_12250);
and U12429 (N_12429,N_12264,N_12140);
and U12430 (N_12430,N_12190,N_12055);
or U12431 (N_12431,N_12266,N_12059);
or U12432 (N_12432,N_12047,N_12247);
and U12433 (N_12433,N_12176,N_12177);
nor U12434 (N_12434,N_12265,N_12258);
nor U12435 (N_12435,N_12098,N_12137);
and U12436 (N_12436,N_12222,N_12044);
xnor U12437 (N_12437,N_12061,N_12248);
xor U12438 (N_12438,N_12087,N_12245);
nor U12439 (N_12439,N_12074,N_12085);
or U12440 (N_12440,N_12273,N_12113);
nor U12441 (N_12441,N_12080,N_12196);
xor U12442 (N_12442,N_12294,N_12260);
nor U12443 (N_12443,N_12192,N_12155);
nand U12444 (N_12444,N_12090,N_12296);
or U12445 (N_12445,N_12283,N_12263);
and U12446 (N_12446,N_12076,N_12274);
nor U12447 (N_12447,N_12111,N_12037);
and U12448 (N_12448,N_12043,N_12053);
xnor U12449 (N_12449,N_12092,N_12216);
nor U12450 (N_12450,N_12171,N_12219);
xnor U12451 (N_12451,N_12272,N_12058);
nor U12452 (N_12452,N_12011,N_12279);
nand U12453 (N_12453,N_12187,N_12294);
nand U12454 (N_12454,N_12285,N_12128);
xnor U12455 (N_12455,N_12143,N_12158);
nand U12456 (N_12456,N_12288,N_12104);
and U12457 (N_12457,N_12096,N_12273);
nor U12458 (N_12458,N_12034,N_12138);
nand U12459 (N_12459,N_12164,N_12136);
and U12460 (N_12460,N_12220,N_12224);
nor U12461 (N_12461,N_12050,N_12245);
nand U12462 (N_12462,N_12128,N_12215);
or U12463 (N_12463,N_12171,N_12109);
xnor U12464 (N_12464,N_12066,N_12021);
and U12465 (N_12465,N_12087,N_12056);
and U12466 (N_12466,N_12136,N_12030);
or U12467 (N_12467,N_12051,N_12066);
nor U12468 (N_12468,N_12288,N_12089);
xnor U12469 (N_12469,N_12216,N_12230);
or U12470 (N_12470,N_12225,N_12075);
nand U12471 (N_12471,N_12295,N_12202);
xor U12472 (N_12472,N_12271,N_12281);
xnor U12473 (N_12473,N_12108,N_12039);
nand U12474 (N_12474,N_12117,N_12297);
nand U12475 (N_12475,N_12041,N_12134);
and U12476 (N_12476,N_12158,N_12165);
xnor U12477 (N_12477,N_12031,N_12101);
and U12478 (N_12478,N_12079,N_12224);
nor U12479 (N_12479,N_12296,N_12259);
nor U12480 (N_12480,N_12042,N_12177);
nand U12481 (N_12481,N_12157,N_12170);
or U12482 (N_12482,N_12154,N_12189);
nor U12483 (N_12483,N_12047,N_12133);
nand U12484 (N_12484,N_12266,N_12114);
or U12485 (N_12485,N_12121,N_12297);
nand U12486 (N_12486,N_12226,N_12032);
nor U12487 (N_12487,N_12110,N_12210);
or U12488 (N_12488,N_12031,N_12273);
and U12489 (N_12489,N_12126,N_12164);
nand U12490 (N_12490,N_12083,N_12085);
xor U12491 (N_12491,N_12066,N_12187);
and U12492 (N_12492,N_12074,N_12299);
and U12493 (N_12493,N_12109,N_12203);
xnor U12494 (N_12494,N_12041,N_12094);
and U12495 (N_12495,N_12137,N_12022);
nand U12496 (N_12496,N_12128,N_12183);
and U12497 (N_12497,N_12097,N_12015);
xnor U12498 (N_12498,N_12226,N_12176);
or U12499 (N_12499,N_12006,N_12063);
xnor U12500 (N_12500,N_12227,N_12034);
or U12501 (N_12501,N_12256,N_12102);
or U12502 (N_12502,N_12158,N_12249);
nand U12503 (N_12503,N_12057,N_12126);
xnor U12504 (N_12504,N_12292,N_12099);
or U12505 (N_12505,N_12050,N_12204);
or U12506 (N_12506,N_12041,N_12256);
nor U12507 (N_12507,N_12082,N_12096);
nand U12508 (N_12508,N_12089,N_12102);
xor U12509 (N_12509,N_12079,N_12249);
nor U12510 (N_12510,N_12114,N_12069);
and U12511 (N_12511,N_12234,N_12099);
or U12512 (N_12512,N_12137,N_12238);
nor U12513 (N_12513,N_12037,N_12298);
or U12514 (N_12514,N_12153,N_12257);
and U12515 (N_12515,N_12229,N_12040);
and U12516 (N_12516,N_12004,N_12296);
nand U12517 (N_12517,N_12246,N_12145);
and U12518 (N_12518,N_12263,N_12108);
or U12519 (N_12519,N_12144,N_12127);
and U12520 (N_12520,N_12030,N_12107);
and U12521 (N_12521,N_12034,N_12280);
xor U12522 (N_12522,N_12173,N_12000);
or U12523 (N_12523,N_12228,N_12046);
nor U12524 (N_12524,N_12041,N_12124);
or U12525 (N_12525,N_12039,N_12213);
xor U12526 (N_12526,N_12138,N_12000);
or U12527 (N_12527,N_12239,N_12049);
xor U12528 (N_12528,N_12256,N_12250);
nor U12529 (N_12529,N_12001,N_12085);
xor U12530 (N_12530,N_12262,N_12202);
nor U12531 (N_12531,N_12053,N_12145);
nor U12532 (N_12532,N_12264,N_12236);
nor U12533 (N_12533,N_12025,N_12178);
xor U12534 (N_12534,N_12206,N_12031);
xnor U12535 (N_12535,N_12242,N_12040);
and U12536 (N_12536,N_12286,N_12277);
and U12537 (N_12537,N_12272,N_12137);
nor U12538 (N_12538,N_12229,N_12060);
and U12539 (N_12539,N_12290,N_12109);
and U12540 (N_12540,N_12131,N_12207);
nor U12541 (N_12541,N_12195,N_12264);
nand U12542 (N_12542,N_12069,N_12062);
and U12543 (N_12543,N_12196,N_12164);
xor U12544 (N_12544,N_12082,N_12283);
xor U12545 (N_12545,N_12068,N_12159);
or U12546 (N_12546,N_12127,N_12228);
nand U12547 (N_12547,N_12140,N_12063);
and U12548 (N_12548,N_12275,N_12236);
or U12549 (N_12549,N_12004,N_12029);
or U12550 (N_12550,N_12101,N_12027);
and U12551 (N_12551,N_12045,N_12000);
nor U12552 (N_12552,N_12198,N_12073);
and U12553 (N_12553,N_12288,N_12135);
nand U12554 (N_12554,N_12064,N_12096);
nor U12555 (N_12555,N_12205,N_12154);
and U12556 (N_12556,N_12076,N_12149);
nor U12557 (N_12557,N_12144,N_12227);
nand U12558 (N_12558,N_12071,N_12077);
and U12559 (N_12559,N_12226,N_12080);
and U12560 (N_12560,N_12065,N_12163);
xor U12561 (N_12561,N_12257,N_12219);
and U12562 (N_12562,N_12052,N_12005);
xnor U12563 (N_12563,N_12155,N_12180);
or U12564 (N_12564,N_12246,N_12015);
and U12565 (N_12565,N_12297,N_12040);
or U12566 (N_12566,N_12164,N_12081);
or U12567 (N_12567,N_12142,N_12026);
nand U12568 (N_12568,N_12134,N_12197);
xnor U12569 (N_12569,N_12023,N_12034);
nor U12570 (N_12570,N_12261,N_12248);
and U12571 (N_12571,N_12241,N_12170);
or U12572 (N_12572,N_12057,N_12194);
xnor U12573 (N_12573,N_12268,N_12106);
and U12574 (N_12574,N_12150,N_12100);
nor U12575 (N_12575,N_12066,N_12152);
and U12576 (N_12576,N_12121,N_12113);
nor U12577 (N_12577,N_12080,N_12045);
xor U12578 (N_12578,N_12290,N_12169);
and U12579 (N_12579,N_12010,N_12221);
nand U12580 (N_12580,N_12134,N_12028);
and U12581 (N_12581,N_12191,N_12187);
nand U12582 (N_12582,N_12013,N_12041);
xor U12583 (N_12583,N_12066,N_12135);
nand U12584 (N_12584,N_12113,N_12177);
nor U12585 (N_12585,N_12036,N_12270);
xnor U12586 (N_12586,N_12096,N_12290);
or U12587 (N_12587,N_12296,N_12035);
xor U12588 (N_12588,N_12128,N_12008);
nor U12589 (N_12589,N_12297,N_12206);
and U12590 (N_12590,N_12227,N_12271);
or U12591 (N_12591,N_12138,N_12109);
nand U12592 (N_12592,N_12113,N_12016);
or U12593 (N_12593,N_12202,N_12273);
nor U12594 (N_12594,N_12068,N_12146);
or U12595 (N_12595,N_12056,N_12094);
nand U12596 (N_12596,N_12285,N_12275);
or U12597 (N_12597,N_12231,N_12074);
nand U12598 (N_12598,N_12141,N_12251);
nor U12599 (N_12599,N_12273,N_12292);
nor U12600 (N_12600,N_12474,N_12561);
nor U12601 (N_12601,N_12354,N_12520);
and U12602 (N_12602,N_12545,N_12502);
nand U12603 (N_12603,N_12459,N_12467);
or U12604 (N_12604,N_12440,N_12344);
nand U12605 (N_12605,N_12300,N_12495);
nor U12606 (N_12606,N_12347,N_12585);
and U12607 (N_12607,N_12444,N_12497);
nor U12608 (N_12608,N_12352,N_12567);
nor U12609 (N_12609,N_12505,N_12499);
and U12610 (N_12610,N_12451,N_12389);
or U12611 (N_12611,N_12583,N_12428);
nor U12612 (N_12612,N_12586,N_12598);
or U12613 (N_12613,N_12446,N_12582);
or U12614 (N_12614,N_12330,N_12532);
nor U12615 (N_12615,N_12388,N_12531);
nor U12616 (N_12616,N_12469,N_12527);
or U12617 (N_12617,N_12595,N_12562);
nor U12618 (N_12618,N_12552,N_12305);
xnor U12619 (N_12619,N_12405,N_12362);
nor U12620 (N_12620,N_12471,N_12336);
or U12621 (N_12621,N_12434,N_12303);
xnor U12622 (N_12622,N_12521,N_12413);
nor U12623 (N_12623,N_12417,N_12569);
xor U12624 (N_12624,N_12316,N_12307);
xnor U12625 (N_12625,N_12309,N_12439);
and U12626 (N_12626,N_12516,N_12327);
xor U12627 (N_12627,N_12512,N_12543);
nand U12628 (N_12628,N_12554,N_12436);
and U12629 (N_12629,N_12523,N_12489);
nor U12630 (N_12630,N_12461,N_12408);
and U12631 (N_12631,N_12482,N_12414);
and U12632 (N_12632,N_12374,N_12429);
nand U12633 (N_12633,N_12478,N_12319);
nand U12634 (N_12634,N_12433,N_12504);
nor U12635 (N_12635,N_12537,N_12490);
xor U12636 (N_12636,N_12403,N_12435);
nand U12637 (N_12637,N_12498,N_12515);
xor U12638 (N_12638,N_12560,N_12481);
nand U12639 (N_12639,N_12301,N_12425);
and U12640 (N_12640,N_12580,N_12556);
nand U12641 (N_12641,N_12501,N_12390);
or U12642 (N_12642,N_12394,N_12525);
nor U12643 (N_12643,N_12360,N_12579);
and U12644 (N_12644,N_12530,N_12575);
or U12645 (N_12645,N_12468,N_12338);
nor U12646 (N_12646,N_12407,N_12308);
nand U12647 (N_12647,N_12540,N_12574);
nand U12648 (N_12648,N_12365,N_12546);
nor U12649 (N_12649,N_12565,N_12438);
or U12650 (N_12650,N_12377,N_12496);
xnor U12651 (N_12651,N_12473,N_12494);
xnor U12652 (N_12652,N_12538,N_12533);
nor U12653 (N_12653,N_12564,N_12470);
and U12654 (N_12654,N_12563,N_12430);
nand U12655 (N_12655,N_12395,N_12375);
or U12656 (N_12656,N_12455,N_12379);
xnor U12657 (N_12657,N_12503,N_12313);
nand U12658 (N_12658,N_12358,N_12590);
nor U12659 (N_12659,N_12306,N_12383);
or U12660 (N_12660,N_12594,N_12559);
xor U12661 (N_12661,N_12572,N_12475);
nor U12662 (N_12662,N_12566,N_12506);
and U12663 (N_12663,N_12348,N_12401);
nand U12664 (N_12664,N_12324,N_12359);
and U12665 (N_12665,N_12568,N_12464);
or U12666 (N_12666,N_12573,N_12542);
xnor U12667 (N_12667,N_12393,N_12380);
nand U12668 (N_12668,N_12320,N_12366);
nand U12669 (N_12669,N_12584,N_12453);
or U12670 (N_12670,N_12526,N_12385);
nand U12671 (N_12671,N_12402,N_12549);
nor U12672 (N_12672,N_12536,N_12491);
or U12673 (N_12673,N_12483,N_12432);
xnor U12674 (N_12674,N_12539,N_12426);
nor U12675 (N_12675,N_12465,N_12371);
and U12676 (N_12676,N_12484,N_12314);
or U12677 (N_12677,N_12353,N_12442);
or U12678 (N_12678,N_12423,N_12399);
nor U12679 (N_12679,N_12384,N_12570);
nor U12680 (N_12680,N_12315,N_12510);
nand U12681 (N_12681,N_12593,N_12418);
nor U12682 (N_12682,N_12553,N_12534);
xnor U12683 (N_12683,N_12304,N_12587);
xnor U12684 (N_12684,N_12441,N_12332);
nor U12685 (N_12685,N_12427,N_12518);
and U12686 (N_12686,N_12477,N_12357);
xor U12687 (N_12687,N_12529,N_12346);
nor U12688 (N_12688,N_12355,N_12488);
and U12689 (N_12689,N_12363,N_12555);
xnor U12690 (N_12690,N_12333,N_12588);
nand U12691 (N_12691,N_12331,N_12487);
or U12692 (N_12692,N_12550,N_12419);
and U12693 (N_12693,N_12581,N_12364);
nor U12694 (N_12694,N_12571,N_12302);
and U12695 (N_12695,N_12528,N_12391);
or U12696 (N_12696,N_12370,N_12524);
or U12697 (N_12697,N_12447,N_12577);
and U12698 (N_12698,N_12493,N_12321);
nor U12699 (N_12699,N_12350,N_12368);
or U12700 (N_12700,N_12596,N_12450);
nand U12701 (N_12701,N_12462,N_12382);
or U12702 (N_12702,N_12509,N_12378);
nor U12703 (N_12703,N_12431,N_12334);
nand U12704 (N_12704,N_12323,N_12597);
and U12705 (N_12705,N_12386,N_12460);
or U12706 (N_12706,N_12373,N_12445);
xor U12707 (N_12707,N_12485,N_12343);
or U12708 (N_12708,N_12342,N_12328);
nand U12709 (N_12709,N_12369,N_12519);
nand U12710 (N_12710,N_12463,N_12511);
nor U12711 (N_12711,N_12479,N_12420);
nor U12712 (N_12712,N_12351,N_12544);
nor U12713 (N_12713,N_12400,N_12557);
and U12714 (N_12714,N_12310,N_12486);
and U12715 (N_12715,N_12410,N_12492);
nor U12716 (N_12716,N_12345,N_12513);
nor U12717 (N_12717,N_12341,N_12335);
and U12718 (N_12718,N_12387,N_12548);
nand U12719 (N_12719,N_12421,N_12340);
or U12720 (N_12720,N_12312,N_12361);
nor U12721 (N_12721,N_12558,N_12576);
xnor U12722 (N_12722,N_12535,N_12422);
nor U12723 (N_12723,N_12339,N_12480);
nand U12724 (N_12724,N_12472,N_12547);
nor U12725 (N_12725,N_12443,N_12424);
and U12726 (N_12726,N_12457,N_12522);
and U12727 (N_12727,N_12476,N_12381);
xor U12728 (N_12728,N_12416,N_12541);
nor U12729 (N_12729,N_12466,N_12454);
nor U12730 (N_12730,N_12411,N_12551);
xor U12731 (N_12731,N_12517,N_12578);
or U12732 (N_12732,N_12591,N_12415);
nor U12733 (N_12733,N_12326,N_12329);
and U12734 (N_12734,N_12507,N_12589);
xnor U12735 (N_12735,N_12317,N_12456);
xor U12736 (N_12736,N_12412,N_12392);
xnor U12737 (N_12737,N_12599,N_12458);
nor U12738 (N_12738,N_12356,N_12406);
and U12739 (N_12739,N_12500,N_12322);
nand U12740 (N_12740,N_12367,N_12452);
nor U12741 (N_12741,N_12325,N_12398);
nor U12742 (N_12742,N_12514,N_12449);
and U12743 (N_12743,N_12372,N_12448);
nor U12744 (N_12744,N_12437,N_12397);
nor U12745 (N_12745,N_12349,N_12404);
nand U12746 (N_12746,N_12396,N_12318);
xor U12747 (N_12747,N_12311,N_12508);
nand U12748 (N_12748,N_12337,N_12592);
and U12749 (N_12749,N_12376,N_12409);
xnor U12750 (N_12750,N_12379,N_12426);
or U12751 (N_12751,N_12526,N_12374);
or U12752 (N_12752,N_12565,N_12566);
nand U12753 (N_12753,N_12507,N_12468);
or U12754 (N_12754,N_12316,N_12496);
nand U12755 (N_12755,N_12477,N_12475);
and U12756 (N_12756,N_12345,N_12529);
xor U12757 (N_12757,N_12593,N_12437);
nor U12758 (N_12758,N_12498,N_12302);
nor U12759 (N_12759,N_12469,N_12480);
nand U12760 (N_12760,N_12546,N_12459);
nor U12761 (N_12761,N_12473,N_12308);
nand U12762 (N_12762,N_12380,N_12542);
or U12763 (N_12763,N_12495,N_12571);
or U12764 (N_12764,N_12594,N_12354);
or U12765 (N_12765,N_12512,N_12486);
and U12766 (N_12766,N_12532,N_12541);
or U12767 (N_12767,N_12386,N_12530);
or U12768 (N_12768,N_12437,N_12478);
or U12769 (N_12769,N_12448,N_12375);
nor U12770 (N_12770,N_12405,N_12314);
or U12771 (N_12771,N_12556,N_12427);
or U12772 (N_12772,N_12374,N_12331);
nand U12773 (N_12773,N_12431,N_12330);
xor U12774 (N_12774,N_12421,N_12318);
nand U12775 (N_12775,N_12438,N_12558);
or U12776 (N_12776,N_12532,N_12319);
nor U12777 (N_12777,N_12319,N_12378);
or U12778 (N_12778,N_12300,N_12591);
nand U12779 (N_12779,N_12533,N_12545);
and U12780 (N_12780,N_12352,N_12444);
xnor U12781 (N_12781,N_12398,N_12402);
xnor U12782 (N_12782,N_12565,N_12413);
xor U12783 (N_12783,N_12553,N_12394);
or U12784 (N_12784,N_12517,N_12336);
nand U12785 (N_12785,N_12336,N_12380);
nand U12786 (N_12786,N_12532,N_12538);
nand U12787 (N_12787,N_12452,N_12364);
xor U12788 (N_12788,N_12335,N_12589);
nand U12789 (N_12789,N_12358,N_12453);
or U12790 (N_12790,N_12403,N_12591);
nor U12791 (N_12791,N_12544,N_12409);
or U12792 (N_12792,N_12551,N_12360);
xnor U12793 (N_12793,N_12411,N_12460);
xor U12794 (N_12794,N_12359,N_12547);
nor U12795 (N_12795,N_12450,N_12470);
nor U12796 (N_12796,N_12400,N_12534);
or U12797 (N_12797,N_12342,N_12505);
xnor U12798 (N_12798,N_12335,N_12313);
xor U12799 (N_12799,N_12310,N_12396);
and U12800 (N_12800,N_12421,N_12417);
or U12801 (N_12801,N_12428,N_12475);
or U12802 (N_12802,N_12568,N_12312);
xor U12803 (N_12803,N_12389,N_12338);
nand U12804 (N_12804,N_12542,N_12429);
nor U12805 (N_12805,N_12530,N_12509);
and U12806 (N_12806,N_12506,N_12520);
and U12807 (N_12807,N_12398,N_12592);
or U12808 (N_12808,N_12511,N_12367);
and U12809 (N_12809,N_12519,N_12439);
and U12810 (N_12810,N_12351,N_12422);
and U12811 (N_12811,N_12562,N_12310);
and U12812 (N_12812,N_12425,N_12307);
nor U12813 (N_12813,N_12542,N_12563);
or U12814 (N_12814,N_12455,N_12445);
or U12815 (N_12815,N_12544,N_12564);
nand U12816 (N_12816,N_12453,N_12589);
or U12817 (N_12817,N_12475,N_12488);
xnor U12818 (N_12818,N_12523,N_12339);
or U12819 (N_12819,N_12518,N_12486);
nand U12820 (N_12820,N_12427,N_12302);
or U12821 (N_12821,N_12496,N_12537);
xnor U12822 (N_12822,N_12566,N_12418);
and U12823 (N_12823,N_12427,N_12376);
xnor U12824 (N_12824,N_12412,N_12521);
xnor U12825 (N_12825,N_12334,N_12419);
xor U12826 (N_12826,N_12470,N_12535);
and U12827 (N_12827,N_12519,N_12535);
nand U12828 (N_12828,N_12595,N_12374);
xor U12829 (N_12829,N_12486,N_12460);
nor U12830 (N_12830,N_12530,N_12355);
nand U12831 (N_12831,N_12471,N_12421);
nand U12832 (N_12832,N_12475,N_12452);
nor U12833 (N_12833,N_12407,N_12439);
nor U12834 (N_12834,N_12543,N_12380);
and U12835 (N_12835,N_12457,N_12404);
and U12836 (N_12836,N_12452,N_12550);
and U12837 (N_12837,N_12371,N_12338);
xor U12838 (N_12838,N_12517,N_12429);
nor U12839 (N_12839,N_12406,N_12434);
or U12840 (N_12840,N_12455,N_12568);
or U12841 (N_12841,N_12410,N_12491);
or U12842 (N_12842,N_12358,N_12435);
xor U12843 (N_12843,N_12474,N_12591);
or U12844 (N_12844,N_12497,N_12422);
xnor U12845 (N_12845,N_12500,N_12453);
nor U12846 (N_12846,N_12424,N_12562);
xnor U12847 (N_12847,N_12583,N_12395);
or U12848 (N_12848,N_12509,N_12320);
and U12849 (N_12849,N_12517,N_12335);
and U12850 (N_12850,N_12462,N_12329);
xor U12851 (N_12851,N_12598,N_12327);
xor U12852 (N_12852,N_12584,N_12532);
and U12853 (N_12853,N_12551,N_12335);
nand U12854 (N_12854,N_12468,N_12543);
xnor U12855 (N_12855,N_12391,N_12460);
nand U12856 (N_12856,N_12326,N_12514);
nand U12857 (N_12857,N_12499,N_12493);
or U12858 (N_12858,N_12589,N_12596);
xnor U12859 (N_12859,N_12379,N_12578);
nor U12860 (N_12860,N_12402,N_12331);
and U12861 (N_12861,N_12410,N_12501);
or U12862 (N_12862,N_12347,N_12578);
nor U12863 (N_12863,N_12473,N_12387);
xor U12864 (N_12864,N_12350,N_12346);
xor U12865 (N_12865,N_12379,N_12555);
xnor U12866 (N_12866,N_12504,N_12334);
nand U12867 (N_12867,N_12449,N_12339);
nand U12868 (N_12868,N_12444,N_12397);
nand U12869 (N_12869,N_12375,N_12548);
nand U12870 (N_12870,N_12382,N_12411);
and U12871 (N_12871,N_12491,N_12522);
xor U12872 (N_12872,N_12468,N_12393);
nor U12873 (N_12873,N_12466,N_12427);
or U12874 (N_12874,N_12582,N_12575);
nor U12875 (N_12875,N_12468,N_12378);
nand U12876 (N_12876,N_12369,N_12401);
nor U12877 (N_12877,N_12533,N_12371);
nor U12878 (N_12878,N_12384,N_12350);
or U12879 (N_12879,N_12490,N_12548);
and U12880 (N_12880,N_12414,N_12445);
nand U12881 (N_12881,N_12461,N_12475);
and U12882 (N_12882,N_12386,N_12566);
or U12883 (N_12883,N_12306,N_12499);
nand U12884 (N_12884,N_12497,N_12407);
or U12885 (N_12885,N_12431,N_12333);
or U12886 (N_12886,N_12392,N_12537);
xor U12887 (N_12887,N_12487,N_12329);
nand U12888 (N_12888,N_12590,N_12438);
or U12889 (N_12889,N_12429,N_12347);
and U12890 (N_12890,N_12356,N_12435);
or U12891 (N_12891,N_12412,N_12546);
xor U12892 (N_12892,N_12518,N_12351);
xor U12893 (N_12893,N_12365,N_12514);
nand U12894 (N_12894,N_12489,N_12522);
and U12895 (N_12895,N_12533,N_12506);
nor U12896 (N_12896,N_12517,N_12379);
nand U12897 (N_12897,N_12578,N_12481);
nor U12898 (N_12898,N_12506,N_12362);
nor U12899 (N_12899,N_12489,N_12531);
and U12900 (N_12900,N_12731,N_12889);
nor U12901 (N_12901,N_12894,N_12839);
or U12902 (N_12902,N_12880,N_12651);
or U12903 (N_12903,N_12716,N_12846);
xor U12904 (N_12904,N_12899,N_12893);
and U12905 (N_12905,N_12744,N_12633);
xnor U12906 (N_12906,N_12660,N_12848);
and U12907 (N_12907,N_12842,N_12810);
and U12908 (N_12908,N_12821,N_12602);
and U12909 (N_12909,N_12876,N_12825);
xnor U12910 (N_12910,N_12708,N_12654);
nand U12911 (N_12911,N_12890,N_12685);
nand U12912 (N_12912,N_12762,N_12702);
nand U12913 (N_12913,N_12745,N_12703);
and U12914 (N_12914,N_12853,N_12618);
nor U12915 (N_12915,N_12729,N_12820);
nor U12916 (N_12916,N_12897,N_12796);
nor U12917 (N_12917,N_12658,N_12807);
and U12918 (N_12918,N_12782,N_12725);
xor U12919 (N_12919,N_12886,N_12608);
nor U12920 (N_12920,N_12833,N_12841);
nand U12921 (N_12921,N_12770,N_12791);
nor U12922 (N_12922,N_12727,N_12746);
and U12923 (N_12923,N_12705,N_12680);
xnor U12924 (N_12924,N_12683,N_12756);
and U12925 (N_12925,N_12775,N_12871);
nand U12926 (N_12926,N_12694,N_12881);
or U12927 (N_12927,N_12664,N_12636);
and U12928 (N_12928,N_12790,N_12778);
and U12929 (N_12929,N_12607,N_12712);
xnor U12930 (N_12930,N_12895,N_12795);
xnor U12931 (N_12931,N_12620,N_12836);
nand U12932 (N_12932,N_12748,N_12780);
nor U12933 (N_12933,N_12860,N_12670);
xnor U12934 (N_12934,N_12774,N_12643);
xnor U12935 (N_12935,N_12630,N_12676);
xor U12936 (N_12936,N_12641,N_12757);
and U12937 (N_12937,N_12678,N_12681);
xor U12938 (N_12938,N_12711,N_12755);
or U12939 (N_12939,N_12814,N_12624);
or U12940 (N_12940,N_12690,N_12609);
or U12941 (N_12941,N_12870,N_12747);
xnor U12942 (N_12942,N_12743,N_12826);
or U12943 (N_12943,N_12614,N_12687);
or U12944 (N_12944,N_12830,N_12793);
and U12945 (N_12945,N_12832,N_12800);
or U12946 (N_12946,N_12753,N_12714);
and U12947 (N_12947,N_12763,N_12816);
xor U12948 (N_12948,N_12722,N_12700);
and U12949 (N_12949,N_12691,N_12809);
or U12950 (N_12950,N_12766,N_12686);
nand U12951 (N_12951,N_12724,N_12612);
and U12952 (N_12952,N_12741,N_12805);
and U12953 (N_12953,N_12781,N_12802);
nand U12954 (N_12954,N_12704,N_12783);
nor U12955 (N_12955,N_12627,N_12642);
and U12956 (N_12956,N_12626,N_12616);
and U12957 (N_12957,N_12752,N_12863);
nor U12958 (N_12958,N_12754,N_12721);
nand U12959 (N_12959,N_12697,N_12872);
xnor U12960 (N_12960,N_12813,N_12845);
nor U12961 (N_12961,N_12885,N_12827);
and U12962 (N_12962,N_12789,N_12615);
nor U12963 (N_12963,N_12888,N_12735);
and U12964 (N_12964,N_12673,N_12662);
nor U12965 (N_12965,N_12606,N_12750);
nor U12966 (N_12966,N_12765,N_12652);
and U12967 (N_12967,N_12764,N_12709);
nand U12968 (N_12968,N_12878,N_12794);
and U12969 (N_12969,N_12603,N_12856);
and U12970 (N_12970,N_12879,N_12773);
nand U12971 (N_12971,N_12682,N_12849);
or U12972 (N_12972,N_12734,N_12733);
nand U12973 (N_12973,N_12883,N_12669);
or U12974 (N_12974,N_12726,N_12874);
or U12975 (N_12975,N_12877,N_12867);
and U12976 (N_12976,N_12869,N_12674);
and U12977 (N_12977,N_12737,N_12657);
nand U12978 (N_12978,N_12646,N_12644);
and U12979 (N_12979,N_12696,N_12840);
or U12980 (N_12980,N_12760,N_12811);
nand U12981 (N_12981,N_12875,N_12613);
and U12982 (N_12982,N_12666,N_12837);
and U12983 (N_12983,N_12767,N_12859);
nor U12984 (N_12984,N_12655,N_12661);
xnor U12985 (N_12985,N_12749,N_12710);
or U12986 (N_12986,N_12647,N_12858);
or U12987 (N_12987,N_12777,N_12617);
or U12988 (N_12988,N_12808,N_12601);
nor U12989 (N_12989,N_12785,N_12882);
xnor U12990 (N_12990,N_12713,N_12701);
and U12991 (N_12991,N_12834,N_12852);
nand U12992 (N_12992,N_12815,N_12865);
or U12993 (N_12993,N_12695,N_12640);
or U12994 (N_12994,N_12844,N_12868);
xor U12995 (N_12995,N_12862,N_12706);
and U12996 (N_12996,N_12797,N_12632);
nand U12997 (N_12997,N_12738,N_12637);
xor U12998 (N_12998,N_12648,N_12671);
xor U12999 (N_12999,N_12887,N_12838);
and U13000 (N_13000,N_12740,N_12635);
nor U13001 (N_13001,N_12653,N_12828);
nand U13002 (N_13002,N_12759,N_12779);
nor U13003 (N_13003,N_12792,N_12786);
nand U13004 (N_13004,N_12776,N_12822);
xnor U13005 (N_13005,N_12667,N_12684);
nand U13006 (N_13006,N_12668,N_12719);
nand U13007 (N_13007,N_12698,N_12730);
xor U13008 (N_13008,N_12656,N_12751);
xor U13009 (N_13009,N_12772,N_12817);
nand U13010 (N_13010,N_12803,N_12768);
nand U13011 (N_13011,N_12679,N_12634);
xor U13012 (N_13012,N_12761,N_12718);
xnor U13013 (N_13013,N_12693,N_12677);
or U13014 (N_13014,N_12861,N_12625);
or U13015 (N_13015,N_12638,N_12788);
xnor U13016 (N_13016,N_12600,N_12843);
xor U13017 (N_13017,N_12896,N_12663);
and U13018 (N_13018,N_12784,N_12739);
nand U13019 (N_13019,N_12728,N_12892);
nand U13020 (N_13020,N_12801,N_12631);
and U13021 (N_13021,N_12645,N_12621);
xnor U13022 (N_13022,N_12699,N_12804);
nand U13023 (N_13023,N_12864,N_12847);
nor U13024 (N_13024,N_12835,N_12799);
nand U13025 (N_13025,N_12732,N_12604);
xor U13026 (N_13026,N_12758,N_12605);
nor U13027 (N_13027,N_12665,N_12742);
nor U13028 (N_13028,N_12692,N_12619);
or U13029 (N_13029,N_12857,N_12689);
and U13030 (N_13030,N_12806,N_12854);
xnor U13031 (N_13031,N_12650,N_12622);
or U13032 (N_13032,N_12823,N_12850);
and U13033 (N_13033,N_12629,N_12723);
xnor U13034 (N_13034,N_12672,N_12898);
or U13035 (N_13035,N_12715,N_12798);
and U13036 (N_13036,N_12623,N_12884);
nand U13037 (N_13037,N_12831,N_12688);
nand U13038 (N_13038,N_12771,N_12717);
xnor U13039 (N_13039,N_12891,N_12628);
and U13040 (N_13040,N_12787,N_12812);
and U13041 (N_13041,N_12873,N_12736);
or U13042 (N_13042,N_12851,N_12818);
xnor U13043 (N_13043,N_12819,N_12611);
nor U13044 (N_13044,N_12649,N_12639);
or U13045 (N_13045,N_12659,N_12866);
nor U13046 (N_13046,N_12855,N_12720);
and U13047 (N_13047,N_12610,N_12829);
or U13048 (N_13048,N_12675,N_12824);
xor U13049 (N_13049,N_12707,N_12769);
xor U13050 (N_13050,N_12750,N_12796);
xor U13051 (N_13051,N_12686,N_12735);
xor U13052 (N_13052,N_12688,N_12675);
and U13053 (N_13053,N_12677,N_12894);
or U13054 (N_13054,N_12682,N_12737);
and U13055 (N_13055,N_12612,N_12814);
nor U13056 (N_13056,N_12843,N_12886);
and U13057 (N_13057,N_12663,N_12854);
and U13058 (N_13058,N_12697,N_12603);
and U13059 (N_13059,N_12819,N_12647);
and U13060 (N_13060,N_12866,N_12806);
xor U13061 (N_13061,N_12700,N_12867);
and U13062 (N_13062,N_12842,N_12632);
and U13063 (N_13063,N_12610,N_12807);
and U13064 (N_13064,N_12814,N_12781);
and U13065 (N_13065,N_12852,N_12841);
and U13066 (N_13066,N_12756,N_12834);
nand U13067 (N_13067,N_12611,N_12623);
xnor U13068 (N_13068,N_12891,N_12893);
nand U13069 (N_13069,N_12882,N_12786);
nand U13070 (N_13070,N_12694,N_12684);
nand U13071 (N_13071,N_12613,N_12695);
or U13072 (N_13072,N_12681,N_12814);
or U13073 (N_13073,N_12727,N_12626);
or U13074 (N_13074,N_12834,N_12605);
or U13075 (N_13075,N_12673,N_12656);
nand U13076 (N_13076,N_12655,N_12754);
and U13077 (N_13077,N_12740,N_12823);
nor U13078 (N_13078,N_12873,N_12746);
xnor U13079 (N_13079,N_12861,N_12661);
nor U13080 (N_13080,N_12649,N_12817);
xnor U13081 (N_13081,N_12854,N_12802);
or U13082 (N_13082,N_12663,N_12807);
xnor U13083 (N_13083,N_12875,N_12714);
xnor U13084 (N_13084,N_12826,N_12797);
xor U13085 (N_13085,N_12610,N_12895);
and U13086 (N_13086,N_12889,N_12704);
and U13087 (N_13087,N_12790,N_12870);
and U13088 (N_13088,N_12636,N_12628);
and U13089 (N_13089,N_12825,N_12892);
nand U13090 (N_13090,N_12616,N_12673);
nand U13091 (N_13091,N_12826,N_12805);
and U13092 (N_13092,N_12802,N_12773);
and U13093 (N_13093,N_12659,N_12785);
xnor U13094 (N_13094,N_12723,N_12830);
nor U13095 (N_13095,N_12814,N_12769);
xor U13096 (N_13096,N_12603,N_12829);
xor U13097 (N_13097,N_12857,N_12802);
xnor U13098 (N_13098,N_12777,N_12673);
xnor U13099 (N_13099,N_12721,N_12795);
and U13100 (N_13100,N_12727,N_12813);
xor U13101 (N_13101,N_12774,N_12857);
and U13102 (N_13102,N_12778,N_12890);
and U13103 (N_13103,N_12640,N_12718);
nand U13104 (N_13104,N_12684,N_12607);
nand U13105 (N_13105,N_12692,N_12655);
nor U13106 (N_13106,N_12751,N_12815);
nand U13107 (N_13107,N_12847,N_12823);
and U13108 (N_13108,N_12746,N_12766);
and U13109 (N_13109,N_12642,N_12628);
or U13110 (N_13110,N_12623,N_12829);
nand U13111 (N_13111,N_12854,N_12863);
xor U13112 (N_13112,N_12643,N_12800);
xnor U13113 (N_13113,N_12692,N_12751);
xor U13114 (N_13114,N_12767,N_12696);
and U13115 (N_13115,N_12708,N_12767);
and U13116 (N_13116,N_12756,N_12625);
xor U13117 (N_13117,N_12692,N_12738);
or U13118 (N_13118,N_12665,N_12802);
xnor U13119 (N_13119,N_12799,N_12607);
nor U13120 (N_13120,N_12669,N_12680);
or U13121 (N_13121,N_12713,N_12862);
xor U13122 (N_13122,N_12850,N_12838);
nand U13123 (N_13123,N_12720,N_12741);
xnor U13124 (N_13124,N_12763,N_12732);
or U13125 (N_13125,N_12878,N_12716);
nand U13126 (N_13126,N_12837,N_12802);
xnor U13127 (N_13127,N_12609,N_12732);
or U13128 (N_13128,N_12827,N_12853);
and U13129 (N_13129,N_12697,N_12667);
or U13130 (N_13130,N_12814,N_12875);
or U13131 (N_13131,N_12758,N_12834);
or U13132 (N_13132,N_12629,N_12608);
and U13133 (N_13133,N_12831,N_12630);
or U13134 (N_13134,N_12675,N_12619);
nor U13135 (N_13135,N_12712,N_12747);
and U13136 (N_13136,N_12756,N_12870);
or U13137 (N_13137,N_12745,N_12684);
and U13138 (N_13138,N_12815,N_12693);
xnor U13139 (N_13139,N_12744,N_12812);
nand U13140 (N_13140,N_12738,N_12850);
xor U13141 (N_13141,N_12834,N_12840);
or U13142 (N_13142,N_12745,N_12761);
xor U13143 (N_13143,N_12656,N_12879);
or U13144 (N_13144,N_12832,N_12728);
nand U13145 (N_13145,N_12839,N_12814);
or U13146 (N_13146,N_12898,N_12642);
nand U13147 (N_13147,N_12884,N_12791);
or U13148 (N_13148,N_12621,N_12616);
nor U13149 (N_13149,N_12635,N_12660);
and U13150 (N_13150,N_12710,N_12646);
nor U13151 (N_13151,N_12862,N_12728);
or U13152 (N_13152,N_12677,N_12647);
nand U13153 (N_13153,N_12658,N_12649);
nand U13154 (N_13154,N_12869,N_12835);
nor U13155 (N_13155,N_12662,N_12625);
xor U13156 (N_13156,N_12732,N_12620);
nor U13157 (N_13157,N_12648,N_12870);
and U13158 (N_13158,N_12889,N_12621);
and U13159 (N_13159,N_12670,N_12703);
or U13160 (N_13160,N_12881,N_12601);
and U13161 (N_13161,N_12603,N_12717);
or U13162 (N_13162,N_12878,N_12686);
nand U13163 (N_13163,N_12837,N_12734);
and U13164 (N_13164,N_12737,N_12738);
or U13165 (N_13165,N_12672,N_12741);
nand U13166 (N_13166,N_12700,N_12803);
nand U13167 (N_13167,N_12674,N_12696);
nor U13168 (N_13168,N_12623,N_12657);
nor U13169 (N_13169,N_12663,N_12676);
nor U13170 (N_13170,N_12813,N_12649);
nand U13171 (N_13171,N_12764,N_12887);
nand U13172 (N_13172,N_12778,N_12613);
nand U13173 (N_13173,N_12666,N_12815);
nand U13174 (N_13174,N_12760,N_12665);
or U13175 (N_13175,N_12802,N_12704);
xor U13176 (N_13176,N_12812,N_12807);
xnor U13177 (N_13177,N_12896,N_12810);
nor U13178 (N_13178,N_12752,N_12640);
and U13179 (N_13179,N_12865,N_12668);
or U13180 (N_13180,N_12814,N_12844);
and U13181 (N_13181,N_12899,N_12696);
and U13182 (N_13182,N_12848,N_12631);
nand U13183 (N_13183,N_12770,N_12711);
nor U13184 (N_13184,N_12608,N_12697);
nor U13185 (N_13185,N_12658,N_12868);
and U13186 (N_13186,N_12678,N_12746);
nor U13187 (N_13187,N_12607,N_12694);
or U13188 (N_13188,N_12867,N_12717);
and U13189 (N_13189,N_12679,N_12892);
or U13190 (N_13190,N_12710,N_12686);
xnor U13191 (N_13191,N_12626,N_12889);
and U13192 (N_13192,N_12873,N_12790);
xor U13193 (N_13193,N_12779,N_12709);
nand U13194 (N_13194,N_12717,N_12724);
xnor U13195 (N_13195,N_12790,N_12863);
nand U13196 (N_13196,N_12847,N_12895);
xnor U13197 (N_13197,N_12625,N_12774);
xor U13198 (N_13198,N_12755,N_12692);
nor U13199 (N_13199,N_12646,N_12747);
or U13200 (N_13200,N_13192,N_13108);
nor U13201 (N_13201,N_12966,N_12951);
nor U13202 (N_13202,N_12971,N_12939);
or U13203 (N_13203,N_12961,N_13132);
and U13204 (N_13204,N_13109,N_13170);
or U13205 (N_13205,N_12912,N_13185);
or U13206 (N_13206,N_12922,N_13139);
and U13207 (N_13207,N_13035,N_12934);
and U13208 (N_13208,N_13018,N_12932);
nor U13209 (N_13209,N_13147,N_13045);
or U13210 (N_13210,N_12938,N_12928);
and U13211 (N_13211,N_13182,N_13187);
and U13212 (N_13212,N_13178,N_12944);
nor U13213 (N_13213,N_13001,N_13127);
and U13214 (N_13214,N_13005,N_12940);
or U13215 (N_13215,N_12995,N_12930);
or U13216 (N_13216,N_13110,N_13145);
xor U13217 (N_13217,N_13113,N_13078);
nor U13218 (N_13218,N_13138,N_13085);
nor U13219 (N_13219,N_13051,N_13006);
and U13220 (N_13220,N_13003,N_13080);
nand U13221 (N_13221,N_12926,N_12972);
xnor U13222 (N_13222,N_13097,N_12987);
or U13223 (N_13223,N_12913,N_12937);
and U13224 (N_13224,N_12978,N_13054);
xor U13225 (N_13225,N_13135,N_12973);
nor U13226 (N_13226,N_13030,N_13086);
nor U13227 (N_13227,N_12908,N_13022);
nor U13228 (N_13228,N_12969,N_13048);
or U13229 (N_13229,N_13026,N_13155);
and U13230 (N_13230,N_13042,N_12960);
xor U13231 (N_13231,N_13146,N_13183);
or U13232 (N_13232,N_12915,N_13133);
and U13233 (N_13233,N_13096,N_12919);
nand U13234 (N_13234,N_13197,N_13164);
nor U13235 (N_13235,N_13055,N_12963);
and U13236 (N_13236,N_12991,N_13065);
nand U13237 (N_13237,N_12947,N_13144);
nand U13238 (N_13238,N_13101,N_12959);
or U13239 (N_13239,N_12952,N_13128);
nand U13240 (N_13240,N_13075,N_12999);
and U13241 (N_13241,N_13041,N_13036);
xor U13242 (N_13242,N_12925,N_13102);
xnor U13243 (N_13243,N_12992,N_13159);
nor U13244 (N_13244,N_12994,N_12968);
xnor U13245 (N_13245,N_13010,N_13149);
xor U13246 (N_13246,N_13126,N_13088);
nor U13247 (N_13247,N_12933,N_13034);
xor U13248 (N_13248,N_13057,N_13194);
xnor U13249 (N_13249,N_13180,N_13062);
or U13250 (N_13250,N_13148,N_13087);
or U13251 (N_13251,N_12984,N_13115);
xnor U13252 (N_13252,N_13019,N_13043);
nand U13253 (N_13253,N_12923,N_12945);
and U13254 (N_13254,N_12900,N_12980);
xnor U13255 (N_13255,N_13025,N_13052);
nand U13256 (N_13256,N_12976,N_12970);
nor U13257 (N_13257,N_12954,N_13039);
xor U13258 (N_13258,N_13123,N_13082);
nor U13259 (N_13259,N_12998,N_13174);
and U13260 (N_13260,N_13131,N_13195);
nor U13261 (N_13261,N_13070,N_12982);
and U13262 (N_13262,N_13084,N_13099);
and U13263 (N_13263,N_12941,N_13157);
nand U13264 (N_13264,N_13176,N_12907);
or U13265 (N_13265,N_12985,N_13112);
and U13266 (N_13266,N_13095,N_13152);
nor U13267 (N_13267,N_13141,N_13023);
xor U13268 (N_13268,N_12901,N_13119);
xor U13269 (N_13269,N_13044,N_13040);
xnor U13270 (N_13270,N_13033,N_12942);
nand U13271 (N_13271,N_12974,N_13014);
nor U13272 (N_13272,N_13004,N_13104);
nand U13273 (N_13273,N_12921,N_12986);
or U13274 (N_13274,N_13177,N_12975);
or U13275 (N_13275,N_13032,N_12967);
xor U13276 (N_13276,N_13071,N_12993);
xnor U13277 (N_13277,N_13013,N_13168);
nand U13278 (N_13278,N_13047,N_13037);
nand U13279 (N_13279,N_13150,N_13163);
nand U13280 (N_13280,N_12958,N_13002);
xor U13281 (N_13281,N_13098,N_12957);
and U13282 (N_13282,N_13077,N_13162);
xor U13283 (N_13283,N_12953,N_12979);
nand U13284 (N_13284,N_13175,N_13016);
nand U13285 (N_13285,N_12943,N_13143);
or U13286 (N_13286,N_13118,N_13009);
and U13287 (N_13287,N_12955,N_12918);
xnor U13288 (N_13288,N_13094,N_13083);
nor U13289 (N_13289,N_13000,N_13167);
nor U13290 (N_13290,N_13153,N_13198);
nor U13291 (N_13291,N_12910,N_13103);
nor U13292 (N_13292,N_13160,N_13166);
nand U13293 (N_13293,N_13184,N_13130);
xnor U13294 (N_13294,N_13079,N_13122);
xnor U13295 (N_13295,N_13116,N_13008);
and U13296 (N_13296,N_13011,N_13121);
nand U13297 (N_13297,N_13069,N_13129);
xnor U13298 (N_13298,N_12988,N_13063);
nand U13299 (N_13299,N_13134,N_13193);
nor U13300 (N_13300,N_13181,N_12929);
nor U13301 (N_13301,N_13024,N_13188);
nor U13302 (N_13302,N_12965,N_12946);
xor U13303 (N_13303,N_13124,N_13093);
nor U13304 (N_13304,N_12911,N_13031);
or U13305 (N_13305,N_13161,N_12902);
and U13306 (N_13306,N_13067,N_13007);
or U13307 (N_13307,N_13050,N_13154);
and U13308 (N_13308,N_13064,N_13117);
xor U13309 (N_13309,N_13046,N_13172);
and U13310 (N_13310,N_13074,N_13199);
nand U13311 (N_13311,N_13106,N_13171);
xnor U13312 (N_13312,N_13073,N_12920);
and U13313 (N_13313,N_13137,N_12977);
nor U13314 (N_13314,N_12904,N_12924);
or U13315 (N_13315,N_12909,N_12950);
xnor U13316 (N_13316,N_13012,N_13100);
xor U13317 (N_13317,N_13089,N_12997);
nor U13318 (N_13318,N_13058,N_13060);
nor U13319 (N_13319,N_13158,N_13068);
nand U13320 (N_13320,N_12949,N_13061);
nand U13321 (N_13321,N_12990,N_12927);
nor U13322 (N_13322,N_13169,N_13020);
nor U13323 (N_13323,N_12906,N_13156);
nand U13324 (N_13324,N_13029,N_13092);
xnor U13325 (N_13325,N_13021,N_13081);
or U13326 (N_13326,N_12905,N_13017);
and U13327 (N_13327,N_13028,N_13105);
and U13328 (N_13328,N_12903,N_13165);
nor U13329 (N_13329,N_13189,N_12964);
nand U13330 (N_13330,N_12981,N_13114);
xnor U13331 (N_13331,N_12916,N_12931);
or U13332 (N_13332,N_12962,N_13140);
nand U13333 (N_13333,N_13059,N_13056);
and U13334 (N_13334,N_13120,N_13038);
xor U13335 (N_13335,N_12935,N_12917);
or U13336 (N_13336,N_12936,N_12948);
nand U13337 (N_13337,N_13190,N_13015);
or U13338 (N_13338,N_12983,N_13125);
nor U13339 (N_13339,N_13066,N_13142);
xor U13340 (N_13340,N_12989,N_13027);
nand U13341 (N_13341,N_12996,N_13091);
nand U13342 (N_13342,N_12956,N_13191);
nor U13343 (N_13343,N_13151,N_13136);
nor U13344 (N_13344,N_13053,N_13072);
or U13345 (N_13345,N_13173,N_13076);
and U13346 (N_13346,N_13186,N_13179);
nand U13347 (N_13347,N_12914,N_13049);
nand U13348 (N_13348,N_13107,N_13111);
nand U13349 (N_13349,N_13090,N_13196);
nand U13350 (N_13350,N_12970,N_13141);
or U13351 (N_13351,N_12943,N_13177);
or U13352 (N_13352,N_12925,N_13096);
xnor U13353 (N_13353,N_13087,N_13167);
nand U13354 (N_13354,N_13126,N_13106);
xor U13355 (N_13355,N_13150,N_13175);
or U13356 (N_13356,N_13198,N_13000);
and U13357 (N_13357,N_13026,N_13129);
nor U13358 (N_13358,N_12991,N_13072);
or U13359 (N_13359,N_13081,N_13173);
xor U13360 (N_13360,N_12924,N_13136);
xnor U13361 (N_13361,N_13083,N_12966);
nand U13362 (N_13362,N_12903,N_12978);
nand U13363 (N_13363,N_13061,N_12951);
nand U13364 (N_13364,N_12920,N_12933);
xnor U13365 (N_13365,N_13128,N_12972);
nand U13366 (N_13366,N_13137,N_13074);
nor U13367 (N_13367,N_13049,N_13078);
or U13368 (N_13368,N_12929,N_13069);
nand U13369 (N_13369,N_12980,N_13128);
and U13370 (N_13370,N_13156,N_12950);
nand U13371 (N_13371,N_12949,N_12981);
xnor U13372 (N_13372,N_13102,N_13119);
nor U13373 (N_13373,N_13153,N_13000);
nor U13374 (N_13374,N_12944,N_13098);
or U13375 (N_13375,N_13137,N_12914);
nor U13376 (N_13376,N_12985,N_12947);
nor U13377 (N_13377,N_13035,N_12930);
nor U13378 (N_13378,N_12959,N_13164);
xor U13379 (N_13379,N_13120,N_12964);
or U13380 (N_13380,N_13107,N_12951);
or U13381 (N_13381,N_12981,N_12950);
or U13382 (N_13382,N_13090,N_13032);
nand U13383 (N_13383,N_12961,N_13013);
nor U13384 (N_13384,N_13128,N_12943);
xnor U13385 (N_13385,N_13083,N_13171);
nor U13386 (N_13386,N_12969,N_13086);
and U13387 (N_13387,N_13128,N_13030);
or U13388 (N_13388,N_12950,N_13073);
nand U13389 (N_13389,N_13076,N_13058);
nor U13390 (N_13390,N_12900,N_13119);
nand U13391 (N_13391,N_13098,N_12965);
nand U13392 (N_13392,N_13007,N_13114);
or U13393 (N_13393,N_13129,N_13019);
nor U13394 (N_13394,N_13121,N_13033);
or U13395 (N_13395,N_12914,N_13004);
nor U13396 (N_13396,N_12984,N_12914);
and U13397 (N_13397,N_13097,N_13142);
xor U13398 (N_13398,N_13136,N_13130);
nand U13399 (N_13399,N_12933,N_13161);
xor U13400 (N_13400,N_13064,N_13148);
or U13401 (N_13401,N_13046,N_13089);
and U13402 (N_13402,N_12957,N_13110);
nor U13403 (N_13403,N_12975,N_13152);
nand U13404 (N_13404,N_13169,N_13151);
nand U13405 (N_13405,N_13166,N_13172);
xor U13406 (N_13406,N_12916,N_13195);
nor U13407 (N_13407,N_13104,N_12926);
and U13408 (N_13408,N_12905,N_13197);
nor U13409 (N_13409,N_13189,N_13198);
xor U13410 (N_13410,N_13150,N_13056);
or U13411 (N_13411,N_12954,N_13104);
nand U13412 (N_13412,N_13135,N_12923);
and U13413 (N_13413,N_12970,N_13087);
or U13414 (N_13414,N_12909,N_13035);
or U13415 (N_13415,N_13014,N_13069);
and U13416 (N_13416,N_13023,N_12970);
nor U13417 (N_13417,N_13017,N_12907);
and U13418 (N_13418,N_12965,N_12978);
or U13419 (N_13419,N_12968,N_13078);
or U13420 (N_13420,N_13017,N_13033);
nor U13421 (N_13421,N_13004,N_13131);
xnor U13422 (N_13422,N_13180,N_13006);
xor U13423 (N_13423,N_13169,N_12990);
xnor U13424 (N_13424,N_13080,N_13082);
nand U13425 (N_13425,N_13118,N_13129);
and U13426 (N_13426,N_13168,N_13080);
or U13427 (N_13427,N_13145,N_12904);
and U13428 (N_13428,N_13162,N_13144);
or U13429 (N_13429,N_12984,N_12940);
or U13430 (N_13430,N_13005,N_12955);
and U13431 (N_13431,N_13015,N_13008);
xnor U13432 (N_13432,N_13111,N_13004);
or U13433 (N_13433,N_13096,N_12963);
and U13434 (N_13434,N_12901,N_13152);
xor U13435 (N_13435,N_13151,N_13077);
or U13436 (N_13436,N_13171,N_13005);
or U13437 (N_13437,N_12969,N_13025);
and U13438 (N_13438,N_13104,N_12970);
xor U13439 (N_13439,N_13052,N_13027);
nor U13440 (N_13440,N_13161,N_13151);
nor U13441 (N_13441,N_13006,N_13000);
nor U13442 (N_13442,N_13179,N_12946);
xnor U13443 (N_13443,N_12961,N_12979);
and U13444 (N_13444,N_13066,N_13064);
nand U13445 (N_13445,N_12986,N_12916);
nor U13446 (N_13446,N_13163,N_13148);
nor U13447 (N_13447,N_13149,N_13016);
xor U13448 (N_13448,N_13116,N_13045);
nor U13449 (N_13449,N_13010,N_13075);
and U13450 (N_13450,N_12947,N_12995);
xor U13451 (N_13451,N_13052,N_12930);
or U13452 (N_13452,N_13083,N_13129);
nor U13453 (N_13453,N_13176,N_13000);
nor U13454 (N_13454,N_12945,N_13011);
nand U13455 (N_13455,N_13166,N_13178);
xnor U13456 (N_13456,N_13008,N_13194);
and U13457 (N_13457,N_12926,N_13055);
nand U13458 (N_13458,N_12916,N_13062);
or U13459 (N_13459,N_13068,N_12977);
nor U13460 (N_13460,N_12941,N_13168);
xnor U13461 (N_13461,N_13109,N_13062);
xor U13462 (N_13462,N_13066,N_12994);
nor U13463 (N_13463,N_12910,N_12981);
nand U13464 (N_13464,N_13040,N_13182);
nand U13465 (N_13465,N_13087,N_13059);
and U13466 (N_13466,N_12937,N_13120);
or U13467 (N_13467,N_13014,N_13065);
nand U13468 (N_13468,N_13188,N_13068);
or U13469 (N_13469,N_12916,N_13086);
nor U13470 (N_13470,N_13181,N_13089);
xnor U13471 (N_13471,N_13098,N_13095);
nor U13472 (N_13472,N_13008,N_13121);
or U13473 (N_13473,N_13063,N_13166);
and U13474 (N_13474,N_13164,N_13096);
or U13475 (N_13475,N_13149,N_13029);
xor U13476 (N_13476,N_12927,N_12969);
nand U13477 (N_13477,N_13079,N_13080);
nor U13478 (N_13478,N_12966,N_13116);
xor U13479 (N_13479,N_12940,N_12914);
xor U13480 (N_13480,N_13120,N_13196);
and U13481 (N_13481,N_13100,N_13114);
nor U13482 (N_13482,N_13043,N_13129);
nor U13483 (N_13483,N_13166,N_13084);
nand U13484 (N_13484,N_13196,N_12927);
nand U13485 (N_13485,N_13172,N_13128);
xor U13486 (N_13486,N_13149,N_12950);
nor U13487 (N_13487,N_13096,N_13138);
and U13488 (N_13488,N_12975,N_13099);
nand U13489 (N_13489,N_12957,N_13031);
or U13490 (N_13490,N_12927,N_13111);
or U13491 (N_13491,N_13172,N_13182);
or U13492 (N_13492,N_12970,N_13150);
nand U13493 (N_13493,N_13195,N_13020);
nor U13494 (N_13494,N_12922,N_12946);
and U13495 (N_13495,N_12976,N_13066);
nand U13496 (N_13496,N_13167,N_13010);
xor U13497 (N_13497,N_13087,N_12927);
or U13498 (N_13498,N_13152,N_12942);
or U13499 (N_13499,N_13048,N_13068);
nor U13500 (N_13500,N_13456,N_13295);
or U13501 (N_13501,N_13241,N_13270);
nor U13502 (N_13502,N_13232,N_13411);
and U13503 (N_13503,N_13415,N_13401);
and U13504 (N_13504,N_13345,N_13200);
and U13505 (N_13505,N_13271,N_13266);
nand U13506 (N_13506,N_13252,N_13227);
nor U13507 (N_13507,N_13349,N_13260);
nor U13508 (N_13508,N_13378,N_13278);
xor U13509 (N_13509,N_13438,N_13485);
xor U13510 (N_13510,N_13394,N_13254);
nand U13511 (N_13511,N_13347,N_13296);
nand U13512 (N_13512,N_13341,N_13372);
or U13513 (N_13513,N_13444,N_13390);
nor U13514 (N_13514,N_13304,N_13328);
or U13515 (N_13515,N_13329,N_13308);
and U13516 (N_13516,N_13332,N_13422);
xnor U13517 (N_13517,N_13206,N_13223);
nor U13518 (N_13518,N_13342,N_13319);
nor U13519 (N_13519,N_13373,N_13307);
and U13520 (N_13520,N_13396,N_13454);
and U13521 (N_13521,N_13478,N_13230);
xor U13522 (N_13522,N_13370,N_13262);
nand U13523 (N_13523,N_13386,N_13312);
nand U13524 (N_13524,N_13413,N_13311);
nand U13525 (N_13525,N_13487,N_13355);
nor U13526 (N_13526,N_13204,N_13461);
or U13527 (N_13527,N_13363,N_13369);
and U13528 (N_13528,N_13491,N_13466);
nor U13529 (N_13529,N_13470,N_13377);
xnor U13530 (N_13530,N_13228,N_13361);
nor U13531 (N_13531,N_13408,N_13250);
nor U13532 (N_13532,N_13337,N_13299);
or U13533 (N_13533,N_13393,N_13240);
and U13534 (N_13534,N_13334,N_13344);
xnor U13535 (N_13535,N_13272,N_13264);
or U13536 (N_13536,N_13467,N_13367);
or U13537 (N_13537,N_13353,N_13446);
or U13538 (N_13538,N_13453,N_13496);
nor U13539 (N_13539,N_13388,N_13483);
or U13540 (N_13540,N_13371,N_13430);
and U13541 (N_13541,N_13225,N_13404);
and U13542 (N_13542,N_13350,N_13448);
xor U13543 (N_13543,N_13450,N_13383);
or U13544 (N_13544,N_13352,N_13479);
nand U13545 (N_13545,N_13406,N_13455);
xor U13546 (N_13546,N_13423,N_13283);
or U13547 (N_13547,N_13417,N_13435);
and U13548 (N_13548,N_13398,N_13309);
nor U13549 (N_13549,N_13480,N_13219);
nand U13550 (N_13550,N_13243,N_13460);
and U13551 (N_13551,N_13387,N_13267);
nor U13552 (N_13552,N_13364,N_13339);
nor U13553 (N_13553,N_13273,N_13358);
nor U13554 (N_13554,N_13284,N_13469);
and U13555 (N_13555,N_13489,N_13488);
nand U13556 (N_13556,N_13294,N_13326);
xor U13557 (N_13557,N_13217,N_13379);
or U13558 (N_13558,N_13324,N_13293);
xor U13559 (N_13559,N_13213,N_13297);
or U13560 (N_13560,N_13202,N_13285);
nor U13561 (N_13561,N_13322,N_13244);
nand U13562 (N_13562,N_13351,N_13286);
and U13563 (N_13563,N_13248,N_13259);
nor U13564 (N_13564,N_13323,N_13320);
nand U13565 (N_13565,N_13424,N_13463);
nand U13566 (N_13566,N_13410,N_13229);
and U13567 (N_13567,N_13333,N_13389);
or U13568 (N_13568,N_13392,N_13427);
nand U13569 (N_13569,N_13476,N_13359);
and U13570 (N_13570,N_13360,N_13346);
xor U13571 (N_13571,N_13269,N_13291);
xnor U13572 (N_13572,N_13428,N_13258);
nor U13573 (N_13573,N_13221,N_13256);
and U13574 (N_13574,N_13318,N_13251);
xor U13575 (N_13575,N_13471,N_13374);
nand U13576 (N_13576,N_13263,N_13368);
nand U13577 (N_13577,N_13305,N_13432);
or U13578 (N_13578,N_13224,N_13357);
or U13579 (N_13579,N_13317,N_13474);
or U13580 (N_13580,N_13282,N_13439);
and U13581 (N_13581,N_13464,N_13209);
nand U13582 (N_13582,N_13433,N_13306);
or U13583 (N_13583,N_13201,N_13313);
nand U13584 (N_13584,N_13459,N_13481);
nor U13585 (N_13585,N_13492,N_13403);
xor U13586 (N_13586,N_13289,N_13255);
nand U13587 (N_13587,N_13298,N_13247);
or U13588 (N_13588,N_13445,N_13416);
nand U13589 (N_13589,N_13443,N_13231);
or U13590 (N_13590,N_13420,N_13376);
or U13591 (N_13591,N_13409,N_13331);
or U13592 (N_13592,N_13465,N_13315);
or U13593 (N_13593,N_13486,N_13280);
or U13594 (N_13594,N_13497,N_13253);
and U13595 (N_13595,N_13407,N_13380);
and U13596 (N_13596,N_13418,N_13375);
nor U13597 (N_13597,N_13400,N_13238);
nor U13598 (N_13598,N_13425,N_13402);
nand U13599 (N_13599,N_13397,N_13327);
or U13600 (N_13600,N_13288,N_13475);
and U13601 (N_13601,N_13381,N_13462);
or U13602 (N_13602,N_13279,N_13281);
xnor U13603 (N_13603,N_13473,N_13211);
or U13604 (N_13604,N_13482,N_13498);
and U13605 (N_13605,N_13440,N_13451);
nand U13606 (N_13606,N_13426,N_13330);
or U13607 (N_13607,N_13233,N_13310);
or U13608 (N_13608,N_13261,N_13356);
or U13609 (N_13609,N_13468,N_13237);
or U13610 (N_13610,N_13421,N_13340);
or U13611 (N_13611,N_13441,N_13316);
nor U13612 (N_13612,N_13385,N_13207);
nand U13613 (N_13613,N_13490,N_13268);
nand U13614 (N_13614,N_13434,N_13234);
nor U13615 (N_13615,N_13499,N_13242);
and U13616 (N_13616,N_13222,N_13212);
nor U13617 (N_13617,N_13236,N_13382);
nor U13618 (N_13618,N_13215,N_13302);
nor U13619 (N_13619,N_13226,N_13208);
nor U13620 (N_13620,N_13301,N_13477);
nor U13621 (N_13621,N_13414,N_13335);
nor U13622 (N_13622,N_13249,N_13354);
xor U13623 (N_13623,N_13274,N_13287);
and U13624 (N_13624,N_13314,N_13391);
nor U13625 (N_13625,N_13235,N_13437);
and U13626 (N_13626,N_13457,N_13405);
xor U13627 (N_13627,N_13348,N_13494);
or U13628 (N_13628,N_13300,N_13325);
nand U13629 (N_13629,N_13336,N_13399);
nand U13630 (N_13630,N_13218,N_13395);
nor U13631 (N_13631,N_13436,N_13203);
nor U13632 (N_13632,N_13419,N_13321);
or U13633 (N_13633,N_13246,N_13214);
and U13634 (N_13634,N_13343,N_13276);
xor U13635 (N_13635,N_13292,N_13412);
xnor U13636 (N_13636,N_13220,N_13365);
xnor U13637 (N_13637,N_13493,N_13447);
and U13638 (N_13638,N_13210,N_13366);
or U13639 (N_13639,N_13290,N_13362);
xnor U13640 (N_13640,N_13257,N_13265);
and U13641 (N_13641,N_13303,N_13449);
xnor U13642 (N_13642,N_13338,N_13429);
and U13643 (N_13643,N_13275,N_13495);
nand U13644 (N_13644,N_13484,N_13431);
and U13645 (N_13645,N_13239,N_13472);
xor U13646 (N_13646,N_13458,N_13442);
xor U13647 (N_13647,N_13452,N_13216);
xnor U13648 (N_13648,N_13384,N_13205);
and U13649 (N_13649,N_13277,N_13245);
nand U13650 (N_13650,N_13338,N_13400);
and U13651 (N_13651,N_13461,N_13441);
and U13652 (N_13652,N_13467,N_13342);
xnor U13653 (N_13653,N_13407,N_13340);
nor U13654 (N_13654,N_13371,N_13372);
or U13655 (N_13655,N_13210,N_13400);
nor U13656 (N_13656,N_13336,N_13231);
nor U13657 (N_13657,N_13466,N_13375);
xor U13658 (N_13658,N_13484,N_13404);
xnor U13659 (N_13659,N_13478,N_13421);
nand U13660 (N_13660,N_13482,N_13329);
or U13661 (N_13661,N_13290,N_13286);
and U13662 (N_13662,N_13347,N_13218);
or U13663 (N_13663,N_13277,N_13291);
and U13664 (N_13664,N_13212,N_13416);
nand U13665 (N_13665,N_13385,N_13476);
nor U13666 (N_13666,N_13485,N_13404);
and U13667 (N_13667,N_13305,N_13293);
xnor U13668 (N_13668,N_13496,N_13370);
nand U13669 (N_13669,N_13414,N_13453);
and U13670 (N_13670,N_13495,N_13355);
nand U13671 (N_13671,N_13329,N_13266);
xor U13672 (N_13672,N_13331,N_13360);
or U13673 (N_13673,N_13282,N_13451);
nand U13674 (N_13674,N_13451,N_13447);
nand U13675 (N_13675,N_13431,N_13302);
nor U13676 (N_13676,N_13403,N_13353);
or U13677 (N_13677,N_13484,N_13368);
or U13678 (N_13678,N_13303,N_13363);
and U13679 (N_13679,N_13479,N_13379);
and U13680 (N_13680,N_13221,N_13209);
and U13681 (N_13681,N_13495,N_13376);
or U13682 (N_13682,N_13258,N_13364);
nand U13683 (N_13683,N_13253,N_13383);
nor U13684 (N_13684,N_13232,N_13215);
xor U13685 (N_13685,N_13313,N_13300);
and U13686 (N_13686,N_13367,N_13359);
nand U13687 (N_13687,N_13402,N_13305);
and U13688 (N_13688,N_13321,N_13409);
xnor U13689 (N_13689,N_13391,N_13399);
or U13690 (N_13690,N_13402,N_13310);
or U13691 (N_13691,N_13361,N_13449);
or U13692 (N_13692,N_13416,N_13441);
or U13693 (N_13693,N_13256,N_13290);
and U13694 (N_13694,N_13396,N_13449);
or U13695 (N_13695,N_13325,N_13299);
xor U13696 (N_13696,N_13438,N_13235);
xnor U13697 (N_13697,N_13238,N_13390);
nor U13698 (N_13698,N_13276,N_13250);
or U13699 (N_13699,N_13355,N_13310);
or U13700 (N_13700,N_13386,N_13472);
nand U13701 (N_13701,N_13349,N_13285);
xnor U13702 (N_13702,N_13225,N_13378);
or U13703 (N_13703,N_13462,N_13486);
and U13704 (N_13704,N_13314,N_13390);
nand U13705 (N_13705,N_13207,N_13258);
and U13706 (N_13706,N_13392,N_13342);
nand U13707 (N_13707,N_13215,N_13308);
or U13708 (N_13708,N_13205,N_13227);
and U13709 (N_13709,N_13246,N_13406);
or U13710 (N_13710,N_13255,N_13471);
nand U13711 (N_13711,N_13355,N_13289);
or U13712 (N_13712,N_13368,N_13370);
and U13713 (N_13713,N_13457,N_13412);
xor U13714 (N_13714,N_13318,N_13432);
and U13715 (N_13715,N_13269,N_13358);
nor U13716 (N_13716,N_13309,N_13254);
nand U13717 (N_13717,N_13494,N_13488);
nand U13718 (N_13718,N_13472,N_13368);
nand U13719 (N_13719,N_13417,N_13490);
nor U13720 (N_13720,N_13248,N_13204);
nand U13721 (N_13721,N_13402,N_13390);
nor U13722 (N_13722,N_13297,N_13317);
nor U13723 (N_13723,N_13274,N_13337);
nand U13724 (N_13724,N_13396,N_13489);
xnor U13725 (N_13725,N_13352,N_13223);
nand U13726 (N_13726,N_13444,N_13208);
and U13727 (N_13727,N_13401,N_13323);
or U13728 (N_13728,N_13215,N_13212);
and U13729 (N_13729,N_13445,N_13284);
xor U13730 (N_13730,N_13379,N_13294);
or U13731 (N_13731,N_13301,N_13384);
or U13732 (N_13732,N_13241,N_13260);
nand U13733 (N_13733,N_13240,N_13488);
or U13734 (N_13734,N_13337,N_13229);
or U13735 (N_13735,N_13497,N_13466);
nor U13736 (N_13736,N_13270,N_13247);
nand U13737 (N_13737,N_13247,N_13364);
or U13738 (N_13738,N_13488,N_13274);
nand U13739 (N_13739,N_13256,N_13458);
xor U13740 (N_13740,N_13436,N_13280);
or U13741 (N_13741,N_13319,N_13323);
or U13742 (N_13742,N_13366,N_13250);
nand U13743 (N_13743,N_13443,N_13498);
or U13744 (N_13744,N_13463,N_13293);
nand U13745 (N_13745,N_13394,N_13345);
and U13746 (N_13746,N_13204,N_13407);
nor U13747 (N_13747,N_13247,N_13441);
xor U13748 (N_13748,N_13432,N_13306);
nor U13749 (N_13749,N_13301,N_13479);
xnor U13750 (N_13750,N_13464,N_13431);
nand U13751 (N_13751,N_13491,N_13273);
nor U13752 (N_13752,N_13205,N_13424);
nor U13753 (N_13753,N_13241,N_13225);
xor U13754 (N_13754,N_13415,N_13423);
nor U13755 (N_13755,N_13277,N_13203);
and U13756 (N_13756,N_13248,N_13470);
nand U13757 (N_13757,N_13470,N_13389);
and U13758 (N_13758,N_13343,N_13389);
xor U13759 (N_13759,N_13224,N_13343);
xor U13760 (N_13760,N_13390,N_13391);
nand U13761 (N_13761,N_13358,N_13207);
nand U13762 (N_13762,N_13450,N_13268);
nor U13763 (N_13763,N_13249,N_13335);
nand U13764 (N_13764,N_13206,N_13465);
nand U13765 (N_13765,N_13263,N_13315);
nand U13766 (N_13766,N_13261,N_13455);
nand U13767 (N_13767,N_13481,N_13344);
and U13768 (N_13768,N_13216,N_13378);
xnor U13769 (N_13769,N_13204,N_13381);
nor U13770 (N_13770,N_13349,N_13278);
and U13771 (N_13771,N_13362,N_13464);
and U13772 (N_13772,N_13407,N_13256);
and U13773 (N_13773,N_13476,N_13224);
or U13774 (N_13774,N_13348,N_13456);
nor U13775 (N_13775,N_13212,N_13388);
nand U13776 (N_13776,N_13257,N_13206);
or U13777 (N_13777,N_13287,N_13494);
nor U13778 (N_13778,N_13377,N_13393);
and U13779 (N_13779,N_13346,N_13374);
xnor U13780 (N_13780,N_13218,N_13271);
or U13781 (N_13781,N_13462,N_13481);
nand U13782 (N_13782,N_13375,N_13353);
and U13783 (N_13783,N_13421,N_13263);
and U13784 (N_13784,N_13457,N_13433);
xnor U13785 (N_13785,N_13415,N_13446);
nand U13786 (N_13786,N_13241,N_13436);
xnor U13787 (N_13787,N_13208,N_13403);
xnor U13788 (N_13788,N_13231,N_13275);
and U13789 (N_13789,N_13312,N_13465);
and U13790 (N_13790,N_13259,N_13480);
and U13791 (N_13791,N_13410,N_13347);
xnor U13792 (N_13792,N_13463,N_13453);
or U13793 (N_13793,N_13392,N_13315);
nor U13794 (N_13794,N_13230,N_13487);
xnor U13795 (N_13795,N_13293,N_13467);
xor U13796 (N_13796,N_13365,N_13202);
xnor U13797 (N_13797,N_13406,N_13319);
nand U13798 (N_13798,N_13271,N_13469);
xnor U13799 (N_13799,N_13484,N_13315);
and U13800 (N_13800,N_13737,N_13503);
or U13801 (N_13801,N_13707,N_13629);
nand U13802 (N_13802,N_13637,N_13730);
or U13803 (N_13803,N_13510,N_13669);
or U13804 (N_13804,N_13766,N_13759);
or U13805 (N_13805,N_13530,N_13745);
or U13806 (N_13806,N_13512,N_13645);
or U13807 (N_13807,N_13580,N_13788);
nor U13808 (N_13808,N_13733,N_13571);
nor U13809 (N_13809,N_13704,N_13721);
or U13810 (N_13810,N_13662,N_13652);
nand U13811 (N_13811,N_13622,N_13750);
or U13812 (N_13812,N_13516,N_13654);
or U13813 (N_13813,N_13584,N_13687);
nor U13814 (N_13814,N_13798,N_13633);
or U13815 (N_13815,N_13736,N_13760);
and U13816 (N_13816,N_13561,N_13656);
or U13817 (N_13817,N_13749,N_13781);
nand U13818 (N_13818,N_13702,N_13794);
xor U13819 (N_13819,N_13641,N_13665);
nor U13820 (N_13820,N_13603,N_13799);
nor U13821 (N_13821,N_13559,N_13536);
nor U13822 (N_13822,N_13617,N_13767);
nor U13823 (N_13823,N_13556,N_13706);
nor U13824 (N_13824,N_13797,N_13661);
and U13825 (N_13825,N_13623,N_13522);
nand U13826 (N_13826,N_13588,N_13548);
nor U13827 (N_13827,N_13775,N_13677);
and U13828 (N_13828,N_13583,N_13500);
nand U13829 (N_13829,N_13607,N_13626);
xnor U13830 (N_13830,N_13533,N_13614);
nand U13831 (N_13831,N_13732,N_13685);
nor U13832 (N_13832,N_13529,N_13589);
nand U13833 (N_13833,N_13710,N_13593);
nor U13834 (N_13834,N_13755,N_13528);
nor U13835 (N_13835,N_13748,N_13783);
nor U13836 (N_13836,N_13776,N_13769);
nand U13837 (N_13837,N_13686,N_13703);
and U13838 (N_13838,N_13586,N_13664);
nand U13839 (N_13839,N_13729,N_13558);
and U13840 (N_13840,N_13765,N_13563);
xnor U13841 (N_13841,N_13609,N_13555);
xor U13842 (N_13842,N_13658,N_13523);
or U13843 (N_13843,N_13735,N_13544);
nand U13844 (N_13844,N_13666,N_13615);
xnor U13845 (N_13845,N_13791,N_13521);
and U13846 (N_13846,N_13597,N_13671);
and U13847 (N_13847,N_13587,N_13722);
xor U13848 (N_13848,N_13624,N_13688);
nor U13849 (N_13849,N_13782,N_13764);
xnor U13850 (N_13850,N_13551,N_13640);
or U13851 (N_13851,N_13660,N_13509);
nor U13852 (N_13852,N_13594,N_13646);
nor U13853 (N_13853,N_13604,N_13742);
nor U13854 (N_13854,N_13634,N_13507);
nor U13855 (N_13855,N_13647,N_13692);
or U13856 (N_13856,N_13743,N_13501);
nand U13857 (N_13857,N_13773,N_13793);
and U13858 (N_13858,N_13600,N_13699);
xor U13859 (N_13859,N_13680,N_13642);
or U13860 (N_13860,N_13540,N_13545);
nand U13861 (N_13861,N_13504,N_13700);
xor U13862 (N_13862,N_13638,N_13569);
and U13863 (N_13863,N_13689,N_13562);
or U13864 (N_13864,N_13630,N_13570);
or U13865 (N_13865,N_13681,N_13649);
or U13866 (N_13866,N_13653,N_13602);
nand U13867 (N_13867,N_13713,N_13711);
nor U13868 (N_13868,N_13754,N_13554);
and U13869 (N_13869,N_13506,N_13717);
nand U13870 (N_13870,N_13605,N_13628);
nor U13871 (N_13871,N_13574,N_13549);
nand U13872 (N_13872,N_13519,N_13596);
nand U13873 (N_13873,N_13655,N_13768);
nand U13874 (N_13874,N_13663,N_13560);
nor U13875 (N_13875,N_13619,N_13673);
and U13876 (N_13876,N_13728,N_13753);
xor U13877 (N_13877,N_13771,N_13705);
nor U13878 (N_13878,N_13632,N_13716);
nand U13879 (N_13879,N_13591,N_13751);
or U13880 (N_13880,N_13547,N_13756);
xor U13881 (N_13881,N_13514,N_13727);
xor U13882 (N_13882,N_13541,N_13770);
xnor U13883 (N_13883,N_13785,N_13608);
nor U13884 (N_13884,N_13650,N_13684);
nand U13885 (N_13885,N_13592,N_13532);
xor U13886 (N_13886,N_13726,N_13724);
xor U13887 (N_13887,N_13772,N_13508);
or U13888 (N_13888,N_13599,N_13696);
nand U13889 (N_13889,N_13675,N_13659);
nand U13890 (N_13890,N_13567,N_13734);
and U13891 (N_13891,N_13566,N_13564);
nor U13892 (N_13892,N_13698,N_13678);
nand U13893 (N_13893,N_13511,N_13635);
and U13894 (N_13894,N_13520,N_13789);
nor U13895 (N_13895,N_13670,N_13505);
and U13896 (N_13896,N_13796,N_13525);
nand U13897 (N_13897,N_13553,N_13513);
or U13898 (N_13898,N_13774,N_13543);
nor U13899 (N_13899,N_13693,N_13568);
or U13900 (N_13900,N_13757,N_13674);
or U13901 (N_13901,N_13601,N_13612);
or U13902 (N_13902,N_13683,N_13777);
nor U13903 (N_13903,N_13731,N_13701);
nor U13904 (N_13904,N_13719,N_13787);
xor U13905 (N_13905,N_13582,N_13744);
nor U13906 (N_13906,N_13578,N_13621);
or U13907 (N_13907,N_13740,N_13778);
or U13908 (N_13908,N_13534,N_13739);
nand U13909 (N_13909,N_13610,N_13723);
xnor U13910 (N_13910,N_13552,N_13780);
or U13911 (N_13911,N_13747,N_13576);
or U13912 (N_13912,N_13682,N_13657);
and U13913 (N_13913,N_13577,N_13531);
nor U13914 (N_13914,N_13679,N_13667);
or U13915 (N_13915,N_13651,N_13518);
and U13916 (N_13916,N_13546,N_13738);
nor U13917 (N_13917,N_13527,N_13515);
or U13918 (N_13918,N_13537,N_13694);
and U13919 (N_13919,N_13572,N_13676);
nor U13920 (N_13920,N_13595,N_13565);
and U13921 (N_13921,N_13590,N_13725);
xor U13922 (N_13922,N_13672,N_13763);
nand U13923 (N_13923,N_13636,N_13535);
nand U13924 (N_13924,N_13720,N_13697);
and U13925 (N_13925,N_13539,N_13585);
xnor U13926 (N_13926,N_13611,N_13538);
and U13927 (N_13927,N_13668,N_13708);
and U13928 (N_13928,N_13639,N_13709);
xor U13929 (N_13929,N_13690,N_13648);
nor U13930 (N_13930,N_13784,N_13598);
and U13931 (N_13931,N_13752,N_13761);
nand U13932 (N_13932,N_13502,N_13550);
xnor U13933 (N_13933,N_13718,N_13762);
nor U13934 (N_13934,N_13695,N_13792);
nand U13935 (N_13935,N_13573,N_13691);
or U13936 (N_13936,N_13631,N_13712);
or U13937 (N_13937,N_13575,N_13715);
and U13938 (N_13938,N_13613,N_13746);
and U13939 (N_13939,N_13790,N_13643);
nand U13940 (N_13940,N_13526,N_13644);
or U13941 (N_13941,N_13581,N_13524);
nor U13942 (N_13942,N_13795,N_13618);
xnor U13943 (N_13943,N_13714,N_13517);
xor U13944 (N_13944,N_13579,N_13758);
or U13945 (N_13945,N_13542,N_13557);
nor U13946 (N_13946,N_13606,N_13625);
or U13947 (N_13947,N_13741,N_13616);
xor U13948 (N_13948,N_13786,N_13620);
nor U13949 (N_13949,N_13627,N_13779);
nand U13950 (N_13950,N_13542,N_13740);
or U13951 (N_13951,N_13518,N_13778);
xor U13952 (N_13952,N_13595,N_13637);
or U13953 (N_13953,N_13610,N_13541);
nand U13954 (N_13954,N_13759,N_13617);
nand U13955 (N_13955,N_13680,N_13787);
and U13956 (N_13956,N_13762,N_13629);
nand U13957 (N_13957,N_13774,N_13756);
xor U13958 (N_13958,N_13627,N_13743);
xnor U13959 (N_13959,N_13634,N_13626);
xnor U13960 (N_13960,N_13518,N_13562);
nand U13961 (N_13961,N_13709,N_13762);
or U13962 (N_13962,N_13750,N_13693);
nor U13963 (N_13963,N_13796,N_13595);
or U13964 (N_13964,N_13635,N_13621);
nor U13965 (N_13965,N_13533,N_13776);
or U13966 (N_13966,N_13605,N_13765);
nor U13967 (N_13967,N_13694,N_13759);
nand U13968 (N_13968,N_13745,N_13514);
xnor U13969 (N_13969,N_13715,N_13589);
nand U13970 (N_13970,N_13658,N_13719);
nand U13971 (N_13971,N_13772,N_13778);
and U13972 (N_13972,N_13552,N_13536);
nand U13973 (N_13973,N_13584,N_13647);
nand U13974 (N_13974,N_13716,N_13697);
or U13975 (N_13975,N_13753,N_13737);
nand U13976 (N_13976,N_13730,N_13608);
nand U13977 (N_13977,N_13614,N_13587);
or U13978 (N_13978,N_13747,N_13666);
nor U13979 (N_13979,N_13547,N_13795);
xnor U13980 (N_13980,N_13607,N_13523);
nand U13981 (N_13981,N_13692,N_13555);
nor U13982 (N_13982,N_13707,N_13660);
nor U13983 (N_13983,N_13656,N_13504);
and U13984 (N_13984,N_13601,N_13639);
and U13985 (N_13985,N_13622,N_13788);
nand U13986 (N_13986,N_13679,N_13614);
and U13987 (N_13987,N_13597,N_13515);
or U13988 (N_13988,N_13547,N_13501);
xnor U13989 (N_13989,N_13693,N_13703);
and U13990 (N_13990,N_13505,N_13760);
nor U13991 (N_13991,N_13611,N_13598);
nand U13992 (N_13992,N_13582,N_13542);
nand U13993 (N_13993,N_13506,N_13711);
nor U13994 (N_13994,N_13637,N_13550);
nor U13995 (N_13995,N_13646,N_13762);
or U13996 (N_13996,N_13613,N_13636);
and U13997 (N_13997,N_13539,N_13776);
xor U13998 (N_13998,N_13640,N_13667);
and U13999 (N_13999,N_13511,N_13577);
xnor U14000 (N_14000,N_13647,N_13753);
or U14001 (N_14001,N_13757,N_13789);
or U14002 (N_14002,N_13598,N_13544);
nand U14003 (N_14003,N_13501,N_13625);
nor U14004 (N_14004,N_13743,N_13629);
and U14005 (N_14005,N_13729,N_13769);
nand U14006 (N_14006,N_13548,N_13693);
or U14007 (N_14007,N_13517,N_13650);
nor U14008 (N_14008,N_13764,N_13574);
xor U14009 (N_14009,N_13719,N_13690);
or U14010 (N_14010,N_13584,N_13595);
xor U14011 (N_14011,N_13509,N_13780);
nand U14012 (N_14012,N_13588,N_13659);
and U14013 (N_14013,N_13798,N_13593);
nand U14014 (N_14014,N_13788,N_13728);
nand U14015 (N_14015,N_13692,N_13652);
and U14016 (N_14016,N_13698,N_13668);
nor U14017 (N_14017,N_13775,N_13779);
xnor U14018 (N_14018,N_13714,N_13775);
xor U14019 (N_14019,N_13587,N_13565);
and U14020 (N_14020,N_13578,N_13525);
and U14021 (N_14021,N_13689,N_13781);
xnor U14022 (N_14022,N_13722,N_13545);
or U14023 (N_14023,N_13752,N_13647);
nand U14024 (N_14024,N_13542,N_13504);
nand U14025 (N_14025,N_13631,N_13779);
nor U14026 (N_14026,N_13518,N_13631);
nand U14027 (N_14027,N_13588,N_13572);
nand U14028 (N_14028,N_13525,N_13598);
or U14029 (N_14029,N_13540,N_13767);
nand U14030 (N_14030,N_13636,N_13562);
nor U14031 (N_14031,N_13788,N_13751);
or U14032 (N_14032,N_13589,N_13647);
xor U14033 (N_14033,N_13509,N_13711);
or U14034 (N_14034,N_13560,N_13606);
and U14035 (N_14035,N_13751,N_13771);
nor U14036 (N_14036,N_13717,N_13764);
xnor U14037 (N_14037,N_13775,N_13623);
or U14038 (N_14038,N_13733,N_13798);
nor U14039 (N_14039,N_13696,N_13685);
and U14040 (N_14040,N_13533,N_13674);
nand U14041 (N_14041,N_13537,N_13632);
nor U14042 (N_14042,N_13664,N_13658);
nor U14043 (N_14043,N_13664,N_13581);
nor U14044 (N_14044,N_13532,N_13570);
nor U14045 (N_14045,N_13749,N_13563);
xor U14046 (N_14046,N_13602,N_13748);
or U14047 (N_14047,N_13768,N_13649);
xnor U14048 (N_14048,N_13766,N_13692);
xor U14049 (N_14049,N_13708,N_13631);
or U14050 (N_14050,N_13520,N_13716);
nor U14051 (N_14051,N_13604,N_13706);
xnor U14052 (N_14052,N_13529,N_13797);
nor U14053 (N_14053,N_13591,N_13755);
and U14054 (N_14054,N_13632,N_13605);
and U14055 (N_14055,N_13714,N_13709);
and U14056 (N_14056,N_13569,N_13767);
and U14057 (N_14057,N_13657,N_13744);
or U14058 (N_14058,N_13631,N_13746);
xnor U14059 (N_14059,N_13714,N_13608);
nor U14060 (N_14060,N_13667,N_13603);
xnor U14061 (N_14061,N_13776,N_13642);
nand U14062 (N_14062,N_13523,N_13651);
and U14063 (N_14063,N_13505,N_13629);
and U14064 (N_14064,N_13612,N_13710);
xor U14065 (N_14065,N_13561,N_13632);
xnor U14066 (N_14066,N_13590,N_13734);
nor U14067 (N_14067,N_13617,N_13628);
nor U14068 (N_14068,N_13678,N_13585);
xor U14069 (N_14069,N_13509,N_13698);
and U14070 (N_14070,N_13717,N_13679);
nor U14071 (N_14071,N_13518,N_13610);
nor U14072 (N_14072,N_13539,N_13728);
and U14073 (N_14073,N_13529,N_13575);
xnor U14074 (N_14074,N_13795,N_13643);
and U14075 (N_14075,N_13620,N_13756);
xor U14076 (N_14076,N_13570,N_13652);
nand U14077 (N_14077,N_13651,N_13693);
nor U14078 (N_14078,N_13772,N_13766);
xnor U14079 (N_14079,N_13603,N_13725);
xnor U14080 (N_14080,N_13734,N_13614);
nor U14081 (N_14081,N_13654,N_13546);
nor U14082 (N_14082,N_13554,N_13750);
xor U14083 (N_14083,N_13677,N_13661);
or U14084 (N_14084,N_13724,N_13621);
xor U14085 (N_14085,N_13663,N_13582);
or U14086 (N_14086,N_13798,N_13758);
nand U14087 (N_14087,N_13675,N_13577);
xor U14088 (N_14088,N_13619,N_13658);
nor U14089 (N_14089,N_13586,N_13593);
nor U14090 (N_14090,N_13737,N_13641);
nand U14091 (N_14091,N_13664,N_13599);
nor U14092 (N_14092,N_13629,N_13721);
nand U14093 (N_14093,N_13641,N_13609);
nor U14094 (N_14094,N_13669,N_13600);
nor U14095 (N_14095,N_13529,N_13642);
nor U14096 (N_14096,N_13788,N_13513);
nor U14097 (N_14097,N_13510,N_13617);
xnor U14098 (N_14098,N_13734,N_13604);
nand U14099 (N_14099,N_13718,N_13713);
nand U14100 (N_14100,N_14091,N_14099);
nand U14101 (N_14101,N_13892,N_13812);
nand U14102 (N_14102,N_13917,N_13807);
xor U14103 (N_14103,N_13888,N_13981);
and U14104 (N_14104,N_13989,N_13958);
or U14105 (N_14105,N_13819,N_13928);
nand U14106 (N_14106,N_13967,N_13953);
or U14107 (N_14107,N_13907,N_13859);
nand U14108 (N_14108,N_14017,N_14065);
or U14109 (N_14109,N_13978,N_13864);
or U14110 (N_14110,N_13988,N_13912);
xor U14111 (N_14111,N_14072,N_13915);
or U14112 (N_14112,N_13946,N_13849);
or U14113 (N_14113,N_13972,N_13830);
or U14114 (N_14114,N_13863,N_14011);
nand U14115 (N_14115,N_14097,N_14003);
or U14116 (N_14116,N_13964,N_13836);
xnor U14117 (N_14117,N_13882,N_14063);
nor U14118 (N_14118,N_13870,N_13889);
or U14119 (N_14119,N_14048,N_14031);
and U14120 (N_14120,N_13977,N_13885);
nand U14121 (N_14121,N_13848,N_13987);
xnor U14122 (N_14122,N_13966,N_13916);
nand U14123 (N_14123,N_13918,N_14037);
nand U14124 (N_14124,N_14002,N_13858);
nand U14125 (N_14125,N_13832,N_14067);
or U14126 (N_14126,N_13890,N_14057);
nor U14127 (N_14127,N_13905,N_13960);
nor U14128 (N_14128,N_13910,N_13996);
and U14129 (N_14129,N_13865,N_13846);
or U14130 (N_14130,N_14073,N_14000);
and U14131 (N_14131,N_14039,N_14047);
or U14132 (N_14132,N_13990,N_13800);
xor U14133 (N_14133,N_13940,N_14081);
nor U14134 (N_14134,N_13976,N_13923);
nand U14135 (N_14135,N_14025,N_14012);
xor U14136 (N_14136,N_14082,N_13901);
nand U14137 (N_14137,N_13852,N_14059);
nand U14138 (N_14138,N_13855,N_13862);
nand U14139 (N_14139,N_13851,N_13929);
or U14140 (N_14140,N_14070,N_14060);
xnor U14141 (N_14141,N_13809,N_14096);
or U14142 (N_14142,N_14071,N_14089);
nand U14143 (N_14143,N_13939,N_14041);
nand U14144 (N_14144,N_13974,N_14093);
xnor U14145 (N_14145,N_13995,N_13844);
xnor U14146 (N_14146,N_13876,N_13970);
and U14147 (N_14147,N_13932,N_13980);
nand U14148 (N_14148,N_14098,N_14054);
xor U14149 (N_14149,N_13948,N_13947);
xor U14150 (N_14150,N_13914,N_14049);
or U14151 (N_14151,N_13934,N_13826);
or U14152 (N_14152,N_14009,N_13810);
xor U14153 (N_14153,N_13897,N_14026);
nor U14154 (N_14154,N_13969,N_13945);
and U14155 (N_14155,N_13881,N_13959);
xor U14156 (N_14156,N_14005,N_14038);
nor U14157 (N_14157,N_13825,N_13823);
nand U14158 (N_14158,N_13839,N_13963);
nor U14159 (N_14159,N_14007,N_13984);
nor U14160 (N_14160,N_14020,N_14004);
and U14161 (N_14161,N_14094,N_13886);
nor U14162 (N_14162,N_13982,N_13931);
nor U14163 (N_14163,N_13815,N_14046);
xor U14164 (N_14164,N_14050,N_13922);
or U14165 (N_14165,N_13942,N_13871);
nor U14166 (N_14166,N_13983,N_13822);
nor U14167 (N_14167,N_13861,N_14058);
and U14168 (N_14168,N_14016,N_13971);
or U14169 (N_14169,N_14064,N_13986);
or U14170 (N_14170,N_13903,N_13944);
or U14171 (N_14171,N_13962,N_13880);
and U14172 (N_14172,N_14092,N_14053);
xor U14173 (N_14173,N_14006,N_13868);
nor U14174 (N_14174,N_14030,N_13821);
and U14175 (N_14175,N_13933,N_13814);
xnor U14176 (N_14176,N_13884,N_14034);
xnor U14177 (N_14177,N_13896,N_13993);
xnor U14178 (N_14178,N_13853,N_13833);
xor U14179 (N_14179,N_14027,N_13921);
nand U14180 (N_14180,N_13919,N_13818);
and U14181 (N_14181,N_14084,N_13999);
nand U14182 (N_14182,N_13994,N_13893);
xor U14183 (N_14183,N_14036,N_14035);
and U14184 (N_14184,N_13911,N_13828);
nor U14185 (N_14185,N_13956,N_13873);
xor U14186 (N_14186,N_13866,N_13951);
xor U14187 (N_14187,N_13834,N_13930);
and U14188 (N_14188,N_13879,N_14066);
xnor U14189 (N_14189,N_14079,N_14023);
xor U14190 (N_14190,N_13829,N_13900);
xnor U14191 (N_14191,N_14010,N_13998);
nand U14192 (N_14192,N_13902,N_14051);
or U14193 (N_14193,N_13992,N_13904);
nor U14194 (N_14194,N_14008,N_13816);
and U14195 (N_14195,N_13968,N_13950);
nor U14196 (N_14196,N_13979,N_13906);
and U14197 (N_14197,N_13935,N_14088);
xor U14198 (N_14198,N_13891,N_13867);
or U14199 (N_14199,N_13831,N_13803);
xor U14200 (N_14200,N_13883,N_13806);
xnor U14201 (N_14201,N_14086,N_13965);
nand U14202 (N_14202,N_13952,N_13874);
nor U14203 (N_14203,N_13899,N_13869);
and U14204 (N_14204,N_14083,N_13924);
nor U14205 (N_14205,N_14078,N_13827);
nand U14206 (N_14206,N_14087,N_13840);
xor U14207 (N_14207,N_13847,N_13801);
and U14208 (N_14208,N_13949,N_13837);
and U14209 (N_14209,N_13813,N_13926);
xor U14210 (N_14210,N_14028,N_13909);
and U14211 (N_14211,N_13887,N_13898);
and U14212 (N_14212,N_14040,N_14077);
nor U14213 (N_14213,N_13843,N_13850);
xor U14214 (N_14214,N_14018,N_13872);
and U14215 (N_14215,N_14085,N_13941);
nor U14216 (N_14216,N_13937,N_13835);
xnor U14217 (N_14217,N_14022,N_13808);
nand U14218 (N_14218,N_14052,N_13811);
nor U14219 (N_14219,N_14042,N_13860);
nor U14220 (N_14220,N_13802,N_14032);
and U14221 (N_14221,N_14068,N_14076);
xor U14222 (N_14222,N_13842,N_14062);
nor U14223 (N_14223,N_13973,N_13854);
and U14224 (N_14224,N_13927,N_13997);
xor U14225 (N_14225,N_14069,N_14090);
xor U14226 (N_14226,N_13943,N_13878);
nand U14227 (N_14227,N_14033,N_14043);
and U14228 (N_14228,N_14013,N_13908);
or U14229 (N_14229,N_14001,N_14045);
or U14230 (N_14230,N_13925,N_13975);
and U14231 (N_14231,N_13985,N_13961);
and U14232 (N_14232,N_13845,N_14095);
nand U14233 (N_14233,N_13838,N_13820);
and U14234 (N_14234,N_13936,N_13920);
xor U14235 (N_14235,N_14014,N_13894);
nor U14236 (N_14236,N_13895,N_13954);
nor U14237 (N_14237,N_13913,N_14055);
or U14238 (N_14238,N_14024,N_14056);
xor U14239 (N_14239,N_13804,N_13955);
and U14240 (N_14240,N_14061,N_14075);
and U14241 (N_14241,N_14029,N_14080);
nand U14242 (N_14242,N_13957,N_13938);
nor U14243 (N_14243,N_13856,N_13824);
nor U14244 (N_14244,N_14015,N_13991);
or U14245 (N_14245,N_13877,N_13857);
xnor U14246 (N_14246,N_14074,N_13805);
xor U14247 (N_14247,N_14021,N_14019);
nand U14248 (N_14248,N_13875,N_13817);
nor U14249 (N_14249,N_13841,N_14044);
or U14250 (N_14250,N_14041,N_14066);
xor U14251 (N_14251,N_13889,N_13930);
or U14252 (N_14252,N_13851,N_13947);
xnor U14253 (N_14253,N_13928,N_13812);
nand U14254 (N_14254,N_13977,N_14052);
nor U14255 (N_14255,N_13911,N_13839);
or U14256 (N_14256,N_13832,N_13916);
and U14257 (N_14257,N_13926,N_13963);
nand U14258 (N_14258,N_13892,N_13934);
nand U14259 (N_14259,N_13838,N_13966);
or U14260 (N_14260,N_14030,N_13843);
and U14261 (N_14261,N_14041,N_14005);
nand U14262 (N_14262,N_13803,N_13887);
nor U14263 (N_14263,N_14096,N_13812);
xor U14264 (N_14264,N_13817,N_13807);
xor U14265 (N_14265,N_13826,N_13834);
or U14266 (N_14266,N_13813,N_13843);
nand U14267 (N_14267,N_14021,N_13946);
or U14268 (N_14268,N_13940,N_13985);
xor U14269 (N_14269,N_14018,N_13831);
and U14270 (N_14270,N_14012,N_13890);
nor U14271 (N_14271,N_13879,N_13828);
or U14272 (N_14272,N_14026,N_14093);
and U14273 (N_14273,N_14063,N_13933);
or U14274 (N_14274,N_14024,N_13990);
nor U14275 (N_14275,N_13994,N_13915);
nand U14276 (N_14276,N_14008,N_13990);
nand U14277 (N_14277,N_13933,N_13857);
and U14278 (N_14278,N_13860,N_13980);
or U14279 (N_14279,N_13928,N_13856);
nor U14280 (N_14280,N_14052,N_13853);
or U14281 (N_14281,N_13819,N_13902);
or U14282 (N_14282,N_14064,N_14009);
nand U14283 (N_14283,N_14069,N_13810);
xor U14284 (N_14284,N_14006,N_13941);
nor U14285 (N_14285,N_14047,N_13985);
and U14286 (N_14286,N_13805,N_13877);
xnor U14287 (N_14287,N_13929,N_13952);
or U14288 (N_14288,N_13875,N_14081);
and U14289 (N_14289,N_14056,N_14077);
nand U14290 (N_14290,N_13973,N_13879);
and U14291 (N_14291,N_13908,N_13807);
or U14292 (N_14292,N_13981,N_14034);
nor U14293 (N_14293,N_14055,N_13999);
xor U14294 (N_14294,N_13912,N_14017);
nor U14295 (N_14295,N_13987,N_13988);
nor U14296 (N_14296,N_13827,N_13936);
xnor U14297 (N_14297,N_13925,N_13828);
or U14298 (N_14298,N_14058,N_14061);
nand U14299 (N_14299,N_14018,N_14094);
nor U14300 (N_14300,N_13941,N_13909);
nand U14301 (N_14301,N_14021,N_14091);
and U14302 (N_14302,N_13818,N_13996);
and U14303 (N_14303,N_13862,N_13903);
or U14304 (N_14304,N_13893,N_13967);
nand U14305 (N_14305,N_13889,N_13822);
or U14306 (N_14306,N_13822,N_13949);
nand U14307 (N_14307,N_13958,N_13839);
xnor U14308 (N_14308,N_14097,N_13971);
or U14309 (N_14309,N_13994,N_13936);
nand U14310 (N_14310,N_14077,N_13871);
xor U14311 (N_14311,N_13813,N_13994);
or U14312 (N_14312,N_14089,N_14016);
nor U14313 (N_14313,N_13810,N_14025);
and U14314 (N_14314,N_13992,N_13917);
or U14315 (N_14315,N_14034,N_13948);
or U14316 (N_14316,N_13811,N_13934);
xnor U14317 (N_14317,N_13914,N_13874);
or U14318 (N_14318,N_13964,N_13911);
xnor U14319 (N_14319,N_13826,N_14043);
nor U14320 (N_14320,N_14005,N_13940);
nand U14321 (N_14321,N_14033,N_14062);
xnor U14322 (N_14322,N_13973,N_14088);
nand U14323 (N_14323,N_13907,N_13890);
nor U14324 (N_14324,N_13990,N_13926);
or U14325 (N_14325,N_13935,N_14028);
or U14326 (N_14326,N_14030,N_14091);
nand U14327 (N_14327,N_14032,N_13822);
nor U14328 (N_14328,N_14001,N_13870);
or U14329 (N_14329,N_14098,N_13838);
or U14330 (N_14330,N_13804,N_13947);
nor U14331 (N_14331,N_14061,N_13821);
or U14332 (N_14332,N_13993,N_13943);
nor U14333 (N_14333,N_13947,N_13872);
or U14334 (N_14334,N_13976,N_13996);
or U14335 (N_14335,N_13990,N_13984);
xor U14336 (N_14336,N_14009,N_14046);
xor U14337 (N_14337,N_13930,N_13925);
or U14338 (N_14338,N_13929,N_13957);
nor U14339 (N_14339,N_13990,N_13855);
or U14340 (N_14340,N_14046,N_13882);
and U14341 (N_14341,N_14050,N_14028);
nand U14342 (N_14342,N_14066,N_13860);
xor U14343 (N_14343,N_13846,N_13864);
or U14344 (N_14344,N_14087,N_13968);
nor U14345 (N_14345,N_13813,N_14093);
xor U14346 (N_14346,N_13948,N_14033);
xnor U14347 (N_14347,N_14029,N_13853);
nand U14348 (N_14348,N_14024,N_13972);
nor U14349 (N_14349,N_14028,N_13858);
xor U14350 (N_14350,N_13900,N_13911);
nor U14351 (N_14351,N_14065,N_13827);
nor U14352 (N_14352,N_14003,N_13933);
nand U14353 (N_14353,N_13816,N_13914);
xor U14354 (N_14354,N_14086,N_13912);
nand U14355 (N_14355,N_13895,N_13877);
nand U14356 (N_14356,N_13830,N_14054);
nor U14357 (N_14357,N_13963,N_13981);
and U14358 (N_14358,N_13955,N_13823);
or U14359 (N_14359,N_14036,N_14092);
or U14360 (N_14360,N_13863,N_13903);
or U14361 (N_14361,N_14062,N_13985);
or U14362 (N_14362,N_13978,N_14027);
or U14363 (N_14363,N_13906,N_13999);
nor U14364 (N_14364,N_13940,N_14002);
and U14365 (N_14365,N_13927,N_14052);
xor U14366 (N_14366,N_14009,N_13931);
nand U14367 (N_14367,N_14023,N_13886);
or U14368 (N_14368,N_13880,N_13819);
nor U14369 (N_14369,N_14073,N_14016);
and U14370 (N_14370,N_13891,N_14002);
nor U14371 (N_14371,N_13812,N_14020);
and U14372 (N_14372,N_14047,N_14019);
nor U14373 (N_14373,N_13946,N_13814);
nand U14374 (N_14374,N_13832,N_14087);
or U14375 (N_14375,N_13820,N_13883);
and U14376 (N_14376,N_13849,N_13831);
and U14377 (N_14377,N_13896,N_14041);
and U14378 (N_14378,N_13816,N_13986);
xnor U14379 (N_14379,N_13994,N_13974);
nand U14380 (N_14380,N_13964,N_13984);
or U14381 (N_14381,N_13859,N_13930);
and U14382 (N_14382,N_13826,N_14054);
and U14383 (N_14383,N_13943,N_14071);
xor U14384 (N_14384,N_13986,N_13971);
or U14385 (N_14385,N_13999,N_14029);
xor U14386 (N_14386,N_13942,N_14095);
and U14387 (N_14387,N_14070,N_14047);
or U14388 (N_14388,N_14071,N_14062);
xor U14389 (N_14389,N_13812,N_14048);
and U14390 (N_14390,N_13852,N_14040);
nor U14391 (N_14391,N_13981,N_14076);
nor U14392 (N_14392,N_13919,N_13839);
xor U14393 (N_14393,N_13971,N_13806);
xnor U14394 (N_14394,N_13945,N_13910);
nand U14395 (N_14395,N_13857,N_14038);
nor U14396 (N_14396,N_13922,N_13872);
xnor U14397 (N_14397,N_13832,N_13899);
nand U14398 (N_14398,N_13809,N_13983);
or U14399 (N_14399,N_14077,N_13964);
and U14400 (N_14400,N_14139,N_14117);
nand U14401 (N_14401,N_14383,N_14263);
or U14402 (N_14402,N_14202,N_14304);
nand U14403 (N_14403,N_14314,N_14367);
nor U14404 (N_14404,N_14363,N_14256);
or U14405 (N_14405,N_14209,N_14357);
or U14406 (N_14406,N_14102,N_14121);
xor U14407 (N_14407,N_14341,N_14328);
xnor U14408 (N_14408,N_14239,N_14258);
nor U14409 (N_14409,N_14307,N_14380);
nor U14410 (N_14410,N_14177,N_14199);
xnor U14411 (N_14411,N_14289,N_14377);
nand U14412 (N_14412,N_14134,N_14116);
nor U14413 (N_14413,N_14143,N_14349);
nor U14414 (N_14414,N_14294,N_14368);
nand U14415 (N_14415,N_14376,N_14128);
or U14416 (N_14416,N_14147,N_14171);
xor U14417 (N_14417,N_14397,N_14130);
or U14418 (N_14418,N_14293,N_14222);
and U14419 (N_14419,N_14246,N_14196);
nand U14420 (N_14420,N_14337,N_14306);
and U14421 (N_14421,N_14124,N_14142);
nor U14422 (N_14422,N_14122,N_14137);
nor U14423 (N_14423,N_14151,N_14141);
and U14424 (N_14424,N_14311,N_14149);
nand U14425 (N_14425,N_14150,N_14182);
or U14426 (N_14426,N_14242,N_14186);
nand U14427 (N_14427,N_14261,N_14131);
nand U14428 (N_14428,N_14206,N_14347);
nand U14429 (N_14429,N_14269,N_14320);
nand U14430 (N_14430,N_14317,N_14332);
xnor U14431 (N_14431,N_14303,N_14253);
or U14432 (N_14432,N_14193,N_14146);
nand U14433 (N_14433,N_14389,N_14158);
xor U14434 (N_14434,N_14174,N_14226);
nand U14435 (N_14435,N_14111,N_14390);
xnor U14436 (N_14436,N_14283,N_14155);
nand U14437 (N_14437,N_14113,N_14361);
nor U14438 (N_14438,N_14278,N_14354);
nand U14439 (N_14439,N_14360,N_14234);
xnor U14440 (N_14440,N_14179,N_14104);
or U14441 (N_14441,N_14244,N_14188);
xnor U14442 (N_14442,N_14135,N_14279);
or U14443 (N_14443,N_14271,N_14250);
xor U14444 (N_14444,N_14212,N_14310);
xnor U14445 (N_14445,N_14379,N_14241);
and U14446 (N_14446,N_14255,N_14210);
xor U14447 (N_14447,N_14191,N_14119);
and U14448 (N_14448,N_14236,N_14308);
and U14449 (N_14449,N_14154,N_14329);
nor U14450 (N_14450,N_14282,N_14275);
or U14451 (N_14451,N_14393,N_14259);
and U14452 (N_14452,N_14160,N_14319);
nand U14453 (N_14453,N_14126,N_14187);
nor U14454 (N_14454,N_14114,N_14112);
nor U14455 (N_14455,N_14331,N_14371);
nand U14456 (N_14456,N_14321,N_14208);
nand U14457 (N_14457,N_14385,N_14254);
xor U14458 (N_14458,N_14298,N_14138);
xnor U14459 (N_14459,N_14281,N_14288);
or U14460 (N_14460,N_14252,N_14339);
and U14461 (N_14461,N_14350,N_14386);
nand U14462 (N_14462,N_14195,N_14238);
nor U14463 (N_14463,N_14276,N_14384);
nand U14464 (N_14464,N_14318,N_14197);
nand U14465 (N_14465,N_14273,N_14219);
and U14466 (N_14466,N_14108,N_14216);
nor U14467 (N_14467,N_14251,N_14233);
and U14468 (N_14468,N_14312,N_14399);
nor U14469 (N_14469,N_14120,N_14277);
nand U14470 (N_14470,N_14133,N_14170);
and U14471 (N_14471,N_14125,N_14237);
nor U14472 (N_14472,N_14145,N_14101);
nand U14473 (N_14473,N_14185,N_14299);
and U14474 (N_14474,N_14220,N_14180);
and U14475 (N_14475,N_14313,N_14204);
or U14476 (N_14476,N_14184,N_14394);
or U14477 (N_14477,N_14148,N_14194);
nand U14478 (N_14478,N_14365,N_14257);
nand U14479 (N_14479,N_14338,N_14245);
or U14480 (N_14480,N_14190,N_14266);
or U14481 (N_14481,N_14364,N_14351);
nor U14482 (N_14482,N_14356,N_14366);
and U14483 (N_14483,N_14300,N_14326);
or U14484 (N_14484,N_14340,N_14213);
nand U14485 (N_14485,N_14382,N_14243);
nor U14486 (N_14486,N_14358,N_14240);
xnor U14487 (N_14487,N_14156,N_14100);
nor U14488 (N_14488,N_14392,N_14374);
nor U14489 (N_14489,N_14181,N_14344);
and U14490 (N_14490,N_14369,N_14224);
and U14491 (N_14491,N_14398,N_14167);
nand U14492 (N_14492,N_14166,N_14302);
xor U14493 (N_14493,N_14391,N_14118);
xnor U14494 (N_14494,N_14109,N_14373);
and U14495 (N_14495,N_14324,N_14173);
xnor U14496 (N_14496,N_14268,N_14262);
and U14497 (N_14497,N_14355,N_14345);
xnor U14498 (N_14498,N_14272,N_14153);
and U14499 (N_14499,N_14172,N_14140);
nor U14500 (N_14500,N_14129,N_14230);
nand U14501 (N_14501,N_14103,N_14284);
nor U14502 (N_14502,N_14161,N_14336);
or U14503 (N_14503,N_14203,N_14292);
and U14504 (N_14504,N_14200,N_14260);
xor U14505 (N_14505,N_14325,N_14265);
nand U14506 (N_14506,N_14296,N_14214);
nand U14507 (N_14507,N_14176,N_14274);
or U14508 (N_14508,N_14205,N_14183);
and U14509 (N_14509,N_14175,N_14267);
and U14510 (N_14510,N_14309,N_14388);
or U14511 (N_14511,N_14395,N_14285);
or U14512 (N_14512,N_14333,N_14348);
or U14513 (N_14513,N_14297,N_14352);
xnor U14514 (N_14514,N_14372,N_14115);
or U14515 (N_14515,N_14359,N_14201);
and U14516 (N_14516,N_14305,N_14168);
xor U14517 (N_14517,N_14106,N_14334);
xor U14518 (N_14518,N_14346,N_14192);
xor U14519 (N_14519,N_14165,N_14132);
xor U14520 (N_14520,N_14248,N_14301);
or U14521 (N_14521,N_14247,N_14218);
nand U14522 (N_14522,N_14362,N_14217);
and U14523 (N_14523,N_14264,N_14295);
nand U14524 (N_14524,N_14211,N_14381);
xnor U14525 (N_14525,N_14159,N_14144);
xor U14526 (N_14526,N_14207,N_14235);
or U14527 (N_14527,N_14270,N_14178);
xnor U14528 (N_14528,N_14327,N_14225);
nor U14529 (N_14529,N_14378,N_14322);
and U14530 (N_14530,N_14290,N_14152);
or U14531 (N_14531,N_14157,N_14280);
xor U14532 (N_14532,N_14105,N_14110);
xnor U14533 (N_14533,N_14353,N_14227);
nor U14534 (N_14534,N_14249,N_14287);
nand U14535 (N_14535,N_14198,N_14221);
nor U14536 (N_14536,N_14123,N_14316);
nand U14537 (N_14537,N_14370,N_14136);
nand U14538 (N_14538,N_14291,N_14223);
and U14539 (N_14539,N_14229,N_14164);
and U14540 (N_14540,N_14343,N_14215);
xor U14541 (N_14541,N_14387,N_14228);
nor U14542 (N_14542,N_14189,N_14163);
nor U14543 (N_14543,N_14162,N_14231);
nand U14544 (N_14544,N_14342,N_14330);
xor U14545 (N_14545,N_14335,N_14396);
and U14546 (N_14546,N_14323,N_14286);
nor U14547 (N_14547,N_14315,N_14232);
or U14548 (N_14548,N_14375,N_14169);
and U14549 (N_14549,N_14107,N_14127);
or U14550 (N_14550,N_14397,N_14124);
or U14551 (N_14551,N_14125,N_14216);
and U14552 (N_14552,N_14125,N_14374);
or U14553 (N_14553,N_14312,N_14368);
nand U14554 (N_14554,N_14136,N_14110);
nor U14555 (N_14555,N_14209,N_14223);
and U14556 (N_14556,N_14276,N_14103);
xor U14557 (N_14557,N_14140,N_14320);
or U14558 (N_14558,N_14214,N_14221);
xnor U14559 (N_14559,N_14142,N_14216);
or U14560 (N_14560,N_14352,N_14244);
nor U14561 (N_14561,N_14117,N_14136);
and U14562 (N_14562,N_14181,N_14114);
and U14563 (N_14563,N_14142,N_14111);
and U14564 (N_14564,N_14364,N_14321);
and U14565 (N_14565,N_14195,N_14387);
and U14566 (N_14566,N_14263,N_14363);
xor U14567 (N_14567,N_14104,N_14270);
nor U14568 (N_14568,N_14383,N_14323);
nor U14569 (N_14569,N_14390,N_14332);
nand U14570 (N_14570,N_14188,N_14237);
nand U14571 (N_14571,N_14111,N_14100);
and U14572 (N_14572,N_14358,N_14293);
nor U14573 (N_14573,N_14357,N_14364);
nand U14574 (N_14574,N_14249,N_14118);
and U14575 (N_14575,N_14379,N_14274);
xnor U14576 (N_14576,N_14273,N_14368);
nand U14577 (N_14577,N_14127,N_14133);
nor U14578 (N_14578,N_14303,N_14111);
or U14579 (N_14579,N_14244,N_14376);
or U14580 (N_14580,N_14254,N_14102);
and U14581 (N_14581,N_14125,N_14256);
or U14582 (N_14582,N_14269,N_14361);
or U14583 (N_14583,N_14386,N_14293);
nor U14584 (N_14584,N_14159,N_14292);
and U14585 (N_14585,N_14297,N_14192);
nor U14586 (N_14586,N_14384,N_14234);
and U14587 (N_14587,N_14205,N_14236);
or U14588 (N_14588,N_14325,N_14235);
nor U14589 (N_14589,N_14373,N_14288);
and U14590 (N_14590,N_14182,N_14258);
or U14591 (N_14591,N_14184,N_14215);
or U14592 (N_14592,N_14343,N_14398);
nor U14593 (N_14593,N_14334,N_14154);
xor U14594 (N_14594,N_14168,N_14105);
nand U14595 (N_14595,N_14209,N_14398);
and U14596 (N_14596,N_14300,N_14252);
or U14597 (N_14597,N_14183,N_14306);
xnor U14598 (N_14598,N_14337,N_14265);
nand U14599 (N_14599,N_14288,N_14396);
xnor U14600 (N_14600,N_14389,N_14297);
nor U14601 (N_14601,N_14254,N_14342);
nand U14602 (N_14602,N_14197,N_14356);
xor U14603 (N_14603,N_14178,N_14391);
or U14604 (N_14604,N_14386,N_14171);
and U14605 (N_14605,N_14195,N_14369);
nor U14606 (N_14606,N_14211,N_14137);
xor U14607 (N_14607,N_14190,N_14289);
xnor U14608 (N_14608,N_14269,N_14196);
nor U14609 (N_14609,N_14385,N_14376);
and U14610 (N_14610,N_14184,N_14313);
xor U14611 (N_14611,N_14132,N_14364);
or U14612 (N_14612,N_14217,N_14216);
or U14613 (N_14613,N_14348,N_14116);
or U14614 (N_14614,N_14381,N_14194);
xnor U14615 (N_14615,N_14364,N_14256);
nor U14616 (N_14616,N_14148,N_14189);
and U14617 (N_14617,N_14343,N_14282);
and U14618 (N_14618,N_14132,N_14184);
xor U14619 (N_14619,N_14201,N_14116);
and U14620 (N_14620,N_14166,N_14113);
nor U14621 (N_14621,N_14211,N_14221);
nor U14622 (N_14622,N_14256,N_14354);
or U14623 (N_14623,N_14169,N_14134);
or U14624 (N_14624,N_14305,N_14121);
nor U14625 (N_14625,N_14102,N_14214);
and U14626 (N_14626,N_14273,N_14331);
nand U14627 (N_14627,N_14294,N_14280);
or U14628 (N_14628,N_14202,N_14152);
and U14629 (N_14629,N_14108,N_14121);
nor U14630 (N_14630,N_14313,N_14308);
xor U14631 (N_14631,N_14328,N_14338);
nor U14632 (N_14632,N_14318,N_14121);
or U14633 (N_14633,N_14222,N_14309);
xor U14634 (N_14634,N_14340,N_14319);
nor U14635 (N_14635,N_14288,N_14152);
and U14636 (N_14636,N_14175,N_14221);
or U14637 (N_14637,N_14351,N_14350);
xnor U14638 (N_14638,N_14144,N_14239);
and U14639 (N_14639,N_14252,N_14109);
xor U14640 (N_14640,N_14244,N_14266);
nand U14641 (N_14641,N_14325,N_14121);
nor U14642 (N_14642,N_14377,N_14310);
nand U14643 (N_14643,N_14395,N_14177);
nor U14644 (N_14644,N_14299,N_14192);
nand U14645 (N_14645,N_14143,N_14297);
or U14646 (N_14646,N_14121,N_14352);
and U14647 (N_14647,N_14249,N_14187);
xnor U14648 (N_14648,N_14125,N_14196);
nor U14649 (N_14649,N_14282,N_14218);
and U14650 (N_14650,N_14237,N_14273);
and U14651 (N_14651,N_14212,N_14368);
or U14652 (N_14652,N_14241,N_14343);
xor U14653 (N_14653,N_14366,N_14211);
and U14654 (N_14654,N_14259,N_14206);
xor U14655 (N_14655,N_14255,N_14382);
nand U14656 (N_14656,N_14345,N_14148);
nor U14657 (N_14657,N_14367,N_14181);
nand U14658 (N_14658,N_14390,N_14396);
or U14659 (N_14659,N_14264,N_14253);
or U14660 (N_14660,N_14229,N_14269);
nor U14661 (N_14661,N_14183,N_14226);
and U14662 (N_14662,N_14207,N_14115);
or U14663 (N_14663,N_14380,N_14351);
xnor U14664 (N_14664,N_14248,N_14170);
nor U14665 (N_14665,N_14273,N_14395);
nor U14666 (N_14666,N_14313,N_14396);
or U14667 (N_14667,N_14148,N_14169);
nand U14668 (N_14668,N_14174,N_14117);
nand U14669 (N_14669,N_14101,N_14381);
and U14670 (N_14670,N_14341,N_14285);
xnor U14671 (N_14671,N_14342,N_14314);
or U14672 (N_14672,N_14111,N_14289);
and U14673 (N_14673,N_14327,N_14318);
or U14674 (N_14674,N_14165,N_14234);
xor U14675 (N_14675,N_14186,N_14272);
xnor U14676 (N_14676,N_14143,N_14137);
nor U14677 (N_14677,N_14328,N_14245);
or U14678 (N_14678,N_14314,N_14191);
and U14679 (N_14679,N_14319,N_14142);
or U14680 (N_14680,N_14312,N_14356);
and U14681 (N_14681,N_14188,N_14229);
nand U14682 (N_14682,N_14386,N_14375);
or U14683 (N_14683,N_14207,N_14203);
nand U14684 (N_14684,N_14217,N_14214);
and U14685 (N_14685,N_14275,N_14292);
nor U14686 (N_14686,N_14391,N_14184);
nand U14687 (N_14687,N_14153,N_14315);
nand U14688 (N_14688,N_14203,N_14142);
and U14689 (N_14689,N_14394,N_14132);
and U14690 (N_14690,N_14279,N_14369);
nand U14691 (N_14691,N_14197,N_14237);
nand U14692 (N_14692,N_14275,N_14375);
and U14693 (N_14693,N_14188,N_14203);
xnor U14694 (N_14694,N_14142,N_14133);
and U14695 (N_14695,N_14216,N_14145);
nand U14696 (N_14696,N_14364,N_14253);
nand U14697 (N_14697,N_14181,N_14152);
and U14698 (N_14698,N_14315,N_14148);
xnor U14699 (N_14699,N_14209,N_14292);
and U14700 (N_14700,N_14690,N_14592);
nand U14701 (N_14701,N_14568,N_14478);
nor U14702 (N_14702,N_14523,N_14441);
nor U14703 (N_14703,N_14404,N_14554);
nor U14704 (N_14704,N_14530,N_14677);
and U14705 (N_14705,N_14503,N_14505);
xnor U14706 (N_14706,N_14442,N_14546);
xnor U14707 (N_14707,N_14619,N_14431);
xnor U14708 (N_14708,N_14580,N_14430);
or U14709 (N_14709,N_14466,N_14538);
xnor U14710 (N_14710,N_14417,N_14635);
nand U14711 (N_14711,N_14632,N_14591);
or U14712 (N_14712,N_14514,N_14612);
nor U14713 (N_14713,N_14551,N_14680);
xor U14714 (N_14714,N_14518,N_14569);
xor U14715 (N_14715,N_14520,N_14429);
nand U14716 (N_14716,N_14552,N_14547);
and U14717 (N_14717,N_14408,N_14698);
nor U14718 (N_14718,N_14402,N_14685);
nor U14719 (N_14719,N_14631,N_14443);
or U14720 (N_14720,N_14629,N_14573);
or U14721 (N_14721,N_14474,N_14473);
nor U14722 (N_14722,N_14485,N_14432);
or U14723 (N_14723,N_14484,N_14601);
and U14724 (N_14724,N_14571,N_14579);
nor U14725 (N_14725,N_14486,N_14658);
xnor U14726 (N_14726,N_14557,N_14684);
and U14727 (N_14727,N_14438,N_14564);
and U14728 (N_14728,N_14614,N_14488);
and U14729 (N_14729,N_14515,N_14605);
nand U14730 (N_14730,N_14433,N_14403);
and U14731 (N_14731,N_14609,N_14480);
xnor U14732 (N_14732,N_14454,N_14511);
or U14733 (N_14733,N_14687,N_14559);
xor U14734 (N_14734,N_14625,N_14418);
and U14735 (N_14735,N_14683,N_14427);
nor U14736 (N_14736,N_14611,N_14587);
nor U14737 (N_14737,N_14641,N_14451);
nand U14738 (N_14738,N_14675,N_14560);
and U14739 (N_14739,N_14562,N_14494);
nor U14740 (N_14740,N_14411,N_14472);
xor U14741 (N_14741,N_14479,N_14495);
nor U14742 (N_14742,N_14656,N_14682);
nor U14743 (N_14743,N_14665,N_14409);
nand U14744 (N_14744,N_14572,N_14540);
nand U14745 (N_14745,N_14651,N_14457);
or U14746 (N_14746,N_14654,N_14519);
or U14747 (N_14747,N_14648,N_14510);
or U14748 (N_14748,N_14553,N_14657);
or U14749 (N_14749,N_14597,N_14421);
nand U14750 (N_14750,N_14558,N_14467);
and U14751 (N_14751,N_14414,N_14444);
xnor U14752 (N_14752,N_14542,N_14585);
xnor U14753 (N_14753,N_14616,N_14477);
xnor U14754 (N_14754,N_14529,N_14499);
xnor U14755 (N_14755,N_14536,N_14561);
or U14756 (N_14756,N_14650,N_14633);
xnor U14757 (N_14757,N_14598,N_14642);
nand U14758 (N_14758,N_14541,N_14527);
nor U14759 (N_14759,N_14671,N_14608);
nor U14760 (N_14760,N_14679,N_14681);
xnor U14761 (N_14761,N_14645,N_14539);
nor U14762 (N_14762,N_14673,N_14575);
and U14763 (N_14763,N_14487,N_14637);
nor U14764 (N_14764,N_14647,N_14581);
nor U14765 (N_14765,N_14506,N_14513);
nor U14766 (N_14766,N_14458,N_14674);
or U14767 (N_14767,N_14618,N_14653);
and U14768 (N_14768,N_14610,N_14422);
nor U14769 (N_14769,N_14576,N_14463);
and U14770 (N_14770,N_14624,N_14525);
or U14771 (N_14771,N_14535,N_14695);
or U14772 (N_14772,N_14584,N_14504);
xnor U14773 (N_14773,N_14588,N_14662);
nand U14774 (N_14774,N_14567,N_14623);
xor U14775 (N_14775,N_14668,N_14602);
nand U14776 (N_14776,N_14507,N_14470);
xnor U14777 (N_14777,N_14666,N_14595);
xnor U14778 (N_14778,N_14522,N_14626);
nand U14779 (N_14779,N_14652,N_14455);
nor U14780 (N_14780,N_14692,N_14694);
nand U14781 (N_14781,N_14672,N_14468);
nand U14782 (N_14782,N_14622,N_14604);
nor U14783 (N_14783,N_14528,N_14563);
and U14784 (N_14784,N_14615,N_14496);
or U14785 (N_14785,N_14440,N_14549);
or U14786 (N_14786,N_14594,N_14586);
and U14787 (N_14787,N_14423,N_14583);
nor U14788 (N_14788,N_14621,N_14426);
and U14789 (N_14789,N_14508,N_14533);
nor U14790 (N_14790,N_14667,N_14460);
nor U14791 (N_14791,N_14696,N_14659);
xor U14792 (N_14792,N_14490,N_14532);
nand U14793 (N_14793,N_14676,N_14456);
nand U14794 (N_14794,N_14464,N_14548);
nand U14795 (N_14795,N_14663,N_14406);
or U14796 (N_14796,N_14512,N_14447);
or U14797 (N_14797,N_14664,N_14450);
or U14798 (N_14798,N_14661,N_14498);
xor U14799 (N_14799,N_14410,N_14446);
nor U14800 (N_14800,N_14646,N_14517);
nand U14801 (N_14801,N_14544,N_14521);
nand U14802 (N_14802,N_14401,N_14531);
and U14803 (N_14803,N_14688,N_14630);
and U14804 (N_14804,N_14415,N_14475);
nand U14805 (N_14805,N_14678,N_14481);
or U14806 (N_14806,N_14634,N_14627);
nor U14807 (N_14807,N_14639,N_14649);
or U14808 (N_14808,N_14492,N_14577);
and U14809 (N_14809,N_14574,N_14603);
or U14810 (N_14810,N_14425,N_14465);
and U14811 (N_14811,N_14669,N_14407);
nor U14812 (N_14812,N_14636,N_14400);
nand U14813 (N_14813,N_14660,N_14471);
nand U14814 (N_14814,N_14524,N_14589);
xor U14815 (N_14815,N_14493,N_14545);
nand U14816 (N_14816,N_14405,N_14643);
xor U14817 (N_14817,N_14491,N_14462);
or U14818 (N_14818,N_14578,N_14550);
nand U14819 (N_14819,N_14502,N_14693);
or U14820 (N_14820,N_14419,N_14606);
and U14821 (N_14821,N_14435,N_14644);
xor U14822 (N_14822,N_14501,N_14691);
and U14823 (N_14823,N_14469,N_14453);
nand U14824 (N_14824,N_14434,N_14413);
and U14825 (N_14825,N_14424,N_14617);
nand U14826 (N_14826,N_14613,N_14500);
and U14827 (N_14827,N_14482,N_14686);
xnor U14828 (N_14828,N_14593,N_14497);
xor U14829 (N_14829,N_14689,N_14590);
nand U14830 (N_14830,N_14670,N_14628);
nor U14831 (N_14831,N_14555,N_14452);
xnor U14832 (N_14832,N_14449,N_14599);
xor U14833 (N_14833,N_14556,N_14420);
nor U14834 (N_14834,N_14476,N_14543);
nor U14835 (N_14835,N_14461,N_14582);
nor U14836 (N_14836,N_14439,N_14697);
or U14837 (N_14837,N_14445,N_14428);
nand U14838 (N_14838,N_14570,N_14483);
and U14839 (N_14839,N_14516,N_14600);
or U14840 (N_14840,N_14640,N_14437);
nor U14841 (N_14841,N_14459,N_14565);
nor U14842 (N_14842,N_14638,N_14448);
and U14843 (N_14843,N_14537,N_14489);
xnor U14844 (N_14844,N_14607,N_14655);
nor U14845 (N_14845,N_14534,N_14526);
and U14846 (N_14846,N_14620,N_14566);
or U14847 (N_14847,N_14509,N_14436);
xnor U14848 (N_14848,N_14412,N_14416);
and U14849 (N_14849,N_14596,N_14699);
xnor U14850 (N_14850,N_14559,N_14446);
xor U14851 (N_14851,N_14589,N_14635);
nor U14852 (N_14852,N_14567,N_14698);
nor U14853 (N_14853,N_14532,N_14400);
nand U14854 (N_14854,N_14583,N_14424);
nand U14855 (N_14855,N_14625,N_14499);
or U14856 (N_14856,N_14614,N_14586);
or U14857 (N_14857,N_14679,N_14593);
and U14858 (N_14858,N_14546,N_14475);
nand U14859 (N_14859,N_14535,N_14538);
xor U14860 (N_14860,N_14504,N_14426);
nor U14861 (N_14861,N_14605,N_14459);
and U14862 (N_14862,N_14473,N_14441);
nor U14863 (N_14863,N_14475,N_14416);
nand U14864 (N_14864,N_14434,N_14420);
nand U14865 (N_14865,N_14457,N_14624);
or U14866 (N_14866,N_14583,N_14655);
or U14867 (N_14867,N_14508,N_14472);
nor U14868 (N_14868,N_14530,N_14678);
xor U14869 (N_14869,N_14645,N_14576);
nand U14870 (N_14870,N_14516,N_14514);
xnor U14871 (N_14871,N_14683,N_14512);
or U14872 (N_14872,N_14440,N_14646);
and U14873 (N_14873,N_14515,N_14610);
nor U14874 (N_14874,N_14412,N_14503);
nand U14875 (N_14875,N_14458,N_14523);
or U14876 (N_14876,N_14499,N_14623);
nand U14877 (N_14877,N_14457,N_14596);
xor U14878 (N_14878,N_14609,N_14431);
xnor U14879 (N_14879,N_14573,N_14692);
and U14880 (N_14880,N_14401,N_14507);
and U14881 (N_14881,N_14421,N_14610);
xnor U14882 (N_14882,N_14408,N_14594);
nor U14883 (N_14883,N_14674,N_14550);
nand U14884 (N_14884,N_14514,N_14691);
or U14885 (N_14885,N_14654,N_14694);
xnor U14886 (N_14886,N_14468,N_14462);
nor U14887 (N_14887,N_14549,N_14678);
nor U14888 (N_14888,N_14423,N_14489);
or U14889 (N_14889,N_14518,N_14492);
nor U14890 (N_14890,N_14585,N_14517);
or U14891 (N_14891,N_14669,N_14474);
xor U14892 (N_14892,N_14601,N_14543);
or U14893 (N_14893,N_14602,N_14598);
and U14894 (N_14894,N_14591,N_14634);
nor U14895 (N_14895,N_14546,N_14654);
nor U14896 (N_14896,N_14411,N_14484);
or U14897 (N_14897,N_14425,N_14554);
and U14898 (N_14898,N_14587,N_14497);
or U14899 (N_14899,N_14545,N_14632);
xor U14900 (N_14900,N_14655,N_14684);
or U14901 (N_14901,N_14412,N_14651);
xor U14902 (N_14902,N_14549,N_14557);
and U14903 (N_14903,N_14699,N_14516);
or U14904 (N_14904,N_14625,N_14471);
and U14905 (N_14905,N_14440,N_14483);
nand U14906 (N_14906,N_14580,N_14435);
nand U14907 (N_14907,N_14525,N_14500);
xor U14908 (N_14908,N_14575,N_14428);
and U14909 (N_14909,N_14590,N_14410);
or U14910 (N_14910,N_14523,N_14583);
and U14911 (N_14911,N_14582,N_14573);
xor U14912 (N_14912,N_14491,N_14561);
nand U14913 (N_14913,N_14404,N_14629);
and U14914 (N_14914,N_14591,N_14668);
xor U14915 (N_14915,N_14645,N_14642);
or U14916 (N_14916,N_14691,N_14566);
and U14917 (N_14917,N_14508,N_14566);
or U14918 (N_14918,N_14457,N_14446);
xnor U14919 (N_14919,N_14698,N_14552);
or U14920 (N_14920,N_14567,N_14681);
nor U14921 (N_14921,N_14413,N_14487);
and U14922 (N_14922,N_14448,N_14590);
nor U14923 (N_14923,N_14620,N_14545);
nor U14924 (N_14924,N_14458,N_14406);
xor U14925 (N_14925,N_14591,N_14471);
and U14926 (N_14926,N_14499,N_14693);
nand U14927 (N_14927,N_14651,N_14575);
or U14928 (N_14928,N_14464,N_14513);
nor U14929 (N_14929,N_14477,N_14615);
or U14930 (N_14930,N_14445,N_14683);
and U14931 (N_14931,N_14522,N_14478);
nor U14932 (N_14932,N_14600,N_14551);
and U14933 (N_14933,N_14541,N_14540);
xnor U14934 (N_14934,N_14430,N_14542);
nand U14935 (N_14935,N_14634,N_14597);
xor U14936 (N_14936,N_14603,N_14695);
nor U14937 (N_14937,N_14611,N_14618);
xor U14938 (N_14938,N_14503,N_14502);
and U14939 (N_14939,N_14679,N_14467);
nor U14940 (N_14940,N_14576,N_14569);
and U14941 (N_14941,N_14509,N_14639);
nand U14942 (N_14942,N_14473,N_14518);
and U14943 (N_14943,N_14403,N_14425);
nand U14944 (N_14944,N_14624,N_14406);
xor U14945 (N_14945,N_14509,N_14562);
nand U14946 (N_14946,N_14474,N_14572);
nand U14947 (N_14947,N_14532,N_14421);
and U14948 (N_14948,N_14485,N_14539);
or U14949 (N_14949,N_14618,N_14507);
nor U14950 (N_14950,N_14467,N_14635);
or U14951 (N_14951,N_14508,N_14423);
nand U14952 (N_14952,N_14559,N_14574);
or U14953 (N_14953,N_14472,N_14652);
nor U14954 (N_14954,N_14686,N_14447);
and U14955 (N_14955,N_14521,N_14529);
xor U14956 (N_14956,N_14576,N_14617);
and U14957 (N_14957,N_14590,N_14419);
xor U14958 (N_14958,N_14439,N_14649);
nand U14959 (N_14959,N_14664,N_14672);
xnor U14960 (N_14960,N_14689,N_14450);
xor U14961 (N_14961,N_14480,N_14569);
or U14962 (N_14962,N_14668,N_14401);
and U14963 (N_14963,N_14666,N_14579);
and U14964 (N_14964,N_14699,N_14534);
and U14965 (N_14965,N_14673,N_14419);
nand U14966 (N_14966,N_14644,N_14412);
and U14967 (N_14967,N_14692,N_14623);
nor U14968 (N_14968,N_14400,N_14639);
and U14969 (N_14969,N_14656,N_14606);
nand U14970 (N_14970,N_14425,N_14693);
or U14971 (N_14971,N_14494,N_14521);
nand U14972 (N_14972,N_14632,N_14526);
nor U14973 (N_14973,N_14659,N_14614);
and U14974 (N_14974,N_14559,N_14680);
and U14975 (N_14975,N_14490,N_14458);
or U14976 (N_14976,N_14620,N_14651);
or U14977 (N_14977,N_14474,N_14699);
nand U14978 (N_14978,N_14582,N_14615);
nand U14979 (N_14979,N_14526,N_14538);
nand U14980 (N_14980,N_14550,N_14457);
xor U14981 (N_14981,N_14608,N_14596);
and U14982 (N_14982,N_14617,N_14513);
or U14983 (N_14983,N_14447,N_14565);
nand U14984 (N_14984,N_14636,N_14678);
and U14985 (N_14985,N_14433,N_14543);
xor U14986 (N_14986,N_14662,N_14436);
and U14987 (N_14987,N_14684,N_14682);
and U14988 (N_14988,N_14632,N_14441);
and U14989 (N_14989,N_14498,N_14621);
xor U14990 (N_14990,N_14687,N_14689);
nor U14991 (N_14991,N_14674,N_14677);
or U14992 (N_14992,N_14635,N_14435);
nand U14993 (N_14993,N_14539,N_14599);
xnor U14994 (N_14994,N_14420,N_14422);
and U14995 (N_14995,N_14620,N_14526);
xnor U14996 (N_14996,N_14428,N_14464);
xnor U14997 (N_14997,N_14637,N_14687);
nand U14998 (N_14998,N_14630,N_14431);
and U14999 (N_14999,N_14624,N_14436);
or UO_0 (O_0,N_14794,N_14904);
or UO_1 (O_1,N_14991,N_14784);
xnor UO_2 (O_2,N_14785,N_14842);
nor UO_3 (O_3,N_14949,N_14830);
nor UO_4 (O_4,N_14778,N_14929);
and UO_5 (O_5,N_14901,N_14770);
and UO_6 (O_6,N_14839,N_14944);
and UO_7 (O_7,N_14907,N_14872);
nor UO_8 (O_8,N_14865,N_14945);
xnor UO_9 (O_9,N_14918,N_14985);
nor UO_10 (O_10,N_14933,N_14957);
or UO_11 (O_11,N_14786,N_14942);
or UO_12 (O_12,N_14810,N_14808);
nor UO_13 (O_13,N_14740,N_14832);
nor UO_14 (O_14,N_14837,N_14887);
xnor UO_15 (O_15,N_14749,N_14713);
nand UO_16 (O_16,N_14843,N_14745);
nor UO_17 (O_17,N_14803,N_14868);
nand UO_18 (O_18,N_14722,N_14921);
or UO_19 (O_19,N_14972,N_14773);
xnor UO_20 (O_20,N_14923,N_14903);
xor UO_21 (O_21,N_14976,N_14978);
and UO_22 (O_22,N_14968,N_14964);
nor UO_23 (O_23,N_14875,N_14847);
or UO_24 (O_24,N_14757,N_14727);
nand UO_25 (O_25,N_14734,N_14767);
nor UO_26 (O_26,N_14946,N_14704);
xor UO_27 (O_27,N_14896,N_14971);
and UO_28 (O_28,N_14851,N_14920);
nor UO_29 (O_29,N_14791,N_14826);
xnor UO_30 (O_30,N_14880,N_14718);
and UO_31 (O_31,N_14715,N_14774);
nor UO_32 (O_32,N_14965,N_14841);
xnor UO_33 (O_33,N_14742,N_14914);
nand UO_34 (O_34,N_14783,N_14838);
nor UO_35 (O_35,N_14994,N_14899);
nor UO_36 (O_36,N_14712,N_14762);
nor UO_37 (O_37,N_14723,N_14828);
xnor UO_38 (O_38,N_14739,N_14995);
xor UO_39 (O_39,N_14768,N_14780);
or UO_40 (O_40,N_14706,N_14754);
nor UO_41 (O_41,N_14703,N_14943);
xor UO_42 (O_42,N_14858,N_14882);
and UO_43 (O_43,N_14714,N_14719);
nand UO_44 (O_44,N_14962,N_14931);
and UO_45 (O_45,N_14910,N_14848);
nor UO_46 (O_46,N_14743,N_14937);
xnor UO_47 (O_47,N_14981,N_14788);
nor UO_48 (O_48,N_14857,N_14974);
xor UO_49 (O_49,N_14824,N_14967);
xor UO_50 (O_50,N_14970,N_14818);
nand UO_51 (O_51,N_14833,N_14732);
and UO_52 (O_52,N_14735,N_14900);
nand UO_53 (O_53,N_14758,N_14908);
or UO_54 (O_54,N_14725,N_14853);
or UO_55 (O_55,N_14804,N_14998);
xnor UO_56 (O_56,N_14856,N_14702);
or UO_57 (O_57,N_14731,N_14936);
xnor UO_58 (O_58,N_14850,N_14924);
or UO_59 (O_59,N_14956,N_14849);
nor UO_60 (O_60,N_14834,N_14797);
or UO_61 (O_61,N_14812,N_14996);
or UO_62 (O_62,N_14835,N_14776);
or UO_63 (O_63,N_14790,N_14930);
nand UO_64 (O_64,N_14869,N_14885);
xor UO_65 (O_65,N_14870,N_14966);
nand UO_66 (O_66,N_14883,N_14905);
or UO_67 (O_67,N_14779,N_14855);
xnor UO_68 (O_68,N_14759,N_14892);
or UO_69 (O_69,N_14819,N_14806);
nand UO_70 (O_70,N_14969,N_14898);
nor UO_71 (O_71,N_14720,N_14982);
nor UO_72 (O_72,N_14795,N_14932);
xnor UO_73 (O_73,N_14705,N_14912);
or UO_74 (O_74,N_14915,N_14955);
or UO_75 (O_75,N_14809,N_14755);
nor UO_76 (O_76,N_14793,N_14708);
or UO_77 (O_77,N_14960,N_14890);
and UO_78 (O_78,N_14893,N_14716);
or UO_79 (O_79,N_14825,N_14983);
nand UO_80 (O_80,N_14884,N_14707);
nand UO_81 (O_81,N_14800,N_14878);
nor UO_82 (O_82,N_14894,N_14730);
nor UO_83 (O_83,N_14895,N_14864);
nand UO_84 (O_84,N_14802,N_14928);
nor UO_85 (O_85,N_14846,N_14750);
or UO_86 (O_86,N_14874,N_14840);
or UO_87 (O_87,N_14744,N_14807);
or UO_88 (O_88,N_14902,N_14726);
xnor UO_89 (O_89,N_14852,N_14909);
nor UO_90 (O_90,N_14709,N_14792);
and UO_91 (O_91,N_14888,N_14741);
xor UO_92 (O_92,N_14879,N_14775);
nand UO_93 (O_93,N_14782,N_14764);
nand UO_94 (O_94,N_14961,N_14777);
nand UO_95 (O_95,N_14861,N_14753);
nand UO_96 (O_96,N_14940,N_14737);
xnor UO_97 (O_97,N_14728,N_14859);
and UO_98 (O_98,N_14987,N_14823);
and UO_99 (O_99,N_14701,N_14766);
xor UO_100 (O_100,N_14950,N_14700);
nand UO_101 (O_101,N_14934,N_14799);
nor UO_102 (O_102,N_14756,N_14917);
nor UO_103 (O_103,N_14787,N_14980);
nor UO_104 (O_104,N_14746,N_14862);
nand UO_105 (O_105,N_14772,N_14729);
nor UO_106 (O_106,N_14736,N_14801);
xnor UO_107 (O_107,N_14916,N_14760);
or UO_108 (O_108,N_14999,N_14889);
or UO_109 (O_109,N_14724,N_14710);
xnor UO_110 (O_110,N_14984,N_14947);
or UO_111 (O_111,N_14711,N_14765);
nand UO_112 (O_112,N_14751,N_14881);
or UO_113 (O_113,N_14988,N_14963);
nand UO_114 (O_114,N_14836,N_14871);
xnor UO_115 (O_115,N_14860,N_14913);
xor UO_116 (O_116,N_14977,N_14876);
nand UO_117 (O_117,N_14844,N_14886);
or UO_118 (O_118,N_14829,N_14939);
and UO_119 (O_119,N_14789,N_14721);
nand UO_120 (O_120,N_14990,N_14816);
nand UO_121 (O_121,N_14781,N_14717);
nor UO_122 (O_122,N_14821,N_14992);
or UO_123 (O_123,N_14752,N_14733);
nand UO_124 (O_124,N_14891,N_14951);
or UO_125 (O_125,N_14938,N_14769);
nand UO_126 (O_126,N_14845,N_14958);
xor UO_127 (O_127,N_14747,N_14997);
xor UO_128 (O_128,N_14827,N_14817);
and UO_129 (O_129,N_14927,N_14897);
xnor UO_130 (O_130,N_14863,N_14796);
nand UO_131 (O_131,N_14738,N_14805);
or UO_132 (O_132,N_14948,N_14867);
nor UO_133 (O_133,N_14926,N_14831);
xor UO_134 (O_134,N_14811,N_14935);
xor UO_135 (O_135,N_14815,N_14906);
xor UO_136 (O_136,N_14813,N_14986);
and UO_137 (O_137,N_14761,N_14748);
and UO_138 (O_138,N_14854,N_14925);
nor UO_139 (O_139,N_14822,N_14771);
or UO_140 (O_140,N_14954,N_14911);
nor UO_141 (O_141,N_14959,N_14989);
and UO_142 (O_142,N_14798,N_14922);
and UO_143 (O_143,N_14973,N_14952);
nand UO_144 (O_144,N_14763,N_14941);
nand UO_145 (O_145,N_14953,N_14919);
or UO_146 (O_146,N_14866,N_14993);
xnor UO_147 (O_147,N_14975,N_14820);
xor UO_148 (O_148,N_14979,N_14877);
or UO_149 (O_149,N_14873,N_14814);
xnor UO_150 (O_150,N_14787,N_14856);
nor UO_151 (O_151,N_14990,N_14919);
xnor UO_152 (O_152,N_14709,N_14895);
and UO_153 (O_153,N_14814,N_14917);
nand UO_154 (O_154,N_14853,N_14923);
nor UO_155 (O_155,N_14751,N_14801);
or UO_156 (O_156,N_14787,N_14741);
and UO_157 (O_157,N_14878,N_14872);
or UO_158 (O_158,N_14828,N_14824);
xnor UO_159 (O_159,N_14858,N_14876);
xor UO_160 (O_160,N_14850,N_14804);
nand UO_161 (O_161,N_14773,N_14803);
nor UO_162 (O_162,N_14856,N_14706);
nor UO_163 (O_163,N_14849,N_14753);
nand UO_164 (O_164,N_14996,N_14964);
nor UO_165 (O_165,N_14842,N_14915);
nand UO_166 (O_166,N_14882,N_14941);
or UO_167 (O_167,N_14741,N_14864);
nand UO_168 (O_168,N_14772,N_14853);
or UO_169 (O_169,N_14836,N_14854);
or UO_170 (O_170,N_14866,N_14877);
nor UO_171 (O_171,N_14820,N_14844);
xnor UO_172 (O_172,N_14887,N_14771);
nand UO_173 (O_173,N_14801,N_14877);
xor UO_174 (O_174,N_14841,N_14731);
xor UO_175 (O_175,N_14824,N_14814);
nand UO_176 (O_176,N_14851,N_14829);
and UO_177 (O_177,N_14964,N_14740);
nand UO_178 (O_178,N_14718,N_14900);
nor UO_179 (O_179,N_14901,N_14904);
and UO_180 (O_180,N_14888,N_14829);
nor UO_181 (O_181,N_14976,N_14871);
nand UO_182 (O_182,N_14839,N_14970);
nor UO_183 (O_183,N_14786,N_14851);
nor UO_184 (O_184,N_14953,N_14707);
xor UO_185 (O_185,N_14803,N_14897);
and UO_186 (O_186,N_14947,N_14872);
and UO_187 (O_187,N_14704,N_14738);
nor UO_188 (O_188,N_14794,N_14850);
xnor UO_189 (O_189,N_14957,N_14894);
and UO_190 (O_190,N_14850,N_14857);
and UO_191 (O_191,N_14892,N_14844);
or UO_192 (O_192,N_14875,N_14882);
or UO_193 (O_193,N_14899,N_14990);
and UO_194 (O_194,N_14778,N_14838);
nor UO_195 (O_195,N_14928,N_14896);
and UO_196 (O_196,N_14909,N_14932);
and UO_197 (O_197,N_14811,N_14768);
and UO_198 (O_198,N_14814,N_14733);
nand UO_199 (O_199,N_14832,N_14958);
or UO_200 (O_200,N_14888,N_14807);
nand UO_201 (O_201,N_14722,N_14746);
nor UO_202 (O_202,N_14830,N_14762);
and UO_203 (O_203,N_14812,N_14980);
xor UO_204 (O_204,N_14988,N_14785);
and UO_205 (O_205,N_14968,N_14886);
nand UO_206 (O_206,N_14913,N_14801);
or UO_207 (O_207,N_14906,N_14700);
nand UO_208 (O_208,N_14858,N_14783);
or UO_209 (O_209,N_14709,N_14887);
and UO_210 (O_210,N_14828,N_14877);
xor UO_211 (O_211,N_14730,N_14972);
nand UO_212 (O_212,N_14728,N_14775);
or UO_213 (O_213,N_14857,N_14953);
or UO_214 (O_214,N_14769,N_14904);
nor UO_215 (O_215,N_14984,N_14855);
nor UO_216 (O_216,N_14848,N_14806);
nand UO_217 (O_217,N_14975,N_14845);
xor UO_218 (O_218,N_14709,N_14950);
nor UO_219 (O_219,N_14957,N_14844);
nor UO_220 (O_220,N_14761,N_14724);
xor UO_221 (O_221,N_14958,N_14773);
nor UO_222 (O_222,N_14908,N_14833);
or UO_223 (O_223,N_14764,N_14744);
nor UO_224 (O_224,N_14708,N_14797);
xnor UO_225 (O_225,N_14853,N_14700);
nor UO_226 (O_226,N_14950,N_14778);
or UO_227 (O_227,N_14923,N_14763);
xnor UO_228 (O_228,N_14994,N_14762);
nand UO_229 (O_229,N_14877,N_14902);
nor UO_230 (O_230,N_14913,N_14823);
and UO_231 (O_231,N_14844,N_14958);
xnor UO_232 (O_232,N_14747,N_14938);
xor UO_233 (O_233,N_14769,N_14891);
and UO_234 (O_234,N_14898,N_14786);
xor UO_235 (O_235,N_14865,N_14762);
xnor UO_236 (O_236,N_14848,N_14722);
or UO_237 (O_237,N_14825,N_14896);
or UO_238 (O_238,N_14744,N_14852);
or UO_239 (O_239,N_14717,N_14986);
nor UO_240 (O_240,N_14700,N_14727);
nand UO_241 (O_241,N_14764,N_14924);
nor UO_242 (O_242,N_14869,N_14907);
or UO_243 (O_243,N_14829,N_14702);
nor UO_244 (O_244,N_14835,N_14725);
nand UO_245 (O_245,N_14755,N_14758);
nand UO_246 (O_246,N_14831,N_14973);
nor UO_247 (O_247,N_14934,N_14875);
or UO_248 (O_248,N_14755,N_14716);
or UO_249 (O_249,N_14898,N_14980);
and UO_250 (O_250,N_14881,N_14736);
and UO_251 (O_251,N_14970,N_14977);
xor UO_252 (O_252,N_14819,N_14784);
and UO_253 (O_253,N_14993,N_14777);
nor UO_254 (O_254,N_14809,N_14800);
or UO_255 (O_255,N_14976,N_14974);
and UO_256 (O_256,N_14806,N_14841);
nor UO_257 (O_257,N_14707,N_14758);
and UO_258 (O_258,N_14728,N_14997);
xor UO_259 (O_259,N_14971,N_14885);
and UO_260 (O_260,N_14977,N_14751);
xnor UO_261 (O_261,N_14881,N_14730);
and UO_262 (O_262,N_14808,N_14730);
nand UO_263 (O_263,N_14841,N_14884);
nand UO_264 (O_264,N_14878,N_14754);
and UO_265 (O_265,N_14775,N_14929);
or UO_266 (O_266,N_14779,N_14879);
xor UO_267 (O_267,N_14985,N_14884);
xnor UO_268 (O_268,N_14874,N_14797);
or UO_269 (O_269,N_14851,N_14718);
nor UO_270 (O_270,N_14855,N_14709);
nand UO_271 (O_271,N_14703,N_14817);
nand UO_272 (O_272,N_14814,N_14855);
or UO_273 (O_273,N_14707,N_14838);
or UO_274 (O_274,N_14933,N_14757);
and UO_275 (O_275,N_14986,N_14861);
nor UO_276 (O_276,N_14782,N_14836);
and UO_277 (O_277,N_14925,N_14903);
nor UO_278 (O_278,N_14824,N_14882);
nor UO_279 (O_279,N_14731,N_14736);
nand UO_280 (O_280,N_14885,N_14884);
and UO_281 (O_281,N_14994,N_14951);
nor UO_282 (O_282,N_14961,N_14864);
nand UO_283 (O_283,N_14800,N_14873);
and UO_284 (O_284,N_14992,N_14839);
and UO_285 (O_285,N_14846,N_14948);
xor UO_286 (O_286,N_14842,N_14980);
nor UO_287 (O_287,N_14973,N_14996);
and UO_288 (O_288,N_14906,N_14849);
nor UO_289 (O_289,N_14748,N_14700);
and UO_290 (O_290,N_14790,N_14779);
xor UO_291 (O_291,N_14779,N_14998);
and UO_292 (O_292,N_14984,N_14707);
nor UO_293 (O_293,N_14738,N_14815);
xnor UO_294 (O_294,N_14703,N_14954);
or UO_295 (O_295,N_14702,N_14954);
or UO_296 (O_296,N_14856,N_14878);
nor UO_297 (O_297,N_14919,N_14767);
xnor UO_298 (O_298,N_14792,N_14819);
or UO_299 (O_299,N_14889,N_14925);
nor UO_300 (O_300,N_14836,N_14896);
nor UO_301 (O_301,N_14903,N_14959);
or UO_302 (O_302,N_14929,N_14984);
and UO_303 (O_303,N_14939,N_14841);
and UO_304 (O_304,N_14849,N_14793);
nand UO_305 (O_305,N_14755,N_14985);
and UO_306 (O_306,N_14883,N_14802);
nand UO_307 (O_307,N_14857,N_14825);
nor UO_308 (O_308,N_14711,N_14967);
and UO_309 (O_309,N_14801,N_14995);
nand UO_310 (O_310,N_14841,N_14941);
xor UO_311 (O_311,N_14803,N_14887);
and UO_312 (O_312,N_14737,N_14872);
or UO_313 (O_313,N_14929,N_14821);
and UO_314 (O_314,N_14787,N_14885);
or UO_315 (O_315,N_14924,N_14704);
nand UO_316 (O_316,N_14703,N_14769);
or UO_317 (O_317,N_14895,N_14759);
or UO_318 (O_318,N_14753,N_14896);
nor UO_319 (O_319,N_14747,N_14791);
nand UO_320 (O_320,N_14851,N_14855);
and UO_321 (O_321,N_14852,N_14960);
and UO_322 (O_322,N_14912,N_14842);
and UO_323 (O_323,N_14960,N_14808);
nor UO_324 (O_324,N_14889,N_14929);
and UO_325 (O_325,N_14991,N_14864);
nor UO_326 (O_326,N_14928,N_14967);
xnor UO_327 (O_327,N_14952,N_14831);
nor UO_328 (O_328,N_14796,N_14968);
and UO_329 (O_329,N_14730,N_14979);
nor UO_330 (O_330,N_14976,N_14729);
nor UO_331 (O_331,N_14712,N_14731);
xor UO_332 (O_332,N_14703,N_14773);
and UO_333 (O_333,N_14781,N_14875);
or UO_334 (O_334,N_14964,N_14975);
xor UO_335 (O_335,N_14914,N_14768);
nand UO_336 (O_336,N_14736,N_14775);
and UO_337 (O_337,N_14991,N_14930);
nand UO_338 (O_338,N_14954,N_14982);
nor UO_339 (O_339,N_14790,N_14803);
or UO_340 (O_340,N_14856,N_14817);
xnor UO_341 (O_341,N_14822,N_14950);
and UO_342 (O_342,N_14846,N_14708);
and UO_343 (O_343,N_14730,N_14833);
nor UO_344 (O_344,N_14761,N_14958);
xor UO_345 (O_345,N_14820,N_14734);
or UO_346 (O_346,N_14736,N_14938);
xnor UO_347 (O_347,N_14906,N_14949);
or UO_348 (O_348,N_14901,N_14805);
nand UO_349 (O_349,N_14939,N_14867);
nand UO_350 (O_350,N_14754,N_14775);
xnor UO_351 (O_351,N_14888,N_14919);
nand UO_352 (O_352,N_14716,N_14837);
and UO_353 (O_353,N_14852,N_14849);
and UO_354 (O_354,N_14720,N_14793);
or UO_355 (O_355,N_14720,N_14755);
nand UO_356 (O_356,N_14867,N_14712);
or UO_357 (O_357,N_14980,N_14732);
xor UO_358 (O_358,N_14988,N_14815);
nand UO_359 (O_359,N_14777,N_14709);
nor UO_360 (O_360,N_14999,N_14794);
nor UO_361 (O_361,N_14879,N_14898);
xnor UO_362 (O_362,N_14703,N_14930);
nor UO_363 (O_363,N_14984,N_14761);
or UO_364 (O_364,N_14779,N_14701);
or UO_365 (O_365,N_14920,N_14836);
and UO_366 (O_366,N_14919,N_14896);
or UO_367 (O_367,N_14743,N_14730);
or UO_368 (O_368,N_14970,N_14821);
xnor UO_369 (O_369,N_14878,N_14901);
xnor UO_370 (O_370,N_14778,N_14897);
nand UO_371 (O_371,N_14893,N_14857);
nand UO_372 (O_372,N_14848,N_14751);
xnor UO_373 (O_373,N_14930,N_14980);
or UO_374 (O_374,N_14983,N_14832);
nand UO_375 (O_375,N_14987,N_14732);
or UO_376 (O_376,N_14923,N_14913);
nor UO_377 (O_377,N_14873,N_14780);
nor UO_378 (O_378,N_14768,N_14700);
nand UO_379 (O_379,N_14964,N_14957);
xnor UO_380 (O_380,N_14838,N_14989);
nand UO_381 (O_381,N_14766,N_14921);
nor UO_382 (O_382,N_14818,N_14788);
nand UO_383 (O_383,N_14866,N_14792);
and UO_384 (O_384,N_14878,N_14909);
nand UO_385 (O_385,N_14976,N_14883);
xor UO_386 (O_386,N_14923,N_14852);
nand UO_387 (O_387,N_14982,N_14876);
nor UO_388 (O_388,N_14946,N_14701);
or UO_389 (O_389,N_14845,N_14844);
xnor UO_390 (O_390,N_14956,N_14751);
or UO_391 (O_391,N_14880,N_14882);
nor UO_392 (O_392,N_14874,N_14748);
and UO_393 (O_393,N_14947,N_14988);
or UO_394 (O_394,N_14745,N_14766);
nand UO_395 (O_395,N_14764,N_14840);
nand UO_396 (O_396,N_14726,N_14747);
and UO_397 (O_397,N_14735,N_14743);
xor UO_398 (O_398,N_14865,N_14819);
and UO_399 (O_399,N_14821,N_14734);
nand UO_400 (O_400,N_14967,N_14924);
and UO_401 (O_401,N_14863,N_14790);
and UO_402 (O_402,N_14997,N_14940);
xnor UO_403 (O_403,N_14767,N_14886);
nand UO_404 (O_404,N_14787,N_14939);
xor UO_405 (O_405,N_14860,N_14962);
and UO_406 (O_406,N_14824,N_14889);
nor UO_407 (O_407,N_14768,N_14979);
and UO_408 (O_408,N_14735,N_14936);
and UO_409 (O_409,N_14924,N_14799);
nor UO_410 (O_410,N_14833,N_14754);
or UO_411 (O_411,N_14987,N_14700);
nand UO_412 (O_412,N_14896,N_14704);
xor UO_413 (O_413,N_14913,N_14944);
and UO_414 (O_414,N_14899,N_14839);
nand UO_415 (O_415,N_14987,N_14904);
nand UO_416 (O_416,N_14978,N_14923);
and UO_417 (O_417,N_14815,N_14756);
nand UO_418 (O_418,N_14722,N_14971);
or UO_419 (O_419,N_14923,N_14822);
and UO_420 (O_420,N_14873,N_14963);
nor UO_421 (O_421,N_14808,N_14926);
nand UO_422 (O_422,N_14776,N_14754);
xor UO_423 (O_423,N_14852,N_14724);
xor UO_424 (O_424,N_14843,N_14706);
and UO_425 (O_425,N_14714,N_14795);
or UO_426 (O_426,N_14878,N_14835);
and UO_427 (O_427,N_14943,N_14988);
or UO_428 (O_428,N_14947,N_14948);
and UO_429 (O_429,N_14733,N_14909);
xnor UO_430 (O_430,N_14948,N_14810);
xnor UO_431 (O_431,N_14702,N_14768);
nand UO_432 (O_432,N_14763,N_14866);
xor UO_433 (O_433,N_14708,N_14748);
or UO_434 (O_434,N_14871,N_14711);
or UO_435 (O_435,N_14723,N_14958);
and UO_436 (O_436,N_14834,N_14761);
or UO_437 (O_437,N_14805,N_14841);
and UO_438 (O_438,N_14989,N_14875);
xor UO_439 (O_439,N_14875,N_14734);
xor UO_440 (O_440,N_14863,N_14953);
nand UO_441 (O_441,N_14943,N_14773);
and UO_442 (O_442,N_14734,N_14811);
and UO_443 (O_443,N_14745,N_14847);
nor UO_444 (O_444,N_14775,N_14770);
and UO_445 (O_445,N_14747,N_14862);
xor UO_446 (O_446,N_14965,N_14711);
xnor UO_447 (O_447,N_14822,N_14889);
and UO_448 (O_448,N_14713,N_14939);
nor UO_449 (O_449,N_14765,N_14973);
and UO_450 (O_450,N_14827,N_14916);
nor UO_451 (O_451,N_14956,N_14771);
xnor UO_452 (O_452,N_14978,N_14755);
xnor UO_453 (O_453,N_14704,N_14840);
nor UO_454 (O_454,N_14932,N_14760);
or UO_455 (O_455,N_14732,N_14721);
and UO_456 (O_456,N_14736,N_14911);
and UO_457 (O_457,N_14714,N_14893);
nor UO_458 (O_458,N_14939,N_14994);
nor UO_459 (O_459,N_14899,N_14834);
or UO_460 (O_460,N_14838,N_14898);
and UO_461 (O_461,N_14800,N_14903);
and UO_462 (O_462,N_14831,N_14959);
xor UO_463 (O_463,N_14908,N_14856);
or UO_464 (O_464,N_14937,N_14756);
nand UO_465 (O_465,N_14920,N_14979);
or UO_466 (O_466,N_14898,N_14897);
nand UO_467 (O_467,N_14975,N_14859);
and UO_468 (O_468,N_14784,N_14968);
and UO_469 (O_469,N_14703,N_14996);
nor UO_470 (O_470,N_14746,N_14850);
and UO_471 (O_471,N_14992,N_14945);
nor UO_472 (O_472,N_14915,N_14720);
and UO_473 (O_473,N_14895,N_14914);
and UO_474 (O_474,N_14989,N_14958);
nor UO_475 (O_475,N_14742,N_14708);
nand UO_476 (O_476,N_14881,N_14965);
or UO_477 (O_477,N_14760,N_14809);
xor UO_478 (O_478,N_14728,N_14959);
xor UO_479 (O_479,N_14949,N_14883);
nor UO_480 (O_480,N_14938,N_14722);
nand UO_481 (O_481,N_14939,N_14880);
or UO_482 (O_482,N_14821,N_14980);
nor UO_483 (O_483,N_14972,N_14835);
or UO_484 (O_484,N_14829,N_14743);
nor UO_485 (O_485,N_14995,N_14917);
nor UO_486 (O_486,N_14864,N_14954);
or UO_487 (O_487,N_14789,N_14719);
nand UO_488 (O_488,N_14955,N_14817);
nor UO_489 (O_489,N_14813,N_14724);
nand UO_490 (O_490,N_14820,N_14827);
and UO_491 (O_491,N_14832,N_14899);
nor UO_492 (O_492,N_14846,N_14862);
xnor UO_493 (O_493,N_14740,N_14989);
nor UO_494 (O_494,N_14831,N_14944);
and UO_495 (O_495,N_14891,N_14803);
or UO_496 (O_496,N_14997,N_14841);
nand UO_497 (O_497,N_14781,N_14941);
nor UO_498 (O_498,N_14814,N_14750);
and UO_499 (O_499,N_14977,N_14728);
nand UO_500 (O_500,N_14976,N_14847);
or UO_501 (O_501,N_14911,N_14915);
nand UO_502 (O_502,N_14800,N_14763);
xnor UO_503 (O_503,N_14944,N_14947);
and UO_504 (O_504,N_14785,N_14977);
nand UO_505 (O_505,N_14865,N_14754);
nor UO_506 (O_506,N_14880,N_14836);
or UO_507 (O_507,N_14782,N_14915);
nor UO_508 (O_508,N_14966,N_14895);
and UO_509 (O_509,N_14822,N_14820);
xor UO_510 (O_510,N_14966,N_14788);
nand UO_511 (O_511,N_14874,N_14779);
nor UO_512 (O_512,N_14720,N_14868);
xor UO_513 (O_513,N_14787,N_14777);
xnor UO_514 (O_514,N_14841,N_14980);
and UO_515 (O_515,N_14937,N_14794);
nand UO_516 (O_516,N_14760,N_14857);
nand UO_517 (O_517,N_14888,N_14939);
and UO_518 (O_518,N_14804,N_14811);
nor UO_519 (O_519,N_14838,N_14965);
nor UO_520 (O_520,N_14872,N_14838);
and UO_521 (O_521,N_14912,N_14712);
nand UO_522 (O_522,N_14791,N_14760);
or UO_523 (O_523,N_14931,N_14879);
nand UO_524 (O_524,N_14712,N_14745);
and UO_525 (O_525,N_14984,N_14970);
or UO_526 (O_526,N_14895,N_14896);
xnor UO_527 (O_527,N_14815,N_14774);
nor UO_528 (O_528,N_14700,N_14977);
xnor UO_529 (O_529,N_14776,N_14966);
nand UO_530 (O_530,N_14982,N_14985);
xnor UO_531 (O_531,N_14896,N_14927);
xor UO_532 (O_532,N_14739,N_14892);
xnor UO_533 (O_533,N_14786,N_14999);
xnor UO_534 (O_534,N_14701,N_14957);
and UO_535 (O_535,N_14839,N_14949);
nand UO_536 (O_536,N_14746,N_14872);
nand UO_537 (O_537,N_14993,N_14700);
nand UO_538 (O_538,N_14716,N_14770);
nand UO_539 (O_539,N_14921,N_14839);
xor UO_540 (O_540,N_14720,N_14818);
nand UO_541 (O_541,N_14924,N_14995);
or UO_542 (O_542,N_14882,N_14819);
or UO_543 (O_543,N_14986,N_14992);
nand UO_544 (O_544,N_14703,N_14940);
nor UO_545 (O_545,N_14912,N_14838);
xor UO_546 (O_546,N_14946,N_14939);
and UO_547 (O_547,N_14764,N_14857);
xor UO_548 (O_548,N_14745,N_14835);
nand UO_549 (O_549,N_14863,N_14848);
xor UO_550 (O_550,N_14875,N_14897);
nand UO_551 (O_551,N_14724,N_14898);
nor UO_552 (O_552,N_14814,N_14911);
or UO_553 (O_553,N_14923,N_14987);
nand UO_554 (O_554,N_14807,N_14794);
xnor UO_555 (O_555,N_14742,N_14845);
xor UO_556 (O_556,N_14726,N_14809);
or UO_557 (O_557,N_14888,N_14867);
nand UO_558 (O_558,N_14956,N_14914);
xor UO_559 (O_559,N_14810,N_14957);
nor UO_560 (O_560,N_14764,N_14711);
or UO_561 (O_561,N_14909,N_14753);
nand UO_562 (O_562,N_14988,N_14857);
nor UO_563 (O_563,N_14779,N_14883);
or UO_564 (O_564,N_14785,N_14717);
nand UO_565 (O_565,N_14995,N_14793);
nor UO_566 (O_566,N_14896,N_14866);
xor UO_567 (O_567,N_14859,N_14979);
xor UO_568 (O_568,N_14819,N_14951);
or UO_569 (O_569,N_14996,N_14909);
nor UO_570 (O_570,N_14812,N_14715);
and UO_571 (O_571,N_14920,N_14814);
or UO_572 (O_572,N_14861,N_14958);
or UO_573 (O_573,N_14760,N_14830);
nand UO_574 (O_574,N_14903,N_14996);
or UO_575 (O_575,N_14937,N_14867);
nand UO_576 (O_576,N_14946,N_14976);
or UO_577 (O_577,N_14766,N_14856);
nand UO_578 (O_578,N_14873,N_14798);
nand UO_579 (O_579,N_14887,N_14880);
or UO_580 (O_580,N_14861,N_14757);
xnor UO_581 (O_581,N_14877,N_14838);
nor UO_582 (O_582,N_14726,N_14955);
and UO_583 (O_583,N_14863,N_14767);
xnor UO_584 (O_584,N_14854,N_14772);
nand UO_585 (O_585,N_14988,N_14751);
xor UO_586 (O_586,N_14725,N_14800);
and UO_587 (O_587,N_14750,N_14974);
or UO_588 (O_588,N_14976,N_14790);
or UO_589 (O_589,N_14905,N_14751);
nor UO_590 (O_590,N_14811,N_14793);
nand UO_591 (O_591,N_14717,N_14716);
or UO_592 (O_592,N_14823,N_14909);
nor UO_593 (O_593,N_14743,N_14817);
xor UO_594 (O_594,N_14704,N_14852);
and UO_595 (O_595,N_14800,N_14832);
xor UO_596 (O_596,N_14944,N_14982);
nand UO_597 (O_597,N_14734,N_14992);
nor UO_598 (O_598,N_14920,N_14809);
xnor UO_599 (O_599,N_14982,N_14702);
or UO_600 (O_600,N_14949,N_14748);
or UO_601 (O_601,N_14993,N_14896);
and UO_602 (O_602,N_14859,N_14834);
nor UO_603 (O_603,N_14773,N_14793);
xor UO_604 (O_604,N_14991,N_14967);
xnor UO_605 (O_605,N_14888,N_14815);
xor UO_606 (O_606,N_14707,N_14858);
and UO_607 (O_607,N_14702,N_14921);
and UO_608 (O_608,N_14775,N_14885);
nand UO_609 (O_609,N_14850,N_14928);
nand UO_610 (O_610,N_14875,N_14725);
and UO_611 (O_611,N_14768,N_14782);
and UO_612 (O_612,N_14736,N_14991);
nand UO_613 (O_613,N_14996,N_14862);
nand UO_614 (O_614,N_14905,N_14853);
nand UO_615 (O_615,N_14722,N_14707);
or UO_616 (O_616,N_14956,N_14822);
or UO_617 (O_617,N_14746,N_14822);
xor UO_618 (O_618,N_14810,N_14742);
nor UO_619 (O_619,N_14837,N_14708);
and UO_620 (O_620,N_14739,N_14867);
xor UO_621 (O_621,N_14937,N_14999);
and UO_622 (O_622,N_14973,N_14956);
or UO_623 (O_623,N_14920,N_14995);
nor UO_624 (O_624,N_14717,N_14831);
and UO_625 (O_625,N_14814,N_14827);
nand UO_626 (O_626,N_14971,N_14920);
nand UO_627 (O_627,N_14875,N_14759);
xor UO_628 (O_628,N_14791,N_14832);
nor UO_629 (O_629,N_14967,N_14730);
or UO_630 (O_630,N_14973,N_14933);
nor UO_631 (O_631,N_14973,N_14948);
and UO_632 (O_632,N_14705,N_14881);
or UO_633 (O_633,N_14761,N_14769);
and UO_634 (O_634,N_14732,N_14762);
xor UO_635 (O_635,N_14909,N_14830);
and UO_636 (O_636,N_14942,N_14835);
xor UO_637 (O_637,N_14832,N_14825);
nand UO_638 (O_638,N_14886,N_14760);
xnor UO_639 (O_639,N_14752,N_14951);
nand UO_640 (O_640,N_14977,N_14755);
nor UO_641 (O_641,N_14863,N_14782);
nor UO_642 (O_642,N_14740,N_14874);
and UO_643 (O_643,N_14704,N_14751);
and UO_644 (O_644,N_14974,N_14774);
and UO_645 (O_645,N_14921,N_14866);
nand UO_646 (O_646,N_14829,N_14744);
nor UO_647 (O_647,N_14758,N_14834);
nand UO_648 (O_648,N_14851,N_14852);
nand UO_649 (O_649,N_14815,N_14916);
nand UO_650 (O_650,N_14913,N_14995);
xor UO_651 (O_651,N_14904,N_14972);
nand UO_652 (O_652,N_14729,N_14760);
nand UO_653 (O_653,N_14756,N_14719);
or UO_654 (O_654,N_14975,N_14984);
or UO_655 (O_655,N_14996,N_14713);
xnor UO_656 (O_656,N_14872,N_14916);
xnor UO_657 (O_657,N_14850,N_14914);
or UO_658 (O_658,N_14810,N_14738);
and UO_659 (O_659,N_14702,N_14901);
xnor UO_660 (O_660,N_14731,N_14855);
nor UO_661 (O_661,N_14984,N_14834);
nand UO_662 (O_662,N_14886,N_14887);
and UO_663 (O_663,N_14935,N_14840);
nand UO_664 (O_664,N_14989,N_14737);
or UO_665 (O_665,N_14897,N_14798);
xnor UO_666 (O_666,N_14795,N_14753);
nand UO_667 (O_667,N_14937,N_14975);
nand UO_668 (O_668,N_14982,N_14923);
nor UO_669 (O_669,N_14918,N_14743);
or UO_670 (O_670,N_14903,N_14941);
or UO_671 (O_671,N_14916,N_14727);
and UO_672 (O_672,N_14744,N_14885);
nor UO_673 (O_673,N_14999,N_14753);
nand UO_674 (O_674,N_14779,N_14764);
xor UO_675 (O_675,N_14967,N_14835);
xor UO_676 (O_676,N_14954,N_14956);
nor UO_677 (O_677,N_14947,N_14708);
xor UO_678 (O_678,N_14742,N_14856);
and UO_679 (O_679,N_14722,N_14754);
nor UO_680 (O_680,N_14978,N_14916);
and UO_681 (O_681,N_14730,N_14824);
nand UO_682 (O_682,N_14996,N_14787);
nor UO_683 (O_683,N_14773,N_14940);
nor UO_684 (O_684,N_14956,N_14860);
or UO_685 (O_685,N_14957,N_14818);
and UO_686 (O_686,N_14719,N_14790);
nor UO_687 (O_687,N_14970,N_14711);
or UO_688 (O_688,N_14726,N_14941);
nand UO_689 (O_689,N_14754,N_14899);
or UO_690 (O_690,N_14884,N_14916);
nor UO_691 (O_691,N_14715,N_14933);
nor UO_692 (O_692,N_14912,N_14775);
nor UO_693 (O_693,N_14753,N_14941);
xor UO_694 (O_694,N_14840,N_14949);
nand UO_695 (O_695,N_14812,N_14757);
or UO_696 (O_696,N_14754,N_14743);
xnor UO_697 (O_697,N_14865,N_14781);
nand UO_698 (O_698,N_14804,N_14741);
and UO_699 (O_699,N_14896,N_14865);
nand UO_700 (O_700,N_14936,N_14905);
nor UO_701 (O_701,N_14919,N_14962);
and UO_702 (O_702,N_14993,N_14762);
nor UO_703 (O_703,N_14849,N_14707);
nor UO_704 (O_704,N_14833,N_14859);
xor UO_705 (O_705,N_14719,N_14936);
nand UO_706 (O_706,N_14860,N_14905);
or UO_707 (O_707,N_14854,N_14774);
and UO_708 (O_708,N_14847,N_14961);
xor UO_709 (O_709,N_14901,N_14898);
xnor UO_710 (O_710,N_14866,N_14778);
or UO_711 (O_711,N_14862,N_14743);
xor UO_712 (O_712,N_14745,N_14809);
xor UO_713 (O_713,N_14917,N_14808);
and UO_714 (O_714,N_14768,N_14869);
nand UO_715 (O_715,N_14713,N_14917);
xor UO_716 (O_716,N_14701,N_14757);
nand UO_717 (O_717,N_14834,N_14828);
xnor UO_718 (O_718,N_14728,N_14916);
nor UO_719 (O_719,N_14974,N_14803);
nand UO_720 (O_720,N_14708,N_14827);
xor UO_721 (O_721,N_14733,N_14783);
nor UO_722 (O_722,N_14863,N_14907);
xnor UO_723 (O_723,N_14955,N_14983);
or UO_724 (O_724,N_14713,N_14901);
xnor UO_725 (O_725,N_14978,N_14702);
xor UO_726 (O_726,N_14941,N_14895);
or UO_727 (O_727,N_14830,N_14783);
and UO_728 (O_728,N_14937,N_14973);
xnor UO_729 (O_729,N_14868,N_14758);
or UO_730 (O_730,N_14855,N_14716);
and UO_731 (O_731,N_14887,N_14799);
xnor UO_732 (O_732,N_14869,N_14957);
nand UO_733 (O_733,N_14827,N_14797);
nand UO_734 (O_734,N_14849,N_14792);
xor UO_735 (O_735,N_14753,N_14884);
nor UO_736 (O_736,N_14906,N_14966);
nand UO_737 (O_737,N_14722,N_14715);
nor UO_738 (O_738,N_14791,N_14861);
and UO_739 (O_739,N_14971,N_14863);
or UO_740 (O_740,N_14960,N_14825);
or UO_741 (O_741,N_14904,N_14989);
or UO_742 (O_742,N_14914,N_14836);
and UO_743 (O_743,N_14773,N_14801);
or UO_744 (O_744,N_14998,N_14773);
xnor UO_745 (O_745,N_14708,N_14780);
and UO_746 (O_746,N_14741,N_14872);
nor UO_747 (O_747,N_14775,N_14715);
or UO_748 (O_748,N_14761,N_14852);
nand UO_749 (O_749,N_14873,N_14911);
xnor UO_750 (O_750,N_14870,N_14788);
nand UO_751 (O_751,N_14719,N_14708);
and UO_752 (O_752,N_14702,N_14923);
xor UO_753 (O_753,N_14722,N_14986);
and UO_754 (O_754,N_14840,N_14937);
nand UO_755 (O_755,N_14902,N_14932);
or UO_756 (O_756,N_14891,N_14862);
or UO_757 (O_757,N_14940,N_14833);
xor UO_758 (O_758,N_14982,N_14902);
or UO_759 (O_759,N_14773,N_14904);
xnor UO_760 (O_760,N_14925,N_14979);
xnor UO_761 (O_761,N_14786,N_14867);
nor UO_762 (O_762,N_14892,N_14716);
xnor UO_763 (O_763,N_14989,N_14931);
and UO_764 (O_764,N_14839,N_14902);
nand UO_765 (O_765,N_14756,N_14743);
nand UO_766 (O_766,N_14807,N_14768);
or UO_767 (O_767,N_14712,N_14911);
or UO_768 (O_768,N_14730,N_14839);
or UO_769 (O_769,N_14775,N_14928);
or UO_770 (O_770,N_14873,N_14883);
or UO_771 (O_771,N_14876,N_14740);
or UO_772 (O_772,N_14825,N_14759);
nor UO_773 (O_773,N_14789,N_14978);
nor UO_774 (O_774,N_14928,N_14752);
nand UO_775 (O_775,N_14779,N_14861);
and UO_776 (O_776,N_14820,N_14825);
nor UO_777 (O_777,N_14849,N_14888);
xnor UO_778 (O_778,N_14877,N_14853);
nand UO_779 (O_779,N_14966,N_14995);
nand UO_780 (O_780,N_14700,N_14960);
nor UO_781 (O_781,N_14927,N_14762);
or UO_782 (O_782,N_14970,N_14778);
or UO_783 (O_783,N_14939,N_14786);
nor UO_784 (O_784,N_14760,N_14956);
nand UO_785 (O_785,N_14914,N_14838);
and UO_786 (O_786,N_14932,N_14764);
xor UO_787 (O_787,N_14723,N_14738);
xor UO_788 (O_788,N_14788,N_14839);
nand UO_789 (O_789,N_14894,N_14979);
xnor UO_790 (O_790,N_14868,N_14765);
xor UO_791 (O_791,N_14940,N_14859);
or UO_792 (O_792,N_14724,N_14883);
nand UO_793 (O_793,N_14767,N_14879);
xnor UO_794 (O_794,N_14903,N_14737);
or UO_795 (O_795,N_14701,N_14751);
nor UO_796 (O_796,N_14733,N_14781);
and UO_797 (O_797,N_14842,N_14947);
and UO_798 (O_798,N_14820,N_14974);
xnor UO_799 (O_799,N_14937,N_14752);
nand UO_800 (O_800,N_14849,N_14798);
or UO_801 (O_801,N_14866,N_14701);
and UO_802 (O_802,N_14786,N_14980);
nand UO_803 (O_803,N_14820,N_14922);
and UO_804 (O_804,N_14887,N_14701);
and UO_805 (O_805,N_14733,N_14764);
nand UO_806 (O_806,N_14845,N_14752);
nand UO_807 (O_807,N_14943,N_14957);
and UO_808 (O_808,N_14752,N_14953);
xor UO_809 (O_809,N_14935,N_14861);
or UO_810 (O_810,N_14738,N_14982);
nor UO_811 (O_811,N_14833,N_14979);
nand UO_812 (O_812,N_14871,N_14748);
or UO_813 (O_813,N_14851,N_14713);
or UO_814 (O_814,N_14780,N_14809);
xnor UO_815 (O_815,N_14742,N_14998);
xor UO_816 (O_816,N_14854,N_14780);
nor UO_817 (O_817,N_14792,N_14783);
nor UO_818 (O_818,N_14845,N_14724);
and UO_819 (O_819,N_14814,N_14811);
and UO_820 (O_820,N_14843,N_14772);
nand UO_821 (O_821,N_14794,N_14834);
xor UO_822 (O_822,N_14711,N_14770);
or UO_823 (O_823,N_14908,N_14781);
and UO_824 (O_824,N_14798,N_14868);
and UO_825 (O_825,N_14708,N_14796);
xnor UO_826 (O_826,N_14902,N_14886);
and UO_827 (O_827,N_14739,N_14792);
nand UO_828 (O_828,N_14877,N_14830);
or UO_829 (O_829,N_14834,N_14722);
or UO_830 (O_830,N_14791,N_14867);
xnor UO_831 (O_831,N_14804,N_14953);
xnor UO_832 (O_832,N_14749,N_14783);
xor UO_833 (O_833,N_14808,N_14800);
and UO_834 (O_834,N_14990,N_14881);
and UO_835 (O_835,N_14920,N_14829);
and UO_836 (O_836,N_14842,N_14833);
nor UO_837 (O_837,N_14783,N_14840);
nor UO_838 (O_838,N_14799,N_14794);
or UO_839 (O_839,N_14712,N_14831);
nor UO_840 (O_840,N_14907,N_14957);
nand UO_841 (O_841,N_14776,N_14964);
and UO_842 (O_842,N_14811,N_14963);
and UO_843 (O_843,N_14961,N_14715);
or UO_844 (O_844,N_14811,N_14859);
and UO_845 (O_845,N_14824,N_14819);
nor UO_846 (O_846,N_14740,N_14802);
nor UO_847 (O_847,N_14851,N_14903);
nand UO_848 (O_848,N_14744,N_14821);
or UO_849 (O_849,N_14843,N_14861);
nor UO_850 (O_850,N_14733,N_14968);
or UO_851 (O_851,N_14807,N_14951);
and UO_852 (O_852,N_14909,N_14789);
nand UO_853 (O_853,N_14794,N_14751);
xnor UO_854 (O_854,N_14765,N_14750);
nand UO_855 (O_855,N_14766,N_14873);
xor UO_856 (O_856,N_14909,N_14971);
nand UO_857 (O_857,N_14928,N_14984);
and UO_858 (O_858,N_14865,N_14709);
and UO_859 (O_859,N_14995,N_14821);
nor UO_860 (O_860,N_14975,N_14752);
and UO_861 (O_861,N_14928,N_14936);
nand UO_862 (O_862,N_14738,N_14816);
nor UO_863 (O_863,N_14823,N_14827);
nor UO_864 (O_864,N_14812,N_14771);
and UO_865 (O_865,N_14862,N_14861);
nor UO_866 (O_866,N_14763,N_14868);
nand UO_867 (O_867,N_14976,N_14848);
or UO_868 (O_868,N_14782,N_14757);
xor UO_869 (O_869,N_14803,N_14989);
or UO_870 (O_870,N_14819,N_14974);
xor UO_871 (O_871,N_14827,N_14705);
nor UO_872 (O_872,N_14892,N_14833);
nor UO_873 (O_873,N_14881,N_14833);
xor UO_874 (O_874,N_14808,N_14981);
nor UO_875 (O_875,N_14960,N_14810);
nor UO_876 (O_876,N_14970,N_14750);
nand UO_877 (O_877,N_14944,N_14879);
or UO_878 (O_878,N_14911,N_14890);
nand UO_879 (O_879,N_14715,N_14782);
nor UO_880 (O_880,N_14773,N_14974);
xor UO_881 (O_881,N_14946,N_14982);
or UO_882 (O_882,N_14800,N_14928);
xor UO_883 (O_883,N_14951,N_14753);
and UO_884 (O_884,N_14927,N_14814);
xor UO_885 (O_885,N_14817,N_14843);
nand UO_886 (O_886,N_14982,N_14931);
nand UO_887 (O_887,N_14951,N_14992);
nor UO_888 (O_888,N_14755,N_14709);
xnor UO_889 (O_889,N_14742,N_14928);
or UO_890 (O_890,N_14811,N_14987);
and UO_891 (O_891,N_14787,N_14708);
or UO_892 (O_892,N_14730,N_14940);
or UO_893 (O_893,N_14890,N_14726);
nor UO_894 (O_894,N_14917,N_14716);
nand UO_895 (O_895,N_14995,N_14816);
or UO_896 (O_896,N_14930,N_14844);
or UO_897 (O_897,N_14822,N_14937);
xor UO_898 (O_898,N_14978,N_14871);
xor UO_899 (O_899,N_14867,N_14938);
and UO_900 (O_900,N_14872,N_14948);
or UO_901 (O_901,N_14984,N_14996);
and UO_902 (O_902,N_14954,N_14932);
or UO_903 (O_903,N_14983,N_14891);
or UO_904 (O_904,N_14753,N_14808);
or UO_905 (O_905,N_14920,N_14953);
nor UO_906 (O_906,N_14933,N_14741);
nor UO_907 (O_907,N_14784,N_14928);
xnor UO_908 (O_908,N_14882,N_14929);
nor UO_909 (O_909,N_14851,N_14841);
nor UO_910 (O_910,N_14734,N_14901);
and UO_911 (O_911,N_14998,N_14912);
and UO_912 (O_912,N_14968,N_14854);
nor UO_913 (O_913,N_14969,N_14751);
and UO_914 (O_914,N_14754,N_14815);
or UO_915 (O_915,N_14788,N_14968);
xor UO_916 (O_916,N_14781,N_14905);
xnor UO_917 (O_917,N_14982,N_14758);
nand UO_918 (O_918,N_14840,N_14806);
nand UO_919 (O_919,N_14824,N_14750);
and UO_920 (O_920,N_14794,N_14897);
and UO_921 (O_921,N_14712,N_14714);
or UO_922 (O_922,N_14958,N_14732);
and UO_923 (O_923,N_14969,N_14992);
xnor UO_924 (O_924,N_14932,N_14965);
xor UO_925 (O_925,N_14821,N_14910);
xnor UO_926 (O_926,N_14884,N_14974);
or UO_927 (O_927,N_14850,N_14720);
or UO_928 (O_928,N_14981,N_14904);
xor UO_929 (O_929,N_14965,N_14877);
or UO_930 (O_930,N_14889,N_14853);
xor UO_931 (O_931,N_14771,N_14933);
xnor UO_932 (O_932,N_14990,N_14981);
and UO_933 (O_933,N_14896,N_14915);
and UO_934 (O_934,N_14925,N_14921);
nand UO_935 (O_935,N_14717,N_14864);
nand UO_936 (O_936,N_14836,N_14954);
or UO_937 (O_937,N_14812,N_14703);
xor UO_938 (O_938,N_14763,N_14874);
xnor UO_939 (O_939,N_14706,N_14958);
nand UO_940 (O_940,N_14968,N_14767);
xnor UO_941 (O_941,N_14744,N_14907);
or UO_942 (O_942,N_14942,N_14707);
nand UO_943 (O_943,N_14886,N_14831);
and UO_944 (O_944,N_14826,N_14806);
and UO_945 (O_945,N_14915,N_14917);
and UO_946 (O_946,N_14703,N_14820);
or UO_947 (O_947,N_14711,N_14931);
nand UO_948 (O_948,N_14764,N_14864);
nand UO_949 (O_949,N_14770,N_14860);
xor UO_950 (O_950,N_14713,N_14823);
and UO_951 (O_951,N_14825,N_14746);
or UO_952 (O_952,N_14720,N_14780);
nor UO_953 (O_953,N_14906,N_14792);
and UO_954 (O_954,N_14795,N_14850);
nor UO_955 (O_955,N_14965,N_14994);
and UO_956 (O_956,N_14965,N_14725);
or UO_957 (O_957,N_14909,N_14910);
nand UO_958 (O_958,N_14708,N_14810);
nand UO_959 (O_959,N_14806,N_14876);
and UO_960 (O_960,N_14991,N_14785);
nor UO_961 (O_961,N_14932,N_14766);
xor UO_962 (O_962,N_14764,N_14865);
or UO_963 (O_963,N_14766,N_14843);
xor UO_964 (O_964,N_14716,N_14852);
xnor UO_965 (O_965,N_14988,N_14744);
or UO_966 (O_966,N_14875,N_14956);
xnor UO_967 (O_967,N_14840,N_14842);
nor UO_968 (O_968,N_14838,N_14936);
and UO_969 (O_969,N_14877,N_14995);
or UO_970 (O_970,N_14819,N_14769);
nor UO_971 (O_971,N_14884,N_14794);
or UO_972 (O_972,N_14844,N_14888);
nand UO_973 (O_973,N_14811,N_14805);
nor UO_974 (O_974,N_14835,N_14890);
nand UO_975 (O_975,N_14857,N_14846);
and UO_976 (O_976,N_14893,N_14777);
nor UO_977 (O_977,N_14796,N_14701);
xor UO_978 (O_978,N_14918,N_14942);
xnor UO_979 (O_979,N_14812,N_14769);
xor UO_980 (O_980,N_14859,N_14903);
nand UO_981 (O_981,N_14745,N_14750);
and UO_982 (O_982,N_14932,N_14836);
xnor UO_983 (O_983,N_14857,N_14717);
or UO_984 (O_984,N_14774,N_14960);
nor UO_985 (O_985,N_14723,N_14936);
nand UO_986 (O_986,N_14952,N_14760);
or UO_987 (O_987,N_14850,N_14925);
xnor UO_988 (O_988,N_14838,N_14889);
nor UO_989 (O_989,N_14816,N_14886);
nor UO_990 (O_990,N_14751,N_14967);
and UO_991 (O_991,N_14964,N_14735);
or UO_992 (O_992,N_14909,N_14772);
xnor UO_993 (O_993,N_14795,N_14991);
or UO_994 (O_994,N_14738,N_14937);
or UO_995 (O_995,N_14721,N_14803);
and UO_996 (O_996,N_14824,N_14726);
nor UO_997 (O_997,N_14900,N_14743);
or UO_998 (O_998,N_14807,N_14727);
or UO_999 (O_999,N_14947,N_14771);
xor UO_1000 (O_1000,N_14768,N_14761);
xor UO_1001 (O_1001,N_14851,N_14948);
and UO_1002 (O_1002,N_14745,N_14705);
and UO_1003 (O_1003,N_14825,N_14821);
or UO_1004 (O_1004,N_14900,N_14977);
xor UO_1005 (O_1005,N_14822,N_14871);
xnor UO_1006 (O_1006,N_14775,N_14843);
or UO_1007 (O_1007,N_14859,N_14765);
nand UO_1008 (O_1008,N_14766,N_14872);
nand UO_1009 (O_1009,N_14714,N_14923);
nand UO_1010 (O_1010,N_14759,N_14848);
nand UO_1011 (O_1011,N_14876,N_14709);
nor UO_1012 (O_1012,N_14805,N_14887);
xnor UO_1013 (O_1013,N_14947,N_14787);
xnor UO_1014 (O_1014,N_14703,N_14960);
nand UO_1015 (O_1015,N_14800,N_14891);
or UO_1016 (O_1016,N_14853,N_14737);
or UO_1017 (O_1017,N_14774,N_14911);
xor UO_1018 (O_1018,N_14867,N_14972);
and UO_1019 (O_1019,N_14936,N_14850);
and UO_1020 (O_1020,N_14788,N_14735);
and UO_1021 (O_1021,N_14859,N_14964);
nor UO_1022 (O_1022,N_14926,N_14809);
nand UO_1023 (O_1023,N_14773,N_14853);
or UO_1024 (O_1024,N_14991,N_14924);
xor UO_1025 (O_1025,N_14977,N_14915);
and UO_1026 (O_1026,N_14911,N_14794);
and UO_1027 (O_1027,N_14893,N_14988);
xor UO_1028 (O_1028,N_14719,N_14709);
or UO_1029 (O_1029,N_14998,N_14827);
nor UO_1030 (O_1030,N_14823,N_14754);
and UO_1031 (O_1031,N_14881,N_14712);
and UO_1032 (O_1032,N_14768,N_14728);
nor UO_1033 (O_1033,N_14988,N_14883);
nand UO_1034 (O_1034,N_14808,N_14703);
or UO_1035 (O_1035,N_14744,N_14938);
nor UO_1036 (O_1036,N_14879,N_14715);
xnor UO_1037 (O_1037,N_14901,N_14741);
or UO_1038 (O_1038,N_14886,N_14855);
xor UO_1039 (O_1039,N_14724,N_14945);
nor UO_1040 (O_1040,N_14773,N_14755);
xnor UO_1041 (O_1041,N_14950,N_14740);
nor UO_1042 (O_1042,N_14922,N_14702);
or UO_1043 (O_1043,N_14736,N_14893);
and UO_1044 (O_1044,N_14787,N_14955);
and UO_1045 (O_1045,N_14802,N_14731);
and UO_1046 (O_1046,N_14836,N_14703);
nand UO_1047 (O_1047,N_14795,N_14825);
nor UO_1048 (O_1048,N_14731,N_14771);
or UO_1049 (O_1049,N_14769,N_14710);
xor UO_1050 (O_1050,N_14700,N_14917);
and UO_1051 (O_1051,N_14967,N_14938);
and UO_1052 (O_1052,N_14765,N_14810);
xnor UO_1053 (O_1053,N_14889,N_14964);
or UO_1054 (O_1054,N_14718,N_14795);
xnor UO_1055 (O_1055,N_14979,N_14769);
nor UO_1056 (O_1056,N_14752,N_14721);
or UO_1057 (O_1057,N_14799,N_14977);
nand UO_1058 (O_1058,N_14851,N_14768);
or UO_1059 (O_1059,N_14774,N_14898);
xnor UO_1060 (O_1060,N_14799,N_14744);
xnor UO_1061 (O_1061,N_14908,N_14772);
or UO_1062 (O_1062,N_14735,N_14907);
nand UO_1063 (O_1063,N_14920,N_14721);
nor UO_1064 (O_1064,N_14926,N_14802);
and UO_1065 (O_1065,N_14759,N_14767);
xor UO_1066 (O_1066,N_14878,N_14730);
nand UO_1067 (O_1067,N_14893,N_14713);
xor UO_1068 (O_1068,N_14910,N_14934);
xnor UO_1069 (O_1069,N_14736,N_14746);
and UO_1070 (O_1070,N_14871,N_14809);
or UO_1071 (O_1071,N_14798,N_14865);
nor UO_1072 (O_1072,N_14844,N_14860);
and UO_1073 (O_1073,N_14823,N_14907);
nor UO_1074 (O_1074,N_14731,N_14816);
nand UO_1075 (O_1075,N_14741,N_14706);
and UO_1076 (O_1076,N_14798,N_14907);
or UO_1077 (O_1077,N_14970,N_14892);
or UO_1078 (O_1078,N_14954,N_14883);
nor UO_1079 (O_1079,N_14717,N_14916);
and UO_1080 (O_1080,N_14934,N_14852);
and UO_1081 (O_1081,N_14823,N_14833);
or UO_1082 (O_1082,N_14868,N_14705);
nand UO_1083 (O_1083,N_14819,N_14860);
and UO_1084 (O_1084,N_14706,N_14775);
nand UO_1085 (O_1085,N_14711,N_14949);
xnor UO_1086 (O_1086,N_14987,N_14749);
xnor UO_1087 (O_1087,N_14700,N_14788);
xor UO_1088 (O_1088,N_14986,N_14869);
nor UO_1089 (O_1089,N_14712,N_14892);
or UO_1090 (O_1090,N_14783,N_14974);
and UO_1091 (O_1091,N_14819,N_14869);
xor UO_1092 (O_1092,N_14952,N_14816);
xor UO_1093 (O_1093,N_14981,N_14847);
nor UO_1094 (O_1094,N_14769,N_14732);
nor UO_1095 (O_1095,N_14995,N_14783);
or UO_1096 (O_1096,N_14857,N_14777);
nor UO_1097 (O_1097,N_14771,N_14790);
or UO_1098 (O_1098,N_14709,N_14756);
or UO_1099 (O_1099,N_14991,N_14781);
xor UO_1100 (O_1100,N_14741,N_14854);
xnor UO_1101 (O_1101,N_14706,N_14866);
nand UO_1102 (O_1102,N_14987,N_14739);
or UO_1103 (O_1103,N_14888,N_14897);
or UO_1104 (O_1104,N_14763,N_14925);
nor UO_1105 (O_1105,N_14815,N_14816);
and UO_1106 (O_1106,N_14913,N_14706);
nand UO_1107 (O_1107,N_14812,N_14761);
and UO_1108 (O_1108,N_14825,N_14814);
nor UO_1109 (O_1109,N_14890,N_14966);
or UO_1110 (O_1110,N_14719,N_14798);
and UO_1111 (O_1111,N_14869,N_14703);
nand UO_1112 (O_1112,N_14962,N_14743);
nand UO_1113 (O_1113,N_14966,N_14797);
and UO_1114 (O_1114,N_14923,N_14855);
and UO_1115 (O_1115,N_14971,N_14887);
xnor UO_1116 (O_1116,N_14862,N_14714);
nand UO_1117 (O_1117,N_14921,N_14874);
nor UO_1118 (O_1118,N_14992,N_14917);
and UO_1119 (O_1119,N_14708,N_14889);
or UO_1120 (O_1120,N_14723,N_14800);
nand UO_1121 (O_1121,N_14844,N_14730);
and UO_1122 (O_1122,N_14947,N_14913);
or UO_1123 (O_1123,N_14935,N_14827);
nor UO_1124 (O_1124,N_14887,N_14825);
nand UO_1125 (O_1125,N_14777,N_14990);
xnor UO_1126 (O_1126,N_14912,N_14911);
xor UO_1127 (O_1127,N_14774,N_14895);
nor UO_1128 (O_1128,N_14952,N_14994);
nand UO_1129 (O_1129,N_14953,N_14895);
xnor UO_1130 (O_1130,N_14749,N_14995);
xor UO_1131 (O_1131,N_14822,N_14765);
or UO_1132 (O_1132,N_14894,N_14910);
and UO_1133 (O_1133,N_14774,N_14768);
or UO_1134 (O_1134,N_14706,N_14717);
nor UO_1135 (O_1135,N_14779,N_14952);
nand UO_1136 (O_1136,N_14972,N_14934);
xor UO_1137 (O_1137,N_14851,N_14797);
nor UO_1138 (O_1138,N_14959,N_14951);
nor UO_1139 (O_1139,N_14961,N_14854);
xor UO_1140 (O_1140,N_14959,N_14790);
or UO_1141 (O_1141,N_14876,N_14980);
or UO_1142 (O_1142,N_14818,N_14804);
nor UO_1143 (O_1143,N_14778,N_14908);
nand UO_1144 (O_1144,N_14927,N_14818);
xor UO_1145 (O_1145,N_14755,N_14704);
and UO_1146 (O_1146,N_14886,N_14843);
nand UO_1147 (O_1147,N_14964,N_14835);
xnor UO_1148 (O_1148,N_14998,N_14780);
nor UO_1149 (O_1149,N_14960,N_14940);
nor UO_1150 (O_1150,N_14947,N_14801);
nand UO_1151 (O_1151,N_14843,N_14933);
or UO_1152 (O_1152,N_14954,N_14777);
and UO_1153 (O_1153,N_14885,N_14710);
xor UO_1154 (O_1154,N_14970,N_14922);
nand UO_1155 (O_1155,N_14880,N_14988);
and UO_1156 (O_1156,N_14898,N_14884);
xnor UO_1157 (O_1157,N_14864,N_14941);
nand UO_1158 (O_1158,N_14740,N_14947);
xor UO_1159 (O_1159,N_14968,N_14992);
nand UO_1160 (O_1160,N_14881,N_14983);
xnor UO_1161 (O_1161,N_14811,N_14864);
or UO_1162 (O_1162,N_14995,N_14982);
xor UO_1163 (O_1163,N_14805,N_14725);
and UO_1164 (O_1164,N_14837,N_14706);
and UO_1165 (O_1165,N_14948,N_14915);
nand UO_1166 (O_1166,N_14985,N_14832);
nand UO_1167 (O_1167,N_14777,N_14981);
nor UO_1168 (O_1168,N_14846,N_14867);
xor UO_1169 (O_1169,N_14856,N_14803);
or UO_1170 (O_1170,N_14751,N_14922);
nand UO_1171 (O_1171,N_14794,N_14786);
nor UO_1172 (O_1172,N_14902,N_14703);
or UO_1173 (O_1173,N_14752,N_14856);
nor UO_1174 (O_1174,N_14941,N_14932);
nand UO_1175 (O_1175,N_14974,N_14936);
or UO_1176 (O_1176,N_14979,N_14935);
and UO_1177 (O_1177,N_14713,N_14841);
nor UO_1178 (O_1178,N_14858,N_14835);
and UO_1179 (O_1179,N_14899,N_14866);
and UO_1180 (O_1180,N_14825,N_14868);
and UO_1181 (O_1181,N_14850,N_14798);
or UO_1182 (O_1182,N_14917,N_14991);
nand UO_1183 (O_1183,N_14815,N_14751);
nand UO_1184 (O_1184,N_14794,N_14753);
and UO_1185 (O_1185,N_14900,N_14833);
nand UO_1186 (O_1186,N_14906,N_14833);
or UO_1187 (O_1187,N_14871,N_14737);
or UO_1188 (O_1188,N_14862,N_14725);
xor UO_1189 (O_1189,N_14941,N_14992);
xor UO_1190 (O_1190,N_14833,N_14971);
xor UO_1191 (O_1191,N_14785,N_14714);
nand UO_1192 (O_1192,N_14906,N_14705);
xnor UO_1193 (O_1193,N_14912,N_14753);
and UO_1194 (O_1194,N_14773,N_14856);
nand UO_1195 (O_1195,N_14941,N_14958);
nor UO_1196 (O_1196,N_14969,N_14815);
or UO_1197 (O_1197,N_14728,N_14719);
and UO_1198 (O_1198,N_14804,N_14906);
and UO_1199 (O_1199,N_14833,N_14963);
or UO_1200 (O_1200,N_14793,N_14902);
and UO_1201 (O_1201,N_14897,N_14946);
nor UO_1202 (O_1202,N_14758,N_14823);
and UO_1203 (O_1203,N_14833,N_14817);
xnor UO_1204 (O_1204,N_14832,N_14948);
and UO_1205 (O_1205,N_14850,N_14950);
or UO_1206 (O_1206,N_14984,N_14824);
nand UO_1207 (O_1207,N_14967,N_14741);
or UO_1208 (O_1208,N_14934,N_14814);
xnor UO_1209 (O_1209,N_14927,N_14962);
nor UO_1210 (O_1210,N_14830,N_14815);
or UO_1211 (O_1211,N_14713,N_14951);
or UO_1212 (O_1212,N_14779,N_14850);
xnor UO_1213 (O_1213,N_14926,N_14943);
xor UO_1214 (O_1214,N_14999,N_14789);
and UO_1215 (O_1215,N_14909,N_14924);
xor UO_1216 (O_1216,N_14939,N_14779);
xnor UO_1217 (O_1217,N_14916,N_14798);
xnor UO_1218 (O_1218,N_14999,N_14865);
xor UO_1219 (O_1219,N_14857,N_14990);
nand UO_1220 (O_1220,N_14943,N_14941);
xnor UO_1221 (O_1221,N_14853,N_14919);
nand UO_1222 (O_1222,N_14967,N_14892);
xnor UO_1223 (O_1223,N_14718,N_14874);
xnor UO_1224 (O_1224,N_14825,N_14979);
nor UO_1225 (O_1225,N_14980,N_14709);
xor UO_1226 (O_1226,N_14747,N_14981);
nand UO_1227 (O_1227,N_14913,N_14894);
and UO_1228 (O_1228,N_14709,N_14961);
and UO_1229 (O_1229,N_14887,N_14774);
nand UO_1230 (O_1230,N_14910,N_14711);
and UO_1231 (O_1231,N_14763,N_14961);
nor UO_1232 (O_1232,N_14836,N_14949);
xnor UO_1233 (O_1233,N_14913,N_14730);
nor UO_1234 (O_1234,N_14738,N_14922);
or UO_1235 (O_1235,N_14805,N_14751);
nand UO_1236 (O_1236,N_14930,N_14736);
xnor UO_1237 (O_1237,N_14922,N_14710);
and UO_1238 (O_1238,N_14749,N_14937);
or UO_1239 (O_1239,N_14959,N_14852);
or UO_1240 (O_1240,N_14839,N_14783);
and UO_1241 (O_1241,N_14804,N_14769);
nor UO_1242 (O_1242,N_14889,N_14789);
nand UO_1243 (O_1243,N_14826,N_14859);
nor UO_1244 (O_1244,N_14803,N_14716);
nor UO_1245 (O_1245,N_14938,N_14729);
xnor UO_1246 (O_1246,N_14946,N_14712);
nor UO_1247 (O_1247,N_14721,N_14877);
nand UO_1248 (O_1248,N_14851,N_14793);
nor UO_1249 (O_1249,N_14874,N_14726);
nor UO_1250 (O_1250,N_14843,N_14754);
nor UO_1251 (O_1251,N_14758,N_14837);
nor UO_1252 (O_1252,N_14882,N_14739);
nand UO_1253 (O_1253,N_14877,N_14831);
xor UO_1254 (O_1254,N_14816,N_14701);
xnor UO_1255 (O_1255,N_14832,N_14976);
nand UO_1256 (O_1256,N_14754,N_14855);
xor UO_1257 (O_1257,N_14998,N_14741);
and UO_1258 (O_1258,N_14920,N_14863);
xnor UO_1259 (O_1259,N_14760,N_14801);
and UO_1260 (O_1260,N_14916,N_14941);
and UO_1261 (O_1261,N_14975,N_14940);
xnor UO_1262 (O_1262,N_14981,N_14899);
xor UO_1263 (O_1263,N_14738,N_14944);
or UO_1264 (O_1264,N_14937,N_14929);
nor UO_1265 (O_1265,N_14782,N_14905);
xor UO_1266 (O_1266,N_14755,N_14787);
nand UO_1267 (O_1267,N_14823,N_14751);
nand UO_1268 (O_1268,N_14859,N_14837);
xor UO_1269 (O_1269,N_14750,N_14778);
xor UO_1270 (O_1270,N_14859,N_14706);
xor UO_1271 (O_1271,N_14911,N_14933);
nand UO_1272 (O_1272,N_14748,N_14853);
nor UO_1273 (O_1273,N_14975,N_14807);
xor UO_1274 (O_1274,N_14837,N_14834);
and UO_1275 (O_1275,N_14943,N_14895);
and UO_1276 (O_1276,N_14739,N_14944);
and UO_1277 (O_1277,N_14837,N_14848);
and UO_1278 (O_1278,N_14901,N_14921);
nand UO_1279 (O_1279,N_14889,N_14805);
xor UO_1280 (O_1280,N_14952,N_14933);
xnor UO_1281 (O_1281,N_14767,N_14839);
nor UO_1282 (O_1282,N_14746,N_14836);
xor UO_1283 (O_1283,N_14994,N_14889);
or UO_1284 (O_1284,N_14764,N_14830);
xnor UO_1285 (O_1285,N_14716,N_14885);
nand UO_1286 (O_1286,N_14832,N_14758);
xnor UO_1287 (O_1287,N_14943,N_14912);
or UO_1288 (O_1288,N_14816,N_14772);
nand UO_1289 (O_1289,N_14764,N_14995);
nor UO_1290 (O_1290,N_14971,N_14933);
and UO_1291 (O_1291,N_14755,N_14934);
nor UO_1292 (O_1292,N_14940,N_14994);
nor UO_1293 (O_1293,N_14783,N_14925);
nor UO_1294 (O_1294,N_14912,N_14709);
or UO_1295 (O_1295,N_14965,N_14811);
or UO_1296 (O_1296,N_14882,N_14735);
xor UO_1297 (O_1297,N_14974,N_14953);
nand UO_1298 (O_1298,N_14878,N_14994);
nand UO_1299 (O_1299,N_14813,N_14855);
xor UO_1300 (O_1300,N_14823,N_14966);
and UO_1301 (O_1301,N_14803,N_14794);
and UO_1302 (O_1302,N_14884,N_14715);
and UO_1303 (O_1303,N_14857,N_14930);
nor UO_1304 (O_1304,N_14819,N_14740);
nor UO_1305 (O_1305,N_14928,N_14974);
nand UO_1306 (O_1306,N_14938,N_14856);
or UO_1307 (O_1307,N_14905,N_14984);
xor UO_1308 (O_1308,N_14853,N_14763);
nor UO_1309 (O_1309,N_14958,N_14909);
or UO_1310 (O_1310,N_14823,N_14733);
nor UO_1311 (O_1311,N_14717,N_14953);
nand UO_1312 (O_1312,N_14937,N_14736);
nand UO_1313 (O_1313,N_14922,N_14884);
and UO_1314 (O_1314,N_14713,N_14706);
nor UO_1315 (O_1315,N_14976,N_14969);
xnor UO_1316 (O_1316,N_14741,N_14853);
xnor UO_1317 (O_1317,N_14920,N_14944);
xnor UO_1318 (O_1318,N_14957,N_14733);
xor UO_1319 (O_1319,N_14935,N_14819);
nor UO_1320 (O_1320,N_14756,N_14847);
or UO_1321 (O_1321,N_14899,N_14714);
nor UO_1322 (O_1322,N_14958,N_14809);
and UO_1323 (O_1323,N_14829,N_14728);
nor UO_1324 (O_1324,N_14785,N_14948);
and UO_1325 (O_1325,N_14891,N_14796);
or UO_1326 (O_1326,N_14882,N_14798);
xnor UO_1327 (O_1327,N_14830,N_14993);
nor UO_1328 (O_1328,N_14802,N_14852);
nand UO_1329 (O_1329,N_14850,N_14876);
or UO_1330 (O_1330,N_14895,N_14806);
nor UO_1331 (O_1331,N_14893,N_14737);
nor UO_1332 (O_1332,N_14851,N_14837);
and UO_1333 (O_1333,N_14847,N_14831);
nand UO_1334 (O_1334,N_14966,N_14701);
nor UO_1335 (O_1335,N_14798,N_14727);
xor UO_1336 (O_1336,N_14790,N_14942);
nor UO_1337 (O_1337,N_14988,N_14858);
nor UO_1338 (O_1338,N_14906,N_14914);
nor UO_1339 (O_1339,N_14741,N_14975);
nand UO_1340 (O_1340,N_14784,N_14913);
or UO_1341 (O_1341,N_14854,N_14782);
or UO_1342 (O_1342,N_14794,N_14755);
xnor UO_1343 (O_1343,N_14725,N_14883);
nand UO_1344 (O_1344,N_14779,N_14870);
nor UO_1345 (O_1345,N_14881,N_14908);
and UO_1346 (O_1346,N_14775,N_14825);
nand UO_1347 (O_1347,N_14707,N_14967);
nor UO_1348 (O_1348,N_14737,N_14736);
nand UO_1349 (O_1349,N_14950,N_14907);
nand UO_1350 (O_1350,N_14729,N_14916);
xor UO_1351 (O_1351,N_14945,N_14975);
or UO_1352 (O_1352,N_14732,N_14811);
and UO_1353 (O_1353,N_14748,N_14877);
and UO_1354 (O_1354,N_14787,N_14793);
or UO_1355 (O_1355,N_14856,N_14911);
xnor UO_1356 (O_1356,N_14863,N_14858);
xor UO_1357 (O_1357,N_14724,N_14903);
nand UO_1358 (O_1358,N_14722,N_14858);
or UO_1359 (O_1359,N_14970,N_14940);
nor UO_1360 (O_1360,N_14819,N_14911);
nand UO_1361 (O_1361,N_14785,N_14838);
and UO_1362 (O_1362,N_14915,N_14746);
or UO_1363 (O_1363,N_14722,N_14764);
xnor UO_1364 (O_1364,N_14933,N_14924);
nand UO_1365 (O_1365,N_14741,N_14952);
xnor UO_1366 (O_1366,N_14920,N_14847);
nor UO_1367 (O_1367,N_14988,N_14713);
and UO_1368 (O_1368,N_14829,N_14802);
nand UO_1369 (O_1369,N_14762,N_14718);
nor UO_1370 (O_1370,N_14713,N_14816);
and UO_1371 (O_1371,N_14994,N_14992);
or UO_1372 (O_1372,N_14805,N_14746);
and UO_1373 (O_1373,N_14806,N_14818);
and UO_1374 (O_1374,N_14821,N_14713);
and UO_1375 (O_1375,N_14938,N_14762);
nand UO_1376 (O_1376,N_14813,N_14745);
or UO_1377 (O_1377,N_14906,N_14974);
xor UO_1378 (O_1378,N_14865,N_14958);
xnor UO_1379 (O_1379,N_14702,N_14979);
or UO_1380 (O_1380,N_14819,N_14709);
and UO_1381 (O_1381,N_14785,N_14826);
nor UO_1382 (O_1382,N_14770,N_14733);
xor UO_1383 (O_1383,N_14890,N_14751);
nand UO_1384 (O_1384,N_14785,N_14718);
nor UO_1385 (O_1385,N_14912,N_14867);
nand UO_1386 (O_1386,N_14942,N_14977);
nor UO_1387 (O_1387,N_14861,N_14940);
and UO_1388 (O_1388,N_14892,N_14848);
nor UO_1389 (O_1389,N_14919,N_14738);
nor UO_1390 (O_1390,N_14845,N_14895);
xnor UO_1391 (O_1391,N_14956,N_14704);
xnor UO_1392 (O_1392,N_14828,N_14707);
nor UO_1393 (O_1393,N_14774,N_14975);
nand UO_1394 (O_1394,N_14933,N_14913);
xnor UO_1395 (O_1395,N_14904,N_14764);
xor UO_1396 (O_1396,N_14869,N_14801);
nand UO_1397 (O_1397,N_14909,N_14806);
nor UO_1398 (O_1398,N_14765,N_14806);
xnor UO_1399 (O_1399,N_14742,N_14773);
or UO_1400 (O_1400,N_14771,N_14795);
or UO_1401 (O_1401,N_14881,N_14931);
or UO_1402 (O_1402,N_14833,N_14776);
nor UO_1403 (O_1403,N_14760,N_14938);
xnor UO_1404 (O_1404,N_14793,N_14803);
or UO_1405 (O_1405,N_14706,N_14829);
nand UO_1406 (O_1406,N_14835,N_14874);
nor UO_1407 (O_1407,N_14915,N_14928);
and UO_1408 (O_1408,N_14805,N_14719);
and UO_1409 (O_1409,N_14884,N_14874);
nand UO_1410 (O_1410,N_14760,N_14996);
nand UO_1411 (O_1411,N_14998,N_14958);
and UO_1412 (O_1412,N_14906,N_14801);
nand UO_1413 (O_1413,N_14777,N_14979);
and UO_1414 (O_1414,N_14928,N_14940);
xnor UO_1415 (O_1415,N_14936,N_14765);
nor UO_1416 (O_1416,N_14890,N_14876);
and UO_1417 (O_1417,N_14807,N_14802);
and UO_1418 (O_1418,N_14756,N_14891);
and UO_1419 (O_1419,N_14775,N_14718);
xnor UO_1420 (O_1420,N_14991,N_14790);
xor UO_1421 (O_1421,N_14704,N_14839);
or UO_1422 (O_1422,N_14720,N_14878);
nor UO_1423 (O_1423,N_14934,N_14801);
nand UO_1424 (O_1424,N_14824,N_14811);
nand UO_1425 (O_1425,N_14998,N_14737);
xnor UO_1426 (O_1426,N_14922,N_14704);
nor UO_1427 (O_1427,N_14760,N_14808);
or UO_1428 (O_1428,N_14736,N_14929);
and UO_1429 (O_1429,N_14958,N_14709);
nand UO_1430 (O_1430,N_14771,N_14938);
and UO_1431 (O_1431,N_14849,N_14900);
nor UO_1432 (O_1432,N_14756,N_14769);
xor UO_1433 (O_1433,N_14766,N_14916);
nand UO_1434 (O_1434,N_14725,N_14741);
and UO_1435 (O_1435,N_14842,N_14941);
or UO_1436 (O_1436,N_14867,N_14737);
or UO_1437 (O_1437,N_14760,N_14810);
nand UO_1438 (O_1438,N_14774,N_14712);
and UO_1439 (O_1439,N_14929,N_14754);
and UO_1440 (O_1440,N_14834,N_14904);
or UO_1441 (O_1441,N_14988,N_14749);
or UO_1442 (O_1442,N_14759,N_14720);
or UO_1443 (O_1443,N_14834,N_14886);
or UO_1444 (O_1444,N_14969,N_14831);
nand UO_1445 (O_1445,N_14774,N_14812);
nand UO_1446 (O_1446,N_14892,N_14996);
or UO_1447 (O_1447,N_14810,N_14789);
and UO_1448 (O_1448,N_14979,N_14881);
and UO_1449 (O_1449,N_14981,N_14970);
xor UO_1450 (O_1450,N_14961,N_14707);
and UO_1451 (O_1451,N_14780,N_14953);
xnor UO_1452 (O_1452,N_14823,N_14701);
and UO_1453 (O_1453,N_14873,N_14981);
nand UO_1454 (O_1454,N_14948,N_14794);
nor UO_1455 (O_1455,N_14892,N_14875);
and UO_1456 (O_1456,N_14817,N_14805);
xnor UO_1457 (O_1457,N_14916,N_14942);
nand UO_1458 (O_1458,N_14772,N_14804);
and UO_1459 (O_1459,N_14773,N_14869);
xnor UO_1460 (O_1460,N_14817,N_14857);
nand UO_1461 (O_1461,N_14797,N_14920);
xor UO_1462 (O_1462,N_14900,N_14963);
xnor UO_1463 (O_1463,N_14990,N_14804);
xnor UO_1464 (O_1464,N_14914,N_14932);
and UO_1465 (O_1465,N_14794,N_14742);
nand UO_1466 (O_1466,N_14987,N_14851);
or UO_1467 (O_1467,N_14787,N_14863);
and UO_1468 (O_1468,N_14962,N_14737);
nand UO_1469 (O_1469,N_14938,N_14998);
and UO_1470 (O_1470,N_14801,N_14904);
and UO_1471 (O_1471,N_14907,N_14827);
nand UO_1472 (O_1472,N_14817,N_14706);
nand UO_1473 (O_1473,N_14932,N_14759);
and UO_1474 (O_1474,N_14763,N_14930);
nand UO_1475 (O_1475,N_14870,N_14745);
nor UO_1476 (O_1476,N_14982,N_14883);
nand UO_1477 (O_1477,N_14794,N_14765);
nor UO_1478 (O_1478,N_14957,N_14920);
or UO_1479 (O_1479,N_14930,N_14734);
or UO_1480 (O_1480,N_14953,N_14701);
nand UO_1481 (O_1481,N_14778,N_14789);
xnor UO_1482 (O_1482,N_14869,N_14850);
or UO_1483 (O_1483,N_14962,N_14934);
or UO_1484 (O_1484,N_14744,N_14760);
and UO_1485 (O_1485,N_14783,N_14955);
nor UO_1486 (O_1486,N_14935,N_14901);
nand UO_1487 (O_1487,N_14901,N_14911);
nor UO_1488 (O_1488,N_14917,N_14819);
or UO_1489 (O_1489,N_14842,N_14730);
nand UO_1490 (O_1490,N_14728,N_14752);
or UO_1491 (O_1491,N_14715,N_14904);
nor UO_1492 (O_1492,N_14831,N_14985);
or UO_1493 (O_1493,N_14750,N_14897);
xor UO_1494 (O_1494,N_14866,N_14952);
nor UO_1495 (O_1495,N_14717,N_14792);
nor UO_1496 (O_1496,N_14961,N_14884);
xnor UO_1497 (O_1497,N_14725,N_14960);
or UO_1498 (O_1498,N_14719,N_14812);
nor UO_1499 (O_1499,N_14922,N_14920);
and UO_1500 (O_1500,N_14709,N_14702);
and UO_1501 (O_1501,N_14944,N_14851);
nor UO_1502 (O_1502,N_14739,N_14713);
or UO_1503 (O_1503,N_14990,N_14948);
nor UO_1504 (O_1504,N_14826,N_14884);
nor UO_1505 (O_1505,N_14760,N_14899);
nor UO_1506 (O_1506,N_14816,N_14960);
nor UO_1507 (O_1507,N_14732,N_14995);
and UO_1508 (O_1508,N_14971,N_14947);
and UO_1509 (O_1509,N_14787,N_14836);
nand UO_1510 (O_1510,N_14712,N_14781);
and UO_1511 (O_1511,N_14942,N_14878);
nor UO_1512 (O_1512,N_14709,N_14810);
or UO_1513 (O_1513,N_14926,N_14788);
xnor UO_1514 (O_1514,N_14764,N_14943);
and UO_1515 (O_1515,N_14875,N_14980);
nand UO_1516 (O_1516,N_14736,N_14773);
and UO_1517 (O_1517,N_14859,N_14734);
and UO_1518 (O_1518,N_14869,N_14946);
xnor UO_1519 (O_1519,N_14869,N_14874);
and UO_1520 (O_1520,N_14882,N_14948);
xnor UO_1521 (O_1521,N_14988,N_14970);
xnor UO_1522 (O_1522,N_14726,N_14810);
and UO_1523 (O_1523,N_14757,N_14895);
nor UO_1524 (O_1524,N_14717,N_14795);
xor UO_1525 (O_1525,N_14979,N_14852);
and UO_1526 (O_1526,N_14961,N_14846);
and UO_1527 (O_1527,N_14769,N_14764);
xor UO_1528 (O_1528,N_14809,N_14989);
nor UO_1529 (O_1529,N_14882,N_14762);
nor UO_1530 (O_1530,N_14932,N_14970);
or UO_1531 (O_1531,N_14875,N_14858);
or UO_1532 (O_1532,N_14781,N_14928);
nor UO_1533 (O_1533,N_14817,N_14908);
and UO_1534 (O_1534,N_14815,N_14990);
or UO_1535 (O_1535,N_14741,N_14723);
nor UO_1536 (O_1536,N_14884,N_14759);
and UO_1537 (O_1537,N_14774,N_14730);
xnor UO_1538 (O_1538,N_14846,N_14715);
xor UO_1539 (O_1539,N_14898,N_14979);
nand UO_1540 (O_1540,N_14783,N_14997);
nand UO_1541 (O_1541,N_14818,N_14946);
or UO_1542 (O_1542,N_14717,N_14722);
and UO_1543 (O_1543,N_14922,N_14878);
nor UO_1544 (O_1544,N_14977,N_14805);
or UO_1545 (O_1545,N_14924,N_14878);
and UO_1546 (O_1546,N_14971,N_14761);
xnor UO_1547 (O_1547,N_14781,N_14951);
nor UO_1548 (O_1548,N_14896,N_14996);
xor UO_1549 (O_1549,N_14790,N_14967);
nand UO_1550 (O_1550,N_14936,N_14943);
xor UO_1551 (O_1551,N_14947,N_14986);
or UO_1552 (O_1552,N_14795,N_14800);
nand UO_1553 (O_1553,N_14811,N_14900);
nor UO_1554 (O_1554,N_14933,N_14972);
or UO_1555 (O_1555,N_14897,N_14869);
and UO_1556 (O_1556,N_14845,N_14775);
nor UO_1557 (O_1557,N_14986,N_14718);
nor UO_1558 (O_1558,N_14802,N_14944);
xnor UO_1559 (O_1559,N_14933,N_14840);
nand UO_1560 (O_1560,N_14919,N_14867);
nand UO_1561 (O_1561,N_14784,N_14897);
or UO_1562 (O_1562,N_14723,N_14866);
or UO_1563 (O_1563,N_14712,N_14908);
or UO_1564 (O_1564,N_14945,N_14957);
nand UO_1565 (O_1565,N_14837,N_14703);
or UO_1566 (O_1566,N_14883,N_14985);
and UO_1567 (O_1567,N_14998,N_14700);
and UO_1568 (O_1568,N_14881,N_14714);
or UO_1569 (O_1569,N_14731,N_14710);
nand UO_1570 (O_1570,N_14966,N_14843);
nor UO_1571 (O_1571,N_14897,N_14905);
or UO_1572 (O_1572,N_14828,N_14785);
nor UO_1573 (O_1573,N_14969,N_14755);
nand UO_1574 (O_1574,N_14871,N_14984);
nor UO_1575 (O_1575,N_14770,N_14998);
nand UO_1576 (O_1576,N_14905,N_14794);
nand UO_1577 (O_1577,N_14770,N_14743);
xnor UO_1578 (O_1578,N_14946,N_14737);
or UO_1579 (O_1579,N_14797,N_14711);
nand UO_1580 (O_1580,N_14880,N_14905);
or UO_1581 (O_1581,N_14780,N_14700);
or UO_1582 (O_1582,N_14900,N_14981);
nor UO_1583 (O_1583,N_14933,N_14918);
nand UO_1584 (O_1584,N_14813,N_14852);
nand UO_1585 (O_1585,N_14947,N_14745);
xor UO_1586 (O_1586,N_14773,N_14791);
xor UO_1587 (O_1587,N_14779,N_14872);
and UO_1588 (O_1588,N_14736,N_14878);
nor UO_1589 (O_1589,N_14985,N_14764);
nand UO_1590 (O_1590,N_14893,N_14938);
and UO_1591 (O_1591,N_14941,N_14718);
xnor UO_1592 (O_1592,N_14834,N_14974);
xnor UO_1593 (O_1593,N_14995,N_14992);
xor UO_1594 (O_1594,N_14969,N_14873);
xor UO_1595 (O_1595,N_14866,N_14837);
nor UO_1596 (O_1596,N_14962,N_14890);
nand UO_1597 (O_1597,N_14808,N_14907);
nor UO_1598 (O_1598,N_14813,N_14884);
and UO_1599 (O_1599,N_14980,N_14818);
or UO_1600 (O_1600,N_14749,N_14821);
nand UO_1601 (O_1601,N_14999,N_14845);
nor UO_1602 (O_1602,N_14742,N_14947);
nor UO_1603 (O_1603,N_14831,N_14893);
nand UO_1604 (O_1604,N_14922,N_14951);
or UO_1605 (O_1605,N_14915,N_14751);
nand UO_1606 (O_1606,N_14703,N_14968);
or UO_1607 (O_1607,N_14743,N_14793);
xnor UO_1608 (O_1608,N_14798,N_14743);
or UO_1609 (O_1609,N_14906,N_14979);
and UO_1610 (O_1610,N_14715,N_14797);
or UO_1611 (O_1611,N_14965,N_14899);
and UO_1612 (O_1612,N_14728,N_14850);
nor UO_1613 (O_1613,N_14980,N_14901);
or UO_1614 (O_1614,N_14981,N_14964);
nand UO_1615 (O_1615,N_14736,N_14949);
xnor UO_1616 (O_1616,N_14938,N_14975);
xnor UO_1617 (O_1617,N_14717,N_14700);
or UO_1618 (O_1618,N_14861,N_14873);
and UO_1619 (O_1619,N_14791,N_14718);
nand UO_1620 (O_1620,N_14850,N_14997);
and UO_1621 (O_1621,N_14884,N_14911);
or UO_1622 (O_1622,N_14922,N_14942);
xnor UO_1623 (O_1623,N_14707,N_14778);
or UO_1624 (O_1624,N_14746,N_14741);
and UO_1625 (O_1625,N_14910,N_14746);
xor UO_1626 (O_1626,N_14972,N_14723);
and UO_1627 (O_1627,N_14730,N_14841);
nand UO_1628 (O_1628,N_14835,N_14783);
or UO_1629 (O_1629,N_14985,N_14751);
nand UO_1630 (O_1630,N_14704,N_14995);
nand UO_1631 (O_1631,N_14837,N_14935);
xor UO_1632 (O_1632,N_14931,N_14813);
or UO_1633 (O_1633,N_14907,N_14853);
or UO_1634 (O_1634,N_14852,N_14843);
xor UO_1635 (O_1635,N_14837,N_14873);
xor UO_1636 (O_1636,N_14811,N_14730);
and UO_1637 (O_1637,N_14817,N_14970);
or UO_1638 (O_1638,N_14845,N_14803);
and UO_1639 (O_1639,N_14837,N_14804);
or UO_1640 (O_1640,N_14820,N_14993);
and UO_1641 (O_1641,N_14930,N_14900);
xor UO_1642 (O_1642,N_14825,N_14956);
nand UO_1643 (O_1643,N_14927,N_14956);
xnor UO_1644 (O_1644,N_14762,N_14800);
xnor UO_1645 (O_1645,N_14805,N_14973);
and UO_1646 (O_1646,N_14989,N_14890);
nand UO_1647 (O_1647,N_14767,N_14842);
nor UO_1648 (O_1648,N_14911,N_14776);
nand UO_1649 (O_1649,N_14930,N_14845);
and UO_1650 (O_1650,N_14705,N_14954);
xor UO_1651 (O_1651,N_14836,N_14910);
or UO_1652 (O_1652,N_14842,N_14999);
nand UO_1653 (O_1653,N_14990,N_14924);
and UO_1654 (O_1654,N_14862,N_14975);
and UO_1655 (O_1655,N_14973,N_14716);
xor UO_1656 (O_1656,N_14882,N_14964);
or UO_1657 (O_1657,N_14802,N_14896);
nor UO_1658 (O_1658,N_14767,N_14713);
nor UO_1659 (O_1659,N_14895,N_14968);
xnor UO_1660 (O_1660,N_14838,N_14941);
nand UO_1661 (O_1661,N_14896,N_14853);
and UO_1662 (O_1662,N_14777,N_14829);
nand UO_1663 (O_1663,N_14889,N_14936);
nand UO_1664 (O_1664,N_14858,N_14905);
nor UO_1665 (O_1665,N_14758,N_14903);
nand UO_1666 (O_1666,N_14827,N_14991);
nand UO_1667 (O_1667,N_14911,N_14718);
nor UO_1668 (O_1668,N_14951,N_14799);
nor UO_1669 (O_1669,N_14792,N_14738);
or UO_1670 (O_1670,N_14900,N_14993);
nand UO_1671 (O_1671,N_14742,N_14921);
nor UO_1672 (O_1672,N_14865,N_14765);
and UO_1673 (O_1673,N_14992,N_14725);
xor UO_1674 (O_1674,N_14811,N_14895);
nand UO_1675 (O_1675,N_14876,N_14734);
nand UO_1676 (O_1676,N_14841,N_14955);
xnor UO_1677 (O_1677,N_14712,N_14793);
nand UO_1678 (O_1678,N_14782,N_14991);
nor UO_1679 (O_1679,N_14932,N_14985);
or UO_1680 (O_1680,N_14773,N_14973);
and UO_1681 (O_1681,N_14927,N_14771);
and UO_1682 (O_1682,N_14839,N_14782);
and UO_1683 (O_1683,N_14799,N_14895);
or UO_1684 (O_1684,N_14955,N_14885);
or UO_1685 (O_1685,N_14909,N_14872);
nand UO_1686 (O_1686,N_14862,N_14870);
and UO_1687 (O_1687,N_14900,N_14939);
or UO_1688 (O_1688,N_14741,N_14739);
nor UO_1689 (O_1689,N_14927,N_14715);
or UO_1690 (O_1690,N_14909,N_14822);
nand UO_1691 (O_1691,N_14727,N_14843);
nand UO_1692 (O_1692,N_14938,N_14819);
nand UO_1693 (O_1693,N_14981,N_14741);
xor UO_1694 (O_1694,N_14721,N_14765);
nor UO_1695 (O_1695,N_14786,N_14956);
or UO_1696 (O_1696,N_14736,N_14749);
xnor UO_1697 (O_1697,N_14905,N_14944);
nand UO_1698 (O_1698,N_14981,N_14888);
and UO_1699 (O_1699,N_14894,N_14939);
and UO_1700 (O_1700,N_14726,N_14965);
and UO_1701 (O_1701,N_14935,N_14969);
nor UO_1702 (O_1702,N_14749,N_14746);
and UO_1703 (O_1703,N_14819,N_14820);
nor UO_1704 (O_1704,N_14760,N_14731);
xnor UO_1705 (O_1705,N_14764,N_14962);
and UO_1706 (O_1706,N_14954,N_14865);
nor UO_1707 (O_1707,N_14887,N_14704);
nor UO_1708 (O_1708,N_14786,N_14755);
xor UO_1709 (O_1709,N_14879,N_14886);
nor UO_1710 (O_1710,N_14882,N_14898);
and UO_1711 (O_1711,N_14842,N_14984);
nand UO_1712 (O_1712,N_14705,N_14809);
or UO_1713 (O_1713,N_14764,N_14745);
xnor UO_1714 (O_1714,N_14977,N_14848);
xor UO_1715 (O_1715,N_14965,N_14761);
xor UO_1716 (O_1716,N_14776,N_14980);
xor UO_1717 (O_1717,N_14949,N_14719);
or UO_1718 (O_1718,N_14833,N_14724);
and UO_1719 (O_1719,N_14748,N_14806);
or UO_1720 (O_1720,N_14951,N_14995);
nand UO_1721 (O_1721,N_14875,N_14913);
xnor UO_1722 (O_1722,N_14785,N_14787);
nand UO_1723 (O_1723,N_14859,N_14712);
xnor UO_1724 (O_1724,N_14942,N_14985);
nand UO_1725 (O_1725,N_14774,N_14773);
nand UO_1726 (O_1726,N_14767,N_14722);
xnor UO_1727 (O_1727,N_14846,N_14879);
or UO_1728 (O_1728,N_14975,N_14768);
nor UO_1729 (O_1729,N_14852,N_14860);
and UO_1730 (O_1730,N_14737,N_14948);
nor UO_1731 (O_1731,N_14977,N_14890);
or UO_1732 (O_1732,N_14788,N_14999);
and UO_1733 (O_1733,N_14728,N_14999);
or UO_1734 (O_1734,N_14870,N_14785);
or UO_1735 (O_1735,N_14737,N_14724);
nand UO_1736 (O_1736,N_14853,N_14815);
nand UO_1737 (O_1737,N_14780,N_14992);
nand UO_1738 (O_1738,N_14700,N_14946);
nor UO_1739 (O_1739,N_14886,N_14715);
nor UO_1740 (O_1740,N_14849,N_14858);
xor UO_1741 (O_1741,N_14721,N_14743);
nor UO_1742 (O_1742,N_14775,N_14768);
nand UO_1743 (O_1743,N_14761,N_14992);
nor UO_1744 (O_1744,N_14701,N_14765);
or UO_1745 (O_1745,N_14749,N_14890);
or UO_1746 (O_1746,N_14773,N_14891);
nor UO_1747 (O_1747,N_14972,N_14911);
or UO_1748 (O_1748,N_14833,N_14866);
nor UO_1749 (O_1749,N_14937,N_14750);
nand UO_1750 (O_1750,N_14957,N_14934);
and UO_1751 (O_1751,N_14858,N_14992);
or UO_1752 (O_1752,N_14752,N_14740);
xor UO_1753 (O_1753,N_14864,N_14773);
or UO_1754 (O_1754,N_14983,N_14855);
and UO_1755 (O_1755,N_14789,N_14946);
nor UO_1756 (O_1756,N_14888,N_14965);
xnor UO_1757 (O_1757,N_14890,N_14999);
and UO_1758 (O_1758,N_14803,N_14862);
or UO_1759 (O_1759,N_14709,N_14884);
xnor UO_1760 (O_1760,N_14952,N_14722);
and UO_1761 (O_1761,N_14706,N_14735);
nand UO_1762 (O_1762,N_14830,N_14739);
or UO_1763 (O_1763,N_14762,N_14921);
and UO_1764 (O_1764,N_14724,N_14868);
and UO_1765 (O_1765,N_14710,N_14907);
xnor UO_1766 (O_1766,N_14839,N_14742);
nor UO_1767 (O_1767,N_14933,N_14852);
and UO_1768 (O_1768,N_14968,N_14877);
and UO_1769 (O_1769,N_14771,N_14766);
xnor UO_1770 (O_1770,N_14974,N_14837);
or UO_1771 (O_1771,N_14922,N_14931);
nor UO_1772 (O_1772,N_14749,N_14721);
and UO_1773 (O_1773,N_14771,N_14862);
and UO_1774 (O_1774,N_14895,N_14831);
or UO_1775 (O_1775,N_14803,N_14960);
and UO_1776 (O_1776,N_14735,N_14856);
nor UO_1777 (O_1777,N_14865,N_14773);
or UO_1778 (O_1778,N_14768,N_14773);
nand UO_1779 (O_1779,N_14804,N_14788);
nand UO_1780 (O_1780,N_14969,N_14917);
nor UO_1781 (O_1781,N_14819,N_14854);
nand UO_1782 (O_1782,N_14837,N_14844);
and UO_1783 (O_1783,N_14707,N_14833);
or UO_1784 (O_1784,N_14882,N_14943);
nor UO_1785 (O_1785,N_14961,N_14869);
or UO_1786 (O_1786,N_14791,N_14730);
nor UO_1787 (O_1787,N_14951,N_14923);
or UO_1788 (O_1788,N_14773,N_14839);
nand UO_1789 (O_1789,N_14706,N_14928);
or UO_1790 (O_1790,N_14811,N_14959);
or UO_1791 (O_1791,N_14816,N_14935);
xnor UO_1792 (O_1792,N_14927,N_14718);
nand UO_1793 (O_1793,N_14937,N_14835);
xnor UO_1794 (O_1794,N_14776,N_14997);
or UO_1795 (O_1795,N_14842,N_14736);
nor UO_1796 (O_1796,N_14844,N_14912);
nor UO_1797 (O_1797,N_14802,N_14786);
nor UO_1798 (O_1798,N_14832,N_14718);
nand UO_1799 (O_1799,N_14776,N_14711);
nand UO_1800 (O_1800,N_14962,N_14816);
xor UO_1801 (O_1801,N_14806,N_14850);
xnor UO_1802 (O_1802,N_14773,N_14731);
nand UO_1803 (O_1803,N_14832,N_14997);
xor UO_1804 (O_1804,N_14798,N_14794);
xnor UO_1805 (O_1805,N_14909,N_14798);
nand UO_1806 (O_1806,N_14709,N_14743);
xor UO_1807 (O_1807,N_14752,N_14779);
nand UO_1808 (O_1808,N_14957,N_14942);
nand UO_1809 (O_1809,N_14984,N_14822);
nand UO_1810 (O_1810,N_14726,N_14940);
xnor UO_1811 (O_1811,N_14839,N_14784);
or UO_1812 (O_1812,N_14883,N_14750);
nor UO_1813 (O_1813,N_14834,N_14815);
nor UO_1814 (O_1814,N_14846,N_14700);
nor UO_1815 (O_1815,N_14944,N_14803);
and UO_1816 (O_1816,N_14798,N_14940);
xor UO_1817 (O_1817,N_14954,N_14887);
or UO_1818 (O_1818,N_14902,N_14916);
or UO_1819 (O_1819,N_14717,N_14770);
and UO_1820 (O_1820,N_14752,N_14769);
xor UO_1821 (O_1821,N_14957,N_14822);
nand UO_1822 (O_1822,N_14702,N_14751);
nor UO_1823 (O_1823,N_14731,N_14965);
xnor UO_1824 (O_1824,N_14781,N_14876);
and UO_1825 (O_1825,N_14853,N_14792);
or UO_1826 (O_1826,N_14719,N_14700);
xnor UO_1827 (O_1827,N_14781,N_14946);
xor UO_1828 (O_1828,N_14709,N_14886);
xnor UO_1829 (O_1829,N_14750,N_14793);
nand UO_1830 (O_1830,N_14766,N_14969);
nand UO_1831 (O_1831,N_14723,N_14934);
nand UO_1832 (O_1832,N_14970,N_14775);
nor UO_1833 (O_1833,N_14967,N_14981);
or UO_1834 (O_1834,N_14940,N_14811);
xor UO_1835 (O_1835,N_14934,N_14787);
and UO_1836 (O_1836,N_14831,N_14787);
or UO_1837 (O_1837,N_14876,N_14901);
and UO_1838 (O_1838,N_14720,N_14778);
nor UO_1839 (O_1839,N_14737,N_14999);
nor UO_1840 (O_1840,N_14983,N_14870);
and UO_1841 (O_1841,N_14922,N_14897);
nand UO_1842 (O_1842,N_14774,N_14747);
nand UO_1843 (O_1843,N_14993,N_14965);
nand UO_1844 (O_1844,N_14991,N_14817);
xnor UO_1845 (O_1845,N_14797,N_14750);
nor UO_1846 (O_1846,N_14713,N_14908);
nand UO_1847 (O_1847,N_14970,N_14934);
nor UO_1848 (O_1848,N_14748,N_14737);
or UO_1849 (O_1849,N_14720,N_14772);
or UO_1850 (O_1850,N_14776,N_14743);
or UO_1851 (O_1851,N_14774,N_14717);
and UO_1852 (O_1852,N_14890,N_14854);
nand UO_1853 (O_1853,N_14804,N_14863);
or UO_1854 (O_1854,N_14834,N_14845);
and UO_1855 (O_1855,N_14794,N_14871);
and UO_1856 (O_1856,N_14960,N_14996);
or UO_1857 (O_1857,N_14754,N_14915);
nor UO_1858 (O_1858,N_14850,N_14821);
nor UO_1859 (O_1859,N_14923,N_14729);
nor UO_1860 (O_1860,N_14873,N_14707);
xor UO_1861 (O_1861,N_14892,N_14988);
nand UO_1862 (O_1862,N_14835,N_14877);
or UO_1863 (O_1863,N_14872,N_14749);
nor UO_1864 (O_1864,N_14769,N_14941);
and UO_1865 (O_1865,N_14939,N_14993);
and UO_1866 (O_1866,N_14780,N_14733);
xor UO_1867 (O_1867,N_14956,N_14975);
nor UO_1868 (O_1868,N_14709,N_14907);
or UO_1869 (O_1869,N_14722,N_14833);
xor UO_1870 (O_1870,N_14770,N_14815);
xor UO_1871 (O_1871,N_14777,N_14969);
and UO_1872 (O_1872,N_14834,N_14830);
xnor UO_1873 (O_1873,N_14856,N_14973);
and UO_1874 (O_1874,N_14753,N_14887);
nand UO_1875 (O_1875,N_14768,N_14786);
nand UO_1876 (O_1876,N_14940,N_14996);
or UO_1877 (O_1877,N_14911,N_14853);
nand UO_1878 (O_1878,N_14705,N_14762);
or UO_1879 (O_1879,N_14809,N_14716);
xnor UO_1880 (O_1880,N_14723,N_14781);
nand UO_1881 (O_1881,N_14954,N_14844);
nor UO_1882 (O_1882,N_14839,N_14929);
or UO_1883 (O_1883,N_14797,N_14700);
xor UO_1884 (O_1884,N_14903,N_14868);
and UO_1885 (O_1885,N_14929,N_14826);
or UO_1886 (O_1886,N_14903,N_14877);
nor UO_1887 (O_1887,N_14968,N_14913);
and UO_1888 (O_1888,N_14716,N_14888);
or UO_1889 (O_1889,N_14968,N_14755);
xor UO_1890 (O_1890,N_14892,N_14709);
xor UO_1891 (O_1891,N_14883,N_14756);
and UO_1892 (O_1892,N_14748,N_14753);
nand UO_1893 (O_1893,N_14845,N_14978);
or UO_1894 (O_1894,N_14960,N_14876);
nand UO_1895 (O_1895,N_14796,N_14966);
or UO_1896 (O_1896,N_14736,N_14989);
xor UO_1897 (O_1897,N_14994,N_14706);
or UO_1898 (O_1898,N_14765,N_14916);
nand UO_1899 (O_1899,N_14860,N_14805);
nor UO_1900 (O_1900,N_14958,N_14790);
nand UO_1901 (O_1901,N_14896,N_14738);
or UO_1902 (O_1902,N_14833,N_14895);
and UO_1903 (O_1903,N_14981,N_14801);
or UO_1904 (O_1904,N_14891,N_14835);
or UO_1905 (O_1905,N_14748,N_14956);
nor UO_1906 (O_1906,N_14743,N_14753);
xor UO_1907 (O_1907,N_14888,N_14723);
xnor UO_1908 (O_1908,N_14779,N_14929);
and UO_1909 (O_1909,N_14885,N_14901);
nand UO_1910 (O_1910,N_14909,N_14983);
and UO_1911 (O_1911,N_14905,N_14841);
and UO_1912 (O_1912,N_14836,N_14890);
and UO_1913 (O_1913,N_14912,N_14721);
xor UO_1914 (O_1914,N_14722,N_14900);
nor UO_1915 (O_1915,N_14977,N_14726);
xor UO_1916 (O_1916,N_14806,N_14929);
nand UO_1917 (O_1917,N_14905,N_14777);
nor UO_1918 (O_1918,N_14790,N_14960);
xnor UO_1919 (O_1919,N_14803,N_14727);
or UO_1920 (O_1920,N_14788,N_14983);
nand UO_1921 (O_1921,N_14918,N_14993);
or UO_1922 (O_1922,N_14761,N_14833);
nand UO_1923 (O_1923,N_14987,N_14938);
nor UO_1924 (O_1924,N_14946,N_14971);
and UO_1925 (O_1925,N_14871,N_14868);
nand UO_1926 (O_1926,N_14701,N_14856);
and UO_1927 (O_1927,N_14801,N_14728);
nand UO_1928 (O_1928,N_14960,N_14895);
nor UO_1929 (O_1929,N_14820,N_14832);
xor UO_1930 (O_1930,N_14752,N_14999);
and UO_1931 (O_1931,N_14804,N_14889);
and UO_1932 (O_1932,N_14969,N_14884);
and UO_1933 (O_1933,N_14748,N_14896);
nand UO_1934 (O_1934,N_14753,N_14841);
nand UO_1935 (O_1935,N_14805,N_14942);
and UO_1936 (O_1936,N_14760,N_14816);
nor UO_1937 (O_1937,N_14873,N_14955);
nor UO_1938 (O_1938,N_14771,N_14936);
or UO_1939 (O_1939,N_14911,N_14861);
nor UO_1940 (O_1940,N_14785,N_14782);
nor UO_1941 (O_1941,N_14790,N_14934);
or UO_1942 (O_1942,N_14861,N_14894);
xor UO_1943 (O_1943,N_14942,N_14712);
or UO_1944 (O_1944,N_14870,N_14724);
nor UO_1945 (O_1945,N_14905,N_14933);
xnor UO_1946 (O_1946,N_14832,N_14874);
nor UO_1947 (O_1947,N_14956,N_14907);
nor UO_1948 (O_1948,N_14741,N_14974);
nor UO_1949 (O_1949,N_14766,N_14879);
xnor UO_1950 (O_1950,N_14983,N_14819);
and UO_1951 (O_1951,N_14791,N_14967);
nor UO_1952 (O_1952,N_14895,N_14763);
xnor UO_1953 (O_1953,N_14789,N_14895);
nor UO_1954 (O_1954,N_14998,N_14902);
nand UO_1955 (O_1955,N_14700,N_14989);
and UO_1956 (O_1956,N_14844,N_14810);
and UO_1957 (O_1957,N_14897,N_14812);
or UO_1958 (O_1958,N_14806,N_14979);
or UO_1959 (O_1959,N_14818,N_14885);
xnor UO_1960 (O_1960,N_14793,N_14832);
xnor UO_1961 (O_1961,N_14894,N_14914);
nand UO_1962 (O_1962,N_14813,N_14845);
nand UO_1963 (O_1963,N_14943,N_14982);
or UO_1964 (O_1964,N_14959,N_14796);
nand UO_1965 (O_1965,N_14852,N_14921);
or UO_1966 (O_1966,N_14784,N_14795);
nand UO_1967 (O_1967,N_14945,N_14999);
xor UO_1968 (O_1968,N_14980,N_14706);
nand UO_1969 (O_1969,N_14816,N_14771);
and UO_1970 (O_1970,N_14867,N_14944);
or UO_1971 (O_1971,N_14781,N_14849);
xor UO_1972 (O_1972,N_14843,N_14823);
or UO_1973 (O_1973,N_14830,N_14710);
or UO_1974 (O_1974,N_14947,N_14707);
nand UO_1975 (O_1975,N_14739,N_14766);
xnor UO_1976 (O_1976,N_14908,N_14959);
or UO_1977 (O_1977,N_14884,N_14835);
and UO_1978 (O_1978,N_14963,N_14786);
and UO_1979 (O_1979,N_14750,N_14843);
nand UO_1980 (O_1980,N_14993,N_14714);
and UO_1981 (O_1981,N_14770,N_14879);
nor UO_1982 (O_1982,N_14918,N_14923);
nor UO_1983 (O_1983,N_14876,N_14741);
and UO_1984 (O_1984,N_14764,N_14895);
nand UO_1985 (O_1985,N_14843,N_14904);
and UO_1986 (O_1986,N_14844,N_14972);
and UO_1987 (O_1987,N_14875,N_14999);
xnor UO_1988 (O_1988,N_14991,N_14749);
nand UO_1989 (O_1989,N_14857,N_14835);
and UO_1990 (O_1990,N_14834,N_14728);
and UO_1991 (O_1991,N_14700,N_14821);
or UO_1992 (O_1992,N_14873,N_14890);
or UO_1993 (O_1993,N_14849,N_14950);
nor UO_1994 (O_1994,N_14841,N_14785);
or UO_1995 (O_1995,N_14934,N_14844);
or UO_1996 (O_1996,N_14973,N_14820);
xnor UO_1997 (O_1997,N_14703,N_14974);
nor UO_1998 (O_1998,N_14726,N_14728);
nor UO_1999 (O_1999,N_14734,N_14760);
endmodule