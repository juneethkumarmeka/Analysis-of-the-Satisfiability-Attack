module basic_750_5000_1000_2_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2506,N_2507,N_2509,N_2510,N_2511,N_2512,N_2514,N_2515,N_2516,N_2517,N_2518,N_2521,N_2522,N_2523,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2540,N_2541,N_2542,N_2544,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2560,N_2561,N_2562,N_2563,N_2564,N_2566,N_2568,N_2569,N_2572,N_2573,N_2574,N_2577,N_2578,N_2579,N_2580,N_2581,N_2584,N_2586,N_2590,N_2593,N_2595,N_2596,N_2597,N_2598,N_2599,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2634,N_2635,N_2636,N_2637,N_2641,N_2642,N_2643,N_2645,N_2647,N_2650,N_2651,N_2652,N_2653,N_2654,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2680,N_2682,N_2684,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2696,N_2697,N_2699,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2725,N_2726,N_2728,N_2729,N_2730,N_2731,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2751,N_2752,N_2753,N_2754,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2783,N_2784,N_2785,N_2787,N_2788,N_2789,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2804,N_2805,N_2806,N_2807,N_2809,N_2810,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2827,N_2828,N_2829,N_2830,N_2831,N_2833,N_2834,N_2836,N_2837,N_2838,N_2839,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2861,N_2862,N_2863,N_2865,N_2866,N_2867,N_2869,N_2870,N_2871,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2893,N_2896,N_2897,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2908,N_2909,N_2910,N_2911,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2923,N_2924,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2939,N_2940,N_2941,N_2943,N_2944,N_2946,N_2947,N_2949,N_2951,N_2952,N_2953,N_2954,N_2955,N_2957,N_2958,N_2960,N_2962,N_2963,N_2964,N_2965,N_2966,N_2968,N_2969,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2992,N_2993,N_2994,N_2995,N_2997,N_2998,N_2999,N_3001,N_3002,N_3004,N_3005,N_3006,N_3007,N_3009,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3024,N_3026,N_3027,N_3029,N_3031,N_3032,N_3034,N_3037,N_3038,N_3040,N_3042,N_3043,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3079,N_3080,N_3081,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3090,N_3091,N_3093,N_3094,N_3095,N_3096,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3154,N_3155,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3186,N_3187,N_3189,N_3190,N_3191,N_3192,N_3193,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3217,N_3218,N_3219,N_3221,N_3222,N_3223,N_3224,N_3225,N_3227,N_3228,N_3229,N_3232,N_3233,N_3234,N_3236,N_3237,N_3238,N_3239,N_3240,N_3242,N_3243,N_3245,N_3247,N_3248,N_3249,N_3250,N_3252,N_3254,N_3256,N_3257,N_3258,N_3259,N_3260,N_3262,N_3264,N_3265,N_3266,N_3268,N_3269,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3279,N_3280,N_3281,N_3282,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3295,N_3296,N_3297,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3307,N_3308,N_3309,N_3311,N_3315,N_3316,N_3317,N_3319,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3361,N_3362,N_3363,N_3364,N_3365,N_3367,N_3368,N_3370,N_3371,N_3372,N_3373,N_3374,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3384,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3395,N_3396,N_3397,N_3398,N_3400,N_3401,N_3402,N_3403,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3417,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3459,N_3460,N_3461,N_3462,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3476,N_3477,N_3479,N_3480,N_3481,N_3482,N_3483,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3494,N_3495,N_3496,N_3497,N_3498,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3524,N_3525,N_3526,N_3527,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3560,N_3563,N_3565,N_3567,N_3568,N_3569,N_3570,N_3572,N_3573,N_3575,N_3577,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3604,N_3605,N_3606,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3623,N_3624,N_3625,N_3626,N_3627,N_3629,N_3632,N_3633,N_3635,N_3636,N_3637,N_3639,N_3640,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3661,N_3662,N_3664,N_3665,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3682,N_3683,N_3684,N_3686,N_3687,N_3688,N_3689,N_3691,N_3692,N_3694,N_3695,N_3696,N_3697,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3729,N_3731,N_3733,N_3734,N_3735,N_3738,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3759,N_3760,N_3762,N_3763,N_3765,N_3766,N_3767,N_3768,N_3769,N_3771,N_3772,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3782,N_3783,N_3785,N_3786,N_3788,N_3789,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3813,N_3815,N_3816,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3846,N_3847,N_3848,N_3849,N_3850,N_3852,N_3853,N_3854,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3885,N_3886,N_3887,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3908,N_3909,N_3910,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3928,N_3929,N_3930,N_3931,N_3933,N_3934,N_3935,N_3936,N_3937,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3969,N_3970,N_3974,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3983,N_3984,N_3985,N_3986,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4005,N_4006,N_4007,N_4009,N_4010,N_4011,N_4012,N_4013,N_4015,N_4016,N_4017,N_4018,N_4019,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4028,N_4030,N_4032,N_4033,N_4035,N_4036,N_4037,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4049,N_4050,N_4051,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4060,N_4062,N_4063,N_4064,N_4065,N_4066,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4078,N_4079,N_4080,N_4081,N_4083,N_4085,N_4087,N_4088,N_4090,N_4093,N_4094,N_4096,N_4097,N_4100,N_4101,N_4102,N_4104,N_4105,N_4106,N_4108,N_4109,N_4111,N_4113,N_4114,N_4115,N_4116,N_4117,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4129,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4141,N_4142,N_4144,N_4147,N_4148,N_4150,N_4152,N_4153,N_4155,N_4157,N_4159,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4173,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4187,N_4189,N_4190,N_4191,N_4192,N_4195,N_4196,N_4197,N_4198,N_4199,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4221,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4239,N_4240,N_4243,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4255,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4265,N_4266,N_4267,N_4269,N_4270,N_4271,N_4274,N_4275,N_4276,N_4279,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4296,N_4298,N_4299,N_4300,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4324,N_4325,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4365,N_4367,N_4368,N_4369,N_4372,N_4373,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4397,N_4398,N_4399,N_4400,N_4402,N_4403,N_4404,N_4407,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4422,N_4424,N_4425,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4434,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4455,N_4456,N_4457,N_4458,N_4459,N_4461,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4471,N_4472,N_4473,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4495,N_4496,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4524,N_4526,N_4527,N_4528,N_4530,N_4531,N_4532,N_4533,N_4534,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4567,N_4568,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4579,N_4582,N_4583,N_4584,N_4585,N_4587,N_4588,N_4591,N_4592,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4632,N_4633,N_4634,N_4635,N_4636,N_4638,N_4640,N_4641,N_4642,N_4644,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4669,N_4670,N_4672,N_4673,N_4675,N_4677,N_4678,N_4679,N_4681,N_4684,N_4685,N_4686,N_4688,N_4689,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4707,N_4709,N_4711,N_4713,N_4715,N_4716,N_4717,N_4718,N_4719,N_4721,N_4722,N_4726,N_4727,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4742,N_4745,N_4746,N_4747,N_4748,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4764,N_4766,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4780,N_4781,N_4782,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4811,N_4812,N_4813,N_4814,N_4815,N_4817,N_4818,N_4820,N_4821,N_4823,N_4824,N_4825,N_4826,N_4828,N_4829,N_4831,N_4832,N_4833,N_4834,N_4835,N_4837,N_4838,N_4839,N_4840,N_4842,N_4843,N_4844,N_4845,N_4847,N_4849,N_4850,N_4852,N_4854,N_4855,N_4857,N_4858,N_4861,N_4862,N_4863,N_4864,N_4866,N_4867,N_4868,N_4869,N_4870,N_4873,N_4874,N_4875,N_4877,N_4878,N_4879,N_4880,N_4881,N_4884,N_4885,N_4887,N_4888,N_4891,N_4893,N_4895,N_4896,N_4898,N_4900,N_4901,N_4902,N_4903,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4913,N_4914,N_4916,N_4917,N_4918,N_4919,N_4921,N_4922,N_4923,N_4926,N_4927,N_4928,N_4932,N_4934,N_4935,N_4936,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4971,N_4972,N_4973,N_4975,N_4976,N_4977,N_4978,N_4980,N_4981,N_4983,N_4985,N_4986,N_4987,N_4988,N_4989,N_4991,N_4992,N_4993,N_4995,N_4996,N_4997,N_4999;
or U0 (N_0,In_289,In_440);
or U1 (N_1,In_14,In_324);
and U2 (N_2,In_633,In_412);
nor U3 (N_3,In_330,In_479);
nand U4 (N_4,In_271,In_32);
nand U5 (N_5,In_735,In_681);
and U6 (N_6,In_409,In_588);
and U7 (N_7,In_403,In_127);
nand U8 (N_8,In_590,In_407);
nand U9 (N_9,In_11,In_653);
nand U10 (N_10,In_656,In_564);
or U11 (N_11,In_577,In_138);
or U12 (N_12,In_563,In_291);
and U13 (N_13,In_628,In_185);
or U14 (N_14,In_355,In_511);
and U15 (N_15,In_370,In_31);
and U16 (N_16,In_384,In_367);
nor U17 (N_17,In_210,In_642);
or U18 (N_18,In_531,In_639);
and U19 (N_19,In_659,In_416);
nand U20 (N_20,In_418,In_431);
or U21 (N_21,In_557,In_448);
or U22 (N_22,In_313,In_264);
nand U23 (N_23,In_13,In_177);
and U24 (N_24,In_404,In_619);
nor U25 (N_25,In_231,In_405);
and U26 (N_26,In_273,In_342);
or U27 (N_27,In_631,In_368);
or U28 (N_28,In_636,In_28);
and U29 (N_29,In_234,In_39);
nand U30 (N_30,In_422,In_574);
and U31 (N_31,In_423,In_3);
and U32 (N_32,In_190,In_340);
or U33 (N_33,In_721,In_672);
or U34 (N_34,In_453,In_372);
xnor U35 (N_35,In_595,In_237);
or U36 (N_36,In_576,In_283);
xor U37 (N_37,In_94,In_137);
nor U38 (N_38,In_5,In_575);
nand U39 (N_39,In_529,In_321);
nor U40 (N_40,In_284,In_637);
nor U41 (N_41,In_720,In_366);
and U42 (N_42,In_38,In_295);
and U43 (N_43,In_105,In_186);
xnor U44 (N_44,In_692,In_430);
nor U45 (N_45,In_740,In_21);
or U46 (N_46,In_374,In_654);
or U47 (N_47,In_40,In_360);
nand U48 (N_48,In_157,In_322);
xor U49 (N_49,In_4,In_457);
nand U50 (N_50,In_468,In_382);
and U51 (N_51,In_334,In_358);
and U52 (N_52,In_81,In_79);
nor U53 (N_53,In_523,In_163);
and U54 (N_54,In_172,In_558);
nor U55 (N_55,In_108,In_580);
and U56 (N_56,In_547,In_287);
and U57 (N_57,In_196,In_215);
or U58 (N_58,In_184,In_128);
nand U59 (N_59,In_549,In_189);
xnor U60 (N_60,In_476,In_593);
nand U61 (N_61,In_98,In_438);
nand U62 (N_62,In_679,In_710);
nor U63 (N_63,In_256,In_59);
nand U64 (N_64,In_408,In_655);
or U65 (N_65,In_22,In_327);
or U66 (N_66,In_214,In_492);
nand U67 (N_67,In_222,In_677);
or U68 (N_68,In_369,In_265);
nor U69 (N_69,In_71,In_160);
nor U70 (N_70,In_396,In_116);
nor U71 (N_71,In_598,In_542);
xnor U72 (N_72,In_742,In_717);
or U73 (N_73,In_586,In_326);
xor U74 (N_74,In_281,In_130);
and U75 (N_75,In_669,In_122);
nor U76 (N_76,In_125,In_725);
or U77 (N_77,In_65,In_341);
and U78 (N_78,In_401,In_18);
and U79 (N_79,In_345,In_303);
nand U80 (N_80,In_695,In_319);
and U81 (N_81,In_191,In_743);
nor U82 (N_82,In_121,In_395);
nand U83 (N_83,In_516,In_328);
nor U84 (N_84,In_51,In_607);
nand U85 (N_85,In_419,In_736);
nand U86 (N_86,In_302,In_131);
xor U87 (N_87,In_635,In_166);
nor U88 (N_88,In_584,In_24);
and U89 (N_89,In_386,In_392);
nand U90 (N_90,In_182,In_680);
nor U91 (N_91,In_747,In_627);
nand U92 (N_92,In_318,In_701);
or U93 (N_93,In_739,In_316);
or U94 (N_94,In_618,In_169);
or U95 (N_95,In_728,In_670);
and U96 (N_96,In_745,In_652);
nor U97 (N_97,In_266,In_624);
nand U98 (N_98,In_645,In_535);
nand U99 (N_99,In_371,In_428);
nor U100 (N_100,In_662,In_391);
nor U101 (N_101,In_362,In_47);
nand U102 (N_102,In_238,In_582);
or U103 (N_103,In_246,In_605);
and U104 (N_104,In_640,In_146);
or U105 (N_105,In_211,In_718);
or U106 (N_106,In_178,In_276);
and U107 (N_107,In_99,In_550);
nand U108 (N_108,In_651,In_235);
and U109 (N_109,In_195,In_219);
nor U110 (N_110,In_16,In_429);
nor U111 (N_111,In_676,In_614);
and U112 (N_112,In_375,In_171);
nand U113 (N_113,In_427,In_152);
nand U114 (N_114,In_441,In_241);
nand U115 (N_115,In_696,In_749);
xor U116 (N_116,In_602,In_707);
nor U117 (N_117,In_539,In_63);
nor U118 (N_118,In_376,In_481);
nand U119 (N_119,In_26,In_27);
nand U120 (N_120,In_261,In_338);
xnor U121 (N_121,In_229,In_57);
nor U122 (N_122,In_454,In_363);
or U123 (N_123,In_364,In_228);
nand U124 (N_124,In_650,In_450);
or U125 (N_125,In_119,In_278);
or U126 (N_126,In_458,In_432);
nand U127 (N_127,In_548,In_33);
nand U128 (N_128,In_232,In_393);
or U129 (N_129,In_663,In_120);
nor U130 (N_130,In_236,In_459);
and U131 (N_131,In_583,In_144);
nor U132 (N_132,In_660,In_478);
nor U133 (N_133,In_630,In_310);
nor U134 (N_134,In_339,In_356);
nor U135 (N_135,In_462,In_361);
xor U136 (N_136,In_202,In_686);
and U137 (N_137,In_267,In_561);
and U138 (N_138,In_684,In_19);
and U139 (N_139,In_406,In_713);
nor U140 (N_140,In_571,In_198);
or U141 (N_141,In_534,In_259);
nor U142 (N_142,In_666,In_45);
nand U143 (N_143,In_390,In_248);
nor U144 (N_144,In_139,In_43);
and U145 (N_145,In_496,In_451);
nor U146 (N_146,In_413,In_223);
nand U147 (N_147,In_294,In_601);
nand U148 (N_148,In_230,In_77);
or U149 (N_149,In_88,In_251);
and U150 (N_150,In_307,In_110);
and U151 (N_151,In_102,In_293);
xnor U152 (N_152,In_277,In_336);
xor U153 (N_153,In_709,In_734);
nand U154 (N_154,In_134,In_722);
or U155 (N_155,In_8,In_425);
xnor U156 (N_156,In_398,In_305);
and U157 (N_157,In_387,In_299);
and U158 (N_158,In_648,In_506);
nand U159 (N_159,In_337,In_643);
and U160 (N_160,In_86,In_187);
nand U161 (N_161,In_56,In_50);
or U162 (N_162,In_262,In_73);
and U163 (N_163,In_80,In_510);
and U164 (N_164,In_706,In_694);
nand U165 (N_165,In_472,In_301);
nand U166 (N_166,In_426,In_239);
or U167 (N_167,In_572,In_221);
xor U168 (N_168,In_194,In_181);
and U169 (N_169,In_17,In_167);
and U170 (N_170,In_66,In_617);
nor U171 (N_171,In_84,In_348);
nor U172 (N_172,In_592,In_480);
nor U173 (N_173,In_179,In_104);
nand U174 (N_174,In_585,In_206);
nand U175 (N_175,In_490,In_514);
nor U176 (N_176,In_70,In_646);
and U177 (N_177,In_526,In_591);
nand U178 (N_178,In_55,In_447);
nor U179 (N_179,In_442,In_699);
and U180 (N_180,In_533,In_200);
nor U181 (N_181,In_520,In_380);
xor U182 (N_182,In_0,In_29);
or U183 (N_183,In_275,In_383);
or U184 (N_184,In_668,In_304);
or U185 (N_185,In_288,In_209);
nor U186 (N_186,In_300,In_46);
nor U187 (N_187,In_483,In_544);
nand U188 (N_188,In_164,In_675);
nand U189 (N_189,In_554,In_467);
and U190 (N_190,In_292,In_297);
nand U191 (N_191,In_60,In_68);
or U192 (N_192,In_159,In_715);
nor U193 (N_193,In_233,In_101);
nand U194 (N_194,In_353,In_314);
nand U195 (N_195,In_258,In_91);
nand U196 (N_196,In_445,In_723);
xor U197 (N_197,In_664,In_513);
nand U198 (N_198,In_205,In_638);
and U199 (N_199,In_192,In_578);
nor U200 (N_200,In_90,In_133);
and U201 (N_201,In_589,In_42);
nand U202 (N_202,In_626,In_731);
nand U203 (N_203,In_702,In_474);
nor U204 (N_204,In_201,In_711);
or U205 (N_205,In_242,In_629);
and U206 (N_206,In_329,In_568);
or U207 (N_207,In_397,In_746);
nor U208 (N_208,In_37,In_315);
nand U209 (N_209,In_213,In_693);
and U210 (N_210,In_488,In_106);
nor U211 (N_211,In_323,In_6);
nor U212 (N_212,In_553,In_730);
nand U213 (N_213,In_269,In_143);
nand U214 (N_214,In_671,In_15);
xor U215 (N_215,In_455,In_683);
xnor U216 (N_216,In_688,In_325);
nand U217 (N_217,In_97,In_597);
and U218 (N_218,In_124,In_446);
nor U219 (N_219,In_537,In_527);
nand U220 (N_220,In_486,In_359);
and U221 (N_221,In_20,In_344);
and U222 (N_222,In_142,In_286);
nor U223 (N_223,In_562,In_744);
and U224 (N_224,In_117,In_543);
nor U225 (N_225,In_417,In_611);
nand U226 (N_226,In_503,In_647);
nor U227 (N_227,In_243,In_487);
nand U228 (N_228,In_320,In_599);
nor U229 (N_229,In_260,In_477);
nor U230 (N_230,In_25,In_634);
nand U231 (N_231,In_30,In_115);
nor U232 (N_232,In_674,In_298);
or U233 (N_233,In_249,In_161);
nor U234 (N_234,In_714,In_697);
nand U235 (N_235,In_312,In_193);
or U236 (N_236,In_493,In_600);
nand U237 (N_237,In_257,In_389);
nor U238 (N_238,In_464,In_421);
nand U239 (N_239,In_10,In_690);
nand U240 (N_240,In_498,In_625);
or U241 (N_241,In_489,In_140);
or U242 (N_242,In_402,In_69);
nor U243 (N_243,In_644,In_536);
nor U244 (N_244,In_606,In_1);
or U245 (N_245,In_373,In_36);
or U246 (N_246,In_180,In_162);
nor U247 (N_247,In_308,In_311);
nor U248 (N_248,In_354,In_658);
or U249 (N_249,In_118,In_204);
nand U250 (N_250,In_461,In_279);
or U251 (N_251,In_158,In_150);
nor U252 (N_252,In_515,In_377);
or U253 (N_253,In_7,In_136);
nor U254 (N_254,In_726,In_518);
and U255 (N_255,In_424,In_132);
nor U256 (N_256,In_85,In_224);
and U257 (N_257,In_466,In_296);
xnor U258 (N_258,In_532,In_456);
or U259 (N_259,In_525,In_175);
and U260 (N_260,In_443,In_176);
xnor U261 (N_261,In_556,In_545);
xor U262 (N_262,In_705,In_280);
nand U263 (N_263,In_34,In_351);
and U264 (N_264,In_112,In_449);
nor U265 (N_265,In_485,In_306);
and U266 (N_266,In_35,In_399);
or U267 (N_267,In_569,In_673);
and U268 (N_268,In_517,In_203);
nand U269 (N_269,In_82,In_507);
xor U270 (N_270,In_540,In_126);
or U271 (N_271,In_49,In_103);
or U272 (N_272,In_565,In_667);
nor U273 (N_273,In_567,In_622);
or U274 (N_274,In_212,In_352);
nor U275 (N_275,In_420,In_560);
or U276 (N_276,In_641,In_350);
or U277 (N_277,In_75,In_74);
or U278 (N_278,In_64,In_632);
and U279 (N_279,In_551,In_388);
nor U280 (N_280,In_147,In_471);
nand U281 (N_281,In_685,In_207);
or U282 (N_282,In_538,In_9);
nor U283 (N_283,In_712,In_621);
xor U284 (N_284,In_436,In_48);
nand U285 (N_285,In_623,In_244);
or U286 (N_286,In_522,In_252);
and U287 (N_287,In_521,In_145);
nor U288 (N_288,In_724,In_444);
nand U289 (N_289,In_379,In_581);
nand U290 (N_290,In_2,In_620);
nor U291 (N_291,In_197,In_394);
xor U292 (N_292,In_733,In_411);
xor U293 (N_293,In_689,In_217);
or U294 (N_294,In_335,In_12);
and U295 (N_295,In_729,In_665);
nand U296 (N_296,In_439,In_470);
nor U297 (N_297,In_255,In_410);
and U298 (N_298,In_272,In_437);
and U299 (N_299,In_153,In_381);
or U300 (N_300,In_41,In_62);
nand U301 (N_301,In_400,In_89);
or U302 (N_302,In_52,In_528);
xor U303 (N_303,In_156,In_151);
nand U304 (N_304,In_282,In_469);
nand U305 (N_305,In_495,In_331);
nor U306 (N_306,In_727,In_475);
nor U307 (N_307,In_433,In_220);
nor U308 (N_308,In_748,In_290);
and U309 (N_309,In_499,In_378);
or U310 (N_310,In_107,In_512);
and U311 (N_311,In_704,In_473);
nor U312 (N_312,In_247,In_716);
nor U313 (N_313,In_268,In_208);
xnor U314 (N_314,In_682,In_505);
nand U315 (N_315,In_155,In_309);
nor U316 (N_316,In_657,In_678);
xor U317 (N_317,In_415,In_123);
xnor U318 (N_318,In_649,In_460);
nor U319 (N_319,In_225,In_732);
nor U320 (N_320,In_465,In_226);
or U321 (N_321,In_559,In_509);
nand U322 (N_322,In_87,In_504);
nand U323 (N_323,In_174,In_566);
nand U324 (N_324,In_508,In_741);
nand U325 (N_325,In_170,In_719);
and U326 (N_326,In_141,In_414);
nand U327 (N_327,In_154,In_491);
nor U328 (N_328,In_698,In_183);
or U329 (N_329,In_113,In_218);
nor U330 (N_330,In_608,In_609);
and U331 (N_331,In_285,In_546);
nor U332 (N_332,In_93,In_61);
nand U333 (N_333,In_435,In_365);
or U334 (N_334,In_579,In_519);
and U335 (N_335,In_594,In_168);
nand U336 (N_336,In_501,In_253);
or U337 (N_337,In_603,In_541);
or U338 (N_338,In_114,In_72);
xnor U339 (N_339,In_199,In_165);
and U340 (N_340,In_343,In_83);
or U341 (N_341,In_661,In_612);
and U342 (N_342,In_227,In_482);
or U343 (N_343,In_708,In_100);
and U344 (N_344,In_616,In_691);
nand U345 (N_345,In_317,In_95);
and U346 (N_346,In_737,In_349);
nand U347 (N_347,In_129,In_385);
and U348 (N_348,In_500,In_703);
or U349 (N_349,In_135,In_332);
nand U350 (N_350,In_615,In_552);
or U351 (N_351,In_587,In_263);
and U352 (N_352,In_76,In_687);
nor U353 (N_353,In_44,In_254);
nor U354 (N_354,In_53,In_452);
nand U355 (N_355,In_58,In_54);
nand U356 (N_356,In_573,In_610);
nor U357 (N_357,In_524,In_270);
and U358 (N_358,In_604,In_216);
or U359 (N_359,In_596,In_570);
nor U360 (N_360,In_555,In_484);
nor U361 (N_361,In_78,In_96);
and U362 (N_362,In_333,In_613);
and U363 (N_363,In_173,In_23);
or U364 (N_364,In_67,In_700);
or U365 (N_365,In_109,In_148);
and U366 (N_366,In_111,In_274);
and U367 (N_367,In_347,In_92);
and U368 (N_368,In_530,In_240);
or U369 (N_369,In_245,In_149);
or U370 (N_370,In_434,In_188);
and U371 (N_371,In_494,In_738);
and U372 (N_372,In_346,In_463);
xor U373 (N_373,In_497,In_357);
or U374 (N_374,In_502,In_250);
nand U375 (N_375,In_714,In_286);
nand U376 (N_376,In_440,In_624);
or U377 (N_377,In_546,In_60);
or U378 (N_378,In_748,In_607);
or U379 (N_379,In_655,In_24);
xor U380 (N_380,In_264,In_281);
or U381 (N_381,In_344,In_123);
and U382 (N_382,In_574,In_16);
and U383 (N_383,In_229,In_221);
and U384 (N_384,In_188,In_645);
or U385 (N_385,In_428,In_159);
or U386 (N_386,In_61,In_228);
xor U387 (N_387,In_348,In_613);
nand U388 (N_388,In_555,In_318);
or U389 (N_389,In_705,In_58);
nand U390 (N_390,In_207,In_748);
nor U391 (N_391,In_538,In_562);
nor U392 (N_392,In_720,In_224);
and U393 (N_393,In_210,In_659);
nand U394 (N_394,In_702,In_705);
nand U395 (N_395,In_300,In_42);
nor U396 (N_396,In_385,In_196);
xor U397 (N_397,In_181,In_574);
nor U398 (N_398,In_413,In_350);
and U399 (N_399,In_250,In_272);
or U400 (N_400,In_434,In_75);
nand U401 (N_401,In_744,In_151);
nand U402 (N_402,In_604,In_79);
and U403 (N_403,In_30,In_449);
or U404 (N_404,In_697,In_702);
or U405 (N_405,In_60,In_623);
nand U406 (N_406,In_375,In_170);
and U407 (N_407,In_256,In_83);
and U408 (N_408,In_246,In_170);
or U409 (N_409,In_293,In_664);
xor U410 (N_410,In_390,In_14);
nand U411 (N_411,In_137,In_66);
or U412 (N_412,In_445,In_538);
and U413 (N_413,In_549,In_419);
or U414 (N_414,In_293,In_53);
nor U415 (N_415,In_376,In_101);
or U416 (N_416,In_666,In_537);
nor U417 (N_417,In_476,In_729);
nand U418 (N_418,In_53,In_157);
or U419 (N_419,In_414,In_611);
nor U420 (N_420,In_186,In_337);
nor U421 (N_421,In_498,In_486);
nor U422 (N_422,In_124,In_245);
and U423 (N_423,In_235,In_485);
and U424 (N_424,In_508,In_78);
nor U425 (N_425,In_456,In_707);
and U426 (N_426,In_275,In_387);
and U427 (N_427,In_421,In_711);
nand U428 (N_428,In_245,In_744);
and U429 (N_429,In_328,In_210);
xor U430 (N_430,In_90,In_333);
nand U431 (N_431,In_39,In_38);
or U432 (N_432,In_264,In_350);
xor U433 (N_433,In_208,In_480);
and U434 (N_434,In_278,In_531);
or U435 (N_435,In_382,In_166);
or U436 (N_436,In_534,In_403);
and U437 (N_437,In_300,In_183);
and U438 (N_438,In_726,In_687);
nor U439 (N_439,In_591,In_236);
or U440 (N_440,In_586,In_392);
or U441 (N_441,In_130,In_237);
nand U442 (N_442,In_688,In_266);
or U443 (N_443,In_63,In_35);
nand U444 (N_444,In_74,In_285);
and U445 (N_445,In_243,In_139);
or U446 (N_446,In_418,In_704);
or U447 (N_447,In_71,In_242);
nand U448 (N_448,In_518,In_247);
nand U449 (N_449,In_672,In_338);
or U450 (N_450,In_382,In_28);
nand U451 (N_451,In_111,In_397);
or U452 (N_452,In_482,In_577);
or U453 (N_453,In_516,In_719);
and U454 (N_454,In_86,In_705);
nor U455 (N_455,In_19,In_235);
or U456 (N_456,In_383,In_17);
nand U457 (N_457,In_505,In_68);
or U458 (N_458,In_522,In_455);
nor U459 (N_459,In_503,In_269);
and U460 (N_460,In_466,In_254);
and U461 (N_461,In_186,In_287);
nand U462 (N_462,In_244,In_577);
nand U463 (N_463,In_67,In_455);
nor U464 (N_464,In_174,In_335);
nor U465 (N_465,In_504,In_337);
and U466 (N_466,In_183,In_525);
and U467 (N_467,In_709,In_600);
or U468 (N_468,In_207,In_68);
and U469 (N_469,In_585,In_360);
and U470 (N_470,In_399,In_74);
or U471 (N_471,In_208,In_342);
nand U472 (N_472,In_658,In_544);
or U473 (N_473,In_285,In_343);
or U474 (N_474,In_518,In_20);
nor U475 (N_475,In_738,In_727);
nor U476 (N_476,In_49,In_309);
and U477 (N_477,In_141,In_584);
or U478 (N_478,In_104,In_708);
and U479 (N_479,In_515,In_567);
or U480 (N_480,In_687,In_91);
or U481 (N_481,In_0,In_532);
nand U482 (N_482,In_689,In_368);
or U483 (N_483,In_565,In_183);
nand U484 (N_484,In_671,In_4);
nand U485 (N_485,In_357,In_94);
nor U486 (N_486,In_486,In_434);
and U487 (N_487,In_367,In_355);
nor U488 (N_488,In_734,In_24);
or U489 (N_489,In_587,In_663);
and U490 (N_490,In_235,In_441);
and U491 (N_491,In_412,In_106);
and U492 (N_492,In_346,In_649);
xnor U493 (N_493,In_564,In_16);
and U494 (N_494,In_441,In_648);
or U495 (N_495,In_560,In_700);
nor U496 (N_496,In_624,In_116);
and U497 (N_497,In_204,In_658);
and U498 (N_498,In_707,In_518);
nand U499 (N_499,In_624,In_658);
nand U500 (N_500,In_732,In_496);
nor U501 (N_501,In_84,In_420);
or U502 (N_502,In_168,In_731);
nor U503 (N_503,In_410,In_349);
nor U504 (N_504,In_662,In_706);
or U505 (N_505,In_232,In_70);
nor U506 (N_506,In_308,In_114);
and U507 (N_507,In_64,In_551);
nand U508 (N_508,In_85,In_17);
and U509 (N_509,In_443,In_677);
nand U510 (N_510,In_62,In_302);
nand U511 (N_511,In_742,In_179);
or U512 (N_512,In_20,In_330);
nand U513 (N_513,In_558,In_234);
and U514 (N_514,In_654,In_211);
and U515 (N_515,In_89,In_260);
nor U516 (N_516,In_688,In_733);
and U517 (N_517,In_625,In_693);
and U518 (N_518,In_453,In_550);
nor U519 (N_519,In_229,In_464);
or U520 (N_520,In_182,In_30);
or U521 (N_521,In_176,In_326);
and U522 (N_522,In_562,In_115);
xor U523 (N_523,In_468,In_680);
xor U524 (N_524,In_229,In_8);
nor U525 (N_525,In_362,In_74);
nand U526 (N_526,In_218,In_468);
or U527 (N_527,In_227,In_609);
nor U528 (N_528,In_123,In_140);
xor U529 (N_529,In_201,In_127);
nand U530 (N_530,In_502,In_3);
nor U531 (N_531,In_203,In_205);
and U532 (N_532,In_220,In_267);
and U533 (N_533,In_438,In_384);
and U534 (N_534,In_567,In_14);
and U535 (N_535,In_504,In_286);
or U536 (N_536,In_404,In_606);
or U537 (N_537,In_478,In_256);
nor U538 (N_538,In_309,In_552);
xnor U539 (N_539,In_375,In_24);
or U540 (N_540,In_617,In_253);
nor U541 (N_541,In_0,In_692);
nand U542 (N_542,In_2,In_541);
or U543 (N_543,In_440,In_352);
nor U544 (N_544,In_677,In_192);
nand U545 (N_545,In_302,In_87);
nand U546 (N_546,In_403,In_366);
nand U547 (N_547,In_16,In_397);
or U548 (N_548,In_457,In_434);
or U549 (N_549,In_560,In_451);
xor U550 (N_550,In_429,In_349);
nand U551 (N_551,In_240,In_472);
nand U552 (N_552,In_629,In_583);
nand U553 (N_553,In_539,In_135);
and U554 (N_554,In_196,In_425);
xnor U555 (N_555,In_348,In_405);
nand U556 (N_556,In_304,In_612);
or U557 (N_557,In_91,In_241);
or U558 (N_558,In_35,In_155);
and U559 (N_559,In_323,In_426);
and U560 (N_560,In_540,In_291);
and U561 (N_561,In_443,In_4);
nand U562 (N_562,In_635,In_278);
nor U563 (N_563,In_92,In_536);
or U564 (N_564,In_68,In_640);
nor U565 (N_565,In_52,In_503);
and U566 (N_566,In_344,In_231);
and U567 (N_567,In_352,In_732);
and U568 (N_568,In_226,In_709);
and U569 (N_569,In_616,In_607);
nor U570 (N_570,In_452,In_247);
or U571 (N_571,In_710,In_313);
or U572 (N_572,In_29,In_38);
and U573 (N_573,In_662,In_5);
nand U574 (N_574,In_598,In_101);
xnor U575 (N_575,In_623,In_711);
nor U576 (N_576,In_238,In_467);
or U577 (N_577,In_421,In_238);
or U578 (N_578,In_32,In_667);
or U579 (N_579,In_136,In_275);
nor U580 (N_580,In_570,In_615);
or U581 (N_581,In_485,In_565);
or U582 (N_582,In_396,In_523);
nor U583 (N_583,In_421,In_149);
or U584 (N_584,In_415,In_56);
nand U585 (N_585,In_685,In_405);
xor U586 (N_586,In_556,In_721);
nand U587 (N_587,In_172,In_159);
xnor U588 (N_588,In_593,In_621);
xor U589 (N_589,In_360,In_497);
nor U590 (N_590,In_629,In_588);
nor U591 (N_591,In_304,In_394);
and U592 (N_592,In_36,In_299);
or U593 (N_593,In_400,In_741);
or U594 (N_594,In_628,In_106);
xnor U595 (N_595,In_98,In_207);
and U596 (N_596,In_294,In_683);
or U597 (N_597,In_642,In_484);
nand U598 (N_598,In_540,In_675);
nor U599 (N_599,In_158,In_679);
and U600 (N_600,In_324,In_99);
nand U601 (N_601,In_608,In_460);
xor U602 (N_602,In_39,In_576);
nand U603 (N_603,In_670,In_522);
or U604 (N_604,In_721,In_248);
or U605 (N_605,In_458,In_250);
nor U606 (N_606,In_243,In_177);
nand U607 (N_607,In_745,In_728);
nand U608 (N_608,In_556,In_436);
and U609 (N_609,In_423,In_562);
or U610 (N_610,In_634,In_277);
nor U611 (N_611,In_480,In_430);
nand U612 (N_612,In_494,In_0);
or U613 (N_613,In_532,In_299);
or U614 (N_614,In_120,In_332);
nand U615 (N_615,In_530,In_10);
and U616 (N_616,In_269,In_649);
or U617 (N_617,In_68,In_342);
and U618 (N_618,In_238,In_715);
and U619 (N_619,In_446,In_552);
and U620 (N_620,In_653,In_395);
nor U621 (N_621,In_587,In_631);
xor U622 (N_622,In_431,In_366);
nor U623 (N_623,In_385,In_351);
nand U624 (N_624,In_638,In_382);
or U625 (N_625,In_516,In_267);
nand U626 (N_626,In_224,In_551);
nand U627 (N_627,In_462,In_266);
nand U628 (N_628,In_641,In_595);
nand U629 (N_629,In_540,In_721);
nor U630 (N_630,In_444,In_175);
nand U631 (N_631,In_359,In_221);
and U632 (N_632,In_74,In_120);
nand U633 (N_633,In_371,In_124);
nor U634 (N_634,In_135,In_648);
nand U635 (N_635,In_221,In_103);
nand U636 (N_636,In_607,In_20);
nand U637 (N_637,In_414,In_110);
nor U638 (N_638,In_251,In_403);
and U639 (N_639,In_701,In_454);
or U640 (N_640,In_134,In_478);
and U641 (N_641,In_84,In_162);
and U642 (N_642,In_439,In_344);
xnor U643 (N_643,In_576,In_394);
xnor U644 (N_644,In_322,In_184);
nor U645 (N_645,In_51,In_649);
nor U646 (N_646,In_46,In_449);
nand U647 (N_647,In_745,In_571);
nand U648 (N_648,In_743,In_115);
nor U649 (N_649,In_179,In_501);
nor U650 (N_650,In_311,In_85);
nor U651 (N_651,In_431,In_479);
or U652 (N_652,In_128,In_31);
and U653 (N_653,In_630,In_383);
xor U654 (N_654,In_457,In_741);
nand U655 (N_655,In_356,In_283);
nand U656 (N_656,In_739,In_237);
nand U657 (N_657,In_368,In_372);
nor U658 (N_658,In_419,In_451);
xnor U659 (N_659,In_196,In_515);
or U660 (N_660,In_472,In_257);
nor U661 (N_661,In_354,In_52);
xor U662 (N_662,In_0,In_309);
nor U663 (N_663,In_310,In_69);
nor U664 (N_664,In_333,In_359);
nor U665 (N_665,In_320,In_345);
and U666 (N_666,In_519,In_237);
xnor U667 (N_667,In_506,In_511);
nor U668 (N_668,In_348,In_569);
xor U669 (N_669,In_157,In_25);
nand U670 (N_670,In_638,In_61);
and U671 (N_671,In_192,In_345);
or U672 (N_672,In_367,In_187);
and U673 (N_673,In_212,In_468);
or U674 (N_674,In_172,In_107);
xnor U675 (N_675,In_409,In_169);
nand U676 (N_676,In_221,In_316);
nor U677 (N_677,In_705,In_188);
and U678 (N_678,In_600,In_732);
or U679 (N_679,In_624,In_231);
or U680 (N_680,In_401,In_620);
or U681 (N_681,In_45,In_106);
xor U682 (N_682,In_75,In_205);
and U683 (N_683,In_49,In_412);
nor U684 (N_684,In_372,In_29);
nand U685 (N_685,In_376,In_243);
xnor U686 (N_686,In_246,In_46);
and U687 (N_687,In_509,In_402);
or U688 (N_688,In_323,In_463);
nor U689 (N_689,In_213,In_544);
or U690 (N_690,In_331,In_747);
or U691 (N_691,In_415,In_462);
and U692 (N_692,In_482,In_303);
nand U693 (N_693,In_514,In_97);
or U694 (N_694,In_522,In_412);
and U695 (N_695,In_562,In_165);
nand U696 (N_696,In_571,In_565);
and U697 (N_697,In_705,In_522);
or U698 (N_698,In_203,In_577);
or U699 (N_699,In_614,In_530);
or U700 (N_700,In_560,In_688);
xor U701 (N_701,In_147,In_459);
and U702 (N_702,In_497,In_36);
nor U703 (N_703,In_85,In_276);
or U704 (N_704,In_230,In_494);
nor U705 (N_705,In_126,In_288);
xor U706 (N_706,In_76,In_524);
or U707 (N_707,In_445,In_505);
and U708 (N_708,In_155,In_551);
or U709 (N_709,In_143,In_359);
nor U710 (N_710,In_56,In_149);
nand U711 (N_711,In_114,In_258);
or U712 (N_712,In_748,In_18);
nor U713 (N_713,In_585,In_455);
or U714 (N_714,In_102,In_741);
nor U715 (N_715,In_205,In_628);
and U716 (N_716,In_519,In_226);
xor U717 (N_717,In_510,In_496);
nand U718 (N_718,In_662,In_495);
nand U719 (N_719,In_7,In_393);
xor U720 (N_720,In_421,In_55);
nor U721 (N_721,In_538,In_408);
or U722 (N_722,In_224,In_418);
xnor U723 (N_723,In_162,In_308);
nand U724 (N_724,In_647,In_506);
nor U725 (N_725,In_226,In_258);
or U726 (N_726,In_64,In_523);
nand U727 (N_727,In_386,In_687);
nand U728 (N_728,In_150,In_686);
and U729 (N_729,In_33,In_286);
xnor U730 (N_730,In_673,In_677);
and U731 (N_731,In_6,In_350);
nand U732 (N_732,In_269,In_544);
or U733 (N_733,In_642,In_313);
nand U734 (N_734,In_284,In_527);
or U735 (N_735,In_452,In_685);
xor U736 (N_736,In_734,In_220);
and U737 (N_737,In_73,In_542);
or U738 (N_738,In_496,In_251);
nand U739 (N_739,In_75,In_333);
xnor U740 (N_740,In_106,In_735);
nand U741 (N_741,In_392,In_455);
nor U742 (N_742,In_292,In_350);
or U743 (N_743,In_510,In_98);
nand U744 (N_744,In_61,In_716);
nand U745 (N_745,In_648,In_287);
nor U746 (N_746,In_593,In_516);
and U747 (N_747,In_634,In_581);
nand U748 (N_748,In_215,In_563);
nor U749 (N_749,In_276,In_324);
nand U750 (N_750,In_125,In_36);
nand U751 (N_751,In_150,In_507);
or U752 (N_752,In_249,In_248);
nor U753 (N_753,In_548,In_501);
or U754 (N_754,In_634,In_533);
nor U755 (N_755,In_686,In_117);
or U756 (N_756,In_665,In_541);
nand U757 (N_757,In_121,In_258);
or U758 (N_758,In_196,In_554);
and U759 (N_759,In_303,In_339);
nor U760 (N_760,In_512,In_433);
nor U761 (N_761,In_138,In_646);
nor U762 (N_762,In_647,In_353);
or U763 (N_763,In_220,In_632);
nand U764 (N_764,In_600,In_339);
and U765 (N_765,In_159,In_629);
and U766 (N_766,In_589,In_459);
nand U767 (N_767,In_56,In_25);
or U768 (N_768,In_48,In_190);
or U769 (N_769,In_583,In_247);
xor U770 (N_770,In_554,In_484);
nor U771 (N_771,In_90,In_681);
nor U772 (N_772,In_421,In_21);
and U773 (N_773,In_469,In_482);
xor U774 (N_774,In_56,In_452);
or U775 (N_775,In_30,In_582);
and U776 (N_776,In_316,In_30);
nor U777 (N_777,In_384,In_2);
nor U778 (N_778,In_81,In_290);
xnor U779 (N_779,In_89,In_461);
nor U780 (N_780,In_648,In_458);
and U781 (N_781,In_330,In_319);
or U782 (N_782,In_482,In_219);
nor U783 (N_783,In_200,In_104);
and U784 (N_784,In_20,In_468);
nor U785 (N_785,In_143,In_746);
or U786 (N_786,In_618,In_390);
nand U787 (N_787,In_295,In_39);
and U788 (N_788,In_335,In_262);
and U789 (N_789,In_142,In_258);
nand U790 (N_790,In_361,In_376);
nand U791 (N_791,In_549,In_158);
and U792 (N_792,In_613,In_425);
and U793 (N_793,In_679,In_526);
and U794 (N_794,In_279,In_631);
and U795 (N_795,In_18,In_194);
nand U796 (N_796,In_376,In_221);
nor U797 (N_797,In_327,In_73);
nand U798 (N_798,In_234,In_98);
nor U799 (N_799,In_260,In_453);
and U800 (N_800,In_359,In_11);
and U801 (N_801,In_314,In_668);
nor U802 (N_802,In_79,In_427);
or U803 (N_803,In_464,In_558);
nor U804 (N_804,In_673,In_581);
nand U805 (N_805,In_32,In_282);
nor U806 (N_806,In_570,In_7);
and U807 (N_807,In_699,In_276);
or U808 (N_808,In_745,In_689);
or U809 (N_809,In_651,In_636);
nand U810 (N_810,In_602,In_645);
xnor U811 (N_811,In_138,In_401);
nand U812 (N_812,In_500,In_589);
nand U813 (N_813,In_156,In_573);
nor U814 (N_814,In_29,In_140);
xnor U815 (N_815,In_404,In_420);
or U816 (N_816,In_624,In_77);
xnor U817 (N_817,In_678,In_377);
and U818 (N_818,In_441,In_706);
and U819 (N_819,In_79,In_295);
nor U820 (N_820,In_290,In_469);
and U821 (N_821,In_579,In_427);
nor U822 (N_822,In_42,In_127);
xor U823 (N_823,In_736,In_686);
and U824 (N_824,In_35,In_665);
and U825 (N_825,In_59,In_209);
nand U826 (N_826,In_102,In_721);
and U827 (N_827,In_94,In_387);
nor U828 (N_828,In_554,In_2);
and U829 (N_829,In_44,In_430);
and U830 (N_830,In_672,In_574);
and U831 (N_831,In_467,In_198);
nand U832 (N_832,In_576,In_685);
or U833 (N_833,In_217,In_105);
or U834 (N_834,In_601,In_482);
and U835 (N_835,In_113,In_395);
and U836 (N_836,In_234,In_501);
xnor U837 (N_837,In_44,In_448);
and U838 (N_838,In_403,In_279);
and U839 (N_839,In_371,In_137);
and U840 (N_840,In_523,In_733);
and U841 (N_841,In_712,In_192);
nand U842 (N_842,In_635,In_221);
and U843 (N_843,In_368,In_21);
nor U844 (N_844,In_172,In_84);
or U845 (N_845,In_116,In_103);
nor U846 (N_846,In_734,In_277);
and U847 (N_847,In_52,In_258);
nor U848 (N_848,In_456,In_449);
nand U849 (N_849,In_545,In_258);
xor U850 (N_850,In_549,In_411);
nand U851 (N_851,In_650,In_152);
or U852 (N_852,In_465,In_691);
and U853 (N_853,In_67,In_248);
nor U854 (N_854,In_629,In_267);
and U855 (N_855,In_722,In_242);
nand U856 (N_856,In_111,In_267);
and U857 (N_857,In_335,In_564);
and U858 (N_858,In_318,In_453);
and U859 (N_859,In_641,In_56);
nor U860 (N_860,In_708,In_546);
or U861 (N_861,In_625,In_208);
xnor U862 (N_862,In_246,In_143);
or U863 (N_863,In_452,In_164);
and U864 (N_864,In_124,In_144);
nor U865 (N_865,In_707,In_19);
nor U866 (N_866,In_602,In_556);
xnor U867 (N_867,In_4,In_148);
nand U868 (N_868,In_553,In_209);
nor U869 (N_869,In_461,In_716);
nand U870 (N_870,In_713,In_34);
nor U871 (N_871,In_142,In_559);
nor U872 (N_872,In_141,In_730);
nand U873 (N_873,In_466,In_305);
nor U874 (N_874,In_297,In_247);
nor U875 (N_875,In_129,In_185);
nor U876 (N_876,In_1,In_464);
nor U877 (N_877,In_723,In_33);
and U878 (N_878,In_120,In_637);
nand U879 (N_879,In_188,In_449);
xnor U880 (N_880,In_402,In_709);
nor U881 (N_881,In_269,In_11);
nor U882 (N_882,In_180,In_359);
xnor U883 (N_883,In_635,In_617);
xor U884 (N_884,In_725,In_544);
and U885 (N_885,In_514,In_130);
nor U886 (N_886,In_314,In_91);
nand U887 (N_887,In_233,In_72);
or U888 (N_888,In_224,In_637);
and U889 (N_889,In_603,In_370);
or U890 (N_890,In_275,In_510);
nor U891 (N_891,In_676,In_429);
nand U892 (N_892,In_39,In_662);
xnor U893 (N_893,In_717,In_401);
and U894 (N_894,In_347,In_640);
nor U895 (N_895,In_608,In_600);
nor U896 (N_896,In_558,In_692);
xnor U897 (N_897,In_102,In_609);
nor U898 (N_898,In_660,In_469);
nand U899 (N_899,In_654,In_52);
and U900 (N_900,In_326,In_170);
and U901 (N_901,In_256,In_565);
nand U902 (N_902,In_492,In_630);
nor U903 (N_903,In_80,In_41);
or U904 (N_904,In_741,In_260);
and U905 (N_905,In_698,In_714);
nor U906 (N_906,In_694,In_673);
or U907 (N_907,In_592,In_610);
nor U908 (N_908,In_438,In_361);
or U909 (N_909,In_81,In_655);
and U910 (N_910,In_35,In_535);
xnor U911 (N_911,In_408,In_476);
and U912 (N_912,In_306,In_54);
and U913 (N_913,In_701,In_694);
nor U914 (N_914,In_440,In_46);
nor U915 (N_915,In_573,In_185);
nand U916 (N_916,In_632,In_43);
or U917 (N_917,In_249,In_364);
and U918 (N_918,In_415,In_427);
and U919 (N_919,In_725,In_310);
and U920 (N_920,In_711,In_229);
nor U921 (N_921,In_105,In_472);
or U922 (N_922,In_611,In_439);
or U923 (N_923,In_471,In_586);
xnor U924 (N_924,In_285,In_53);
or U925 (N_925,In_510,In_580);
nand U926 (N_926,In_278,In_191);
or U927 (N_927,In_53,In_586);
nor U928 (N_928,In_80,In_629);
nand U929 (N_929,In_72,In_666);
or U930 (N_930,In_485,In_273);
nand U931 (N_931,In_427,In_154);
nand U932 (N_932,In_541,In_240);
nor U933 (N_933,In_131,In_430);
nand U934 (N_934,In_482,In_453);
nand U935 (N_935,In_261,In_669);
or U936 (N_936,In_659,In_241);
nor U937 (N_937,In_411,In_509);
and U938 (N_938,In_693,In_745);
nand U939 (N_939,In_442,In_661);
nor U940 (N_940,In_128,In_613);
nor U941 (N_941,In_477,In_453);
or U942 (N_942,In_199,In_446);
nor U943 (N_943,In_695,In_568);
nor U944 (N_944,In_58,In_241);
xor U945 (N_945,In_671,In_200);
nand U946 (N_946,In_618,In_446);
or U947 (N_947,In_370,In_704);
nand U948 (N_948,In_634,In_319);
and U949 (N_949,In_533,In_585);
and U950 (N_950,In_206,In_240);
xnor U951 (N_951,In_608,In_633);
and U952 (N_952,In_277,In_316);
nand U953 (N_953,In_95,In_507);
nor U954 (N_954,In_398,In_377);
or U955 (N_955,In_392,In_584);
xor U956 (N_956,In_132,In_585);
and U957 (N_957,In_641,In_472);
or U958 (N_958,In_253,In_621);
nor U959 (N_959,In_178,In_35);
and U960 (N_960,In_75,In_580);
nand U961 (N_961,In_590,In_265);
and U962 (N_962,In_195,In_311);
nand U963 (N_963,In_275,In_121);
nor U964 (N_964,In_408,In_20);
xnor U965 (N_965,In_143,In_139);
nor U966 (N_966,In_226,In_291);
nand U967 (N_967,In_54,In_69);
nand U968 (N_968,In_207,In_241);
and U969 (N_969,In_600,In_352);
nor U970 (N_970,In_96,In_609);
nor U971 (N_971,In_21,In_13);
and U972 (N_972,In_323,In_584);
nor U973 (N_973,In_226,In_593);
or U974 (N_974,In_228,In_154);
or U975 (N_975,In_326,In_469);
nor U976 (N_976,In_284,In_445);
xor U977 (N_977,In_573,In_172);
xnor U978 (N_978,In_388,In_145);
nand U979 (N_979,In_483,In_265);
and U980 (N_980,In_453,In_153);
or U981 (N_981,In_635,In_252);
and U982 (N_982,In_392,In_728);
nor U983 (N_983,In_631,In_288);
nor U984 (N_984,In_527,In_390);
xnor U985 (N_985,In_453,In_225);
or U986 (N_986,In_215,In_552);
or U987 (N_987,In_556,In_363);
nand U988 (N_988,In_672,In_164);
xor U989 (N_989,In_141,In_402);
and U990 (N_990,In_221,In_690);
and U991 (N_991,In_489,In_111);
or U992 (N_992,In_122,In_279);
nand U993 (N_993,In_227,In_202);
or U994 (N_994,In_743,In_77);
nor U995 (N_995,In_481,In_494);
nor U996 (N_996,In_599,In_102);
and U997 (N_997,In_661,In_297);
nor U998 (N_998,In_646,In_636);
nor U999 (N_999,In_481,In_117);
nor U1000 (N_1000,In_572,In_35);
nor U1001 (N_1001,In_395,In_463);
or U1002 (N_1002,In_632,In_191);
nor U1003 (N_1003,In_423,In_235);
nand U1004 (N_1004,In_489,In_694);
or U1005 (N_1005,In_110,In_534);
nor U1006 (N_1006,In_212,In_298);
xor U1007 (N_1007,In_389,In_284);
and U1008 (N_1008,In_404,In_154);
nand U1009 (N_1009,In_424,In_319);
or U1010 (N_1010,In_279,In_672);
nand U1011 (N_1011,In_522,In_85);
and U1012 (N_1012,In_75,In_408);
or U1013 (N_1013,In_442,In_344);
nor U1014 (N_1014,In_475,In_6);
nor U1015 (N_1015,In_737,In_266);
nor U1016 (N_1016,In_421,In_334);
nand U1017 (N_1017,In_179,In_7);
nand U1018 (N_1018,In_531,In_68);
nand U1019 (N_1019,In_30,In_54);
nand U1020 (N_1020,In_619,In_31);
and U1021 (N_1021,In_613,In_210);
or U1022 (N_1022,In_255,In_172);
nor U1023 (N_1023,In_22,In_505);
or U1024 (N_1024,In_397,In_273);
nand U1025 (N_1025,In_690,In_611);
xor U1026 (N_1026,In_388,In_129);
nor U1027 (N_1027,In_375,In_71);
and U1028 (N_1028,In_682,In_316);
nand U1029 (N_1029,In_62,In_215);
nand U1030 (N_1030,In_437,In_722);
nand U1031 (N_1031,In_546,In_637);
nor U1032 (N_1032,In_207,In_49);
nand U1033 (N_1033,In_519,In_471);
or U1034 (N_1034,In_641,In_447);
or U1035 (N_1035,In_98,In_624);
and U1036 (N_1036,In_461,In_606);
nand U1037 (N_1037,In_250,In_587);
and U1038 (N_1038,In_99,In_106);
or U1039 (N_1039,In_406,In_199);
nor U1040 (N_1040,In_78,In_655);
and U1041 (N_1041,In_563,In_488);
nor U1042 (N_1042,In_380,In_287);
nor U1043 (N_1043,In_443,In_397);
nor U1044 (N_1044,In_479,In_707);
nor U1045 (N_1045,In_477,In_562);
nor U1046 (N_1046,In_586,In_83);
and U1047 (N_1047,In_245,In_64);
nand U1048 (N_1048,In_623,In_486);
or U1049 (N_1049,In_631,In_450);
nor U1050 (N_1050,In_447,In_528);
nor U1051 (N_1051,In_296,In_246);
or U1052 (N_1052,In_502,In_652);
or U1053 (N_1053,In_201,In_379);
xnor U1054 (N_1054,In_198,In_207);
and U1055 (N_1055,In_285,In_421);
nand U1056 (N_1056,In_406,In_218);
or U1057 (N_1057,In_210,In_484);
and U1058 (N_1058,In_137,In_449);
nand U1059 (N_1059,In_30,In_87);
and U1060 (N_1060,In_210,In_253);
nor U1061 (N_1061,In_280,In_407);
nand U1062 (N_1062,In_289,In_530);
nor U1063 (N_1063,In_249,In_261);
xor U1064 (N_1064,In_494,In_250);
or U1065 (N_1065,In_496,In_680);
xor U1066 (N_1066,In_704,In_151);
nand U1067 (N_1067,In_557,In_382);
or U1068 (N_1068,In_186,In_208);
or U1069 (N_1069,In_556,In_27);
nand U1070 (N_1070,In_708,In_215);
and U1071 (N_1071,In_653,In_602);
and U1072 (N_1072,In_445,In_636);
or U1073 (N_1073,In_732,In_105);
nand U1074 (N_1074,In_707,In_11);
or U1075 (N_1075,In_607,In_234);
or U1076 (N_1076,In_415,In_245);
and U1077 (N_1077,In_270,In_644);
xnor U1078 (N_1078,In_576,In_535);
nand U1079 (N_1079,In_89,In_494);
xor U1080 (N_1080,In_720,In_537);
and U1081 (N_1081,In_45,In_584);
nor U1082 (N_1082,In_324,In_141);
and U1083 (N_1083,In_605,In_7);
or U1084 (N_1084,In_137,In_501);
nor U1085 (N_1085,In_687,In_367);
nor U1086 (N_1086,In_571,In_248);
or U1087 (N_1087,In_701,In_627);
or U1088 (N_1088,In_222,In_113);
or U1089 (N_1089,In_241,In_9);
and U1090 (N_1090,In_622,In_497);
and U1091 (N_1091,In_103,In_205);
nand U1092 (N_1092,In_692,In_554);
and U1093 (N_1093,In_746,In_570);
nor U1094 (N_1094,In_680,In_133);
and U1095 (N_1095,In_624,In_357);
and U1096 (N_1096,In_345,In_473);
nand U1097 (N_1097,In_436,In_152);
and U1098 (N_1098,In_233,In_327);
nor U1099 (N_1099,In_671,In_582);
or U1100 (N_1100,In_338,In_742);
or U1101 (N_1101,In_126,In_376);
nor U1102 (N_1102,In_574,In_455);
nor U1103 (N_1103,In_573,In_70);
nand U1104 (N_1104,In_170,In_3);
and U1105 (N_1105,In_322,In_237);
xnor U1106 (N_1106,In_49,In_448);
xnor U1107 (N_1107,In_529,In_217);
or U1108 (N_1108,In_158,In_227);
or U1109 (N_1109,In_604,In_507);
and U1110 (N_1110,In_310,In_358);
and U1111 (N_1111,In_643,In_207);
xor U1112 (N_1112,In_342,In_139);
and U1113 (N_1113,In_178,In_507);
nand U1114 (N_1114,In_1,In_12);
nand U1115 (N_1115,In_42,In_317);
nor U1116 (N_1116,In_31,In_741);
nor U1117 (N_1117,In_525,In_36);
xor U1118 (N_1118,In_248,In_438);
nor U1119 (N_1119,In_403,In_387);
nor U1120 (N_1120,In_417,In_486);
or U1121 (N_1121,In_307,In_491);
and U1122 (N_1122,In_659,In_725);
or U1123 (N_1123,In_129,In_610);
and U1124 (N_1124,In_470,In_552);
or U1125 (N_1125,In_519,In_403);
nand U1126 (N_1126,In_476,In_538);
nand U1127 (N_1127,In_400,In_695);
or U1128 (N_1128,In_719,In_144);
nor U1129 (N_1129,In_727,In_110);
nor U1130 (N_1130,In_240,In_648);
or U1131 (N_1131,In_238,In_675);
xnor U1132 (N_1132,In_49,In_516);
nor U1133 (N_1133,In_613,In_655);
or U1134 (N_1134,In_413,In_384);
nor U1135 (N_1135,In_340,In_616);
and U1136 (N_1136,In_244,In_552);
or U1137 (N_1137,In_664,In_670);
nand U1138 (N_1138,In_124,In_27);
nand U1139 (N_1139,In_328,In_245);
nand U1140 (N_1140,In_742,In_503);
nor U1141 (N_1141,In_176,In_660);
and U1142 (N_1142,In_688,In_334);
xor U1143 (N_1143,In_205,In_285);
or U1144 (N_1144,In_104,In_725);
nor U1145 (N_1145,In_177,In_193);
nor U1146 (N_1146,In_613,In_147);
nand U1147 (N_1147,In_564,In_321);
nand U1148 (N_1148,In_577,In_165);
or U1149 (N_1149,In_441,In_687);
nor U1150 (N_1150,In_162,In_189);
or U1151 (N_1151,In_333,In_37);
or U1152 (N_1152,In_127,In_553);
nand U1153 (N_1153,In_659,In_583);
and U1154 (N_1154,In_35,In_267);
nor U1155 (N_1155,In_641,In_91);
nor U1156 (N_1156,In_663,In_554);
nor U1157 (N_1157,In_182,In_384);
and U1158 (N_1158,In_378,In_108);
nand U1159 (N_1159,In_221,In_94);
nand U1160 (N_1160,In_212,In_306);
or U1161 (N_1161,In_91,In_119);
nand U1162 (N_1162,In_646,In_238);
nand U1163 (N_1163,In_71,In_406);
or U1164 (N_1164,In_165,In_670);
or U1165 (N_1165,In_495,In_105);
and U1166 (N_1166,In_461,In_197);
or U1167 (N_1167,In_682,In_184);
nand U1168 (N_1168,In_536,In_139);
or U1169 (N_1169,In_189,In_577);
nor U1170 (N_1170,In_194,In_27);
nand U1171 (N_1171,In_426,In_94);
nand U1172 (N_1172,In_565,In_622);
nand U1173 (N_1173,In_245,In_645);
nand U1174 (N_1174,In_397,In_57);
and U1175 (N_1175,In_44,In_327);
or U1176 (N_1176,In_460,In_535);
xor U1177 (N_1177,In_746,In_711);
and U1178 (N_1178,In_149,In_91);
nor U1179 (N_1179,In_418,In_63);
or U1180 (N_1180,In_144,In_249);
nor U1181 (N_1181,In_179,In_252);
and U1182 (N_1182,In_141,In_534);
nand U1183 (N_1183,In_151,In_195);
nand U1184 (N_1184,In_741,In_198);
or U1185 (N_1185,In_541,In_493);
nor U1186 (N_1186,In_479,In_538);
or U1187 (N_1187,In_423,In_144);
or U1188 (N_1188,In_398,In_600);
xnor U1189 (N_1189,In_707,In_312);
and U1190 (N_1190,In_439,In_115);
nor U1191 (N_1191,In_275,In_138);
and U1192 (N_1192,In_266,In_206);
nand U1193 (N_1193,In_325,In_88);
nor U1194 (N_1194,In_387,In_330);
nor U1195 (N_1195,In_448,In_501);
nand U1196 (N_1196,In_174,In_29);
xnor U1197 (N_1197,In_195,In_526);
and U1198 (N_1198,In_465,In_227);
nor U1199 (N_1199,In_111,In_215);
xor U1200 (N_1200,In_597,In_125);
or U1201 (N_1201,In_715,In_394);
xnor U1202 (N_1202,In_282,In_513);
or U1203 (N_1203,In_577,In_710);
nor U1204 (N_1204,In_338,In_703);
and U1205 (N_1205,In_376,In_382);
nor U1206 (N_1206,In_435,In_537);
and U1207 (N_1207,In_329,In_253);
nor U1208 (N_1208,In_2,In_361);
or U1209 (N_1209,In_300,In_694);
and U1210 (N_1210,In_84,In_52);
nor U1211 (N_1211,In_129,In_257);
or U1212 (N_1212,In_114,In_736);
or U1213 (N_1213,In_139,In_554);
and U1214 (N_1214,In_125,In_674);
and U1215 (N_1215,In_344,In_280);
nand U1216 (N_1216,In_60,In_36);
xor U1217 (N_1217,In_237,In_540);
and U1218 (N_1218,In_68,In_496);
nor U1219 (N_1219,In_55,In_98);
or U1220 (N_1220,In_188,In_345);
or U1221 (N_1221,In_440,In_132);
nor U1222 (N_1222,In_364,In_297);
or U1223 (N_1223,In_587,In_640);
or U1224 (N_1224,In_163,In_184);
and U1225 (N_1225,In_283,In_290);
and U1226 (N_1226,In_137,In_648);
nor U1227 (N_1227,In_70,In_333);
nand U1228 (N_1228,In_300,In_25);
or U1229 (N_1229,In_714,In_372);
nand U1230 (N_1230,In_488,In_287);
or U1231 (N_1231,In_143,In_30);
and U1232 (N_1232,In_78,In_353);
nor U1233 (N_1233,In_595,In_428);
nor U1234 (N_1234,In_480,In_466);
and U1235 (N_1235,In_428,In_381);
and U1236 (N_1236,In_103,In_391);
nor U1237 (N_1237,In_349,In_710);
nand U1238 (N_1238,In_573,In_31);
and U1239 (N_1239,In_427,In_116);
nor U1240 (N_1240,In_357,In_428);
nor U1241 (N_1241,In_571,In_563);
nor U1242 (N_1242,In_433,In_700);
nor U1243 (N_1243,In_520,In_18);
and U1244 (N_1244,In_304,In_366);
and U1245 (N_1245,In_546,In_66);
or U1246 (N_1246,In_327,In_108);
or U1247 (N_1247,In_270,In_157);
or U1248 (N_1248,In_171,In_422);
nand U1249 (N_1249,In_428,In_257);
nor U1250 (N_1250,In_592,In_290);
and U1251 (N_1251,In_299,In_108);
and U1252 (N_1252,In_55,In_389);
nor U1253 (N_1253,In_528,In_284);
or U1254 (N_1254,In_491,In_642);
nand U1255 (N_1255,In_529,In_607);
and U1256 (N_1256,In_137,In_70);
nand U1257 (N_1257,In_44,In_239);
and U1258 (N_1258,In_195,In_82);
or U1259 (N_1259,In_720,In_565);
nand U1260 (N_1260,In_258,In_269);
nand U1261 (N_1261,In_176,In_156);
nand U1262 (N_1262,In_602,In_154);
nor U1263 (N_1263,In_249,In_72);
nor U1264 (N_1264,In_593,In_421);
nor U1265 (N_1265,In_306,In_353);
nor U1266 (N_1266,In_576,In_293);
nand U1267 (N_1267,In_94,In_102);
or U1268 (N_1268,In_611,In_331);
and U1269 (N_1269,In_277,In_612);
nand U1270 (N_1270,In_663,In_635);
xnor U1271 (N_1271,In_601,In_321);
nand U1272 (N_1272,In_40,In_623);
nor U1273 (N_1273,In_665,In_568);
and U1274 (N_1274,In_297,In_68);
or U1275 (N_1275,In_531,In_432);
or U1276 (N_1276,In_677,In_117);
nand U1277 (N_1277,In_460,In_334);
or U1278 (N_1278,In_680,In_612);
or U1279 (N_1279,In_556,In_483);
xnor U1280 (N_1280,In_702,In_103);
and U1281 (N_1281,In_544,In_530);
nand U1282 (N_1282,In_482,In_411);
nand U1283 (N_1283,In_590,In_408);
nor U1284 (N_1284,In_203,In_327);
or U1285 (N_1285,In_52,In_213);
xor U1286 (N_1286,In_437,In_625);
and U1287 (N_1287,In_79,In_652);
nor U1288 (N_1288,In_201,In_309);
nor U1289 (N_1289,In_534,In_54);
nor U1290 (N_1290,In_204,In_537);
nand U1291 (N_1291,In_447,In_617);
and U1292 (N_1292,In_239,In_342);
nand U1293 (N_1293,In_364,In_41);
or U1294 (N_1294,In_639,In_627);
nand U1295 (N_1295,In_256,In_449);
and U1296 (N_1296,In_175,In_681);
xnor U1297 (N_1297,In_137,In_583);
or U1298 (N_1298,In_296,In_712);
nor U1299 (N_1299,In_697,In_665);
or U1300 (N_1300,In_592,In_715);
nor U1301 (N_1301,In_669,In_518);
nor U1302 (N_1302,In_167,In_72);
nor U1303 (N_1303,In_315,In_503);
or U1304 (N_1304,In_353,In_47);
xor U1305 (N_1305,In_204,In_264);
nor U1306 (N_1306,In_77,In_15);
or U1307 (N_1307,In_743,In_55);
xor U1308 (N_1308,In_570,In_613);
and U1309 (N_1309,In_128,In_499);
and U1310 (N_1310,In_494,In_81);
nor U1311 (N_1311,In_267,In_725);
and U1312 (N_1312,In_682,In_581);
nor U1313 (N_1313,In_600,In_361);
xor U1314 (N_1314,In_684,In_416);
nand U1315 (N_1315,In_578,In_342);
nand U1316 (N_1316,In_23,In_385);
or U1317 (N_1317,In_363,In_42);
nand U1318 (N_1318,In_729,In_575);
and U1319 (N_1319,In_410,In_532);
nand U1320 (N_1320,In_58,In_597);
and U1321 (N_1321,In_116,In_166);
or U1322 (N_1322,In_228,In_43);
nor U1323 (N_1323,In_470,In_654);
nor U1324 (N_1324,In_630,In_260);
nand U1325 (N_1325,In_64,In_2);
nand U1326 (N_1326,In_126,In_430);
nor U1327 (N_1327,In_497,In_495);
nor U1328 (N_1328,In_217,In_267);
nor U1329 (N_1329,In_370,In_281);
or U1330 (N_1330,In_202,In_38);
nor U1331 (N_1331,In_686,In_200);
or U1332 (N_1332,In_189,In_706);
nor U1333 (N_1333,In_414,In_308);
xor U1334 (N_1334,In_32,In_157);
or U1335 (N_1335,In_622,In_44);
nand U1336 (N_1336,In_14,In_352);
and U1337 (N_1337,In_719,In_350);
or U1338 (N_1338,In_111,In_440);
nand U1339 (N_1339,In_508,In_584);
nand U1340 (N_1340,In_90,In_601);
nor U1341 (N_1341,In_377,In_615);
xnor U1342 (N_1342,In_264,In_199);
nand U1343 (N_1343,In_612,In_674);
nor U1344 (N_1344,In_125,In_570);
or U1345 (N_1345,In_150,In_742);
nor U1346 (N_1346,In_327,In_670);
nor U1347 (N_1347,In_724,In_658);
and U1348 (N_1348,In_712,In_240);
and U1349 (N_1349,In_237,In_388);
and U1350 (N_1350,In_88,In_554);
nand U1351 (N_1351,In_336,In_57);
nor U1352 (N_1352,In_170,In_688);
or U1353 (N_1353,In_373,In_462);
and U1354 (N_1354,In_400,In_652);
or U1355 (N_1355,In_8,In_223);
and U1356 (N_1356,In_718,In_379);
or U1357 (N_1357,In_339,In_201);
and U1358 (N_1358,In_526,In_6);
nor U1359 (N_1359,In_118,In_462);
nor U1360 (N_1360,In_674,In_704);
xor U1361 (N_1361,In_560,In_86);
xor U1362 (N_1362,In_590,In_626);
or U1363 (N_1363,In_276,In_743);
nand U1364 (N_1364,In_24,In_722);
nand U1365 (N_1365,In_479,In_21);
nor U1366 (N_1366,In_692,In_663);
nor U1367 (N_1367,In_450,In_730);
nor U1368 (N_1368,In_601,In_610);
nor U1369 (N_1369,In_409,In_229);
nor U1370 (N_1370,In_603,In_638);
xor U1371 (N_1371,In_50,In_508);
nand U1372 (N_1372,In_548,In_506);
and U1373 (N_1373,In_546,In_241);
nor U1374 (N_1374,In_77,In_555);
nor U1375 (N_1375,In_408,In_66);
nor U1376 (N_1376,In_650,In_636);
nand U1377 (N_1377,In_121,In_459);
or U1378 (N_1378,In_479,In_204);
and U1379 (N_1379,In_426,In_636);
or U1380 (N_1380,In_693,In_729);
nor U1381 (N_1381,In_614,In_197);
nand U1382 (N_1382,In_270,In_260);
nor U1383 (N_1383,In_397,In_50);
or U1384 (N_1384,In_512,In_504);
or U1385 (N_1385,In_558,In_184);
nor U1386 (N_1386,In_225,In_637);
xor U1387 (N_1387,In_290,In_677);
or U1388 (N_1388,In_320,In_13);
and U1389 (N_1389,In_457,In_8);
nor U1390 (N_1390,In_553,In_222);
nand U1391 (N_1391,In_534,In_270);
or U1392 (N_1392,In_173,In_560);
xor U1393 (N_1393,In_304,In_310);
or U1394 (N_1394,In_68,In_236);
nand U1395 (N_1395,In_632,In_224);
or U1396 (N_1396,In_681,In_155);
nand U1397 (N_1397,In_408,In_121);
and U1398 (N_1398,In_67,In_468);
xor U1399 (N_1399,In_720,In_31);
xor U1400 (N_1400,In_382,In_40);
or U1401 (N_1401,In_701,In_310);
nand U1402 (N_1402,In_543,In_417);
nor U1403 (N_1403,In_647,In_244);
nand U1404 (N_1404,In_579,In_61);
xor U1405 (N_1405,In_263,In_338);
nand U1406 (N_1406,In_174,In_727);
nand U1407 (N_1407,In_131,In_710);
nor U1408 (N_1408,In_188,In_578);
nand U1409 (N_1409,In_169,In_39);
and U1410 (N_1410,In_442,In_654);
nor U1411 (N_1411,In_530,In_552);
or U1412 (N_1412,In_675,In_83);
nor U1413 (N_1413,In_544,In_405);
or U1414 (N_1414,In_185,In_121);
or U1415 (N_1415,In_159,In_536);
xor U1416 (N_1416,In_701,In_623);
and U1417 (N_1417,In_55,In_604);
nor U1418 (N_1418,In_591,In_732);
nand U1419 (N_1419,In_149,In_481);
or U1420 (N_1420,In_305,In_9);
xnor U1421 (N_1421,In_10,In_621);
nor U1422 (N_1422,In_738,In_630);
and U1423 (N_1423,In_585,In_594);
xor U1424 (N_1424,In_464,In_244);
or U1425 (N_1425,In_419,In_539);
and U1426 (N_1426,In_467,In_94);
or U1427 (N_1427,In_459,In_556);
or U1428 (N_1428,In_270,In_304);
nor U1429 (N_1429,In_354,In_168);
nand U1430 (N_1430,In_461,In_104);
and U1431 (N_1431,In_314,In_257);
or U1432 (N_1432,In_295,In_545);
or U1433 (N_1433,In_690,In_544);
or U1434 (N_1434,In_1,In_619);
nand U1435 (N_1435,In_720,In_49);
or U1436 (N_1436,In_662,In_269);
or U1437 (N_1437,In_231,In_123);
nor U1438 (N_1438,In_554,In_334);
nand U1439 (N_1439,In_265,In_371);
xnor U1440 (N_1440,In_123,In_376);
nor U1441 (N_1441,In_64,In_366);
nand U1442 (N_1442,In_359,In_664);
nor U1443 (N_1443,In_629,In_712);
or U1444 (N_1444,In_83,In_691);
nor U1445 (N_1445,In_630,In_98);
nor U1446 (N_1446,In_375,In_688);
and U1447 (N_1447,In_93,In_228);
or U1448 (N_1448,In_420,In_274);
or U1449 (N_1449,In_56,In_692);
nor U1450 (N_1450,In_159,In_255);
or U1451 (N_1451,In_330,In_713);
nand U1452 (N_1452,In_653,In_153);
xnor U1453 (N_1453,In_713,In_145);
nor U1454 (N_1454,In_21,In_185);
and U1455 (N_1455,In_153,In_400);
nor U1456 (N_1456,In_115,In_132);
nor U1457 (N_1457,In_692,In_710);
nor U1458 (N_1458,In_639,In_380);
nor U1459 (N_1459,In_257,In_661);
or U1460 (N_1460,In_457,In_46);
or U1461 (N_1461,In_667,In_746);
nand U1462 (N_1462,In_682,In_557);
or U1463 (N_1463,In_343,In_358);
nor U1464 (N_1464,In_239,In_693);
or U1465 (N_1465,In_582,In_152);
or U1466 (N_1466,In_138,In_258);
and U1467 (N_1467,In_259,In_121);
and U1468 (N_1468,In_199,In_597);
and U1469 (N_1469,In_172,In_165);
nor U1470 (N_1470,In_31,In_499);
xor U1471 (N_1471,In_188,In_99);
or U1472 (N_1472,In_718,In_386);
xnor U1473 (N_1473,In_669,In_749);
and U1474 (N_1474,In_434,In_403);
and U1475 (N_1475,In_249,In_60);
and U1476 (N_1476,In_96,In_177);
nor U1477 (N_1477,In_696,In_590);
nor U1478 (N_1478,In_708,In_667);
nand U1479 (N_1479,In_264,In_708);
or U1480 (N_1480,In_182,In_551);
xnor U1481 (N_1481,In_389,In_239);
nor U1482 (N_1482,In_420,In_333);
xnor U1483 (N_1483,In_110,In_145);
nand U1484 (N_1484,In_264,In_294);
nand U1485 (N_1485,In_1,In_663);
or U1486 (N_1486,In_354,In_364);
nor U1487 (N_1487,In_638,In_485);
nor U1488 (N_1488,In_496,In_346);
nand U1489 (N_1489,In_470,In_202);
and U1490 (N_1490,In_565,In_419);
nor U1491 (N_1491,In_702,In_671);
or U1492 (N_1492,In_369,In_19);
or U1493 (N_1493,In_475,In_690);
xnor U1494 (N_1494,In_197,In_124);
nor U1495 (N_1495,In_185,In_593);
and U1496 (N_1496,In_238,In_568);
or U1497 (N_1497,In_154,In_747);
xor U1498 (N_1498,In_437,In_669);
or U1499 (N_1499,In_133,In_81);
and U1500 (N_1500,In_583,In_387);
nand U1501 (N_1501,In_294,In_640);
nor U1502 (N_1502,In_186,In_379);
nand U1503 (N_1503,In_396,In_127);
or U1504 (N_1504,In_139,In_541);
xor U1505 (N_1505,In_344,In_289);
or U1506 (N_1506,In_218,In_458);
and U1507 (N_1507,In_320,In_380);
and U1508 (N_1508,In_645,In_470);
nor U1509 (N_1509,In_432,In_416);
nand U1510 (N_1510,In_606,In_234);
or U1511 (N_1511,In_212,In_483);
nand U1512 (N_1512,In_685,In_22);
nand U1513 (N_1513,In_57,In_456);
nor U1514 (N_1514,In_447,In_572);
xnor U1515 (N_1515,In_542,In_415);
nor U1516 (N_1516,In_45,In_263);
and U1517 (N_1517,In_56,In_501);
and U1518 (N_1518,In_110,In_117);
xor U1519 (N_1519,In_273,In_410);
nand U1520 (N_1520,In_138,In_36);
nor U1521 (N_1521,In_131,In_153);
nor U1522 (N_1522,In_28,In_632);
nand U1523 (N_1523,In_100,In_316);
or U1524 (N_1524,In_248,In_246);
xnor U1525 (N_1525,In_505,In_21);
nand U1526 (N_1526,In_373,In_515);
nand U1527 (N_1527,In_499,In_210);
and U1528 (N_1528,In_36,In_64);
nor U1529 (N_1529,In_8,In_117);
nand U1530 (N_1530,In_736,In_409);
nand U1531 (N_1531,In_624,In_436);
nand U1532 (N_1532,In_597,In_610);
or U1533 (N_1533,In_250,In_27);
xnor U1534 (N_1534,In_97,In_537);
nor U1535 (N_1535,In_216,In_537);
and U1536 (N_1536,In_260,In_361);
xor U1537 (N_1537,In_174,In_688);
xor U1538 (N_1538,In_456,In_490);
or U1539 (N_1539,In_57,In_685);
nand U1540 (N_1540,In_351,In_7);
and U1541 (N_1541,In_217,In_639);
nor U1542 (N_1542,In_675,In_449);
and U1543 (N_1543,In_539,In_155);
nor U1544 (N_1544,In_317,In_521);
nand U1545 (N_1545,In_448,In_594);
nand U1546 (N_1546,In_359,In_501);
nor U1547 (N_1547,In_728,In_364);
nor U1548 (N_1548,In_258,In_657);
nor U1549 (N_1549,In_98,In_732);
and U1550 (N_1550,In_0,In_414);
and U1551 (N_1551,In_284,In_688);
and U1552 (N_1552,In_80,In_700);
xor U1553 (N_1553,In_585,In_80);
nand U1554 (N_1554,In_673,In_114);
and U1555 (N_1555,In_365,In_15);
nand U1556 (N_1556,In_653,In_353);
nor U1557 (N_1557,In_251,In_318);
and U1558 (N_1558,In_628,In_432);
or U1559 (N_1559,In_665,In_664);
nor U1560 (N_1560,In_631,In_417);
xor U1561 (N_1561,In_479,In_131);
nand U1562 (N_1562,In_427,In_326);
or U1563 (N_1563,In_23,In_500);
nand U1564 (N_1564,In_555,In_113);
nand U1565 (N_1565,In_624,In_201);
and U1566 (N_1566,In_693,In_400);
nand U1567 (N_1567,In_666,In_56);
or U1568 (N_1568,In_209,In_669);
nand U1569 (N_1569,In_746,In_62);
or U1570 (N_1570,In_156,In_640);
and U1571 (N_1571,In_272,In_737);
or U1572 (N_1572,In_367,In_627);
nand U1573 (N_1573,In_113,In_509);
xor U1574 (N_1574,In_312,In_655);
and U1575 (N_1575,In_14,In_230);
and U1576 (N_1576,In_434,In_628);
xor U1577 (N_1577,In_207,In_725);
nor U1578 (N_1578,In_678,In_132);
nand U1579 (N_1579,In_164,In_465);
or U1580 (N_1580,In_747,In_633);
and U1581 (N_1581,In_134,In_429);
and U1582 (N_1582,In_590,In_716);
xor U1583 (N_1583,In_409,In_671);
nand U1584 (N_1584,In_715,In_285);
nand U1585 (N_1585,In_511,In_663);
and U1586 (N_1586,In_147,In_99);
nand U1587 (N_1587,In_155,In_543);
or U1588 (N_1588,In_405,In_132);
nor U1589 (N_1589,In_249,In_258);
xor U1590 (N_1590,In_174,In_294);
or U1591 (N_1591,In_161,In_631);
or U1592 (N_1592,In_654,In_542);
or U1593 (N_1593,In_133,In_663);
and U1594 (N_1594,In_212,In_300);
nand U1595 (N_1595,In_352,In_355);
and U1596 (N_1596,In_52,In_341);
nor U1597 (N_1597,In_491,In_143);
or U1598 (N_1598,In_601,In_5);
nor U1599 (N_1599,In_383,In_547);
nor U1600 (N_1600,In_12,In_644);
or U1601 (N_1601,In_604,In_126);
or U1602 (N_1602,In_100,In_212);
nand U1603 (N_1603,In_630,In_366);
and U1604 (N_1604,In_528,In_347);
nor U1605 (N_1605,In_292,In_542);
nand U1606 (N_1606,In_747,In_726);
and U1607 (N_1607,In_302,In_36);
nor U1608 (N_1608,In_162,In_236);
and U1609 (N_1609,In_192,In_539);
or U1610 (N_1610,In_361,In_289);
and U1611 (N_1611,In_594,In_515);
nor U1612 (N_1612,In_209,In_470);
nor U1613 (N_1613,In_59,In_568);
or U1614 (N_1614,In_451,In_169);
or U1615 (N_1615,In_261,In_312);
nand U1616 (N_1616,In_86,In_14);
and U1617 (N_1617,In_332,In_353);
and U1618 (N_1618,In_525,In_65);
nor U1619 (N_1619,In_198,In_116);
or U1620 (N_1620,In_381,In_419);
nand U1621 (N_1621,In_223,In_568);
and U1622 (N_1622,In_296,In_473);
or U1623 (N_1623,In_52,In_97);
nor U1624 (N_1624,In_543,In_194);
nor U1625 (N_1625,In_638,In_459);
xor U1626 (N_1626,In_233,In_629);
and U1627 (N_1627,In_187,In_398);
nand U1628 (N_1628,In_166,In_13);
nor U1629 (N_1629,In_204,In_541);
or U1630 (N_1630,In_649,In_205);
nor U1631 (N_1631,In_321,In_607);
xor U1632 (N_1632,In_662,In_487);
nand U1633 (N_1633,In_293,In_531);
nand U1634 (N_1634,In_469,In_295);
nand U1635 (N_1635,In_559,In_384);
nor U1636 (N_1636,In_304,In_174);
or U1637 (N_1637,In_463,In_494);
xnor U1638 (N_1638,In_372,In_421);
nand U1639 (N_1639,In_112,In_201);
nand U1640 (N_1640,In_58,In_446);
and U1641 (N_1641,In_610,In_21);
and U1642 (N_1642,In_599,In_88);
and U1643 (N_1643,In_726,In_624);
xnor U1644 (N_1644,In_367,In_66);
nand U1645 (N_1645,In_606,In_703);
nand U1646 (N_1646,In_520,In_1);
or U1647 (N_1647,In_221,In_19);
or U1648 (N_1648,In_39,In_614);
nor U1649 (N_1649,In_25,In_37);
and U1650 (N_1650,In_152,In_184);
nor U1651 (N_1651,In_116,In_220);
and U1652 (N_1652,In_69,In_204);
and U1653 (N_1653,In_530,In_129);
or U1654 (N_1654,In_585,In_109);
nand U1655 (N_1655,In_678,In_519);
nor U1656 (N_1656,In_127,In_209);
xor U1657 (N_1657,In_433,In_679);
nand U1658 (N_1658,In_364,In_281);
xnor U1659 (N_1659,In_261,In_418);
or U1660 (N_1660,In_269,In_288);
xor U1661 (N_1661,In_367,In_248);
nand U1662 (N_1662,In_0,In_356);
and U1663 (N_1663,In_297,In_184);
and U1664 (N_1664,In_114,In_149);
nand U1665 (N_1665,In_376,In_400);
or U1666 (N_1666,In_657,In_212);
nor U1667 (N_1667,In_605,In_360);
or U1668 (N_1668,In_621,In_574);
nor U1669 (N_1669,In_259,In_532);
xor U1670 (N_1670,In_643,In_493);
nand U1671 (N_1671,In_55,In_267);
xnor U1672 (N_1672,In_614,In_507);
nor U1673 (N_1673,In_445,In_644);
or U1674 (N_1674,In_186,In_185);
nand U1675 (N_1675,In_153,In_562);
and U1676 (N_1676,In_609,In_516);
or U1677 (N_1677,In_125,In_679);
xnor U1678 (N_1678,In_368,In_229);
nand U1679 (N_1679,In_53,In_104);
nor U1680 (N_1680,In_471,In_352);
nand U1681 (N_1681,In_482,In_367);
nand U1682 (N_1682,In_171,In_686);
or U1683 (N_1683,In_482,In_529);
and U1684 (N_1684,In_459,In_542);
xnor U1685 (N_1685,In_362,In_660);
nor U1686 (N_1686,In_659,In_140);
nor U1687 (N_1687,In_438,In_386);
nor U1688 (N_1688,In_135,In_146);
nand U1689 (N_1689,In_331,In_239);
nor U1690 (N_1690,In_629,In_178);
nand U1691 (N_1691,In_275,In_27);
nor U1692 (N_1692,In_334,In_471);
nor U1693 (N_1693,In_268,In_131);
nor U1694 (N_1694,In_323,In_45);
nand U1695 (N_1695,In_464,In_471);
nor U1696 (N_1696,In_563,In_494);
or U1697 (N_1697,In_186,In_363);
or U1698 (N_1698,In_741,In_99);
nor U1699 (N_1699,In_641,In_70);
nor U1700 (N_1700,In_23,In_360);
nand U1701 (N_1701,In_450,In_132);
xor U1702 (N_1702,In_727,In_21);
nand U1703 (N_1703,In_202,In_312);
or U1704 (N_1704,In_335,In_311);
or U1705 (N_1705,In_528,In_97);
xor U1706 (N_1706,In_571,In_680);
nand U1707 (N_1707,In_266,In_676);
nor U1708 (N_1708,In_524,In_498);
and U1709 (N_1709,In_5,In_396);
and U1710 (N_1710,In_549,In_389);
nor U1711 (N_1711,In_550,In_162);
nand U1712 (N_1712,In_170,In_502);
nand U1713 (N_1713,In_114,In_481);
and U1714 (N_1714,In_367,In_736);
or U1715 (N_1715,In_404,In_402);
or U1716 (N_1716,In_497,In_233);
or U1717 (N_1717,In_441,In_84);
or U1718 (N_1718,In_613,In_391);
xnor U1719 (N_1719,In_19,In_137);
or U1720 (N_1720,In_181,In_460);
or U1721 (N_1721,In_611,In_380);
xnor U1722 (N_1722,In_739,In_274);
and U1723 (N_1723,In_207,In_590);
xnor U1724 (N_1724,In_159,In_408);
nor U1725 (N_1725,In_273,In_156);
nor U1726 (N_1726,In_195,In_703);
or U1727 (N_1727,In_146,In_172);
nand U1728 (N_1728,In_317,In_164);
and U1729 (N_1729,In_573,In_566);
nand U1730 (N_1730,In_259,In_674);
nand U1731 (N_1731,In_705,In_204);
nand U1732 (N_1732,In_501,In_191);
or U1733 (N_1733,In_238,In_392);
or U1734 (N_1734,In_376,In_80);
nand U1735 (N_1735,In_476,In_80);
xnor U1736 (N_1736,In_259,In_580);
nor U1737 (N_1737,In_196,In_201);
nand U1738 (N_1738,In_497,In_468);
or U1739 (N_1739,In_114,In_120);
and U1740 (N_1740,In_673,In_580);
or U1741 (N_1741,In_47,In_229);
or U1742 (N_1742,In_483,In_487);
or U1743 (N_1743,In_538,In_431);
nand U1744 (N_1744,In_194,In_62);
or U1745 (N_1745,In_237,In_8);
nand U1746 (N_1746,In_538,In_327);
or U1747 (N_1747,In_473,In_666);
nor U1748 (N_1748,In_334,In_61);
nor U1749 (N_1749,In_9,In_108);
nand U1750 (N_1750,In_601,In_266);
nor U1751 (N_1751,In_482,In_448);
nand U1752 (N_1752,In_610,In_416);
and U1753 (N_1753,In_111,In_708);
nor U1754 (N_1754,In_734,In_208);
nor U1755 (N_1755,In_642,In_465);
nor U1756 (N_1756,In_356,In_313);
nand U1757 (N_1757,In_638,In_548);
nand U1758 (N_1758,In_139,In_234);
nor U1759 (N_1759,In_5,In_687);
nor U1760 (N_1760,In_372,In_577);
and U1761 (N_1761,In_225,In_630);
or U1762 (N_1762,In_726,In_207);
and U1763 (N_1763,In_26,In_668);
or U1764 (N_1764,In_124,In_456);
or U1765 (N_1765,In_267,In_469);
xor U1766 (N_1766,In_78,In_173);
nor U1767 (N_1767,In_233,In_486);
and U1768 (N_1768,In_67,In_97);
nand U1769 (N_1769,In_94,In_364);
nor U1770 (N_1770,In_44,In_230);
or U1771 (N_1771,In_37,In_701);
xnor U1772 (N_1772,In_697,In_10);
or U1773 (N_1773,In_702,In_112);
or U1774 (N_1774,In_297,In_697);
nor U1775 (N_1775,In_472,In_36);
and U1776 (N_1776,In_739,In_440);
nand U1777 (N_1777,In_530,In_356);
or U1778 (N_1778,In_81,In_651);
nand U1779 (N_1779,In_343,In_435);
nand U1780 (N_1780,In_251,In_436);
and U1781 (N_1781,In_727,In_350);
nand U1782 (N_1782,In_450,In_140);
and U1783 (N_1783,In_712,In_433);
and U1784 (N_1784,In_545,In_572);
nand U1785 (N_1785,In_299,In_528);
or U1786 (N_1786,In_301,In_578);
nand U1787 (N_1787,In_231,In_681);
nor U1788 (N_1788,In_24,In_268);
and U1789 (N_1789,In_437,In_423);
nand U1790 (N_1790,In_658,In_545);
or U1791 (N_1791,In_538,In_204);
or U1792 (N_1792,In_403,In_416);
nand U1793 (N_1793,In_219,In_9);
and U1794 (N_1794,In_97,In_1);
nor U1795 (N_1795,In_93,In_634);
nor U1796 (N_1796,In_83,In_705);
nand U1797 (N_1797,In_375,In_206);
nor U1798 (N_1798,In_293,In_77);
xor U1799 (N_1799,In_749,In_434);
nand U1800 (N_1800,In_599,In_305);
and U1801 (N_1801,In_726,In_509);
nor U1802 (N_1802,In_665,In_567);
nand U1803 (N_1803,In_638,In_376);
nor U1804 (N_1804,In_339,In_586);
or U1805 (N_1805,In_432,In_564);
nor U1806 (N_1806,In_257,In_152);
and U1807 (N_1807,In_194,In_446);
or U1808 (N_1808,In_251,In_95);
nand U1809 (N_1809,In_82,In_736);
and U1810 (N_1810,In_501,In_578);
nor U1811 (N_1811,In_250,In_400);
nor U1812 (N_1812,In_98,In_532);
or U1813 (N_1813,In_587,In_232);
nor U1814 (N_1814,In_734,In_291);
or U1815 (N_1815,In_686,In_547);
nand U1816 (N_1816,In_687,In_219);
nor U1817 (N_1817,In_41,In_397);
or U1818 (N_1818,In_20,In_139);
or U1819 (N_1819,In_446,In_479);
nor U1820 (N_1820,In_748,In_72);
and U1821 (N_1821,In_509,In_345);
nor U1822 (N_1822,In_316,In_722);
and U1823 (N_1823,In_696,In_650);
nor U1824 (N_1824,In_729,In_231);
and U1825 (N_1825,In_72,In_403);
nor U1826 (N_1826,In_475,In_126);
nor U1827 (N_1827,In_387,In_685);
nor U1828 (N_1828,In_121,In_650);
and U1829 (N_1829,In_652,In_376);
or U1830 (N_1830,In_204,In_256);
xor U1831 (N_1831,In_163,In_622);
or U1832 (N_1832,In_734,In_150);
and U1833 (N_1833,In_600,In_267);
and U1834 (N_1834,In_46,In_233);
or U1835 (N_1835,In_372,In_620);
xnor U1836 (N_1836,In_717,In_699);
nor U1837 (N_1837,In_70,In_269);
or U1838 (N_1838,In_244,In_499);
nand U1839 (N_1839,In_407,In_67);
xor U1840 (N_1840,In_327,In_152);
and U1841 (N_1841,In_604,In_742);
and U1842 (N_1842,In_192,In_70);
or U1843 (N_1843,In_49,In_112);
nor U1844 (N_1844,In_692,In_676);
xor U1845 (N_1845,In_360,In_197);
xor U1846 (N_1846,In_732,In_285);
or U1847 (N_1847,In_269,In_135);
xor U1848 (N_1848,In_177,In_708);
nand U1849 (N_1849,In_243,In_525);
nand U1850 (N_1850,In_14,In_360);
nor U1851 (N_1851,In_121,In_685);
or U1852 (N_1852,In_123,In_26);
and U1853 (N_1853,In_432,In_198);
nand U1854 (N_1854,In_360,In_694);
or U1855 (N_1855,In_603,In_565);
or U1856 (N_1856,In_679,In_698);
nand U1857 (N_1857,In_205,In_476);
nand U1858 (N_1858,In_657,In_581);
and U1859 (N_1859,In_294,In_589);
nor U1860 (N_1860,In_168,In_328);
nor U1861 (N_1861,In_282,In_386);
and U1862 (N_1862,In_193,In_52);
and U1863 (N_1863,In_485,In_504);
nor U1864 (N_1864,In_305,In_218);
nor U1865 (N_1865,In_361,In_714);
nor U1866 (N_1866,In_329,In_323);
or U1867 (N_1867,In_283,In_155);
and U1868 (N_1868,In_682,In_60);
xnor U1869 (N_1869,In_737,In_423);
and U1870 (N_1870,In_366,In_241);
and U1871 (N_1871,In_591,In_242);
and U1872 (N_1872,In_30,In_603);
nand U1873 (N_1873,In_659,In_514);
and U1874 (N_1874,In_70,In_623);
and U1875 (N_1875,In_267,In_307);
or U1876 (N_1876,In_544,In_444);
xor U1877 (N_1877,In_421,In_570);
xnor U1878 (N_1878,In_354,In_163);
nor U1879 (N_1879,In_269,In_478);
and U1880 (N_1880,In_738,In_551);
nor U1881 (N_1881,In_187,In_513);
nor U1882 (N_1882,In_387,In_580);
nand U1883 (N_1883,In_159,In_110);
xnor U1884 (N_1884,In_10,In_192);
nor U1885 (N_1885,In_648,In_108);
xnor U1886 (N_1886,In_208,In_735);
or U1887 (N_1887,In_415,In_17);
nand U1888 (N_1888,In_595,In_671);
or U1889 (N_1889,In_73,In_110);
and U1890 (N_1890,In_279,In_287);
or U1891 (N_1891,In_305,In_669);
nand U1892 (N_1892,In_508,In_277);
or U1893 (N_1893,In_340,In_684);
or U1894 (N_1894,In_349,In_551);
and U1895 (N_1895,In_632,In_399);
nand U1896 (N_1896,In_476,In_384);
nand U1897 (N_1897,In_656,In_115);
nor U1898 (N_1898,In_528,In_355);
and U1899 (N_1899,In_641,In_347);
nor U1900 (N_1900,In_723,In_385);
or U1901 (N_1901,In_76,In_654);
nand U1902 (N_1902,In_731,In_427);
or U1903 (N_1903,In_685,In_231);
nand U1904 (N_1904,In_248,In_391);
and U1905 (N_1905,In_135,In_51);
xnor U1906 (N_1906,In_528,In_469);
or U1907 (N_1907,In_113,In_691);
nand U1908 (N_1908,In_36,In_161);
nor U1909 (N_1909,In_391,In_252);
and U1910 (N_1910,In_533,In_630);
nor U1911 (N_1911,In_520,In_291);
nand U1912 (N_1912,In_446,In_100);
and U1913 (N_1913,In_554,In_30);
and U1914 (N_1914,In_574,In_267);
or U1915 (N_1915,In_382,In_538);
nor U1916 (N_1916,In_250,In_665);
nor U1917 (N_1917,In_475,In_275);
nor U1918 (N_1918,In_234,In_420);
and U1919 (N_1919,In_211,In_642);
or U1920 (N_1920,In_683,In_286);
nand U1921 (N_1921,In_726,In_737);
or U1922 (N_1922,In_567,In_274);
nor U1923 (N_1923,In_240,In_469);
and U1924 (N_1924,In_672,In_549);
nor U1925 (N_1925,In_344,In_308);
xor U1926 (N_1926,In_685,In_708);
nand U1927 (N_1927,In_361,In_115);
nor U1928 (N_1928,In_297,In_601);
or U1929 (N_1929,In_563,In_597);
or U1930 (N_1930,In_551,In_10);
and U1931 (N_1931,In_18,In_58);
or U1932 (N_1932,In_31,In_675);
nor U1933 (N_1933,In_20,In_442);
nor U1934 (N_1934,In_199,In_671);
nor U1935 (N_1935,In_497,In_593);
nor U1936 (N_1936,In_2,In_662);
and U1937 (N_1937,In_505,In_739);
nand U1938 (N_1938,In_210,In_218);
and U1939 (N_1939,In_239,In_254);
nand U1940 (N_1940,In_468,In_205);
nand U1941 (N_1941,In_46,In_595);
nand U1942 (N_1942,In_711,In_576);
or U1943 (N_1943,In_126,In_41);
or U1944 (N_1944,In_647,In_66);
nand U1945 (N_1945,In_569,In_743);
nand U1946 (N_1946,In_268,In_398);
xnor U1947 (N_1947,In_705,In_21);
nand U1948 (N_1948,In_377,In_424);
nand U1949 (N_1949,In_712,In_146);
and U1950 (N_1950,In_727,In_184);
nand U1951 (N_1951,In_694,In_395);
or U1952 (N_1952,In_573,In_621);
xor U1953 (N_1953,In_532,In_607);
or U1954 (N_1954,In_305,In_221);
and U1955 (N_1955,In_310,In_300);
nor U1956 (N_1956,In_87,In_650);
nand U1957 (N_1957,In_59,In_708);
nand U1958 (N_1958,In_631,In_690);
or U1959 (N_1959,In_179,In_516);
nand U1960 (N_1960,In_722,In_253);
nand U1961 (N_1961,In_390,In_323);
nand U1962 (N_1962,In_569,In_198);
or U1963 (N_1963,In_339,In_508);
nand U1964 (N_1964,In_97,In_285);
and U1965 (N_1965,In_595,In_483);
and U1966 (N_1966,In_725,In_197);
nand U1967 (N_1967,In_562,In_663);
nor U1968 (N_1968,In_103,In_461);
and U1969 (N_1969,In_244,In_433);
nor U1970 (N_1970,In_699,In_610);
nand U1971 (N_1971,In_277,In_31);
nand U1972 (N_1972,In_164,In_538);
xor U1973 (N_1973,In_104,In_15);
xnor U1974 (N_1974,In_597,In_253);
nand U1975 (N_1975,In_275,In_244);
or U1976 (N_1976,In_583,In_433);
and U1977 (N_1977,In_483,In_686);
and U1978 (N_1978,In_623,In_318);
and U1979 (N_1979,In_279,In_728);
and U1980 (N_1980,In_645,In_543);
nand U1981 (N_1981,In_407,In_324);
or U1982 (N_1982,In_684,In_404);
nand U1983 (N_1983,In_36,In_410);
or U1984 (N_1984,In_145,In_555);
and U1985 (N_1985,In_728,In_415);
nand U1986 (N_1986,In_303,In_639);
and U1987 (N_1987,In_206,In_470);
or U1988 (N_1988,In_478,In_412);
or U1989 (N_1989,In_373,In_319);
and U1990 (N_1990,In_564,In_278);
or U1991 (N_1991,In_8,In_381);
xnor U1992 (N_1992,In_698,In_685);
nor U1993 (N_1993,In_500,In_438);
or U1994 (N_1994,In_196,In_519);
or U1995 (N_1995,In_420,In_190);
nand U1996 (N_1996,In_165,In_94);
nand U1997 (N_1997,In_211,In_431);
nand U1998 (N_1998,In_641,In_138);
or U1999 (N_1999,In_64,In_360);
nor U2000 (N_2000,In_532,In_243);
nor U2001 (N_2001,In_314,In_266);
nand U2002 (N_2002,In_483,In_76);
or U2003 (N_2003,In_223,In_14);
nand U2004 (N_2004,In_683,In_71);
nand U2005 (N_2005,In_729,In_309);
or U2006 (N_2006,In_48,In_99);
nand U2007 (N_2007,In_361,In_423);
and U2008 (N_2008,In_146,In_106);
nand U2009 (N_2009,In_284,In_299);
or U2010 (N_2010,In_262,In_238);
nand U2011 (N_2011,In_400,In_101);
nor U2012 (N_2012,In_726,In_264);
xor U2013 (N_2013,In_95,In_642);
and U2014 (N_2014,In_412,In_133);
xor U2015 (N_2015,In_82,In_153);
nor U2016 (N_2016,In_87,In_637);
xnor U2017 (N_2017,In_739,In_712);
nand U2018 (N_2018,In_636,In_44);
and U2019 (N_2019,In_594,In_306);
or U2020 (N_2020,In_596,In_372);
nand U2021 (N_2021,In_210,In_246);
nor U2022 (N_2022,In_558,In_45);
or U2023 (N_2023,In_360,In_615);
or U2024 (N_2024,In_569,In_708);
or U2025 (N_2025,In_625,In_20);
or U2026 (N_2026,In_449,In_658);
nand U2027 (N_2027,In_138,In_334);
or U2028 (N_2028,In_714,In_194);
and U2029 (N_2029,In_606,In_175);
and U2030 (N_2030,In_500,In_185);
and U2031 (N_2031,In_119,In_121);
nor U2032 (N_2032,In_582,In_497);
and U2033 (N_2033,In_745,In_285);
xnor U2034 (N_2034,In_579,In_55);
or U2035 (N_2035,In_725,In_460);
nand U2036 (N_2036,In_479,In_384);
nand U2037 (N_2037,In_417,In_484);
and U2038 (N_2038,In_572,In_318);
and U2039 (N_2039,In_19,In_503);
xor U2040 (N_2040,In_53,In_418);
or U2041 (N_2041,In_13,In_698);
nand U2042 (N_2042,In_483,In_25);
or U2043 (N_2043,In_507,In_635);
nand U2044 (N_2044,In_733,In_535);
or U2045 (N_2045,In_293,In_535);
nor U2046 (N_2046,In_667,In_642);
xor U2047 (N_2047,In_286,In_679);
or U2048 (N_2048,In_636,In_123);
xnor U2049 (N_2049,In_161,In_622);
nor U2050 (N_2050,In_586,In_328);
or U2051 (N_2051,In_89,In_683);
nor U2052 (N_2052,In_706,In_416);
or U2053 (N_2053,In_452,In_373);
nand U2054 (N_2054,In_559,In_740);
and U2055 (N_2055,In_560,In_685);
and U2056 (N_2056,In_517,In_87);
nand U2057 (N_2057,In_696,In_289);
and U2058 (N_2058,In_410,In_236);
nor U2059 (N_2059,In_587,In_148);
and U2060 (N_2060,In_544,In_324);
or U2061 (N_2061,In_210,In_295);
nor U2062 (N_2062,In_28,In_311);
nand U2063 (N_2063,In_706,In_50);
nand U2064 (N_2064,In_503,In_226);
or U2065 (N_2065,In_585,In_25);
nand U2066 (N_2066,In_284,In_171);
xnor U2067 (N_2067,In_665,In_523);
and U2068 (N_2068,In_200,In_730);
nor U2069 (N_2069,In_157,In_576);
and U2070 (N_2070,In_472,In_644);
nand U2071 (N_2071,In_361,In_675);
nor U2072 (N_2072,In_125,In_217);
and U2073 (N_2073,In_152,In_654);
nor U2074 (N_2074,In_679,In_173);
nor U2075 (N_2075,In_695,In_549);
or U2076 (N_2076,In_216,In_359);
or U2077 (N_2077,In_495,In_531);
nand U2078 (N_2078,In_247,In_160);
and U2079 (N_2079,In_229,In_190);
and U2080 (N_2080,In_14,In_655);
nor U2081 (N_2081,In_520,In_554);
nand U2082 (N_2082,In_503,In_374);
and U2083 (N_2083,In_516,In_156);
nand U2084 (N_2084,In_384,In_13);
and U2085 (N_2085,In_283,In_152);
nand U2086 (N_2086,In_635,In_352);
and U2087 (N_2087,In_404,In_258);
or U2088 (N_2088,In_150,In_354);
and U2089 (N_2089,In_619,In_142);
and U2090 (N_2090,In_659,In_420);
nor U2091 (N_2091,In_157,In_27);
nor U2092 (N_2092,In_419,In_505);
or U2093 (N_2093,In_79,In_368);
xor U2094 (N_2094,In_655,In_455);
nor U2095 (N_2095,In_647,In_271);
nand U2096 (N_2096,In_692,In_228);
nand U2097 (N_2097,In_258,In_92);
nand U2098 (N_2098,In_406,In_747);
and U2099 (N_2099,In_622,In_522);
and U2100 (N_2100,In_271,In_592);
xnor U2101 (N_2101,In_10,In_695);
nor U2102 (N_2102,In_586,In_584);
or U2103 (N_2103,In_96,In_42);
nand U2104 (N_2104,In_352,In_65);
nand U2105 (N_2105,In_436,In_137);
or U2106 (N_2106,In_64,In_251);
and U2107 (N_2107,In_124,In_25);
and U2108 (N_2108,In_617,In_79);
and U2109 (N_2109,In_150,In_30);
and U2110 (N_2110,In_644,In_281);
and U2111 (N_2111,In_248,In_399);
nand U2112 (N_2112,In_407,In_158);
nor U2113 (N_2113,In_27,In_289);
and U2114 (N_2114,In_88,In_207);
nor U2115 (N_2115,In_536,In_670);
or U2116 (N_2116,In_636,In_54);
nand U2117 (N_2117,In_597,In_115);
or U2118 (N_2118,In_421,In_343);
and U2119 (N_2119,In_697,In_288);
nand U2120 (N_2120,In_67,In_136);
or U2121 (N_2121,In_190,In_192);
nor U2122 (N_2122,In_223,In_57);
or U2123 (N_2123,In_394,In_605);
nand U2124 (N_2124,In_29,In_132);
nand U2125 (N_2125,In_652,In_549);
nand U2126 (N_2126,In_45,In_374);
nor U2127 (N_2127,In_738,In_181);
nand U2128 (N_2128,In_419,In_59);
or U2129 (N_2129,In_738,In_280);
nor U2130 (N_2130,In_168,In_266);
or U2131 (N_2131,In_283,In_307);
xor U2132 (N_2132,In_271,In_45);
nor U2133 (N_2133,In_3,In_341);
xor U2134 (N_2134,In_437,In_98);
nor U2135 (N_2135,In_3,In_18);
and U2136 (N_2136,In_143,In_352);
nand U2137 (N_2137,In_289,In_1);
nand U2138 (N_2138,In_335,In_231);
nor U2139 (N_2139,In_578,In_382);
and U2140 (N_2140,In_159,In_625);
xnor U2141 (N_2141,In_682,In_440);
and U2142 (N_2142,In_334,In_214);
nor U2143 (N_2143,In_509,In_293);
or U2144 (N_2144,In_75,In_304);
nor U2145 (N_2145,In_624,In_525);
nand U2146 (N_2146,In_430,In_479);
and U2147 (N_2147,In_75,In_722);
and U2148 (N_2148,In_347,In_300);
nand U2149 (N_2149,In_534,In_325);
nor U2150 (N_2150,In_591,In_97);
nand U2151 (N_2151,In_285,In_408);
or U2152 (N_2152,In_316,In_179);
nor U2153 (N_2153,In_10,In_683);
and U2154 (N_2154,In_378,In_391);
or U2155 (N_2155,In_268,In_273);
and U2156 (N_2156,In_617,In_25);
and U2157 (N_2157,In_371,In_592);
nor U2158 (N_2158,In_482,In_140);
or U2159 (N_2159,In_109,In_620);
or U2160 (N_2160,In_409,In_128);
and U2161 (N_2161,In_374,In_58);
and U2162 (N_2162,In_284,In_390);
nand U2163 (N_2163,In_305,In_252);
nand U2164 (N_2164,In_705,In_635);
nand U2165 (N_2165,In_283,In_86);
nand U2166 (N_2166,In_443,In_456);
or U2167 (N_2167,In_215,In_167);
or U2168 (N_2168,In_645,In_273);
nand U2169 (N_2169,In_206,In_80);
or U2170 (N_2170,In_74,In_265);
and U2171 (N_2171,In_252,In_636);
nand U2172 (N_2172,In_523,In_231);
xor U2173 (N_2173,In_44,In_556);
nand U2174 (N_2174,In_625,In_333);
and U2175 (N_2175,In_373,In_46);
nor U2176 (N_2176,In_229,In_491);
and U2177 (N_2177,In_223,In_172);
and U2178 (N_2178,In_355,In_264);
and U2179 (N_2179,In_542,In_691);
or U2180 (N_2180,In_489,In_157);
and U2181 (N_2181,In_730,In_19);
and U2182 (N_2182,In_630,In_202);
and U2183 (N_2183,In_705,In_275);
and U2184 (N_2184,In_60,In_471);
or U2185 (N_2185,In_697,In_380);
or U2186 (N_2186,In_535,In_422);
nand U2187 (N_2187,In_69,In_608);
nand U2188 (N_2188,In_11,In_667);
nand U2189 (N_2189,In_192,In_711);
nor U2190 (N_2190,In_117,In_525);
and U2191 (N_2191,In_462,In_1);
and U2192 (N_2192,In_232,In_410);
nor U2193 (N_2193,In_365,In_682);
nor U2194 (N_2194,In_42,In_435);
nand U2195 (N_2195,In_342,In_680);
or U2196 (N_2196,In_26,In_32);
nand U2197 (N_2197,In_94,In_64);
xor U2198 (N_2198,In_13,In_363);
xor U2199 (N_2199,In_452,In_276);
or U2200 (N_2200,In_82,In_496);
and U2201 (N_2201,In_495,In_509);
nand U2202 (N_2202,In_699,In_734);
or U2203 (N_2203,In_60,In_719);
and U2204 (N_2204,In_639,In_744);
nor U2205 (N_2205,In_474,In_347);
nand U2206 (N_2206,In_530,In_632);
and U2207 (N_2207,In_617,In_730);
nor U2208 (N_2208,In_11,In_632);
nor U2209 (N_2209,In_52,In_74);
nor U2210 (N_2210,In_362,In_401);
nor U2211 (N_2211,In_644,In_222);
nand U2212 (N_2212,In_6,In_287);
nor U2213 (N_2213,In_509,In_73);
nor U2214 (N_2214,In_37,In_403);
or U2215 (N_2215,In_71,In_299);
nor U2216 (N_2216,In_443,In_701);
and U2217 (N_2217,In_649,In_384);
xnor U2218 (N_2218,In_434,In_242);
or U2219 (N_2219,In_525,In_348);
nand U2220 (N_2220,In_235,In_726);
xnor U2221 (N_2221,In_547,In_477);
or U2222 (N_2222,In_413,In_720);
or U2223 (N_2223,In_616,In_571);
nand U2224 (N_2224,In_517,In_619);
nand U2225 (N_2225,In_295,In_269);
nand U2226 (N_2226,In_292,In_559);
or U2227 (N_2227,In_18,In_521);
nand U2228 (N_2228,In_445,In_189);
and U2229 (N_2229,In_257,In_87);
or U2230 (N_2230,In_393,In_736);
and U2231 (N_2231,In_391,In_13);
nand U2232 (N_2232,In_693,In_630);
and U2233 (N_2233,In_344,In_502);
and U2234 (N_2234,In_315,In_431);
nor U2235 (N_2235,In_313,In_610);
xor U2236 (N_2236,In_283,In_561);
nor U2237 (N_2237,In_577,In_187);
nor U2238 (N_2238,In_406,In_547);
or U2239 (N_2239,In_574,In_375);
nor U2240 (N_2240,In_45,In_301);
xor U2241 (N_2241,In_206,In_100);
nand U2242 (N_2242,In_392,In_174);
nand U2243 (N_2243,In_631,In_443);
or U2244 (N_2244,In_298,In_24);
xnor U2245 (N_2245,In_70,In_91);
nand U2246 (N_2246,In_680,In_397);
nand U2247 (N_2247,In_233,In_493);
nor U2248 (N_2248,In_632,In_466);
xnor U2249 (N_2249,In_692,In_671);
nand U2250 (N_2250,In_548,In_187);
xor U2251 (N_2251,In_701,In_542);
nor U2252 (N_2252,In_612,In_620);
or U2253 (N_2253,In_507,In_390);
nor U2254 (N_2254,In_218,In_11);
nand U2255 (N_2255,In_28,In_510);
and U2256 (N_2256,In_682,In_167);
nor U2257 (N_2257,In_26,In_37);
nor U2258 (N_2258,In_740,In_609);
xnor U2259 (N_2259,In_667,In_239);
and U2260 (N_2260,In_634,In_295);
or U2261 (N_2261,In_273,In_137);
nand U2262 (N_2262,In_203,In_72);
and U2263 (N_2263,In_618,In_123);
nand U2264 (N_2264,In_200,In_93);
nor U2265 (N_2265,In_276,In_463);
nand U2266 (N_2266,In_296,In_457);
or U2267 (N_2267,In_402,In_287);
and U2268 (N_2268,In_6,In_455);
xor U2269 (N_2269,In_334,In_309);
nand U2270 (N_2270,In_451,In_145);
nand U2271 (N_2271,In_388,In_110);
and U2272 (N_2272,In_555,In_653);
nor U2273 (N_2273,In_505,In_376);
nand U2274 (N_2274,In_359,In_546);
and U2275 (N_2275,In_713,In_132);
and U2276 (N_2276,In_347,In_703);
or U2277 (N_2277,In_413,In_247);
nor U2278 (N_2278,In_153,In_236);
nor U2279 (N_2279,In_377,In_136);
nor U2280 (N_2280,In_617,In_722);
and U2281 (N_2281,In_93,In_607);
and U2282 (N_2282,In_264,In_106);
or U2283 (N_2283,In_719,In_609);
and U2284 (N_2284,In_737,In_655);
nand U2285 (N_2285,In_90,In_695);
nor U2286 (N_2286,In_109,In_270);
and U2287 (N_2287,In_703,In_235);
nor U2288 (N_2288,In_319,In_152);
and U2289 (N_2289,In_660,In_554);
nand U2290 (N_2290,In_514,In_656);
nor U2291 (N_2291,In_306,In_711);
nor U2292 (N_2292,In_614,In_328);
or U2293 (N_2293,In_645,In_310);
or U2294 (N_2294,In_6,In_609);
xnor U2295 (N_2295,In_401,In_628);
nor U2296 (N_2296,In_440,In_116);
xor U2297 (N_2297,In_393,In_298);
nand U2298 (N_2298,In_679,In_335);
nor U2299 (N_2299,In_441,In_264);
or U2300 (N_2300,In_588,In_396);
nor U2301 (N_2301,In_683,In_525);
nor U2302 (N_2302,In_148,In_665);
nand U2303 (N_2303,In_169,In_732);
nand U2304 (N_2304,In_263,In_698);
nor U2305 (N_2305,In_325,In_285);
xor U2306 (N_2306,In_540,In_198);
and U2307 (N_2307,In_522,In_669);
nand U2308 (N_2308,In_132,In_706);
nor U2309 (N_2309,In_556,In_733);
or U2310 (N_2310,In_126,In_557);
nor U2311 (N_2311,In_389,In_417);
and U2312 (N_2312,In_6,In_548);
or U2313 (N_2313,In_634,In_481);
nand U2314 (N_2314,In_613,In_527);
nand U2315 (N_2315,In_649,In_152);
nor U2316 (N_2316,In_147,In_58);
nor U2317 (N_2317,In_622,In_551);
nor U2318 (N_2318,In_363,In_145);
xnor U2319 (N_2319,In_388,In_615);
nor U2320 (N_2320,In_479,In_53);
or U2321 (N_2321,In_474,In_231);
xor U2322 (N_2322,In_293,In_311);
nor U2323 (N_2323,In_283,In_266);
and U2324 (N_2324,In_177,In_390);
nand U2325 (N_2325,In_438,In_68);
or U2326 (N_2326,In_747,In_42);
or U2327 (N_2327,In_477,In_685);
nor U2328 (N_2328,In_706,In_478);
and U2329 (N_2329,In_724,In_587);
and U2330 (N_2330,In_99,In_543);
or U2331 (N_2331,In_233,In_478);
and U2332 (N_2332,In_458,In_34);
xor U2333 (N_2333,In_643,In_458);
and U2334 (N_2334,In_588,In_24);
nand U2335 (N_2335,In_688,In_510);
and U2336 (N_2336,In_325,In_565);
nand U2337 (N_2337,In_688,In_386);
nor U2338 (N_2338,In_446,In_346);
xor U2339 (N_2339,In_509,In_701);
nand U2340 (N_2340,In_579,In_65);
nor U2341 (N_2341,In_12,In_170);
nor U2342 (N_2342,In_686,In_413);
or U2343 (N_2343,In_584,In_322);
nor U2344 (N_2344,In_44,In_537);
nor U2345 (N_2345,In_410,In_643);
nand U2346 (N_2346,In_508,In_438);
or U2347 (N_2347,In_552,In_272);
or U2348 (N_2348,In_354,In_164);
nand U2349 (N_2349,In_497,In_571);
nor U2350 (N_2350,In_140,In_80);
or U2351 (N_2351,In_686,In_57);
and U2352 (N_2352,In_647,In_92);
nor U2353 (N_2353,In_23,In_738);
nor U2354 (N_2354,In_612,In_481);
and U2355 (N_2355,In_19,In_605);
or U2356 (N_2356,In_9,In_410);
nor U2357 (N_2357,In_461,In_405);
xor U2358 (N_2358,In_385,In_220);
nand U2359 (N_2359,In_392,In_509);
and U2360 (N_2360,In_80,In_652);
nor U2361 (N_2361,In_250,In_127);
or U2362 (N_2362,In_118,In_716);
or U2363 (N_2363,In_564,In_48);
nor U2364 (N_2364,In_318,In_189);
and U2365 (N_2365,In_441,In_305);
nor U2366 (N_2366,In_326,In_178);
nand U2367 (N_2367,In_574,In_40);
xnor U2368 (N_2368,In_261,In_4);
xnor U2369 (N_2369,In_601,In_9);
or U2370 (N_2370,In_347,In_418);
and U2371 (N_2371,In_137,In_652);
nand U2372 (N_2372,In_626,In_406);
and U2373 (N_2373,In_1,In_501);
and U2374 (N_2374,In_304,In_57);
nor U2375 (N_2375,In_674,In_94);
or U2376 (N_2376,In_150,In_123);
nand U2377 (N_2377,In_3,In_11);
nand U2378 (N_2378,In_390,In_139);
nand U2379 (N_2379,In_365,In_286);
nand U2380 (N_2380,In_241,In_81);
nor U2381 (N_2381,In_450,In_632);
nand U2382 (N_2382,In_724,In_736);
nand U2383 (N_2383,In_147,In_36);
nand U2384 (N_2384,In_696,In_648);
nand U2385 (N_2385,In_43,In_87);
nor U2386 (N_2386,In_121,In_639);
or U2387 (N_2387,In_412,In_85);
xor U2388 (N_2388,In_359,In_699);
and U2389 (N_2389,In_439,In_255);
xnor U2390 (N_2390,In_575,In_255);
and U2391 (N_2391,In_61,In_384);
or U2392 (N_2392,In_522,In_532);
nor U2393 (N_2393,In_749,In_90);
or U2394 (N_2394,In_494,In_695);
and U2395 (N_2395,In_55,In_577);
nand U2396 (N_2396,In_444,In_522);
xor U2397 (N_2397,In_704,In_104);
and U2398 (N_2398,In_373,In_289);
and U2399 (N_2399,In_341,In_339);
nand U2400 (N_2400,In_287,In_565);
or U2401 (N_2401,In_452,In_309);
nor U2402 (N_2402,In_590,In_549);
nor U2403 (N_2403,In_568,In_166);
or U2404 (N_2404,In_319,In_412);
nor U2405 (N_2405,In_545,In_208);
xor U2406 (N_2406,In_274,In_49);
nand U2407 (N_2407,In_223,In_453);
nor U2408 (N_2408,In_103,In_452);
xnor U2409 (N_2409,In_53,In_29);
nor U2410 (N_2410,In_697,In_0);
or U2411 (N_2411,In_366,In_286);
and U2412 (N_2412,In_69,In_408);
or U2413 (N_2413,In_17,In_670);
or U2414 (N_2414,In_58,In_508);
and U2415 (N_2415,In_27,In_110);
or U2416 (N_2416,In_463,In_59);
nor U2417 (N_2417,In_68,In_617);
nand U2418 (N_2418,In_359,In_667);
nor U2419 (N_2419,In_275,In_339);
xnor U2420 (N_2420,In_252,In_287);
xor U2421 (N_2421,In_158,In_477);
nand U2422 (N_2422,In_249,In_405);
or U2423 (N_2423,In_419,In_373);
or U2424 (N_2424,In_117,In_527);
nand U2425 (N_2425,In_18,In_20);
or U2426 (N_2426,In_129,In_4);
and U2427 (N_2427,In_685,In_203);
or U2428 (N_2428,In_164,In_228);
and U2429 (N_2429,In_357,In_637);
nor U2430 (N_2430,In_248,In_316);
nor U2431 (N_2431,In_741,In_352);
xnor U2432 (N_2432,In_69,In_221);
nand U2433 (N_2433,In_156,In_21);
nor U2434 (N_2434,In_87,In_180);
and U2435 (N_2435,In_632,In_251);
nand U2436 (N_2436,In_265,In_276);
and U2437 (N_2437,In_88,In_138);
nand U2438 (N_2438,In_498,In_309);
nand U2439 (N_2439,In_376,In_74);
nor U2440 (N_2440,In_53,In_131);
and U2441 (N_2441,In_419,In_127);
nand U2442 (N_2442,In_667,In_331);
nand U2443 (N_2443,In_499,In_394);
nor U2444 (N_2444,In_159,In_268);
xor U2445 (N_2445,In_167,In_709);
or U2446 (N_2446,In_59,In_435);
nor U2447 (N_2447,In_519,In_598);
xnor U2448 (N_2448,In_186,In_110);
xnor U2449 (N_2449,In_54,In_458);
nand U2450 (N_2450,In_10,In_148);
nand U2451 (N_2451,In_541,In_172);
xor U2452 (N_2452,In_240,In_209);
nand U2453 (N_2453,In_9,In_109);
xnor U2454 (N_2454,In_661,In_684);
nand U2455 (N_2455,In_298,In_68);
and U2456 (N_2456,In_511,In_174);
or U2457 (N_2457,In_426,In_379);
nor U2458 (N_2458,In_156,In_294);
or U2459 (N_2459,In_614,In_453);
xnor U2460 (N_2460,In_164,In_328);
nor U2461 (N_2461,In_713,In_32);
nor U2462 (N_2462,In_696,In_600);
or U2463 (N_2463,In_497,In_441);
nand U2464 (N_2464,In_306,In_489);
and U2465 (N_2465,In_56,In_658);
nand U2466 (N_2466,In_335,In_43);
or U2467 (N_2467,In_604,In_526);
or U2468 (N_2468,In_41,In_327);
or U2469 (N_2469,In_634,In_445);
or U2470 (N_2470,In_495,In_621);
and U2471 (N_2471,In_717,In_606);
and U2472 (N_2472,In_365,In_511);
nand U2473 (N_2473,In_549,In_631);
and U2474 (N_2474,In_214,In_319);
or U2475 (N_2475,In_220,In_730);
nand U2476 (N_2476,In_28,In_81);
xor U2477 (N_2477,In_730,In_511);
and U2478 (N_2478,In_317,In_150);
or U2479 (N_2479,In_4,In_584);
nor U2480 (N_2480,In_308,In_624);
nand U2481 (N_2481,In_510,In_210);
nor U2482 (N_2482,In_262,In_374);
or U2483 (N_2483,In_408,In_38);
and U2484 (N_2484,In_395,In_303);
nor U2485 (N_2485,In_561,In_70);
xor U2486 (N_2486,In_669,In_270);
nand U2487 (N_2487,In_127,In_498);
nor U2488 (N_2488,In_226,In_505);
nand U2489 (N_2489,In_641,In_729);
xor U2490 (N_2490,In_432,In_331);
and U2491 (N_2491,In_109,In_434);
or U2492 (N_2492,In_615,In_22);
nand U2493 (N_2493,In_324,In_162);
nor U2494 (N_2494,In_518,In_288);
and U2495 (N_2495,In_483,In_410);
xor U2496 (N_2496,In_460,In_453);
or U2497 (N_2497,In_664,In_100);
nand U2498 (N_2498,In_237,In_507);
or U2499 (N_2499,In_586,In_112);
nor U2500 (N_2500,N_1181,N_191);
nor U2501 (N_2501,N_803,N_1722);
or U2502 (N_2502,N_473,N_659);
nor U2503 (N_2503,N_792,N_116);
and U2504 (N_2504,N_1785,N_1411);
or U2505 (N_2505,N_1644,N_912);
nand U2506 (N_2506,N_1145,N_1499);
and U2507 (N_2507,N_1897,N_1718);
nor U2508 (N_2508,N_1613,N_787);
or U2509 (N_2509,N_1929,N_513);
nand U2510 (N_2510,N_254,N_1941);
nand U2511 (N_2511,N_2119,N_570);
or U2512 (N_2512,N_2124,N_2228);
and U2513 (N_2513,N_1231,N_263);
or U2514 (N_2514,N_802,N_1899);
or U2515 (N_2515,N_1174,N_1825);
or U2516 (N_2516,N_1671,N_1434);
nand U2517 (N_2517,N_557,N_703);
or U2518 (N_2518,N_1924,N_2164);
and U2519 (N_2519,N_692,N_267);
nor U2520 (N_2520,N_1773,N_2410);
nand U2521 (N_2521,N_452,N_35);
nand U2522 (N_2522,N_598,N_610);
nand U2523 (N_2523,N_1221,N_2297);
nor U2524 (N_2524,N_704,N_2427);
and U2525 (N_2525,N_970,N_1707);
or U2526 (N_2526,N_1334,N_261);
or U2527 (N_2527,N_2203,N_418);
nor U2528 (N_2528,N_1206,N_1954);
nor U2529 (N_2529,N_638,N_1564);
and U2530 (N_2530,N_238,N_1703);
and U2531 (N_2531,N_743,N_2070);
nor U2532 (N_2532,N_2281,N_1368);
nand U2533 (N_2533,N_2393,N_662);
nor U2534 (N_2534,N_2007,N_1634);
nand U2535 (N_2535,N_1042,N_204);
or U2536 (N_2536,N_1255,N_1905);
nor U2537 (N_2537,N_1400,N_2457);
nor U2538 (N_2538,N_2463,N_1957);
nor U2539 (N_2539,N_274,N_290);
nand U2540 (N_2540,N_748,N_1316);
nand U2541 (N_2541,N_2091,N_251);
and U2542 (N_2542,N_1688,N_1521);
nor U2543 (N_2543,N_1534,N_1939);
and U2544 (N_2544,N_790,N_1951);
xnor U2545 (N_2545,N_1758,N_1120);
nor U2546 (N_2546,N_282,N_353);
nor U2547 (N_2547,N_2063,N_2148);
nor U2548 (N_2548,N_785,N_1458);
and U2549 (N_2549,N_2411,N_1178);
nand U2550 (N_2550,N_62,N_1639);
and U2551 (N_2551,N_1457,N_91);
nor U2552 (N_2552,N_306,N_928);
or U2553 (N_2553,N_1071,N_1708);
nand U2554 (N_2554,N_444,N_2183);
nor U2555 (N_2555,N_1354,N_1784);
or U2556 (N_2556,N_636,N_377);
nand U2557 (N_2557,N_2377,N_1973);
and U2558 (N_2558,N_1418,N_615);
and U2559 (N_2559,N_1234,N_917);
and U2560 (N_2560,N_75,N_1161);
or U2561 (N_2561,N_305,N_2420);
or U2562 (N_2562,N_966,N_442);
nor U2563 (N_2563,N_284,N_214);
xnor U2564 (N_2564,N_941,N_390);
nor U2565 (N_2565,N_2485,N_1168);
or U2566 (N_2566,N_97,N_666);
nor U2567 (N_2567,N_276,N_118);
nor U2568 (N_2568,N_721,N_2199);
or U2569 (N_2569,N_890,N_1753);
nand U2570 (N_2570,N_2376,N_985);
nor U2571 (N_2571,N_2288,N_430);
or U2572 (N_2572,N_1982,N_732);
nor U2573 (N_2573,N_1863,N_455);
nand U2574 (N_2574,N_2122,N_2469);
or U2575 (N_2575,N_893,N_1467);
or U2576 (N_2576,N_1369,N_222);
xnor U2577 (N_2577,N_438,N_1324);
nor U2578 (N_2578,N_70,N_1387);
or U2579 (N_2579,N_462,N_1682);
xor U2580 (N_2580,N_1648,N_411);
or U2581 (N_2581,N_1110,N_544);
and U2582 (N_2582,N_867,N_1995);
nand U2583 (N_2583,N_1967,N_2419);
nor U2584 (N_2584,N_1841,N_2165);
xnor U2585 (N_2585,N_1332,N_229);
nand U2586 (N_2586,N_246,N_1422);
nor U2587 (N_2587,N_609,N_1069);
or U2588 (N_2588,N_599,N_2035);
nor U2589 (N_2589,N_1143,N_577);
nand U2590 (N_2590,N_853,N_866);
or U2591 (N_2591,N_990,N_2027);
xnor U2592 (N_2592,N_82,N_2193);
nor U2593 (N_2593,N_1030,N_1625);
and U2594 (N_2594,N_877,N_142);
nand U2595 (N_2595,N_1050,N_2430);
nand U2596 (N_2596,N_1920,N_1796);
nor U2597 (N_2597,N_387,N_1646);
nand U2598 (N_2598,N_687,N_1937);
and U2599 (N_2599,N_769,N_2102);
nand U2600 (N_2600,N_2251,N_1686);
xnor U2601 (N_2601,N_889,N_818);
nor U2602 (N_2602,N_1872,N_1138);
xor U2603 (N_2603,N_73,N_407);
nor U2604 (N_2604,N_911,N_2213);
xnor U2605 (N_2605,N_2409,N_2138);
and U2606 (N_2606,N_838,N_2317);
and U2607 (N_2607,N_240,N_1609);
and U2608 (N_2608,N_1352,N_1163);
and U2609 (N_2609,N_2058,N_1478);
and U2610 (N_2610,N_1590,N_1011);
or U2611 (N_2611,N_695,N_1070);
nor U2612 (N_2612,N_1159,N_1019);
nor U2613 (N_2613,N_1105,N_1198);
nor U2614 (N_2614,N_232,N_1520);
or U2615 (N_2615,N_1531,N_1342);
and U2616 (N_2616,N_2338,N_1808);
and U2617 (N_2617,N_2214,N_194);
nand U2618 (N_2618,N_1051,N_1428);
and U2619 (N_2619,N_1752,N_2466);
or U2620 (N_2620,N_1782,N_1235);
nor U2621 (N_2621,N_804,N_129);
or U2622 (N_2622,N_78,N_1705);
and U2623 (N_2623,N_1474,N_1472);
nor U2624 (N_2624,N_2490,N_1371);
nand U2625 (N_2625,N_961,N_1853);
nor U2626 (N_2626,N_625,N_2118);
or U2627 (N_2627,N_2090,N_1035);
xnor U2628 (N_2628,N_1612,N_56);
and U2629 (N_2629,N_588,N_1603);
nor U2630 (N_2630,N_2342,N_2097);
nand U2631 (N_2631,N_134,N_1485);
nand U2632 (N_2632,N_656,N_2416);
nor U2633 (N_2633,N_1282,N_1783);
or U2634 (N_2634,N_1015,N_1965);
or U2635 (N_2635,N_117,N_712);
nor U2636 (N_2636,N_929,N_189);
nand U2637 (N_2637,N_664,N_1092);
nand U2638 (N_2638,N_2237,N_2182);
nor U2639 (N_2639,N_1495,N_1569);
nand U2640 (N_2640,N_1542,N_1621);
nor U2641 (N_2641,N_1618,N_356);
nor U2642 (N_2642,N_1194,N_2352);
or U2643 (N_2643,N_1366,N_2139);
or U2644 (N_2644,N_1777,N_2101);
or U2645 (N_2645,N_1873,N_1728);
nor U2646 (N_2646,N_809,N_706);
and U2647 (N_2647,N_650,N_46);
xnor U2648 (N_2648,N_1774,N_1806);
xnor U2649 (N_2649,N_1741,N_1242);
and U2650 (N_2650,N_2059,N_2045);
nand U2651 (N_2651,N_1433,N_566);
or U2652 (N_2652,N_1879,N_2057);
nand U2653 (N_2653,N_1341,N_1560);
xnor U2654 (N_2654,N_124,N_1479);
and U2655 (N_2655,N_1701,N_2405);
nor U2656 (N_2656,N_318,N_741);
xnor U2657 (N_2657,N_1126,N_1057);
or U2658 (N_2658,N_2181,N_11);
nor U2659 (N_2659,N_707,N_2191);
or U2660 (N_2660,N_474,N_791);
nor U2661 (N_2661,N_2412,N_206);
nand U2662 (N_2662,N_2019,N_1160);
or U2663 (N_2663,N_1635,N_1622);
or U2664 (N_2664,N_2304,N_1518);
nand U2665 (N_2665,N_2061,N_2459);
or U2666 (N_2666,N_1236,N_1606);
nor U2667 (N_2667,N_59,N_1153);
nor U2668 (N_2668,N_2255,N_17);
and U2669 (N_2669,N_1880,N_1944);
or U2670 (N_2670,N_775,N_1616);
and U2671 (N_2671,N_199,N_80);
and U2672 (N_2672,N_1575,N_1482);
or U2673 (N_2673,N_44,N_516);
xor U2674 (N_2674,N_810,N_1347);
nand U2675 (N_2675,N_1619,N_1127);
or U2676 (N_2676,N_1488,N_2468);
nand U2677 (N_2677,N_1059,N_1135);
nand U2678 (N_2678,N_312,N_2062);
nor U2679 (N_2679,N_1310,N_1481);
nor U2680 (N_2680,N_605,N_628);
and U2681 (N_2681,N_942,N_724);
nand U2682 (N_2682,N_1591,N_1241);
or U2683 (N_2683,N_1933,N_2290);
nand U2684 (N_2684,N_107,N_1441);
xnor U2685 (N_2685,N_383,N_937);
nand U2686 (N_2686,N_1854,N_1208);
nand U2687 (N_2687,N_244,N_1102);
and U2688 (N_2688,N_76,N_1810);
and U2689 (N_2689,N_1798,N_266);
nor U2690 (N_2690,N_1089,N_537);
or U2691 (N_2691,N_956,N_1516);
nor U2692 (N_2692,N_376,N_54);
nand U2693 (N_2693,N_1514,N_977);
and U2694 (N_2694,N_1245,N_2403);
xor U2695 (N_2695,N_1480,N_2074);
or U2696 (N_2696,N_705,N_1857);
and U2697 (N_2697,N_1771,N_906);
and U2698 (N_2698,N_1367,N_2355);
nand U2699 (N_2699,N_1763,N_2060);
xor U2700 (N_2700,N_1453,N_972);
or U2701 (N_2701,N_1142,N_1739);
xnor U2702 (N_2702,N_984,N_1445);
and U2703 (N_2703,N_1865,N_763);
nor U2704 (N_2704,N_137,N_1350);
nor U2705 (N_2705,N_2155,N_1577);
nand U2706 (N_2706,N_1169,N_1121);
nand U2707 (N_2707,N_1313,N_1526);
xnor U2708 (N_2708,N_34,N_1058);
nand U2709 (N_2709,N_2445,N_784);
nor U2710 (N_2710,N_1389,N_1195);
nor U2711 (N_2711,N_1617,N_1980);
and U2712 (N_2712,N_1451,N_24);
nand U2713 (N_2713,N_2323,N_1250);
nor U2714 (N_2714,N_2022,N_2429);
nor U2715 (N_2715,N_48,N_829);
or U2716 (N_2716,N_1395,N_963);
and U2717 (N_2717,N_1079,N_1755);
nor U2718 (N_2718,N_1704,N_1421);
nor U2719 (N_2719,N_2086,N_753);
nor U2720 (N_2720,N_427,N_1861);
or U2721 (N_2721,N_1695,N_2021);
nand U2722 (N_2722,N_641,N_2235);
nor U2723 (N_2723,N_2049,N_173);
nor U2724 (N_2724,N_2351,N_2006);
nand U2725 (N_2725,N_2220,N_378);
xor U2726 (N_2726,N_1775,N_945);
xor U2727 (N_2727,N_2284,N_1734);
nand U2728 (N_2728,N_611,N_1394);
and U2729 (N_2729,N_1826,N_2134);
or U2730 (N_2730,N_478,N_2083);
nor U2731 (N_2731,N_1111,N_1118);
nor U2732 (N_2732,N_2280,N_749);
nor U2733 (N_2733,N_1768,N_1925);
nor U2734 (N_2734,N_329,N_660);
and U2735 (N_2735,N_429,N_677);
nor U2736 (N_2736,N_2349,N_1620);
nor U2737 (N_2737,N_551,N_25);
xnor U2738 (N_2738,N_1788,N_690);
nand U2739 (N_2739,N_2225,N_2383);
and U2740 (N_2740,N_2115,N_903);
or U2741 (N_2741,N_169,N_668);
nand U2742 (N_2742,N_856,N_409);
and U2743 (N_2743,N_236,N_2363);
nor U2744 (N_2744,N_1333,N_1259);
xor U2745 (N_2745,N_1657,N_1228);
nor U2746 (N_2746,N_1288,N_1845);
or U2747 (N_2747,N_1296,N_88);
or U2748 (N_2748,N_164,N_591);
nand U2749 (N_2749,N_1476,N_110);
nor U2750 (N_2750,N_2464,N_152);
nand U2751 (N_2751,N_2286,N_1889);
and U2752 (N_2752,N_1253,N_2334);
nand U2753 (N_2753,N_899,N_959);
nor U2754 (N_2754,N_65,N_505);
nor U2755 (N_2755,N_1958,N_751);
nor U2756 (N_2756,N_823,N_256);
nor U2757 (N_2757,N_2067,N_1116);
and U2758 (N_2758,N_1427,N_279);
and U2759 (N_2759,N_1563,N_1263);
or U2760 (N_2760,N_2096,N_1468);
nand U2761 (N_2761,N_1824,N_686);
nand U2762 (N_2762,N_2396,N_141);
nor U2763 (N_2763,N_919,N_1884);
nand U2764 (N_2764,N_456,N_976);
nand U2765 (N_2765,N_1247,N_1483);
nor U2766 (N_2766,N_808,N_996);
and U2767 (N_2767,N_2448,N_488);
nand U2768 (N_2768,N_547,N_1869);
xnor U2769 (N_2769,N_1172,N_382);
nand U2770 (N_2770,N_1327,N_1054);
xor U2771 (N_2771,N_127,N_674);
xnor U2772 (N_2772,N_716,N_420);
nor U2773 (N_2773,N_559,N_2497);
or U2774 (N_2774,N_2229,N_616);
nand U2775 (N_2775,N_1960,N_1238);
or U2776 (N_2776,N_19,N_1171);
nand U2777 (N_2777,N_1740,N_1000);
or U2778 (N_2778,N_337,N_2394);
nor U2779 (N_2779,N_475,N_316);
nand U2780 (N_2780,N_2367,N_1456);
and U2781 (N_2781,N_1381,N_1589);
and U2782 (N_2782,N_1340,N_89);
and U2783 (N_2783,N_549,N_1436);
nand U2784 (N_2784,N_77,N_933);
xor U2785 (N_2785,N_2152,N_2343);
nor U2786 (N_2786,N_797,N_1535);
or U2787 (N_2787,N_1985,N_1556);
nand U2788 (N_2788,N_2492,N_1216);
nand U2789 (N_2789,N_2345,N_640);
or U2790 (N_2790,N_1203,N_723);
or U2791 (N_2791,N_375,N_79);
nor U2792 (N_2792,N_459,N_1404);
xnor U2793 (N_2793,N_2262,N_1225);
or U2794 (N_2794,N_2095,N_898);
and U2795 (N_2795,N_179,N_1399);
or U2796 (N_2796,N_449,N_1979);
and U2797 (N_2797,N_613,N_725);
nand U2798 (N_2798,N_1790,N_1412);
or U2799 (N_2799,N_1280,N_340);
and U2800 (N_2800,N_397,N_1338);
or U2801 (N_2801,N_2037,N_1878);
or U2802 (N_2802,N_271,N_2076);
or U2803 (N_2803,N_1191,N_2157);
nor U2804 (N_2804,N_1358,N_216);
or U2805 (N_2805,N_669,N_582);
or U2806 (N_2806,N_2285,N_2404);
xnor U2807 (N_2807,N_2054,N_1762);
nand U2808 (N_2808,N_243,N_61);
and U2809 (N_2809,N_2350,N_341);
nor U2810 (N_2810,N_103,N_421);
xnor U2811 (N_2811,N_500,N_2141);
nor U2812 (N_2812,N_1165,N_1385);
or U2813 (N_2813,N_1572,N_494);
or U2814 (N_2814,N_2269,N_857);
or U2815 (N_2815,N_1673,N_1156);
or U2816 (N_2816,N_1438,N_322);
or U2817 (N_2817,N_342,N_339);
nor U2818 (N_2818,N_1176,N_175);
and U2819 (N_2819,N_2175,N_231);
and U2820 (N_2820,N_900,N_1917);
nor U2821 (N_2821,N_998,N_2145);
nand U2822 (N_2822,N_396,N_359);
and U2823 (N_2823,N_2346,N_190);
xnor U2824 (N_2824,N_1681,N_1510);
nand U2825 (N_2825,N_1281,N_534);
or U2826 (N_2826,N_973,N_737);
nor U2827 (N_2827,N_532,N_1570);
and U2828 (N_2828,N_1230,N_181);
and U2829 (N_2829,N_1527,N_1866);
and U2830 (N_2830,N_675,N_1950);
nand U2831 (N_2831,N_1239,N_1098);
nand U2832 (N_2832,N_257,N_1522);
and U2833 (N_2833,N_2208,N_1328);
nand U2834 (N_2834,N_2489,N_719);
or U2835 (N_2835,N_83,N_527);
and U2836 (N_2836,N_1345,N_1723);
or U2837 (N_2837,N_962,N_672);
nor U2838 (N_2838,N_2261,N_1013);
or U2839 (N_2839,N_311,N_2369);
and U2840 (N_2840,N_1099,N_2008);
or U2841 (N_2841,N_2081,N_1470);
nand U2842 (N_2842,N_1061,N_1945);
nand U2843 (N_2843,N_149,N_589);
nor U2844 (N_2844,N_1698,N_1066);
nor U2845 (N_2845,N_2186,N_289);
and U2846 (N_2846,N_1858,N_386);
nor U2847 (N_2847,N_1193,N_2392);
nand U2848 (N_2848,N_1760,N_57);
nand U2849 (N_2849,N_496,N_1076);
nand U2850 (N_2850,N_224,N_634);
or U2851 (N_2851,N_1379,N_1048);
or U2852 (N_2852,N_1595,N_183);
xor U2853 (N_2853,N_2472,N_2458);
nor U2854 (N_2854,N_2402,N_2263);
xor U2855 (N_2855,N_151,N_2250);
and U2856 (N_2856,N_1182,N_1601);
nor U2857 (N_2857,N_2426,N_2205);
or U2858 (N_2858,N_2105,N_1793);
or U2859 (N_2859,N_1525,N_2123);
xnor U2860 (N_2860,N_1439,N_1977);
nor U2861 (N_2861,N_1638,N_177);
nand U2862 (N_2862,N_303,N_1930);
nand U2863 (N_2863,N_1666,N_1357);
nand U2864 (N_2864,N_2391,N_1506);
nand U2865 (N_2865,N_673,N_852);
and U2866 (N_2866,N_1931,N_2116);
or U2867 (N_2867,N_925,N_2480);
nand U2868 (N_2868,N_835,N_255);
or U2869 (N_2869,N_1665,N_1084);
nand U2870 (N_2870,N_1713,N_2310);
nor U2871 (N_2871,N_132,N_1383);
nand U2872 (N_2872,N_1746,N_1712);
nor U2873 (N_2873,N_2434,N_780);
nand U2874 (N_2874,N_680,N_36);
nand U2875 (N_2875,N_2011,N_623);
nor U2876 (N_2876,N_1815,N_49);
and U2877 (N_2877,N_1576,N_26);
and U2878 (N_2878,N_1492,N_1106);
and U2879 (N_2879,N_1139,N_272);
xnor U2880 (N_2880,N_125,N_230);
xnor U2881 (N_2881,N_1124,N_606);
or U2882 (N_2882,N_2357,N_2162);
nand U2883 (N_2883,N_1305,N_2340);
or U2884 (N_2884,N_874,N_400);
and U2885 (N_2885,N_55,N_1487);
or U2886 (N_2886,N_1087,N_1370);
nor U2887 (N_2887,N_902,N_1093);
or U2888 (N_2888,N_463,N_2364);
nor U2889 (N_2889,N_1088,N_2386);
or U2890 (N_2890,N_72,N_1033);
and U2891 (N_2891,N_93,N_2380);
nand U2892 (N_2892,N_2299,N_847);
and U2893 (N_2893,N_60,N_2337);
nand U2894 (N_2894,N_543,N_99);
nor U2895 (N_2895,N_495,N_458);
or U2896 (N_2896,N_321,N_1262);
and U2897 (N_2897,N_1107,N_1002);
and U2898 (N_2898,N_720,N_1805);
and U2899 (N_2899,N_381,N_31);
nor U2900 (N_2900,N_1991,N_112);
or U2901 (N_2901,N_975,N_1025);
nor U2902 (N_2902,N_1565,N_1814);
xnor U2903 (N_2903,N_860,N_319);
nand U2904 (N_2904,N_2414,N_1849);
nand U2905 (N_2905,N_286,N_1373);
and U2906 (N_2906,N_1538,N_66);
nand U2907 (N_2907,N_1044,N_176);
and U2908 (N_2908,N_101,N_374);
or U2909 (N_2909,N_71,N_1992);
nand U2910 (N_2910,N_2065,N_2483);
nor U2911 (N_2911,N_536,N_540);
and U2912 (N_2912,N_627,N_1598);
and U2913 (N_2913,N_21,N_1730);
and U2914 (N_2914,N_1402,N_2204);
nor U2915 (N_2915,N_363,N_2108);
or U2916 (N_2916,N_868,N_1668);
xnor U2917 (N_2917,N_1726,N_38);
and U2918 (N_2918,N_888,N_2189);
and U2919 (N_2919,N_924,N_197);
nor U2920 (N_2920,N_2137,N_670);
nor U2921 (N_2921,N_521,N_327);
and U2922 (N_2922,N_2014,N_1505);
or U2923 (N_2923,N_1710,N_742);
and U2924 (N_2924,N_1844,N_1818);
or U2925 (N_2925,N_2314,N_1949);
and U2926 (N_2926,N_750,N_200);
nand U2927 (N_2927,N_1154,N_1401);
nor U2928 (N_2928,N_172,N_1993);
nor U2929 (N_2929,N_1656,N_1765);
nand U2930 (N_2930,N_1137,N_1706);
nor U2931 (N_2931,N_1677,N_815);
nand U2932 (N_2932,N_1988,N_824);
xnor U2933 (N_2933,N_1754,N_793);
nor U2934 (N_2934,N_2303,N_1691);
nand U2935 (N_2935,N_1173,N_2477);
xnor U2936 (N_2936,N_2153,N_1817);
and U2937 (N_2937,N_762,N_1109);
and U2938 (N_2938,N_2400,N_113);
xnor U2939 (N_2939,N_930,N_2217);
nand U2940 (N_2940,N_980,N_2293);
nor U2941 (N_2941,N_1278,N_947);
or U2942 (N_2942,N_2234,N_2329);
and U2943 (N_2943,N_502,N_2399);
nand U2944 (N_2944,N_1183,N_1942);
xor U2945 (N_2945,N_2029,N_1297);
nor U2946 (N_2946,N_424,N_1749);
nand U2947 (N_2947,N_512,N_1122);
or U2948 (N_2948,N_1643,N_2318);
or U2949 (N_2949,N_2036,N_2253);
or U2950 (N_2950,N_145,N_1588);
and U2951 (N_2951,N_2238,N_1264);
and U2952 (N_2952,N_504,N_395);
nand U2953 (N_2953,N_317,N_1318);
nor U2954 (N_2954,N_1291,N_1331);
and U2955 (N_2955,N_1348,N_2302);
or U2956 (N_2956,N_294,N_287);
or U2957 (N_2957,N_2406,N_1764);
or U2958 (N_2958,N_135,N_1852);
nand U2959 (N_2959,N_58,N_1396);
xnor U2960 (N_2960,N_2192,N_1955);
and U2961 (N_2961,N_548,N_2471);
nand U2962 (N_2962,N_935,N_603);
nor U2963 (N_2963,N_349,N_439);
or U2964 (N_2964,N_2000,N_842);
nand U2965 (N_2965,N_85,N_195);
or U2966 (N_2966,N_2106,N_92);
nor U2967 (N_2967,N_2136,N_2498);
nand U2968 (N_2968,N_414,N_1587);
nor U2969 (N_2969,N_2247,N_635);
or U2970 (N_2970,N_1851,N_2442);
or U2971 (N_2971,N_1675,N_1398);
nand U2972 (N_2972,N_1811,N_350);
nor U2973 (N_2973,N_1876,N_1792);
and U2974 (N_2974,N_1660,N_1607);
and U2975 (N_2975,N_192,N_2366);
and U2976 (N_2976,N_466,N_1406);
xnor U2977 (N_2977,N_830,N_208);
nor U2978 (N_2978,N_367,N_1883);
xnor U2979 (N_2979,N_69,N_2439);
or U2980 (N_2980,N_1286,N_1983);
nor U2981 (N_2981,N_2018,N_211);
nand U2982 (N_2982,N_1166,N_2093);
nor U2983 (N_2983,N_530,N_2195);
xnor U2984 (N_2984,N_2215,N_302);
and U2985 (N_2985,N_1224,N_2407);
nand U2986 (N_2986,N_604,N_944);
and U2987 (N_2987,N_710,N_837);
and U2988 (N_2988,N_174,N_1874);
or U2989 (N_2989,N_1254,N_3);
and U2990 (N_2990,N_1486,N_1081);
nor U2991 (N_2991,N_2425,N_1839);
or U2992 (N_2992,N_1028,N_2158);
or U2993 (N_2993,N_2210,N_2179);
nor U2994 (N_2994,N_1658,N_795);
and U2995 (N_2995,N_1921,N_826);
nand U2996 (N_2996,N_533,N_1994);
nor U2997 (N_2997,N_1295,N_334);
nor U2998 (N_2998,N_1032,N_1149);
or U2999 (N_2999,N_1838,N_564);
xnor U3000 (N_3000,N_827,N_736);
nand U3001 (N_3001,N_2089,N_1714);
nor U3002 (N_3002,N_1232,N_45);
nor U3003 (N_3003,N_460,N_170);
nor U3004 (N_3004,N_691,N_2099);
and U3005 (N_3005,N_850,N_1902);
nor U3006 (N_3006,N_596,N_832);
nand U3007 (N_3007,N_1888,N_1094);
nor U3008 (N_3008,N_1012,N_683);
and U3009 (N_3009,N_590,N_1336);
nand U3010 (N_3010,N_1157,N_1539);
or U3011 (N_3011,N_2015,N_1319);
and U3012 (N_3012,N_1747,N_592);
and U3013 (N_3013,N_831,N_1192);
or U3014 (N_3014,N_1375,N_1493);
or U3015 (N_3015,N_1963,N_1240);
xnor U3016 (N_3016,N_2112,N_1503);
nand U3017 (N_3017,N_1339,N_1557);
nor U3018 (N_3018,N_965,N_1045);
nand U3019 (N_3019,N_1210,N_1130);
nand U3020 (N_3020,N_1894,N_1407);
nor U3021 (N_3021,N_209,N_2233);
or U3022 (N_3022,N_1132,N_729);
nand U3023 (N_3023,N_468,N_128);
nor U3024 (N_3024,N_187,N_820);
nor U3025 (N_3025,N_2388,N_587);
and U3026 (N_3026,N_997,N_1721);
nor U3027 (N_3027,N_1355,N_484);
and U3028 (N_3028,N_1885,N_1699);
nor U3029 (N_3029,N_1346,N_479);
nor U3030 (N_3030,N_2040,N_2339);
or U3031 (N_3031,N_2451,N_520);
xor U3032 (N_3032,N_1948,N_7);
and U3033 (N_3033,N_196,N_2474);
and U3034 (N_3034,N_817,N_1276);
and U3035 (N_3035,N_584,N_1700);
nand U3036 (N_3036,N_968,N_1578);
and U3037 (N_3037,N_2249,N_1757);
nand U3038 (N_3038,N_2431,N_2360);
or U3039 (N_3039,N_2232,N_940);
or U3040 (N_3040,N_1414,N_2421);
and U3041 (N_3041,N_1997,N_2413);
nand U3042 (N_3042,N_630,N_896);
nand U3043 (N_3043,N_806,N_2449);
or U3044 (N_3044,N_1926,N_2025);
nand U3045 (N_3045,N_226,N_1964);
nor U3046 (N_3046,N_1215,N_2159);
and U3047 (N_3047,N_1261,N_1080);
and U3048 (N_3048,N_617,N_2375);
and U3049 (N_3049,N_40,N_1243);
xnor U3050 (N_3050,N_165,N_2331);
xnor U3051 (N_3051,N_1791,N_845);
nand U3052 (N_3052,N_120,N_878);
and U3053 (N_3053,N_2194,N_2163);
xnor U3054 (N_3054,N_718,N_1962);
or U3055 (N_3055,N_1830,N_1196);
nand U3056 (N_3056,N_1068,N_1162);
nor U3057 (N_3057,N_535,N_50);
or U3058 (N_3058,N_764,N_307);
nand U3059 (N_3059,N_18,N_435);
nand U3060 (N_3060,N_1461,N_354);
nor U3061 (N_3061,N_2166,N_529);
nor U3062 (N_3062,N_987,N_1614);
or U3063 (N_3063,N_239,N_469);
or U3064 (N_3064,N_1725,N_2488);
and U3065 (N_3065,N_2142,N_1680);
nor U3066 (N_3066,N_1463,N_949);
or U3067 (N_3067,N_2440,N_1789);
nor U3068 (N_3068,N_2294,N_2026);
and U3069 (N_3069,N_1413,N_955);
nand U3070 (N_3070,N_665,N_884);
and U3071 (N_3071,N_1256,N_2456);
and U3072 (N_3072,N_2344,N_1390);
nand U3073 (N_3073,N_782,N_918);
nor U3074 (N_3074,N_733,N_854);
or U3075 (N_3075,N_967,N_1786);
and U3076 (N_3076,N_1836,N_1226);
and U3077 (N_3077,N_227,N_182);
nor U3078 (N_3078,N_2265,N_140);
nand U3079 (N_3079,N_1175,N_1023);
nor U3080 (N_3080,N_497,N_265);
nand U3081 (N_3081,N_1056,N_2087);
and U3082 (N_3082,N_1750,N_2185);
or U3083 (N_3083,N_562,N_506);
and U3084 (N_3084,N_1213,N_1821);
xor U3085 (N_3085,N_556,N_567);
nand U3086 (N_3086,N_1662,N_1447);
or U3087 (N_3087,N_417,N_81);
nor U3088 (N_3088,N_1329,N_1751);
or U3089 (N_3089,N_2252,N_1694);
nand U3090 (N_3090,N_1446,N_1464);
and U3091 (N_3091,N_1914,N_682);
nor U3092 (N_3092,N_1197,N_1915);
or U3093 (N_3093,N_499,N_1626);
or U3094 (N_3094,N_361,N_581);
or U3095 (N_3095,N_2268,N_799);
nor U3096 (N_3096,N_573,N_297);
nor U3097 (N_3097,N_2438,N_1146);
and U3098 (N_3098,N_859,N_657);
nand U3099 (N_3099,N_624,N_801);
nor U3100 (N_3100,N_32,N_268);
or U3101 (N_3101,N_2336,N_347);
nand U3102 (N_3102,N_583,N_600);
nor U3103 (N_3103,N_1448,N_1437);
xor U3104 (N_3104,N_767,N_1970);
nor U3105 (N_3105,N_2196,N_2169);
or U3106 (N_3106,N_482,N_2499);
xnor U3107 (N_3107,N_1010,N_1907);
nand U3108 (N_3108,N_2371,N_1641);
nor U3109 (N_3109,N_150,N_2446);
nand U3110 (N_3110,N_2177,N_1776);
nor U3111 (N_3111,N_816,N_1544);
or U3112 (N_3112,N_1005,N_1756);
and U3113 (N_3113,N_1365,N_905);
and U3114 (N_3114,N_957,N_1582);
and U3115 (N_3115,N_1833,N_1189);
nand U3116 (N_3116,N_813,N_1214);
and U3117 (N_3117,N_1523,N_1610);
or U3118 (N_3118,N_1152,N_631);
nor U3119 (N_3119,N_493,N_2151);
xor U3120 (N_3120,N_1496,N_2452);
nor U3121 (N_3121,N_2170,N_2223);
and U3122 (N_3122,N_1709,N_445);
nand U3123 (N_3123,N_1440,N_1207);
nor U3124 (N_3124,N_639,N_1301);
and U3125 (N_3125,N_1500,N_578);
and U3126 (N_3126,N_1947,N_291);
xor U3127 (N_3127,N_486,N_1652);
nand U3128 (N_3128,N_542,N_186);
nor U3129 (N_3129,N_1684,N_2031);
and U3130 (N_3130,N_221,N_722);
nand U3131 (N_3131,N_403,N_2052);
and U3132 (N_3132,N_1104,N_734);
and U3133 (N_3133,N_999,N_2023);
or U3134 (N_3134,N_2126,N_1968);
xnor U3135 (N_3135,N_2272,N_676);
and U3136 (N_3136,N_786,N_1584);
nor U3137 (N_3137,N_419,N_2129);
nand U3138 (N_3138,N_2212,N_392);
nand U3139 (N_3139,N_633,N_2259);
nand U3140 (N_3140,N_343,N_20);
nor U3141 (N_3141,N_910,N_1583);
nor U3142 (N_3142,N_2361,N_1976);
nand U3143 (N_3143,N_1063,N_858);
nor U3144 (N_3144,N_745,N_2432);
or U3145 (N_3145,N_2094,N_1119);
or U3146 (N_3146,N_1653,N_447);
or U3147 (N_3147,N_948,N_1562);
or U3148 (N_3148,N_621,N_517);
or U3149 (N_3149,N_1549,N_2);
nor U3150 (N_3150,N_154,N_2222);
and U3151 (N_3151,N_776,N_2465);
or U3152 (N_3152,N_1167,N_552);
nand U3153 (N_3153,N_1819,N_1031);
or U3154 (N_3154,N_1409,N_344);
nand U3155 (N_3155,N_932,N_41);
or U3156 (N_3156,N_1891,N_388);
nand U3157 (N_3157,N_1835,N_2254);
and U3158 (N_3158,N_836,N_1551);
nor U3159 (N_3159,N_52,N_1566);
nand U3160 (N_3160,N_1302,N_2327);
nand U3161 (N_3161,N_663,N_538);
nand U3162 (N_3162,N_1140,N_2278);
or U3163 (N_3163,N_2493,N_415);
nor U3164 (N_3164,N_514,N_1211);
or U3165 (N_3165,N_1855,N_39);
and U3166 (N_3166,N_871,N_1667);
and U3167 (N_3167,N_365,N_369);
and U3168 (N_3168,N_2467,N_1637);
and U3169 (N_3169,N_649,N_1277);
and U3170 (N_3170,N_247,N_1972);
nand U3171 (N_3171,N_2197,N_53);
or U3172 (N_3172,N_1016,N_2012);
nand U3173 (N_3173,N_1384,N_2312);
and U3174 (N_3174,N_1290,N_1910);
or U3175 (N_3175,N_1927,N_1125);
and U3176 (N_3176,N_1220,N_2024);
nand U3177 (N_3177,N_1155,N_2418);
or U3178 (N_3178,N_2374,N_760);
and U3179 (N_3179,N_2154,N_410);
nand U3180 (N_3180,N_467,N_425);
or U3181 (N_3181,N_1133,N_2168);
xnor U3182 (N_3182,N_2047,N_658);
xnor U3183 (N_3183,N_1454,N_2082);
nand U3184 (N_3184,N_144,N_422);
nor U3185 (N_3185,N_1881,N_1943);
and U3186 (N_3186,N_260,N_1374);
nor U3187 (N_3187,N_2130,N_1738);
or U3188 (N_3188,N_2075,N_1596);
nor U3189 (N_3189,N_2032,N_1744);
nor U3190 (N_3190,N_1892,N_2071);
nand U3191 (N_3191,N_223,N_2020);
and U3192 (N_3192,N_1901,N_215);
nand U3193 (N_3193,N_1420,N_485);
or U3194 (N_3194,N_2201,N_880);
nand U3195 (N_3195,N_1761,N_708);
or U3196 (N_3196,N_2347,N_193);
and U3197 (N_3197,N_1903,N_844);
or U3198 (N_3198,N_1898,N_1693);
and U3199 (N_3199,N_1990,N_1640);
xor U3200 (N_3200,N_1018,N_218);
or U3201 (N_3201,N_654,N_1008);
or U3202 (N_3202,N_1027,N_28);
nor U3203 (N_3203,N_2227,N_233);
nand U3204 (N_3204,N_471,N_296);
and U3205 (N_3205,N_357,N_2013);
or U3206 (N_3206,N_1376,N_1101);
nor U3207 (N_3207,N_2378,N_1403);
or U3208 (N_3208,N_2478,N_2275);
nor U3209 (N_3209,N_1987,N_1364);
or U3210 (N_3210,N_2044,N_1683);
nand U3211 (N_3211,N_558,N_432);
nand U3212 (N_3212,N_1223,N_2160);
and U3213 (N_3213,N_1410,N_1559);
nand U3214 (N_3214,N_755,N_1219);
and U3215 (N_3215,N_1909,N_1735);
and U3216 (N_3216,N_772,N_153);
nand U3217 (N_3217,N_108,N_259);
nand U3218 (N_3218,N_1200,N_15);
nor U3219 (N_3219,N_2239,N_2309);
nor U3220 (N_3220,N_273,N_1465);
and U3221 (N_3221,N_2273,N_2033);
nand U3222 (N_3222,N_1047,N_974);
xor U3223 (N_3223,N_696,N_981);
nand U3224 (N_3224,N_237,N_373);
and U3225 (N_3225,N_825,N_1359);
and U3226 (N_3226,N_51,N_406);
nor U3227 (N_3227,N_1906,N_2300);
nor U3228 (N_3228,N_907,N_2370);
nor U3229 (N_3229,N_1307,N_2002);
nor U3230 (N_3230,N_2080,N_1627);
nand U3231 (N_3231,N_926,N_872);
nor U3232 (N_3232,N_2368,N_234);
nand U3233 (N_3233,N_1314,N_2190);
or U3234 (N_3234,N_1444,N_1335);
nor U3235 (N_3235,N_642,N_2333);
nor U3236 (N_3236,N_938,N_300);
or U3237 (N_3237,N_920,N_384);
or U3238 (N_3238,N_2077,N_205);
and U3239 (N_3239,N_1248,N_756);
nor U3240 (N_3240,N_1308,N_1021);
nor U3241 (N_3241,N_245,N_331);
nand U3242 (N_3242,N_2295,N_1585);
nor U3243 (N_3243,N_579,N_2365);
and U3244 (N_3244,N_1647,N_1843);
nand U3245 (N_3245,N_1797,N_2306);
and U3246 (N_3246,N_2324,N_2171);
or U3247 (N_3247,N_1727,N_1325);
and U3248 (N_3248,N_269,N_1600);
nand U3249 (N_3249,N_1416,N_1813);
and U3250 (N_3250,N_1770,N_412);
or U3251 (N_3251,N_332,N_2260);
and U3252 (N_3252,N_1004,N_133);
nand U3253 (N_3253,N_2384,N_519);
nor U3254 (N_3254,N_2009,N_1184);
or U3255 (N_3255,N_895,N_960);
and U3256 (N_3256,N_483,N_1131);
and U3257 (N_3257,N_1524,N_2140);
and U3258 (N_3258,N_1809,N_1599);
or U3259 (N_3259,N_2453,N_1630);
or U3260 (N_3260,N_620,N_2476);
and U3261 (N_3261,N_1594,N_180);
xnor U3262 (N_3262,N_295,N_1604);
and U3263 (N_3263,N_1123,N_426);
and U3264 (N_3264,N_1636,N_1502);
xnor U3265 (N_3265,N_702,N_235);
and U3266 (N_3266,N_1073,N_1337);
nor U3267 (N_3267,N_653,N_29);
and U3268 (N_3268,N_1919,N_2051);
nor U3269 (N_3269,N_2200,N_1459);
nand U3270 (N_3270,N_1148,N_1309);
nand U3271 (N_3271,N_523,N_913);
nor U3272 (N_3272,N_2325,N_1266);
nand U3273 (N_3273,N_646,N_428);
or U3274 (N_3274,N_2241,N_1246);
or U3275 (N_3275,N_2207,N_1517);
and U3276 (N_3276,N_979,N_1780);
xnor U3277 (N_3277,N_921,N_2161);
or U3278 (N_3278,N_1936,N_851);
nor U3279 (N_3279,N_954,N_727);
and U3280 (N_3280,N_927,N_385);
nor U3281 (N_3281,N_526,N_309);
and U3282 (N_3282,N_5,N_711);
nand U3283 (N_3283,N_2172,N_1904);
or U3284 (N_3284,N_794,N_522);
nand U3285 (N_3285,N_971,N_220);
nand U3286 (N_3286,N_1151,N_1868);
and U3287 (N_3287,N_2379,N_1651);
nand U3288 (N_3288,N_671,N_1581);
nor U3289 (N_3289,N_2354,N_699);
and U3290 (N_3290,N_453,N_1179);
and U3291 (N_3291,N_614,N_413);
or U3292 (N_3292,N_1060,N_796);
and U3293 (N_3293,N_2358,N_1017);
nor U3294 (N_3294,N_2455,N_2428);
and U3295 (N_3295,N_207,N_1432);
nand U3296 (N_3296,N_1431,N_576);
nand U3297 (N_3297,N_2231,N_2276);
nor U3298 (N_3298,N_580,N_2372);
nor U3299 (N_3299,N_1077,N_1455);
nand U3300 (N_3300,N_2030,N_441);
nand U3301 (N_3301,N_1989,N_1190);
nor U3302 (N_3302,N_1961,N_839);
or U3303 (N_3303,N_1923,N_1001);
nor U3304 (N_3304,N_90,N_768);
nor U3305 (N_3305,N_923,N_1848);
nand U3306 (N_3306,N_1846,N_2330);
nor U3307 (N_3307,N_398,N_2264);
nand U3308 (N_3308,N_511,N_561);
nand U3309 (N_3309,N_1512,N_402);
xor U3310 (N_3310,N_2266,N_2311);
nor U3311 (N_3311,N_121,N_1096);
and U3312 (N_3312,N_1078,N_30);
or U3313 (N_3313,N_253,N_1847);
nor U3314 (N_3314,N_1022,N_2156);
xor U3315 (N_3315,N_1912,N_84);
and U3316 (N_3316,N_2257,N_2443);
nor U3317 (N_3317,N_104,N_346);
nor U3318 (N_3318,N_210,N_1289);
nor U3319 (N_3319,N_1180,N_1561);
xor U3320 (N_3320,N_1733,N_994);
or U3321 (N_3321,N_1343,N_679);
or U3322 (N_3322,N_1330,N_1471);
nor U3323 (N_3323,N_156,N_2450);
xor U3324 (N_3324,N_1946,N_1592);
nor U3325 (N_3325,N_454,N_162);
nor U3326 (N_3326,N_380,N_2398);
nand U3327 (N_3327,N_1676,N_1405);
nand U3328 (N_3328,N_2046,N_1469);
or U3329 (N_3329,N_1271,N_2321);
xor U3330 (N_3330,N_571,N_1530);
nor U3331 (N_3331,N_1998,N_171);
and U3332 (N_3332,N_607,N_1632);
nand U3333 (N_3333,N_1204,N_1423);
xor U3334 (N_3334,N_1270,N_1711);
and U3335 (N_3335,N_541,N_16);
or U3336 (N_3336,N_472,N_1745);
xor U3337 (N_3337,N_612,N_43);
and U3338 (N_3338,N_2435,N_23);
nand U3339 (N_3339,N_371,N_320);
xor U3340 (N_3340,N_1186,N_1349);
or U3341 (N_3341,N_1966,N_1862);
nor U3342 (N_3342,N_841,N_1091);
and U3343 (N_3343,N_1064,N_1362);
or U3344 (N_3344,N_2073,N_883);
nand U3345 (N_3345,N_887,N_1547);
and U3346 (N_3346,N_4,N_811);
nor U3347 (N_3347,N_1678,N_2017);
nand U3348 (N_3348,N_1928,N_2113);
and U3349 (N_3349,N_490,N_1498);
or U3350 (N_3350,N_1046,N_389);
and U3351 (N_3351,N_694,N_2326);
nor U3352 (N_3352,N_1822,N_2041);
nor U3353 (N_3353,N_372,N_159);
nor U3354 (N_3354,N_1940,N_539);
or U3355 (N_3355,N_1724,N_876);
xor U3356 (N_3356,N_1075,N_555);
and U3357 (N_3357,N_969,N_689);
nand U3358 (N_3358,N_299,N_2167);
or U3359 (N_3359,N_593,N_434);
or U3360 (N_3360,N_1424,N_840);
nor U3361 (N_3361,N_1743,N_833);
nor U3362 (N_3362,N_1719,N_1567);
nand U3363 (N_3363,N_416,N_746);
nor U3364 (N_3364,N_446,N_1085);
or U3365 (N_3365,N_2230,N_2390);
nor U3366 (N_3366,N_1426,N_470);
and U3367 (N_3367,N_277,N_2287);
nand U3368 (N_3368,N_2462,N_862);
nor U3369 (N_3369,N_394,N_217);
nand U3370 (N_3370,N_717,N_2245);
and U3371 (N_3371,N_405,N_643);
or U3372 (N_3372,N_1654,N_915);
and U3373 (N_3373,N_1697,N_2437);
nand U3374 (N_3374,N_2144,N_2359);
and U3375 (N_3375,N_2098,N_629);
nand U3376 (N_3376,N_1217,N_2258);
nor U3377 (N_3377,N_1537,N_752);
or U3378 (N_3378,N_1491,N_1269);
nor U3379 (N_3379,N_1759,N_1134);
nand U3380 (N_3380,N_292,N_2319);
nand U3381 (N_3381,N_778,N_126);
or U3382 (N_3382,N_1602,N_518);
or U3383 (N_3383,N_492,N_2289);
or U3384 (N_3384,N_1890,N_1952);
or U3385 (N_3385,N_2486,N_2461);
and U3386 (N_3386,N_27,N_451);
nor U3387 (N_3387,N_515,N_939);
or U3388 (N_3388,N_2292,N_568);
or U3389 (N_3389,N_1177,N_1669);
xor U3390 (N_3390,N_201,N_1322);
and U3391 (N_3391,N_1272,N_1860);
or U3392 (N_3392,N_1209,N_1429);
nor U3393 (N_3393,N_166,N_1974);
or U3394 (N_3394,N_2496,N_684);
nor U3395 (N_3395,N_619,N_651);
nor U3396 (N_3396,N_203,N_2072);
and U3397 (N_3397,N_988,N_546);
nor U3398 (N_3398,N_1642,N_111);
xor U3399 (N_3399,N_715,N_1244);
nor U3400 (N_3400,N_1742,N_2382);
and U3401 (N_3401,N_1185,N_298);
xnor U3402 (N_3402,N_1515,N_1956);
nand U3403 (N_3403,N_2050,N_507);
nor U3404 (N_3404,N_1435,N_1150);
xor U3405 (N_3405,N_2110,N_1674);
nand U3406 (N_3406,N_1144,N_1300);
or U3407 (N_3407,N_1624,N_1494);
nor U3408 (N_3408,N_2085,N_185);
and U3409 (N_3409,N_1893,N_821);
nor U3410 (N_3410,N_94,N_2315);
or U3411 (N_3411,N_1812,N_1392);
xor U3412 (N_3412,N_1114,N_457);
nand U3413 (N_3413,N_1552,N_1415);
and U3414 (N_3414,N_524,N_248);
xor U3415 (N_3415,N_602,N_358);
nor U3416 (N_3416,N_2221,N_1475);
and U3417 (N_3417,N_2242,N_1233);
and U3418 (N_3418,N_399,N_1315);
or U3419 (N_3419,N_1450,N_1938);
or U3420 (N_3420,N_891,N_115);
nor U3421 (N_3421,N_1953,N_1593);
and U3422 (N_3422,N_1283,N_744);
nor U3423 (N_3423,N_1827,N_2240);
nand U3424 (N_3424,N_1679,N_2274);
nor U3425 (N_3425,N_693,N_487);
or U3426 (N_3426,N_1801,N_1009);
xor U3427 (N_3427,N_68,N_618);
or U3428 (N_3428,N_1586,N_423);
or U3429 (N_3429,N_1,N_433);
nand U3430 (N_3430,N_2066,N_1212);
and U3431 (N_3431,N_0,N_2373);
and U3432 (N_3432,N_1922,N_8);
nor U3433 (N_3433,N_6,N_2109);
nand U3434 (N_3434,N_1380,N_105);
nor U3435 (N_3435,N_1504,N_528);
and U3436 (N_3436,N_1840,N_1864);
xnor U3437 (N_3437,N_2188,N_601);
xor U3438 (N_3438,N_774,N_740);
and U3439 (N_3439,N_393,N_739);
and U3440 (N_3440,N_437,N_1649);
or U3441 (N_3441,N_914,N_700);
xor U3442 (N_3442,N_13,N_301);
nor U3443 (N_3443,N_1293,N_1579);
or U3444 (N_3444,N_1026,N_983);
or U3445 (N_3445,N_2103,N_2004);
nand U3446 (N_3446,N_477,N_1611);
or U3447 (N_3447,N_123,N_1103);
and U3448 (N_3448,N_1716,N_1580);
and U3449 (N_3449,N_1170,N_160);
and U3450 (N_3450,N_2068,N_213);
and U3451 (N_3451,N_1696,N_882);
nor U3452 (N_3452,N_798,N_1935);
and U3453 (N_3453,N_2436,N_310);
nor U3454 (N_3454,N_678,N_1100);
and U3455 (N_3455,N_1918,N_95);
nand U3456 (N_3456,N_1408,N_324);
nor U3457 (N_3457,N_819,N_1911);
nor U3458 (N_3458,N_96,N_1528);
xnor U3459 (N_3459,N_800,N_2353);
or U3460 (N_3460,N_184,N_2042);
nor U3461 (N_3461,N_167,N_1320);
or U3462 (N_3462,N_1779,N_37);
nand U3463 (N_3463,N_1490,N_1275);
xor U3464 (N_3464,N_2127,N_1690);
or U3465 (N_3465,N_783,N_1043);
nor U3466 (N_3466,N_1882,N_391);
or U3467 (N_3467,N_1687,N_87);
and U3468 (N_3468,N_102,N_1615);
and U3469 (N_3469,N_1548,N_9);
and U3470 (N_3470,N_2056,N_2131);
nor U3471 (N_3471,N_1908,N_1298);
nand U3472 (N_3472,N_461,N_1268);
nand U3473 (N_3473,N_2187,N_1052);
or U3474 (N_3474,N_2494,N_2005);
nor U3475 (N_3475,N_1108,N_1041);
nor U3476 (N_3476,N_345,N_1507);
and U3477 (N_3477,N_849,N_1344);
nor U3478 (N_3478,N_554,N_2246);
and U3479 (N_3479,N_2055,N_1978);
or U3480 (N_3480,N_757,N_336);
nor U3481 (N_3481,N_2389,N_252);
or U3482 (N_3482,N_1720,N_812);
xor U3483 (N_3483,N_1356,N_1717);
nand U3484 (N_3484,N_1748,N_139);
nor U3485 (N_3485,N_1650,N_67);
and U3486 (N_3486,N_2305,N_1554);
nand U3487 (N_3487,N_936,N_281);
and U3488 (N_3488,N_685,N_1284);
nor U3489 (N_3489,N_681,N_885);
xor U3490 (N_3490,N_1769,N_464);
nand U3491 (N_3491,N_138,N_330);
nor U3492 (N_3492,N_1689,N_1113);
or U3493 (N_3493,N_881,N_697);
nand U3494 (N_3494,N_2218,N_2282);
and U3495 (N_3495,N_1129,N_863);
nor U3496 (N_3496,N_1969,N_1633);
xor U3497 (N_3497,N_1842,N_834);
nor U3498 (N_3498,N_2078,N_22);
nor U3499 (N_3499,N_1252,N_1053);
and U3500 (N_3500,N_1090,N_2211);
nand U3501 (N_3501,N_2149,N_726);
nor U3502 (N_3502,N_1003,N_943);
nor U3503 (N_3503,N_777,N_157);
and U3504 (N_3504,N_498,N_1829);
nand U3505 (N_3505,N_1006,N_879);
nand U3506 (N_3506,N_1803,N_1326);
or U3507 (N_3507,N_1361,N_2397);
or U3508 (N_3508,N_951,N_158);
nor U3509 (N_3509,N_953,N_241);
nor U3510 (N_3510,N_848,N_1877);
nand U3511 (N_3511,N_713,N_1659);
nor U3512 (N_3512,N_1425,N_143);
nor U3513 (N_3513,N_2387,N_2173);
nor U3514 (N_3514,N_632,N_1007);
or U3515 (N_3515,N_2341,N_731);
nand U3516 (N_3516,N_42,N_946);
xor U3517 (N_3517,N_2043,N_2322);
nand U3518 (N_3518,N_2146,N_1158);
and U3519 (N_3519,N_2332,N_1729);
nor U3520 (N_3520,N_323,N_2277);
nor U3521 (N_3521,N_1097,N_2133);
and U3522 (N_3522,N_730,N_1317);
nand U3523 (N_3523,N_146,N_1285);
and U3524 (N_3524,N_2048,N_1895);
or U3525 (N_3525,N_1536,N_314);
and U3526 (N_3526,N_1072,N_2064);
and U3527 (N_3527,N_1702,N_861);
nor U3528 (N_3528,N_333,N_293);
nand U3529 (N_3529,N_219,N_1558);
and U3530 (N_3530,N_1260,N_2034);
or U3531 (N_3531,N_2248,N_728);
nor U3532 (N_3532,N_2143,N_2356);
and U3533 (N_3533,N_481,N_805);
nor U3534 (N_3534,N_2135,N_304);
nor U3535 (N_3535,N_875,N_645);
nand U3536 (N_3536,N_2283,N_1778);
nor U3537 (N_3537,N_1229,N_1597);
or U3538 (N_3538,N_1820,N_2441);
nand U3539 (N_3539,N_2224,N_1772);
or U3540 (N_3540,N_843,N_1222);
nor U3541 (N_3541,N_1489,N_258);
nand U3542 (N_3542,N_1417,N_2016);
nand U3543 (N_3543,N_608,N_98);
nand U3544 (N_3544,N_109,N_904);
and U3545 (N_3545,N_2291,N_1886);
or U3546 (N_3546,N_2092,N_1251);
or U3547 (N_3547,N_2209,N_869);
xnor U3548 (N_3548,N_1568,N_909);
nor U3549 (N_3549,N_1932,N_508);
nor U3550 (N_3550,N_1095,N_1391);
nand U3551 (N_3551,N_74,N_1837);
nor U3552 (N_3552,N_338,N_275);
xnor U3553 (N_3553,N_2128,N_2150);
or U3554 (N_3554,N_991,N_1732);
and U3555 (N_3555,N_1082,N_1971);
nand U3556 (N_3556,N_114,N_822);
nand U3557 (N_3557,N_2117,N_934);
or U3558 (N_3558,N_1360,N_572);
and U3559 (N_3559,N_647,N_1292);
or U3560 (N_3560,N_1136,N_2039);
and U3561 (N_3561,N_2454,N_550);
and U3562 (N_3562,N_278,N_1442);
and U3563 (N_3563,N_1249,N_1299);
nand U3564 (N_3564,N_1067,N_1608);
nor U3565 (N_3565,N_766,N_661);
nor U3566 (N_3566,N_1767,N_1083);
and U3567 (N_3567,N_2313,N_2491);
nor U3568 (N_3568,N_1832,N_262);
nand U3569 (N_3569,N_1685,N_1532);
nor U3570 (N_3570,N_1287,N_249);
or U3571 (N_3571,N_351,N_765);
nor U3572 (N_3572,N_644,N_1363);
and U3573 (N_3573,N_901,N_368);
xnor U3574 (N_3574,N_1141,N_352);
nor U3575 (N_3575,N_2202,N_892);
and U3576 (N_3576,N_622,N_595);
or U3577 (N_3577,N_2114,N_1913);
or U3578 (N_3578,N_1513,N_1443);
or U3579 (N_3579,N_2244,N_2475);
nor U3580 (N_3580,N_2320,N_2470);
nor U3581 (N_3581,N_2460,N_2198);
nand U3582 (N_3582,N_652,N_1258);
nor U3583 (N_3583,N_491,N_2335);
nand U3584 (N_3584,N_1631,N_1128);
and U3585 (N_3585,N_1372,N_2482);
and U3586 (N_3586,N_1294,N_315);
or U3587 (N_3587,N_379,N_1550);
nand U3588 (N_3588,N_761,N_1304);
and U3589 (N_3589,N_2267,N_950);
nand U3590 (N_3590,N_119,N_1164);
or U3591 (N_3591,N_637,N_308);
nand U3592 (N_3592,N_2125,N_1460);
and U3593 (N_3593,N_2107,N_575);
and U3594 (N_3594,N_1802,N_1807);
nand U3595 (N_3595,N_2236,N_995);
and U3596 (N_3596,N_1999,N_1188);
xor U3597 (N_3597,N_2120,N_1870);
nor U3598 (N_3598,N_1074,N_2495);
nor U3599 (N_3599,N_264,N_1736);
nor U3600 (N_3600,N_1896,N_986);
or U3601 (N_3601,N_1393,N_155);
and U3602 (N_3602,N_2316,N_1804);
and U3603 (N_3603,N_2408,N_2296);
and U3604 (N_3604,N_2219,N_1573);
nor U3605 (N_3605,N_1279,N_1731);
and U3606 (N_3606,N_202,N_1553);
nor U3607 (N_3607,N_594,N_147);
nor U3608 (N_3608,N_807,N_759);
nor U3609 (N_3609,N_1859,N_476);
nor U3610 (N_3610,N_1795,N_597);
nand U3611 (N_3611,N_2433,N_448);
or U3612 (N_3612,N_2423,N_2104);
and U3613 (N_3613,N_489,N_667);
and U3614 (N_3614,N_770,N_1382);
xnor U3615 (N_3615,N_2473,N_1541);
nand U3616 (N_3616,N_1227,N_922);
nor U3617 (N_3617,N_465,N_1311);
and U3618 (N_3618,N_1661,N_855);
nor U3619 (N_3619,N_1040,N_1062);
nand U3620 (N_3620,N_1529,N_1543);
nor U3621 (N_3621,N_982,N_1540);
nand U3622 (N_3622,N_714,N_758);
nor U3623 (N_3623,N_864,N_1147);
or U3624 (N_3624,N_1020,N_1900);
nor U3625 (N_3625,N_12,N_64);
nor U3626 (N_3626,N_964,N_2100);
nand U3627 (N_3627,N_1115,N_1306);
nand U3628 (N_3628,N_1975,N_2424);
nor U3629 (N_3629,N_1555,N_2348);
and U3630 (N_3630,N_1273,N_362);
or U3631 (N_3631,N_2053,N_1692);
or U3632 (N_3632,N_1397,N_1834);
nand U3633 (N_3633,N_2184,N_2395);
or U3634 (N_3634,N_626,N_443);
and U3635 (N_3635,N_1831,N_553);
and U3636 (N_3636,N_1670,N_952);
and U3637 (N_3637,N_2279,N_2176);
and U3638 (N_3638,N_1039,N_1038);
xor U3639 (N_3639,N_355,N_131);
nand U3640 (N_3640,N_688,N_1187);
and U3641 (N_3641,N_161,N_136);
nor U3642 (N_3642,N_436,N_1501);
and U3643 (N_3643,N_1519,N_1257);
nor U3644 (N_3644,N_1477,N_440);
nand U3645 (N_3645,N_509,N_1029);
and U3646 (N_3646,N_565,N_1377);
nor U3647 (N_3647,N_1887,N_1629);
nor U3648 (N_3648,N_1828,N_188);
and U3649 (N_3649,N_2307,N_1737);
or U3650 (N_3650,N_1664,N_1959);
nor U3651 (N_3651,N_1430,N_1065);
or U3652 (N_3652,N_1508,N_2422);
and U3653 (N_3653,N_779,N_886);
nand U3654 (N_3654,N_1353,N_408);
or U3655 (N_3655,N_754,N_2216);
nor U3656 (N_3656,N_2415,N_992);
and U3657 (N_3657,N_280,N_1303);
or U3658 (N_3658,N_709,N_283);
or U3659 (N_3659,N_1875,N_1055);
nand U3660 (N_3660,N_2487,N_1623);
and U3661 (N_3661,N_2132,N_1321);
and U3662 (N_3662,N_1800,N_560);
or U3663 (N_3663,N_1996,N_1037);
or U3664 (N_3664,N_1816,N_897);
and U3665 (N_3665,N_1871,N_242);
or U3666 (N_3666,N_212,N_1645);
nand U3667 (N_3667,N_1351,N_1605);
xor U3668 (N_3668,N_148,N_1237);
and U3669 (N_3669,N_586,N_2206);
nand U3670 (N_3670,N_1856,N_958);
or U3671 (N_3671,N_873,N_63);
or U3672 (N_3672,N_1462,N_2243);
nand U3673 (N_3673,N_1034,N_789);
or U3674 (N_3674,N_198,N_325);
nand U3675 (N_3675,N_2174,N_285);
nor U3676 (N_3676,N_335,N_348);
or U3677 (N_3677,N_270,N_525);
nor U3678 (N_3678,N_1452,N_510);
and U3679 (N_3679,N_1787,N_648);
nor U3680 (N_3680,N_931,N_978);
nand U3681 (N_3681,N_47,N_1201);
xor U3682 (N_3682,N_2079,N_1545);
or U3683 (N_3683,N_1205,N_1934);
and U3684 (N_3684,N_2328,N_168);
and U3685 (N_3685,N_2180,N_1766);
xnor U3686 (N_3686,N_2417,N_993);
nor U3687 (N_3687,N_122,N_480);
xnor U3688 (N_3688,N_1497,N_401);
xor U3689 (N_3689,N_1655,N_2178);
and U3690 (N_3690,N_106,N_1024);
nand U3691 (N_3691,N_2121,N_328);
nor U3692 (N_3692,N_747,N_2401);
and U3693 (N_3693,N_1036,N_2270);
and U3694 (N_3694,N_14,N_781);
nand U3695 (N_3695,N_2003,N_1267);
and U3696 (N_3696,N_1419,N_1867);
or U3697 (N_3697,N_2385,N_431);
or U3698 (N_3698,N_326,N_1672);
and U3699 (N_3699,N_10,N_178);
or U3700 (N_3700,N_1388,N_2084);
or U3701 (N_3701,N_2447,N_1199);
or U3702 (N_3702,N_1014,N_1086);
nand U3703 (N_3703,N_2038,N_2481);
or U3704 (N_3704,N_916,N_1571);
or U3705 (N_3705,N_250,N_1794);
nand U3706 (N_3706,N_1916,N_735);
and U3707 (N_3707,N_2069,N_2111);
nand U3708 (N_3708,N_569,N_2301);
or U3709 (N_3709,N_698,N_828);
and U3710 (N_3710,N_2256,N_1473);
xor U3711 (N_3711,N_130,N_1202);
and U3712 (N_3712,N_2088,N_1781);
or U3713 (N_3713,N_773,N_2444);
xor U3714 (N_3714,N_1323,N_771);
nor U3715 (N_3715,N_163,N_1823);
and U3716 (N_3716,N_814,N_1663);
xnor U3717 (N_3717,N_865,N_1466);
xor U3718 (N_3718,N_1484,N_2147);
or U3719 (N_3719,N_701,N_503);
nor U3720 (N_3720,N_1546,N_228);
nor U3721 (N_3721,N_1509,N_1981);
nand U3722 (N_3722,N_531,N_100);
and U3723 (N_3723,N_2010,N_2484);
or U3724 (N_3724,N_1574,N_574);
nand U3725 (N_3725,N_2381,N_1984);
nand U3726 (N_3726,N_1312,N_870);
and U3727 (N_3727,N_1378,N_86);
and U3728 (N_3728,N_404,N_1274);
and U3729 (N_3729,N_1117,N_2362);
nand U3730 (N_3730,N_1449,N_2308);
and U3731 (N_3731,N_1511,N_1986);
or U3732 (N_3732,N_370,N_1850);
and U3733 (N_3733,N_2298,N_655);
nand U3734 (N_3734,N_2226,N_1265);
or U3735 (N_3735,N_788,N_364);
xnor U3736 (N_3736,N_360,N_1715);
or U3737 (N_3737,N_2271,N_908);
or U3738 (N_3738,N_33,N_738);
or U3739 (N_3739,N_989,N_1799);
and U3740 (N_3740,N_313,N_2479);
nor U3741 (N_3741,N_894,N_545);
nor U3742 (N_3742,N_225,N_366);
nor U3743 (N_3743,N_2001,N_1533);
and U3744 (N_3744,N_846,N_585);
nor U3745 (N_3745,N_1112,N_2028);
and U3746 (N_3746,N_1386,N_501);
nor U3747 (N_3747,N_1628,N_288);
and U3748 (N_3748,N_450,N_1218);
and U3749 (N_3749,N_563,N_1049);
nor U3750 (N_3750,N_1051,N_191);
or U3751 (N_3751,N_1337,N_1777);
and U3752 (N_3752,N_467,N_2176);
or U3753 (N_3753,N_1135,N_1477);
or U3754 (N_3754,N_916,N_1462);
nor U3755 (N_3755,N_1534,N_1502);
nand U3756 (N_3756,N_1950,N_1868);
and U3757 (N_3757,N_223,N_1740);
or U3758 (N_3758,N_2134,N_362);
nand U3759 (N_3759,N_436,N_717);
nand U3760 (N_3760,N_2386,N_2195);
nand U3761 (N_3761,N_1022,N_1727);
nor U3762 (N_3762,N_2012,N_1419);
nor U3763 (N_3763,N_1979,N_2029);
nor U3764 (N_3764,N_1229,N_1267);
and U3765 (N_3765,N_1803,N_1914);
and U3766 (N_3766,N_2070,N_697);
nor U3767 (N_3767,N_1120,N_1497);
nor U3768 (N_3768,N_883,N_1142);
nor U3769 (N_3769,N_1382,N_1934);
or U3770 (N_3770,N_2330,N_1479);
and U3771 (N_3771,N_269,N_1540);
nand U3772 (N_3772,N_2314,N_1867);
or U3773 (N_3773,N_25,N_796);
nand U3774 (N_3774,N_2133,N_1674);
nand U3775 (N_3775,N_289,N_1440);
and U3776 (N_3776,N_2482,N_600);
or U3777 (N_3777,N_960,N_190);
nor U3778 (N_3778,N_332,N_1568);
and U3779 (N_3779,N_542,N_2381);
nand U3780 (N_3780,N_403,N_1297);
or U3781 (N_3781,N_453,N_2055);
nand U3782 (N_3782,N_686,N_476);
xor U3783 (N_3783,N_1078,N_1671);
nor U3784 (N_3784,N_710,N_376);
and U3785 (N_3785,N_1337,N_118);
and U3786 (N_3786,N_998,N_1433);
and U3787 (N_3787,N_999,N_2188);
xnor U3788 (N_3788,N_893,N_243);
or U3789 (N_3789,N_1066,N_1143);
or U3790 (N_3790,N_630,N_215);
or U3791 (N_3791,N_2113,N_1380);
xor U3792 (N_3792,N_192,N_2495);
nor U3793 (N_3793,N_2364,N_2002);
and U3794 (N_3794,N_2004,N_168);
or U3795 (N_3795,N_2319,N_1893);
nor U3796 (N_3796,N_1568,N_2051);
nand U3797 (N_3797,N_151,N_593);
and U3798 (N_3798,N_1119,N_292);
nand U3799 (N_3799,N_108,N_2097);
nand U3800 (N_3800,N_190,N_1244);
nor U3801 (N_3801,N_657,N_436);
and U3802 (N_3802,N_283,N_1391);
xnor U3803 (N_3803,N_452,N_502);
or U3804 (N_3804,N_1096,N_298);
and U3805 (N_3805,N_2101,N_1526);
or U3806 (N_3806,N_1869,N_136);
nand U3807 (N_3807,N_753,N_2026);
and U3808 (N_3808,N_1874,N_887);
nand U3809 (N_3809,N_1709,N_2017);
or U3810 (N_3810,N_783,N_1797);
or U3811 (N_3811,N_366,N_2045);
xnor U3812 (N_3812,N_1641,N_1972);
or U3813 (N_3813,N_1017,N_1881);
nor U3814 (N_3814,N_2074,N_913);
xor U3815 (N_3815,N_2035,N_952);
nor U3816 (N_3816,N_1818,N_161);
xor U3817 (N_3817,N_1433,N_2122);
or U3818 (N_3818,N_1407,N_1252);
and U3819 (N_3819,N_901,N_1220);
nor U3820 (N_3820,N_1232,N_917);
and U3821 (N_3821,N_899,N_1087);
nand U3822 (N_3822,N_1160,N_495);
nand U3823 (N_3823,N_1466,N_1164);
or U3824 (N_3824,N_1147,N_1173);
or U3825 (N_3825,N_104,N_1374);
and U3826 (N_3826,N_1276,N_1190);
or U3827 (N_3827,N_2055,N_967);
xnor U3828 (N_3828,N_1967,N_1642);
or U3829 (N_3829,N_544,N_1970);
and U3830 (N_3830,N_306,N_1949);
nand U3831 (N_3831,N_2451,N_1873);
nor U3832 (N_3832,N_526,N_501);
or U3833 (N_3833,N_1101,N_27);
and U3834 (N_3834,N_520,N_2363);
nand U3835 (N_3835,N_1046,N_1537);
or U3836 (N_3836,N_367,N_1488);
nand U3837 (N_3837,N_840,N_1745);
nor U3838 (N_3838,N_2394,N_1090);
nor U3839 (N_3839,N_1316,N_171);
or U3840 (N_3840,N_1623,N_2357);
or U3841 (N_3841,N_201,N_1262);
nand U3842 (N_3842,N_2127,N_633);
and U3843 (N_3843,N_1681,N_856);
and U3844 (N_3844,N_767,N_841);
or U3845 (N_3845,N_2358,N_2256);
or U3846 (N_3846,N_1079,N_2277);
and U3847 (N_3847,N_1837,N_658);
nor U3848 (N_3848,N_2097,N_422);
or U3849 (N_3849,N_2375,N_1091);
nand U3850 (N_3850,N_2440,N_932);
and U3851 (N_3851,N_2192,N_2234);
or U3852 (N_3852,N_104,N_614);
and U3853 (N_3853,N_1637,N_924);
or U3854 (N_3854,N_1121,N_401);
and U3855 (N_3855,N_7,N_1272);
and U3856 (N_3856,N_1726,N_919);
or U3857 (N_3857,N_604,N_2381);
and U3858 (N_3858,N_2086,N_848);
and U3859 (N_3859,N_1973,N_1729);
nor U3860 (N_3860,N_802,N_1108);
xor U3861 (N_3861,N_511,N_71);
or U3862 (N_3862,N_345,N_698);
and U3863 (N_3863,N_160,N_22);
nand U3864 (N_3864,N_802,N_25);
nor U3865 (N_3865,N_2210,N_1618);
nor U3866 (N_3866,N_145,N_98);
or U3867 (N_3867,N_2000,N_592);
nor U3868 (N_3868,N_1150,N_1297);
nand U3869 (N_3869,N_464,N_642);
nor U3870 (N_3870,N_196,N_458);
and U3871 (N_3871,N_2025,N_242);
xnor U3872 (N_3872,N_1360,N_454);
and U3873 (N_3873,N_1415,N_292);
and U3874 (N_3874,N_530,N_1369);
nand U3875 (N_3875,N_2227,N_1259);
nand U3876 (N_3876,N_2136,N_387);
nand U3877 (N_3877,N_509,N_160);
or U3878 (N_3878,N_585,N_956);
nand U3879 (N_3879,N_2374,N_1438);
nor U3880 (N_3880,N_481,N_769);
nand U3881 (N_3881,N_1162,N_1157);
nand U3882 (N_3882,N_548,N_829);
and U3883 (N_3883,N_1064,N_1146);
nand U3884 (N_3884,N_1235,N_855);
or U3885 (N_3885,N_1713,N_482);
nand U3886 (N_3886,N_2325,N_250);
nor U3887 (N_3887,N_1951,N_1344);
nor U3888 (N_3888,N_628,N_141);
and U3889 (N_3889,N_695,N_1678);
xor U3890 (N_3890,N_225,N_789);
nor U3891 (N_3891,N_1684,N_1575);
and U3892 (N_3892,N_962,N_2286);
xor U3893 (N_3893,N_2171,N_985);
nand U3894 (N_3894,N_1336,N_223);
and U3895 (N_3895,N_63,N_1891);
or U3896 (N_3896,N_264,N_664);
nor U3897 (N_3897,N_342,N_846);
nor U3898 (N_3898,N_1699,N_2243);
nand U3899 (N_3899,N_2442,N_2313);
nor U3900 (N_3900,N_240,N_1172);
xnor U3901 (N_3901,N_2080,N_187);
and U3902 (N_3902,N_2139,N_1799);
nor U3903 (N_3903,N_1945,N_82);
or U3904 (N_3904,N_2281,N_1160);
and U3905 (N_3905,N_2433,N_2389);
or U3906 (N_3906,N_1458,N_6);
and U3907 (N_3907,N_726,N_1277);
and U3908 (N_3908,N_1901,N_35);
and U3909 (N_3909,N_2470,N_1881);
xor U3910 (N_3910,N_1806,N_771);
or U3911 (N_3911,N_273,N_1253);
or U3912 (N_3912,N_247,N_2183);
nand U3913 (N_3913,N_1403,N_1620);
nand U3914 (N_3914,N_151,N_75);
or U3915 (N_3915,N_1066,N_484);
nor U3916 (N_3916,N_1198,N_1974);
nand U3917 (N_3917,N_2104,N_1941);
nor U3918 (N_3918,N_2181,N_2490);
xor U3919 (N_3919,N_2129,N_257);
and U3920 (N_3920,N_1974,N_2249);
nand U3921 (N_3921,N_217,N_1123);
nor U3922 (N_3922,N_1307,N_2304);
or U3923 (N_3923,N_2317,N_275);
xor U3924 (N_3924,N_920,N_1552);
xor U3925 (N_3925,N_1589,N_218);
nor U3926 (N_3926,N_913,N_2048);
nand U3927 (N_3927,N_1420,N_189);
and U3928 (N_3928,N_245,N_1875);
nand U3929 (N_3929,N_1650,N_163);
nand U3930 (N_3930,N_618,N_606);
nor U3931 (N_3931,N_1210,N_1569);
nor U3932 (N_3932,N_1952,N_2249);
nor U3933 (N_3933,N_2244,N_766);
or U3934 (N_3934,N_2258,N_2241);
and U3935 (N_3935,N_2147,N_2463);
nand U3936 (N_3936,N_2163,N_2359);
nor U3937 (N_3937,N_511,N_713);
nand U3938 (N_3938,N_270,N_577);
and U3939 (N_3939,N_1178,N_2044);
and U3940 (N_3940,N_859,N_623);
nor U3941 (N_3941,N_1571,N_810);
and U3942 (N_3942,N_603,N_1468);
nor U3943 (N_3943,N_932,N_1263);
nor U3944 (N_3944,N_745,N_1300);
nor U3945 (N_3945,N_1670,N_87);
or U3946 (N_3946,N_2167,N_196);
or U3947 (N_3947,N_66,N_242);
nand U3948 (N_3948,N_138,N_2316);
or U3949 (N_3949,N_2023,N_2479);
and U3950 (N_3950,N_1713,N_1379);
nand U3951 (N_3951,N_1186,N_2359);
nor U3952 (N_3952,N_2443,N_1540);
and U3953 (N_3953,N_1197,N_613);
xnor U3954 (N_3954,N_1451,N_166);
or U3955 (N_3955,N_97,N_517);
or U3956 (N_3956,N_1542,N_135);
or U3957 (N_3957,N_1277,N_1812);
nor U3958 (N_3958,N_1616,N_1267);
nand U3959 (N_3959,N_572,N_989);
or U3960 (N_3960,N_1324,N_1133);
and U3961 (N_3961,N_1122,N_1207);
nand U3962 (N_3962,N_395,N_736);
and U3963 (N_3963,N_28,N_2266);
nor U3964 (N_3964,N_249,N_1789);
nor U3965 (N_3965,N_1647,N_2292);
nor U3966 (N_3966,N_1986,N_938);
and U3967 (N_3967,N_2486,N_652);
and U3968 (N_3968,N_1839,N_1547);
nor U3969 (N_3969,N_1938,N_1013);
or U3970 (N_3970,N_1594,N_1363);
xnor U3971 (N_3971,N_2072,N_2346);
and U3972 (N_3972,N_1175,N_257);
nand U3973 (N_3973,N_1996,N_128);
nand U3974 (N_3974,N_873,N_584);
or U3975 (N_3975,N_2241,N_2319);
and U3976 (N_3976,N_1246,N_1219);
and U3977 (N_3977,N_350,N_2498);
nor U3978 (N_3978,N_2478,N_1206);
or U3979 (N_3979,N_1257,N_1399);
and U3980 (N_3980,N_2028,N_735);
and U3981 (N_3981,N_184,N_2162);
nor U3982 (N_3982,N_419,N_1132);
and U3983 (N_3983,N_1144,N_1632);
and U3984 (N_3984,N_857,N_763);
nor U3985 (N_3985,N_1134,N_1899);
or U3986 (N_3986,N_390,N_1933);
and U3987 (N_3987,N_1029,N_634);
and U3988 (N_3988,N_1697,N_2122);
nand U3989 (N_3989,N_70,N_2364);
and U3990 (N_3990,N_1537,N_1410);
or U3991 (N_3991,N_815,N_1908);
nand U3992 (N_3992,N_2462,N_1851);
nand U3993 (N_3993,N_1185,N_313);
nor U3994 (N_3994,N_2113,N_1108);
nand U3995 (N_3995,N_1867,N_29);
and U3996 (N_3996,N_1981,N_693);
xor U3997 (N_3997,N_345,N_2374);
nor U3998 (N_3998,N_1466,N_623);
nor U3999 (N_3999,N_192,N_1282);
and U4000 (N_4000,N_1728,N_387);
nor U4001 (N_4001,N_1791,N_1118);
and U4002 (N_4002,N_2392,N_1581);
nor U4003 (N_4003,N_1233,N_1866);
or U4004 (N_4004,N_2211,N_429);
or U4005 (N_4005,N_1331,N_624);
xnor U4006 (N_4006,N_575,N_531);
nand U4007 (N_4007,N_2491,N_2253);
nand U4008 (N_4008,N_1269,N_623);
and U4009 (N_4009,N_2202,N_2248);
and U4010 (N_4010,N_1387,N_712);
nor U4011 (N_4011,N_703,N_1937);
or U4012 (N_4012,N_1327,N_76);
nor U4013 (N_4013,N_1014,N_1615);
or U4014 (N_4014,N_707,N_2478);
nand U4015 (N_4015,N_532,N_2404);
nand U4016 (N_4016,N_745,N_1575);
xor U4017 (N_4017,N_585,N_1570);
or U4018 (N_4018,N_1072,N_528);
nand U4019 (N_4019,N_1644,N_735);
or U4020 (N_4020,N_260,N_1270);
nor U4021 (N_4021,N_1935,N_716);
or U4022 (N_4022,N_1406,N_252);
nand U4023 (N_4023,N_2029,N_1712);
or U4024 (N_4024,N_147,N_1211);
nor U4025 (N_4025,N_2125,N_1161);
or U4026 (N_4026,N_2188,N_1664);
and U4027 (N_4027,N_1858,N_2030);
nor U4028 (N_4028,N_2178,N_1918);
nor U4029 (N_4029,N_1828,N_1449);
nor U4030 (N_4030,N_1938,N_567);
nor U4031 (N_4031,N_1947,N_820);
xnor U4032 (N_4032,N_2409,N_438);
or U4033 (N_4033,N_1986,N_2140);
or U4034 (N_4034,N_27,N_1660);
and U4035 (N_4035,N_1167,N_1602);
nand U4036 (N_4036,N_1592,N_1362);
or U4037 (N_4037,N_1872,N_1457);
or U4038 (N_4038,N_1787,N_1164);
xor U4039 (N_4039,N_215,N_913);
and U4040 (N_4040,N_934,N_87);
nor U4041 (N_4041,N_443,N_631);
nand U4042 (N_4042,N_1290,N_561);
nor U4043 (N_4043,N_352,N_77);
nor U4044 (N_4044,N_1842,N_2229);
nor U4045 (N_4045,N_840,N_2175);
nand U4046 (N_4046,N_909,N_34);
nand U4047 (N_4047,N_815,N_1956);
and U4048 (N_4048,N_371,N_2174);
nor U4049 (N_4049,N_1650,N_1577);
or U4050 (N_4050,N_1095,N_1178);
nand U4051 (N_4051,N_151,N_1522);
nand U4052 (N_4052,N_1444,N_1152);
nand U4053 (N_4053,N_1456,N_131);
and U4054 (N_4054,N_1531,N_2237);
and U4055 (N_4055,N_525,N_1696);
or U4056 (N_4056,N_2197,N_1102);
xnor U4057 (N_4057,N_1501,N_2498);
or U4058 (N_4058,N_1462,N_910);
or U4059 (N_4059,N_1456,N_1298);
nor U4060 (N_4060,N_1288,N_655);
nor U4061 (N_4061,N_1206,N_529);
and U4062 (N_4062,N_247,N_2082);
xor U4063 (N_4063,N_1660,N_1076);
or U4064 (N_4064,N_488,N_713);
nor U4065 (N_4065,N_144,N_606);
nor U4066 (N_4066,N_2485,N_723);
nand U4067 (N_4067,N_1864,N_262);
nor U4068 (N_4068,N_39,N_1443);
nand U4069 (N_4069,N_2446,N_887);
xor U4070 (N_4070,N_2183,N_1490);
nor U4071 (N_4071,N_1129,N_1585);
nor U4072 (N_4072,N_2490,N_2054);
nor U4073 (N_4073,N_156,N_622);
nor U4074 (N_4074,N_521,N_323);
nor U4075 (N_4075,N_1910,N_797);
nor U4076 (N_4076,N_108,N_1859);
nor U4077 (N_4077,N_949,N_1324);
or U4078 (N_4078,N_1362,N_1731);
or U4079 (N_4079,N_1333,N_2318);
or U4080 (N_4080,N_1826,N_1808);
nor U4081 (N_4081,N_2106,N_572);
nor U4082 (N_4082,N_1395,N_1487);
nor U4083 (N_4083,N_981,N_284);
nor U4084 (N_4084,N_1883,N_833);
nor U4085 (N_4085,N_2313,N_715);
and U4086 (N_4086,N_1707,N_110);
nor U4087 (N_4087,N_173,N_691);
nand U4088 (N_4088,N_1290,N_806);
xor U4089 (N_4089,N_2202,N_177);
and U4090 (N_4090,N_813,N_1642);
xor U4091 (N_4091,N_178,N_2213);
nor U4092 (N_4092,N_1965,N_2166);
or U4093 (N_4093,N_1119,N_2262);
or U4094 (N_4094,N_1598,N_1586);
or U4095 (N_4095,N_678,N_1057);
or U4096 (N_4096,N_413,N_2225);
nor U4097 (N_4097,N_21,N_2176);
nor U4098 (N_4098,N_1872,N_92);
and U4099 (N_4099,N_391,N_20);
nor U4100 (N_4100,N_2059,N_1997);
nor U4101 (N_4101,N_2000,N_1571);
nor U4102 (N_4102,N_1319,N_1562);
nor U4103 (N_4103,N_87,N_412);
and U4104 (N_4104,N_1485,N_98);
nor U4105 (N_4105,N_24,N_1440);
nand U4106 (N_4106,N_66,N_389);
nor U4107 (N_4107,N_875,N_1115);
and U4108 (N_4108,N_59,N_130);
nor U4109 (N_4109,N_336,N_138);
nor U4110 (N_4110,N_1154,N_435);
nand U4111 (N_4111,N_1278,N_529);
nor U4112 (N_4112,N_353,N_2275);
nand U4113 (N_4113,N_1176,N_2158);
or U4114 (N_4114,N_1777,N_210);
nor U4115 (N_4115,N_527,N_258);
nand U4116 (N_4116,N_1771,N_2487);
nand U4117 (N_4117,N_2446,N_873);
nor U4118 (N_4118,N_2012,N_1617);
or U4119 (N_4119,N_655,N_904);
nand U4120 (N_4120,N_2149,N_1337);
nor U4121 (N_4121,N_1834,N_309);
or U4122 (N_4122,N_1017,N_1064);
and U4123 (N_4123,N_1710,N_1630);
and U4124 (N_4124,N_855,N_1153);
nand U4125 (N_4125,N_1511,N_951);
nor U4126 (N_4126,N_2052,N_372);
nand U4127 (N_4127,N_496,N_43);
nor U4128 (N_4128,N_1076,N_2320);
or U4129 (N_4129,N_928,N_1784);
and U4130 (N_4130,N_30,N_802);
xnor U4131 (N_4131,N_870,N_878);
nand U4132 (N_4132,N_490,N_2207);
and U4133 (N_4133,N_446,N_1346);
nand U4134 (N_4134,N_128,N_543);
nor U4135 (N_4135,N_350,N_995);
and U4136 (N_4136,N_2387,N_966);
xor U4137 (N_4137,N_1616,N_1910);
nor U4138 (N_4138,N_1609,N_2012);
and U4139 (N_4139,N_2362,N_782);
or U4140 (N_4140,N_1314,N_1390);
nand U4141 (N_4141,N_1669,N_682);
and U4142 (N_4142,N_1675,N_456);
nor U4143 (N_4143,N_1818,N_1731);
nor U4144 (N_4144,N_2094,N_2271);
and U4145 (N_4145,N_601,N_1197);
nor U4146 (N_4146,N_861,N_1668);
nor U4147 (N_4147,N_1514,N_2186);
nand U4148 (N_4148,N_276,N_899);
or U4149 (N_4149,N_87,N_44);
and U4150 (N_4150,N_1200,N_1801);
or U4151 (N_4151,N_1308,N_2157);
and U4152 (N_4152,N_2352,N_192);
nand U4153 (N_4153,N_1359,N_546);
nand U4154 (N_4154,N_1291,N_2480);
or U4155 (N_4155,N_17,N_1661);
and U4156 (N_4156,N_610,N_618);
nand U4157 (N_4157,N_1621,N_1023);
nor U4158 (N_4158,N_1313,N_2095);
and U4159 (N_4159,N_1886,N_1171);
nor U4160 (N_4160,N_1836,N_1215);
and U4161 (N_4161,N_1708,N_1735);
or U4162 (N_4162,N_1708,N_1258);
nor U4163 (N_4163,N_652,N_297);
nor U4164 (N_4164,N_1551,N_2163);
xor U4165 (N_4165,N_976,N_2465);
nor U4166 (N_4166,N_1909,N_524);
xnor U4167 (N_4167,N_1435,N_1156);
nor U4168 (N_4168,N_1420,N_713);
and U4169 (N_4169,N_1578,N_1317);
and U4170 (N_4170,N_154,N_2259);
or U4171 (N_4171,N_445,N_1759);
and U4172 (N_4172,N_524,N_2310);
and U4173 (N_4173,N_2315,N_209);
or U4174 (N_4174,N_2183,N_2414);
or U4175 (N_4175,N_467,N_1468);
nor U4176 (N_4176,N_119,N_1411);
nor U4177 (N_4177,N_2071,N_1095);
nand U4178 (N_4178,N_1342,N_674);
nand U4179 (N_4179,N_689,N_1183);
xnor U4180 (N_4180,N_1796,N_2012);
nand U4181 (N_4181,N_527,N_1877);
or U4182 (N_4182,N_1718,N_2205);
nor U4183 (N_4183,N_1024,N_97);
nor U4184 (N_4184,N_253,N_2324);
and U4185 (N_4185,N_837,N_1119);
and U4186 (N_4186,N_2181,N_505);
xnor U4187 (N_4187,N_552,N_1429);
and U4188 (N_4188,N_2494,N_1960);
and U4189 (N_4189,N_2257,N_1427);
nor U4190 (N_4190,N_1031,N_1774);
xnor U4191 (N_4191,N_1876,N_2319);
or U4192 (N_4192,N_1274,N_2043);
nor U4193 (N_4193,N_92,N_772);
nor U4194 (N_4194,N_1323,N_2433);
nand U4195 (N_4195,N_2245,N_1250);
xnor U4196 (N_4196,N_524,N_455);
or U4197 (N_4197,N_1187,N_1743);
xnor U4198 (N_4198,N_962,N_779);
or U4199 (N_4199,N_2305,N_827);
nor U4200 (N_4200,N_1296,N_2398);
nand U4201 (N_4201,N_2272,N_629);
nor U4202 (N_4202,N_1212,N_982);
or U4203 (N_4203,N_1128,N_61);
nor U4204 (N_4204,N_2253,N_1188);
and U4205 (N_4205,N_361,N_1070);
nor U4206 (N_4206,N_1445,N_1674);
or U4207 (N_4207,N_1978,N_725);
or U4208 (N_4208,N_41,N_1655);
nor U4209 (N_4209,N_1236,N_74);
or U4210 (N_4210,N_1424,N_677);
nand U4211 (N_4211,N_1213,N_2418);
or U4212 (N_4212,N_1368,N_2350);
nand U4213 (N_4213,N_2499,N_960);
or U4214 (N_4214,N_2156,N_998);
nand U4215 (N_4215,N_1920,N_176);
or U4216 (N_4216,N_819,N_1813);
and U4217 (N_4217,N_1025,N_1544);
or U4218 (N_4218,N_1861,N_2043);
nand U4219 (N_4219,N_627,N_2471);
and U4220 (N_4220,N_768,N_970);
or U4221 (N_4221,N_228,N_604);
or U4222 (N_4222,N_568,N_1348);
nor U4223 (N_4223,N_635,N_403);
or U4224 (N_4224,N_292,N_1107);
and U4225 (N_4225,N_1721,N_1083);
and U4226 (N_4226,N_498,N_1637);
nor U4227 (N_4227,N_1700,N_610);
xnor U4228 (N_4228,N_2313,N_2156);
or U4229 (N_4229,N_1383,N_1772);
nor U4230 (N_4230,N_1443,N_991);
nand U4231 (N_4231,N_1630,N_569);
nor U4232 (N_4232,N_979,N_725);
nor U4233 (N_4233,N_925,N_1038);
nor U4234 (N_4234,N_1693,N_437);
nand U4235 (N_4235,N_1002,N_1792);
or U4236 (N_4236,N_918,N_1766);
or U4237 (N_4237,N_1854,N_2454);
or U4238 (N_4238,N_2044,N_876);
nor U4239 (N_4239,N_770,N_1543);
or U4240 (N_4240,N_1431,N_1399);
or U4241 (N_4241,N_987,N_1835);
and U4242 (N_4242,N_2461,N_2101);
nand U4243 (N_4243,N_1246,N_1197);
nor U4244 (N_4244,N_721,N_1602);
or U4245 (N_4245,N_1089,N_1239);
nor U4246 (N_4246,N_557,N_180);
nor U4247 (N_4247,N_2275,N_1215);
nor U4248 (N_4248,N_1816,N_385);
nor U4249 (N_4249,N_512,N_1081);
nor U4250 (N_4250,N_1209,N_1503);
and U4251 (N_4251,N_1448,N_116);
and U4252 (N_4252,N_798,N_822);
or U4253 (N_4253,N_1051,N_2448);
nor U4254 (N_4254,N_1174,N_1856);
xor U4255 (N_4255,N_28,N_1565);
or U4256 (N_4256,N_1382,N_937);
nor U4257 (N_4257,N_50,N_934);
nand U4258 (N_4258,N_521,N_2085);
nor U4259 (N_4259,N_179,N_440);
or U4260 (N_4260,N_562,N_647);
and U4261 (N_4261,N_14,N_110);
nand U4262 (N_4262,N_1466,N_795);
or U4263 (N_4263,N_1335,N_1607);
and U4264 (N_4264,N_753,N_97);
and U4265 (N_4265,N_1514,N_2123);
and U4266 (N_4266,N_1846,N_868);
and U4267 (N_4267,N_873,N_1238);
or U4268 (N_4268,N_1512,N_1638);
or U4269 (N_4269,N_277,N_1310);
xor U4270 (N_4270,N_1842,N_2414);
nor U4271 (N_4271,N_436,N_1560);
xnor U4272 (N_4272,N_179,N_1998);
nor U4273 (N_4273,N_1585,N_2194);
and U4274 (N_4274,N_2032,N_1352);
nor U4275 (N_4275,N_979,N_740);
xnor U4276 (N_4276,N_173,N_499);
nor U4277 (N_4277,N_48,N_201);
nand U4278 (N_4278,N_871,N_2326);
or U4279 (N_4279,N_811,N_1437);
and U4280 (N_4280,N_136,N_1759);
and U4281 (N_4281,N_1615,N_1186);
nor U4282 (N_4282,N_1039,N_755);
and U4283 (N_4283,N_286,N_1248);
nor U4284 (N_4284,N_666,N_2369);
and U4285 (N_4285,N_346,N_2016);
nand U4286 (N_4286,N_1072,N_663);
or U4287 (N_4287,N_2113,N_846);
and U4288 (N_4288,N_566,N_2108);
or U4289 (N_4289,N_2252,N_477);
xnor U4290 (N_4290,N_2150,N_256);
xor U4291 (N_4291,N_1188,N_2067);
nand U4292 (N_4292,N_1012,N_476);
and U4293 (N_4293,N_108,N_2126);
or U4294 (N_4294,N_1476,N_1432);
and U4295 (N_4295,N_20,N_1644);
nand U4296 (N_4296,N_1187,N_1970);
nor U4297 (N_4297,N_2416,N_1728);
xor U4298 (N_4298,N_861,N_1732);
nor U4299 (N_4299,N_899,N_1696);
or U4300 (N_4300,N_278,N_367);
nand U4301 (N_4301,N_826,N_876);
nor U4302 (N_4302,N_253,N_1580);
nand U4303 (N_4303,N_2368,N_342);
and U4304 (N_4304,N_1259,N_2049);
and U4305 (N_4305,N_91,N_650);
and U4306 (N_4306,N_1084,N_778);
or U4307 (N_4307,N_2425,N_1977);
and U4308 (N_4308,N_73,N_1856);
nand U4309 (N_4309,N_1988,N_2336);
nand U4310 (N_4310,N_874,N_1443);
nand U4311 (N_4311,N_648,N_1015);
and U4312 (N_4312,N_957,N_1657);
nand U4313 (N_4313,N_962,N_1343);
or U4314 (N_4314,N_1299,N_1089);
nor U4315 (N_4315,N_1418,N_768);
and U4316 (N_4316,N_438,N_70);
and U4317 (N_4317,N_1588,N_951);
or U4318 (N_4318,N_2157,N_2448);
nor U4319 (N_4319,N_367,N_1184);
or U4320 (N_4320,N_30,N_99);
and U4321 (N_4321,N_1243,N_1460);
xnor U4322 (N_4322,N_958,N_487);
and U4323 (N_4323,N_808,N_50);
nor U4324 (N_4324,N_826,N_620);
nor U4325 (N_4325,N_1603,N_2036);
and U4326 (N_4326,N_1356,N_2051);
and U4327 (N_4327,N_2125,N_135);
nand U4328 (N_4328,N_1442,N_1966);
nor U4329 (N_4329,N_2370,N_1725);
nand U4330 (N_4330,N_1761,N_1419);
and U4331 (N_4331,N_1394,N_424);
and U4332 (N_4332,N_89,N_543);
and U4333 (N_4333,N_338,N_19);
nand U4334 (N_4334,N_322,N_783);
and U4335 (N_4335,N_2030,N_2489);
nor U4336 (N_4336,N_885,N_1481);
nand U4337 (N_4337,N_1047,N_812);
nor U4338 (N_4338,N_1875,N_629);
nand U4339 (N_4339,N_772,N_1807);
nor U4340 (N_4340,N_1844,N_1704);
or U4341 (N_4341,N_1314,N_815);
and U4342 (N_4342,N_1349,N_1750);
and U4343 (N_4343,N_1423,N_955);
nor U4344 (N_4344,N_266,N_676);
and U4345 (N_4345,N_1627,N_2160);
nor U4346 (N_4346,N_1029,N_1419);
or U4347 (N_4347,N_2170,N_177);
nand U4348 (N_4348,N_798,N_1655);
xor U4349 (N_4349,N_763,N_2312);
nand U4350 (N_4350,N_1772,N_931);
nand U4351 (N_4351,N_765,N_378);
nor U4352 (N_4352,N_1421,N_1208);
and U4353 (N_4353,N_1466,N_335);
and U4354 (N_4354,N_1654,N_2206);
and U4355 (N_4355,N_187,N_2287);
nand U4356 (N_4356,N_1589,N_1766);
or U4357 (N_4357,N_983,N_32);
nor U4358 (N_4358,N_833,N_1188);
or U4359 (N_4359,N_938,N_1740);
xnor U4360 (N_4360,N_496,N_462);
or U4361 (N_4361,N_1817,N_933);
nor U4362 (N_4362,N_9,N_435);
nand U4363 (N_4363,N_867,N_164);
xnor U4364 (N_4364,N_2203,N_1346);
nand U4365 (N_4365,N_1150,N_1788);
and U4366 (N_4366,N_581,N_2288);
nand U4367 (N_4367,N_1667,N_1564);
nand U4368 (N_4368,N_1416,N_155);
and U4369 (N_4369,N_481,N_1674);
or U4370 (N_4370,N_2290,N_228);
or U4371 (N_4371,N_1225,N_1399);
and U4372 (N_4372,N_88,N_545);
or U4373 (N_4373,N_530,N_906);
or U4374 (N_4374,N_867,N_410);
and U4375 (N_4375,N_2083,N_1259);
nor U4376 (N_4376,N_768,N_2361);
or U4377 (N_4377,N_538,N_20);
nor U4378 (N_4378,N_32,N_2061);
nand U4379 (N_4379,N_834,N_765);
and U4380 (N_4380,N_1916,N_1573);
nor U4381 (N_4381,N_817,N_2244);
or U4382 (N_4382,N_1476,N_1757);
nor U4383 (N_4383,N_838,N_1304);
nor U4384 (N_4384,N_2339,N_881);
xnor U4385 (N_4385,N_2126,N_2240);
nand U4386 (N_4386,N_49,N_1098);
nor U4387 (N_4387,N_260,N_2130);
and U4388 (N_4388,N_66,N_1913);
and U4389 (N_4389,N_1129,N_1036);
and U4390 (N_4390,N_1845,N_765);
or U4391 (N_4391,N_2108,N_767);
or U4392 (N_4392,N_398,N_2060);
and U4393 (N_4393,N_2446,N_1599);
or U4394 (N_4394,N_1948,N_1927);
nor U4395 (N_4395,N_1891,N_546);
xnor U4396 (N_4396,N_851,N_708);
nand U4397 (N_4397,N_1811,N_74);
or U4398 (N_4398,N_1194,N_1259);
or U4399 (N_4399,N_1847,N_1886);
nor U4400 (N_4400,N_531,N_161);
and U4401 (N_4401,N_1389,N_513);
and U4402 (N_4402,N_1854,N_112);
or U4403 (N_4403,N_1870,N_1923);
and U4404 (N_4404,N_1787,N_2049);
and U4405 (N_4405,N_497,N_996);
nand U4406 (N_4406,N_1673,N_232);
nor U4407 (N_4407,N_348,N_1686);
nor U4408 (N_4408,N_742,N_303);
and U4409 (N_4409,N_2417,N_2477);
xor U4410 (N_4410,N_264,N_1580);
or U4411 (N_4411,N_1604,N_1629);
or U4412 (N_4412,N_845,N_619);
nand U4413 (N_4413,N_807,N_1717);
and U4414 (N_4414,N_905,N_1405);
and U4415 (N_4415,N_229,N_1377);
or U4416 (N_4416,N_76,N_1392);
nor U4417 (N_4417,N_1102,N_445);
nor U4418 (N_4418,N_1828,N_2194);
and U4419 (N_4419,N_1370,N_1692);
or U4420 (N_4420,N_801,N_1703);
or U4421 (N_4421,N_2076,N_1415);
nand U4422 (N_4422,N_1498,N_746);
nand U4423 (N_4423,N_1706,N_241);
and U4424 (N_4424,N_899,N_1631);
and U4425 (N_4425,N_2195,N_987);
nand U4426 (N_4426,N_32,N_2137);
or U4427 (N_4427,N_684,N_952);
or U4428 (N_4428,N_2432,N_1135);
or U4429 (N_4429,N_180,N_2283);
or U4430 (N_4430,N_1528,N_77);
nor U4431 (N_4431,N_113,N_626);
nor U4432 (N_4432,N_690,N_966);
or U4433 (N_4433,N_1816,N_486);
or U4434 (N_4434,N_1553,N_1923);
nand U4435 (N_4435,N_550,N_2485);
nor U4436 (N_4436,N_1084,N_1994);
or U4437 (N_4437,N_875,N_148);
xor U4438 (N_4438,N_1361,N_2206);
nand U4439 (N_4439,N_2467,N_1068);
and U4440 (N_4440,N_1846,N_2145);
or U4441 (N_4441,N_2288,N_1982);
or U4442 (N_4442,N_2304,N_506);
nor U4443 (N_4443,N_1872,N_1466);
and U4444 (N_4444,N_2453,N_533);
and U4445 (N_4445,N_857,N_2224);
nand U4446 (N_4446,N_50,N_792);
nand U4447 (N_4447,N_1345,N_27);
nor U4448 (N_4448,N_2185,N_1565);
and U4449 (N_4449,N_767,N_1842);
nand U4450 (N_4450,N_1988,N_36);
or U4451 (N_4451,N_817,N_2450);
and U4452 (N_4452,N_1280,N_2390);
or U4453 (N_4453,N_894,N_1310);
nor U4454 (N_4454,N_580,N_1206);
and U4455 (N_4455,N_707,N_999);
and U4456 (N_4456,N_1426,N_878);
and U4457 (N_4457,N_1392,N_2248);
nand U4458 (N_4458,N_1153,N_2163);
nand U4459 (N_4459,N_887,N_1559);
or U4460 (N_4460,N_79,N_571);
xnor U4461 (N_4461,N_2477,N_1362);
or U4462 (N_4462,N_1662,N_2136);
nand U4463 (N_4463,N_390,N_631);
nor U4464 (N_4464,N_56,N_2085);
and U4465 (N_4465,N_154,N_1337);
and U4466 (N_4466,N_64,N_2124);
or U4467 (N_4467,N_1495,N_529);
nand U4468 (N_4468,N_1852,N_264);
or U4469 (N_4469,N_608,N_1266);
nor U4470 (N_4470,N_1587,N_779);
or U4471 (N_4471,N_1466,N_2136);
nand U4472 (N_4472,N_1175,N_2306);
nor U4473 (N_4473,N_876,N_2251);
and U4474 (N_4474,N_593,N_1145);
nor U4475 (N_4475,N_2008,N_2372);
nand U4476 (N_4476,N_1291,N_36);
nor U4477 (N_4477,N_1265,N_183);
nand U4478 (N_4478,N_1941,N_1784);
or U4479 (N_4479,N_803,N_1887);
and U4480 (N_4480,N_1991,N_621);
xnor U4481 (N_4481,N_126,N_444);
nand U4482 (N_4482,N_2093,N_1846);
nor U4483 (N_4483,N_619,N_1186);
nor U4484 (N_4484,N_1426,N_1877);
nand U4485 (N_4485,N_793,N_923);
and U4486 (N_4486,N_2398,N_31);
nor U4487 (N_4487,N_510,N_868);
or U4488 (N_4488,N_750,N_29);
xnor U4489 (N_4489,N_1708,N_234);
nand U4490 (N_4490,N_396,N_2218);
xnor U4491 (N_4491,N_273,N_717);
or U4492 (N_4492,N_362,N_1448);
nor U4493 (N_4493,N_1944,N_1753);
nand U4494 (N_4494,N_2061,N_1574);
or U4495 (N_4495,N_469,N_683);
nand U4496 (N_4496,N_300,N_367);
and U4497 (N_4497,N_62,N_1237);
nand U4498 (N_4498,N_36,N_858);
or U4499 (N_4499,N_1254,N_2258);
nand U4500 (N_4500,N_1827,N_2346);
xor U4501 (N_4501,N_744,N_1711);
nor U4502 (N_4502,N_926,N_801);
nand U4503 (N_4503,N_492,N_2349);
and U4504 (N_4504,N_1783,N_2409);
and U4505 (N_4505,N_1914,N_17);
nand U4506 (N_4506,N_1191,N_2027);
or U4507 (N_4507,N_1298,N_2016);
or U4508 (N_4508,N_501,N_2095);
xor U4509 (N_4509,N_1114,N_2223);
and U4510 (N_4510,N_1509,N_1935);
and U4511 (N_4511,N_1038,N_400);
and U4512 (N_4512,N_16,N_1719);
or U4513 (N_4513,N_2464,N_1853);
nand U4514 (N_4514,N_940,N_2408);
or U4515 (N_4515,N_575,N_1897);
xor U4516 (N_4516,N_138,N_1292);
nor U4517 (N_4517,N_1688,N_1141);
or U4518 (N_4518,N_2223,N_185);
or U4519 (N_4519,N_641,N_1016);
and U4520 (N_4520,N_1657,N_1178);
xnor U4521 (N_4521,N_469,N_385);
nand U4522 (N_4522,N_128,N_769);
and U4523 (N_4523,N_737,N_1779);
nand U4524 (N_4524,N_1631,N_608);
nand U4525 (N_4525,N_1544,N_1244);
nand U4526 (N_4526,N_1406,N_1116);
nor U4527 (N_4527,N_2193,N_440);
or U4528 (N_4528,N_495,N_2392);
nor U4529 (N_4529,N_326,N_2);
and U4530 (N_4530,N_192,N_1076);
nand U4531 (N_4531,N_1632,N_288);
xnor U4532 (N_4532,N_32,N_1025);
nand U4533 (N_4533,N_1796,N_1883);
and U4534 (N_4534,N_1414,N_2183);
nor U4535 (N_4535,N_1531,N_1317);
xnor U4536 (N_4536,N_819,N_210);
xnor U4537 (N_4537,N_248,N_936);
nor U4538 (N_4538,N_1955,N_2102);
nor U4539 (N_4539,N_808,N_689);
nand U4540 (N_4540,N_1059,N_769);
or U4541 (N_4541,N_1532,N_159);
nand U4542 (N_4542,N_872,N_1315);
nor U4543 (N_4543,N_693,N_2299);
xnor U4544 (N_4544,N_721,N_966);
and U4545 (N_4545,N_549,N_420);
or U4546 (N_4546,N_2399,N_468);
and U4547 (N_4547,N_1804,N_2324);
and U4548 (N_4548,N_396,N_113);
nand U4549 (N_4549,N_2147,N_346);
or U4550 (N_4550,N_1343,N_799);
or U4551 (N_4551,N_1866,N_514);
xnor U4552 (N_4552,N_2376,N_999);
and U4553 (N_4553,N_1707,N_17);
nor U4554 (N_4554,N_774,N_1690);
or U4555 (N_4555,N_790,N_2391);
xor U4556 (N_4556,N_640,N_2120);
and U4557 (N_4557,N_2023,N_2032);
nor U4558 (N_4558,N_1483,N_1992);
and U4559 (N_4559,N_415,N_2124);
xnor U4560 (N_4560,N_1738,N_160);
nor U4561 (N_4561,N_494,N_879);
xnor U4562 (N_4562,N_981,N_1350);
nor U4563 (N_4563,N_2292,N_794);
nor U4564 (N_4564,N_450,N_1701);
nor U4565 (N_4565,N_801,N_1332);
or U4566 (N_4566,N_412,N_1918);
nor U4567 (N_4567,N_1003,N_2210);
or U4568 (N_4568,N_355,N_1578);
or U4569 (N_4569,N_438,N_194);
and U4570 (N_4570,N_2294,N_1233);
nor U4571 (N_4571,N_1572,N_801);
and U4572 (N_4572,N_600,N_1220);
xnor U4573 (N_4573,N_1961,N_1916);
and U4574 (N_4574,N_1044,N_2358);
nor U4575 (N_4575,N_1412,N_1884);
xor U4576 (N_4576,N_1001,N_369);
nor U4577 (N_4577,N_2058,N_1663);
and U4578 (N_4578,N_997,N_1177);
nand U4579 (N_4579,N_2164,N_2223);
nand U4580 (N_4580,N_923,N_1283);
and U4581 (N_4581,N_502,N_786);
or U4582 (N_4582,N_2313,N_2229);
nor U4583 (N_4583,N_1009,N_747);
nand U4584 (N_4584,N_640,N_768);
or U4585 (N_4585,N_2287,N_959);
nor U4586 (N_4586,N_2216,N_1543);
nor U4587 (N_4587,N_1006,N_632);
and U4588 (N_4588,N_66,N_1659);
nand U4589 (N_4589,N_1910,N_2342);
and U4590 (N_4590,N_1350,N_2194);
nor U4591 (N_4591,N_207,N_646);
and U4592 (N_4592,N_397,N_1034);
nor U4593 (N_4593,N_33,N_2243);
nor U4594 (N_4594,N_354,N_748);
xor U4595 (N_4595,N_1199,N_2028);
or U4596 (N_4596,N_477,N_1576);
and U4597 (N_4597,N_805,N_419);
or U4598 (N_4598,N_1386,N_2233);
or U4599 (N_4599,N_1801,N_459);
nand U4600 (N_4600,N_718,N_1123);
nor U4601 (N_4601,N_2142,N_1284);
and U4602 (N_4602,N_1438,N_1924);
or U4603 (N_4603,N_362,N_395);
nor U4604 (N_4604,N_853,N_555);
nor U4605 (N_4605,N_2307,N_2344);
or U4606 (N_4606,N_294,N_890);
and U4607 (N_4607,N_392,N_1970);
nor U4608 (N_4608,N_2339,N_1393);
nand U4609 (N_4609,N_1326,N_2474);
or U4610 (N_4610,N_1358,N_362);
and U4611 (N_4611,N_1294,N_1864);
nor U4612 (N_4612,N_2195,N_690);
or U4613 (N_4613,N_2202,N_1614);
or U4614 (N_4614,N_342,N_1709);
and U4615 (N_4615,N_1493,N_1946);
nand U4616 (N_4616,N_1107,N_1315);
nand U4617 (N_4617,N_2229,N_1742);
and U4618 (N_4618,N_2205,N_1151);
or U4619 (N_4619,N_1402,N_602);
xor U4620 (N_4620,N_181,N_184);
nor U4621 (N_4621,N_653,N_1950);
and U4622 (N_4622,N_1696,N_2280);
and U4623 (N_4623,N_867,N_1034);
and U4624 (N_4624,N_2348,N_1900);
nand U4625 (N_4625,N_275,N_1587);
and U4626 (N_4626,N_270,N_2188);
xor U4627 (N_4627,N_2093,N_125);
and U4628 (N_4628,N_2412,N_975);
and U4629 (N_4629,N_1092,N_2376);
or U4630 (N_4630,N_2097,N_1617);
and U4631 (N_4631,N_600,N_1081);
nand U4632 (N_4632,N_1000,N_1941);
nand U4633 (N_4633,N_374,N_2331);
nor U4634 (N_4634,N_2034,N_1299);
and U4635 (N_4635,N_846,N_2150);
or U4636 (N_4636,N_2020,N_1730);
and U4637 (N_4637,N_1305,N_741);
and U4638 (N_4638,N_1042,N_604);
nor U4639 (N_4639,N_2487,N_373);
nand U4640 (N_4640,N_2207,N_1172);
nor U4641 (N_4641,N_2496,N_1063);
and U4642 (N_4642,N_2181,N_2296);
nand U4643 (N_4643,N_1975,N_2347);
nor U4644 (N_4644,N_1577,N_1388);
or U4645 (N_4645,N_2384,N_2024);
or U4646 (N_4646,N_793,N_1894);
or U4647 (N_4647,N_41,N_1404);
nor U4648 (N_4648,N_942,N_2353);
xnor U4649 (N_4649,N_443,N_1368);
xnor U4650 (N_4650,N_591,N_1296);
nand U4651 (N_4651,N_698,N_2234);
and U4652 (N_4652,N_52,N_1823);
nand U4653 (N_4653,N_1283,N_1278);
nand U4654 (N_4654,N_1836,N_179);
nor U4655 (N_4655,N_1588,N_207);
nand U4656 (N_4656,N_2034,N_110);
and U4657 (N_4657,N_1067,N_344);
or U4658 (N_4658,N_1473,N_1732);
or U4659 (N_4659,N_206,N_2068);
nor U4660 (N_4660,N_1516,N_1030);
nor U4661 (N_4661,N_1228,N_2280);
nand U4662 (N_4662,N_2491,N_10);
nor U4663 (N_4663,N_907,N_1164);
and U4664 (N_4664,N_2163,N_2183);
nand U4665 (N_4665,N_1869,N_618);
nor U4666 (N_4666,N_1163,N_260);
xor U4667 (N_4667,N_929,N_2257);
nor U4668 (N_4668,N_2210,N_798);
or U4669 (N_4669,N_22,N_530);
or U4670 (N_4670,N_2410,N_1010);
nand U4671 (N_4671,N_160,N_273);
nor U4672 (N_4672,N_980,N_251);
nand U4673 (N_4673,N_275,N_1522);
or U4674 (N_4674,N_2037,N_1744);
nor U4675 (N_4675,N_2009,N_450);
and U4676 (N_4676,N_1179,N_423);
or U4677 (N_4677,N_996,N_625);
nand U4678 (N_4678,N_915,N_2155);
or U4679 (N_4679,N_1827,N_857);
or U4680 (N_4680,N_1250,N_456);
or U4681 (N_4681,N_293,N_1551);
nand U4682 (N_4682,N_1303,N_605);
nand U4683 (N_4683,N_2192,N_1356);
and U4684 (N_4684,N_410,N_123);
nor U4685 (N_4685,N_1416,N_29);
or U4686 (N_4686,N_1327,N_334);
and U4687 (N_4687,N_1138,N_881);
xnor U4688 (N_4688,N_1813,N_1568);
nand U4689 (N_4689,N_161,N_832);
nand U4690 (N_4690,N_568,N_188);
nor U4691 (N_4691,N_2142,N_592);
nand U4692 (N_4692,N_2314,N_236);
and U4693 (N_4693,N_1552,N_2468);
xnor U4694 (N_4694,N_23,N_138);
xnor U4695 (N_4695,N_1598,N_2184);
or U4696 (N_4696,N_1088,N_1433);
and U4697 (N_4697,N_1104,N_815);
nor U4698 (N_4698,N_1104,N_2471);
or U4699 (N_4699,N_518,N_854);
nand U4700 (N_4700,N_283,N_2450);
and U4701 (N_4701,N_2194,N_264);
or U4702 (N_4702,N_1154,N_1920);
xor U4703 (N_4703,N_13,N_1222);
nor U4704 (N_4704,N_2399,N_1861);
nor U4705 (N_4705,N_1897,N_1064);
and U4706 (N_4706,N_1748,N_1542);
nor U4707 (N_4707,N_695,N_1689);
or U4708 (N_4708,N_1364,N_822);
or U4709 (N_4709,N_585,N_1694);
nand U4710 (N_4710,N_1269,N_31);
nor U4711 (N_4711,N_719,N_127);
or U4712 (N_4712,N_1380,N_2265);
nand U4713 (N_4713,N_1372,N_2476);
and U4714 (N_4714,N_2240,N_1086);
or U4715 (N_4715,N_236,N_1024);
nor U4716 (N_4716,N_1927,N_1500);
and U4717 (N_4717,N_188,N_1950);
nor U4718 (N_4718,N_48,N_2421);
xor U4719 (N_4719,N_1683,N_1903);
and U4720 (N_4720,N_2388,N_1028);
or U4721 (N_4721,N_539,N_1696);
and U4722 (N_4722,N_1268,N_927);
xnor U4723 (N_4723,N_1276,N_557);
nand U4724 (N_4724,N_1576,N_2375);
nor U4725 (N_4725,N_1913,N_723);
or U4726 (N_4726,N_2235,N_328);
nand U4727 (N_4727,N_1206,N_2464);
or U4728 (N_4728,N_249,N_600);
nand U4729 (N_4729,N_1169,N_529);
and U4730 (N_4730,N_1968,N_1641);
nand U4731 (N_4731,N_1339,N_1108);
nand U4732 (N_4732,N_2332,N_446);
nor U4733 (N_4733,N_1348,N_2045);
and U4734 (N_4734,N_1383,N_2341);
nand U4735 (N_4735,N_503,N_585);
nand U4736 (N_4736,N_1987,N_1848);
or U4737 (N_4737,N_348,N_1274);
or U4738 (N_4738,N_579,N_2324);
or U4739 (N_4739,N_1746,N_840);
xnor U4740 (N_4740,N_2137,N_2219);
and U4741 (N_4741,N_1329,N_830);
xnor U4742 (N_4742,N_1746,N_528);
nor U4743 (N_4743,N_1333,N_1161);
nand U4744 (N_4744,N_1454,N_664);
and U4745 (N_4745,N_2301,N_2135);
or U4746 (N_4746,N_704,N_1854);
and U4747 (N_4747,N_1475,N_528);
and U4748 (N_4748,N_687,N_950);
and U4749 (N_4749,N_2412,N_692);
or U4750 (N_4750,N_1806,N_972);
nor U4751 (N_4751,N_166,N_2341);
nor U4752 (N_4752,N_1443,N_164);
nand U4753 (N_4753,N_1437,N_280);
nand U4754 (N_4754,N_1603,N_280);
and U4755 (N_4755,N_1832,N_540);
and U4756 (N_4756,N_1532,N_1337);
or U4757 (N_4757,N_993,N_2452);
or U4758 (N_4758,N_470,N_2016);
nor U4759 (N_4759,N_93,N_1066);
nand U4760 (N_4760,N_1872,N_1807);
or U4761 (N_4761,N_1336,N_2381);
or U4762 (N_4762,N_1612,N_172);
and U4763 (N_4763,N_975,N_2430);
nand U4764 (N_4764,N_2156,N_1916);
nand U4765 (N_4765,N_442,N_2360);
nand U4766 (N_4766,N_680,N_1720);
and U4767 (N_4767,N_1649,N_1416);
and U4768 (N_4768,N_1380,N_2379);
or U4769 (N_4769,N_1085,N_1509);
and U4770 (N_4770,N_1866,N_1947);
xnor U4771 (N_4771,N_1770,N_2405);
or U4772 (N_4772,N_1731,N_1862);
nor U4773 (N_4773,N_1760,N_98);
and U4774 (N_4774,N_142,N_1592);
nand U4775 (N_4775,N_473,N_866);
or U4776 (N_4776,N_2018,N_149);
or U4777 (N_4777,N_93,N_1266);
nor U4778 (N_4778,N_2025,N_1499);
and U4779 (N_4779,N_1171,N_2125);
xnor U4780 (N_4780,N_60,N_1398);
or U4781 (N_4781,N_1477,N_1861);
and U4782 (N_4782,N_1668,N_134);
nand U4783 (N_4783,N_2333,N_575);
or U4784 (N_4784,N_1088,N_2198);
nor U4785 (N_4785,N_1093,N_231);
nand U4786 (N_4786,N_1061,N_477);
or U4787 (N_4787,N_1447,N_2000);
nor U4788 (N_4788,N_2425,N_1263);
xor U4789 (N_4789,N_131,N_94);
or U4790 (N_4790,N_1310,N_633);
xnor U4791 (N_4791,N_255,N_1045);
nand U4792 (N_4792,N_2044,N_2105);
or U4793 (N_4793,N_921,N_2374);
nor U4794 (N_4794,N_1813,N_968);
and U4795 (N_4795,N_2124,N_1272);
or U4796 (N_4796,N_866,N_177);
nand U4797 (N_4797,N_706,N_2405);
and U4798 (N_4798,N_2391,N_2382);
nor U4799 (N_4799,N_1172,N_1297);
nor U4800 (N_4800,N_102,N_781);
or U4801 (N_4801,N_947,N_1622);
or U4802 (N_4802,N_809,N_2295);
xnor U4803 (N_4803,N_190,N_786);
and U4804 (N_4804,N_1236,N_232);
or U4805 (N_4805,N_2488,N_1285);
and U4806 (N_4806,N_1394,N_352);
xor U4807 (N_4807,N_936,N_2299);
xor U4808 (N_4808,N_2375,N_781);
nand U4809 (N_4809,N_2149,N_2092);
nor U4810 (N_4810,N_2129,N_521);
xor U4811 (N_4811,N_423,N_1283);
or U4812 (N_4812,N_106,N_879);
nor U4813 (N_4813,N_174,N_739);
or U4814 (N_4814,N_1818,N_197);
or U4815 (N_4815,N_1765,N_1741);
nor U4816 (N_4816,N_1941,N_472);
nand U4817 (N_4817,N_2462,N_1391);
nor U4818 (N_4818,N_2416,N_1356);
nand U4819 (N_4819,N_673,N_199);
nor U4820 (N_4820,N_1975,N_275);
nor U4821 (N_4821,N_2230,N_1374);
nor U4822 (N_4822,N_1470,N_1001);
or U4823 (N_4823,N_174,N_424);
and U4824 (N_4824,N_219,N_2018);
nor U4825 (N_4825,N_989,N_105);
xor U4826 (N_4826,N_1517,N_1178);
xnor U4827 (N_4827,N_852,N_538);
nand U4828 (N_4828,N_1154,N_28);
nor U4829 (N_4829,N_513,N_1450);
and U4830 (N_4830,N_766,N_1792);
nor U4831 (N_4831,N_1317,N_1937);
nand U4832 (N_4832,N_1339,N_2273);
nand U4833 (N_4833,N_1016,N_1827);
or U4834 (N_4834,N_231,N_327);
nor U4835 (N_4835,N_742,N_1998);
nor U4836 (N_4836,N_2336,N_113);
nor U4837 (N_4837,N_2030,N_1896);
and U4838 (N_4838,N_1878,N_30);
or U4839 (N_4839,N_336,N_1624);
nand U4840 (N_4840,N_2259,N_774);
and U4841 (N_4841,N_1993,N_1415);
nor U4842 (N_4842,N_1100,N_58);
xnor U4843 (N_4843,N_1754,N_237);
or U4844 (N_4844,N_1858,N_569);
nand U4845 (N_4845,N_1555,N_1920);
and U4846 (N_4846,N_1922,N_1776);
or U4847 (N_4847,N_202,N_2165);
or U4848 (N_4848,N_1700,N_1217);
or U4849 (N_4849,N_2223,N_757);
or U4850 (N_4850,N_1441,N_923);
nand U4851 (N_4851,N_1626,N_1114);
and U4852 (N_4852,N_1842,N_197);
and U4853 (N_4853,N_1000,N_2007);
or U4854 (N_4854,N_2071,N_542);
nor U4855 (N_4855,N_1430,N_581);
nor U4856 (N_4856,N_2074,N_1393);
nand U4857 (N_4857,N_764,N_2454);
and U4858 (N_4858,N_221,N_2099);
xor U4859 (N_4859,N_977,N_2073);
or U4860 (N_4860,N_771,N_2313);
xnor U4861 (N_4861,N_185,N_1184);
or U4862 (N_4862,N_636,N_1321);
nor U4863 (N_4863,N_1357,N_1317);
and U4864 (N_4864,N_145,N_2486);
nand U4865 (N_4865,N_2232,N_1028);
or U4866 (N_4866,N_1968,N_603);
or U4867 (N_4867,N_806,N_1637);
and U4868 (N_4868,N_37,N_2224);
xor U4869 (N_4869,N_1980,N_1491);
or U4870 (N_4870,N_34,N_664);
or U4871 (N_4871,N_2412,N_1875);
xor U4872 (N_4872,N_892,N_1219);
or U4873 (N_4873,N_828,N_1267);
or U4874 (N_4874,N_457,N_710);
nand U4875 (N_4875,N_1033,N_810);
or U4876 (N_4876,N_2397,N_1718);
nor U4877 (N_4877,N_2327,N_869);
nand U4878 (N_4878,N_1671,N_1404);
nand U4879 (N_4879,N_1020,N_1280);
and U4880 (N_4880,N_1958,N_2085);
nor U4881 (N_4881,N_595,N_1217);
nand U4882 (N_4882,N_292,N_228);
and U4883 (N_4883,N_1685,N_1558);
and U4884 (N_4884,N_2452,N_266);
nor U4885 (N_4885,N_453,N_564);
nor U4886 (N_4886,N_392,N_190);
or U4887 (N_4887,N_1156,N_88);
nand U4888 (N_4888,N_2299,N_1444);
nand U4889 (N_4889,N_1277,N_1947);
nand U4890 (N_4890,N_1395,N_2269);
and U4891 (N_4891,N_2110,N_1483);
nand U4892 (N_4892,N_1349,N_2196);
or U4893 (N_4893,N_864,N_533);
and U4894 (N_4894,N_2451,N_1474);
and U4895 (N_4895,N_191,N_1557);
nand U4896 (N_4896,N_638,N_403);
or U4897 (N_4897,N_1876,N_748);
and U4898 (N_4898,N_48,N_1551);
or U4899 (N_4899,N_276,N_2324);
or U4900 (N_4900,N_432,N_1593);
and U4901 (N_4901,N_1281,N_1103);
nand U4902 (N_4902,N_2332,N_595);
or U4903 (N_4903,N_2329,N_1211);
or U4904 (N_4904,N_1881,N_1073);
or U4905 (N_4905,N_1819,N_35);
and U4906 (N_4906,N_1264,N_1000);
nand U4907 (N_4907,N_116,N_859);
and U4908 (N_4908,N_484,N_1401);
nand U4909 (N_4909,N_1305,N_484);
nand U4910 (N_4910,N_184,N_1372);
and U4911 (N_4911,N_22,N_1402);
nand U4912 (N_4912,N_595,N_2193);
nand U4913 (N_4913,N_1799,N_2259);
nand U4914 (N_4914,N_2166,N_525);
xor U4915 (N_4915,N_1999,N_415);
nand U4916 (N_4916,N_1469,N_1553);
nor U4917 (N_4917,N_2495,N_923);
xor U4918 (N_4918,N_563,N_1850);
nand U4919 (N_4919,N_1227,N_855);
nor U4920 (N_4920,N_282,N_923);
or U4921 (N_4921,N_792,N_403);
xnor U4922 (N_4922,N_257,N_101);
nand U4923 (N_4923,N_1807,N_1048);
or U4924 (N_4924,N_540,N_666);
xnor U4925 (N_4925,N_1264,N_2365);
and U4926 (N_4926,N_2127,N_2152);
nand U4927 (N_4927,N_69,N_549);
nor U4928 (N_4928,N_1628,N_894);
nand U4929 (N_4929,N_899,N_1330);
nor U4930 (N_4930,N_1144,N_187);
nand U4931 (N_4931,N_2434,N_2423);
nor U4932 (N_4932,N_2318,N_1044);
nand U4933 (N_4933,N_1476,N_1191);
xor U4934 (N_4934,N_407,N_746);
and U4935 (N_4935,N_2313,N_211);
nor U4936 (N_4936,N_1728,N_1260);
or U4937 (N_4937,N_1850,N_1011);
xor U4938 (N_4938,N_1666,N_527);
and U4939 (N_4939,N_1701,N_1340);
and U4940 (N_4940,N_888,N_854);
or U4941 (N_4941,N_1436,N_1269);
nand U4942 (N_4942,N_1875,N_339);
nor U4943 (N_4943,N_2188,N_507);
or U4944 (N_4944,N_2097,N_146);
nor U4945 (N_4945,N_590,N_1992);
and U4946 (N_4946,N_1004,N_1065);
or U4947 (N_4947,N_1287,N_1208);
or U4948 (N_4948,N_1365,N_2225);
and U4949 (N_4949,N_2021,N_919);
or U4950 (N_4950,N_515,N_1408);
nor U4951 (N_4951,N_227,N_1823);
nand U4952 (N_4952,N_1710,N_944);
nand U4953 (N_4953,N_1011,N_813);
nor U4954 (N_4954,N_57,N_492);
and U4955 (N_4955,N_1979,N_1827);
and U4956 (N_4956,N_219,N_118);
or U4957 (N_4957,N_2105,N_1213);
nor U4958 (N_4958,N_190,N_2270);
nor U4959 (N_4959,N_1564,N_1083);
nor U4960 (N_4960,N_1726,N_841);
nand U4961 (N_4961,N_837,N_1145);
and U4962 (N_4962,N_682,N_231);
nand U4963 (N_4963,N_493,N_875);
nor U4964 (N_4964,N_1879,N_1816);
nor U4965 (N_4965,N_975,N_1548);
or U4966 (N_4966,N_390,N_757);
or U4967 (N_4967,N_1134,N_421);
and U4968 (N_4968,N_427,N_1083);
nand U4969 (N_4969,N_2373,N_1088);
or U4970 (N_4970,N_838,N_25);
nor U4971 (N_4971,N_37,N_12);
and U4972 (N_4972,N_1791,N_1805);
or U4973 (N_4973,N_2204,N_1785);
nor U4974 (N_4974,N_1755,N_1524);
nand U4975 (N_4975,N_510,N_322);
nor U4976 (N_4976,N_2256,N_99);
or U4977 (N_4977,N_2475,N_430);
or U4978 (N_4978,N_1337,N_1200);
nand U4979 (N_4979,N_716,N_2220);
nand U4980 (N_4980,N_1450,N_1462);
and U4981 (N_4981,N_2358,N_688);
xnor U4982 (N_4982,N_2210,N_521);
nor U4983 (N_4983,N_396,N_477);
nand U4984 (N_4984,N_563,N_812);
nand U4985 (N_4985,N_965,N_34);
nand U4986 (N_4986,N_1915,N_678);
nor U4987 (N_4987,N_394,N_95);
and U4988 (N_4988,N_971,N_408);
nand U4989 (N_4989,N_66,N_2491);
and U4990 (N_4990,N_1939,N_1501);
and U4991 (N_4991,N_394,N_1052);
nor U4992 (N_4992,N_1592,N_2381);
and U4993 (N_4993,N_1679,N_378);
nand U4994 (N_4994,N_966,N_514);
and U4995 (N_4995,N_2389,N_2180);
and U4996 (N_4996,N_2162,N_1587);
xor U4997 (N_4997,N_585,N_1684);
and U4998 (N_4998,N_161,N_116);
nand U4999 (N_4999,N_1172,N_1272);
nor UO_0 (O_0,N_4987,N_4884);
or UO_1 (O_1,N_4459,N_2955);
nor UO_2 (O_2,N_4359,N_4949);
nor UO_3 (O_3,N_3882,N_2767);
and UO_4 (O_4,N_3319,N_2817);
nor UO_5 (O_5,N_2602,N_2997);
and UO_6 (O_6,N_3215,N_2599);
or UO_7 (O_7,N_4261,N_2890);
or UO_8 (O_8,N_3203,N_4814);
nand UO_9 (O_9,N_4378,N_3901);
xnor UO_10 (O_10,N_4207,N_3050);
or UO_11 (O_11,N_4431,N_3204);
nand UO_12 (O_12,N_3114,N_3077);
and UO_13 (O_13,N_4199,N_3783);
or UO_14 (O_14,N_3130,N_4153);
nand UO_15 (O_15,N_2972,N_2707);
or UO_16 (O_16,N_3886,N_4248);
or UO_17 (O_17,N_3307,N_4766);
nor UO_18 (O_18,N_4666,N_2549);
xnor UO_19 (O_19,N_3533,N_4686);
nand UO_20 (O_20,N_2926,N_3980);
nand UO_21 (O_21,N_3161,N_3326);
nor UO_22 (O_22,N_4923,N_3429);
and UO_23 (O_23,N_2823,N_4721);
or UO_24 (O_24,N_2537,N_4942);
or UO_25 (O_25,N_3676,N_4833);
and UO_26 (O_26,N_4781,N_3795);
xnor UO_27 (O_27,N_3611,N_3191);
nand UO_28 (O_28,N_3895,N_3745);
and UO_29 (O_29,N_4219,N_4075);
or UO_30 (O_30,N_3433,N_4893);
xor UO_31 (O_31,N_3428,N_4438);
nand UO_32 (O_32,N_2527,N_3826);
xnor UO_33 (O_33,N_2722,N_4928);
and UO_34 (O_34,N_3877,N_4735);
xnor UO_35 (O_35,N_3684,N_3274);
nand UO_36 (O_36,N_4520,N_3504);
nor UO_37 (O_37,N_2561,N_3472);
or UO_38 (O_38,N_3380,N_4450);
nor UO_39 (O_39,N_4346,N_3487);
nor UO_40 (O_40,N_3675,N_4618);
or UO_41 (O_41,N_2999,N_4357);
and UO_42 (O_42,N_3657,N_2851);
nor UO_43 (O_43,N_4304,N_3146);
or UO_44 (O_44,N_4279,N_3444);
nand UO_45 (O_45,N_4491,N_2848);
nor UO_46 (O_46,N_4670,N_3060);
and UO_47 (O_47,N_3621,N_4345);
or UO_48 (O_48,N_2740,N_3774);
xor UO_49 (O_49,N_2614,N_4550);
or UO_50 (O_50,N_4541,N_4672);
or UO_51 (O_51,N_2837,N_4715);
or UO_52 (O_52,N_2522,N_2719);
xnor UO_53 (O_53,N_3042,N_4478);
nor UO_54 (O_54,N_2866,N_3085);
nor UO_55 (O_55,N_2758,N_4999);
nor UO_56 (O_56,N_4141,N_3296);
and UO_57 (O_57,N_4512,N_4325);
nor UO_58 (O_58,N_4247,N_2966);
or UO_59 (O_59,N_3206,N_3521);
nor UO_60 (O_60,N_2664,N_4239);
and UO_61 (O_61,N_3766,N_4429);
nor UO_62 (O_62,N_4201,N_3391);
or UO_63 (O_63,N_4561,N_3368);
and UO_64 (O_64,N_4591,N_3421);
nand UO_65 (O_65,N_3308,N_2535);
nand UO_66 (O_66,N_3565,N_3771);
xor UO_67 (O_67,N_2515,N_3789);
nand UO_68 (O_68,N_4916,N_3515);
nor UO_69 (O_69,N_4064,N_4962);
nor UO_70 (O_70,N_4619,N_3126);
or UO_71 (O_71,N_4640,N_3821);
nand UO_72 (O_72,N_3379,N_2985);
or UO_73 (O_73,N_3259,N_3960);
and UO_74 (O_74,N_3696,N_4677);
nand UO_75 (O_75,N_4125,N_2525);
nor UO_76 (O_76,N_3412,N_2981);
nor UO_77 (O_77,N_2828,N_3854);
nor UO_78 (O_78,N_2834,N_4213);
or UO_79 (O_79,N_3999,N_4961);
or UO_80 (O_80,N_4722,N_4960);
nor UO_81 (O_81,N_3543,N_2869);
xnor UO_82 (O_82,N_2547,N_3589);
and UO_83 (O_83,N_2856,N_2951);
nor UO_84 (O_84,N_2944,N_4265);
and UO_85 (O_85,N_3568,N_4204);
nand UO_86 (O_86,N_4675,N_3422);
xnor UO_87 (O_87,N_4787,N_2729);
nand UO_88 (O_88,N_4117,N_3407);
nor UO_89 (O_89,N_2544,N_3051);
nor UO_90 (O_90,N_3301,N_2717);
xnor UO_91 (O_91,N_4854,N_2503);
xor UO_92 (O_92,N_2609,N_3942);
nand UO_93 (O_93,N_2538,N_4245);
and UO_94 (O_94,N_3133,N_3718);
xor UO_95 (O_95,N_3748,N_4855);
and UO_96 (O_96,N_4567,N_2936);
nor UO_97 (O_97,N_2831,N_3058);
nand UO_98 (O_98,N_3460,N_3572);
or UO_99 (O_99,N_2775,N_4161);
or UO_100 (O_100,N_4695,N_4985);
or UO_101 (O_101,N_2770,N_4602);
nor UO_102 (O_102,N_3833,N_3554);
or UO_103 (O_103,N_2718,N_4094);
or UO_104 (O_104,N_4114,N_2780);
nand UO_105 (O_105,N_4100,N_2556);
or UO_106 (O_106,N_4654,N_4548);
and UO_107 (O_107,N_2501,N_2911);
or UO_108 (O_108,N_3386,N_4362);
or UO_109 (O_109,N_4636,N_4964);
or UO_110 (O_110,N_3569,N_2716);
nand UO_111 (O_111,N_3922,N_4321);
xnor UO_112 (O_112,N_2839,N_4790);
and UO_113 (O_113,N_3755,N_4108);
nand UO_114 (O_114,N_3234,N_2968);
or UO_115 (O_115,N_4414,N_3029);
or UO_116 (O_116,N_4629,N_4701);
and UO_117 (O_117,N_3909,N_4214);
and UO_118 (O_118,N_4372,N_4185);
and UO_119 (O_119,N_3329,N_4457);
and UO_120 (O_120,N_4797,N_3358);
and UO_121 (O_121,N_3513,N_2858);
and UO_122 (O_122,N_3687,N_4991);
nor UO_123 (O_123,N_4041,N_2975);
and UO_124 (O_124,N_4564,N_4390);
nand UO_125 (O_125,N_3807,N_3182);
and UO_126 (O_126,N_3443,N_3908);
and UO_127 (O_127,N_4129,N_3176);
and UO_128 (O_128,N_3004,N_4407);
xor UO_129 (O_129,N_4224,N_3483);
nor UO_130 (O_130,N_4824,N_3136);
nand UO_131 (O_131,N_3527,N_3957);
or UO_132 (O_132,N_4235,N_4503);
and UO_133 (O_133,N_3944,N_4980);
and UO_134 (O_134,N_3476,N_3725);
nor UO_135 (O_135,N_2563,N_4626);
or UO_136 (O_136,N_4656,N_3705);
xnor UO_137 (O_137,N_2578,N_3678);
and UO_138 (O_138,N_4389,N_2743);
and UO_139 (O_139,N_4699,N_2863);
or UO_140 (O_140,N_3929,N_3275);
nor UO_141 (O_141,N_4354,N_2957);
and UO_142 (O_142,N_3546,N_3813);
or UO_143 (O_143,N_4298,N_4397);
nor UO_144 (O_144,N_4333,N_2794);
nor UO_145 (O_145,N_3926,N_4641);
or UO_146 (O_146,N_3323,N_4542);
nand UO_147 (O_147,N_4463,N_3614);
or UO_148 (O_148,N_3816,N_3059);
nand UO_149 (O_149,N_3376,N_4183);
nand UO_150 (O_150,N_4169,N_2663);
and UO_151 (O_151,N_2841,N_3896);
nand UO_152 (O_152,N_4003,N_4565);
and UO_153 (O_153,N_3081,N_3517);
or UO_154 (O_154,N_2779,N_4394);
or UO_155 (O_155,N_3852,N_3257);
nand UO_156 (O_156,N_2730,N_3891);
or UO_157 (O_157,N_2827,N_2932);
xor UO_158 (O_158,N_3266,N_4085);
nand UO_159 (O_159,N_4012,N_2785);
or UO_160 (O_160,N_4922,N_4237);
xnor UO_161 (O_161,N_3034,N_3145);
nor UO_162 (O_162,N_3302,N_3289);
nand UO_163 (O_163,N_2523,N_2983);
or UO_164 (O_164,N_3342,N_3017);
nor UO_165 (O_165,N_2674,N_4662);
or UO_166 (O_166,N_4761,N_2577);
and UO_167 (O_167,N_3961,N_4612);
xnor UO_168 (O_168,N_3337,N_2753);
or UO_169 (O_169,N_2878,N_4732);
and UO_170 (O_170,N_4352,N_3183);
nor UO_171 (O_171,N_4948,N_4793);
xor UO_172 (O_172,N_4274,N_4415);
or UO_173 (O_173,N_2789,N_3121);
nand UO_174 (O_174,N_4587,N_4726);
xnor UO_175 (O_175,N_4908,N_3967);
nand UO_176 (O_176,N_2896,N_2720);
nor UO_177 (O_177,N_3388,N_4804);
nand UO_178 (O_178,N_4025,N_4455);
or UO_179 (O_179,N_3168,N_4330);
and UO_180 (O_180,N_3871,N_3876);
and UO_181 (O_181,N_2888,N_3742);
nor UO_182 (O_182,N_4770,N_2875);
nand UO_183 (O_183,N_2843,N_4057);
or UO_184 (O_184,N_3954,N_4750);
or UO_185 (O_185,N_3112,N_4039);
or UO_186 (O_186,N_3759,N_2939);
or UO_187 (O_187,N_4166,N_3155);
xor UO_188 (O_188,N_3064,N_3951);
nand UO_189 (O_189,N_3471,N_2784);
nand UO_190 (O_190,N_4831,N_3462);
xor UO_191 (O_191,N_4549,N_3398);
xnor UO_192 (O_192,N_2853,N_2608);
and UO_193 (O_193,N_3806,N_3560);
nand UO_194 (O_194,N_3500,N_4327);
nor UO_195 (O_195,N_4303,N_4951);
nor UO_196 (O_196,N_4035,N_2555);
or UO_197 (O_197,N_3461,N_2887);
nor UO_198 (O_198,N_2598,N_4023);
and UO_199 (O_199,N_4427,N_3710);
and UO_200 (O_200,N_2978,N_4538);
and UO_201 (O_201,N_4788,N_4016);
and UO_202 (O_202,N_4492,N_4152);
nor UO_203 (O_203,N_3322,N_4243);
and UO_204 (O_204,N_4163,N_4707);
or UO_205 (O_205,N_4689,N_4425);
or UO_206 (O_206,N_2621,N_3227);
nand UO_207 (O_207,N_2971,N_3309);
and UO_208 (O_208,N_3767,N_3211);
nand UO_209 (O_209,N_4685,N_3445);
and UO_210 (O_210,N_3733,N_4206);
nor UO_211 (O_211,N_2529,N_2586);
or UO_212 (O_212,N_4608,N_2667);
xnor UO_213 (O_213,N_2914,N_3820);
or UO_214 (O_214,N_4338,N_3067);
xnor UO_215 (O_215,N_2745,N_3150);
xnor UO_216 (O_216,N_3866,N_3496);
nand UO_217 (O_217,N_4127,N_3522);
and UO_218 (O_218,N_3184,N_3958);
nand UO_219 (O_219,N_4234,N_2994);
xor UO_220 (O_220,N_2798,N_4919);
or UO_221 (O_221,N_2656,N_3545);
and UO_222 (O_222,N_4424,N_2710);
and UO_223 (O_223,N_4877,N_4339);
nand UO_224 (O_224,N_3963,N_3073);
or UO_225 (O_225,N_3514,N_3343);
nor UO_226 (O_226,N_3099,N_3520);
nor UO_227 (O_227,N_3361,N_3535);
nand UO_228 (O_228,N_4506,N_2581);
nor UO_229 (O_229,N_2733,N_2696);
xor UO_230 (O_230,N_3237,N_3108);
xnor UO_231 (O_231,N_4349,N_4162);
nor UO_232 (O_232,N_3180,N_4875);
nand UO_233 (O_233,N_4773,N_3950);
or UO_234 (O_234,N_3297,N_3363);
xnor UO_235 (O_235,N_4746,N_3768);
and UO_236 (O_236,N_3594,N_4251);
or UO_237 (O_237,N_3452,N_4719);
and UO_238 (O_238,N_2879,N_2783);
nor UO_239 (O_239,N_2712,N_4124);
and UO_240 (O_240,N_3086,N_4539);
nand UO_241 (O_241,N_3586,N_4486);
nand UO_242 (O_242,N_4441,N_3238);
nor UO_243 (O_243,N_4954,N_3832);
and UO_244 (O_244,N_3626,N_3187);
or UO_245 (O_245,N_2654,N_2850);
and UO_246 (O_246,N_3276,N_2993);
nand UO_247 (O_247,N_3135,N_4903);
nand UO_248 (O_248,N_2631,N_4444);
xnor UO_249 (O_249,N_2830,N_3819);
or UO_250 (O_250,N_4009,N_2736);
and UO_251 (O_251,N_3392,N_4742);
or UO_252 (O_252,N_2605,N_3062);
nand UO_253 (O_253,N_4795,N_2870);
and UO_254 (O_254,N_4568,N_3162);
nand UO_255 (O_255,N_4927,N_4028);
xnor UO_256 (O_256,N_2516,N_3378);
nand UO_257 (O_257,N_3691,N_4386);
or UO_258 (O_258,N_2781,N_4032);
or UO_259 (O_259,N_3579,N_3466);
or UO_260 (O_260,N_2532,N_4800);
nor UO_261 (O_261,N_3292,N_4493);
and UO_262 (O_262,N_4399,N_2747);
nor UO_263 (O_263,N_3377,N_2897);
xnor UO_264 (O_264,N_4652,N_2610);
nand UO_265 (O_265,N_3897,N_2772);
xnor UO_266 (O_266,N_3870,N_3602);
nand UO_267 (O_267,N_3955,N_3526);
nand UO_268 (O_268,N_3446,N_3205);
and UO_269 (O_269,N_3419,N_3752);
or UO_270 (O_270,N_3101,N_3055);
or UO_271 (O_271,N_3116,N_2766);
and UO_272 (O_272,N_4202,N_4164);
or UO_273 (O_273,N_2512,N_4344);
and UO_274 (O_274,N_4484,N_3974);
and UO_275 (O_275,N_4458,N_3727);
nor UO_276 (O_276,N_2660,N_4521);
and UO_277 (O_277,N_4476,N_2818);
nand UO_278 (O_278,N_3716,N_2806);
nor UO_279 (O_279,N_2998,N_4902);
nand UO_280 (O_280,N_4921,N_4296);
or UO_281 (O_281,N_3334,N_4885);
nand UO_282 (O_282,N_3134,N_2676);
xnor UO_283 (O_283,N_2845,N_2995);
and UO_284 (O_284,N_3047,N_4005);
and UO_285 (O_285,N_4861,N_4208);
nor UO_286 (O_286,N_3953,N_3793);
or UO_287 (O_287,N_3822,N_4053);
and UO_288 (O_288,N_2825,N_3489);
or UO_289 (O_289,N_2731,N_2548);
nand UO_290 (O_290,N_3581,N_2690);
nor UO_291 (O_291,N_3470,N_3245);
or UO_292 (O_292,N_4178,N_4530);
nand UO_293 (O_293,N_4316,N_4465);
or UO_294 (O_294,N_4412,N_3260);
nand UO_295 (O_295,N_2821,N_4398);
nand UO_296 (O_296,N_4605,N_3420);
and UO_297 (O_297,N_2682,N_3615);
and UO_298 (O_298,N_4471,N_3485);
nand UO_299 (O_299,N_4528,N_2657);
and UO_300 (O_300,N_4437,N_3702);
or UO_301 (O_301,N_4751,N_3438);
nor UO_302 (O_302,N_2751,N_4416);
or UO_303 (O_303,N_2816,N_2533);
or UO_304 (O_304,N_4655,N_3490);
nand UO_305 (O_305,N_2637,N_3415);
or UO_306 (O_306,N_3879,N_3936);
and UO_307 (O_307,N_3223,N_4332);
xnor UO_308 (O_308,N_3328,N_4446);
xor UO_309 (O_309,N_4289,N_3503);
or UO_310 (O_310,N_3915,N_3624);
nor UO_311 (O_311,N_3537,N_4181);
nand UO_312 (O_312,N_4144,N_4260);
and UO_313 (O_313,N_4262,N_2634);
nand UO_314 (O_314,N_4037,N_3859);
xnor UO_315 (O_315,N_3549,N_3913);
and UO_316 (O_316,N_3582,N_3998);
nand UO_317 (O_317,N_3762,N_4452);
or UO_318 (O_318,N_2723,N_3288);
or UO_319 (O_319,N_4663,N_4001);
or UO_320 (O_320,N_3949,N_4519);
and UO_321 (O_321,N_3843,N_3207);
and UO_322 (O_322,N_3536,N_4950);
and UO_323 (O_323,N_4650,N_4290);
and UO_324 (O_324,N_3119,N_3616);
nor UO_325 (O_325,N_4047,N_3906);
or UO_326 (O_326,N_4341,N_4080);
or UO_327 (O_327,N_3904,N_3148);
nor UO_328 (O_328,N_4905,N_4050);
or UO_329 (O_329,N_4583,N_3542);
or UO_330 (O_330,N_3959,N_3287);
nor UO_331 (O_331,N_4996,N_3076);
nor UO_332 (O_332,N_4319,N_4355);
and UO_333 (O_333,N_2518,N_3068);
xnor UO_334 (O_334,N_4315,N_3894);
or UO_335 (O_335,N_3159,N_3341);
or UO_336 (O_336,N_2917,N_4292);
and UO_337 (O_337,N_2625,N_3414);
and UO_338 (O_338,N_4002,N_4653);
or UO_339 (O_339,N_3746,N_3262);
nand UO_340 (O_340,N_3124,N_2511);
nand UO_341 (O_341,N_2680,N_4229);
and UO_342 (O_342,N_4635,N_4522);
nor UO_343 (O_343,N_4445,N_3919);
or UO_344 (O_344,N_3734,N_2619);
xor UO_345 (O_345,N_4759,N_4678);
nand UO_346 (O_346,N_4944,N_3709);
or UO_347 (O_347,N_3141,N_2765);
or UO_348 (O_348,N_3338,N_4070);
nor UO_349 (O_349,N_3738,N_4240);
nor UO_350 (O_350,N_3865,N_3492);
and UO_351 (O_351,N_3930,N_4291);
and UO_352 (O_352,N_4588,N_3088);
nor UO_353 (O_353,N_2615,N_4659);
nor UO_354 (O_354,N_4418,N_4620);
xnor UO_355 (O_355,N_4259,N_4963);
or UO_356 (O_356,N_3848,N_3584);
xor UO_357 (O_357,N_3860,N_2923);
or UO_358 (O_358,N_2778,N_4617);
nor UO_359 (O_359,N_4495,N_4180);
nand UO_360 (O_360,N_2611,N_4451);
or UO_361 (O_361,N_3962,N_4624);
nor UO_362 (O_362,N_2540,N_3592);
and UO_363 (O_363,N_2916,N_4713);
xor UO_364 (O_364,N_3688,N_3846);
or UO_365 (O_365,N_3610,N_4829);
nor UO_366 (O_366,N_4776,N_2886);
nand UO_367 (O_367,N_4560,N_4524);
or UO_368 (O_368,N_2692,N_4361);
nor UO_369 (O_369,N_4832,N_3005);
nand UO_370 (O_370,N_4615,N_3189);
nand UO_371 (O_371,N_2881,N_4584);
or UO_372 (O_372,N_3811,N_4209);
nor UO_373 (O_373,N_4377,N_3563);
or UO_374 (O_374,N_4040,N_4842);
and UO_375 (O_375,N_3792,N_4036);
nand UO_376 (O_376,N_4850,N_4013);
nand UO_377 (O_377,N_3606,N_3916);
nand UO_378 (O_378,N_4148,N_2946);
nor UO_379 (O_379,N_3080,N_2502);
nor UO_380 (O_380,N_4083,N_2584);
nand UO_381 (O_381,N_3834,N_4688);
and UO_382 (O_382,N_4123,N_2919);
nor UO_383 (O_383,N_3889,N_4147);
xor UO_384 (O_384,N_2606,N_2773);
and UO_385 (O_385,N_3785,N_3113);
xnor UO_386 (O_386,N_3530,N_3439);
and UO_387 (O_387,N_3729,N_4269);
or UO_388 (O_388,N_3111,N_4825);
nand UO_389 (O_389,N_3651,N_2509);
and UO_390 (O_390,N_4952,N_3132);
nand UO_391 (O_391,N_4496,N_4977);
nor UO_392 (O_392,N_2973,N_3928);
and UO_393 (O_393,N_4343,N_4932);
xnor UO_394 (O_394,N_3713,N_4294);
and UO_395 (O_395,N_4953,N_3286);
nor UO_396 (O_396,N_2641,N_4380);
xor UO_397 (O_397,N_4536,N_3623);
xor UO_398 (O_398,N_4993,N_4758);
xor UO_399 (O_399,N_4111,N_2901);
or UO_400 (O_400,N_4342,N_3095);
xor UO_401 (O_401,N_4997,N_4079);
and UO_402 (O_402,N_3519,N_3648);
xor UO_403 (O_403,N_3031,N_3152);
xor UO_404 (O_404,N_3903,N_4696);
nand UO_405 (O_405,N_3937,N_4225);
nor UO_406 (O_406,N_2833,N_3346);
or UO_407 (O_407,N_2802,N_3154);
nor UO_408 (O_408,N_4698,N_2920);
or UO_409 (O_409,N_4011,N_4281);
and UO_410 (O_410,N_3284,N_3473);
and UO_411 (O_411,N_3305,N_3588);
xnor UO_412 (O_412,N_2760,N_4413);
nand UO_413 (O_413,N_4197,N_3477);
and UO_414 (O_414,N_3340,N_3664);
and UO_415 (O_415,N_4918,N_3977);
or UO_416 (O_416,N_4774,N_4328);
nand UO_417 (O_417,N_4717,N_4562);
and UO_418 (O_418,N_4900,N_2536);
nor UO_419 (O_419,N_3679,N_4060);
and UO_420 (O_420,N_3726,N_2809);
nand UO_421 (O_421,N_4468,N_3529);
nor UO_422 (O_422,N_2861,N_3127);
nor UO_423 (O_423,N_4467,N_2550);
nor UO_424 (O_424,N_4411,N_4607);
xor UO_425 (O_425,N_2603,N_2650);
nor UO_426 (O_426,N_4400,N_4782);
and UO_427 (O_427,N_3665,N_3910);
or UO_428 (O_428,N_3642,N_3747);
nor UO_429 (O_429,N_2815,N_3335);
and UO_430 (O_430,N_4896,N_4891);
and UO_431 (O_431,N_2735,N_3351);
and UO_432 (O_432,N_4137,N_4447);
and UO_433 (O_433,N_4058,N_4760);
or UO_434 (O_434,N_4901,N_2801);
xnor UO_435 (O_435,N_4592,N_3658);
nand UO_436 (O_436,N_4967,N_3001);
nand UO_437 (O_437,N_2969,N_4317);
xnor UO_438 (O_438,N_3195,N_4285);
or UO_439 (O_439,N_3355,N_4898);
or UO_440 (O_440,N_4017,N_3769);
and UO_441 (O_441,N_2659,N_3779);
nand UO_442 (O_442,N_3804,N_3170);
nor UO_443 (O_443,N_3362,N_4518);
and UO_444 (O_444,N_3844,N_3173);
nand UO_445 (O_445,N_3715,N_2947);
xnor UO_446 (O_446,N_3636,N_3371);
nor UO_447 (O_447,N_4212,N_2814);
or UO_448 (O_448,N_3570,N_3070);
nor UO_449 (O_449,N_2759,N_4109);
and UO_450 (O_450,N_4667,N_4275);
xnor UO_451 (O_451,N_4252,N_2930);
nor UO_452 (O_452,N_3878,N_3976);
nor UO_453 (O_453,N_3435,N_3827);
nor UO_454 (O_454,N_2708,N_4019);
and UO_455 (O_455,N_3012,N_3885);
nor UO_456 (O_456,N_4681,N_3171);
nand UO_457 (O_457,N_3352,N_3652);
or UO_458 (O_458,N_2908,N_2687);
nand UO_459 (O_459,N_2909,N_2665);
or UO_460 (O_460,N_4818,N_4926);
nand UO_461 (O_461,N_3079,N_4632);
nor UO_462 (O_462,N_4988,N_3763);
and UO_463 (O_463,N_3629,N_4557);
nor UO_464 (O_464,N_2987,N_4500);
and UO_465 (O_465,N_3243,N_3947);
xnor UO_466 (O_466,N_3158,N_4318);
and UO_467 (O_467,N_3518,N_3707);
or UO_468 (O_468,N_2928,N_4887);
and UO_469 (O_469,N_3838,N_4651);
nand UO_470 (O_470,N_3697,N_4941);
and UO_471 (O_471,N_2777,N_2645);
nor UO_472 (O_472,N_3045,N_4946);
and UO_473 (O_473,N_3772,N_3788);
nor UO_474 (O_474,N_2635,N_3923);
xor UO_475 (O_475,N_3847,N_3109);
or UO_476 (O_476,N_3451,N_2883);
nand UO_477 (O_477,N_2697,N_4360);
or UO_478 (O_478,N_3842,N_2627);
and UO_479 (O_479,N_4228,N_4288);
nor UO_480 (O_480,N_4055,N_2865);
or UO_481 (O_481,N_4839,N_4329);
or UO_482 (O_482,N_4311,N_4483);
nand UO_483 (O_483,N_3704,N_3791);
nor UO_484 (O_484,N_3853,N_3945);
or UO_485 (O_485,N_3021,N_3450);
nor UO_486 (O_486,N_4232,N_3254);
and UO_487 (O_487,N_4981,N_4874);
or UO_488 (O_488,N_2728,N_2824);
and UO_489 (O_489,N_4381,N_3874);
nand UO_490 (O_490,N_3502,N_2558);
nor UO_491 (O_491,N_3409,N_4965);
nand UO_492 (O_492,N_4844,N_3303);
or UO_493 (O_493,N_3862,N_3890);
nand UO_494 (O_494,N_4718,N_4066);
nor UO_495 (O_495,N_4867,N_3777);
and UO_496 (O_496,N_3285,N_3053);
or UO_497 (O_497,N_3873,N_4442);
or UO_498 (O_498,N_3347,N_4449);
nand UO_499 (O_499,N_4807,N_4504);
nor UO_500 (O_500,N_3250,N_3264);
nand UO_501 (O_501,N_3057,N_4537);
nand UO_502 (O_502,N_2541,N_2562);
and UO_503 (O_503,N_4772,N_4157);
nor UO_504 (O_504,N_4585,N_3662);
or UO_505 (O_505,N_3271,N_3741);
nand UO_506 (O_506,N_2788,N_4868);
xor UO_507 (O_507,N_3384,N_4502);
xor UO_508 (O_508,N_2607,N_3316);
xnor UO_509 (O_509,N_4579,N_4820);
and UO_510 (O_510,N_4516,N_3222);
nand UO_511 (O_511,N_4150,N_2854);
or UO_512 (O_512,N_4097,N_3943);
and UO_513 (O_513,N_2593,N_3281);
or UO_514 (O_514,N_3128,N_3199);
nor UO_515 (O_515,N_3233,N_3353);
nor UO_516 (O_516,N_3090,N_4935);
and UO_517 (O_517,N_3332,N_3049);
and UO_518 (O_518,N_3540,N_4312);
xnor UO_519 (O_519,N_2902,N_3583);
xnor UO_520 (O_520,N_4369,N_4513);
or UO_521 (O_521,N_4791,N_2702);
or UO_522 (O_522,N_3757,N_4309);
and UO_523 (O_523,N_4170,N_4784);
or UO_524 (O_524,N_3986,N_4026);
or UO_525 (O_525,N_4866,N_2800);
xnor UO_526 (O_526,N_2867,N_3699);
and UO_527 (O_527,N_3459,N_4488);
xor UO_528 (O_528,N_2742,N_2754);
and UO_529 (O_529,N_3228,N_4132);
or UO_530 (O_530,N_3557,N_4558);
xnor UO_531 (O_531,N_2705,N_3674);
and UO_532 (O_532,N_4363,N_3032);
xnor UO_533 (O_533,N_3612,N_3117);
nor UO_534 (O_534,N_2507,N_3731);
and UO_535 (O_535,N_2855,N_2988);
nand UO_536 (O_536,N_4286,N_3985);
nand UO_537 (O_537,N_4198,N_4074);
xnor UO_538 (O_538,N_3645,N_3075);
nand UO_539 (O_539,N_4805,N_4598);
nor UO_540 (O_540,N_4551,N_4864);
xor UO_541 (O_541,N_3007,N_3442);
nand UO_542 (O_542,N_4563,N_3236);
nand UO_543 (O_543,N_3799,N_4176);
xnor UO_544 (O_544,N_3382,N_2965);
and UO_545 (O_545,N_2842,N_2871);
or UO_546 (O_546,N_3258,N_4056);
xnor UO_547 (O_547,N_4226,N_4306);
nand UO_548 (O_548,N_3669,N_4434);
or UO_549 (O_549,N_4489,N_3280);
and UO_550 (O_550,N_3800,N_4532);
nor UO_551 (O_551,N_4878,N_4798);
nor UO_552 (O_552,N_2974,N_4122);
xor UO_553 (O_553,N_3103,N_3349);
xor UO_554 (O_554,N_4852,N_4448);
xor UO_555 (O_555,N_4508,N_4464);
nand UO_556 (O_556,N_3939,N_3456);
nand UO_557 (O_557,N_4811,N_3861);
xor UO_558 (O_558,N_4837,N_3782);
nor UO_559 (O_559,N_3802,N_3455);
nor UO_560 (O_560,N_3268,N_4623);
and UO_561 (O_561,N_2521,N_4989);
nand UO_562 (O_562,N_3632,N_3925);
nor UO_563 (O_563,N_3934,N_4410);
or UO_564 (O_564,N_4227,N_3381);
xor UO_565 (O_565,N_2979,N_4757);
nand UO_566 (O_566,N_4913,N_2553);
nor UO_567 (O_567,N_3065,N_2836);
or UO_568 (O_568,N_2706,N_4601);
nand UO_569 (O_569,N_2880,N_4487);
nand UO_570 (O_570,N_2799,N_3984);
xnor UO_571 (O_571,N_3749,N_4134);
or UO_572 (O_572,N_2962,N_3598);
or UO_573 (O_573,N_2807,N_3640);
nor UO_574 (O_574,N_4709,N_4133);
nor UO_575 (O_575,N_3933,N_3740);
xnor UO_576 (O_576,N_2618,N_3617);
nand UO_577 (O_577,N_4081,N_3857);
or UO_578 (O_578,N_2572,N_4255);
nand UO_579 (O_579,N_3242,N_3992);
or UO_580 (O_580,N_2672,N_3722);
xnor UO_581 (O_581,N_3315,N_4582);
nand UO_582 (O_582,N_4051,N_4046);
xor UO_583 (O_583,N_4570,N_3655);
or UO_584 (O_584,N_4729,N_4106);
and UO_585 (O_585,N_4403,N_4293);
xnor UO_586 (O_586,N_4845,N_3186);
nand UO_587 (O_587,N_4007,N_3593);
or UO_588 (O_588,N_4391,N_2506);
nand UO_589 (O_589,N_3613,N_3850);
xnor UO_590 (O_590,N_3330,N_2675);
and UO_591 (O_591,N_4096,N_4078);
nor UO_592 (O_592,N_2612,N_4044);
nor UO_593 (O_593,N_4828,N_3118);
nor UO_594 (O_594,N_4179,N_3516);
nand UO_595 (O_595,N_4940,N_4514);
nand UO_596 (O_596,N_4167,N_4910);
and UO_597 (O_597,N_3139,N_2691);
and UO_598 (O_598,N_2757,N_3498);
or UO_599 (O_599,N_4205,N_4835);
or UO_600 (O_600,N_3653,N_4184);
nor UO_601 (O_601,N_4276,N_4223);
or UO_602 (O_602,N_2797,N_3336);
and UO_603 (O_603,N_2734,N_3009);
and UO_604 (O_604,N_3300,N_3256);
or UO_605 (O_605,N_3448,N_4600);
or UO_606 (O_606,N_3591,N_3643);
and UO_607 (O_607,N_2822,N_3331);
xor UO_608 (O_608,N_2616,N_3620);
xnor UO_609 (O_609,N_2918,N_3724);
nor UO_610 (O_610,N_4307,N_3509);
or UO_611 (O_611,N_3956,N_4748);
nor UO_612 (O_612,N_3619,N_4432);
nand UO_613 (O_613,N_3488,N_3575);
nand UO_614 (O_614,N_3160,N_3823);
xnor UO_615 (O_615,N_4606,N_4808);
or UO_616 (O_616,N_4849,N_3867);
nor UO_617 (O_617,N_4806,N_3174);
or UO_618 (O_618,N_4613,N_2651);
nor UO_619 (O_619,N_3482,N_4266);
nor UO_620 (O_620,N_3453,N_3538);
or UO_621 (O_621,N_3417,N_2514);
nand UO_622 (O_622,N_3864,N_4189);
nand UO_623 (O_623,N_3140,N_3011);
and UO_624 (O_624,N_2590,N_4101);
and UO_625 (O_625,N_4745,N_3430);
or UO_626 (O_626,N_4673,N_2738);
nor UO_627 (O_627,N_4794,N_2714);
nor UO_628 (O_628,N_3567,N_4022);
xnor UO_629 (O_629,N_3825,N_4510);
or UO_630 (O_630,N_3760,N_3304);
xnor UO_631 (O_631,N_4614,N_3753);
or UO_632 (O_632,N_2741,N_3102);
and UO_633 (O_633,N_3695,N_2636);
or UO_634 (O_634,N_4138,N_2658);
nand UO_635 (O_635,N_3694,N_3282);
or UO_636 (O_636,N_4210,N_2643);
xnor UO_637 (O_637,N_2630,N_2669);
or UO_638 (O_638,N_4365,N_4348);
and UO_639 (O_639,N_3410,N_4975);
xnor UO_640 (O_640,N_3087,N_2652);
nand UO_641 (O_641,N_4657,N_4625);
nand UO_642 (O_642,N_2903,N_3656);
nand UO_643 (O_643,N_4694,N_3370);
or UO_644 (O_644,N_3016,N_3181);
or UO_645 (O_645,N_4597,N_4440);
or UO_646 (O_646,N_3365,N_4559);
and UO_647 (O_647,N_3393,N_3618);
or UO_648 (O_648,N_4917,N_2952);
and UO_649 (O_649,N_4088,N_4015);
nand UO_650 (O_650,N_3151,N_3364);
or UO_651 (O_651,N_4644,N_4165);
nor UO_652 (O_652,N_4393,N_4527);
and UO_653 (O_653,N_3711,N_2673);
and UO_654 (O_654,N_4553,N_4472);
nor UO_655 (O_655,N_3027,N_3018);
and UO_656 (O_656,N_3703,N_4443);
and UO_657 (O_657,N_4526,N_2768);
nand UO_658 (O_658,N_2604,N_4972);
nor UO_659 (O_659,N_2904,N_3966);
nor UO_660 (O_660,N_3397,N_4604);
nand UO_661 (O_661,N_3175,N_3868);
or UO_662 (O_662,N_3374,N_4379);
nor UO_663 (O_663,N_3510,N_3147);
nor UO_664 (O_664,N_3599,N_3544);
nor UO_665 (O_665,N_3094,N_2873);
or UO_666 (O_666,N_2531,N_4422);
or UO_667 (O_667,N_4572,N_4731);
and UO_668 (O_668,N_3708,N_2628);
nand UO_669 (O_669,N_2704,N_2874);
and UO_670 (O_670,N_4646,N_4809);
xor UO_671 (O_671,N_3014,N_4073);
nand UO_672 (O_672,N_3810,N_2862);
or UO_673 (O_673,N_3480,N_4368);
nor UO_674 (O_674,N_3144,N_4622);
nor UO_675 (O_675,N_3006,N_3573);
nor UO_676 (O_676,N_2569,N_4509);
and UO_677 (O_677,N_3577,N_3454);
nand UO_678 (O_678,N_3683,N_3465);
and UO_679 (O_679,N_4258,N_3295);
xor UO_680 (O_680,N_2671,N_3639);
xor UO_681 (O_681,N_3437,N_4439);
nand UO_682 (O_682,N_4649,N_4402);
nand UO_683 (O_683,N_3212,N_3805);
nand UO_684 (O_684,N_3163,N_3935);
nor UO_685 (O_685,N_4554,N_3311);
nand UO_686 (O_686,N_3072,N_4771);
nor UO_687 (O_687,N_4621,N_4490);
nor UO_688 (O_688,N_4873,N_2953);
or UO_689 (O_689,N_3178,N_3048);
nand UO_690 (O_690,N_3701,N_4616);
nand UO_691 (O_691,N_3902,N_4203);
nor UO_692 (O_692,N_4367,N_3143);
or UO_693 (O_693,N_4351,N_4973);
nor UO_694 (O_694,N_3056,N_3650);
xnor UO_695 (O_695,N_2666,N_4190);
and UO_696 (O_696,N_2771,N_2642);
or UO_697 (O_697,N_2574,N_3129);
nor UO_698 (O_698,N_2884,N_3672);
and UO_699 (O_699,N_3202,N_3321);
and UO_700 (O_700,N_2984,N_4155);
nand UO_701 (O_701,N_4847,N_3605);
and UO_702 (O_702,N_3002,N_4764);
or UO_703 (O_703,N_2510,N_3210);
nor UO_704 (O_704,N_4556,N_4018);
and UO_705 (O_705,N_3040,N_3348);
nor UO_706 (O_706,N_3948,N_3647);
nor UO_707 (O_707,N_4063,N_3037);
or UO_708 (O_708,N_3600,N_3277);
nand UO_709 (O_709,N_3373,N_3165);
xnor UO_710 (O_710,N_3744,N_3479);
or UO_711 (O_711,N_4936,N_4826);
nor UO_712 (O_712,N_3809,N_4436);
or UO_713 (O_713,N_2934,N_2713);
nand UO_714 (O_714,N_4802,N_2613);
and UO_715 (O_715,N_3356,N_3869);
xnor UO_716 (O_716,N_3291,N_2900);
nand UO_717 (O_717,N_3218,N_4283);
nor UO_718 (O_718,N_4308,N_3043);
xor UO_719 (O_719,N_4895,N_3367);
xor UO_720 (O_720,N_4076,N_2626);
nor UO_721 (O_721,N_2977,N_4461);
nor UO_722 (O_722,N_4909,N_3796);
or UO_723 (O_723,N_2560,N_4270);
and UO_724 (O_724,N_4376,N_3252);
nand UO_725 (O_725,N_4762,N_3635);
nand UO_726 (O_726,N_4139,N_4499);
or UO_727 (O_727,N_3756,N_2564);
and UO_728 (O_728,N_3402,N_4395);
or UO_729 (O_729,N_2829,N_4177);
and UO_730 (O_730,N_4658,N_4995);
or UO_731 (O_731,N_4577,N_4337);
nor UO_732 (O_732,N_3508,N_4633);
or UO_733 (O_733,N_3100,N_4531);
or UO_734 (O_734,N_3512,N_2795);
nand UO_735 (O_735,N_3411,N_3024);
and UO_736 (O_736,N_3372,N_3213);
nand UO_737 (O_737,N_3912,N_3671);
or UO_738 (O_738,N_4473,N_2976);
and UO_739 (O_739,N_2528,N_2963);
nand UO_740 (O_740,N_3644,N_4113);
nand UO_741 (O_741,N_4817,N_3849);
and UO_742 (O_742,N_3325,N_3765);
and UO_743 (O_743,N_3071,N_3190);
xnor UO_744 (O_744,N_2596,N_3142);
xor UO_745 (O_745,N_3604,N_2761);
nand UO_746 (O_746,N_4628,N_4485);
and UO_747 (O_747,N_4753,N_2551);
and UO_748 (O_748,N_4115,N_2752);
xnor UO_749 (O_749,N_3983,N_4727);
nand UO_750 (O_750,N_4545,N_4684);
nand UO_751 (O_751,N_3201,N_4627);
nor UO_752 (O_752,N_3667,N_3721);
and UO_753 (O_753,N_3551,N_4175);
and UO_754 (O_754,N_3164,N_4815);
and UO_755 (O_755,N_3539,N_2670);
xor UO_756 (O_756,N_4388,N_3249);
nor UO_757 (O_757,N_3524,N_3240);
or UO_758 (O_758,N_4314,N_3046);
nor UO_759 (O_759,N_3661,N_4477);
and UO_760 (O_760,N_4126,N_3387);
nand UO_761 (O_761,N_4978,N_3649);
or UO_762 (O_762,N_4880,N_3970);
and UO_763 (O_763,N_4823,N_3467);
or UO_764 (O_764,N_2899,N_4573);
and UO_765 (O_765,N_4456,N_4575);
nand UO_766 (O_766,N_2885,N_3875);
and UO_767 (O_767,N_4021,N_3423);
xor UO_768 (O_768,N_4062,N_3083);
or UO_769 (O_769,N_3829,N_3627);
nor UO_770 (O_770,N_3988,N_4838);
xnor UO_771 (O_771,N_3022,N_3900);
nor UO_772 (O_772,N_3969,N_2557);
nand UO_773 (O_773,N_2711,N_4257);
nor UO_774 (O_774,N_4121,N_3917);
and UO_775 (O_775,N_2622,N_3670);
and UO_776 (O_776,N_3720,N_3511);
or UO_777 (O_777,N_3837,N_2810);
or UO_778 (O_778,N_4033,N_4754);
nor UO_779 (O_779,N_3013,N_3265);
or UO_780 (O_780,N_4267,N_2715);
nor UO_781 (O_781,N_4702,N_3893);
nor UO_782 (O_782,N_4843,N_3179);
or UO_783 (O_783,N_4609,N_2762);
and UO_784 (O_784,N_3880,N_2804);
nor UO_785 (O_785,N_3431,N_3952);
nand UO_786 (O_786,N_4282,N_4093);
xnor UO_787 (O_787,N_4869,N_3225);
or UO_788 (O_788,N_3506,N_4045);
or UO_789 (O_789,N_4642,N_2852);
xor UO_790 (O_790,N_3905,N_3997);
nand UO_791 (O_791,N_2542,N_4335);
and UO_792 (O_792,N_3723,N_4799);
or UO_793 (O_793,N_4196,N_2964);
nand UO_794 (O_794,N_3122,N_3389);
nor UO_795 (O_795,N_3093,N_4065);
nor UO_796 (O_796,N_3798,N_3587);
or UO_797 (O_797,N_2889,N_4087);
nand UO_798 (O_798,N_2943,N_3637);
nand UO_799 (O_799,N_3400,N_3026);
xor UO_800 (O_800,N_3198,N_2986);
or UO_801 (O_801,N_4216,N_3743);
or UO_802 (O_802,N_3390,N_3299);
nor UO_803 (O_803,N_4385,N_4030);
nor UO_804 (O_804,N_2915,N_4049);
nand UO_805 (O_805,N_4054,N_3835);
nor UO_806 (O_806,N_2694,N_3714);
nor UO_807 (O_807,N_2620,N_3091);
nor UO_808 (O_808,N_4976,N_3149);
and UO_809 (O_809,N_4544,N_3217);
xor UO_810 (O_810,N_3995,N_2597);
xor UO_811 (O_811,N_3269,N_4480);
and UO_812 (O_812,N_3801,N_3601);
or UO_813 (O_813,N_3863,N_3403);
xor UO_814 (O_814,N_2500,N_3532);
nand UO_815 (O_815,N_3219,N_2954);
nand UO_816 (O_816,N_2623,N_4336);
nor UO_817 (O_817,N_4834,N_4934);
xor UO_818 (O_818,N_3831,N_2684);
nor UO_819 (O_819,N_3841,N_4373);
or UO_820 (O_820,N_3497,N_4135);
nand UO_821 (O_821,N_4195,N_4287);
nand UO_822 (O_822,N_3735,N_3200);
nand UO_823 (O_823,N_4971,N_2805);
or UO_824 (O_824,N_2791,N_3556);
and UO_825 (O_825,N_4911,N_2813);
and UO_826 (O_826,N_2905,N_3924);
xor UO_827 (O_827,N_2647,N_3501);
nand UO_828 (O_828,N_3494,N_3836);
and UO_829 (O_829,N_2534,N_4733);
nand UO_830 (O_830,N_2526,N_4547);
nand UO_831 (O_831,N_3290,N_4507);
or UO_832 (O_832,N_4812,N_2726);
nand UO_833 (O_833,N_2721,N_2744);
or UO_834 (O_834,N_4552,N_4983);
or UO_835 (O_835,N_2517,N_3344);
xnor UO_836 (O_836,N_3110,N_2725);
nor UO_837 (O_837,N_3797,N_2678);
nor UO_838 (O_838,N_2921,N_3700);
and UO_839 (O_839,N_3682,N_4322);
or UO_840 (O_840,N_2653,N_2661);
nor UO_841 (O_841,N_3775,N_3668);
nand UO_842 (O_842,N_2546,N_3345);
or UO_843 (O_843,N_4914,N_3786);
and UO_844 (O_844,N_3481,N_4634);
nor UO_845 (O_845,N_2960,N_3828);
nor UO_846 (O_846,N_3405,N_2737);
or UO_847 (O_847,N_4700,N_2776);
nand UO_848 (O_848,N_4043,N_2787);
xnor UO_849 (O_849,N_3940,N_3525);
xnor UO_850 (O_850,N_4236,N_2756);
nand UO_851 (O_851,N_2632,N_4752);
nand UO_852 (O_852,N_3754,N_3413);
xor UO_853 (O_853,N_3468,N_4693);
xnor UO_854 (O_854,N_3625,N_4469);
or UO_855 (O_855,N_4780,N_3633);
and UO_856 (O_856,N_4071,N_4801);
nor UO_857 (O_857,N_2820,N_4755);
or UO_858 (O_858,N_4576,N_3585);
or UO_859 (O_859,N_4785,N_4610);
nand UO_860 (O_860,N_4511,N_3595);
nand UO_861 (O_861,N_3751,N_4159);
and UO_862 (O_862,N_3979,N_2677);
nand UO_863 (O_863,N_4555,N_3858);
nor UO_864 (O_864,N_4665,N_3555);
nor UO_865 (O_865,N_3247,N_3447);
nor UO_866 (O_866,N_4072,N_3432);
nor UO_867 (O_867,N_4679,N_4331);
or UO_868 (O_868,N_4543,N_4638);
nor UO_869 (O_869,N_2629,N_4534);
nand UO_870 (O_870,N_2699,N_3534);
nand UO_871 (O_871,N_2941,N_4173);
xor UO_872 (O_872,N_4888,N_4375);
and UO_873 (O_873,N_3596,N_3654);
and UO_874 (O_874,N_4404,N_4313);
or UO_875 (O_875,N_2992,N_4870);
or UO_876 (O_876,N_3052,N_4090);
nor UO_877 (O_877,N_2982,N_4187);
nand UO_878 (O_878,N_4171,N_3357);
and UO_879 (O_879,N_2566,N_3339);
or UO_880 (O_880,N_4945,N_3548);
nor UO_881 (O_881,N_2580,N_3892);
nor UO_882 (O_882,N_2958,N_2924);
nor UO_883 (O_883,N_4102,N_3778);
or UO_884 (O_884,N_3965,N_3192);
or UO_885 (O_885,N_3541,N_3084);
or UO_886 (O_886,N_4215,N_3272);
nor UO_887 (O_887,N_4611,N_3921);
xnor UO_888 (O_888,N_3239,N_2877);
or UO_889 (O_889,N_3712,N_3689);
or UO_890 (O_890,N_4703,N_4353);
and UO_891 (O_891,N_4300,N_2935);
and UO_892 (O_892,N_2933,N_3815);
nand UO_893 (O_893,N_3038,N_4863);
or UO_894 (O_894,N_3401,N_4943);
xnor UO_895 (O_895,N_4747,N_4191);
nor UO_896 (O_896,N_3066,N_3659);
or UO_897 (O_897,N_3978,N_4221);
nor UO_898 (O_898,N_4142,N_4907);
or UO_899 (O_899,N_3063,N_4862);
xor UO_900 (O_900,N_3396,N_4324);
nor UO_901 (O_901,N_4250,N_4691);
nand UO_902 (O_902,N_3354,N_3964);
or UO_903 (O_903,N_3221,N_2989);
nand UO_904 (O_904,N_3408,N_2530);
or UO_905 (O_905,N_4358,N_3830);
nor UO_906 (O_906,N_4574,N_4992);
nor UO_907 (O_907,N_4417,N_4906);
xnor UO_908 (O_908,N_2668,N_3425);
and UO_909 (O_909,N_3324,N_2763);
nand UO_910 (O_910,N_4000,N_3673);
and UO_911 (O_911,N_4959,N_3172);
or UO_912 (O_912,N_3794,N_4182);
or UO_913 (O_913,N_4786,N_4217);
and UO_914 (O_914,N_3990,N_3550);
xnor UO_915 (O_915,N_3229,N_3646);
and UO_916 (O_916,N_4475,N_2819);
xnor UO_917 (O_917,N_4010,N_4192);
nand UO_918 (O_918,N_3898,N_4879);
and UO_919 (O_919,N_3232,N_4737);
nand UO_920 (O_920,N_3317,N_3918);
and UO_921 (O_921,N_3197,N_2893);
and UO_922 (O_922,N_4716,N_4858);
nand UO_923 (O_923,N_4840,N_3686);
xnor UO_924 (O_924,N_4104,N_3920);
nand UO_925 (O_925,N_3248,N_4599);
nor UO_926 (O_926,N_4769,N_3677);
or UO_927 (O_927,N_4955,N_4246);
xor UO_928 (O_928,N_3273,N_4320);
nand UO_929 (O_929,N_2568,N_4006);
nor UO_930 (O_930,N_4734,N_4305);
or UO_931 (O_931,N_3692,N_4736);
or UO_932 (O_932,N_3427,N_3981);
nor UO_933 (O_933,N_3327,N_2554);
xor UO_934 (O_934,N_4116,N_2847);
and UO_935 (O_935,N_3406,N_2949);
and UO_936 (O_936,N_3169,N_2573);
or UO_937 (O_937,N_2595,N_3993);
nor UO_938 (O_938,N_4501,N_2688);
nor UO_939 (O_939,N_2793,N_4647);
and UO_940 (O_940,N_4857,N_4466);
xnor UO_941 (O_941,N_4249,N_3531);
or UO_942 (O_942,N_3074,N_4730);
or UO_943 (O_943,N_2579,N_4387);
or UO_944 (O_944,N_3104,N_3941);
or UO_945 (O_945,N_4595,N_2693);
and UO_946 (O_946,N_3680,N_3505);
nor UO_947 (O_947,N_4382,N_3020);
and UO_948 (O_948,N_3434,N_4310);
and UO_949 (O_949,N_4648,N_4136);
and UO_950 (O_950,N_4821,N_3931);
or UO_951 (O_951,N_4350,N_3137);
nand UO_952 (O_952,N_3019,N_4347);
and UO_953 (O_953,N_4775,N_3883);
nand UO_954 (O_954,N_3279,N_2910);
nand UO_955 (O_955,N_3994,N_3424);
and UO_956 (O_956,N_2844,N_3839);
nor UO_957 (O_957,N_4704,N_2838);
nor UO_958 (O_958,N_4813,N_4540);
nor UO_959 (O_959,N_4789,N_3840);
nand UO_960 (O_960,N_4881,N_2931);
or UO_961 (O_961,N_2792,N_3872);
nand UO_962 (O_962,N_3464,N_3776);
nand UO_963 (O_963,N_4664,N_3553);
and UO_964 (O_964,N_4271,N_3495);
or UO_965 (O_965,N_4966,N_3989);
and UO_966 (O_966,N_2940,N_2703);
nand UO_967 (O_967,N_3717,N_4792);
or UO_968 (O_968,N_3469,N_3125);
nand UO_969 (O_969,N_4479,N_4777);
or UO_970 (O_970,N_4669,N_4596);
nand UO_971 (O_971,N_4986,N_4105);
nand UO_972 (O_972,N_3214,N_2769);
and UO_973 (O_973,N_3991,N_3486);
or UO_974 (O_974,N_3098,N_4705);
nor UO_975 (O_975,N_2846,N_4042);
nor UO_976 (O_976,N_4505,N_4233);
and UO_977 (O_977,N_3015,N_4024);
and UO_978 (O_978,N_3824,N_2857);
xor UO_979 (O_979,N_4211,N_3818);
or UO_980 (O_980,N_3395,N_3914);
and UO_981 (O_981,N_4168,N_2746);
nand UO_982 (O_982,N_4392,N_3166);
nand UO_983 (O_983,N_2876,N_3881);
nor UO_984 (O_984,N_3609,N_3196);
nand UO_985 (O_985,N_4409,N_3436);
nor UO_986 (O_986,N_3580,N_3096);
nor UO_987 (O_987,N_3224,N_4778);
or UO_988 (O_988,N_3552,N_4711);
and UO_989 (O_989,N_4428,N_4697);
nand UO_990 (O_990,N_4334,N_3491);
or UO_991 (O_991,N_3120,N_2689);
or UO_992 (O_992,N_4481,N_2504);
xor UO_993 (O_993,N_3193,N_4299);
nand UO_994 (O_994,N_3887,N_4692);
nor UO_995 (O_995,N_4533,N_4517);
or UO_996 (O_996,N_2990,N_4284);
xor UO_997 (O_997,N_4430,N_3808);
nor UO_998 (O_998,N_2739,N_2796);
nand UO_999 (O_999,N_4947,N_2929);
endmodule