module basic_750_5000_1000_5_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_722,In_635);
nor U1 (N_1,In_511,In_185);
nand U2 (N_2,In_9,In_564);
and U3 (N_3,In_705,In_547);
or U4 (N_4,In_42,In_278);
and U5 (N_5,In_420,In_574);
or U6 (N_6,In_177,In_436);
nand U7 (N_7,In_597,In_634);
and U8 (N_8,In_71,In_224);
nand U9 (N_9,In_54,In_405);
or U10 (N_10,In_304,In_173);
nor U11 (N_11,In_65,In_676);
nor U12 (N_12,In_552,In_95);
or U13 (N_13,In_711,In_736);
xor U14 (N_14,In_656,In_460);
nand U15 (N_15,In_56,In_260);
or U16 (N_16,In_474,In_67);
and U17 (N_17,In_629,In_164);
or U18 (N_18,In_165,In_307);
or U19 (N_19,In_333,In_653);
and U20 (N_20,In_465,In_598);
or U21 (N_21,In_674,In_24);
nand U22 (N_22,In_317,In_84);
nor U23 (N_23,In_223,In_663);
nor U24 (N_24,In_619,In_251);
nand U25 (N_25,In_275,In_428);
or U26 (N_26,In_562,In_162);
xor U27 (N_27,In_581,In_683);
nor U28 (N_28,In_369,In_612);
nor U29 (N_29,In_521,In_27);
and U30 (N_30,In_684,In_253);
and U31 (N_31,In_572,In_394);
or U32 (N_32,In_126,In_397);
or U33 (N_33,In_345,In_290);
and U34 (N_34,In_77,In_380);
nor U35 (N_35,In_403,In_323);
nor U36 (N_36,In_549,In_396);
and U37 (N_37,In_152,In_376);
or U38 (N_38,In_678,In_721);
nor U39 (N_39,In_603,In_608);
nand U40 (N_40,In_500,In_208);
nor U41 (N_41,In_681,In_669);
nor U42 (N_42,In_391,In_207);
or U43 (N_43,In_2,In_483);
nand U44 (N_44,In_337,In_433);
nor U45 (N_45,In_194,In_386);
and U46 (N_46,In_110,In_475);
nand U47 (N_47,In_144,In_692);
nand U48 (N_48,In_216,In_537);
or U49 (N_49,In_593,In_719);
and U50 (N_50,In_335,In_256);
or U51 (N_51,In_180,In_648);
nor U52 (N_52,In_363,In_170);
nor U53 (N_53,In_244,In_248);
and U54 (N_54,In_489,In_49);
or U55 (N_55,In_638,In_133);
and U56 (N_56,In_390,In_192);
or U57 (N_57,In_37,In_577);
nor U58 (N_58,In_236,In_136);
nand U59 (N_59,In_375,In_111);
and U60 (N_60,In_688,In_350);
or U61 (N_61,In_617,In_140);
and U62 (N_62,In_568,In_195);
and U63 (N_63,In_621,In_199);
nor U64 (N_64,In_543,In_203);
nand U65 (N_65,In_353,In_519);
and U66 (N_66,In_263,In_11);
or U67 (N_67,In_70,In_163);
or U68 (N_68,In_252,In_540);
and U69 (N_69,In_690,In_423);
xnor U70 (N_70,In_698,In_295);
nor U71 (N_71,In_633,In_576);
nand U72 (N_72,In_28,In_230);
and U73 (N_73,In_117,In_132);
or U74 (N_74,In_35,In_109);
nand U75 (N_75,In_33,In_101);
nand U76 (N_76,In_286,In_639);
nor U77 (N_77,In_416,In_366);
nand U78 (N_78,In_455,In_298);
or U79 (N_79,In_351,In_343);
nand U80 (N_80,In_348,In_266);
nand U81 (N_81,In_495,In_349);
nand U82 (N_82,In_127,In_580);
nand U83 (N_83,In_419,In_399);
and U84 (N_84,In_148,In_505);
or U85 (N_85,In_478,In_518);
nand U86 (N_86,In_594,In_229);
xor U87 (N_87,In_430,In_691);
and U88 (N_88,In_701,In_299);
or U89 (N_89,In_389,In_385);
and U90 (N_90,In_280,In_513);
nor U91 (N_91,In_329,In_440);
nor U92 (N_92,In_661,In_586);
nor U93 (N_93,In_636,In_291);
and U94 (N_94,In_306,In_325);
or U95 (N_95,In_447,In_502);
nand U96 (N_96,In_544,In_590);
and U97 (N_97,In_398,In_143);
or U98 (N_98,In_310,In_113);
nor U99 (N_99,In_288,In_167);
nor U100 (N_100,In_431,In_340);
or U101 (N_101,In_331,In_441);
nor U102 (N_102,In_240,In_239);
and U103 (N_103,In_206,In_178);
and U104 (N_104,In_3,In_130);
nand U105 (N_105,In_166,In_566);
nor U106 (N_106,In_293,In_91);
or U107 (N_107,In_411,In_472);
nand U108 (N_108,In_85,In_425);
or U109 (N_109,In_467,In_709);
nand U110 (N_110,In_55,In_749);
and U111 (N_111,In_102,In_13);
and U112 (N_112,In_4,In_451);
xnor U113 (N_113,In_517,In_641);
or U114 (N_114,In_623,In_402);
nor U115 (N_115,In_699,In_99);
or U116 (N_116,In_745,In_614);
or U117 (N_117,In_655,In_535);
nor U118 (N_118,In_90,In_370);
and U119 (N_119,In_695,In_46);
nor U120 (N_120,In_740,In_196);
nand U121 (N_121,In_365,In_625);
nor U122 (N_122,In_606,In_190);
xor U123 (N_123,In_39,In_485);
nand U124 (N_124,In_536,In_7);
xnor U125 (N_125,In_346,In_654);
nor U126 (N_126,In_401,In_727);
nor U127 (N_127,In_22,In_748);
and U128 (N_128,In_120,In_412);
and U129 (N_129,In_480,In_642);
or U130 (N_130,In_496,In_315);
and U131 (N_131,In_245,In_172);
and U132 (N_132,In_332,In_108);
nor U133 (N_133,In_255,In_584);
nand U134 (N_134,In_174,In_358);
and U135 (N_135,In_274,In_19);
nand U136 (N_136,In_632,In_242);
nand U137 (N_137,In_728,In_62);
xor U138 (N_138,In_490,In_508);
and U139 (N_139,In_601,In_339);
nand U140 (N_140,In_732,In_408);
nand U141 (N_141,In_198,In_156);
nor U142 (N_142,In_147,In_302);
and U143 (N_143,In_258,In_418);
and U144 (N_144,In_512,In_637);
nand U145 (N_145,In_539,In_115);
or U146 (N_146,In_462,In_657);
nor U147 (N_147,In_209,In_432);
nand U148 (N_148,In_320,In_344);
or U149 (N_149,In_422,In_80);
nor U150 (N_150,In_383,In_437);
or U151 (N_151,In_600,In_650);
and U152 (N_152,In_526,In_563);
and U153 (N_153,In_300,In_316);
and U154 (N_154,In_289,In_26);
and U155 (N_155,In_527,In_96);
nor U156 (N_156,In_92,In_557);
nor U157 (N_157,In_616,In_741);
nand U158 (N_158,In_371,In_624);
and U159 (N_159,In_682,In_357);
nand U160 (N_160,In_29,In_267);
nand U161 (N_161,In_509,In_730);
nor U162 (N_162,In_538,In_532);
nor U163 (N_163,In_227,In_159);
or U164 (N_164,In_491,In_744);
nor U165 (N_165,In_103,In_469);
nor U166 (N_166,In_622,In_60);
and U167 (N_167,In_43,In_171);
nor U168 (N_168,In_666,In_222);
and U169 (N_169,In_646,In_610);
nor U170 (N_170,In_546,In_555);
nor U171 (N_171,In_314,In_64);
nand U172 (N_172,In_51,In_492);
or U173 (N_173,In_292,In_599);
nor U174 (N_174,In_352,In_561);
nand U175 (N_175,In_107,In_279);
nand U176 (N_176,In_188,In_94);
nor U177 (N_177,In_439,In_149);
nor U178 (N_178,In_76,In_680);
or U179 (N_179,In_146,In_318);
or U180 (N_180,In_78,In_82);
nand U181 (N_181,In_225,In_212);
xor U182 (N_182,In_742,In_201);
and U183 (N_183,In_157,In_651);
and U184 (N_184,In_15,In_98);
xnor U185 (N_185,In_217,In_356);
nand U186 (N_186,In_668,In_720);
and U187 (N_187,In_334,In_313);
or U188 (N_188,In_123,In_183);
and U189 (N_189,In_367,In_501);
and U190 (N_190,In_336,In_360);
and U191 (N_191,In_305,In_435);
or U192 (N_192,In_504,In_382);
and U193 (N_193,In_287,In_724);
nor U194 (N_194,In_457,In_285);
or U195 (N_195,In_712,In_122);
and U196 (N_196,In_541,In_83);
or U197 (N_197,In_393,In_421);
nor U198 (N_198,In_613,In_232);
nor U199 (N_199,In_739,In_114);
and U200 (N_200,In_8,In_182);
nor U201 (N_201,In_718,In_643);
and U202 (N_202,In_707,In_734);
nor U203 (N_203,In_415,In_249);
or U204 (N_204,In_570,In_168);
and U205 (N_205,In_205,In_481);
and U206 (N_206,In_628,In_717);
nand U207 (N_207,In_466,In_630);
nand U208 (N_208,In_246,In_534);
or U209 (N_209,In_254,In_100);
and U210 (N_210,In_677,In_283);
or U211 (N_211,In_671,In_434);
nor U212 (N_212,In_571,In_694);
or U213 (N_213,In_464,In_450);
nor U214 (N_214,In_220,In_342);
or U215 (N_215,In_567,In_296);
nand U216 (N_216,In_73,In_409);
or U217 (N_217,In_530,In_670);
or U218 (N_218,In_587,In_14);
nand U219 (N_219,In_226,In_618);
or U220 (N_220,In_609,In_233);
nor U221 (N_221,In_44,In_326);
and U222 (N_222,In_10,In_551);
nand U223 (N_223,In_506,In_377);
and U224 (N_224,In_262,In_673);
nor U225 (N_225,In_738,In_241);
and U226 (N_226,In_602,In_658);
and U227 (N_227,In_477,In_514);
and U228 (N_228,In_387,In_160);
and U229 (N_229,In_424,In_589);
nor U230 (N_230,In_737,In_235);
nor U231 (N_231,In_347,In_200);
nor U232 (N_232,In_175,In_381);
nor U233 (N_233,In_309,In_40);
or U234 (N_234,In_197,In_213);
nor U235 (N_235,In_221,In_1);
nand U236 (N_236,In_36,In_458);
nand U237 (N_237,In_79,In_75);
and U238 (N_238,In_686,In_259);
nor U239 (N_239,In_118,In_550);
and U240 (N_240,In_311,In_72);
or U241 (N_241,In_583,In_533);
or U242 (N_242,In_58,In_607);
nor U243 (N_243,In_238,In_141);
and U244 (N_244,In_364,In_189);
xnor U245 (N_245,In_372,In_479);
nor U246 (N_246,In_520,In_700);
and U247 (N_247,In_384,In_498);
and U248 (N_248,In_0,In_32);
nand U249 (N_249,In_338,In_124);
nor U250 (N_250,In_88,In_57);
or U251 (N_251,In_575,In_308);
nand U252 (N_252,In_626,In_476);
and U253 (N_253,In_716,In_665);
nor U254 (N_254,In_487,In_703);
xnor U255 (N_255,In_128,In_693);
xnor U256 (N_256,In_17,In_611);
xor U257 (N_257,In_459,In_516);
nand U258 (N_258,In_87,In_303);
or U259 (N_259,In_134,In_214);
nand U260 (N_260,In_560,In_445);
nor U261 (N_261,In_81,In_373);
nor U262 (N_262,In_404,In_247);
nand U263 (N_263,In_158,In_378);
xnor U264 (N_264,In_588,In_228);
or U265 (N_265,In_556,In_294);
or U266 (N_266,In_74,In_47);
nand U267 (N_267,In_406,In_12);
or U268 (N_268,In_438,In_545);
nor U269 (N_269,In_620,In_59);
or U270 (N_270,In_155,In_664);
nand U271 (N_271,In_297,In_470);
nand U272 (N_272,In_585,In_644);
nand U273 (N_273,In_605,In_627);
nand U274 (N_274,In_66,In_282);
and U275 (N_275,In_354,In_368);
and U276 (N_276,In_631,In_503);
nor U277 (N_277,In_204,In_507);
or U278 (N_278,In_142,In_219);
nand U279 (N_279,In_135,In_31);
nand U280 (N_280,In_139,In_548);
nand U281 (N_281,In_672,In_116);
nor U282 (N_282,In_647,In_161);
and U283 (N_283,In_388,In_50);
and U284 (N_284,In_330,In_524);
or U285 (N_285,In_362,In_272);
xor U286 (N_286,In_497,In_5);
or U287 (N_287,In_121,In_592);
or U288 (N_288,In_16,In_689);
nand U289 (N_289,In_687,In_319);
and U290 (N_290,In_429,In_176);
or U291 (N_291,In_34,In_522);
or U292 (N_292,In_93,In_30);
or U293 (N_293,In_270,In_186);
nor U294 (N_294,In_735,In_446);
nand U295 (N_295,In_53,In_486);
or U296 (N_296,In_515,In_410);
and U297 (N_297,In_129,In_97);
nand U298 (N_298,In_324,In_604);
or U299 (N_299,In_708,In_591);
nor U300 (N_300,In_23,In_596);
nand U301 (N_301,In_531,In_104);
nand U302 (N_302,In_181,In_52);
xnor U303 (N_303,In_125,In_105);
or U304 (N_304,In_443,In_442);
or U305 (N_305,In_61,In_106);
nor U306 (N_306,In_528,In_573);
and U307 (N_307,In_456,In_234);
nand U308 (N_308,In_559,In_202);
xnor U309 (N_309,In_355,In_659);
or U310 (N_310,In_321,In_18);
xor U311 (N_311,In_747,In_468);
nor U312 (N_312,In_154,In_112);
nand U313 (N_313,In_427,In_273);
or U314 (N_314,In_257,In_565);
nand U315 (N_315,In_138,In_284);
and U316 (N_316,In_237,In_453);
nor U317 (N_317,In_264,In_696);
and U318 (N_318,In_454,In_704);
nor U319 (N_319,In_269,In_726);
nand U320 (N_320,In_250,In_649);
nand U321 (N_321,In_731,In_471);
or U322 (N_322,In_265,In_729);
and U323 (N_323,In_448,In_452);
or U324 (N_324,In_68,In_675);
xnor U325 (N_325,In_449,In_119);
xnor U326 (N_326,In_400,In_179);
nor U327 (N_327,In_89,In_392);
or U328 (N_328,In_510,In_150);
and U329 (N_329,In_702,In_529);
nor U330 (N_330,In_667,In_341);
or U331 (N_331,In_725,In_25);
and U332 (N_332,In_231,In_281);
and U333 (N_333,In_710,In_714);
or U334 (N_334,In_417,In_322);
nand U335 (N_335,In_268,In_301);
and U336 (N_336,In_215,In_21);
and U337 (N_337,In_407,In_484);
nand U338 (N_338,In_706,In_169);
and U339 (N_339,In_210,In_482);
and U340 (N_340,In_327,In_652);
xnor U341 (N_341,In_271,In_685);
nand U342 (N_342,In_558,In_640);
or U343 (N_343,In_137,In_193);
nand U344 (N_344,In_723,In_697);
xnor U345 (N_345,In_488,In_523);
nand U346 (N_346,In_444,In_645);
and U347 (N_347,In_463,In_595);
nand U348 (N_348,In_542,In_746);
xnor U349 (N_349,In_86,In_277);
and U350 (N_350,In_582,In_374);
and U351 (N_351,In_715,In_379);
and U352 (N_352,In_662,In_493);
and U353 (N_353,In_48,In_243);
or U354 (N_354,In_312,In_395);
nor U355 (N_355,In_131,In_660);
nor U356 (N_356,In_276,In_554);
and U357 (N_357,In_151,In_733);
and U358 (N_358,In_41,In_184);
and U359 (N_359,In_579,In_569);
xor U360 (N_360,In_525,In_218);
or U361 (N_361,In_20,In_145);
and U362 (N_362,In_191,In_187);
nand U363 (N_363,In_38,In_615);
nor U364 (N_364,In_713,In_328);
or U365 (N_365,In_499,In_426);
or U366 (N_366,In_361,In_413);
nand U367 (N_367,In_6,In_473);
nor U368 (N_368,In_743,In_211);
xor U369 (N_369,In_553,In_679);
nand U370 (N_370,In_261,In_69);
or U371 (N_371,In_414,In_63);
nor U372 (N_372,In_494,In_578);
nor U373 (N_373,In_461,In_359);
xnor U374 (N_374,In_153,In_45);
nand U375 (N_375,In_347,In_634);
nand U376 (N_376,In_727,In_121);
nand U377 (N_377,In_515,In_241);
nor U378 (N_378,In_269,In_648);
and U379 (N_379,In_48,In_626);
and U380 (N_380,In_540,In_490);
and U381 (N_381,In_646,In_89);
nor U382 (N_382,In_237,In_372);
nor U383 (N_383,In_563,In_425);
or U384 (N_384,In_153,In_663);
or U385 (N_385,In_596,In_343);
and U386 (N_386,In_516,In_278);
nor U387 (N_387,In_232,In_600);
nand U388 (N_388,In_700,In_432);
or U389 (N_389,In_297,In_717);
nand U390 (N_390,In_53,In_216);
and U391 (N_391,In_573,In_339);
or U392 (N_392,In_215,In_398);
and U393 (N_393,In_225,In_611);
nand U394 (N_394,In_573,In_685);
or U395 (N_395,In_259,In_683);
nand U396 (N_396,In_105,In_168);
and U397 (N_397,In_725,In_3);
nor U398 (N_398,In_641,In_436);
xor U399 (N_399,In_679,In_110);
xnor U400 (N_400,In_453,In_621);
nand U401 (N_401,In_370,In_415);
nand U402 (N_402,In_643,In_572);
nor U403 (N_403,In_687,In_621);
or U404 (N_404,In_68,In_92);
xnor U405 (N_405,In_523,In_665);
or U406 (N_406,In_745,In_198);
or U407 (N_407,In_456,In_441);
xor U408 (N_408,In_584,In_151);
xor U409 (N_409,In_147,In_167);
nand U410 (N_410,In_40,In_216);
or U411 (N_411,In_71,In_677);
or U412 (N_412,In_19,In_88);
nor U413 (N_413,In_53,In_67);
nand U414 (N_414,In_369,In_637);
or U415 (N_415,In_79,In_185);
nand U416 (N_416,In_591,In_651);
xnor U417 (N_417,In_597,In_335);
and U418 (N_418,In_282,In_612);
nand U419 (N_419,In_490,In_331);
nor U420 (N_420,In_162,In_687);
nor U421 (N_421,In_106,In_519);
or U422 (N_422,In_183,In_407);
nor U423 (N_423,In_396,In_713);
nand U424 (N_424,In_179,In_738);
and U425 (N_425,In_553,In_149);
xor U426 (N_426,In_371,In_5);
nand U427 (N_427,In_566,In_43);
and U428 (N_428,In_183,In_529);
xnor U429 (N_429,In_280,In_451);
and U430 (N_430,In_195,In_435);
nand U431 (N_431,In_563,In_135);
or U432 (N_432,In_683,In_291);
nor U433 (N_433,In_689,In_298);
nor U434 (N_434,In_91,In_673);
xnor U435 (N_435,In_144,In_572);
or U436 (N_436,In_644,In_205);
or U437 (N_437,In_480,In_287);
and U438 (N_438,In_69,In_435);
xor U439 (N_439,In_561,In_263);
nand U440 (N_440,In_38,In_486);
xor U441 (N_441,In_573,In_658);
or U442 (N_442,In_313,In_409);
and U443 (N_443,In_703,In_612);
or U444 (N_444,In_272,In_130);
and U445 (N_445,In_589,In_58);
nor U446 (N_446,In_412,In_272);
nand U447 (N_447,In_8,In_658);
nand U448 (N_448,In_700,In_226);
or U449 (N_449,In_660,In_559);
or U450 (N_450,In_467,In_702);
nand U451 (N_451,In_343,In_378);
nand U452 (N_452,In_524,In_350);
or U453 (N_453,In_501,In_623);
and U454 (N_454,In_55,In_696);
and U455 (N_455,In_170,In_111);
and U456 (N_456,In_739,In_687);
or U457 (N_457,In_131,In_592);
nand U458 (N_458,In_376,In_437);
nor U459 (N_459,In_742,In_303);
nand U460 (N_460,In_494,In_557);
nor U461 (N_461,In_523,In_6);
nand U462 (N_462,In_569,In_89);
nand U463 (N_463,In_91,In_559);
and U464 (N_464,In_125,In_131);
xor U465 (N_465,In_5,In_108);
or U466 (N_466,In_466,In_657);
and U467 (N_467,In_349,In_572);
nand U468 (N_468,In_328,In_460);
nor U469 (N_469,In_461,In_306);
nand U470 (N_470,In_464,In_313);
nor U471 (N_471,In_9,In_93);
and U472 (N_472,In_11,In_642);
nand U473 (N_473,In_314,In_322);
nand U474 (N_474,In_722,In_729);
or U475 (N_475,In_432,In_167);
or U476 (N_476,In_295,In_666);
nand U477 (N_477,In_236,In_190);
or U478 (N_478,In_637,In_174);
nor U479 (N_479,In_400,In_24);
nand U480 (N_480,In_140,In_385);
nand U481 (N_481,In_246,In_541);
or U482 (N_482,In_360,In_362);
and U483 (N_483,In_45,In_246);
or U484 (N_484,In_11,In_499);
and U485 (N_485,In_233,In_334);
and U486 (N_486,In_637,In_167);
nor U487 (N_487,In_735,In_668);
nand U488 (N_488,In_257,In_719);
and U489 (N_489,In_282,In_428);
or U490 (N_490,In_420,In_88);
and U491 (N_491,In_171,In_647);
nor U492 (N_492,In_317,In_245);
or U493 (N_493,In_401,In_246);
nor U494 (N_494,In_12,In_244);
or U495 (N_495,In_317,In_241);
nor U496 (N_496,In_431,In_749);
nor U497 (N_497,In_236,In_381);
nor U498 (N_498,In_688,In_561);
nand U499 (N_499,In_688,In_659);
nand U500 (N_500,In_672,In_635);
or U501 (N_501,In_475,In_495);
and U502 (N_502,In_346,In_745);
nand U503 (N_503,In_601,In_434);
nor U504 (N_504,In_540,In_476);
xnor U505 (N_505,In_423,In_126);
and U506 (N_506,In_572,In_253);
nor U507 (N_507,In_274,In_288);
nand U508 (N_508,In_604,In_35);
or U509 (N_509,In_571,In_425);
nor U510 (N_510,In_98,In_314);
and U511 (N_511,In_660,In_282);
nand U512 (N_512,In_202,In_67);
nand U513 (N_513,In_18,In_301);
xor U514 (N_514,In_555,In_221);
nand U515 (N_515,In_7,In_565);
and U516 (N_516,In_642,In_194);
nand U517 (N_517,In_103,In_345);
nor U518 (N_518,In_464,In_675);
nand U519 (N_519,In_634,In_99);
and U520 (N_520,In_260,In_454);
nor U521 (N_521,In_722,In_701);
xnor U522 (N_522,In_685,In_39);
nor U523 (N_523,In_103,In_71);
nor U524 (N_524,In_667,In_13);
or U525 (N_525,In_549,In_370);
nor U526 (N_526,In_442,In_586);
and U527 (N_527,In_92,In_56);
xnor U528 (N_528,In_612,In_133);
nor U529 (N_529,In_615,In_537);
nand U530 (N_530,In_429,In_433);
and U531 (N_531,In_17,In_493);
or U532 (N_532,In_186,In_55);
xnor U533 (N_533,In_151,In_684);
or U534 (N_534,In_699,In_170);
nor U535 (N_535,In_172,In_26);
and U536 (N_536,In_425,In_633);
nand U537 (N_537,In_343,In_728);
and U538 (N_538,In_282,In_360);
xor U539 (N_539,In_149,In_334);
nand U540 (N_540,In_724,In_566);
nand U541 (N_541,In_121,In_435);
and U542 (N_542,In_622,In_220);
or U543 (N_543,In_674,In_299);
nand U544 (N_544,In_686,In_417);
or U545 (N_545,In_622,In_300);
nor U546 (N_546,In_306,In_485);
nand U547 (N_547,In_604,In_206);
nand U548 (N_548,In_118,In_242);
nand U549 (N_549,In_578,In_105);
nor U550 (N_550,In_49,In_222);
or U551 (N_551,In_78,In_546);
or U552 (N_552,In_300,In_695);
nor U553 (N_553,In_17,In_40);
xnor U554 (N_554,In_278,In_492);
nand U555 (N_555,In_388,In_311);
nor U556 (N_556,In_184,In_106);
xor U557 (N_557,In_283,In_395);
nor U558 (N_558,In_349,In_164);
or U559 (N_559,In_596,In_570);
xnor U560 (N_560,In_250,In_309);
or U561 (N_561,In_587,In_246);
nor U562 (N_562,In_265,In_726);
xnor U563 (N_563,In_580,In_151);
xor U564 (N_564,In_377,In_554);
nand U565 (N_565,In_204,In_725);
xnor U566 (N_566,In_418,In_170);
or U567 (N_567,In_457,In_46);
nor U568 (N_568,In_572,In_571);
or U569 (N_569,In_572,In_45);
or U570 (N_570,In_521,In_336);
xnor U571 (N_571,In_367,In_313);
nor U572 (N_572,In_567,In_503);
nor U573 (N_573,In_446,In_267);
nor U574 (N_574,In_572,In_161);
and U575 (N_575,In_354,In_388);
nor U576 (N_576,In_272,In_676);
nor U577 (N_577,In_543,In_8);
and U578 (N_578,In_283,In_101);
or U579 (N_579,In_416,In_96);
nor U580 (N_580,In_376,In_346);
nand U581 (N_581,In_13,In_577);
or U582 (N_582,In_484,In_33);
and U583 (N_583,In_511,In_421);
and U584 (N_584,In_72,In_57);
and U585 (N_585,In_544,In_378);
and U586 (N_586,In_57,In_575);
nor U587 (N_587,In_444,In_106);
nor U588 (N_588,In_742,In_171);
or U589 (N_589,In_440,In_62);
nand U590 (N_590,In_592,In_138);
nor U591 (N_591,In_725,In_517);
nand U592 (N_592,In_586,In_9);
and U593 (N_593,In_738,In_29);
and U594 (N_594,In_506,In_584);
nand U595 (N_595,In_354,In_356);
and U596 (N_596,In_282,In_593);
nand U597 (N_597,In_310,In_605);
and U598 (N_598,In_205,In_89);
or U599 (N_599,In_567,In_300);
nand U600 (N_600,In_276,In_256);
and U601 (N_601,In_286,In_414);
nor U602 (N_602,In_241,In_499);
nor U603 (N_603,In_93,In_580);
or U604 (N_604,In_327,In_541);
nor U605 (N_605,In_167,In_563);
or U606 (N_606,In_497,In_83);
nand U607 (N_607,In_531,In_294);
and U608 (N_608,In_302,In_20);
nor U609 (N_609,In_518,In_1);
and U610 (N_610,In_371,In_114);
and U611 (N_611,In_421,In_279);
nand U612 (N_612,In_502,In_674);
and U613 (N_613,In_367,In_736);
nor U614 (N_614,In_135,In_94);
nand U615 (N_615,In_602,In_596);
nand U616 (N_616,In_475,In_385);
nor U617 (N_617,In_467,In_723);
or U618 (N_618,In_213,In_529);
or U619 (N_619,In_431,In_712);
and U620 (N_620,In_478,In_143);
nand U621 (N_621,In_160,In_617);
or U622 (N_622,In_719,In_611);
nor U623 (N_623,In_657,In_519);
or U624 (N_624,In_284,In_664);
and U625 (N_625,In_370,In_743);
nand U626 (N_626,In_379,In_648);
nor U627 (N_627,In_19,In_124);
and U628 (N_628,In_179,In_174);
nor U629 (N_629,In_520,In_605);
nor U630 (N_630,In_498,In_428);
nor U631 (N_631,In_592,In_443);
nor U632 (N_632,In_534,In_323);
nor U633 (N_633,In_89,In_122);
nand U634 (N_634,In_252,In_633);
nor U635 (N_635,In_20,In_97);
or U636 (N_636,In_385,In_640);
nand U637 (N_637,In_381,In_163);
and U638 (N_638,In_367,In_106);
and U639 (N_639,In_695,In_65);
and U640 (N_640,In_527,In_742);
and U641 (N_641,In_577,In_138);
nor U642 (N_642,In_561,In_589);
or U643 (N_643,In_21,In_488);
and U644 (N_644,In_475,In_67);
nand U645 (N_645,In_703,In_706);
nand U646 (N_646,In_202,In_355);
nor U647 (N_647,In_435,In_78);
and U648 (N_648,In_436,In_290);
and U649 (N_649,In_695,In_211);
and U650 (N_650,In_193,In_147);
nor U651 (N_651,In_639,In_656);
and U652 (N_652,In_274,In_247);
and U653 (N_653,In_479,In_674);
and U654 (N_654,In_482,In_729);
xnor U655 (N_655,In_183,In_85);
nand U656 (N_656,In_663,In_716);
xnor U657 (N_657,In_614,In_134);
or U658 (N_658,In_176,In_451);
nor U659 (N_659,In_306,In_386);
nand U660 (N_660,In_485,In_325);
or U661 (N_661,In_708,In_147);
and U662 (N_662,In_282,In_449);
nand U663 (N_663,In_69,In_280);
and U664 (N_664,In_556,In_734);
or U665 (N_665,In_426,In_51);
nand U666 (N_666,In_617,In_631);
xnor U667 (N_667,In_454,In_717);
nor U668 (N_668,In_65,In_583);
xor U669 (N_669,In_43,In_75);
nand U670 (N_670,In_406,In_381);
nand U671 (N_671,In_691,In_190);
or U672 (N_672,In_499,In_379);
or U673 (N_673,In_604,In_308);
and U674 (N_674,In_537,In_154);
nand U675 (N_675,In_17,In_569);
xor U676 (N_676,In_674,In_346);
and U677 (N_677,In_729,In_547);
nor U678 (N_678,In_341,In_471);
nand U679 (N_679,In_184,In_40);
and U680 (N_680,In_680,In_259);
and U681 (N_681,In_475,In_662);
xnor U682 (N_682,In_458,In_740);
or U683 (N_683,In_499,In_484);
and U684 (N_684,In_558,In_689);
or U685 (N_685,In_20,In_151);
xor U686 (N_686,In_32,In_316);
or U687 (N_687,In_721,In_472);
nand U688 (N_688,In_199,In_450);
and U689 (N_689,In_368,In_518);
xnor U690 (N_690,In_88,In_261);
nand U691 (N_691,In_459,In_72);
nand U692 (N_692,In_405,In_380);
nor U693 (N_693,In_119,In_89);
xnor U694 (N_694,In_11,In_523);
and U695 (N_695,In_325,In_239);
nand U696 (N_696,In_631,In_209);
xnor U697 (N_697,In_140,In_13);
nor U698 (N_698,In_503,In_252);
and U699 (N_699,In_255,In_627);
nor U700 (N_700,In_387,In_242);
nand U701 (N_701,In_280,In_243);
nor U702 (N_702,In_702,In_390);
and U703 (N_703,In_321,In_372);
nand U704 (N_704,In_189,In_352);
xor U705 (N_705,In_158,In_463);
or U706 (N_706,In_319,In_372);
nor U707 (N_707,In_54,In_562);
and U708 (N_708,In_142,In_322);
nor U709 (N_709,In_384,In_710);
nand U710 (N_710,In_562,In_275);
xnor U711 (N_711,In_635,In_463);
nand U712 (N_712,In_481,In_9);
xor U713 (N_713,In_710,In_149);
and U714 (N_714,In_350,In_747);
xor U715 (N_715,In_175,In_414);
nand U716 (N_716,In_597,In_505);
nor U717 (N_717,In_668,In_507);
nor U718 (N_718,In_572,In_706);
or U719 (N_719,In_477,In_648);
nand U720 (N_720,In_137,In_239);
or U721 (N_721,In_682,In_17);
nor U722 (N_722,In_608,In_712);
or U723 (N_723,In_284,In_586);
xnor U724 (N_724,In_664,In_105);
nand U725 (N_725,In_746,In_105);
nor U726 (N_726,In_747,In_645);
nor U727 (N_727,In_176,In_409);
xor U728 (N_728,In_302,In_445);
nand U729 (N_729,In_305,In_321);
nor U730 (N_730,In_694,In_499);
or U731 (N_731,In_575,In_109);
or U732 (N_732,In_195,In_579);
nor U733 (N_733,In_729,In_576);
or U734 (N_734,In_490,In_24);
nor U735 (N_735,In_94,In_286);
nand U736 (N_736,In_743,In_282);
nor U737 (N_737,In_589,In_47);
nand U738 (N_738,In_316,In_181);
or U739 (N_739,In_340,In_723);
nor U740 (N_740,In_706,In_241);
nand U741 (N_741,In_369,In_306);
and U742 (N_742,In_153,In_368);
or U743 (N_743,In_703,In_233);
or U744 (N_744,In_643,In_258);
nand U745 (N_745,In_176,In_534);
or U746 (N_746,In_426,In_36);
and U747 (N_747,In_622,In_436);
nor U748 (N_748,In_731,In_581);
nand U749 (N_749,In_290,In_618);
nor U750 (N_750,In_11,In_91);
xor U751 (N_751,In_150,In_61);
and U752 (N_752,In_654,In_605);
and U753 (N_753,In_443,In_486);
and U754 (N_754,In_586,In_731);
xnor U755 (N_755,In_608,In_442);
xor U756 (N_756,In_332,In_675);
or U757 (N_757,In_531,In_662);
or U758 (N_758,In_324,In_109);
nand U759 (N_759,In_377,In_215);
and U760 (N_760,In_68,In_428);
and U761 (N_761,In_414,In_94);
and U762 (N_762,In_535,In_190);
xor U763 (N_763,In_397,In_76);
xnor U764 (N_764,In_660,In_335);
nand U765 (N_765,In_563,In_520);
or U766 (N_766,In_301,In_648);
and U767 (N_767,In_185,In_2);
nor U768 (N_768,In_629,In_1);
nor U769 (N_769,In_478,In_404);
nor U770 (N_770,In_309,In_226);
nor U771 (N_771,In_504,In_42);
xor U772 (N_772,In_253,In_167);
nand U773 (N_773,In_504,In_476);
nor U774 (N_774,In_518,In_360);
or U775 (N_775,In_555,In_140);
or U776 (N_776,In_323,In_488);
nor U777 (N_777,In_6,In_107);
and U778 (N_778,In_443,In_17);
nor U779 (N_779,In_455,In_411);
and U780 (N_780,In_226,In_290);
nor U781 (N_781,In_358,In_462);
nor U782 (N_782,In_332,In_323);
nor U783 (N_783,In_392,In_419);
nand U784 (N_784,In_253,In_175);
nand U785 (N_785,In_351,In_710);
and U786 (N_786,In_574,In_456);
and U787 (N_787,In_611,In_227);
and U788 (N_788,In_485,In_20);
and U789 (N_789,In_434,In_397);
or U790 (N_790,In_430,In_568);
nand U791 (N_791,In_97,In_573);
nor U792 (N_792,In_217,In_617);
xor U793 (N_793,In_63,In_614);
xor U794 (N_794,In_560,In_361);
and U795 (N_795,In_498,In_100);
and U796 (N_796,In_210,In_452);
and U797 (N_797,In_280,In_230);
and U798 (N_798,In_595,In_262);
nand U799 (N_799,In_700,In_680);
nor U800 (N_800,In_261,In_231);
and U801 (N_801,In_417,In_373);
nand U802 (N_802,In_727,In_431);
and U803 (N_803,In_336,In_164);
nand U804 (N_804,In_633,In_87);
or U805 (N_805,In_495,In_260);
and U806 (N_806,In_426,In_460);
nand U807 (N_807,In_433,In_527);
and U808 (N_808,In_370,In_44);
xnor U809 (N_809,In_448,In_238);
or U810 (N_810,In_347,In_397);
nor U811 (N_811,In_139,In_644);
nand U812 (N_812,In_167,In_281);
and U813 (N_813,In_572,In_398);
or U814 (N_814,In_551,In_498);
nand U815 (N_815,In_402,In_422);
and U816 (N_816,In_211,In_712);
nor U817 (N_817,In_183,In_241);
nor U818 (N_818,In_116,In_126);
nand U819 (N_819,In_722,In_178);
nor U820 (N_820,In_499,In_743);
xor U821 (N_821,In_738,In_557);
and U822 (N_822,In_56,In_579);
or U823 (N_823,In_443,In_252);
or U824 (N_824,In_369,In_495);
or U825 (N_825,In_703,In_67);
or U826 (N_826,In_386,In_185);
nand U827 (N_827,In_619,In_185);
or U828 (N_828,In_660,In_625);
nor U829 (N_829,In_664,In_440);
and U830 (N_830,In_408,In_349);
and U831 (N_831,In_458,In_700);
or U832 (N_832,In_510,In_597);
or U833 (N_833,In_659,In_362);
and U834 (N_834,In_653,In_599);
nand U835 (N_835,In_679,In_405);
and U836 (N_836,In_148,In_412);
nand U837 (N_837,In_723,In_7);
nor U838 (N_838,In_279,In_566);
nand U839 (N_839,In_343,In_230);
nor U840 (N_840,In_526,In_605);
nor U841 (N_841,In_170,In_348);
or U842 (N_842,In_513,In_166);
nor U843 (N_843,In_214,In_714);
nor U844 (N_844,In_30,In_536);
nor U845 (N_845,In_265,In_50);
nand U846 (N_846,In_214,In_310);
and U847 (N_847,In_547,In_473);
nor U848 (N_848,In_142,In_362);
xnor U849 (N_849,In_165,In_591);
and U850 (N_850,In_738,In_150);
xnor U851 (N_851,In_443,In_132);
or U852 (N_852,In_495,In_81);
or U853 (N_853,In_384,In_172);
or U854 (N_854,In_130,In_612);
nand U855 (N_855,In_521,In_17);
or U856 (N_856,In_541,In_488);
nor U857 (N_857,In_729,In_221);
xor U858 (N_858,In_653,In_370);
nor U859 (N_859,In_83,In_648);
xor U860 (N_860,In_63,In_302);
nand U861 (N_861,In_295,In_464);
or U862 (N_862,In_264,In_3);
and U863 (N_863,In_388,In_239);
and U864 (N_864,In_278,In_183);
or U865 (N_865,In_452,In_749);
xnor U866 (N_866,In_290,In_118);
nor U867 (N_867,In_50,In_6);
and U868 (N_868,In_550,In_153);
and U869 (N_869,In_341,In_567);
and U870 (N_870,In_238,In_103);
nor U871 (N_871,In_389,In_508);
or U872 (N_872,In_97,In_367);
nand U873 (N_873,In_98,In_330);
xor U874 (N_874,In_264,In_78);
and U875 (N_875,In_408,In_559);
and U876 (N_876,In_510,In_270);
nand U877 (N_877,In_316,In_200);
nand U878 (N_878,In_453,In_661);
xnor U879 (N_879,In_159,In_741);
and U880 (N_880,In_748,In_137);
nor U881 (N_881,In_543,In_214);
and U882 (N_882,In_333,In_345);
nand U883 (N_883,In_305,In_482);
nor U884 (N_884,In_544,In_213);
nand U885 (N_885,In_323,In_267);
and U886 (N_886,In_381,In_611);
nand U887 (N_887,In_400,In_267);
nand U888 (N_888,In_493,In_519);
or U889 (N_889,In_350,In_365);
or U890 (N_890,In_376,In_101);
xnor U891 (N_891,In_345,In_734);
nand U892 (N_892,In_135,In_47);
nor U893 (N_893,In_472,In_625);
and U894 (N_894,In_709,In_718);
nand U895 (N_895,In_172,In_178);
and U896 (N_896,In_404,In_190);
or U897 (N_897,In_373,In_707);
or U898 (N_898,In_644,In_182);
nor U899 (N_899,In_49,In_2);
and U900 (N_900,In_578,In_462);
or U901 (N_901,In_24,In_423);
nor U902 (N_902,In_331,In_68);
or U903 (N_903,In_673,In_121);
nand U904 (N_904,In_151,In_381);
nand U905 (N_905,In_567,In_590);
or U906 (N_906,In_113,In_64);
nand U907 (N_907,In_45,In_693);
nor U908 (N_908,In_393,In_32);
nor U909 (N_909,In_592,In_23);
nor U910 (N_910,In_476,In_352);
and U911 (N_911,In_668,In_181);
nor U912 (N_912,In_556,In_296);
nand U913 (N_913,In_155,In_286);
and U914 (N_914,In_401,In_541);
nand U915 (N_915,In_86,In_316);
or U916 (N_916,In_572,In_211);
nor U917 (N_917,In_602,In_446);
nor U918 (N_918,In_266,In_180);
nand U919 (N_919,In_456,In_632);
nor U920 (N_920,In_588,In_532);
and U921 (N_921,In_689,In_268);
xor U922 (N_922,In_124,In_499);
nor U923 (N_923,In_629,In_654);
or U924 (N_924,In_691,In_157);
nor U925 (N_925,In_86,In_514);
and U926 (N_926,In_93,In_136);
nor U927 (N_927,In_319,In_286);
nor U928 (N_928,In_638,In_32);
nor U929 (N_929,In_630,In_717);
and U930 (N_930,In_594,In_394);
nor U931 (N_931,In_250,In_610);
nor U932 (N_932,In_454,In_149);
and U933 (N_933,In_85,In_524);
nand U934 (N_934,In_745,In_411);
nand U935 (N_935,In_725,In_359);
or U936 (N_936,In_444,In_350);
or U937 (N_937,In_155,In_396);
nor U938 (N_938,In_116,In_170);
nand U939 (N_939,In_598,In_476);
nor U940 (N_940,In_290,In_306);
or U941 (N_941,In_37,In_66);
and U942 (N_942,In_599,In_407);
or U943 (N_943,In_498,In_430);
nor U944 (N_944,In_488,In_709);
nand U945 (N_945,In_748,In_253);
and U946 (N_946,In_376,In_583);
xnor U947 (N_947,In_40,In_514);
and U948 (N_948,In_150,In_20);
or U949 (N_949,In_117,In_65);
nor U950 (N_950,In_99,In_395);
nand U951 (N_951,In_295,In_401);
or U952 (N_952,In_589,In_464);
or U953 (N_953,In_681,In_465);
or U954 (N_954,In_231,In_639);
or U955 (N_955,In_579,In_742);
or U956 (N_956,In_704,In_655);
xnor U957 (N_957,In_656,In_107);
nor U958 (N_958,In_89,In_193);
or U959 (N_959,In_396,In_366);
xnor U960 (N_960,In_29,In_659);
xor U961 (N_961,In_342,In_334);
or U962 (N_962,In_4,In_637);
nor U963 (N_963,In_139,In_80);
xor U964 (N_964,In_655,In_300);
nand U965 (N_965,In_409,In_598);
nand U966 (N_966,In_118,In_283);
and U967 (N_967,In_111,In_369);
nor U968 (N_968,In_598,In_639);
nor U969 (N_969,In_632,In_26);
nor U970 (N_970,In_297,In_480);
and U971 (N_971,In_707,In_694);
nand U972 (N_972,In_77,In_158);
nand U973 (N_973,In_582,In_371);
and U974 (N_974,In_601,In_247);
nand U975 (N_975,In_371,In_639);
nor U976 (N_976,In_650,In_511);
nor U977 (N_977,In_65,In_429);
or U978 (N_978,In_164,In_293);
and U979 (N_979,In_520,In_18);
and U980 (N_980,In_200,In_663);
xnor U981 (N_981,In_692,In_37);
and U982 (N_982,In_389,In_544);
and U983 (N_983,In_155,In_405);
nor U984 (N_984,In_362,In_286);
nand U985 (N_985,In_378,In_574);
nor U986 (N_986,In_252,In_650);
nor U987 (N_987,In_511,In_273);
and U988 (N_988,In_171,In_70);
nand U989 (N_989,In_81,In_561);
and U990 (N_990,In_518,In_341);
nor U991 (N_991,In_351,In_144);
and U992 (N_992,In_72,In_369);
nand U993 (N_993,In_516,In_183);
nor U994 (N_994,In_307,In_411);
or U995 (N_995,In_727,In_567);
nand U996 (N_996,In_695,In_590);
and U997 (N_997,In_573,In_239);
nand U998 (N_998,In_284,In_566);
nor U999 (N_999,In_159,In_177);
xnor U1000 (N_1000,N_466,N_104);
nand U1001 (N_1001,N_877,N_858);
xor U1002 (N_1002,N_584,N_324);
and U1003 (N_1003,N_248,N_317);
and U1004 (N_1004,N_538,N_9);
or U1005 (N_1005,N_790,N_894);
nor U1006 (N_1006,N_167,N_788);
xor U1007 (N_1007,N_920,N_10);
and U1008 (N_1008,N_614,N_767);
nand U1009 (N_1009,N_604,N_744);
and U1010 (N_1010,N_683,N_859);
nand U1011 (N_1011,N_738,N_183);
or U1012 (N_1012,N_840,N_350);
nand U1013 (N_1013,N_14,N_641);
and U1014 (N_1014,N_161,N_616);
or U1015 (N_1015,N_133,N_694);
and U1016 (N_1016,N_776,N_356);
nand U1017 (N_1017,N_366,N_217);
or U1018 (N_1018,N_897,N_433);
nor U1019 (N_1019,N_743,N_745);
and U1020 (N_1020,N_841,N_158);
nor U1021 (N_1021,N_799,N_832);
nor U1022 (N_1022,N_652,N_467);
and U1023 (N_1023,N_32,N_51);
and U1024 (N_1024,N_27,N_146);
nand U1025 (N_1025,N_59,N_68);
nand U1026 (N_1026,N_885,N_239);
nand U1027 (N_1027,N_477,N_876);
or U1028 (N_1028,N_479,N_657);
nand U1029 (N_1029,N_670,N_564);
and U1030 (N_1030,N_560,N_934);
nand U1031 (N_1031,N_110,N_638);
and U1032 (N_1032,N_322,N_570);
nand U1033 (N_1033,N_706,N_160);
and U1034 (N_1034,N_275,N_251);
nand U1035 (N_1035,N_7,N_634);
or U1036 (N_1036,N_144,N_709);
nand U1037 (N_1037,N_880,N_524);
nor U1038 (N_1038,N_819,N_782);
nor U1039 (N_1039,N_296,N_320);
nand U1040 (N_1040,N_891,N_949);
and U1041 (N_1041,N_105,N_688);
nand U1042 (N_1042,N_729,N_932);
and U1043 (N_1043,N_310,N_583);
or U1044 (N_1044,N_974,N_884);
and U1045 (N_1045,N_504,N_265);
or U1046 (N_1046,N_807,N_287);
nand U1047 (N_1047,N_510,N_730);
nand U1048 (N_1048,N_966,N_390);
nand U1049 (N_1049,N_689,N_74);
and U1050 (N_1050,N_123,N_778);
and U1051 (N_1051,N_842,N_406);
or U1052 (N_1052,N_243,N_575);
nor U1053 (N_1053,N_644,N_16);
nor U1054 (N_1054,N_758,N_921);
nor U1055 (N_1055,N_441,N_553);
xnor U1056 (N_1056,N_215,N_847);
or U1057 (N_1057,N_773,N_574);
nor U1058 (N_1058,N_209,N_806);
and U1059 (N_1059,N_326,N_337);
nor U1060 (N_1060,N_501,N_623);
nor U1061 (N_1061,N_855,N_572);
or U1062 (N_1062,N_976,N_514);
nand U1063 (N_1063,N_517,N_12);
and U1064 (N_1064,N_454,N_761);
and U1065 (N_1065,N_965,N_896);
nand U1066 (N_1066,N_672,N_389);
or U1067 (N_1067,N_409,N_973);
nand U1068 (N_1068,N_78,N_810);
or U1069 (N_1069,N_618,N_901);
or U1070 (N_1070,N_230,N_591);
xor U1071 (N_1071,N_967,N_667);
nand U1072 (N_1072,N_888,N_463);
xnor U1073 (N_1073,N_686,N_386);
or U1074 (N_1074,N_978,N_804);
or U1075 (N_1075,N_168,N_281);
and U1076 (N_1076,N_696,N_165);
nor U1077 (N_1077,N_526,N_132);
or U1078 (N_1078,N_475,N_291);
nor U1079 (N_1079,N_330,N_443);
and U1080 (N_1080,N_771,N_802);
and U1081 (N_1081,N_297,N_292);
and U1082 (N_1082,N_61,N_923);
nor U1083 (N_1083,N_756,N_969);
or U1084 (N_1084,N_38,N_55);
or U1085 (N_1085,N_252,N_627);
nand U1086 (N_1086,N_30,N_660);
nor U1087 (N_1087,N_376,N_836);
nand U1088 (N_1088,N_953,N_49);
and U1089 (N_1089,N_54,N_786);
nor U1090 (N_1090,N_726,N_4);
or U1091 (N_1091,N_380,N_601);
nand U1092 (N_1092,N_299,N_813);
and U1093 (N_1093,N_935,N_502);
and U1094 (N_1094,N_527,N_218);
xnor U1095 (N_1095,N_88,N_182);
nand U1096 (N_1096,N_882,N_692);
or U1097 (N_1097,N_590,N_610);
nand U1098 (N_1098,N_750,N_752);
nand U1099 (N_1099,N_302,N_425);
or U1100 (N_1100,N_668,N_404);
nand U1101 (N_1101,N_582,N_488);
nand U1102 (N_1102,N_163,N_300);
and U1103 (N_1103,N_201,N_731);
or U1104 (N_1104,N_342,N_81);
nor U1105 (N_1105,N_86,N_474);
nor U1106 (N_1106,N_747,N_860);
or U1107 (N_1107,N_753,N_64);
xor U1108 (N_1108,N_343,N_60);
nand U1109 (N_1109,N_795,N_67);
nand U1110 (N_1110,N_863,N_805);
or U1111 (N_1111,N_955,N_988);
nor U1112 (N_1112,N_844,N_2);
nor U1113 (N_1113,N_116,N_924);
nor U1114 (N_1114,N_846,N_147);
or U1115 (N_1115,N_185,N_196);
or U1116 (N_1116,N_25,N_437);
xor U1117 (N_1117,N_46,N_41);
nand U1118 (N_1118,N_315,N_108);
nand U1119 (N_1119,N_312,N_496);
nor U1120 (N_1120,N_453,N_303);
or U1121 (N_1121,N_367,N_448);
nor U1122 (N_1122,N_140,N_725);
nor U1123 (N_1123,N_58,N_370);
nor U1124 (N_1124,N_371,N_930);
nor U1125 (N_1125,N_495,N_336);
or U1126 (N_1126,N_940,N_255);
nand U1127 (N_1127,N_199,N_621);
nand U1128 (N_1128,N_344,N_981);
nand U1129 (N_1129,N_349,N_276);
nor U1130 (N_1130,N_485,N_830);
nand U1131 (N_1131,N_794,N_698);
nand U1132 (N_1132,N_868,N_760);
or U1133 (N_1133,N_650,N_159);
and U1134 (N_1134,N_914,N_415);
nor U1135 (N_1135,N_798,N_115);
or U1136 (N_1136,N_869,N_279);
nand U1137 (N_1137,N_62,N_763);
xor U1138 (N_1138,N_557,N_831);
nor U1139 (N_1139,N_879,N_498);
xnor U1140 (N_1140,N_261,N_325);
nand U1141 (N_1141,N_613,N_234);
nand U1142 (N_1142,N_91,N_272);
or U1143 (N_1143,N_647,N_908);
and U1144 (N_1144,N_142,N_164);
nor U1145 (N_1145,N_203,N_693);
or U1146 (N_1146,N_664,N_284);
nand U1147 (N_1147,N_340,N_681);
nand U1148 (N_1148,N_460,N_509);
nand U1149 (N_1149,N_338,N_961);
nand U1150 (N_1150,N_679,N_33);
or U1151 (N_1151,N_461,N_331);
and U1152 (N_1152,N_493,N_233);
and U1153 (N_1153,N_399,N_121);
nand U1154 (N_1154,N_23,N_742);
nand U1155 (N_1155,N_143,N_515);
and U1156 (N_1156,N_103,N_837);
or U1157 (N_1157,N_241,N_952);
and U1158 (N_1158,N_224,N_907);
or U1159 (N_1159,N_552,N_216);
and U1160 (N_1160,N_355,N_434);
xnor U1161 (N_1161,N_112,N_89);
or U1162 (N_1162,N_52,N_536);
nor U1163 (N_1163,N_705,N_665);
nand U1164 (N_1164,N_918,N_449);
nand U1165 (N_1165,N_17,N_669);
and U1166 (N_1166,N_362,N_414);
or U1167 (N_1167,N_954,N_202);
nor U1168 (N_1168,N_700,N_676);
or U1169 (N_1169,N_1,N_962);
nor U1170 (N_1170,N_633,N_178);
nand U1171 (N_1171,N_643,N_93);
or U1172 (N_1172,N_24,N_600);
nor U1173 (N_1173,N_438,N_492);
nand U1174 (N_1174,N_436,N_977);
or U1175 (N_1175,N_569,N_0);
nor U1176 (N_1176,N_851,N_191);
nor U1177 (N_1177,N_608,N_662);
and U1178 (N_1178,N_379,N_958);
nor U1179 (N_1179,N_779,N_938);
nor U1180 (N_1180,N_6,N_917);
nand U1181 (N_1181,N_648,N_179);
nor U1182 (N_1182,N_581,N_781);
or U1183 (N_1183,N_120,N_939);
nand U1184 (N_1184,N_586,N_598);
or U1185 (N_1185,N_695,N_603);
nand U1186 (N_1186,N_153,N_173);
nand U1187 (N_1187,N_549,N_459);
nor U1188 (N_1188,N_174,N_566);
and U1189 (N_1189,N_780,N_546);
nor U1190 (N_1190,N_188,N_358);
nor U1191 (N_1191,N_473,N_889);
nand U1192 (N_1192,N_341,N_875);
nand U1193 (N_1193,N_521,N_152);
xnor U1194 (N_1194,N_100,N_381);
nand U1195 (N_1195,N_413,N_701);
nand U1196 (N_1196,N_469,N_345);
and U1197 (N_1197,N_484,N_393);
and U1198 (N_1198,N_150,N_190);
nor U1199 (N_1199,N_50,N_220);
nor U1200 (N_1200,N_928,N_411);
or U1201 (N_1201,N_470,N_937);
xor U1202 (N_1202,N_204,N_687);
and U1203 (N_1203,N_361,N_391);
nor U1204 (N_1204,N_445,N_135);
or U1205 (N_1205,N_294,N_36);
nor U1206 (N_1206,N_503,N_214);
and U1207 (N_1207,N_378,N_571);
or U1208 (N_1208,N_431,N_711);
or U1209 (N_1209,N_480,N_192);
and U1210 (N_1210,N_262,N_775);
nand U1211 (N_1211,N_124,N_993);
and U1212 (N_1212,N_594,N_442);
nor U1213 (N_1213,N_177,N_733);
nand U1214 (N_1214,N_593,N_432);
or U1215 (N_1215,N_290,N_533);
nor U1216 (N_1216,N_871,N_96);
nor U1217 (N_1217,N_339,N_332);
xor U1218 (N_1218,N_826,N_768);
and U1219 (N_1219,N_348,N_931);
nand U1220 (N_1220,N_374,N_316);
or U1221 (N_1221,N_606,N_865);
or U1222 (N_1222,N_22,N_267);
nand U1223 (N_1223,N_987,N_360);
nand U1224 (N_1224,N_746,N_945);
nor U1225 (N_1225,N_559,N_645);
nand U1226 (N_1226,N_690,N_646);
xnor U1227 (N_1227,N_114,N_346);
nand U1228 (N_1228,N_785,N_456);
and U1229 (N_1229,N_53,N_718);
nor U1230 (N_1230,N_223,N_968);
or U1231 (N_1231,N_180,N_511);
nand U1232 (N_1232,N_853,N_856);
or U1233 (N_1233,N_890,N_979);
and U1234 (N_1234,N_365,N_151);
or U1235 (N_1235,N_403,N_95);
or U1236 (N_1236,N_713,N_715);
xor U1237 (N_1237,N_430,N_991);
xnor U1238 (N_1238,N_671,N_548);
nand U1239 (N_1239,N_109,N_8);
nand U1240 (N_1240,N_673,N_44);
nor U1241 (N_1241,N_465,N_472);
nor U1242 (N_1242,N_71,N_866);
xnor U1243 (N_1243,N_857,N_83);
or U1244 (N_1244,N_892,N_257);
nor U1245 (N_1245,N_809,N_225);
or U1246 (N_1246,N_149,N_423);
and U1247 (N_1247,N_800,N_900);
or U1248 (N_1248,N_568,N_812);
xnor U1249 (N_1249,N_169,N_424);
nor U1250 (N_1250,N_471,N_893);
and U1251 (N_1251,N_999,N_678);
and U1252 (N_1252,N_351,N_626);
or U1253 (N_1253,N_208,N_410);
nor U1254 (N_1254,N_545,N_285);
or U1255 (N_1255,N_596,N_491);
nor U1256 (N_1256,N_998,N_400);
and U1257 (N_1257,N_102,N_237);
or U1258 (N_1258,N_427,N_301);
and U1259 (N_1259,N_905,N_499);
or U1260 (N_1260,N_588,N_682);
or U1261 (N_1261,N_770,N_555);
xor U1262 (N_1262,N_845,N_986);
or U1263 (N_1263,N_21,N_578);
or U1264 (N_1264,N_323,N_254);
or U1265 (N_1265,N_304,N_661);
nor U1266 (N_1266,N_872,N_653);
or U1267 (N_1267,N_57,N_561);
nand U1268 (N_1268,N_922,N_567);
or U1269 (N_1269,N_929,N_490);
xnor U1270 (N_1270,N_605,N_597);
and U1271 (N_1271,N_925,N_226);
and U1272 (N_1272,N_659,N_273);
or U1273 (N_1273,N_874,N_867);
or U1274 (N_1274,N_630,N_959);
nand U1275 (N_1275,N_772,N_629);
xor U1276 (N_1276,N_505,N_373);
nand U1277 (N_1277,N_808,N_79);
and U1278 (N_1278,N_915,N_306);
nor U1279 (N_1279,N_244,N_784);
nor U1280 (N_1280,N_573,N_523);
nor U1281 (N_1281,N_268,N_684);
nand U1282 (N_1282,N_117,N_43);
nand U1283 (N_1283,N_801,N_862);
xor U1284 (N_1284,N_446,N_126);
nand U1285 (N_1285,N_394,N_75);
nand U1286 (N_1286,N_211,N_213);
nand U1287 (N_1287,N_422,N_704);
or U1288 (N_1288,N_429,N_625);
nor U1289 (N_1289,N_850,N_904);
xor U1290 (N_1290,N_912,N_383);
nand U1291 (N_1291,N_375,N_451);
nor U1292 (N_1292,N_899,N_293);
and U1293 (N_1293,N_944,N_843);
nor U1294 (N_1294,N_184,N_269);
and U1295 (N_1295,N_654,N_195);
and U1296 (N_1296,N_487,N_642);
nor U1297 (N_1297,N_984,N_270);
nand U1298 (N_1298,N_65,N_820);
nand U1299 (N_1299,N_947,N_996);
and U1300 (N_1300,N_395,N_861);
nor U1301 (N_1301,N_878,N_118);
nor U1302 (N_1302,N_397,N_82);
nand U1303 (N_1303,N_516,N_864);
nor U1304 (N_1304,N_823,N_535);
or U1305 (N_1305,N_817,N_881);
or U1306 (N_1306,N_421,N_739);
nand U1307 (N_1307,N_540,N_525);
or U1308 (N_1308,N_834,N_428);
or U1309 (N_1309,N_387,N_960);
xor U1310 (N_1310,N_541,N_3);
nor U1311 (N_1311,N_353,N_766);
xor U1312 (N_1312,N_455,N_227);
xor U1313 (N_1313,N_417,N_816);
nor U1314 (N_1314,N_15,N_699);
or U1315 (N_1315,N_171,N_87);
nor U1316 (N_1316,N_727,N_119);
nor U1317 (N_1317,N_550,N_335);
and U1318 (N_1318,N_611,N_822);
nand U1319 (N_1319,N_580,N_895);
nand U1320 (N_1320,N_392,N_482);
xnor U1321 (N_1321,N_250,N_92);
xnor U1322 (N_1322,N_728,N_481);
or U1323 (N_1323,N_274,N_507);
nand U1324 (N_1324,N_827,N_278);
and U1325 (N_1325,N_995,N_754);
nor U1326 (N_1326,N_266,N_90);
nor U1327 (N_1327,N_228,N_762);
and U1328 (N_1328,N_18,N_200);
nor U1329 (N_1329,N_186,N_249);
nor U1330 (N_1330,N_280,N_520);
or U1331 (N_1331,N_352,N_612);
or U1332 (N_1332,N_839,N_619);
xnor U1333 (N_1333,N_385,N_631);
nand U1334 (N_1334,N_757,N_941);
nor U1335 (N_1335,N_926,N_364);
and U1336 (N_1336,N_854,N_764);
and U1337 (N_1337,N_368,N_458);
or U1338 (N_1338,N_136,N_898);
nand U1339 (N_1339,N_263,N_447);
xor U1340 (N_1340,N_289,N_222);
nand U1341 (N_1341,N_655,N_295);
and U1342 (N_1342,N_811,N_85);
xnor U1343 (N_1343,N_288,N_137);
and U1344 (N_1344,N_283,N_909);
nand U1345 (N_1345,N_970,N_412);
or U1346 (N_1346,N_628,N_777);
nor U1347 (N_1347,N_334,N_194);
nand U1348 (N_1348,N_989,N_635);
or U1349 (N_1349,N_131,N_401);
or U1350 (N_1350,N_791,N_259);
nand U1351 (N_1351,N_680,N_500);
nor U1352 (N_1352,N_416,N_565);
nor U1353 (N_1353,N_129,N_755);
and U1354 (N_1354,N_717,N_483);
nor U1355 (N_1355,N_253,N_408);
or U1356 (N_1356,N_537,N_5);
nand U1357 (N_1357,N_637,N_723);
and U1358 (N_1358,N_741,N_814);
nor U1359 (N_1359,N_797,N_796);
nor U1360 (N_1360,N_286,N_489);
nand U1361 (N_1361,N_789,N_522);
and U1362 (N_1362,N_37,N_592);
and U1363 (N_1363,N_11,N_702);
nand U1364 (N_1364,N_542,N_77);
nand U1365 (N_1365,N_157,N_997);
nor U1366 (N_1366,N_369,N_585);
xor U1367 (N_1367,N_906,N_26);
nor U1368 (N_1368,N_240,N_632);
or U1369 (N_1369,N_155,N_236);
and U1370 (N_1370,N_388,N_321);
and U1371 (N_1371,N_111,N_734);
nor U1372 (N_1372,N_554,N_838);
or U1373 (N_1373,N_452,N_319);
or U1374 (N_1374,N_219,N_707);
nand U1375 (N_1375,N_402,N_913);
nand U1376 (N_1376,N_198,N_130);
or U1377 (N_1377,N_181,N_19);
nand U1378 (N_1378,N_205,N_691);
and U1379 (N_1379,N_982,N_587);
nand U1380 (N_1380,N_99,N_439);
nand U1381 (N_1381,N_506,N_35);
and U1382 (N_1382,N_712,N_94);
and U1383 (N_1383,N_80,N_210);
and U1384 (N_1384,N_235,N_282);
or U1385 (N_1385,N_615,N_34);
or U1386 (N_1386,N_736,N_551);
or U1387 (N_1387,N_308,N_873);
nor U1388 (N_1388,N_708,N_426);
nor U1389 (N_1389,N_478,N_29);
and U1390 (N_1390,N_141,N_547);
nor U1391 (N_1391,N_848,N_724);
or U1392 (N_1392,N_663,N_639);
or U1393 (N_1393,N_494,N_229);
nor U1394 (N_1394,N_72,N_207);
nand U1395 (N_1395,N_419,N_956);
xor U1396 (N_1396,N_42,N_197);
nand U1397 (N_1397,N_333,N_936);
or U1398 (N_1398,N_983,N_309);
nand U1399 (N_1399,N_48,N_539);
and U1400 (N_1400,N_792,N_769);
and U1401 (N_1401,N_45,N_543);
and U1402 (N_1402,N_902,N_911);
and U1403 (N_1403,N_529,N_531);
or U1404 (N_1404,N_476,N_793);
nor U1405 (N_1405,N_113,N_148);
and U1406 (N_1406,N_73,N_607);
and U1407 (N_1407,N_833,N_589);
nor U1408 (N_1408,N_307,N_457);
nor U1409 (N_1409,N_990,N_787);
nand U1410 (N_1410,N_311,N_530);
nand U1411 (N_1411,N_579,N_189);
and U1412 (N_1412,N_162,N_824);
nand U1413 (N_1413,N_363,N_714);
nand U1414 (N_1414,N_577,N_740);
and U1415 (N_1415,N_563,N_719);
nor U1416 (N_1416,N_145,N_260);
and U1417 (N_1417,N_508,N_450);
nand U1418 (N_1418,N_245,N_398);
nor U1419 (N_1419,N_624,N_258);
or U1420 (N_1420,N_595,N_84);
nand U1421 (N_1421,N_951,N_238);
and U1422 (N_1422,N_435,N_154);
nand U1423 (N_1423,N_532,N_97);
and U1424 (N_1424,N_994,N_697);
xnor U1425 (N_1425,N_13,N_405);
nand U1426 (N_1426,N_948,N_674);
nor U1427 (N_1427,N_464,N_685);
nand U1428 (N_1428,N_518,N_134);
and U1429 (N_1429,N_101,N_318);
nand U1430 (N_1430,N_640,N_829);
or U1431 (N_1431,N_328,N_242);
nand U1432 (N_1432,N_576,N_964);
and U1433 (N_1433,N_127,N_852);
nand U1434 (N_1434,N_327,N_206);
and U1435 (N_1435,N_818,N_396);
xnor U1436 (N_1436,N_815,N_382);
or U1437 (N_1437,N_440,N_828);
nor U1438 (N_1438,N_675,N_39);
and U1439 (N_1439,N_957,N_710);
nor U1440 (N_1440,N_128,N_359);
and U1441 (N_1441,N_849,N_31);
nor U1442 (N_1442,N_468,N_649);
nor U1443 (N_1443,N_246,N_651);
and U1444 (N_1444,N_910,N_950);
or U1445 (N_1445,N_20,N_602);
or U1446 (N_1446,N_166,N_722);
or U1447 (N_1447,N_992,N_329);
nor U1448 (N_1448,N_212,N_264);
nor U1449 (N_1449,N_903,N_887);
nor U1450 (N_1450,N_122,N_751);
nand U1451 (N_1451,N_63,N_963);
nor U1452 (N_1452,N_193,N_656);
and U1453 (N_1453,N_774,N_314);
and U1454 (N_1454,N_617,N_305);
nand U1455 (N_1455,N_636,N_354);
and U1456 (N_1456,N_835,N_783);
and U1457 (N_1457,N_156,N_28);
xor U1458 (N_1458,N_886,N_377);
nor U1459 (N_1459,N_737,N_277);
nand U1460 (N_1460,N_138,N_971);
nand U1461 (N_1461,N_170,N_444);
nand U1462 (N_1462,N_66,N_825);
or U1463 (N_1463,N_972,N_519);
nor U1464 (N_1464,N_721,N_271);
nand U1465 (N_1465,N_172,N_125);
or U1466 (N_1466,N_916,N_558);
nand U1467 (N_1467,N_716,N_56);
and U1468 (N_1468,N_975,N_40);
xor U1469 (N_1469,N_720,N_749);
and U1470 (N_1470,N_175,N_139);
and U1471 (N_1471,N_556,N_943);
or U1472 (N_1472,N_298,N_187);
and U1473 (N_1473,N_107,N_927);
or U1474 (N_1474,N_933,N_47);
nor U1475 (N_1475,N_620,N_407);
nand U1476 (N_1476,N_622,N_562);
nand U1477 (N_1477,N_384,N_609);
xor U1478 (N_1478,N_418,N_69);
and U1479 (N_1479,N_803,N_512);
nand U1480 (N_1480,N_946,N_420);
and U1481 (N_1481,N_221,N_759);
nand U1482 (N_1482,N_232,N_513);
nand U1483 (N_1483,N_870,N_883);
nand U1484 (N_1484,N_544,N_247);
and U1485 (N_1485,N_765,N_462);
nand U1486 (N_1486,N_666,N_486);
nor U1487 (N_1487,N_70,N_919);
nand U1488 (N_1488,N_76,N_497);
and U1489 (N_1489,N_256,N_748);
and U1490 (N_1490,N_231,N_313);
nand U1491 (N_1491,N_357,N_732);
or U1492 (N_1492,N_677,N_735);
nand U1493 (N_1493,N_980,N_821);
xnor U1494 (N_1494,N_176,N_534);
xnor U1495 (N_1495,N_528,N_703);
nand U1496 (N_1496,N_658,N_98);
or U1497 (N_1497,N_106,N_372);
and U1498 (N_1498,N_599,N_985);
or U1499 (N_1499,N_942,N_347);
or U1500 (N_1500,N_446,N_598);
nand U1501 (N_1501,N_640,N_662);
nor U1502 (N_1502,N_743,N_546);
and U1503 (N_1503,N_618,N_941);
and U1504 (N_1504,N_234,N_221);
and U1505 (N_1505,N_535,N_411);
or U1506 (N_1506,N_230,N_93);
or U1507 (N_1507,N_545,N_882);
or U1508 (N_1508,N_576,N_222);
nand U1509 (N_1509,N_19,N_289);
nor U1510 (N_1510,N_429,N_643);
nand U1511 (N_1511,N_89,N_658);
nand U1512 (N_1512,N_21,N_771);
and U1513 (N_1513,N_430,N_464);
and U1514 (N_1514,N_795,N_426);
nand U1515 (N_1515,N_803,N_386);
xnor U1516 (N_1516,N_581,N_328);
or U1517 (N_1517,N_955,N_674);
and U1518 (N_1518,N_813,N_171);
and U1519 (N_1519,N_602,N_222);
or U1520 (N_1520,N_459,N_113);
or U1521 (N_1521,N_59,N_126);
or U1522 (N_1522,N_969,N_913);
xnor U1523 (N_1523,N_750,N_255);
and U1524 (N_1524,N_322,N_161);
or U1525 (N_1525,N_699,N_350);
nand U1526 (N_1526,N_91,N_938);
and U1527 (N_1527,N_528,N_639);
or U1528 (N_1528,N_717,N_387);
or U1529 (N_1529,N_615,N_661);
nand U1530 (N_1530,N_401,N_799);
and U1531 (N_1531,N_119,N_343);
and U1532 (N_1532,N_522,N_128);
and U1533 (N_1533,N_260,N_329);
xor U1534 (N_1534,N_687,N_539);
xor U1535 (N_1535,N_542,N_31);
or U1536 (N_1536,N_415,N_115);
nor U1537 (N_1537,N_991,N_375);
and U1538 (N_1538,N_161,N_325);
and U1539 (N_1539,N_735,N_65);
or U1540 (N_1540,N_380,N_243);
nand U1541 (N_1541,N_451,N_974);
nor U1542 (N_1542,N_519,N_455);
nor U1543 (N_1543,N_470,N_293);
and U1544 (N_1544,N_339,N_870);
nand U1545 (N_1545,N_352,N_785);
and U1546 (N_1546,N_778,N_473);
nor U1547 (N_1547,N_295,N_443);
or U1548 (N_1548,N_368,N_569);
and U1549 (N_1549,N_370,N_135);
nor U1550 (N_1550,N_990,N_955);
nor U1551 (N_1551,N_66,N_135);
or U1552 (N_1552,N_249,N_993);
nand U1553 (N_1553,N_19,N_589);
and U1554 (N_1554,N_752,N_396);
nand U1555 (N_1555,N_204,N_343);
or U1556 (N_1556,N_434,N_526);
nand U1557 (N_1557,N_539,N_268);
and U1558 (N_1558,N_298,N_511);
or U1559 (N_1559,N_689,N_855);
and U1560 (N_1560,N_295,N_868);
nor U1561 (N_1561,N_44,N_24);
or U1562 (N_1562,N_740,N_113);
nor U1563 (N_1563,N_225,N_3);
and U1564 (N_1564,N_194,N_118);
nor U1565 (N_1565,N_248,N_597);
nor U1566 (N_1566,N_995,N_710);
or U1567 (N_1567,N_870,N_614);
and U1568 (N_1568,N_48,N_345);
xor U1569 (N_1569,N_52,N_466);
and U1570 (N_1570,N_722,N_434);
or U1571 (N_1571,N_358,N_66);
nor U1572 (N_1572,N_966,N_707);
nand U1573 (N_1573,N_859,N_892);
nor U1574 (N_1574,N_137,N_22);
and U1575 (N_1575,N_89,N_738);
and U1576 (N_1576,N_437,N_556);
nand U1577 (N_1577,N_904,N_296);
nand U1578 (N_1578,N_790,N_935);
nand U1579 (N_1579,N_232,N_727);
xnor U1580 (N_1580,N_495,N_831);
nor U1581 (N_1581,N_960,N_902);
and U1582 (N_1582,N_480,N_30);
nand U1583 (N_1583,N_697,N_963);
nand U1584 (N_1584,N_852,N_645);
or U1585 (N_1585,N_102,N_403);
nor U1586 (N_1586,N_524,N_768);
nand U1587 (N_1587,N_124,N_320);
or U1588 (N_1588,N_453,N_205);
xor U1589 (N_1589,N_346,N_143);
or U1590 (N_1590,N_555,N_767);
or U1591 (N_1591,N_289,N_624);
nand U1592 (N_1592,N_471,N_722);
and U1593 (N_1593,N_869,N_562);
nand U1594 (N_1594,N_190,N_623);
nand U1595 (N_1595,N_926,N_427);
nor U1596 (N_1596,N_198,N_910);
and U1597 (N_1597,N_662,N_465);
nand U1598 (N_1598,N_722,N_705);
xnor U1599 (N_1599,N_300,N_736);
nor U1600 (N_1600,N_496,N_62);
and U1601 (N_1601,N_233,N_458);
nor U1602 (N_1602,N_472,N_259);
nand U1603 (N_1603,N_267,N_444);
or U1604 (N_1604,N_475,N_431);
and U1605 (N_1605,N_915,N_252);
or U1606 (N_1606,N_246,N_242);
nand U1607 (N_1607,N_905,N_533);
nor U1608 (N_1608,N_252,N_487);
and U1609 (N_1609,N_665,N_504);
nand U1610 (N_1610,N_764,N_332);
nand U1611 (N_1611,N_418,N_284);
and U1612 (N_1612,N_215,N_522);
and U1613 (N_1613,N_174,N_693);
and U1614 (N_1614,N_939,N_139);
and U1615 (N_1615,N_255,N_983);
and U1616 (N_1616,N_11,N_976);
and U1617 (N_1617,N_266,N_415);
or U1618 (N_1618,N_30,N_625);
or U1619 (N_1619,N_384,N_478);
nor U1620 (N_1620,N_765,N_692);
xnor U1621 (N_1621,N_255,N_154);
nand U1622 (N_1622,N_281,N_570);
or U1623 (N_1623,N_852,N_818);
and U1624 (N_1624,N_618,N_175);
and U1625 (N_1625,N_151,N_795);
nor U1626 (N_1626,N_149,N_150);
nor U1627 (N_1627,N_667,N_208);
nor U1628 (N_1628,N_692,N_486);
nand U1629 (N_1629,N_958,N_747);
nand U1630 (N_1630,N_660,N_0);
nand U1631 (N_1631,N_760,N_192);
nor U1632 (N_1632,N_57,N_513);
or U1633 (N_1633,N_963,N_943);
nand U1634 (N_1634,N_442,N_197);
nor U1635 (N_1635,N_622,N_80);
nand U1636 (N_1636,N_477,N_561);
and U1637 (N_1637,N_680,N_485);
and U1638 (N_1638,N_321,N_544);
nand U1639 (N_1639,N_173,N_833);
nor U1640 (N_1640,N_413,N_715);
nor U1641 (N_1641,N_563,N_19);
and U1642 (N_1642,N_819,N_42);
or U1643 (N_1643,N_330,N_515);
nand U1644 (N_1644,N_161,N_645);
or U1645 (N_1645,N_644,N_166);
or U1646 (N_1646,N_274,N_701);
nor U1647 (N_1647,N_261,N_932);
nand U1648 (N_1648,N_859,N_315);
and U1649 (N_1649,N_157,N_833);
nand U1650 (N_1650,N_559,N_287);
nor U1651 (N_1651,N_501,N_949);
nand U1652 (N_1652,N_491,N_34);
or U1653 (N_1653,N_594,N_547);
xor U1654 (N_1654,N_163,N_601);
nor U1655 (N_1655,N_524,N_838);
and U1656 (N_1656,N_524,N_256);
nand U1657 (N_1657,N_773,N_397);
or U1658 (N_1658,N_424,N_332);
or U1659 (N_1659,N_515,N_614);
and U1660 (N_1660,N_373,N_138);
nand U1661 (N_1661,N_440,N_187);
nor U1662 (N_1662,N_785,N_271);
nor U1663 (N_1663,N_290,N_459);
nand U1664 (N_1664,N_429,N_135);
nor U1665 (N_1665,N_328,N_576);
nand U1666 (N_1666,N_908,N_416);
and U1667 (N_1667,N_316,N_88);
or U1668 (N_1668,N_706,N_993);
or U1669 (N_1669,N_872,N_926);
nand U1670 (N_1670,N_543,N_205);
xor U1671 (N_1671,N_662,N_186);
nor U1672 (N_1672,N_384,N_28);
or U1673 (N_1673,N_615,N_648);
and U1674 (N_1674,N_841,N_323);
or U1675 (N_1675,N_989,N_142);
or U1676 (N_1676,N_774,N_329);
and U1677 (N_1677,N_511,N_54);
nor U1678 (N_1678,N_579,N_967);
or U1679 (N_1679,N_917,N_521);
and U1680 (N_1680,N_857,N_207);
and U1681 (N_1681,N_820,N_71);
or U1682 (N_1682,N_360,N_820);
or U1683 (N_1683,N_352,N_347);
nor U1684 (N_1684,N_890,N_571);
and U1685 (N_1685,N_405,N_875);
and U1686 (N_1686,N_756,N_511);
nor U1687 (N_1687,N_520,N_453);
nor U1688 (N_1688,N_676,N_442);
xnor U1689 (N_1689,N_234,N_458);
xor U1690 (N_1690,N_305,N_83);
nor U1691 (N_1691,N_809,N_379);
nand U1692 (N_1692,N_635,N_836);
xnor U1693 (N_1693,N_6,N_264);
nand U1694 (N_1694,N_737,N_356);
or U1695 (N_1695,N_310,N_385);
or U1696 (N_1696,N_456,N_123);
nor U1697 (N_1697,N_829,N_392);
xnor U1698 (N_1698,N_214,N_148);
or U1699 (N_1699,N_405,N_130);
nand U1700 (N_1700,N_948,N_124);
or U1701 (N_1701,N_855,N_3);
xor U1702 (N_1702,N_233,N_681);
nor U1703 (N_1703,N_481,N_611);
and U1704 (N_1704,N_503,N_437);
or U1705 (N_1705,N_495,N_645);
and U1706 (N_1706,N_218,N_246);
nor U1707 (N_1707,N_17,N_652);
or U1708 (N_1708,N_436,N_887);
nor U1709 (N_1709,N_705,N_895);
and U1710 (N_1710,N_731,N_658);
xnor U1711 (N_1711,N_60,N_685);
xor U1712 (N_1712,N_415,N_369);
and U1713 (N_1713,N_244,N_379);
nand U1714 (N_1714,N_490,N_793);
nor U1715 (N_1715,N_310,N_806);
and U1716 (N_1716,N_866,N_915);
nand U1717 (N_1717,N_620,N_315);
nand U1718 (N_1718,N_782,N_260);
or U1719 (N_1719,N_921,N_224);
and U1720 (N_1720,N_568,N_246);
or U1721 (N_1721,N_737,N_10);
or U1722 (N_1722,N_226,N_215);
nor U1723 (N_1723,N_940,N_917);
or U1724 (N_1724,N_504,N_694);
and U1725 (N_1725,N_289,N_489);
nand U1726 (N_1726,N_294,N_629);
and U1727 (N_1727,N_133,N_558);
nand U1728 (N_1728,N_654,N_960);
nand U1729 (N_1729,N_439,N_887);
and U1730 (N_1730,N_79,N_465);
and U1731 (N_1731,N_673,N_723);
nor U1732 (N_1732,N_832,N_204);
nand U1733 (N_1733,N_46,N_400);
or U1734 (N_1734,N_972,N_89);
and U1735 (N_1735,N_295,N_871);
nor U1736 (N_1736,N_901,N_178);
xnor U1737 (N_1737,N_131,N_723);
nor U1738 (N_1738,N_899,N_797);
nor U1739 (N_1739,N_406,N_39);
nor U1740 (N_1740,N_607,N_47);
and U1741 (N_1741,N_307,N_333);
and U1742 (N_1742,N_958,N_276);
and U1743 (N_1743,N_422,N_959);
or U1744 (N_1744,N_524,N_771);
and U1745 (N_1745,N_414,N_952);
nand U1746 (N_1746,N_415,N_168);
nor U1747 (N_1747,N_678,N_803);
nand U1748 (N_1748,N_869,N_437);
and U1749 (N_1749,N_597,N_878);
and U1750 (N_1750,N_958,N_652);
and U1751 (N_1751,N_823,N_55);
and U1752 (N_1752,N_873,N_607);
and U1753 (N_1753,N_44,N_517);
and U1754 (N_1754,N_520,N_902);
and U1755 (N_1755,N_791,N_570);
and U1756 (N_1756,N_994,N_872);
nand U1757 (N_1757,N_211,N_2);
xnor U1758 (N_1758,N_120,N_454);
and U1759 (N_1759,N_598,N_767);
or U1760 (N_1760,N_965,N_479);
nor U1761 (N_1761,N_633,N_133);
and U1762 (N_1762,N_1,N_839);
and U1763 (N_1763,N_454,N_694);
or U1764 (N_1764,N_600,N_712);
nand U1765 (N_1765,N_587,N_750);
or U1766 (N_1766,N_421,N_263);
nand U1767 (N_1767,N_695,N_876);
nor U1768 (N_1768,N_790,N_60);
nor U1769 (N_1769,N_546,N_167);
nand U1770 (N_1770,N_802,N_25);
or U1771 (N_1771,N_469,N_119);
or U1772 (N_1772,N_629,N_837);
or U1773 (N_1773,N_790,N_70);
nor U1774 (N_1774,N_313,N_688);
nor U1775 (N_1775,N_592,N_365);
nand U1776 (N_1776,N_587,N_177);
and U1777 (N_1777,N_751,N_885);
or U1778 (N_1778,N_907,N_492);
nor U1779 (N_1779,N_66,N_946);
or U1780 (N_1780,N_324,N_127);
nand U1781 (N_1781,N_627,N_631);
nor U1782 (N_1782,N_848,N_742);
or U1783 (N_1783,N_659,N_392);
or U1784 (N_1784,N_844,N_762);
nand U1785 (N_1785,N_183,N_524);
and U1786 (N_1786,N_193,N_578);
and U1787 (N_1787,N_204,N_425);
or U1788 (N_1788,N_151,N_17);
and U1789 (N_1789,N_73,N_464);
and U1790 (N_1790,N_571,N_906);
and U1791 (N_1791,N_538,N_281);
or U1792 (N_1792,N_578,N_480);
nor U1793 (N_1793,N_720,N_515);
and U1794 (N_1794,N_969,N_812);
and U1795 (N_1795,N_740,N_900);
nor U1796 (N_1796,N_890,N_955);
nor U1797 (N_1797,N_78,N_494);
nor U1798 (N_1798,N_850,N_314);
and U1799 (N_1799,N_837,N_218);
nand U1800 (N_1800,N_373,N_811);
and U1801 (N_1801,N_754,N_818);
nor U1802 (N_1802,N_269,N_785);
xnor U1803 (N_1803,N_177,N_594);
and U1804 (N_1804,N_668,N_209);
nand U1805 (N_1805,N_589,N_313);
nand U1806 (N_1806,N_478,N_332);
xnor U1807 (N_1807,N_582,N_443);
nor U1808 (N_1808,N_448,N_171);
xnor U1809 (N_1809,N_130,N_63);
and U1810 (N_1810,N_542,N_676);
or U1811 (N_1811,N_127,N_782);
or U1812 (N_1812,N_417,N_112);
or U1813 (N_1813,N_356,N_636);
xnor U1814 (N_1814,N_729,N_264);
nor U1815 (N_1815,N_322,N_883);
nand U1816 (N_1816,N_144,N_15);
xnor U1817 (N_1817,N_649,N_539);
or U1818 (N_1818,N_312,N_623);
nand U1819 (N_1819,N_3,N_64);
or U1820 (N_1820,N_681,N_222);
or U1821 (N_1821,N_344,N_500);
or U1822 (N_1822,N_377,N_35);
nor U1823 (N_1823,N_179,N_221);
or U1824 (N_1824,N_458,N_427);
nand U1825 (N_1825,N_932,N_573);
nand U1826 (N_1826,N_613,N_372);
xnor U1827 (N_1827,N_662,N_62);
or U1828 (N_1828,N_988,N_852);
nand U1829 (N_1829,N_282,N_760);
nor U1830 (N_1830,N_469,N_940);
nand U1831 (N_1831,N_400,N_567);
nor U1832 (N_1832,N_852,N_618);
nor U1833 (N_1833,N_13,N_206);
or U1834 (N_1834,N_428,N_669);
and U1835 (N_1835,N_221,N_706);
nor U1836 (N_1836,N_358,N_793);
nor U1837 (N_1837,N_169,N_72);
nand U1838 (N_1838,N_824,N_768);
nor U1839 (N_1839,N_305,N_572);
nand U1840 (N_1840,N_84,N_569);
xnor U1841 (N_1841,N_516,N_645);
nor U1842 (N_1842,N_584,N_249);
or U1843 (N_1843,N_425,N_912);
or U1844 (N_1844,N_595,N_412);
nor U1845 (N_1845,N_21,N_311);
nor U1846 (N_1846,N_345,N_453);
or U1847 (N_1847,N_218,N_556);
nand U1848 (N_1848,N_926,N_589);
or U1849 (N_1849,N_825,N_313);
nor U1850 (N_1850,N_279,N_313);
and U1851 (N_1851,N_3,N_359);
nand U1852 (N_1852,N_817,N_992);
and U1853 (N_1853,N_25,N_715);
nor U1854 (N_1854,N_586,N_342);
and U1855 (N_1855,N_628,N_28);
nand U1856 (N_1856,N_752,N_876);
nand U1857 (N_1857,N_596,N_136);
nor U1858 (N_1858,N_489,N_77);
and U1859 (N_1859,N_415,N_407);
or U1860 (N_1860,N_707,N_60);
xnor U1861 (N_1861,N_238,N_507);
or U1862 (N_1862,N_58,N_73);
nor U1863 (N_1863,N_9,N_723);
nor U1864 (N_1864,N_654,N_862);
or U1865 (N_1865,N_827,N_290);
nor U1866 (N_1866,N_196,N_280);
and U1867 (N_1867,N_317,N_62);
or U1868 (N_1868,N_624,N_637);
or U1869 (N_1869,N_383,N_78);
and U1870 (N_1870,N_279,N_207);
nor U1871 (N_1871,N_105,N_935);
or U1872 (N_1872,N_71,N_99);
nor U1873 (N_1873,N_151,N_319);
and U1874 (N_1874,N_430,N_711);
nor U1875 (N_1875,N_194,N_518);
or U1876 (N_1876,N_543,N_93);
nand U1877 (N_1877,N_754,N_183);
nand U1878 (N_1878,N_916,N_508);
and U1879 (N_1879,N_31,N_937);
nor U1880 (N_1880,N_244,N_387);
and U1881 (N_1881,N_377,N_470);
and U1882 (N_1882,N_971,N_109);
nor U1883 (N_1883,N_551,N_350);
or U1884 (N_1884,N_769,N_15);
nand U1885 (N_1885,N_765,N_205);
nor U1886 (N_1886,N_334,N_102);
and U1887 (N_1887,N_145,N_905);
or U1888 (N_1888,N_886,N_957);
nand U1889 (N_1889,N_787,N_472);
or U1890 (N_1890,N_8,N_397);
nand U1891 (N_1891,N_443,N_146);
nand U1892 (N_1892,N_988,N_939);
and U1893 (N_1893,N_581,N_295);
or U1894 (N_1894,N_516,N_931);
or U1895 (N_1895,N_269,N_419);
or U1896 (N_1896,N_81,N_377);
or U1897 (N_1897,N_628,N_828);
and U1898 (N_1898,N_986,N_1);
xor U1899 (N_1899,N_163,N_90);
xor U1900 (N_1900,N_151,N_446);
and U1901 (N_1901,N_23,N_614);
or U1902 (N_1902,N_858,N_218);
or U1903 (N_1903,N_537,N_78);
nand U1904 (N_1904,N_178,N_357);
nand U1905 (N_1905,N_729,N_858);
nor U1906 (N_1906,N_13,N_27);
and U1907 (N_1907,N_241,N_295);
or U1908 (N_1908,N_596,N_872);
and U1909 (N_1909,N_409,N_459);
and U1910 (N_1910,N_683,N_235);
and U1911 (N_1911,N_332,N_487);
nor U1912 (N_1912,N_964,N_965);
and U1913 (N_1913,N_815,N_297);
and U1914 (N_1914,N_723,N_808);
and U1915 (N_1915,N_371,N_403);
nand U1916 (N_1916,N_801,N_591);
nand U1917 (N_1917,N_529,N_776);
nand U1918 (N_1918,N_403,N_988);
and U1919 (N_1919,N_130,N_535);
and U1920 (N_1920,N_667,N_502);
nor U1921 (N_1921,N_560,N_183);
nor U1922 (N_1922,N_129,N_398);
nor U1923 (N_1923,N_700,N_402);
xnor U1924 (N_1924,N_65,N_292);
or U1925 (N_1925,N_859,N_553);
nand U1926 (N_1926,N_348,N_952);
xnor U1927 (N_1927,N_922,N_505);
nor U1928 (N_1928,N_759,N_132);
nand U1929 (N_1929,N_666,N_444);
xnor U1930 (N_1930,N_468,N_143);
nand U1931 (N_1931,N_783,N_226);
and U1932 (N_1932,N_634,N_949);
nand U1933 (N_1933,N_397,N_335);
nor U1934 (N_1934,N_583,N_3);
and U1935 (N_1935,N_783,N_882);
nor U1936 (N_1936,N_470,N_628);
and U1937 (N_1937,N_212,N_33);
nand U1938 (N_1938,N_42,N_600);
nand U1939 (N_1939,N_299,N_827);
nor U1940 (N_1940,N_319,N_510);
nand U1941 (N_1941,N_694,N_839);
nor U1942 (N_1942,N_769,N_456);
and U1943 (N_1943,N_820,N_400);
and U1944 (N_1944,N_715,N_86);
and U1945 (N_1945,N_318,N_6);
nor U1946 (N_1946,N_307,N_784);
nand U1947 (N_1947,N_457,N_879);
or U1948 (N_1948,N_42,N_132);
or U1949 (N_1949,N_515,N_486);
or U1950 (N_1950,N_669,N_125);
and U1951 (N_1951,N_56,N_368);
or U1952 (N_1952,N_600,N_332);
and U1953 (N_1953,N_600,N_917);
or U1954 (N_1954,N_98,N_140);
or U1955 (N_1955,N_727,N_717);
nor U1956 (N_1956,N_43,N_108);
nand U1957 (N_1957,N_657,N_812);
xor U1958 (N_1958,N_266,N_291);
or U1959 (N_1959,N_94,N_179);
nor U1960 (N_1960,N_43,N_811);
or U1961 (N_1961,N_191,N_243);
and U1962 (N_1962,N_243,N_200);
nand U1963 (N_1963,N_942,N_382);
nand U1964 (N_1964,N_679,N_617);
nor U1965 (N_1965,N_544,N_599);
nor U1966 (N_1966,N_380,N_80);
or U1967 (N_1967,N_629,N_377);
nand U1968 (N_1968,N_427,N_666);
nor U1969 (N_1969,N_532,N_188);
nand U1970 (N_1970,N_938,N_200);
and U1971 (N_1971,N_52,N_405);
nor U1972 (N_1972,N_883,N_877);
nor U1973 (N_1973,N_964,N_482);
or U1974 (N_1974,N_434,N_282);
xor U1975 (N_1975,N_754,N_225);
xnor U1976 (N_1976,N_890,N_215);
nor U1977 (N_1977,N_703,N_472);
nand U1978 (N_1978,N_745,N_255);
xor U1979 (N_1979,N_612,N_847);
nand U1980 (N_1980,N_414,N_767);
xor U1981 (N_1981,N_793,N_292);
xor U1982 (N_1982,N_550,N_730);
or U1983 (N_1983,N_952,N_748);
nor U1984 (N_1984,N_826,N_93);
nand U1985 (N_1985,N_661,N_852);
or U1986 (N_1986,N_248,N_816);
nand U1987 (N_1987,N_189,N_367);
or U1988 (N_1988,N_580,N_396);
and U1989 (N_1989,N_11,N_372);
nor U1990 (N_1990,N_948,N_139);
nand U1991 (N_1991,N_308,N_408);
and U1992 (N_1992,N_234,N_842);
nand U1993 (N_1993,N_664,N_313);
nor U1994 (N_1994,N_292,N_163);
nand U1995 (N_1995,N_503,N_254);
nor U1996 (N_1996,N_427,N_624);
nor U1997 (N_1997,N_659,N_664);
xor U1998 (N_1998,N_536,N_789);
or U1999 (N_1999,N_922,N_23);
nor U2000 (N_2000,N_1502,N_1879);
nor U2001 (N_2001,N_1573,N_1032);
nor U2002 (N_2002,N_1805,N_1344);
or U2003 (N_2003,N_1629,N_1345);
nand U2004 (N_2004,N_1818,N_1135);
xor U2005 (N_2005,N_1668,N_1029);
or U2006 (N_2006,N_1289,N_1428);
nand U2007 (N_2007,N_1496,N_1855);
or U2008 (N_2008,N_1710,N_1619);
nand U2009 (N_2009,N_1579,N_1305);
nand U2010 (N_2010,N_1337,N_1241);
and U2011 (N_2011,N_1012,N_1625);
and U2012 (N_2012,N_1764,N_1633);
and U2013 (N_2013,N_1970,N_1533);
and U2014 (N_2014,N_1176,N_1596);
and U2015 (N_2015,N_1813,N_1831);
or U2016 (N_2016,N_1525,N_1228);
nor U2017 (N_2017,N_1508,N_1900);
nand U2018 (N_2018,N_1954,N_1922);
nor U2019 (N_2019,N_1258,N_1053);
and U2020 (N_2020,N_1595,N_1203);
and U2021 (N_2021,N_1683,N_1482);
nand U2022 (N_2022,N_1811,N_1038);
or U2023 (N_2023,N_1156,N_1812);
nand U2024 (N_2024,N_1751,N_1070);
or U2025 (N_2025,N_1055,N_1988);
nand U2026 (N_2026,N_1732,N_1825);
and U2027 (N_2027,N_1715,N_1202);
nand U2028 (N_2028,N_1528,N_1438);
and U2029 (N_2029,N_1653,N_1192);
nand U2030 (N_2030,N_1948,N_1404);
or U2031 (N_2031,N_1475,N_1309);
and U2032 (N_2032,N_1935,N_1356);
or U2033 (N_2033,N_1762,N_1031);
xor U2034 (N_2034,N_1924,N_1105);
nor U2035 (N_2035,N_1355,N_1590);
xor U2036 (N_2036,N_1999,N_1223);
nand U2037 (N_2037,N_1981,N_1326);
nand U2038 (N_2038,N_1374,N_1684);
nor U2039 (N_2039,N_1681,N_1616);
or U2040 (N_2040,N_1214,N_1276);
xor U2041 (N_2041,N_1285,N_1361);
or U2042 (N_2042,N_1154,N_1264);
nor U2043 (N_2043,N_1772,N_1101);
nand U2044 (N_2044,N_1499,N_1645);
nor U2045 (N_2045,N_1942,N_1898);
and U2046 (N_2046,N_1737,N_1410);
nor U2047 (N_2047,N_1092,N_1717);
and U2048 (N_2048,N_1474,N_1709);
or U2049 (N_2049,N_1048,N_1399);
and U2050 (N_2050,N_1876,N_1023);
or U2051 (N_2051,N_1511,N_1131);
nor U2052 (N_2052,N_1330,N_1087);
and U2053 (N_2053,N_1507,N_1538);
nor U2054 (N_2054,N_1464,N_1632);
or U2055 (N_2055,N_1465,N_1166);
xor U2056 (N_2056,N_1054,N_1072);
nor U2057 (N_2057,N_1789,N_1130);
or U2058 (N_2058,N_1125,N_1868);
xnor U2059 (N_2059,N_1771,N_1980);
nand U2060 (N_2060,N_1147,N_1841);
and U2061 (N_2061,N_1586,N_1901);
nor U2062 (N_2062,N_1765,N_1743);
and U2063 (N_2063,N_1052,N_1910);
or U2064 (N_2064,N_1444,N_1251);
nor U2065 (N_2065,N_1049,N_1421);
nor U2066 (N_2066,N_1115,N_1484);
or U2067 (N_2067,N_1576,N_1673);
and U2068 (N_2068,N_1918,N_1102);
nor U2069 (N_2069,N_1895,N_1057);
nor U2070 (N_2070,N_1697,N_1015);
nor U2071 (N_2071,N_1550,N_1318);
and U2072 (N_2072,N_1729,N_1845);
xor U2073 (N_2073,N_1553,N_1187);
or U2074 (N_2074,N_1298,N_1140);
nand U2075 (N_2075,N_1617,N_1614);
nand U2076 (N_2076,N_1201,N_1299);
and U2077 (N_2077,N_1725,N_1064);
nor U2078 (N_2078,N_1395,N_1069);
nand U2079 (N_2079,N_1852,N_1363);
nor U2080 (N_2080,N_1408,N_1396);
and U2081 (N_2081,N_1104,N_1992);
and U2082 (N_2082,N_1001,N_1951);
and U2083 (N_2083,N_1445,N_1664);
and U2084 (N_2084,N_1008,N_1422);
and U2085 (N_2085,N_1768,N_1557);
and U2086 (N_2086,N_1136,N_1711);
nor U2087 (N_2087,N_1184,N_1262);
and U2088 (N_2088,N_1928,N_1229);
nor U2089 (N_2089,N_1007,N_1562);
or U2090 (N_2090,N_1675,N_1490);
nor U2091 (N_2091,N_1952,N_1893);
nand U2092 (N_2092,N_1979,N_1220);
nor U2093 (N_2093,N_1856,N_1416);
nand U2094 (N_2094,N_1036,N_1721);
or U2095 (N_2095,N_1787,N_1760);
xnor U2096 (N_2096,N_1584,N_1969);
or U2097 (N_2097,N_1107,N_1839);
nand U2098 (N_2098,N_1338,N_1836);
or U2099 (N_2099,N_1034,N_1545);
or U2100 (N_2100,N_1110,N_1466);
nand U2101 (N_2101,N_1854,N_1727);
nand U2102 (N_2102,N_1733,N_1714);
and U2103 (N_2103,N_1062,N_1837);
nor U2104 (N_2104,N_1148,N_1091);
xor U2105 (N_2105,N_1934,N_1244);
nand U2106 (N_2106,N_1660,N_1539);
nand U2107 (N_2107,N_1128,N_1249);
nand U2108 (N_2108,N_1866,N_1367);
nand U2109 (N_2109,N_1358,N_1761);
nor U2110 (N_2110,N_1132,N_1405);
or U2111 (N_2111,N_1861,N_1937);
nand U2112 (N_2112,N_1044,N_1779);
nand U2113 (N_2113,N_1067,N_1529);
nand U2114 (N_2114,N_1526,N_1234);
and U2115 (N_2115,N_1256,N_1118);
or U2116 (N_2116,N_1548,N_1078);
nor U2117 (N_2117,N_1293,N_1639);
or U2118 (N_2118,N_1902,N_1303);
xor U2119 (N_2119,N_1409,N_1597);
nor U2120 (N_2120,N_1261,N_1674);
nor U2121 (N_2121,N_1860,N_1844);
nor U2122 (N_2122,N_1068,N_1752);
nor U2123 (N_2123,N_1749,N_1437);
nor U2124 (N_2124,N_1495,N_1759);
and U2125 (N_2125,N_1349,N_1451);
and U2126 (N_2126,N_1987,N_1050);
nor U2127 (N_2127,N_1966,N_1609);
nor U2128 (N_2128,N_1277,N_1603);
nor U2129 (N_2129,N_1065,N_1534);
or U2130 (N_2130,N_1366,N_1955);
nor U2131 (N_2131,N_1699,N_1317);
nor U2132 (N_2132,N_1212,N_1731);
and U2133 (N_2133,N_1155,N_1327);
and U2134 (N_2134,N_1191,N_1167);
nand U2135 (N_2135,N_1378,N_1630);
or U2136 (N_2136,N_1141,N_1708);
nand U2137 (N_2137,N_1635,N_1060);
or U2138 (N_2138,N_1306,N_1843);
nor U2139 (N_2139,N_1835,N_1041);
and U2140 (N_2140,N_1111,N_1369);
nand U2141 (N_2141,N_1613,N_1758);
and U2142 (N_2142,N_1195,N_1800);
xor U2143 (N_2143,N_1546,N_1564);
nor U2144 (N_2144,N_1292,N_1974);
nand U2145 (N_2145,N_1583,N_1996);
or U2146 (N_2146,N_1077,N_1314);
nor U2147 (N_2147,N_1447,N_1903);
nand U2148 (N_2148,N_1936,N_1393);
nand U2149 (N_2149,N_1139,N_1657);
and U2150 (N_2150,N_1436,N_1585);
nor U2151 (N_2151,N_1061,N_1706);
nand U2152 (N_2152,N_1501,N_1198);
nand U2153 (N_2153,N_1472,N_1875);
nand U2154 (N_2154,N_1341,N_1990);
and U2155 (N_2155,N_1331,N_1536);
nand U2156 (N_2156,N_1100,N_1368);
nor U2157 (N_2157,N_1527,N_1089);
or U2158 (N_2158,N_1186,N_1209);
xor U2159 (N_2159,N_1857,N_1371);
or U2160 (N_2160,N_1450,N_1888);
nand U2161 (N_2161,N_1975,N_1178);
or U2162 (N_2162,N_1941,N_1607);
nand U2163 (N_2163,N_1667,N_1082);
or U2164 (N_2164,N_1566,N_1881);
nor U2165 (N_2165,N_1321,N_1809);
nand U2166 (N_2166,N_1871,N_1016);
nand U2167 (N_2167,N_1917,N_1252);
and U2168 (N_2168,N_1134,N_1976);
or U2169 (N_2169,N_1763,N_1340);
or U2170 (N_2170,N_1865,N_1365);
or U2171 (N_2171,N_1608,N_1520);
or U2172 (N_2172,N_1690,N_1773);
or U2173 (N_2173,N_1913,N_1040);
xor U2174 (N_2174,N_1420,N_1322);
nand U2175 (N_2175,N_1046,N_1686);
or U2176 (N_2176,N_1215,N_1523);
nand U2177 (N_2177,N_1803,N_1886);
and U2178 (N_2178,N_1470,N_1418);
xnor U2179 (N_2179,N_1682,N_1424);
or U2180 (N_2180,N_1850,N_1204);
xor U2181 (N_2181,N_1869,N_1076);
or U2182 (N_2182,N_1827,N_1138);
nand U2183 (N_2183,N_1612,N_1571);
xor U2184 (N_2184,N_1964,N_1766);
nor U2185 (N_2185,N_1904,N_1381);
or U2186 (N_2186,N_1647,N_1672);
or U2187 (N_2187,N_1940,N_1830);
nor U2188 (N_2188,N_1042,N_1119);
and U2189 (N_2189,N_1792,N_1093);
nand U2190 (N_2190,N_1582,N_1026);
and U2191 (N_2191,N_1781,N_1921);
and U2192 (N_2192,N_1847,N_1696);
nand U2193 (N_2193,N_1649,N_1103);
nand U2194 (N_2194,N_1384,N_1601);
and U2195 (N_2195,N_1808,N_1221);
nor U2196 (N_2196,N_1775,N_1943);
nand U2197 (N_2197,N_1059,N_1972);
and U2198 (N_2198,N_1926,N_1636);
or U2199 (N_2199,N_1821,N_1098);
nand U2200 (N_2200,N_1577,N_1503);
nor U2201 (N_2201,N_1905,N_1513);
nor U2202 (N_2202,N_1694,N_1494);
nand U2203 (N_2203,N_1920,N_1021);
nor U2204 (N_2204,N_1419,N_1750);
xnor U2205 (N_2205,N_1112,N_1791);
and U2206 (N_2206,N_1572,N_1307);
and U2207 (N_2207,N_1480,N_1829);
nand U2208 (N_2208,N_1310,N_1073);
or U2209 (N_2209,N_1174,N_1376);
nand U2210 (N_2210,N_1932,N_1730);
or U2211 (N_2211,N_1887,N_1810);
or U2212 (N_2212,N_1379,N_1250);
nor U2213 (N_2213,N_1628,N_1896);
nand U2214 (N_2214,N_1488,N_1144);
and U2215 (N_2215,N_1084,N_1991);
xnor U2216 (N_2216,N_1334,N_1149);
nor U2217 (N_2217,N_1017,N_1978);
nor U2218 (N_2218,N_1965,N_1207);
and U2219 (N_2219,N_1531,N_1815);
nand U2220 (N_2220,N_1517,N_1554);
nand U2221 (N_2221,N_1137,N_1197);
nor U2222 (N_2222,N_1817,N_1161);
and U2223 (N_2223,N_1985,N_1315);
xnor U2224 (N_2224,N_1169,N_1086);
and U2225 (N_2225,N_1736,N_1183);
and U2226 (N_2226,N_1287,N_1801);
nor U2227 (N_2227,N_1689,N_1891);
nor U2228 (N_2228,N_1459,N_1916);
and U2229 (N_2229,N_1339,N_1784);
nor U2230 (N_2230,N_1179,N_1485);
or U2231 (N_2231,N_1514,N_1414);
or U2232 (N_2232,N_1497,N_1823);
nor U2233 (N_2233,N_1279,N_1593);
or U2234 (N_2234,N_1117,N_1782);
nand U2235 (N_2235,N_1716,N_1142);
or U2236 (N_2236,N_1362,N_1938);
nor U2237 (N_2237,N_1642,N_1551);
xnor U2238 (N_2238,N_1219,N_1862);
or U2239 (N_2239,N_1807,N_1320);
and U2240 (N_2240,N_1670,N_1615);
and U2241 (N_2241,N_1863,N_1930);
nand U2242 (N_2242,N_1385,N_1492);
or U2243 (N_2243,N_1346,N_1109);
nor U2244 (N_2244,N_1208,N_1217);
nor U2245 (N_2245,N_1650,N_1448);
nor U2246 (N_2246,N_1908,N_1561);
nand U2247 (N_2247,N_1491,N_1434);
and U2248 (N_2248,N_1039,N_1159);
or U2249 (N_2249,N_1372,N_1892);
and U2250 (N_2250,N_1592,N_1022);
xnor U2251 (N_2251,N_1833,N_1740);
xor U2252 (N_2252,N_1798,N_1542);
nor U2253 (N_2253,N_1185,N_1849);
xnor U2254 (N_2254,N_1348,N_1297);
nor U2255 (N_2255,N_1559,N_1544);
nor U2256 (N_2256,N_1027,N_1272);
nand U2257 (N_2257,N_1864,N_1691);
or U2258 (N_2258,N_1200,N_1243);
nand U2259 (N_2259,N_1909,N_1211);
nor U2260 (N_2260,N_1867,N_1259);
or U2261 (N_2261,N_1375,N_1599);
or U2262 (N_2262,N_1602,N_1788);
nor U2263 (N_2263,N_1594,N_1890);
and U2264 (N_2264,N_1712,N_1143);
nor U2265 (N_2265,N_1426,N_1840);
nand U2266 (N_2266,N_1894,N_1006);
nand U2267 (N_2267,N_1610,N_1402);
nor U2268 (N_2268,N_1164,N_1493);
and U2269 (N_2269,N_1578,N_1172);
and U2270 (N_2270,N_1695,N_1035);
nand U2271 (N_2271,N_1030,N_1796);
nand U2272 (N_2272,N_1270,N_1218);
and U2273 (N_2273,N_1265,N_1859);
nand U2274 (N_2274,N_1343,N_1193);
or U2275 (N_2275,N_1842,N_1353);
nand U2276 (N_2276,N_1477,N_1406);
and U2277 (N_2277,N_1713,N_1519);
nand U2278 (N_2278,N_1671,N_1967);
nor U2279 (N_2279,N_1273,N_1411);
nor U2280 (N_2280,N_1165,N_1205);
and U2281 (N_2281,N_1877,N_1024);
and U2282 (N_2282,N_1120,N_1648);
and U2283 (N_2283,N_1382,N_1939);
or U2284 (N_2284,N_1814,N_1962);
nor U2285 (N_2285,N_1194,N_1415);
nand U2286 (N_2286,N_1242,N_1720);
nand U2287 (N_2287,N_1388,N_1832);
or U2288 (N_2288,N_1189,N_1227);
nand U2289 (N_2289,N_1020,N_1263);
and U2290 (N_2290,N_1957,N_1944);
nor U2291 (N_2291,N_1780,N_1504);
or U2292 (N_2292,N_1741,N_1746);
or U2293 (N_2293,N_1676,N_1268);
or U2294 (N_2294,N_1257,N_1460);
or U2295 (N_2295,N_1688,N_1605);
nor U2296 (N_2296,N_1515,N_1947);
nor U2297 (N_2297,N_1565,N_1802);
and U2298 (N_2298,N_1755,N_1816);
and U2299 (N_2299,N_1449,N_1190);
or U2300 (N_2300,N_1747,N_1173);
and U2301 (N_2301,N_1638,N_1654);
nor U2302 (N_2302,N_1230,N_1457);
nand U2303 (N_2303,N_1960,N_1288);
and U2304 (N_2304,N_1013,N_1516);
or U2305 (N_2305,N_1977,N_1181);
nand U2306 (N_2306,N_1774,N_1483);
nand U2307 (N_2307,N_1300,N_1794);
nor U2308 (N_2308,N_1398,N_1247);
xor U2309 (N_2309,N_1453,N_1777);
or U2310 (N_2310,N_1010,N_1984);
xor U2311 (N_2311,N_1387,N_1925);
nor U2312 (N_2312,N_1308,N_1662);
nor U2313 (N_2313,N_1646,N_1004);
nand U2314 (N_2314,N_1995,N_1931);
or U2315 (N_2315,N_1656,N_1328);
nand U2316 (N_2316,N_1580,N_1769);
or U2317 (N_2317,N_1088,N_1626);
nor U2318 (N_2318,N_1175,N_1822);
nor U2319 (N_2319,N_1336,N_1883);
and U2320 (N_2320,N_1734,N_1567);
and U2321 (N_2321,N_1240,N_1213);
or U2322 (N_2322,N_1563,N_1168);
nand U2323 (N_2323,N_1748,N_1652);
and U2324 (N_2324,N_1873,N_1705);
or U2325 (N_2325,N_1989,N_1698);
nor U2326 (N_2326,N_1160,N_1591);
nand U2327 (N_2327,N_1724,N_1973);
xor U2328 (N_2328,N_1025,N_1430);
or U2329 (N_2329,N_1342,N_1742);
nand U2330 (N_2330,N_1804,N_1911);
and U2331 (N_2331,N_1019,N_1239);
nor U2332 (N_2332,N_1506,N_1018);
xnor U2333 (N_2333,N_1116,N_1377);
nor U2334 (N_2334,N_1260,N_1296);
nor U2335 (N_2335,N_1754,N_1199);
nand U2336 (N_2336,N_1425,N_1651);
and U2337 (N_2337,N_1350,N_1108);
nand U2338 (N_2338,N_1735,N_1568);
xnor U2339 (N_2339,N_1413,N_1463);
nor U2340 (N_2340,N_1598,N_1627);
nand U2341 (N_2341,N_1728,N_1704);
xor U2342 (N_2342,N_1543,N_1530);
nor U2343 (N_2343,N_1433,N_1329);
or U2344 (N_2344,N_1510,N_1225);
and U2345 (N_2345,N_1226,N_1958);
nor U2346 (N_2346,N_1870,N_1826);
or U2347 (N_2347,N_1094,N_1392);
or U2348 (N_2348,N_1919,N_1518);
and U2349 (N_2349,N_1687,N_1180);
and U2350 (N_2350,N_1290,N_1719);
or U2351 (N_2351,N_1956,N_1075);
or U2352 (N_2352,N_1767,N_1373);
nor U2353 (N_2353,N_1487,N_1456);
or U2354 (N_2354,N_1083,N_1702);
nand U2355 (N_2355,N_1498,N_1106);
and U2356 (N_2356,N_1524,N_1469);
xor U2357 (N_2357,N_1401,N_1882);
nor U2358 (N_2358,N_1071,N_1047);
nor U2359 (N_2359,N_1095,N_1797);
or U2360 (N_2360,N_1558,N_1899);
and U2361 (N_2361,N_1963,N_1216);
or U2362 (N_2362,N_1968,N_1961);
xor U2363 (N_2363,N_1246,N_1114);
nor U2364 (N_2364,N_1574,N_1245);
and U2365 (N_2365,N_1885,N_1045);
nor U2366 (N_2366,N_1945,N_1986);
nor U2367 (N_2367,N_1274,N_1644);
or U2368 (N_2368,N_1848,N_1581);
nand U2369 (N_2369,N_1443,N_1163);
nor U2370 (N_2370,N_1471,N_1560);
nor U2371 (N_2371,N_1878,N_1604);
or U2372 (N_2372,N_1757,N_1291);
nand U2373 (N_2373,N_1014,N_1933);
or U2374 (N_2374,N_1806,N_1123);
nor U2375 (N_2375,N_1003,N_1982);
nor U2376 (N_2376,N_1403,N_1145);
or U2377 (N_2377,N_1631,N_1454);
and U2378 (N_2378,N_1462,N_1043);
or U2379 (N_2379,N_1623,N_1011);
nor U2380 (N_2380,N_1738,N_1589);
and U2381 (N_2381,N_1744,N_1085);
and U2382 (N_2382,N_1884,N_1770);
nand U2383 (N_2383,N_1127,N_1000);
xnor U2384 (N_2384,N_1611,N_1452);
and U2385 (N_2385,N_1254,N_1005);
nor U2386 (N_2386,N_1678,N_1233);
nor U2387 (N_2387,N_1325,N_1824);
and U2388 (N_2388,N_1693,N_1858);
and U2389 (N_2389,N_1090,N_1231);
and U2390 (N_2390,N_1618,N_1467);
nor U2391 (N_2391,N_1994,N_1423);
nand U2392 (N_2392,N_1037,N_1313);
nor U2393 (N_2393,N_1906,N_1606);
and U2394 (N_2394,N_1634,N_1838);
nor U2395 (N_2395,N_1441,N_1324);
nand U2396 (N_2396,N_1872,N_1210);
and U2397 (N_2397,N_1846,N_1489);
and U2398 (N_2398,N_1509,N_1283);
nor U2399 (N_2399,N_1622,N_1248);
and U2400 (N_2400,N_1679,N_1993);
or U2401 (N_2401,N_1182,N_1785);
and U2402 (N_2402,N_1051,N_1232);
nand U2403 (N_2403,N_1282,N_1971);
or U2404 (N_2404,N_1521,N_1124);
nand U2405 (N_2405,N_1304,N_1701);
or U2406 (N_2406,N_1547,N_1319);
nand U2407 (N_2407,N_1665,N_1162);
nor U2408 (N_2408,N_1912,N_1235);
and U2409 (N_2409,N_1620,N_1532);
and U2410 (N_2410,N_1786,N_1351);
nand U2411 (N_2411,N_1312,N_1286);
nand U2412 (N_2412,N_1468,N_1096);
and U2413 (N_2413,N_1442,N_1158);
xnor U2414 (N_2414,N_1146,N_1357);
and U2415 (N_2415,N_1429,N_1271);
nand U2416 (N_2416,N_1455,N_1397);
nor U2417 (N_2417,N_1680,N_1549);
nor U2418 (N_2418,N_1575,N_1157);
and U2419 (N_2419,N_1959,N_1851);
nand U2420 (N_2420,N_1659,N_1280);
or U2421 (N_2421,N_1756,N_1793);
or U2422 (N_2422,N_1080,N_1058);
nand U2423 (N_2423,N_1739,N_1081);
nand U2424 (N_2424,N_1238,N_1440);
nor U2425 (N_2425,N_1316,N_1897);
xor U2426 (N_2426,N_1359,N_1275);
and U2427 (N_2427,N_1587,N_1370);
nand U2428 (N_2428,N_1505,N_1643);
nand U2429 (N_2429,N_1431,N_1196);
or U2430 (N_2430,N_1700,N_1953);
nand U2431 (N_2431,N_1323,N_1133);
nand U2432 (N_2432,N_1658,N_1669);
nor U2433 (N_2433,N_1540,N_1820);
nor U2434 (N_2434,N_1552,N_1889);
nor U2435 (N_2435,N_1129,N_1481);
and U2436 (N_2436,N_1266,N_1500);
nor U2437 (N_2437,N_1347,N_1311);
xor U2438 (N_2438,N_1389,N_1555);
nor U2439 (N_2439,N_1386,N_1188);
nor U2440 (N_2440,N_1819,N_1417);
nor U2441 (N_2441,N_1458,N_1224);
xor U2442 (N_2442,N_1461,N_1028);
or U2443 (N_2443,N_1360,N_1783);
nor U2444 (N_2444,N_1790,N_1745);
nand U2445 (N_2445,N_1874,N_1412);
nor U2446 (N_2446,N_1927,N_1853);
or U2447 (N_2447,N_1661,N_1113);
nand U2448 (N_2448,N_1391,N_1099);
and U2449 (N_2449,N_1914,N_1364);
and U2450 (N_2450,N_1478,N_1284);
or U2451 (N_2451,N_1400,N_1983);
nor U2452 (N_2452,N_1427,N_1880);
nand U2453 (N_2453,N_1294,N_1949);
or U2454 (N_2454,N_1333,N_1778);
or U2455 (N_2455,N_1222,N_1473);
nand U2456 (N_2456,N_1063,N_1352);
and U2457 (N_2457,N_1177,N_1600);
nor U2458 (N_2458,N_1153,N_1267);
or U2459 (N_2459,N_1269,N_1718);
nor U2460 (N_2460,N_1432,N_1569);
and U2461 (N_2461,N_1152,N_1390);
xnor U2462 (N_2462,N_1726,N_1723);
nor U2463 (N_2463,N_1122,N_1556);
or U2464 (N_2464,N_1439,N_1950);
and U2465 (N_2465,N_1541,N_1795);
or U2466 (N_2466,N_1302,N_1255);
and U2467 (N_2467,N_1479,N_1074);
xor U2468 (N_2468,N_1380,N_1435);
nand U2469 (N_2469,N_1066,N_1637);
nand U2470 (N_2470,N_1640,N_1009);
nand U2471 (N_2471,N_1753,N_1281);
and U2472 (N_2472,N_1170,N_1121);
or U2473 (N_2473,N_1171,N_1666);
or U2474 (N_2474,N_1923,N_1655);
and U2475 (N_2475,N_1624,N_1512);
or U2476 (N_2476,N_1394,N_1486);
and U2477 (N_2477,N_1621,N_1537);
xor U2478 (N_2478,N_1998,N_1641);
nand U2479 (N_2479,N_1236,N_1056);
nand U2480 (N_2480,N_1677,N_1079);
nand U2481 (N_2481,N_1332,N_1354);
nand U2482 (N_2482,N_1834,N_1126);
nand U2483 (N_2483,N_1301,N_1570);
nor U2484 (N_2484,N_1253,N_1097);
and U2485 (N_2485,N_1828,N_1002);
nand U2486 (N_2486,N_1776,N_1929);
and U2487 (N_2487,N_1446,N_1707);
and U2488 (N_2488,N_1722,N_1907);
and U2489 (N_2489,N_1703,N_1476);
xor U2490 (N_2490,N_1206,N_1685);
or U2491 (N_2491,N_1799,N_1335);
nor U2492 (N_2492,N_1692,N_1407);
and U2493 (N_2493,N_1588,N_1278);
xor U2494 (N_2494,N_1946,N_1663);
xnor U2495 (N_2495,N_1522,N_1915);
and U2496 (N_2496,N_1150,N_1237);
nand U2497 (N_2497,N_1535,N_1383);
nor U2498 (N_2498,N_1033,N_1997);
nor U2499 (N_2499,N_1295,N_1151);
and U2500 (N_2500,N_1584,N_1618);
and U2501 (N_2501,N_1070,N_1067);
nor U2502 (N_2502,N_1950,N_1433);
nor U2503 (N_2503,N_1895,N_1880);
or U2504 (N_2504,N_1069,N_1004);
or U2505 (N_2505,N_1625,N_1765);
nor U2506 (N_2506,N_1645,N_1427);
and U2507 (N_2507,N_1059,N_1946);
nor U2508 (N_2508,N_1840,N_1828);
or U2509 (N_2509,N_1338,N_1318);
nand U2510 (N_2510,N_1269,N_1014);
and U2511 (N_2511,N_1729,N_1574);
nand U2512 (N_2512,N_1455,N_1810);
nor U2513 (N_2513,N_1954,N_1548);
nor U2514 (N_2514,N_1172,N_1826);
and U2515 (N_2515,N_1094,N_1911);
nor U2516 (N_2516,N_1866,N_1403);
and U2517 (N_2517,N_1096,N_1556);
nand U2518 (N_2518,N_1405,N_1379);
or U2519 (N_2519,N_1541,N_1115);
nor U2520 (N_2520,N_1469,N_1997);
nand U2521 (N_2521,N_1061,N_1537);
nand U2522 (N_2522,N_1495,N_1007);
nand U2523 (N_2523,N_1317,N_1007);
nor U2524 (N_2524,N_1779,N_1824);
or U2525 (N_2525,N_1804,N_1129);
nor U2526 (N_2526,N_1702,N_1394);
or U2527 (N_2527,N_1138,N_1171);
and U2528 (N_2528,N_1275,N_1738);
or U2529 (N_2529,N_1873,N_1468);
nor U2530 (N_2530,N_1547,N_1247);
and U2531 (N_2531,N_1499,N_1495);
and U2532 (N_2532,N_1902,N_1786);
xnor U2533 (N_2533,N_1207,N_1744);
nand U2534 (N_2534,N_1463,N_1765);
nand U2535 (N_2535,N_1318,N_1732);
or U2536 (N_2536,N_1739,N_1656);
or U2537 (N_2537,N_1900,N_1035);
and U2538 (N_2538,N_1112,N_1676);
and U2539 (N_2539,N_1241,N_1334);
nor U2540 (N_2540,N_1944,N_1524);
nor U2541 (N_2541,N_1185,N_1184);
nor U2542 (N_2542,N_1187,N_1866);
or U2543 (N_2543,N_1509,N_1677);
and U2544 (N_2544,N_1657,N_1868);
xor U2545 (N_2545,N_1180,N_1882);
xor U2546 (N_2546,N_1316,N_1386);
nor U2547 (N_2547,N_1595,N_1606);
or U2548 (N_2548,N_1280,N_1163);
nor U2549 (N_2549,N_1817,N_1644);
nand U2550 (N_2550,N_1959,N_1452);
and U2551 (N_2551,N_1496,N_1592);
nand U2552 (N_2552,N_1028,N_1268);
nand U2553 (N_2553,N_1130,N_1602);
or U2554 (N_2554,N_1006,N_1031);
or U2555 (N_2555,N_1492,N_1246);
nand U2556 (N_2556,N_1845,N_1279);
or U2557 (N_2557,N_1070,N_1527);
nand U2558 (N_2558,N_1734,N_1305);
nand U2559 (N_2559,N_1430,N_1665);
nor U2560 (N_2560,N_1850,N_1151);
nand U2561 (N_2561,N_1720,N_1285);
nand U2562 (N_2562,N_1504,N_1191);
nor U2563 (N_2563,N_1674,N_1643);
or U2564 (N_2564,N_1220,N_1142);
nor U2565 (N_2565,N_1503,N_1289);
xor U2566 (N_2566,N_1139,N_1836);
xnor U2567 (N_2567,N_1871,N_1578);
or U2568 (N_2568,N_1073,N_1467);
nor U2569 (N_2569,N_1003,N_1884);
nor U2570 (N_2570,N_1604,N_1656);
nand U2571 (N_2571,N_1766,N_1245);
nand U2572 (N_2572,N_1016,N_1055);
nor U2573 (N_2573,N_1639,N_1725);
nand U2574 (N_2574,N_1907,N_1089);
nor U2575 (N_2575,N_1218,N_1619);
nand U2576 (N_2576,N_1939,N_1736);
xnor U2577 (N_2577,N_1248,N_1610);
and U2578 (N_2578,N_1906,N_1507);
xnor U2579 (N_2579,N_1025,N_1803);
nor U2580 (N_2580,N_1758,N_1914);
nand U2581 (N_2581,N_1919,N_1764);
nor U2582 (N_2582,N_1323,N_1590);
nand U2583 (N_2583,N_1841,N_1048);
nor U2584 (N_2584,N_1802,N_1899);
nor U2585 (N_2585,N_1654,N_1609);
nand U2586 (N_2586,N_1868,N_1008);
nor U2587 (N_2587,N_1110,N_1468);
nand U2588 (N_2588,N_1580,N_1635);
or U2589 (N_2589,N_1024,N_1370);
nand U2590 (N_2590,N_1687,N_1741);
nand U2591 (N_2591,N_1502,N_1797);
or U2592 (N_2592,N_1000,N_1510);
or U2593 (N_2593,N_1768,N_1578);
nand U2594 (N_2594,N_1638,N_1321);
nor U2595 (N_2595,N_1732,N_1206);
xnor U2596 (N_2596,N_1023,N_1940);
nand U2597 (N_2597,N_1072,N_1338);
and U2598 (N_2598,N_1226,N_1916);
nor U2599 (N_2599,N_1743,N_1251);
nor U2600 (N_2600,N_1372,N_1036);
nand U2601 (N_2601,N_1183,N_1167);
nand U2602 (N_2602,N_1376,N_1194);
and U2603 (N_2603,N_1503,N_1314);
and U2604 (N_2604,N_1048,N_1527);
nand U2605 (N_2605,N_1266,N_1345);
nor U2606 (N_2606,N_1809,N_1477);
nor U2607 (N_2607,N_1928,N_1039);
xor U2608 (N_2608,N_1275,N_1662);
or U2609 (N_2609,N_1157,N_1919);
nor U2610 (N_2610,N_1053,N_1882);
or U2611 (N_2611,N_1222,N_1116);
and U2612 (N_2612,N_1892,N_1548);
nand U2613 (N_2613,N_1100,N_1007);
and U2614 (N_2614,N_1445,N_1937);
or U2615 (N_2615,N_1479,N_1119);
nor U2616 (N_2616,N_1189,N_1600);
and U2617 (N_2617,N_1236,N_1590);
nand U2618 (N_2618,N_1897,N_1265);
or U2619 (N_2619,N_1339,N_1801);
xnor U2620 (N_2620,N_1557,N_1133);
nand U2621 (N_2621,N_1721,N_1558);
xnor U2622 (N_2622,N_1550,N_1952);
nor U2623 (N_2623,N_1481,N_1487);
xnor U2624 (N_2624,N_1722,N_1447);
nand U2625 (N_2625,N_1291,N_1370);
or U2626 (N_2626,N_1106,N_1780);
and U2627 (N_2627,N_1690,N_1298);
nor U2628 (N_2628,N_1963,N_1650);
nor U2629 (N_2629,N_1857,N_1294);
nor U2630 (N_2630,N_1261,N_1830);
nor U2631 (N_2631,N_1505,N_1965);
nand U2632 (N_2632,N_1517,N_1799);
nor U2633 (N_2633,N_1558,N_1207);
xor U2634 (N_2634,N_1519,N_1649);
xnor U2635 (N_2635,N_1721,N_1711);
nor U2636 (N_2636,N_1861,N_1651);
nor U2637 (N_2637,N_1092,N_1854);
or U2638 (N_2638,N_1611,N_1911);
nor U2639 (N_2639,N_1236,N_1605);
or U2640 (N_2640,N_1215,N_1061);
and U2641 (N_2641,N_1678,N_1708);
nor U2642 (N_2642,N_1799,N_1917);
and U2643 (N_2643,N_1182,N_1580);
nand U2644 (N_2644,N_1642,N_1289);
xor U2645 (N_2645,N_1911,N_1901);
nand U2646 (N_2646,N_1721,N_1593);
or U2647 (N_2647,N_1177,N_1923);
and U2648 (N_2648,N_1700,N_1278);
and U2649 (N_2649,N_1799,N_1248);
nand U2650 (N_2650,N_1222,N_1374);
nand U2651 (N_2651,N_1019,N_1716);
nor U2652 (N_2652,N_1527,N_1716);
nand U2653 (N_2653,N_1526,N_1751);
nand U2654 (N_2654,N_1954,N_1597);
and U2655 (N_2655,N_1281,N_1702);
and U2656 (N_2656,N_1289,N_1329);
or U2657 (N_2657,N_1227,N_1942);
nor U2658 (N_2658,N_1429,N_1171);
and U2659 (N_2659,N_1134,N_1631);
or U2660 (N_2660,N_1295,N_1118);
and U2661 (N_2661,N_1149,N_1510);
nor U2662 (N_2662,N_1978,N_1361);
nor U2663 (N_2663,N_1759,N_1211);
nor U2664 (N_2664,N_1990,N_1248);
and U2665 (N_2665,N_1552,N_1414);
xor U2666 (N_2666,N_1327,N_1344);
nor U2667 (N_2667,N_1766,N_1079);
nor U2668 (N_2668,N_1227,N_1322);
and U2669 (N_2669,N_1171,N_1679);
and U2670 (N_2670,N_1746,N_1407);
and U2671 (N_2671,N_1476,N_1056);
nor U2672 (N_2672,N_1351,N_1785);
nor U2673 (N_2673,N_1104,N_1364);
nor U2674 (N_2674,N_1470,N_1983);
nor U2675 (N_2675,N_1183,N_1261);
and U2676 (N_2676,N_1179,N_1984);
nand U2677 (N_2677,N_1020,N_1984);
nand U2678 (N_2678,N_1103,N_1642);
and U2679 (N_2679,N_1348,N_1553);
nor U2680 (N_2680,N_1386,N_1520);
xor U2681 (N_2681,N_1483,N_1462);
nand U2682 (N_2682,N_1615,N_1540);
or U2683 (N_2683,N_1578,N_1135);
nor U2684 (N_2684,N_1233,N_1929);
nand U2685 (N_2685,N_1513,N_1922);
nand U2686 (N_2686,N_1239,N_1875);
and U2687 (N_2687,N_1653,N_1004);
or U2688 (N_2688,N_1484,N_1583);
nor U2689 (N_2689,N_1801,N_1510);
or U2690 (N_2690,N_1854,N_1586);
nor U2691 (N_2691,N_1137,N_1864);
or U2692 (N_2692,N_1338,N_1734);
nand U2693 (N_2693,N_1253,N_1645);
and U2694 (N_2694,N_1373,N_1001);
nor U2695 (N_2695,N_1657,N_1742);
and U2696 (N_2696,N_1696,N_1582);
nor U2697 (N_2697,N_1178,N_1686);
and U2698 (N_2698,N_1831,N_1663);
and U2699 (N_2699,N_1209,N_1932);
nand U2700 (N_2700,N_1628,N_1342);
nand U2701 (N_2701,N_1407,N_1072);
and U2702 (N_2702,N_1106,N_1839);
or U2703 (N_2703,N_1363,N_1531);
and U2704 (N_2704,N_1488,N_1503);
nor U2705 (N_2705,N_1857,N_1456);
or U2706 (N_2706,N_1273,N_1541);
and U2707 (N_2707,N_1057,N_1867);
or U2708 (N_2708,N_1767,N_1549);
and U2709 (N_2709,N_1958,N_1512);
or U2710 (N_2710,N_1500,N_1345);
xor U2711 (N_2711,N_1341,N_1815);
or U2712 (N_2712,N_1558,N_1406);
and U2713 (N_2713,N_1770,N_1606);
and U2714 (N_2714,N_1237,N_1905);
xor U2715 (N_2715,N_1295,N_1071);
or U2716 (N_2716,N_1195,N_1370);
xnor U2717 (N_2717,N_1811,N_1647);
and U2718 (N_2718,N_1844,N_1682);
and U2719 (N_2719,N_1482,N_1563);
nor U2720 (N_2720,N_1325,N_1721);
nand U2721 (N_2721,N_1022,N_1799);
nor U2722 (N_2722,N_1569,N_1220);
nand U2723 (N_2723,N_1830,N_1007);
and U2724 (N_2724,N_1834,N_1037);
or U2725 (N_2725,N_1578,N_1218);
or U2726 (N_2726,N_1084,N_1827);
or U2727 (N_2727,N_1186,N_1737);
and U2728 (N_2728,N_1739,N_1002);
and U2729 (N_2729,N_1873,N_1700);
or U2730 (N_2730,N_1651,N_1998);
and U2731 (N_2731,N_1201,N_1664);
or U2732 (N_2732,N_1518,N_1259);
and U2733 (N_2733,N_1808,N_1224);
or U2734 (N_2734,N_1830,N_1082);
or U2735 (N_2735,N_1788,N_1693);
and U2736 (N_2736,N_1794,N_1946);
or U2737 (N_2737,N_1716,N_1553);
and U2738 (N_2738,N_1120,N_1097);
and U2739 (N_2739,N_1237,N_1338);
nor U2740 (N_2740,N_1693,N_1848);
nor U2741 (N_2741,N_1484,N_1166);
or U2742 (N_2742,N_1605,N_1868);
xnor U2743 (N_2743,N_1594,N_1200);
nand U2744 (N_2744,N_1796,N_1086);
xnor U2745 (N_2745,N_1461,N_1217);
and U2746 (N_2746,N_1669,N_1527);
nand U2747 (N_2747,N_1534,N_1716);
or U2748 (N_2748,N_1685,N_1213);
nor U2749 (N_2749,N_1894,N_1316);
nor U2750 (N_2750,N_1279,N_1539);
nor U2751 (N_2751,N_1072,N_1910);
nand U2752 (N_2752,N_1110,N_1050);
or U2753 (N_2753,N_1521,N_1833);
and U2754 (N_2754,N_1785,N_1663);
nand U2755 (N_2755,N_1118,N_1671);
nand U2756 (N_2756,N_1183,N_1184);
nor U2757 (N_2757,N_1164,N_1885);
or U2758 (N_2758,N_1813,N_1055);
and U2759 (N_2759,N_1037,N_1332);
and U2760 (N_2760,N_1318,N_1814);
nor U2761 (N_2761,N_1001,N_1070);
and U2762 (N_2762,N_1279,N_1938);
xnor U2763 (N_2763,N_1799,N_1395);
or U2764 (N_2764,N_1495,N_1595);
nand U2765 (N_2765,N_1076,N_1380);
xor U2766 (N_2766,N_1999,N_1117);
xor U2767 (N_2767,N_1548,N_1894);
nand U2768 (N_2768,N_1648,N_1360);
xnor U2769 (N_2769,N_1583,N_1470);
nand U2770 (N_2770,N_1296,N_1498);
and U2771 (N_2771,N_1701,N_1640);
and U2772 (N_2772,N_1371,N_1708);
and U2773 (N_2773,N_1071,N_1461);
nand U2774 (N_2774,N_1682,N_1642);
xnor U2775 (N_2775,N_1953,N_1395);
or U2776 (N_2776,N_1335,N_1213);
xnor U2777 (N_2777,N_1736,N_1537);
xor U2778 (N_2778,N_1615,N_1285);
nor U2779 (N_2779,N_1137,N_1866);
nand U2780 (N_2780,N_1323,N_1435);
nor U2781 (N_2781,N_1346,N_1844);
or U2782 (N_2782,N_1698,N_1408);
or U2783 (N_2783,N_1318,N_1093);
and U2784 (N_2784,N_1003,N_1545);
or U2785 (N_2785,N_1851,N_1515);
and U2786 (N_2786,N_1186,N_1843);
nand U2787 (N_2787,N_1783,N_1790);
or U2788 (N_2788,N_1924,N_1922);
xor U2789 (N_2789,N_1362,N_1332);
and U2790 (N_2790,N_1364,N_1437);
nor U2791 (N_2791,N_1628,N_1117);
and U2792 (N_2792,N_1739,N_1076);
or U2793 (N_2793,N_1419,N_1504);
and U2794 (N_2794,N_1203,N_1430);
nor U2795 (N_2795,N_1057,N_1948);
nand U2796 (N_2796,N_1783,N_1182);
nor U2797 (N_2797,N_1352,N_1964);
and U2798 (N_2798,N_1841,N_1495);
nor U2799 (N_2799,N_1736,N_1762);
and U2800 (N_2800,N_1741,N_1705);
and U2801 (N_2801,N_1923,N_1134);
nor U2802 (N_2802,N_1310,N_1546);
or U2803 (N_2803,N_1792,N_1446);
and U2804 (N_2804,N_1750,N_1113);
nand U2805 (N_2805,N_1424,N_1692);
nand U2806 (N_2806,N_1637,N_1672);
and U2807 (N_2807,N_1658,N_1697);
or U2808 (N_2808,N_1172,N_1361);
nand U2809 (N_2809,N_1681,N_1653);
or U2810 (N_2810,N_1331,N_1613);
nand U2811 (N_2811,N_1777,N_1629);
xnor U2812 (N_2812,N_1699,N_1837);
or U2813 (N_2813,N_1262,N_1193);
nor U2814 (N_2814,N_1407,N_1166);
and U2815 (N_2815,N_1312,N_1997);
or U2816 (N_2816,N_1455,N_1578);
nand U2817 (N_2817,N_1881,N_1044);
nor U2818 (N_2818,N_1639,N_1563);
or U2819 (N_2819,N_1330,N_1958);
and U2820 (N_2820,N_1639,N_1034);
nand U2821 (N_2821,N_1472,N_1029);
xnor U2822 (N_2822,N_1200,N_1400);
xnor U2823 (N_2823,N_1448,N_1462);
and U2824 (N_2824,N_1115,N_1221);
or U2825 (N_2825,N_1674,N_1858);
nand U2826 (N_2826,N_1015,N_1236);
or U2827 (N_2827,N_1898,N_1160);
nand U2828 (N_2828,N_1586,N_1364);
nand U2829 (N_2829,N_1638,N_1714);
nor U2830 (N_2830,N_1423,N_1512);
nor U2831 (N_2831,N_1518,N_1730);
nand U2832 (N_2832,N_1615,N_1037);
and U2833 (N_2833,N_1709,N_1471);
or U2834 (N_2834,N_1658,N_1684);
xnor U2835 (N_2835,N_1866,N_1438);
and U2836 (N_2836,N_1242,N_1028);
xnor U2837 (N_2837,N_1517,N_1939);
nand U2838 (N_2838,N_1552,N_1954);
nand U2839 (N_2839,N_1591,N_1240);
xnor U2840 (N_2840,N_1218,N_1324);
nand U2841 (N_2841,N_1463,N_1652);
and U2842 (N_2842,N_1593,N_1381);
xnor U2843 (N_2843,N_1498,N_1729);
or U2844 (N_2844,N_1707,N_1177);
nand U2845 (N_2845,N_1722,N_1817);
or U2846 (N_2846,N_1706,N_1770);
nor U2847 (N_2847,N_1965,N_1843);
xor U2848 (N_2848,N_1564,N_1585);
and U2849 (N_2849,N_1427,N_1396);
nor U2850 (N_2850,N_1984,N_1769);
nor U2851 (N_2851,N_1163,N_1449);
and U2852 (N_2852,N_1281,N_1539);
nand U2853 (N_2853,N_1062,N_1412);
nor U2854 (N_2854,N_1635,N_1850);
or U2855 (N_2855,N_1396,N_1576);
xnor U2856 (N_2856,N_1126,N_1071);
nor U2857 (N_2857,N_1367,N_1795);
nand U2858 (N_2858,N_1160,N_1431);
or U2859 (N_2859,N_1974,N_1743);
nor U2860 (N_2860,N_1300,N_1159);
and U2861 (N_2861,N_1308,N_1818);
nand U2862 (N_2862,N_1447,N_1192);
nand U2863 (N_2863,N_1632,N_1090);
nand U2864 (N_2864,N_1168,N_1034);
and U2865 (N_2865,N_1585,N_1061);
nor U2866 (N_2866,N_1157,N_1268);
xnor U2867 (N_2867,N_1122,N_1193);
and U2868 (N_2868,N_1881,N_1115);
nor U2869 (N_2869,N_1601,N_1764);
nor U2870 (N_2870,N_1394,N_1636);
nor U2871 (N_2871,N_1933,N_1268);
and U2872 (N_2872,N_1253,N_1488);
and U2873 (N_2873,N_1926,N_1546);
xnor U2874 (N_2874,N_1984,N_1193);
and U2875 (N_2875,N_1740,N_1196);
nand U2876 (N_2876,N_1244,N_1547);
nor U2877 (N_2877,N_1303,N_1296);
nand U2878 (N_2878,N_1793,N_1274);
or U2879 (N_2879,N_1346,N_1386);
nand U2880 (N_2880,N_1620,N_1350);
nor U2881 (N_2881,N_1397,N_1551);
and U2882 (N_2882,N_1015,N_1410);
or U2883 (N_2883,N_1251,N_1262);
nand U2884 (N_2884,N_1984,N_1886);
nor U2885 (N_2885,N_1784,N_1110);
or U2886 (N_2886,N_1210,N_1931);
or U2887 (N_2887,N_1899,N_1145);
or U2888 (N_2888,N_1509,N_1687);
and U2889 (N_2889,N_1568,N_1679);
nand U2890 (N_2890,N_1885,N_1388);
and U2891 (N_2891,N_1721,N_1512);
and U2892 (N_2892,N_1219,N_1609);
and U2893 (N_2893,N_1330,N_1924);
or U2894 (N_2894,N_1359,N_1282);
and U2895 (N_2895,N_1188,N_1371);
nor U2896 (N_2896,N_1144,N_1339);
xor U2897 (N_2897,N_1874,N_1582);
xnor U2898 (N_2898,N_1516,N_1303);
nand U2899 (N_2899,N_1135,N_1223);
and U2900 (N_2900,N_1913,N_1587);
nand U2901 (N_2901,N_1297,N_1129);
nand U2902 (N_2902,N_1141,N_1570);
nand U2903 (N_2903,N_1170,N_1595);
or U2904 (N_2904,N_1357,N_1383);
nand U2905 (N_2905,N_1379,N_1940);
nor U2906 (N_2906,N_1394,N_1006);
nand U2907 (N_2907,N_1955,N_1980);
nor U2908 (N_2908,N_1971,N_1621);
and U2909 (N_2909,N_1949,N_1877);
nand U2910 (N_2910,N_1809,N_1419);
xnor U2911 (N_2911,N_1801,N_1670);
or U2912 (N_2912,N_1281,N_1671);
nand U2913 (N_2913,N_1505,N_1658);
and U2914 (N_2914,N_1056,N_1280);
and U2915 (N_2915,N_1502,N_1791);
nor U2916 (N_2916,N_1099,N_1837);
nand U2917 (N_2917,N_1333,N_1946);
nand U2918 (N_2918,N_1366,N_1388);
and U2919 (N_2919,N_1261,N_1302);
or U2920 (N_2920,N_1845,N_1425);
or U2921 (N_2921,N_1915,N_1715);
and U2922 (N_2922,N_1923,N_1665);
nor U2923 (N_2923,N_1726,N_1076);
and U2924 (N_2924,N_1118,N_1904);
xnor U2925 (N_2925,N_1810,N_1740);
or U2926 (N_2926,N_1682,N_1766);
or U2927 (N_2927,N_1971,N_1230);
and U2928 (N_2928,N_1742,N_1238);
and U2929 (N_2929,N_1783,N_1982);
nand U2930 (N_2930,N_1192,N_1939);
or U2931 (N_2931,N_1627,N_1772);
xnor U2932 (N_2932,N_1304,N_1690);
and U2933 (N_2933,N_1828,N_1597);
or U2934 (N_2934,N_1561,N_1006);
nand U2935 (N_2935,N_1371,N_1161);
or U2936 (N_2936,N_1001,N_1713);
and U2937 (N_2937,N_1456,N_1898);
nor U2938 (N_2938,N_1963,N_1774);
nor U2939 (N_2939,N_1728,N_1602);
nor U2940 (N_2940,N_1565,N_1862);
xor U2941 (N_2941,N_1933,N_1993);
xor U2942 (N_2942,N_1114,N_1238);
nand U2943 (N_2943,N_1107,N_1386);
xor U2944 (N_2944,N_1411,N_1915);
nor U2945 (N_2945,N_1504,N_1988);
and U2946 (N_2946,N_1549,N_1709);
nand U2947 (N_2947,N_1988,N_1758);
nand U2948 (N_2948,N_1673,N_1726);
and U2949 (N_2949,N_1904,N_1563);
nand U2950 (N_2950,N_1260,N_1428);
and U2951 (N_2951,N_1072,N_1540);
nor U2952 (N_2952,N_1452,N_1989);
nand U2953 (N_2953,N_1323,N_1038);
and U2954 (N_2954,N_1312,N_1002);
or U2955 (N_2955,N_1738,N_1684);
xor U2956 (N_2956,N_1353,N_1594);
and U2957 (N_2957,N_1977,N_1795);
and U2958 (N_2958,N_1512,N_1482);
and U2959 (N_2959,N_1010,N_1554);
nor U2960 (N_2960,N_1544,N_1533);
and U2961 (N_2961,N_1656,N_1003);
nand U2962 (N_2962,N_1105,N_1011);
or U2963 (N_2963,N_1383,N_1076);
or U2964 (N_2964,N_1023,N_1473);
nor U2965 (N_2965,N_1232,N_1669);
xnor U2966 (N_2966,N_1296,N_1535);
nand U2967 (N_2967,N_1259,N_1082);
nor U2968 (N_2968,N_1046,N_1414);
nand U2969 (N_2969,N_1251,N_1226);
nand U2970 (N_2970,N_1620,N_1927);
and U2971 (N_2971,N_1306,N_1736);
nand U2972 (N_2972,N_1575,N_1202);
nor U2973 (N_2973,N_1589,N_1617);
and U2974 (N_2974,N_1256,N_1615);
and U2975 (N_2975,N_1589,N_1817);
nor U2976 (N_2976,N_1134,N_1606);
nand U2977 (N_2977,N_1719,N_1678);
nor U2978 (N_2978,N_1419,N_1824);
nor U2979 (N_2979,N_1719,N_1442);
and U2980 (N_2980,N_1861,N_1383);
nor U2981 (N_2981,N_1352,N_1855);
nor U2982 (N_2982,N_1072,N_1288);
nand U2983 (N_2983,N_1985,N_1157);
or U2984 (N_2984,N_1183,N_1732);
or U2985 (N_2985,N_1522,N_1258);
and U2986 (N_2986,N_1276,N_1736);
nor U2987 (N_2987,N_1713,N_1594);
or U2988 (N_2988,N_1167,N_1452);
and U2989 (N_2989,N_1847,N_1257);
or U2990 (N_2990,N_1392,N_1340);
nor U2991 (N_2991,N_1335,N_1148);
and U2992 (N_2992,N_1950,N_1720);
nor U2993 (N_2993,N_1757,N_1388);
nand U2994 (N_2994,N_1085,N_1636);
nor U2995 (N_2995,N_1826,N_1318);
and U2996 (N_2996,N_1575,N_1147);
nand U2997 (N_2997,N_1159,N_1708);
xnor U2998 (N_2998,N_1879,N_1526);
nand U2999 (N_2999,N_1498,N_1849);
nand U3000 (N_3000,N_2966,N_2533);
nor U3001 (N_3001,N_2945,N_2706);
nor U3002 (N_3002,N_2215,N_2852);
nor U3003 (N_3003,N_2965,N_2885);
nor U3004 (N_3004,N_2336,N_2057);
nand U3005 (N_3005,N_2012,N_2402);
nor U3006 (N_3006,N_2924,N_2120);
nor U3007 (N_3007,N_2708,N_2812);
nand U3008 (N_3008,N_2566,N_2937);
nand U3009 (N_3009,N_2488,N_2356);
xnor U3010 (N_3010,N_2574,N_2483);
nor U3011 (N_3011,N_2561,N_2037);
nor U3012 (N_3012,N_2839,N_2844);
xor U3013 (N_3013,N_2276,N_2711);
and U3014 (N_3014,N_2605,N_2280);
and U3015 (N_3015,N_2415,N_2775);
nand U3016 (N_3016,N_2648,N_2505);
or U3017 (N_3017,N_2727,N_2870);
nor U3018 (N_3018,N_2218,N_2432);
or U3019 (N_3019,N_2419,N_2498);
and U3020 (N_3020,N_2657,N_2075);
xor U3021 (N_3021,N_2278,N_2100);
and U3022 (N_3022,N_2284,N_2990);
xnor U3023 (N_3023,N_2859,N_2548);
and U3024 (N_3024,N_2763,N_2472);
or U3025 (N_3025,N_2320,N_2433);
xor U3026 (N_3026,N_2802,N_2459);
nand U3027 (N_3027,N_2537,N_2429);
and U3028 (N_3028,N_2880,N_2510);
nor U3029 (N_3029,N_2744,N_2204);
or U3030 (N_3030,N_2492,N_2974);
and U3031 (N_3031,N_2266,N_2261);
xnor U3032 (N_3032,N_2017,N_2868);
and U3033 (N_3033,N_2239,N_2353);
or U3034 (N_3034,N_2248,N_2555);
and U3035 (N_3035,N_2940,N_2287);
nand U3036 (N_3036,N_2993,N_2190);
nor U3037 (N_3037,N_2560,N_2346);
and U3038 (N_3038,N_2211,N_2442);
or U3039 (N_3039,N_2947,N_2213);
or U3040 (N_3040,N_2138,N_2318);
and U3041 (N_3041,N_2831,N_2104);
or U3042 (N_3042,N_2473,N_2665);
and U3043 (N_3043,N_2748,N_2692);
nor U3044 (N_3044,N_2541,N_2134);
nand U3045 (N_3045,N_2717,N_2712);
nor U3046 (N_3046,N_2165,N_2203);
and U3047 (N_3047,N_2809,N_2580);
and U3048 (N_3048,N_2932,N_2301);
or U3049 (N_3049,N_2998,N_2002);
nor U3050 (N_3050,N_2450,N_2506);
or U3051 (N_3051,N_2316,N_2615);
nor U3052 (N_3052,N_2270,N_2073);
xor U3053 (N_3053,N_2245,N_2293);
and U3054 (N_3054,N_2798,N_2901);
or U3055 (N_3055,N_2647,N_2520);
xor U3056 (N_3056,N_2854,N_2801);
or U3057 (N_3057,N_2166,N_2761);
or U3058 (N_3058,N_2867,N_2219);
and U3059 (N_3059,N_2011,N_2919);
and U3060 (N_3060,N_2311,N_2992);
nand U3061 (N_3061,N_2837,N_2710);
and U3062 (N_3062,N_2500,N_2179);
or U3063 (N_3063,N_2289,N_2093);
and U3064 (N_3064,N_2395,N_2968);
and U3065 (N_3065,N_2825,N_2034);
nand U3066 (N_3066,N_2110,N_2550);
or U3067 (N_3067,N_2299,N_2896);
xor U3068 (N_3068,N_2344,N_2341);
and U3069 (N_3069,N_2645,N_2600);
and U3070 (N_3070,N_2026,N_2015);
nor U3071 (N_3071,N_2222,N_2479);
and U3072 (N_3072,N_2961,N_2051);
or U3073 (N_3073,N_2391,N_2599);
or U3074 (N_3074,N_2610,N_2258);
xnor U3075 (N_3075,N_2275,N_2879);
nand U3076 (N_3076,N_2379,N_2206);
or U3077 (N_3077,N_2791,N_2770);
or U3078 (N_3078,N_2742,N_2092);
nand U3079 (N_3079,N_2119,N_2697);
nor U3080 (N_3080,N_2385,N_2753);
nor U3081 (N_3081,N_2991,N_2928);
nand U3082 (N_3082,N_2660,N_2514);
and U3083 (N_3083,N_2833,N_2490);
and U3084 (N_3084,N_2070,N_2489);
or U3085 (N_3085,N_2519,N_2944);
and U3086 (N_3086,N_2412,N_2332);
nor U3087 (N_3087,N_2659,N_2914);
nor U3088 (N_3088,N_2970,N_2564);
nand U3089 (N_3089,N_2283,N_2487);
and U3090 (N_3090,N_2513,N_2670);
or U3091 (N_3091,N_2797,N_2237);
and U3092 (N_3092,N_2951,N_2458);
or U3093 (N_3093,N_2535,N_2756);
or U3094 (N_3094,N_2335,N_2116);
nor U3095 (N_3095,N_2875,N_2155);
nor U3096 (N_3096,N_2463,N_2277);
xor U3097 (N_3097,N_2347,N_2524);
nor U3098 (N_3098,N_2794,N_2829);
or U3099 (N_3099,N_2554,N_2713);
or U3100 (N_3100,N_2707,N_2021);
nand U3101 (N_3101,N_2027,N_2673);
nor U3102 (N_3102,N_2403,N_2269);
nand U3103 (N_3103,N_2509,N_2544);
and U3104 (N_3104,N_2962,N_2095);
xnor U3105 (N_3105,N_2633,N_2913);
nand U3106 (N_3106,N_2781,N_2004);
and U3107 (N_3107,N_2296,N_2008);
and U3108 (N_3108,N_2223,N_2687);
nand U3109 (N_3109,N_2969,N_2820);
xnor U3110 (N_3110,N_2139,N_2741);
and U3111 (N_3111,N_2934,N_2150);
and U3112 (N_3112,N_2367,N_2661);
nand U3113 (N_3113,N_2076,N_2387);
xor U3114 (N_3114,N_2251,N_2634);
nand U3115 (N_3115,N_2842,N_2495);
or U3116 (N_3116,N_2586,N_2153);
or U3117 (N_3117,N_2396,N_2098);
nor U3118 (N_3118,N_2899,N_2230);
nand U3119 (N_3119,N_2579,N_2405);
or U3120 (N_3120,N_2639,N_2699);
or U3121 (N_3121,N_2131,N_2516);
nor U3122 (N_3122,N_2908,N_2694);
or U3123 (N_3123,N_2935,N_2654);
nor U3124 (N_3124,N_2570,N_2136);
xor U3125 (N_3125,N_2228,N_2421);
xnor U3126 (N_3126,N_2752,N_2771);
and U3127 (N_3127,N_2815,N_2983);
and U3128 (N_3128,N_2994,N_2351);
nand U3129 (N_3129,N_2929,N_2381);
nor U3130 (N_3130,N_2760,N_2822);
nor U3131 (N_3131,N_2024,N_2973);
or U3132 (N_3132,N_2397,N_2900);
or U3133 (N_3133,N_2613,N_2091);
nand U3134 (N_3134,N_2588,N_2321);
nand U3135 (N_3135,N_2111,N_2077);
nor U3136 (N_3136,N_2804,N_2740);
xor U3137 (N_3137,N_2172,N_2591);
or U3138 (N_3138,N_2894,N_2679);
and U3139 (N_3139,N_2714,N_2467);
and U3140 (N_3140,N_2193,N_2062);
and U3141 (N_3141,N_2089,N_2511);
nand U3142 (N_3142,N_2902,N_2486);
xor U3143 (N_3143,N_2413,N_2049);
or U3144 (N_3144,N_2036,N_2773);
nor U3145 (N_3145,N_2194,N_2658);
and U3146 (N_3146,N_2572,N_2468);
nand U3147 (N_3147,N_2959,N_2783);
nand U3148 (N_3148,N_2365,N_2662);
nor U3149 (N_3149,N_2217,N_2984);
or U3150 (N_3150,N_2010,N_2841);
and U3151 (N_3151,N_2149,N_2264);
nor U3152 (N_3152,N_2762,N_2102);
or U3153 (N_3153,N_2071,N_2078);
nand U3154 (N_3154,N_2227,N_2652);
nor U3155 (N_3155,N_2543,N_2826);
or U3156 (N_3156,N_2305,N_2766);
and U3157 (N_3157,N_2986,N_2602);
or U3158 (N_3158,N_2151,N_2470);
or U3159 (N_3159,N_2478,N_2922);
nor U3160 (N_3160,N_2109,N_2627);
xnor U3161 (N_3161,N_2518,N_2680);
or U3162 (N_3162,N_2437,N_2238);
or U3163 (N_3163,N_2916,N_2858);
and U3164 (N_3164,N_2087,N_2625);
nor U3165 (N_3165,N_2001,N_2253);
nand U3166 (N_3166,N_2496,N_2823);
or U3167 (N_3167,N_2866,N_2265);
and U3168 (N_3168,N_2977,N_2569);
nor U3169 (N_3169,N_2754,N_2814);
and U3170 (N_3170,N_2485,N_2632);
nor U3171 (N_3171,N_2236,N_2549);
or U3172 (N_3172,N_2864,N_2274);
and U3173 (N_3173,N_2371,N_2090);
nor U3174 (N_3174,N_2988,N_2624);
nand U3175 (N_3175,N_2884,N_2290);
or U3176 (N_3176,N_2398,N_2592);
nand U3177 (N_3177,N_2214,N_2933);
xor U3178 (N_3178,N_2608,N_2406);
xor U3179 (N_3179,N_2856,N_2512);
or U3180 (N_3180,N_2263,N_2006);
nor U3181 (N_3181,N_2031,N_2016);
nand U3182 (N_3182,N_2127,N_2857);
or U3183 (N_3183,N_2428,N_2246);
and U3184 (N_3184,N_2799,N_2200);
nor U3185 (N_3185,N_2538,N_2949);
and U3186 (N_3186,N_2331,N_2334);
nand U3187 (N_3187,N_2009,N_2782);
nand U3188 (N_3188,N_2898,N_2597);
or U3189 (N_3189,N_2309,N_2701);
or U3190 (N_3190,N_2154,N_2609);
nand U3191 (N_3191,N_2388,N_2147);
nand U3192 (N_3192,N_2435,N_2641);
and U3193 (N_3193,N_2022,N_2018);
or U3194 (N_3194,N_2129,N_2271);
nand U3195 (N_3195,N_2835,N_2521);
nor U3196 (N_3196,N_2803,N_2546);
and U3197 (N_3197,N_2925,N_2558);
xnor U3198 (N_3198,N_2503,N_2065);
nor U3199 (N_3199,N_2917,N_2923);
and U3200 (N_3200,N_2019,N_2040);
and U3201 (N_3201,N_2431,N_2052);
nand U3202 (N_3202,N_2229,N_2596);
or U3203 (N_3203,N_2989,N_2169);
or U3204 (N_3204,N_2501,N_2860);
or U3205 (N_3205,N_2730,N_2853);
xnor U3206 (N_3206,N_2313,N_2855);
nor U3207 (N_3207,N_2173,N_2603);
nor U3208 (N_3208,N_2637,N_2000);
xor U3209 (N_3209,N_2948,N_2436);
or U3210 (N_3210,N_2410,N_2664);
and U3211 (N_3211,N_2577,N_2348);
nand U3212 (N_3212,N_2465,N_2455);
nand U3213 (N_3213,N_2630,N_2618);
nor U3214 (N_3214,N_2359,N_2681);
nor U3215 (N_3215,N_2617,N_2372);
and U3216 (N_3216,N_2553,N_2882);
and U3217 (N_3217,N_2921,N_2210);
nand U3218 (N_3218,N_2556,N_2806);
nor U3219 (N_3219,N_2584,N_2441);
nor U3220 (N_3220,N_2715,N_2863);
nand U3221 (N_3221,N_2593,N_2982);
nor U3222 (N_3222,N_2851,N_2082);
or U3223 (N_3223,N_2281,N_2446);
xnor U3224 (N_3224,N_2423,N_2861);
and U3225 (N_3225,N_2786,N_2523);
nor U3226 (N_3226,N_2143,N_2113);
xor U3227 (N_3227,N_2758,N_2819);
or U3228 (N_3228,N_2105,N_2199);
nand U3229 (N_3229,N_2374,N_2881);
nand U3230 (N_3230,N_2889,N_2705);
nand U3231 (N_3231,N_2207,N_2790);
xnor U3232 (N_3232,N_2757,N_2621);
xor U3233 (N_3233,N_2085,N_2972);
and U3234 (N_3234,N_2045,N_2407);
or U3235 (N_3235,N_2163,N_2643);
nor U3236 (N_3236,N_2747,N_2118);
nand U3237 (N_3237,N_2716,N_2848);
nor U3238 (N_3238,N_2507,N_2152);
and U3239 (N_3239,N_2125,N_2475);
and U3240 (N_3240,N_2447,N_2457);
and U3241 (N_3241,N_2862,N_2130);
nand U3242 (N_3242,N_2912,N_2522);
or U3243 (N_3243,N_2080,N_2267);
nor U3244 (N_3244,N_2499,N_2843);
and U3245 (N_3245,N_2704,N_2939);
nand U3246 (N_3246,N_2640,N_2612);
nand U3247 (N_3247,N_2954,N_2755);
nor U3248 (N_3248,N_2529,N_2517);
and U3249 (N_3249,N_2845,N_2767);
and U3250 (N_3250,N_2997,N_2291);
or U3251 (N_3251,N_2449,N_2128);
or U3252 (N_3252,N_2573,N_2732);
nand U3253 (N_3253,N_2987,N_2191);
xnor U3254 (N_3254,N_2865,N_2849);
nor U3255 (N_3255,N_2482,N_2197);
or U3256 (N_3256,N_2084,N_2174);
or U3257 (N_3257,N_2684,N_2774);
or U3258 (N_3258,N_2779,N_2838);
and U3259 (N_3259,N_2426,N_2349);
nor U3260 (N_3260,N_2025,N_2377);
nand U3261 (N_3261,N_2056,N_2187);
nor U3262 (N_3262,N_2326,N_2375);
and U3263 (N_3263,N_2370,N_2247);
and U3264 (N_3264,N_2067,N_2903);
or U3265 (N_3265,N_2186,N_2185);
nor U3266 (N_3266,N_2133,N_2023);
and U3267 (N_3267,N_2722,N_2038);
nor U3268 (N_3268,N_2642,N_2890);
nor U3269 (N_3269,N_2698,N_2399);
or U3270 (N_3270,N_2832,N_2619);
nor U3271 (N_3271,N_2389,N_2343);
and U3272 (N_3272,N_2156,N_2614);
nor U3273 (N_3273,N_2910,N_2357);
and U3274 (N_3274,N_2672,N_2339);
or U3275 (N_3275,N_2252,N_2552);
nor U3276 (N_3276,N_2623,N_2526);
or U3277 (N_3277,N_2719,N_2481);
nand U3278 (N_3278,N_2562,N_2733);
nor U3279 (N_3279,N_2107,N_2244);
nor U3280 (N_3280,N_2691,N_2836);
nand U3281 (N_3281,N_2099,N_2378);
nand U3282 (N_3282,N_2751,N_2678);
xor U3283 (N_3283,N_2534,N_2655);
nor U3284 (N_3284,N_2392,N_2117);
and U3285 (N_3285,N_2996,N_2976);
xor U3286 (N_3286,N_2995,N_2053);
nor U3287 (N_3287,N_2314,N_2720);
and U3288 (N_3288,N_2587,N_2141);
nand U3289 (N_3289,N_2821,N_2373);
nor U3290 (N_3290,N_2477,N_2693);
xnor U3291 (N_3291,N_2840,N_2279);
nand U3292 (N_3292,N_2094,N_2830);
nand U3293 (N_3293,N_2626,N_2805);
nor U3294 (N_3294,N_2887,N_2338);
nand U3295 (N_3295,N_2536,N_2493);
xnor U3296 (N_3296,N_2622,N_2765);
nor U3297 (N_3297,N_2273,N_2616);
or U3298 (N_3298,N_2323,N_2904);
nand U3299 (N_3299,N_2721,N_2776);
nand U3300 (N_3300,N_2302,N_2003);
and U3301 (N_3301,N_2772,N_2793);
or U3302 (N_3302,N_2736,N_2883);
and U3303 (N_3303,N_2941,N_2649);
and U3304 (N_3304,N_2952,N_2304);
nand U3305 (N_3305,N_2474,N_2257);
nor U3306 (N_3306,N_2540,N_2088);
nor U3307 (N_3307,N_2709,N_2906);
nor U3308 (N_3308,N_2362,N_2328);
and U3309 (N_3309,N_2877,N_2160);
or U3310 (N_3310,N_2956,N_2525);
nand U3311 (N_3311,N_2101,N_2764);
and U3312 (N_3312,N_2508,N_2176);
nand U3313 (N_3313,N_2425,N_2743);
nor U3314 (N_3314,N_2888,N_2096);
and U3315 (N_3315,N_2878,N_2817);
and U3316 (N_3316,N_2083,N_2184);
and U3317 (N_3317,N_2297,N_2629);
or U3318 (N_3318,N_2177,N_2869);
nand U3319 (N_3319,N_2192,N_2241);
nor U3320 (N_3320,N_2559,N_2589);
nand U3321 (N_3321,N_2542,N_2785);
nand U3322 (N_3322,N_2703,N_2233);
xnor U3323 (N_3323,N_2137,N_2386);
and U3324 (N_3324,N_2960,N_2303);
nand U3325 (N_3325,N_2827,N_2445);
nand U3326 (N_3326,N_2943,N_2161);
nand U3327 (N_3327,N_2312,N_2234);
nor U3328 (N_3328,N_2074,N_2063);
or U3329 (N_3329,N_2749,N_2739);
nor U3330 (N_3330,N_2702,N_2581);
nor U3331 (N_3331,N_2050,N_2350);
or U3332 (N_3332,N_2295,N_2690);
and U3333 (N_3333,N_2695,N_2007);
xor U3334 (N_3334,N_2810,N_2180);
nor U3335 (N_3335,N_2568,N_2545);
nand U3336 (N_3336,N_2201,N_2656);
or U3337 (N_3337,N_2847,N_2417);
and U3338 (N_3338,N_2444,N_2604);
nand U3339 (N_3339,N_2033,N_2606);
and U3340 (N_3340,N_2055,N_2850);
nand U3341 (N_3341,N_2121,N_2635);
and U3342 (N_3342,N_2325,N_2807);
nand U3343 (N_3343,N_2380,N_2285);
and U3344 (N_3344,N_2920,N_2737);
or U3345 (N_3345,N_2811,N_2333);
xor U3346 (N_3346,N_2427,N_2808);
or U3347 (N_3347,N_2469,N_2158);
or U3348 (N_3348,N_2162,N_2759);
or U3349 (N_3349,N_2307,N_2726);
nand U3350 (N_3350,N_2787,N_2582);
and U3351 (N_3351,N_2462,N_2746);
and U3352 (N_3352,N_2254,N_2683);
and U3353 (N_3353,N_2300,N_2735);
nor U3354 (N_3354,N_2675,N_2286);
nand U3355 (N_3355,N_2895,N_2931);
nand U3356 (N_3356,N_2813,N_2183);
nor U3357 (N_3357,N_2212,N_2936);
and U3358 (N_3358,N_2926,N_2718);
xor U3359 (N_3359,N_2685,N_2975);
or U3360 (N_3360,N_2409,N_2324);
or U3361 (N_3361,N_2886,N_2985);
nand U3362 (N_3362,N_2414,N_2064);
xor U3363 (N_3363,N_2557,N_2682);
or U3364 (N_3364,N_2393,N_2188);
and U3365 (N_3365,N_2607,N_2368);
nor U3366 (N_3366,N_2376,N_2769);
or U3367 (N_3367,N_2108,N_2337);
or U3368 (N_3368,N_2620,N_2262);
nand U3369 (N_3369,N_2724,N_2216);
and U3370 (N_3370,N_2438,N_2461);
nand U3371 (N_3371,N_2651,N_2358);
nand U3372 (N_3372,N_2310,N_2530);
or U3373 (N_3373,N_2565,N_2443);
nand U3374 (N_3374,N_2598,N_2927);
and U3375 (N_3375,N_2340,N_2964);
nand U3376 (N_3376,N_2824,N_2689);
xor U3377 (N_3377,N_2590,N_2464);
nor U3378 (N_3378,N_2126,N_2272);
and U3379 (N_3379,N_2778,N_2072);
nand U3380 (N_3380,N_2122,N_2322);
or U3381 (N_3381,N_2725,N_2048);
nand U3382 (N_3382,N_2032,N_2114);
or U3383 (N_3383,N_2364,N_2950);
and U3384 (N_3384,N_2221,N_2159);
and U3385 (N_3385,N_2400,N_2170);
or U3386 (N_3386,N_2144,N_2745);
or U3387 (N_3387,N_2422,N_2196);
and U3388 (N_3388,N_2644,N_2575);
and U3389 (N_3389,N_2563,N_2220);
nand U3390 (N_3390,N_2734,N_2355);
or U3391 (N_3391,N_2958,N_2123);
nand U3392 (N_3392,N_2532,N_2167);
xnor U3393 (N_3393,N_2352,N_2384);
nor U3394 (N_3394,N_2918,N_2750);
and U3395 (N_3395,N_2892,N_2366);
or U3396 (N_3396,N_2979,N_2955);
and U3397 (N_3397,N_2306,N_2594);
nand U3398 (N_3398,N_2020,N_2980);
nand U3399 (N_3399,N_2729,N_2484);
nand U3400 (N_3400,N_2646,N_2930);
nor U3401 (N_3401,N_2547,N_2345);
and U3402 (N_3402,N_2891,N_2638);
nor U3403 (N_3403,N_2818,N_2667);
nor U3404 (N_3404,N_2874,N_2595);
nand U3405 (N_3405,N_2728,N_2068);
nand U3406 (N_3406,N_2124,N_2330);
xnor U3407 (N_3407,N_2515,N_2669);
and U3408 (N_3408,N_2873,N_2846);
nor U3409 (N_3409,N_2585,N_2480);
nand U3410 (N_3410,N_2013,N_2157);
or U3411 (N_3411,N_2476,N_2676);
xnor U3412 (N_3412,N_2834,N_2142);
and U3413 (N_3413,N_2394,N_2789);
or U3414 (N_3414,N_2448,N_2942);
nor U3415 (N_3415,N_2209,N_2504);
nand U3416 (N_3416,N_2106,N_2893);
nor U3417 (N_3417,N_2571,N_2058);
nand U3418 (N_3418,N_2567,N_2631);
and U3419 (N_3419,N_2042,N_2451);
nor U3420 (N_3420,N_2416,N_2527);
or U3421 (N_3421,N_2800,N_2653);
nand U3422 (N_3422,N_2418,N_2282);
nor U3423 (N_3423,N_2700,N_2382);
nor U3424 (N_3424,N_2360,N_2601);
or U3425 (N_3425,N_2005,N_2308);
nor U3426 (N_3426,N_2039,N_2576);
nand U3427 (N_3427,N_2046,N_2182);
or U3428 (N_3428,N_2171,N_2029);
and U3429 (N_3429,N_2225,N_2208);
and U3430 (N_3430,N_2872,N_2456);
or U3431 (N_3431,N_2981,N_2369);
and U3432 (N_3432,N_2404,N_2198);
or U3433 (N_3433,N_2240,N_2226);
nand U3434 (N_3434,N_2663,N_2411);
and U3435 (N_3435,N_2784,N_2420);
or U3436 (N_3436,N_2768,N_2361);
and U3437 (N_3437,N_2471,N_2259);
or U3438 (N_3438,N_2909,N_2181);
nor U3439 (N_3439,N_2668,N_2907);
or U3440 (N_3440,N_2401,N_2430);
or U3441 (N_3441,N_2342,N_2650);
xor U3442 (N_3442,N_2828,N_2132);
or U3443 (N_3443,N_2583,N_2439);
nand U3444 (N_3444,N_2168,N_2963);
xor U3445 (N_3445,N_2363,N_2298);
nor U3446 (N_3446,N_2317,N_2636);
nor U3447 (N_3447,N_2175,N_2205);
nor U3448 (N_3448,N_2957,N_2315);
nand U3449 (N_3449,N_2871,N_2014);
and U3450 (N_3450,N_2294,N_2202);
nand U3451 (N_3451,N_2030,N_2466);
or U3452 (N_3452,N_2905,N_2189);
nand U3453 (N_3453,N_2135,N_2971);
nor U3454 (N_3454,N_2059,N_2531);
and U3455 (N_3455,N_2231,N_2319);
or U3456 (N_3456,N_2967,N_2140);
and U3457 (N_3457,N_2723,N_2054);
or U3458 (N_3458,N_2329,N_2383);
xor U3459 (N_3459,N_2164,N_2528);
and U3460 (N_3460,N_2671,N_2060);
nand U3461 (N_3461,N_2677,N_2044);
and U3462 (N_3462,N_2738,N_2497);
nand U3463 (N_3463,N_2327,N_2688);
or U3464 (N_3464,N_2494,N_2103);
or U3465 (N_3465,N_2460,N_2696);
nor U3466 (N_3466,N_2292,N_2453);
xor U3467 (N_3467,N_2674,N_2260);
or U3468 (N_3468,N_2551,N_2146);
and U3469 (N_3469,N_2145,N_2041);
or U3470 (N_3470,N_2081,N_2816);
nor U3471 (N_3471,N_2086,N_2242);
nor U3472 (N_3472,N_2354,N_2491);
nor U3473 (N_3473,N_2796,N_2539);
or U3474 (N_3474,N_2578,N_2978);
or U3475 (N_3475,N_2256,N_2243);
and U3476 (N_3476,N_2946,N_2061);
or U3477 (N_3477,N_2938,N_2148);
nor U3478 (N_3478,N_2731,N_2502);
xor U3479 (N_3479,N_2788,N_2288);
and U3480 (N_3480,N_2452,N_2953);
xnor U3481 (N_3481,N_2043,N_2255);
or U3482 (N_3482,N_2112,N_2795);
nand U3483 (N_3483,N_2047,N_2454);
and U3484 (N_3484,N_2235,N_2408);
xor U3485 (N_3485,N_2232,N_2666);
nor U3486 (N_3486,N_2028,N_2224);
nor U3487 (N_3487,N_2268,N_2440);
xor U3488 (N_3488,N_2178,N_2250);
xnor U3489 (N_3489,N_2876,N_2777);
or U3490 (N_3490,N_2686,N_2628);
and U3491 (N_3491,N_2249,N_2999);
and U3492 (N_3492,N_2035,N_2424);
xor U3493 (N_3493,N_2780,N_2390);
and U3494 (N_3494,N_2079,N_2195);
xnor U3495 (N_3495,N_2097,N_2066);
or U3496 (N_3496,N_2069,N_2115);
xnor U3497 (N_3497,N_2792,N_2434);
nand U3498 (N_3498,N_2915,N_2611);
xor U3499 (N_3499,N_2897,N_2911);
nor U3500 (N_3500,N_2607,N_2970);
nand U3501 (N_3501,N_2339,N_2239);
and U3502 (N_3502,N_2808,N_2803);
nand U3503 (N_3503,N_2298,N_2064);
xor U3504 (N_3504,N_2143,N_2424);
nand U3505 (N_3505,N_2538,N_2257);
nand U3506 (N_3506,N_2163,N_2068);
or U3507 (N_3507,N_2298,N_2159);
or U3508 (N_3508,N_2468,N_2255);
nor U3509 (N_3509,N_2671,N_2537);
nor U3510 (N_3510,N_2335,N_2123);
or U3511 (N_3511,N_2226,N_2281);
nand U3512 (N_3512,N_2137,N_2056);
xor U3513 (N_3513,N_2551,N_2805);
nand U3514 (N_3514,N_2393,N_2992);
or U3515 (N_3515,N_2183,N_2909);
xor U3516 (N_3516,N_2697,N_2133);
or U3517 (N_3517,N_2096,N_2226);
or U3518 (N_3518,N_2927,N_2132);
and U3519 (N_3519,N_2404,N_2191);
xor U3520 (N_3520,N_2213,N_2581);
xnor U3521 (N_3521,N_2897,N_2248);
and U3522 (N_3522,N_2234,N_2837);
and U3523 (N_3523,N_2789,N_2997);
and U3524 (N_3524,N_2197,N_2717);
or U3525 (N_3525,N_2409,N_2980);
and U3526 (N_3526,N_2263,N_2563);
xor U3527 (N_3527,N_2602,N_2997);
nor U3528 (N_3528,N_2673,N_2799);
nor U3529 (N_3529,N_2039,N_2995);
and U3530 (N_3530,N_2927,N_2523);
xor U3531 (N_3531,N_2797,N_2698);
nand U3532 (N_3532,N_2128,N_2834);
nor U3533 (N_3533,N_2733,N_2101);
xnor U3534 (N_3534,N_2060,N_2837);
xor U3535 (N_3535,N_2903,N_2378);
nand U3536 (N_3536,N_2366,N_2772);
and U3537 (N_3537,N_2101,N_2184);
nand U3538 (N_3538,N_2271,N_2911);
nor U3539 (N_3539,N_2736,N_2225);
nand U3540 (N_3540,N_2060,N_2524);
nand U3541 (N_3541,N_2527,N_2906);
and U3542 (N_3542,N_2618,N_2143);
or U3543 (N_3543,N_2133,N_2210);
and U3544 (N_3544,N_2759,N_2268);
nor U3545 (N_3545,N_2237,N_2442);
and U3546 (N_3546,N_2096,N_2123);
and U3547 (N_3547,N_2113,N_2060);
and U3548 (N_3548,N_2902,N_2844);
xor U3549 (N_3549,N_2214,N_2853);
nand U3550 (N_3550,N_2070,N_2602);
and U3551 (N_3551,N_2199,N_2590);
nand U3552 (N_3552,N_2976,N_2572);
nor U3553 (N_3553,N_2577,N_2465);
or U3554 (N_3554,N_2063,N_2325);
nand U3555 (N_3555,N_2172,N_2361);
nand U3556 (N_3556,N_2035,N_2586);
and U3557 (N_3557,N_2258,N_2978);
nand U3558 (N_3558,N_2564,N_2639);
or U3559 (N_3559,N_2740,N_2022);
and U3560 (N_3560,N_2630,N_2981);
or U3561 (N_3561,N_2582,N_2559);
and U3562 (N_3562,N_2773,N_2823);
or U3563 (N_3563,N_2751,N_2006);
nor U3564 (N_3564,N_2941,N_2067);
and U3565 (N_3565,N_2399,N_2981);
nor U3566 (N_3566,N_2425,N_2289);
or U3567 (N_3567,N_2439,N_2872);
and U3568 (N_3568,N_2907,N_2945);
and U3569 (N_3569,N_2693,N_2130);
xor U3570 (N_3570,N_2274,N_2529);
nor U3571 (N_3571,N_2615,N_2934);
nand U3572 (N_3572,N_2582,N_2710);
or U3573 (N_3573,N_2903,N_2636);
xor U3574 (N_3574,N_2641,N_2568);
and U3575 (N_3575,N_2907,N_2393);
and U3576 (N_3576,N_2912,N_2833);
nand U3577 (N_3577,N_2840,N_2064);
and U3578 (N_3578,N_2358,N_2728);
nand U3579 (N_3579,N_2880,N_2371);
and U3580 (N_3580,N_2508,N_2107);
nor U3581 (N_3581,N_2709,N_2021);
or U3582 (N_3582,N_2530,N_2427);
nor U3583 (N_3583,N_2208,N_2065);
nand U3584 (N_3584,N_2120,N_2464);
or U3585 (N_3585,N_2603,N_2038);
or U3586 (N_3586,N_2494,N_2250);
nor U3587 (N_3587,N_2915,N_2157);
and U3588 (N_3588,N_2382,N_2283);
xor U3589 (N_3589,N_2273,N_2035);
nor U3590 (N_3590,N_2432,N_2980);
or U3591 (N_3591,N_2993,N_2925);
nand U3592 (N_3592,N_2626,N_2550);
nand U3593 (N_3593,N_2354,N_2718);
and U3594 (N_3594,N_2518,N_2940);
and U3595 (N_3595,N_2821,N_2013);
or U3596 (N_3596,N_2372,N_2155);
xor U3597 (N_3597,N_2615,N_2047);
or U3598 (N_3598,N_2936,N_2801);
nor U3599 (N_3599,N_2648,N_2761);
nor U3600 (N_3600,N_2242,N_2172);
and U3601 (N_3601,N_2233,N_2396);
nand U3602 (N_3602,N_2661,N_2890);
or U3603 (N_3603,N_2792,N_2402);
xnor U3604 (N_3604,N_2245,N_2050);
nand U3605 (N_3605,N_2002,N_2051);
or U3606 (N_3606,N_2052,N_2803);
nand U3607 (N_3607,N_2765,N_2680);
and U3608 (N_3608,N_2258,N_2917);
nand U3609 (N_3609,N_2316,N_2954);
nand U3610 (N_3610,N_2743,N_2764);
nand U3611 (N_3611,N_2299,N_2977);
xnor U3612 (N_3612,N_2370,N_2308);
or U3613 (N_3613,N_2166,N_2167);
or U3614 (N_3614,N_2423,N_2574);
nor U3615 (N_3615,N_2763,N_2368);
and U3616 (N_3616,N_2568,N_2985);
and U3617 (N_3617,N_2339,N_2496);
nor U3618 (N_3618,N_2712,N_2537);
xnor U3619 (N_3619,N_2341,N_2705);
or U3620 (N_3620,N_2852,N_2625);
nand U3621 (N_3621,N_2656,N_2308);
nand U3622 (N_3622,N_2832,N_2371);
or U3623 (N_3623,N_2472,N_2504);
and U3624 (N_3624,N_2034,N_2101);
xnor U3625 (N_3625,N_2260,N_2681);
nor U3626 (N_3626,N_2177,N_2815);
xnor U3627 (N_3627,N_2118,N_2942);
xor U3628 (N_3628,N_2221,N_2216);
nor U3629 (N_3629,N_2352,N_2533);
or U3630 (N_3630,N_2085,N_2994);
or U3631 (N_3631,N_2591,N_2767);
or U3632 (N_3632,N_2058,N_2095);
nand U3633 (N_3633,N_2981,N_2438);
or U3634 (N_3634,N_2627,N_2133);
and U3635 (N_3635,N_2649,N_2446);
or U3636 (N_3636,N_2782,N_2323);
and U3637 (N_3637,N_2789,N_2479);
nor U3638 (N_3638,N_2585,N_2287);
nand U3639 (N_3639,N_2545,N_2409);
xnor U3640 (N_3640,N_2183,N_2602);
nor U3641 (N_3641,N_2848,N_2736);
or U3642 (N_3642,N_2491,N_2988);
or U3643 (N_3643,N_2273,N_2362);
and U3644 (N_3644,N_2321,N_2753);
or U3645 (N_3645,N_2430,N_2029);
nor U3646 (N_3646,N_2371,N_2287);
or U3647 (N_3647,N_2698,N_2062);
nand U3648 (N_3648,N_2502,N_2317);
or U3649 (N_3649,N_2171,N_2556);
xnor U3650 (N_3650,N_2834,N_2879);
and U3651 (N_3651,N_2307,N_2762);
or U3652 (N_3652,N_2205,N_2386);
nand U3653 (N_3653,N_2346,N_2970);
or U3654 (N_3654,N_2538,N_2184);
nand U3655 (N_3655,N_2475,N_2086);
nor U3656 (N_3656,N_2293,N_2716);
nor U3657 (N_3657,N_2397,N_2180);
nand U3658 (N_3658,N_2773,N_2666);
nor U3659 (N_3659,N_2476,N_2618);
nand U3660 (N_3660,N_2212,N_2539);
and U3661 (N_3661,N_2492,N_2629);
and U3662 (N_3662,N_2033,N_2930);
or U3663 (N_3663,N_2836,N_2249);
xor U3664 (N_3664,N_2408,N_2897);
or U3665 (N_3665,N_2965,N_2420);
nor U3666 (N_3666,N_2823,N_2992);
nand U3667 (N_3667,N_2847,N_2065);
nand U3668 (N_3668,N_2285,N_2376);
nor U3669 (N_3669,N_2497,N_2918);
nor U3670 (N_3670,N_2108,N_2386);
or U3671 (N_3671,N_2425,N_2579);
nand U3672 (N_3672,N_2722,N_2774);
or U3673 (N_3673,N_2165,N_2118);
and U3674 (N_3674,N_2908,N_2976);
and U3675 (N_3675,N_2476,N_2930);
nand U3676 (N_3676,N_2863,N_2675);
nand U3677 (N_3677,N_2880,N_2698);
and U3678 (N_3678,N_2770,N_2363);
and U3679 (N_3679,N_2181,N_2706);
nand U3680 (N_3680,N_2071,N_2060);
xnor U3681 (N_3681,N_2879,N_2326);
nand U3682 (N_3682,N_2742,N_2307);
xnor U3683 (N_3683,N_2425,N_2162);
nand U3684 (N_3684,N_2792,N_2290);
and U3685 (N_3685,N_2591,N_2707);
nand U3686 (N_3686,N_2395,N_2401);
nor U3687 (N_3687,N_2084,N_2666);
nand U3688 (N_3688,N_2629,N_2659);
and U3689 (N_3689,N_2452,N_2294);
nand U3690 (N_3690,N_2305,N_2967);
or U3691 (N_3691,N_2179,N_2722);
and U3692 (N_3692,N_2393,N_2083);
or U3693 (N_3693,N_2178,N_2595);
or U3694 (N_3694,N_2501,N_2781);
nand U3695 (N_3695,N_2284,N_2235);
xor U3696 (N_3696,N_2986,N_2414);
nor U3697 (N_3697,N_2716,N_2354);
and U3698 (N_3698,N_2565,N_2468);
nor U3699 (N_3699,N_2845,N_2600);
nor U3700 (N_3700,N_2807,N_2558);
nor U3701 (N_3701,N_2076,N_2600);
or U3702 (N_3702,N_2678,N_2415);
or U3703 (N_3703,N_2044,N_2943);
nor U3704 (N_3704,N_2035,N_2184);
and U3705 (N_3705,N_2019,N_2950);
and U3706 (N_3706,N_2846,N_2120);
and U3707 (N_3707,N_2949,N_2813);
nand U3708 (N_3708,N_2963,N_2151);
and U3709 (N_3709,N_2818,N_2362);
or U3710 (N_3710,N_2925,N_2206);
nor U3711 (N_3711,N_2292,N_2708);
and U3712 (N_3712,N_2762,N_2866);
or U3713 (N_3713,N_2832,N_2485);
or U3714 (N_3714,N_2308,N_2116);
and U3715 (N_3715,N_2736,N_2229);
nor U3716 (N_3716,N_2193,N_2738);
or U3717 (N_3717,N_2325,N_2990);
nand U3718 (N_3718,N_2309,N_2716);
nand U3719 (N_3719,N_2926,N_2488);
nor U3720 (N_3720,N_2833,N_2704);
and U3721 (N_3721,N_2547,N_2282);
xor U3722 (N_3722,N_2086,N_2148);
xor U3723 (N_3723,N_2401,N_2854);
and U3724 (N_3724,N_2741,N_2170);
and U3725 (N_3725,N_2769,N_2895);
xnor U3726 (N_3726,N_2353,N_2369);
or U3727 (N_3727,N_2802,N_2990);
nand U3728 (N_3728,N_2969,N_2117);
nand U3729 (N_3729,N_2287,N_2895);
or U3730 (N_3730,N_2808,N_2685);
or U3731 (N_3731,N_2728,N_2360);
nor U3732 (N_3732,N_2317,N_2163);
nor U3733 (N_3733,N_2282,N_2724);
and U3734 (N_3734,N_2706,N_2226);
nand U3735 (N_3735,N_2857,N_2340);
or U3736 (N_3736,N_2971,N_2646);
and U3737 (N_3737,N_2301,N_2252);
or U3738 (N_3738,N_2349,N_2543);
or U3739 (N_3739,N_2629,N_2979);
nor U3740 (N_3740,N_2133,N_2560);
nor U3741 (N_3741,N_2225,N_2508);
or U3742 (N_3742,N_2149,N_2277);
nor U3743 (N_3743,N_2158,N_2496);
nor U3744 (N_3744,N_2904,N_2934);
or U3745 (N_3745,N_2284,N_2918);
nand U3746 (N_3746,N_2241,N_2516);
and U3747 (N_3747,N_2875,N_2012);
or U3748 (N_3748,N_2528,N_2981);
nor U3749 (N_3749,N_2723,N_2123);
nand U3750 (N_3750,N_2274,N_2699);
or U3751 (N_3751,N_2294,N_2352);
nand U3752 (N_3752,N_2881,N_2755);
and U3753 (N_3753,N_2702,N_2038);
nand U3754 (N_3754,N_2599,N_2263);
and U3755 (N_3755,N_2715,N_2082);
xnor U3756 (N_3756,N_2013,N_2187);
and U3757 (N_3757,N_2252,N_2547);
and U3758 (N_3758,N_2290,N_2796);
or U3759 (N_3759,N_2595,N_2660);
nor U3760 (N_3760,N_2064,N_2059);
and U3761 (N_3761,N_2339,N_2616);
and U3762 (N_3762,N_2696,N_2529);
xor U3763 (N_3763,N_2529,N_2336);
nor U3764 (N_3764,N_2365,N_2324);
or U3765 (N_3765,N_2356,N_2274);
nand U3766 (N_3766,N_2662,N_2520);
and U3767 (N_3767,N_2250,N_2169);
nand U3768 (N_3768,N_2043,N_2284);
nor U3769 (N_3769,N_2012,N_2028);
nor U3770 (N_3770,N_2592,N_2191);
or U3771 (N_3771,N_2913,N_2059);
nand U3772 (N_3772,N_2270,N_2714);
or U3773 (N_3773,N_2966,N_2246);
nand U3774 (N_3774,N_2702,N_2658);
nor U3775 (N_3775,N_2471,N_2138);
and U3776 (N_3776,N_2641,N_2507);
and U3777 (N_3777,N_2671,N_2993);
and U3778 (N_3778,N_2032,N_2400);
nor U3779 (N_3779,N_2591,N_2481);
nor U3780 (N_3780,N_2928,N_2542);
and U3781 (N_3781,N_2384,N_2541);
nor U3782 (N_3782,N_2924,N_2400);
nand U3783 (N_3783,N_2670,N_2238);
and U3784 (N_3784,N_2691,N_2812);
and U3785 (N_3785,N_2958,N_2678);
nor U3786 (N_3786,N_2059,N_2136);
nand U3787 (N_3787,N_2079,N_2896);
or U3788 (N_3788,N_2983,N_2207);
xor U3789 (N_3789,N_2944,N_2278);
and U3790 (N_3790,N_2720,N_2727);
xor U3791 (N_3791,N_2117,N_2450);
nand U3792 (N_3792,N_2804,N_2319);
nand U3793 (N_3793,N_2002,N_2134);
xor U3794 (N_3794,N_2901,N_2250);
and U3795 (N_3795,N_2295,N_2223);
nor U3796 (N_3796,N_2618,N_2557);
nor U3797 (N_3797,N_2327,N_2318);
nor U3798 (N_3798,N_2575,N_2426);
nand U3799 (N_3799,N_2371,N_2353);
or U3800 (N_3800,N_2714,N_2417);
and U3801 (N_3801,N_2278,N_2614);
and U3802 (N_3802,N_2870,N_2946);
xnor U3803 (N_3803,N_2062,N_2935);
nor U3804 (N_3804,N_2536,N_2562);
and U3805 (N_3805,N_2406,N_2684);
or U3806 (N_3806,N_2578,N_2119);
nand U3807 (N_3807,N_2174,N_2533);
or U3808 (N_3808,N_2054,N_2134);
nor U3809 (N_3809,N_2748,N_2812);
and U3810 (N_3810,N_2762,N_2361);
nand U3811 (N_3811,N_2416,N_2302);
nor U3812 (N_3812,N_2286,N_2631);
nand U3813 (N_3813,N_2604,N_2058);
nor U3814 (N_3814,N_2380,N_2818);
xnor U3815 (N_3815,N_2360,N_2779);
nand U3816 (N_3816,N_2536,N_2135);
nor U3817 (N_3817,N_2092,N_2799);
nand U3818 (N_3818,N_2895,N_2693);
nor U3819 (N_3819,N_2535,N_2993);
or U3820 (N_3820,N_2033,N_2325);
nand U3821 (N_3821,N_2898,N_2414);
or U3822 (N_3822,N_2481,N_2889);
and U3823 (N_3823,N_2385,N_2089);
and U3824 (N_3824,N_2113,N_2024);
nand U3825 (N_3825,N_2632,N_2123);
and U3826 (N_3826,N_2096,N_2337);
nand U3827 (N_3827,N_2247,N_2045);
nand U3828 (N_3828,N_2787,N_2492);
or U3829 (N_3829,N_2941,N_2001);
xor U3830 (N_3830,N_2828,N_2023);
or U3831 (N_3831,N_2169,N_2304);
and U3832 (N_3832,N_2906,N_2163);
or U3833 (N_3833,N_2803,N_2592);
and U3834 (N_3834,N_2975,N_2514);
and U3835 (N_3835,N_2700,N_2579);
or U3836 (N_3836,N_2139,N_2673);
nor U3837 (N_3837,N_2464,N_2546);
nor U3838 (N_3838,N_2666,N_2728);
and U3839 (N_3839,N_2721,N_2652);
nand U3840 (N_3840,N_2781,N_2283);
or U3841 (N_3841,N_2218,N_2878);
nor U3842 (N_3842,N_2630,N_2958);
nand U3843 (N_3843,N_2199,N_2085);
and U3844 (N_3844,N_2995,N_2415);
nor U3845 (N_3845,N_2235,N_2325);
and U3846 (N_3846,N_2837,N_2681);
nand U3847 (N_3847,N_2468,N_2348);
and U3848 (N_3848,N_2878,N_2776);
or U3849 (N_3849,N_2037,N_2670);
and U3850 (N_3850,N_2472,N_2633);
nor U3851 (N_3851,N_2374,N_2880);
and U3852 (N_3852,N_2406,N_2206);
nor U3853 (N_3853,N_2109,N_2600);
and U3854 (N_3854,N_2387,N_2684);
or U3855 (N_3855,N_2164,N_2451);
nor U3856 (N_3856,N_2618,N_2580);
or U3857 (N_3857,N_2083,N_2487);
and U3858 (N_3858,N_2519,N_2595);
and U3859 (N_3859,N_2408,N_2475);
nand U3860 (N_3860,N_2724,N_2832);
xor U3861 (N_3861,N_2991,N_2898);
nor U3862 (N_3862,N_2516,N_2896);
nand U3863 (N_3863,N_2369,N_2553);
or U3864 (N_3864,N_2140,N_2733);
nand U3865 (N_3865,N_2869,N_2187);
and U3866 (N_3866,N_2886,N_2332);
and U3867 (N_3867,N_2976,N_2936);
or U3868 (N_3868,N_2948,N_2380);
and U3869 (N_3869,N_2225,N_2397);
or U3870 (N_3870,N_2415,N_2226);
nor U3871 (N_3871,N_2671,N_2454);
xor U3872 (N_3872,N_2231,N_2347);
and U3873 (N_3873,N_2589,N_2218);
nor U3874 (N_3874,N_2824,N_2893);
xor U3875 (N_3875,N_2434,N_2369);
or U3876 (N_3876,N_2120,N_2342);
nand U3877 (N_3877,N_2471,N_2316);
and U3878 (N_3878,N_2056,N_2029);
or U3879 (N_3879,N_2034,N_2403);
and U3880 (N_3880,N_2004,N_2951);
nor U3881 (N_3881,N_2328,N_2347);
nand U3882 (N_3882,N_2075,N_2835);
or U3883 (N_3883,N_2784,N_2487);
or U3884 (N_3884,N_2100,N_2319);
nand U3885 (N_3885,N_2237,N_2937);
nor U3886 (N_3886,N_2593,N_2396);
and U3887 (N_3887,N_2906,N_2842);
or U3888 (N_3888,N_2247,N_2770);
or U3889 (N_3889,N_2763,N_2292);
or U3890 (N_3890,N_2098,N_2642);
nand U3891 (N_3891,N_2686,N_2960);
xnor U3892 (N_3892,N_2104,N_2984);
xor U3893 (N_3893,N_2195,N_2902);
and U3894 (N_3894,N_2945,N_2757);
or U3895 (N_3895,N_2496,N_2820);
nor U3896 (N_3896,N_2581,N_2007);
nand U3897 (N_3897,N_2088,N_2583);
xnor U3898 (N_3898,N_2039,N_2735);
nor U3899 (N_3899,N_2184,N_2804);
nand U3900 (N_3900,N_2066,N_2497);
nor U3901 (N_3901,N_2706,N_2729);
or U3902 (N_3902,N_2560,N_2748);
or U3903 (N_3903,N_2888,N_2205);
nand U3904 (N_3904,N_2188,N_2530);
nand U3905 (N_3905,N_2510,N_2453);
nor U3906 (N_3906,N_2845,N_2612);
and U3907 (N_3907,N_2306,N_2214);
nor U3908 (N_3908,N_2753,N_2165);
and U3909 (N_3909,N_2032,N_2430);
nor U3910 (N_3910,N_2659,N_2884);
nor U3911 (N_3911,N_2072,N_2698);
or U3912 (N_3912,N_2908,N_2769);
nor U3913 (N_3913,N_2012,N_2380);
nor U3914 (N_3914,N_2062,N_2554);
or U3915 (N_3915,N_2766,N_2208);
nor U3916 (N_3916,N_2633,N_2997);
nand U3917 (N_3917,N_2157,N_2736);
and U3918 (N_3918,N_2564,N_2413);
or U3919 (N_3919,N_2834,N_2252);
and U3920 (N_3920,N_2846,N_2091);
nand U3921 (N_3921,N_2804,N_2886);
or U3922 (N_3922,N_2196,N_2165);
and U3923 (N_3923,N_2460,N_2175);
and U3924 (N_3924,N_2690,N_2549);
nor U3925 (N_3925,N_2403,N_2715);
and U3926 (N_3926,N_2791,N_2641);
xor U3927 (N_3927,N_2988,N_2946);
and U3928 (N_3928,N_2027,N_2734);
and U3929 (N_3929,N_2814,N_2671);
nand U3930 (N_3930,N_2651,N_2948);
nor U3931 (N_3931,N_2257,N_2073);
or U3932 (N_3932,N_2054,N_2498);
or U3933 (N_3933,N_2932,N_2523);
nand U3934 (N_3934,N_2873,N_2553);
or U3935 (N_3935,N_2424,N_2699);
xnor U3936 (N_3936,N_2621,N_2879);
or U3937 (N_3937,N_2837,N_2848);
and U3938 (N_3938,N_2694,N_2656);
xnor U3939 (N_3939,N_2158,N_2430);
and U3940 (N_3940,N_2342,N_2500);
and U3941 (N_3941,N_2366,N_2659);
and U3942 (N_3942,N_2975,N_2290);
nand U3943 (N_3943,N_2182,N_2197);
and U3944 (N_3944,N_2791,N_2274);
and U3945 (N_3945,N_2751,N_2728);
or U3946 (N_3946,N_2419,N_2854);
nor U3947 (N_3947,N_2438,N_2816);
nor U3948 (N_3948,N_2419,N_2773);
nand U3949 (N_3949,N_2140,N_2503);
or U3950 (N_3950,N_2300,N_2136);
nor U3951 (N_3951,N_2907,N_2089);
and U3952 (N_3952,N_2151,N_2612);
nand U3953 (N_3953,N_2839,N_2619);
and U3954 (N_3954,N_2661,N_2925);
xnor U3955 (N_3955,N_2274,N_2185);
and U3956 (N_3956,N_2919,N_2759);
and U3957 (N_3957,N_2537,N_2896);
nand U3958 (N_3958,N_2351,N_2914);
nand U3959 (N_3959,N_2148,N_2111);
nand U3960 (N_3960,N_2952,N_2608);
nand U3961 (N_3961,N_2708,N_2046);
nand U3962 (N_3962,N_2863,N_2457);
xnor U3963 (N_3963,N_2980,N_2411);
nand U3964 (N_3964,N_2573,N_2699);
nor U3965 (N_3965,N_2033,N_2659);
or U3966 (N_3966,N_2663,N_2484);
and U3967 (N_3967,N_2783,N_2141);
nand U3968 (N_3968,N_2007,N_2735);
or U3969 (N_3969,N_2156,N_2479);
nor U3970 (N_3970,N_2139,N_2645);
or U3971 (N_3971,N_2970,N_2338);
and U3972 (N_3972,N_2250,N_2609);
or U3973 (N_3973,N_2886,N_2359);
or U3974 (N_3974,N_2673,N_2028);
nand U3975 (N_3975,N_2631,N_2330);
nor U3976 (N_3976,N_2977,N_2073);
or U3977 (N_3977,N_2170,N_2757);
nor U3978 (N_3978,N_2284,N_2372);
or U3979 (N_3979,N_2053,N_2256);
and U3980 (N_3980,N_2417,N_2616);
and U3981 (N_3981,N_2808,N_2331);
nor U3982 (N_3982,N_2443,N_2756);
or U3983 (N_3983,N_2411,N_2213);
xor U3984 (N_3984,N_2549,N_2044);
or U3985 (N_3985,N_2732,N_2253);
nor U3986 (N_3986,N_2185,N_2620);
nand U3987 (N_3987,N_2387,N_2674);
or U3988 (N_3988,N_2348,N_2284);
and U3989 (N_3989,N_2305,N_2483);
nand U3990 (N_3990,N_2056,N_2552);
and U3991 (N_3991,N_2713,N_2114);
nand U3992 (N_3992,N_2792,N_2135);
or U3993 (N_3993,N_2376,N_2972);
nand U3994 (N_3994,N_2820,N_2690);
nand U3995 (N_3995,N_2934,N_2104);
xor U3996 (N_3996,N_2492,N_2894);
and U3997 (N_3997,N_2202,N_2459);
nor U3998 (N_3998,N_2516,N_2583);
xor U3999 (N_3999,N_2895,N_2108);
or U4000 (N_4000,N_3357,N_3324);
xnor U4001 (N_4001,N_3215,N_3256);
nand U4002 (N_4002,N_3009,N_3580);
nand U4003 (N_4003,N_3113,N_3822);
and U4004 (N_4004,N_3348,N_3501);
or U4005 (N_4005,N_3549,N_3763);
and U4006 (N_4006,N_3230,N_3940);
xnor U4007 (N_4007,N_3091,N_3169);
nor U4008 (N_4008,N_3359,N_3967);
nand U4009 (N_4009,N_3863,N_3366);
nand U4010 (N_4010,N_3685,N_3221);
nor U4011 (N_4011,N_3669,N_3275);
or U4012 (N_4012,N_3400,N_3854);
nor U4013 (N_4013,N_3878,N_3417);
or U4014 (N_4014,N_3869,N_3175);
nor U4015 (N_4015,N_3646,N_3194);
nand U4016 (N_4016,N_3054,N_3949);
nand U4017 (N_4017,N_3942,N_3701);
or U4018 (N_4018,N_3453,N_3068);
nand U4019 (N_4019,N_3190,N_3441);
and U4020 (N_4020,N_3868,N_3493);
and U4021 (N_4021,N_3595,N_3153);
nor U4022 (N_4022,N_3399,N_3533);
xnor U4023 (N_4023,N_3197,N_3810);
xnor U4024 (N_4024,N_3142,N_3261);
and U4025 (N_4025,N_3048,N_3136);
nand U4026 (N_4026,N_3691,N_3771);
nand U4027 (N_4027,N_3069,N_3220);
xnor U4028 (N_4028,N_3515,N_3895);
or U4029 (N_4029,N_3788,N_3758);
nor U4030 (N_4030,N_3634,N_3893);
nor U4031 (N_4031,N_3316,N_3222);
xnor U4032 (N_4032,N_3250,N_3428);
nor U4033 (N_4033,N_3335,N_3704);
nor U4034 (N_4034,N_3997,N_3527);
xnor U4035 (N_4035,N_3747,N_3782);
nor U4036 (N_4036,N_3905,N_3717);
and U4037 (N_4037,N_3920,N_3645);
xnor U4038 (N_4038,N_3539,N_3017);
nor U4039 (N_4039,N_3235,N_3579);
nand U4040 (N_4040,N_3584,N_3554);
and U4041 (N_4041,N_3706,N_3476);
nand U4042 (N_4042,N_3187,N_3380);
or U4043 (N_4043,N_3756,N_3360);
nor U4044 (N_4044,N_3877,N_3793);
nand U4045 (N_4045,N_3448,N_3563);
nand U4046 (N_4046,N_3383,N_3847);
xor U4047 (N_4047,N_3770,N_3519);
nand U4048 (N_4048,N_3486,N_3376);
and U4049 (N_4049,N_3974,N_3491);
or U4050 (N_4050,N_3059,N_3223);
nor U4051 (N_4051,N_3299,N_3056);
and U4052 (N_4052,N_3978,N_3991);
or U4053 (N_4053,N_3729,N_3590);
nand U4054 (N_4054,N_3842,N_3667);
nand U4055 (N_4055,N_3690,N_3640);
nor U4056 (N_4056,N_3405,N_3787);
and U4057 (N_4057,N_3814,N_3266);
nand U4058 (N_4058,N_3638,N_3098);
nand U4059 (N_4059,N_3733,N_3676);
or U4060 (N_4060,N_3444,N_3093);
nor U4061 (N_4061,N_3523,N_3530);
xnor U4062 (N_4062,N_3970,N_3532);
nand U4063 (N_4063,N_3425,N_3154);
or U4064 (N_4064,N_3671,N_3838);
or U4065 (N_4065,N_3976,N_3458);
nand U4066 (N_4066,N_3742,N_3705);
or U4067 (N_4067,N_3981,N_3962);
xor U4068 (N_4068,N_3648,N_3343);
and U4069 (N_4069,N_3713,N_3754);
and U4070 (N_4070,N_3079,N_3118);
and U4071 (N_4071,N_3484,N_3662);
nor U4072 (N_4072,N_3427,N_3435);
or U4073 (N_4073,N_3172,N_3278);
nor U4074 (N_4074,N_3524,N_3636);
and U4075 (N_4075,N_3833,N_3642);
xnor U4076 (N_4076,N_3625,N_3020);
or U4077 (N_4077,N_3109,N_3857);
and U4078 (N_4078,N_3319,N_3851);
or U4079 (N_4079,N_3916,N_3389);
nor U4080 (N_4080,N_3065,N_3332);
or U4081 (N_4081,N_3908,N_3875);
nor U4082 (N_4082,N_3798,N_3687);
nor U4083 (N_4083,N_3150,N_3252);
nand U4084 (N_4084,N_3621,N_3070);
nor U4085 (N_4085,N_3693,N_3200);
and U4086 (N_4086,N_3748,N_3732);
nand U4087 (N_4087,N_3209,N_3945);
xor U4088 (N_4088,N_3585,N_3609);
nand U4089 (N_4089,N_3024,N_3503);
nand U4090 (N_4090,N_3921,N_3925);
and U4091 (N_4091,N_3617,N_3802);
nor U4092 (N_4092,N_3510,N_3689);
and U4093 (N_4093,N_3149,N_3882);
nand U4094 (N_4094,N_3795,N_3816);
nand U4095 (N_4095,N_3482,N_3078);
or U4096 (N_4096,N_3635,N_3651);
nand U4097 (N_4097,N_3047,N_3544);
nor U4098 (N_4098,N_3591,N_3198);
nor U4099 (N_4099,N_3783,N_3211);
xnor U4100 (N_4100,N_3233,N_3718);
and U4101 (N_4101,N_3144,N_3112);
and U4102 (N_4102,N_3917,N_3295);
nor U4103 (N_4103,N_3856,N_3883);
nand U4104 (N_4104,N_3298,N_3182);
or U4105 (N_4105,N_3821,N_3774);
or U4106 (N_4106,N_3650,N_3099);
xnor U4107 (N_4107,N_3294,N_3464);
and U4108 (N_4108,N_3518,N_3156);
or U4109 (N_4109,N_3002,N_3203);
nand U4110 (N_4110,N_3269,N_3352);
nand U4111 (N_4111,N_3206,N_3664);
nor U4112 (N_4112,N_3291,N_3864);
nand U4113 (N_4113,N_3305,N_3710);
or U4114 (N_4114,N_3353,N_3499);
and U4115 (N_4115,N_3089,N_3548);
xnor U4116 (N_4116,N_3328,N_3557);
nand U4117 (N_4117,N_3236,N_3268);
or U4118 (N_4118,N_3722,N_3263);
xor U4119 (N_4119,N_3684,N_3589);
nor U4120 (N_4120,N_3440,N_3108);
or U4121 (N_4121,N_3026,N_3016);
and U4122 (N_4122,N_3892,N_3364);
and U4123 (N_4123,N_3556,N_3979);
or U4124 (N_4124,N_3547,N_3057);
xor U4125 (N_4125,N_3932,N_3536);
nor U4126 (N_4126,N_3654,N_3596);
xor U4127 (N_4127,N_3682,N_3008);
nor U4128 (N_4128,N_3429,N_3937);
or U4129 (N_4129,N_3067,N_3210);
nand U4130 (N_4130,N_3204,N_3337);
nand U4131 (N_4131,N_3034,N_3260);
xor U4132 (N_4132,N_3046,N_3082);
or U4133 (N_4133,N_3568,N_3708);
nor U4134 (N_4134,N_3987,N_3051);
xnor U4135 (N_4135,N_3692,N_3426);
nand U4136 (N_4136,N_3373,N_3117);
or U4137 (N_4137,N_3846,N_3829);
nor U4138 (N_4138,N_3355,N_3290);
or U4139 (N_4139,N_3124,N_3422);
or U4140 (N_4140,N_3354,N_3721);
nand U4141 (N_4141,N_3021,N_3575);
nor U4142 (N_4142,N_3063,N_3028);
and U4143 (N_4143,N_3811,N_3943);
and U4144 (N_4144,N_3660,N_3672);
and U4145 (N_4145,N_3673,N_3891);
nor U4146 (N_4146,N_3623,N_3968);
xnor U4147 (N_4147,N_3189,N_3447);
nand U4148 (N_4148,N_3132,N_3870);
nor U4149 (N_4149,N_3966,N_3151);
or U4150 (N_4150,N_3762,N_3504);
xor U4151 (N_4151,N_3094,N_3349);
nand U4152 (N_4152,N_3367,N_3781);
nor U4153 (N_4153,N_3066,N_3724);
nor U4154 (N_4154,N_3728,N_3488);
nand U4155 (N_4155,N_3449,N_3903);
xor U4156 (N_4156,N_3351,N_3871);
and U4157 (N_4157,N_3277,N_3387);
and U4158 (N_4158,N_3508,N_3471);
nor U4159 (N_4159,N_3247,N_3894);
xor U4160 (N_4160,N_3304,N_3392);
and U4161 (N_4161,N_3700,N_3941);
and U4162 (N_4162,N_3490,N_3831);
nor U4163 (N_4163,N_3889,N_3919);
or U4164 (N_4164,N_3924,N_3786);
nor U4165 (N_4165,N_3385,N_3765);
xnor U4166 (N_4166,N_3329,N_3844);
and U4167 (N_4167,N_3961,N_3887);
nor U4168 (N_4168,N_3027,N_3282);
nor U4169 (N_4169,N_3639,N_3271);
nand U4170 (N_4170,N_3657,N_3307);
or U4171 (N_4171,N_3752,N_3288);
nor U4172 (N_4172,N_3993,N_3292);
xor U4173 (N_4173,N_3293,N_3165);
and U4174 (N_4174,N_3181,N_3627);
nor U4175 (N_4175,N_3995,N_3217);
nor U4176 (N_4176,N_3365,N_3064);
and U4177 (N_4177,N_3287,N_3450);
nand U4178 (N_4178,N_3564,N_3884);
or U4179 (N_4179,N_3661,N_3817);
and U4180 (N_4180,N_3577,N_3773);
nand U4181 (N_4181,N_3622,N_3982);
nand U4182 (N_4182,N_3567,N_3980);
nand U4183 (N_4183,N_3478,N_3192);
xnor U4184 (N_4184,N_3445,N_3258);
and U4185 (N_4185,N_3439,N_3601);
nand U4186 (N_4186,N_3990,N_3741);
nor U4187 (N_4187,N_3302,N_3558);
or U4188 (N_4188,N_3096,N_3725);
and U4189 (N_4189,N_3423,N_3963);
and U4190 (N_4190,N_3517,N_3163);
and U4191 (N_4191,N_3614,N_3456);
nor U4192 (N_4192,N_3679,N_3767);
and U4193 (N_4193,N_3309,N_3242);
nand U4194 (N_4194,N_3576,N_3018);
nor U4195 (N_4195,N_3106,N_3931);
and U4196 (N_4196,N_3137,N_3855);
nand U4197 (N_4197,N_3415,N_3935);
and U4198 (N_4198,N_3393,N_3301);
nand U4199 (N_4199,N_3600,N_3371);
nand U4200 (N_4200,N_3837,N_3485);
xor U4201 (N_4201,N_3396,N_3280);
nand U4202 (N_4202,N_3356,N_3226);
nor U4203 (N_4203,N_3133,N_3985);
nand U4204 (N_4204,N_3193,N_3947);
nor U4205 (N_4205,N_3246,N_3284);
or U4206 (N_4206,N_3414,N_3633);
nand U4207 (N_4207,N_3755,N_3602);
xor U4208 (N_4208,N_3326,N_3031);
nor U4209 (N_4209,N_3898,N_3500);
nand U4210 (N_4210,N_3806,N_3241);
nand U4211 (N_4211,N_3964,N_3224);
nand U4212 (N_4212,N_3570,N_3404);
xnor U4213 (N_4213,N_3668,N_3043);
or U4214 (N_4214,N_3946,N_3922);
or U4215 (N_4215,N_3680,N_3746);
nor U4216 (N_4216,N_3597,N_3134);
nand U4217 (N_4217,N_3587,N_3088);
and U4218 (N_4218,N_3726,N_3419);
and U4219 (N_4219,N_3513,N_3442);
nor U4220 (N_4220,N_3338,N_3716);
nand U4221 (N_4221,N_3528,N_3095);
nand U4222 (N_4222,N_3703,N_3757);
and U4223 (N_4223,N_3331,N_3073);
nand U4224 (N_4224,N_3053,N_3382);
nand U4225 (N_4225,N_3583,N_3216);
nand U4226 (N_4226,N_3044,N_3205);
and U4227 (N_4227,N_3092,N_3911);
nor U4228 (N_4228,N_3372,N_3255);
and U4229 (N_4229,N_3731,N_3801);
and U4230 (N_4230,N_3267,N_3804);
nand U4231 (N_4231,N_3835,N_3511);
or U4232 (N_4232,N_3123,N_3121);
nor U4233 (N_4233,N_3229,N_3828);
nor U4234 (N_4234,N_3674,N_3011);
nor U4235 (N_4235,N_3466,N_3861);
and U4236 (N_4236,N_3115,N_3789);
or U4237 (N_4237,N_3727,N_3202);
xnor U4238 (N_4238,N_3735,N_3397);
nand U4239 (N_4239,N_3753,N_3760);
or U4240 (N_4240,N_3670,N_3412);
nor U4241 (N_4241,N_3166,N_3714);
nor U4242 (N_4242,N_3652,N_3446);
nand U4243 (N_4243,N_3346,N_3629);
nand U4244 (N_4244,N_3232,N_3249);
xor U4245 (N_4245,N_3688,N_3873);
nand U4246 (N_4246,N_3314,N_3418);
nand U4247 (N_4247,N_3483,N_3105);
and U4248 (N_4248,N_3167,N_3715);
and U4249 (N_4249,N_3384,N_3948);
and U4250 (N_4250,N_3698,N_3998);
and U4251 (N_4251,N_3743,N_3084);
nor U4252 (N_4252,N_3100,N_3984);
nand U4253 (N_4253,N_3666,N_3038);
and U4254 (N_4254,N_3929,N_3540);
or U4255 (N_4255,N_3406,N_3431);
and U4256 (N_4256,N_3253,N_3474);
nor U4257 (N_4257,N_3712,N_3345);
xor U4258 (N_4258,N_3928,N_3101);
or U4259 (N_4259,N_3543,N_3644);
nand U4260 (N_4260,N_3286,N_3045);
nand U4261 (N_4261,N_3516,N_3325);
nor U4262 (N_4262,N_3296,N_3107);
nand U4263 (N_4263,N_3604,N_3323);
nor U4264 (N_4264,N_3228,N_3308);
or U4265 (N_4265,N_3174,N_3522);
nor U4266 (N_4266,N_3244,N_3749);
nor U4267 (N_4267,N_3000,N_3049);
and U4268 (N_4268,N_3632,N_3561);
nor U4269 (N_4269,N_3014,N_3283);
and U4270 (N_4270,N_3463,N_3058);
or U4271 (N_4271,N_3465,N_3157);
and U4272 (N_4272,N_3502,N_3853);
nor U4273 (N_4273,N_3090,N_3512);
nand U4274 (N_4274,N_3487,N_3766);
and U4275 (N_4275,N_3850,N_3347);
or U4276 (N_4276,N_3039,N_3784);
nor U4277 (N_4277,N_3608,N_3610);
nand U4278 (N_4278,N_3312,N_3184);
and U4279 (N_4279,N_3907,N_3083);
or U4280 (N_4280,N_3158,N_3938);
nor U4281 (N_4281,N_3697,N_3819);
or U4282 (N_4282,N_3265,N_3479);
xnor U4283 (N_4283,N_3033,N_3339);
nand U4284 (N_4284,N_3103,N_3778);
nand U4285 (N_4285,N_3129,N_3824);
nand U4286 (N_4286,N_3649,N_3188);
and U4287 (N_4287,N_3720,N_3888);
or U4288 (N_4288,N_3497,N_3436);
nor U4289 (N_4289,N_3912,N_3832);
nor U4290 (N_4290,N_3251,N_3906);
or U4291 (N_4291,N_3035,N_3665);
nand U4292 (N_4292,N_3128,N_3245);
nand U4293 (N_4293,N_3276,N_3433);
nand U4294 (N_4294,N_3398,N_3734);
nor U4295 (N_4295,N_3272,N_3469);
or U4296 (N_4296,N_3183,N_3185);
xnor U4297 (N_4297,N_3022,N_3553);
and U4298 (N_4298,N_3195,N_3358);
or U4299 (N_4299,N_3139,N_3986);
or U4300 (N_4300,N_3212,N_3826);
and U4301 (N_4301,N_3881,N_3102);
and U4302 (N_4302,N_3201,N_3334);
nand U4303 (N_4303,N_3135,N_3333);
nor U4304 (N_4304,N_3240,N_3848);
xnor U4305 (N_4305,N_3876,N_3213);
nor U4306 (N_4306,N_3159,N_3840);
nand U4307 (N_4307,N_3506,N_3274);
xnor U4308 (N_4308,N_3815,N_3413);
nor U4309 (N_4309,N_3297,N_3694);
or U4310 (N_4310,N_3866,N_3707);
or U4311 (N_4311,N_3030,N_3231);
nand U4312 (N_4312,N_3958,N_3173);
nor U4313 (N_4313,N_3807,N_3001);
nand U4314 (N_4314,N_3475,N_3569);
or U4315 (N_4315,N_3141,N_3592);
and U4316 (N_4316,N_3775,N_3960);
nor U4317 (N_4317,N_3927,N_3534);
and U4318 (N_4318,N_3546,N_3790);
or U4319 (N_4319,N_3900,N_3571);
nor U4320 (N_4320,N_3408,N_3588);
and U4321 (N_4321,N_3492,N_3969);
or U4322 (N_4322,N_3125,N_3473);
nor U4323 (N_4323,N_3097,N_3010);
nand U4324 (N_4324,N_3859,N_3207);
and U4325 (N_4325,N_3498,N_3075);
and U4326 (N_4326,N_3061,N_3273);
and U4327 (N_4327,N_3138,N_3751);
or U4328 (N_4328,N_3971,N_3130);
nand U4329 (N_4329,N_3378,N_3999);
and U4330 (N_4330,N_3886,N_3023);
nor U4331 (N_4331,N_3825,N_3972);
nor U4332 (N_4332,N_3841,N_3171);
xor U4333 (N_4333,N_3989,N_3164);
nand U4334 (N_4334,N_3535,N_3003);
nand U4335 (N_4335,N_3738,N_3179);
nand U4336 (N_4336,N_3438,N_3890);
nor U4337 (N_4337,N_3119,N_3072);
nand U4338 (N_4338,N_3311,N_3495);
nand U4339 (N_4339,N_3797,N_3531);
nand U4340 (N_4340,N_3430,N_3696);
or U4341 (N_4341,N_3081,N_3681);
nand U4342 (N_4342,N_3306,N_3451);
and U4343 (N_4343,N_3818,N_3586);
nor U4344 (N_4344,N_3013,N_3191);
and U4345 (N_4345,N_3437,N_3566);
or U4346 (N_4346,N_3470,N_3526);
nor U4347 (N_4347,N_3975,N_3514);
and U4348 (N_4348,N_3318,N_3630);
and U4349 (N_4349,N_3381,N_3340);
nor U4350 (N_4350,N_3029,N_3390);
nand U4351 (N_4351,N_3973,N_3086);
and U4352 (N_4352,N_3699,N_3140);
and U4353 (N_4353,N_3409,N_3062);
or U4354 (N_4354,N_3525,N_3055);
nor U4355 (N_4355,N_3910,N_3394);
nand U4356 (N_4356,N_3168,N_3953);
or U4357 (N_4357,N_3076,N_3410);
xnor U4358 (N_4358,N_3836,N_3736);
nor U4359 (N_4359,N_3452,N_3042);
or U4360 (N_4360,N_3880,N_3799);
or U4361 (N_4361,N_3780,N_3341);
or U4362 (N_4362,N_3032,N_3915);
xor U4363 (N_4363,N_3234,N_3737);
nand U4364 (N_4364,N_3370,N_3007);
nand U4365 (N_4365,N_3730,N_3885);
nand U4366 (N_4366,N_3992,N_3214);
nor U4367 (N_4367,N_3126,N_3776);
nor U4368 (N_4368,N_3186,N_3006);
and U4369 (N_4369,N_3424,N_3374);
or U4370 (N_4370,N_3239,N_3300);
or U4371 (N_4371,N_3865,N_3122);
or U4372 (N_4372,N_3805,N_3369);
and U4373 (N_4373,N_3930,N_3845);
nor U4374 (N_4374,N_3952,N_3677);
nor U4375 (N_4375,N_3104,N_3143);
and U4376 (N_4376,N_3606,N_3812);
and U4377 (N_4377,N_3489,N_3709);
nor U4378 (N_4378,N_3264,N_3545);
nor U4379 (N_4379,N_3160,N_3950);
nand U4380 (N_4380,N_3977,N_3037);
nand U4381 (N_4381,N_3658,N_3116);
or U4382 (N_4382,N_3120,N_3285);
nor U4383 (N_4383,N_3270,N_3618);
nand U4384 (N_4384,N_3322,N_3852);
nor U4385 (N_4385,N_3769,N_3918);
nand U4386 (N_4386,N_3611,N_3114);
nand U4387 (N_4387,N_3897,N_3155);
and U4388 (N_4388,N_3462,N_3573);
nor U4389 (N_4389,N_3641,N_3914);
xnor U4390 (N_4390,N_3403,N_3581);
or U4391 (N_4391,N_3454,N_3607);
and U4392 (N_4392,N_3310,N_3363);
xnor U4393 (N_4393,N_3827,N_3050);
xor U4394 (N_4394,N_3529,N_3004);
or U4395 (N_4395,N_3507,N_3289);
nor U4396 (N_4396,N_3131,N_3823);
xnor U4397 (N_4397,N_3178,N_3443);
or U4398 (N_4398,N_3259,N_3792);
nand U4399 (N_4399,N_3330,N_3199);
and U4400 (N_4400,N_3628,N_3936);
nor U4401 (N_4401,N_3653,N_3820);
xor U4402 (N_4402,N_3574,N_3631);
and U4403 (N_4403,N_3541,N_3605);
nor U4404 (N_4404,N_3362,N_3281);
xnor U4405 (N_4405,N_3036,N_3896);
and U4406 (N_4406,N_3723,N_3785);
and U4407 (N_4407,N_3663,N_3933);
nand U4408 (N_4408,N_3996,N_3542);
nor U4409 (N_4409,N_3565,N_3772);
nor U4410 (N_4410,N_3719,N_3603);
and U4411 (N_4411,N_3407,N_3420);
and U4412 (N_4412,N_3254,N_3678);
nand U4413 (N_4413,N_3262,N_3647);
or U4414 (N_4414,N_3005,N_3147);
nand U4415 (N_4415,N_3218,N_3052);
nand U4416 (N_4416,N_3434,N_3336);
nand U4417 (N_4417,N_3496,N_3379);
and U4418 (N_4418,N_3208,N_3416);
nor U4419 (N_4419,N_3809,N_3237);
or U4420 (N_4420,N_3521,N_3560);
nand U4421 (N_4421,N_3350,N_3459);
nor U4422 (N_4422,N_3796,N_3480);
nor U4423 (N_4423,N_3598,N_3800);
nand U4424 (N_4424,N_3219,N_3934);
or U4425 (N_4425,N_3537,N_3803);
nor U4426 (N_4426,N_3675,N_3012);
xor U4427 (N_4427,N_3361,N_3040);
and U4428 (N_4428,N_3957,N_3965);
xnor U4429 (N_4429,N_3599,N_3954);
nor U4430 (N_4430,N_3494,N_3509);
nand U4431 (N_4431,N_3320,N_3152);
or U4432 (N_4432,N_3879,N_3071);
xor U4433 (N_4433,N_3626,N_3904);
or U4434 (N_4434,N_3744,N_3148);
nor U4435 (N_4435,N_3145,N_3375);
nand U4436 (N_4436,N_3616,N_3391);
nand U4437 (N_4437,N_3074,N_3620);
and U4438 (N_4438,N_3740,N_3578);
xnor U4439 (N_4439,N_3768,N_3467);
nor U4440 (N_4440,N_3902,N_3761);
nand U4441 (N_4441,N_3401,N_3656);
or U4442 (N_4442,N_3421,N_3739);
nand U4443 (N_4443,N_3327,N_3315);
or U4444 (N_4444,N_3552,N_3659);
or U4445 (N_4445,N_3111,N_3764);
and U4446 (N_4446,N_3745,N_3959);
nor U4447 (N_4447,N_3901,N_3248);
nand U4448 (N_4448,N_3468,N_3015);
or U4449 (N_4449,N_3702,N_3411);
or U4450 (N_4450,N_3227,N_3913);
nor U4451 (N_4451,N_3983,N_3460);
nand U4452 (N_4452,N_3994,N_3344);
or U4453 (N_4453,N_3926,N_3582);
nand U4454 (N_4454,N_3481,N_3843);
and U4455 (N_4455,N_3955,N_3457);
and U4456 (N_4456,N_3085,N_3317);
and U4457 (N_4457,N_3455,N_3619);
or U4458 (N_4458,N_3777,N_3279);
and U4459 (N_4459,N_3862,N_3572);
nor U4460 (N_4460,N_3643,N_3477);
and U4461 (N_4461,N_3813,N_3613);
nor U4462 (N_4462,N_3461,N_3395);
nor U4463 (N_4463,N_3593,N_3041);
and U4464 (N_4464,N_3550,N_3060);
or U4465 (N_4465,N_3655,N_3594);
xnor U4466 (N_4466,N_3196,N_3779);
xnor U4467 (N_4467,N_3860,N_3791);
nor U4468 (N_4468,N_3615,N_3988);
nand U4469 (N_4469,N_3909,N_3808);
nor U4470 (N_4470,N_3472,N_3243);
and U4471 (N_4471,N_3695,N_3874);
or U4472 (N_4472,N_3683,N_3559);
nor U4473 (N_4473,N_3162,N_3313);
and U4474 (N_4474,N_3939,N_3923);
or U4475 (N_4475,N_3019,N_3538);
nor U4476 (N_4476,N_3505,N_3170);
and U4477 (N_4477,N_3303,N_3951);
nor U4478 (N_4478,N_3686,N_3612);
xnor U4479 (N_4479,N_3080,N_3176);
xnor U4480 (N_4480,N_3759,N_3368);
nor U4481 (N_4481,N_3944,N_3257);
nand U4482 (N_4482,N_3127,N_3872);
nor U4483 (N_4483,N_3087,N_3750);
and U4484 (N_4484,N_3899,N_3146);
nor U4485 (N_4485,N_3551,N_3180);
nor U4486 (N_4486,N_3711,N_3624);
or U4487 (N_4487,N_3238,N_3321);
nand U4488 (N_4488,N_3177,N_3834);
xnor U4489 (N_4489,N_3377,N_3386);
nand U4490 (N_4490,N_3077,N_3225);
nand U4491 (N_4491,N_3867,N_3858);
nor U4492 (N_4492,N_3342,N_3555);
nor U4493 (N_4493,N_3637,N_3839);
nor U4494 (N_4494,N_3562,N_3025);
nand U4495 (N_4495,N_3849,N_3432);
or U4496 (N_4496,N_3110,N_3956);
xnor U4497 (N_4497,N_3161,N_3388);
nor U4498 (N_4498,N_3402,N_3520);
or U4499 (N_4499,N_3830,N_3794);
nand U4500 (N_4500,N_3634,N_3176);
nor U4501 (N_4501,N_3645,N_3728);
nor U4502 (N_4502,N_3658,N_3951);
xnor U4503 (N_4503,N_3862,N_3855);
and U4504 (N_4504,N_3600,N_3374);
nand U4505 (N_4505,N_3596,N_3697);
nor U4506 (N_4506,N_3706,N_3354);
and U4507 (N_4507,N_3925,N_3410);
and U4508 (N_4508,N_3076,N_3981);
xor U4509 (N_4509,N_3829,N_3350);
and U4510 (N_4510,N_3001,N_3774);
or U4511 (N_4511,N_3852,N_3425);
and U4512 (N_4512,N_3414,N_3250);
or U4513 (N_4513,N_3972,N_3649);
and U4514 (N_4514,N_3846,N_3154);
nor U4515 (N_4515,N_3536,N_3251);
nand U4516 (N_4516,N_3820,N_3591);
or U4517 (N_4517,N_3112,N_3841);
and U4518 (N_4518,N_3040,N_3619);
nor U4519 (N_4519,N_3432,N_3896);
or U4520 (N_4520,N_3550,N_3723);
xor U4521 (N_4521,N_3833,N_3732);
nor U4522 (N_4522,N_3574,N_3974);
and U4523 (N_4523,N_3059,N_3565);
or U4524 (N_4524,N_3632,N_3998);
or U4525 (N_4525,N_3366,N_3083);
and U4526 (N_4526,N_3850,N_3373);
nand U4527 (N_4527,N_3189,N_3286);
nor U4528 (N_4528,N_3769,N_3015);
or U4529 (N_4529,N_3729,N_3915);
and U4530 (N_4530,N_3037,N_3022);
nand U4531 (N_4531,N_3702,N_3901);
nor U4532 (N_4532,N_3671,N_3297);
nor U4533 (N_4533,N_3749,N_3995);
nor U4534 (N_4534,N_3119,N_3536);
nand U4535 (N_4535,N_3878,N_3611);
and U4536 (N_4536,N_3295,N_3498);
or U4537 (N_4537,N_3664,N_3345);
nand U4538 (N_4538,N_3669,N_3861);
or U4539 (N_4539,N_3760,N_3622);
nand U4540 (N_4540,N_3434,N_3254);
nand U4541 (N_4541,N_3367,N_3380);
nor U4542 (N_4542,N_3319,N_3541);
and U4543 (N_4543,N_3012,N_3533);
or U4544 (N_4544,N_3097,N_3530);
and U4545 (N_4545,N_3677,N_3986);
or U4546 (N_4546,N_3399,N_3032);
or U4547 (N_4547,N_3351,N_3252);
nand U4548 (N_4548,N_3075,N_3356);
or U4549 (N_4549,N_3758,N_3415);
nor U4550 (N_4550,N_3547,N_3137);
and U4551 (N_4551,N_3514,N_3991);
nor U4552 (N_4552,N_3833,N_3280);
or U4553 (N_4553,N_3359,N_3225);
and U4554 (N_4554,N_3658,N_3656);
nor U4555 (N_4555,N_3035,N_3296);
and U4556 (N_4556,N_3439,N_3490);
or U4557 (N_4557,N_3998,N_3436);
or U4558 (N_4558,N_3621,N_3736);
or U4559 (N_4559,N_3204,N_3729);
nor U4560 (N_4560,N_3369,N_3684);
nand U4561 (N_4561,N_3677,N_3830);
or U4562 (N_4562,N_3945,N_3384);
nor U4563 (N_4563,N_3814,N_3207);
and U4564 (N_4564,N_3186,N_3145);
nand U4565 (N_4565,N_3448,N_3339);
nor U4566 (N_4566,N_3755,N_3250);
nor U4567 (N_4567,N_3341,N_3717);
and U4568 (N_4568,N_3002,N_3789);
nand U4569 (N_4569,N_3974,N_3438);
xor U4570 (N_4570,N_3222,N_3068);
nand U4571 (N_4571,N_3410,N_3821);
and U4572 (N_4572,N_3049,N_3169);
and U4573 (N_4573,N_3097,N_3778);
nor U4574 (N_4574,N_3073,N_3628);
nand U4575 (N_4575,N_3579,N_3464);
or U4576 (N_4576,N_3254,N_3095);
nor U4577 (N_4577,N_3873,N_3127);
or U4578 (N_4578,N_3872,N_3663);
nand U4579 (N_4579,N_3115,N_3738);
or U4580 (N_4580,N_3860,N_3033);
nor U4581 (N_4581,N_3269,N_3591);
or U4582 (N_4582,N_3064,N_3652);
or U4583 (N_4583,N_3492,N_3968);
nand U4584 (N_4584,N_3163,N_3432);
nand U4585 (N_4585,N_3480,N_3833);
nand U4586 (N_4586,N_3357,N_3155);
nor U4587 (N_4587,N_3673,N_3058);
and U4588 (N_4588,N_3822,N_3091);
nor U4589 (N_4589,N_3754,N_3449);
nand U4590 (N_4590,N_3055,N_3630);
nor U4591 (N_4591,N_3328,N_3107);
nand U4592 (N_4592,N_3527,N_3538);
and U4593 (N_4593,N_3212,N_3271);
nor U4594 (N_4594,N_3353,N_3506);
and U4595 (N_4595,N_3352,N_3786);
xnor U4596 (N_4596,N_3859,N_3422);
nand U4597 (N_4597,N_3462,N_3979);
or U4598 (N_4598,N_3995,N_3031);
xor U4599 (N_4599,N_3777,N_3088);
or U4600 (N_4600,N_3233,N_3299);
xor U4601 (N_4601,N_3832,N_3490);
or U4602 (N_4602,N_3355,N_3914);
nor U4603 (N_4603,N_3565,N_3256);
and U4604 (N_4604,N_3834,N_3776);
or U4605 (N_4605,N_3674,N_3437);
xnor U4606 (N_4606,N_3846,N_3735);
or U4607 (N_4607,N_3007,N_3878);
xor U4608 (N_4608,N_3299,N_3920);
nand U4609 (N_4609,N_3588,N_3580);
xnor U4610 (N_4610,N_3896,N_3907);
nand U4611 (N_4611,N_3664,N_3521);
nand U4612 (N_4612,N_3549,N_3125);
and U4613 (N_4613,N_3612,N_3045);
or U4614 (N_4614,N_3478,N_3391);
nor U4615 (N_4615,N_3619,N_3651);
nor U4616 (N_4616,N_3778,N_3593);
or U4617 (N_4617,N_3713,N_3387);
and U4618 (N_4618,N_3329,N_3736);
nand U4619 (N_4619,N_3140,N_3147);
xor U4620 (N_4620,N_3128,N_3754);
or U4621 (N_4621,N_3773,N_3235);
and U4622 (N_4622,N_3545,N_3638);
or U4623 (N_4623,N_3614,N_3080);
or U4624 (N_4624,N_3247,N_3461);
or U4625 (N_4625,N_3888,N_3586);
nand U4626 (N_4626,N_3265,N_3803);
nor U4627 (N_4627,N_3803,N_3291);
or U4628 (N_4628,N_3337,N_3839);
xnor U4629 (N_4629,N_3578,N_3152);
and U4630 (N_4630,N_3005,N_3087);
or U4631 (N_4631,N_3723,N_3190);
and U4632 (N_4632,N_3297,N_3714);
and U4633 (N_4633,N_3010,N_3266);
or U4634 (N_4634,N_3162,N_3962);
and U4635 (N_4635,N_3828,N_3184);
nand U4636 (N_4636,N_3876,N_3880);
nand U4637 (N_4637,N_3978,N_3693);
nand U4638 (N_4638,N_3396,N_3817);
and U4639 (N_4639,N_3308,N_3572);
nor U4640 (N_4640,N_3993,N_3949);
xnor U4641 (N_4641,N_3646,N_3095);
xnor U4642 (N_4642,N_3748,N_3285);
nor U4643 (N_4643,N_3740,N_3003);
and U4644 (N_4644,N_3312,N_3326);
nand U4645 (N_4645,N_3388,N_3344);
nor U4646 (N_4646,N_3057,N_3156);
nand U4647 (N_4647,N_3987,N_3916);
nor U4648 (N_4648,N_3617,N_3908);
and U4649 (N_4649,N_3638,N_3977);
or U4650 (N_4650,N_3527,N_3654);
nor U4651 (N_4651,N_3793,N_3925);
and U4652 (N_4652,N_3447,N_3497);
or U4653 (N_4653,N_3956,N_3267);
and U4654 (N_4654,N_3752,N_3657);
and U4655 (N_4655,N_3368,N_3848);
and U4656 (N_4656,N_3480,N_3783);
or U4657 (N_4657,N_3040,N_3267);
xor U4658 (N_4658,N_3535,N_3996);
nand U4659 (N_4659,N_3944,N_3887);
xor U4660 (N_4660,N_3662,N_3314);
or U4661 (N_4661,N_3977,N_3128);
nand U4662 (N_4662,N_3509,N_3515);
nand U4663 (N_4663,N_3811,N_3465);
and U4664 (N_4664,N_3382,N_3318);
and U4665 (N_4665,N_3624,N_3333);
nor U4666 (N_4666,N_3363,N_3671);
xnor U4667 (N_4667,N_3365,N_3715);
nand U4668 (N_4668,N_3839,N_3881);
xnor U4669 (N_4669,N_3480,N_3752);
nand U4670 (N_4670,N_3739,N_3192);
and U4671 (N_4671,N_3301,N_3410);
nor U4672 (N_4672,N_3304,N_3264);
or U4673 (N_4673,N_3957,N_3893);
nand U4674 (N_4674,N_3372,N_3932);
or U4675 (N_4675,N_3746,N_3705);
or U4676 (N_4676,N_3103,N_3914);
nand U4677 (N_4677,N_3702,N_3329);
and U4678 (N_4678,N_3713,N_3745);
or U4679 (N_4679,N_3320,N_3603);
nand U4680 (N_4680,N_3735,N_3937);
or U4681 (N_4681,N_3335,N_3920);
or U4682 (N_4682,N_3048,N_3637);
nor U4683 (N_4683,N_3793,N_3478);
and U4684 (N_4684,N_3139,N_3411);
and U4685 (N_4685,N_3989,N_3191);
nor U4686 (N_4686,N_3684,N_3650);
nor U4687 (N_4687,N_3451,N_3522);
or U4688 (N_4688,N_3378,N_3300);
and U4689 (N_4689,N_3748,N_3738);
xnor U4690 (N_4690,N_3342,N_3529);
xor U4691 (N_4691,N_3196,N_3137);
and U4692 (N_4692,N_3913,N_3927);
nand U4693 (N_4693,N_3582,N_3543);
nand U4694 (N_4694,N_3428,N_3457);
and U4695 (N_4695,N_3392,N_3411);
nor U4696 (N_4696,N_3768,N_3900);
or U4697 (N_4697,N_3232,N_3066);
or U4698 (N_4698,N_3475,N_3711);
nand U4699 (N_4699,N_3787,N_3121);
or U4700 (N_4700,N_3910,N_3058);
or U4701 (N_4701,N_3703,N_3334);
and U4702 (N_4702,N_3190,N_3135);
nand U4703 (N_4703,N_3412,N_3007);
and U4704 (N_4704,N_3330,N_3777);
or U4705 (N_4705,N_3774,N_3154);
or U4706 (N_4706,N_3983,N_3655);
nor U4707 (N_4707,N_3659,N_3004);
xnor U4708 (N_4708,N_3423,N_3188);
xnor U4709 (N_4709,N_3479,N_3821);
nand U4710 (N_4710,N_3573,N_3460);
or U4711 (N_4711,N_3363,N_3883);
nor U4712 (N_4712,N_3084,N_3310);
nand U4713 (N_4713,N_3680,N_3957);
nor U4714 (N_4714,N_3176,N_3717);
and U4715 (N_4715,N_3441,N_3526);
or U4716 (N_4716,N_3411,N_3593);
nand U4717 (N_4717,N_3891,N_3857);
and U4718 (N_4718,N_3650,N_3247);
and U4719 (N_4719,N_3346,N_3744);
and U4720 (N_4720,N_3749,N_3198);
xor U4721 (N_4721,N_3579,N_3021);
or U4722 (N_4722,N_3866,N_3777);
and U4723 (N_4723,N_3417,N_3654);
xor U4724 (N_4724,N_3695,N_3128);
xnor U4725 (N_4725,N_3756,N_3939);
xor U4726 (N_4726,N_3409,N_3864);
and U4727 (N_4727,N_3450,N_3797);
nor U4728 (N_4728,N_3131,N_3277);
and U4729 (N_4729,N_3496,N_3641);
nor U4730 (N_4730,N_3657,N_3285);
nand U4731 (N_4731,N_3740,N_3926);
and U4732 (N_4732,N_3259,N_3980);
or U4733 (N_4733,N_3628,N_3426);
nand U4734 (N_4734,N_3935,N_3746);
nand U4735 (N_4735,N_3057,N_3691);
nor U4736 (N_4736,N_3334,N_3058);
nand U4737 (N_4737,N_3940,N_3651);
or U4738 (N_4738,N_3989,N_3091);
nand U4739 (N_4739,N_3342,N_3381);
or U4740 (N_4740,N_3969,N_3407);
or U4741 (N_4741,N_3671,N_3451);
nand U4742 (N_4742,N_3814,N_3214);
and U4743 (N_4743,N_3347,N_3628);
nor U4744 (N_4744,N_3451,N_3920);
and U4745 (N_4745,N_3589,N_3692);
nand U4746 (N_4746,N_3023,N_3099);
and U4747 (N_4747,N_3896,N_3220);
nor U4748 (N_4748,N_3810,N_3119);
nor U4749 (N_4749,N_3581,N_3666);
and U4750 (N_4750,N_3784,N_3151);
and U4751 (N_4751,N_3912,N_3436);
nor U4752 (N_4752,N_3085,N_3816);
and U4753 (N_4753,N_3269,N_3905);
or U4754 (N_4754,N_3274,N_3337);
nor U4755 (N_4755,N_3394,N_3523);
or U4756 (N_4756,N_3430,N_3159);
nor U4757 (N_4757,N_3078,N_3270);
and U4758 (N_4758,N_3956,N_3241);
nand U4759 (N_4759,N_3553,N_3650);
xor U4760 (N_4760,N_3709,N_3447);
nor U4761 (N_4761,N_3639,N_3368);
nor U4762 (N_4762,N_3123,N_3762);
nand U4763 (N_4763,N_3101,N_3181);
or U4764 (N_4764,N_3171,N_3641);
or U4765 (N_4765,N_3607,N_3447);
or U4766 (N_4766,N_3174,N_3530);
nor U4767 (N_4767,N_3526,N_3698);
nor U4768 (N_4768,N_3468,N_3684);
nand U4769 (N_4769,N_3602,N_3278);
xor U4770 (N_4770,N_3785,N_3452);
nand U4771 (N_4771,N_3521,N_3580);
nor U4772 (N_4772,N_3735,N_3522);
or U4773 (N_4773,N_3514,N_3216);
xor U4774 (N_4774,N_3996,N_3789);
xor U4775 (N_4775,N_3491,N_3447);
or U4776 (N_4776,N_3278,N_3398);
nand U4777 (N_4777,N_3896,N_3323);
and U4778 (N_4778,N_3608,N_3501);
nand U4779 (N_4779,N_3152,N_3736);
nor U4780 (N_4780,N_3361,N_3600);
and U4781 (N_4781,N_3233,N_3284);
or U4782 (N_4782,N_3867,N_3769);
and U4783 (N_4783,N_3704,N_3858);
or U4784 (N_4784,N_3324,N_3525);
and U4785 (N_4785,N_3020,N_3218);
nor U4786 (N_4786,N_3915,N_3670);
nand U4787 (N_4787,N_3628,N_3300);
or U4788 (N_4788,N_3313,N_3056);
nand U4789 (N_4789,N_3264,N_3548);
and U4790 (N_4790,N_3057,N_3075);
or U4791 (N_4791,N_3869,N_3468);
nand U4792 (N_4792,N_3725,N_3987);
and U4793 (N_4793,N_3681,N_3801);
nor U4794 (N_4794,N_3038,N_3562);
nor U4795 (N_4795,N_3796,N_3247);
nand U4796 (N_4796,N_3008,N_3190);
and U4797 (N_4797,N_3325,N_3746);
nand U4798 (N_4798,N_3297,N_3778);
nand U4799 (N_4799,N_3873,N_3685);
nand U4800 (N_4800,N_3610,N_3374);
nand U4801 (N_4801,N_3335,N_3047);
nand U4802 (N_4802,N_3580,N_3530);
and U4803 (N_4803,N_3155,N_3413);
or U4804 (N_4804,N_3944,N_3889);
nor U4805 (N_4805,N_3245,N_3742);
nor U4806 (N_4806,N_3143,N_3110);
nor U4807 (N_4807,N_3144,N_3086);
or U4808 (N_4808,N_3598,N_3331);
or U4809 (N_4809,N_3463,N_3006);
nand U4810 (N_4810,N_3227,N_3687);
and U4811 (N_4811,N_3875,N_3379);
nor U4812 (N_4812,N_3581,N_3431);
nor U4813 (N_4813,N_3241,N_3275);
nor U4814 (N_4814,N_3563,N_3282);
or U4815 (N_4815,N_3251,N_3600);
nand U4816 (N_4816,N_3411,N_3364);
nor U4817 (N_4817,N_3812,N_3053);
xnor U4818 (N_4818,N_3267,N_3979);
and U4819 (N_4819,N_3254,N_3047);
nand U4820 (N_4820,N_3481,N_3403);
and U4821 (N_4821,N_3240,N_3476);
nand U4822 (N_4822,N_3329,N_3321);
or U4823 (N_4823,N_3982,N_3816);
nand U4824 (N_4824,N_3167,N_3349);
nor U4825 (N_4825,N_3639,N_3443);
nor U4826 (N_4826,N_3799,N_3238);
nor U4827 (N_4827,N_3056,N_3533);
nor U4828 (N_4828,N_3970,N_3915);
xor U4829 (N_4829,N_3905,N_3342);
nand U4830 (N_4830,N_3314,N_3050);
xnor U4831 (N_4831,N_3436,N_3457);
nor U4832 (N_4832,N_3368,N_3769);
nor U4833 (N_4833,N_3569,N_3458);
and U4834 (N_4834,N_3535,N_3949);
nor U4835 (N_4835,N_3854,N_3149);
nand U4836 (N_4836,N_3154,N_3692);
or U4837 (N_4837,N_3722,N_3747);
nor U4838 (N_4838,N_3491,N_3888);
and U4839 (N_4839,N_3507,N_3774);
or U4840 (N_4840,N_3721,N_3327);
nand U4841 (N_4841,N_3128,N_3544);
nand U4842 (N_4842,N_3795,N_3420);
nand U4843 (N_4843,N_3844,N_3641);
or U4844 (N_4844,N_3362,N_3674);
xor U4845 (N_4845,N_3418,N_3523);
nand U4846 (N_4846,N_3044,N_3232);
or U4847 (N_4847,N_3705,N_3836);
and U4848 (N_4848,N_3735,N_3091);
xor U4849 (N_4849,N_3134,N_3705);
xnor U4850 (N_4850,N_3859,N_3378);
and U4851 (N_4851,N_3515,N_3392);
xnor U4852 (N_4852,N_3334,N_3142);
xnor U4853 (N_4853,N_3715,N_3448);
nor U4854 (N_4854,N_3448,N_3367);
nor U4855 (N_4855,N_3057,N_3559);
nor U4856 (N_4856,N_3343,N_3616);
nand U4857 (N_4857,N_3284,N_3736);
nand U4858 (N_4858,N_3614,N_3874);
nand U4859 (N_4859,N_3881,N_3212);
nor U4860 (N_4860,N_3736,N_3296);
and U4861 (N_4861,N_3671,N_3477);
nand U4862 (N_4862,N_3155,N_3080);
or U4863 (N_4863,N_3233,N_3961);
or U4864 (N_4864,N_3516,N_3360);
nand U4865 (N_4865,N_3138,N_3774);
and U4866 (N_4866,N_3072,N_3223);
nand U4867 (N_4867,N_3683,N_3125);
or U4868 (N_4868,N_3459,N_3025);
and U4869 (N_4869,N_3652,N_3354);
and U4870 (N_4870,N_3809,N_3750);
and U4871 (N_4871,N_3478,N_3104);
nor U4872 (N_4872,N_3142,N_3387);
or U4873 (N_4873,N_3163,N_3451);
and U4874 (N_4874,N_3796,N_3696);
nor U4875 (N_4875,N_3343,N_3421);
or U4876 (N_4876,N_3096,N_3900);
xnor U4877 (N_4877,N_3520,N_3881);
nand U4878 (N_4878,N_3870,N_3089);
nand U4879 (N_4879,N_3583,N_3856);
or U4880 (N_4880,N_3443,N_3309);
nand U4881 (N_4881,N_3484,N_3908);
and U4882 (N_4882,N_3164,N_3960);
nand U4883 (N_4883,N_3542,N_3210);
xnor U4884 (N_4884,N_3366,N_3552);
and U4885 (N_4885,N_3576,N_3822);
or U4886 (N_4886,N_3924,N_3197);
nand U4887 (N_4887,N_3021,N_3905);
or U4888 (N_4888,N_3360,N_3299);
nor U4889 (N_4889,N_3584,N_3965);
xnor U4890 (N_4890,N_3862,N_3391);
and U4891 (N_4891,N_3526,N_3694);
nor U4892 (N_4892,N_3216,N_3852);
xnor U4893 (N_4893,N_3880,N_3050);
nor U4894 (N_4894,N_3605,N_3630);
nand U4895 (N_4895,N_3982,N_3004);
and U4896 (N_4896,N_3127,N_3621);
xor U4897 (N_4897,N_3172,N_3066);
and U4898 (N_4898,N_3890,N_3743);
or U4899 (N_4899,N_3246,N_3691);
or U4900 (N_4900,N_3997,N_3855);
and U4901 (N_4901,N_3131,N_3993);
nor U4902 (N_4902,N_3179,N_3389);
or U4903 (N_4903,N_3572,N_3972);
nand U4904 (N_4904,N_3952,N_3820);
nor U4905 (N_4905,N_3708,N_3090);
nor U4906 (N_4906,N_3902,N_3065);
or U4907 (N_4907,N_3267,N_3628);
nor U4908 (N_4908,N_3223,N_3999);
nor U4909 (N_4909,N_3206,N_3975);
nor U4910 (N_4910,N_3009,N_3593);
nand U4911 (N_4911,N_3223,N_3827);
nor U4912 (N_4912,N_3189,N_3246);
or U4913 (N_4913,N_3944,N_3911);
xor U4914 (N_4914,N_3082,N_3072);
nor U4915 (N_4915,N_3451,N_3612);
or U4916 (N_4916,N_3424,N_3410);
and U4917 (N_4917,N_3202,N_3599);
or U4918 (N_4918,N_3218,N_3054);
nor U4919 (N_4919,N_3976,N_3796);
nand U4920 (N_4920,N_3164,N_3204);
or U4921 (N_4921,N_3453,N_3340);
or U4922 (N_4922,N_3037,N_3728);
nor U4923 (N_4923,N_3995,N_3522);
nor U4924 (N_4924,N_3958,N_3333);
and U4925 (N_4925,N_3668,N_3315);
or U4926 (N_4926,N_3077,N_3668);
xor U4927 (N_4927,N_3970,N_3855);
and U4928 (N_4928,N_3889,N_3471);
nand U4929 (N_4929,N_3206,N_3835);
xor U4930 (N_4930,N_3107,N_3765);
nand U4931 (N_4931,N_3282,N_3168);
nand U4932 (N_4932,N_3290,N_3020);
xor U4933 (N_4933,N_3339,N_3512);
nor U4934 (N_4934,N_3021,N_3580);
and U4935 (N_4935,N_3818,N_3043);
or U4936 (N_4936,N_3775,N_3900);
xor U4937 (N_4937,N_3590,N_3990);
nor U4938 (N_4938,N_3927,N_3660);
nand U4939 (N_4939,N_3162,N_3135);
nand U4940 (N_4940,N_3619,N_3928);
and U4941 (N_4941,N_3755,N_3915);
xor U4942 (N_4942,N_3961,N_3765);
nor U4943 (N_4943,N_3881,N_3609);
xnor U4944 (N_4944,N_3146,N_3449);
nor U4945 (N_4945,N_3576,N_3400);
or U4946 (N_4946,N_3178,N_3647);
or U4947 (N_4947,N_3404,N_3643);
or U4948 (N_4948,N_3877,N_3569);
nor U4949 (N_4949,N_3956,N_3651);
and U4950 (N_4950,N_3205,N_3278);
nor U4951 (N_4951,N_3727,N_3374);
nor U4952 (N_4952,N_3347,N_3234);
and U4953 (N_4953,N_3396,N_3825);
and U4954 (N_4954,N_3206,N_3877);
nand U4955 (N_4955,N_3889,N_3632);
xor U4956 (N_4956,N_3910,N_3793);
and U4957 (N_4957,N_3359,N_3577);
and U4958 (N_4958,N_3996,N_3017);
or U4959 (N_4959,N_3919,N_3876);
xor U4960 (N_4960,N_3892,N_3490);
and U4961 (N_4961,N_3724,N_3450);
or U4962 (N_4962,N_3860,N_3425);
nand U4963 (N_4963,N_3925,N_3880);
and U4964 (N_4964,N_3485,N_3619);
nor U4965 (N_4965,N_3870,N_3379);
and U4966 (N_4966,N_3786,N_3647);
and U4967 (N_4967,N_3305,N_3892);
nor U4968 (N_4968,N_3532,N_3049);
nand U4969 (N_4969,N_3206,N_3926);
xor U4970 (N_4970,N_3182,N_3322);
nand U4971 (N_4971,N_3974,N_3929);
and U4972 (N_4972,N_3757,N_3584);
nand U4973 (N_4973,N_3591,N_3078);
nor U4974 (N_4974,N_3120,N_3167);
or U4975 (N_4975,N_3633,N_3975);
xnor U4976 (N_4976,N_3970,N_3941);
or U4977 (N_4977,N_3590,N_3501);
or U4978 (N_4978,N_3661,N_3014);
and U4979 (N_4979,N_3297,N_3614);
nand U4980 (N_4980,N_3927,N_3901);
nor U4981 (N_4981,N_3421,N_3001);
or U4982 (N_4982,N_3776,N_3769);
or U4983 (N_4983,N_3713,N_3453);
nand U4984 (N_4984,N_3604,N_3186);
and U4985 (N_4985,N_3338,N_3284);
or U4986 (N_4986,N_3506,N_3101);
nand U4987 (N_4987,N_3964,N_3228);
xor U4988 (N_4988,N_3733,N_3383);
or U4989 (N_4989,N_3082,N_3388);
xor U4990 (N_4990,N_3864,N_3139);
nand U4991 (N_4991,N_3865,N_3498);
nor U4992 (N_4992,N_3662,N_3328);
nor U4993 (N_4993,N_3231,N_3232);
nor U4994 (N_4994,N_3993,N_3777);
nor U4995 (N_4995,N_3040,N_3237);
nand U4996 (N_4996,N_3079,N_3846);
xor U4997 (N_4997,N_3648,N_3628);
and U4998 (N_4998,N_3078,N_3198);
xor U4999 (N_4999,N_3549,N_3870);
nor UO_0 (O_0,N_4621,N_4484);
and UO_1 (O_1,N_4222,N_4155);
or UO_2 (O_2,N_4661,N_4398);
and UO_3 (O_3,N_4157,N_4032);
or UO_4 (O_4,N_4173,N_4938);
nand UO_5 (O_5,N_4952,N_4551);
xnor UO_6 (O_6,N_4322,N_4646);
nand UO_7 (O_7,N_4994,N_4557);
nor UO_8 (O_8,N_4019,N_4345);
nor UO_9 (O_9,N_4587,N_4811);
and UO_10 (O_10,N_4654,N_4995);
nand UO_11 (O_11,N_4614,N_4919);
nand UO_12 (O_12,N_4888,N_4151);
and UO_13 (O_13,N_4179,N_4884);
and UO_14 (O_14,N_4441,N_4357);
and UO_15 (O_15,N_4000,N_4846);
nor UO_16 (O_16,N_4803,N_4918);
and UO_17 (O_17,N_4027,N_4148);
nand UO_18 (O_18,N_4313,N_4762);
xor UO_19 (O_19,N_4801,N_4527);
nor UO_20 (O_20,N_4407,N_4715);
xor UO_21 (O_21,N_4930,N_4867);
xor UO_22 (O_22,N_4003,N_4556);
nand UO_23 (O_23,N_4181,N_4028);
or UO_24 (O_24,N_4100,N_4649);
nand UO_25 (O_25,N_4102,N_4237);
nor UO_26 (O_26,N_4008,N_4010);
or UO_27 (O_27,N_4460,N_4143);
xnor UO_28 (O_28,N_4545,N_4477);
nor UO_29 (O_29,N_4030,N_4087);
nor UO_30 (O_30,N_4560,N_4285);
nor UO_31 (O_31,N_4754,N_4763);
nor UO_32 (O_32,N_4134,N_4929);
nand UO_33 (O_33,N_4933,N_4240);
nand UO_34 (O_34,N_4721,N_4057);
xor UO_35 (O_35,N_4203,N_4388);
and UO_36 (O_36,N_4841,N_4936);
xor UO_37 (O_37,N_4164,N_4312);
nand UO_38 (O_38,N_4116,N_4332);
or UO_39 (O_39,N_4080,N_4466);
nor UO_40 (O_40,N_4139,N_4049);
or UO_41 (O_41,N_4468,N_4140);
nand UO_42 (O_42,N_4603,N_4448);
or UO_43 (O_43,N_4656,N_4483);
xor UO_44 (O_44,N_4061,N_4768);
nand UO_45 (O_45,N_4463,N_4426);
xnor UO_46 (O_46,N_4009,N_4177);
nand UO_47 (O_47,N_4992,N_4074);
and UO_48 (O_48,N_4403,N_4439);
and UO_49 (O_49,N_4026,N_4373);
nand UO_50 (O_50,N_4872,N_4892);
xnor UO_51 (O_51,N_4590,N_4889);
nor UO_52 (O_52,N_4939,N_4834);
and UO_53 (O_53,N_4899,N_4200);
nand UO_54 (O_54,N_4982,N_4396);
or UO_55 (O_55,N_4437,N_4209);
or UO_56 (O_56,N_4178,N_4981);
nand UO_57 (O_57,N_4001,N_4276);
and UO_58 (O_58,N_4714,N_4537);
nor UO_59 (O_59,N_4683,N_4362);
or UO_60 (O_60,N_4904,N_4651);
nand UO_61 (O_61,N_4898,N_4883);
nor UO_62 (O_62,N_4152,N_4130);
nor UO_63 (O_63,N_4894,N_4381);
nand UO_64 (O_64,N_4252,N_4171);
and UO_65 (O_65,N_4789,N_4137);
or UO_66 (O_66,N_4999,N_4135);
and UO_67 (O_67,N_4795,N_4820);
nand UO_68 (O_68,N_4214,N_4832);
nor UO_69 (O_69,N_4607,N_4355);
nand UO_70 (O_70,N_4953,N_4695);
nand UO_71 (O_71,N_4062,N_4085);
or UO_72 (O_72,N_4827,N_4497);
nand UO_73 (O_73,N_4895,N_4666);
or UO_74 (O_74,N_4329,N_4605);
nand UO_75 (O_75,N_4572,N_4415);
and UO_76 (O_76,N_4273,N_4977);
nor UO_77 (O_77,N_4160,N_4422);
or UO_78 (O_78,N_4502,N_4594);
or UO_79 (O_79,N_4309,N_4948);
and UO_80 (O_80,N_4735,N_4413);
nor UO_81 (O_81,N_4186,N_4903);
nand UO_82 (O_82,N_4119,N_4772);
and UO_83 (O_83,N_4491,N_4984);
nor UO_84 (O_84,N_4519,N_4391);
xnor UO_85 (O_85,N_4574,N_4686);
nor UO_86 (O_86,N_4769,N_4593);
nor UO_87 (O_87,N_4700,N_4089);
nand UO_88 (O_88,N_4395,N_4427);
or UO_89 (O_89,N_4558,N_4434);
nand UO_90 (O_90,N_4779,N_4744);
and UO_91 (O_91,N_4464,N_4311);
nand UO_92 (O_92,N_4238,N_4333);
nor UO_93 (O_93,N_4138,N_4166);
or UO_94 (O_94,N_4923,N_4927);
nor UO_95 (O_95,N_4577,N_4124);
nor UO_96 (O_96,N_4792,N_4047);
or UO_97 (O_97,N_4696,N_4011);
xnor UO_98 (O_98,N_4882,N_4924);
or UO_99 (O_99,N_4813,N_4455);
nor UO_100 (O_100,N_4153,N_4486);
or UO_101 (O_101,N_4053,N_4900);
nand UO_102 (O_102,N_4839,N_4886);
or UO_103 (O_103,N_4111,N_4370);
and UO_104 (O_104,N_4891,N_4728);
nor UO_105 (O_105,N_4824,N_4347);
or UO_106 (O_106,N_4255,N_4976);
or UO_107 (O_107,N_4665,N_4679);
nor UO_108 (O_108,N_4295,N_4267);
and UO_109 (O_109,N_4669,N_4073);
nor UO_110 (O_110,N_4514,N_4759);
nand UO_111 (O_111,N_4419,N_4726);
nand UO_112 (O_112,N_4299,N_4488);
or UO_113 (O_113,N_4457,N_4809);
and UO_114 (O_114,N_4020,N_4873);
and UO_115 (O_115,N_4453,N_4851);
or UO_116 (O_116,N_4505,N_4440);
xor UO_117 (O_117,N_4647,N_4349);
or UO_118 (O_118,N_4132,N_4243);
xnor UO_119 (O_119,N_4829,N_4423);
or UO_120 (O_120,N_4787,N_4245);
and UO_121 (O_121,N_4580,N_4499);
and UO_122 (O_122,N_4893,N_4231);
nand UO_123 (O_123,N_4296,N_4302);
or UO_124 (O_124,N_4861,N_4376);
xor UO_125 (O_125,N_4268,N_4401);
or UO_126 (O_126,N_4781,N_4432);
nor UO_127 (O_127,N_4664,N_4963);
nand UO_128 (O_128,N_4293,N_4371);
nor UO_129 (O_129,N_4251,N_4390);
nor UO_130 (O_130,N_4562,N_4622);
nor UO_131 (O_131,N_4420,N_4775);
nor UO_132 (O_132,N_4879,N_4778);
nand UO_133 (O_133,N_4458,N_4967);
nand UO_134 (O_134,N_4636,N_4798);
or UO_135 (O_135,N_4288,N_4335);
xnor UO_136 (O_136,N_4504,N_4360);
nand UO_137 (O_137,N_4914,N_4814);
nor UO_138 (O_138,N_4777,N_4599);
nand UO_139 (O_139,N_4123,N_4785);
nor UO_140 (O_140,N_4986,N_4041);
nor UO_141 (O_141,N_4091,N_4910);
and UO_142 (O_142,N_4985,N_4474);
and UO_143 (O_143,N_4732,N_4961);
and UO_144 (O_144,N_4857,N_4808);
and UO_145 (O_145,N_4642,N_4624);
nand UO_146 (O_146,N_4196,N_4328);
xnor UO_147 (O_147,N_4536,N_4430);
nor UO_148 (O_148,N_4084,N_4175);
or UO_149 (O_149,N_4561,N_4418);
xnor UO_150 (O_150,N_4366,N_4617);
or UO_151 (O_151,N_4416,N_4860);
nor UO_152 (O_152,N_4090,N_4611);
or UO_153 (O_153,N_4589,N_4467);
nand UO_154 (O_154,N_4826,N_4690);
and UO_155 (O_155,N_4350,N_4257);
nor UO_156 (O_156,N_4048,N_4385);
xnor UO_157 (O_157,N_4109,N_4653);
nand UO_158 (O_158,N_4670,N_4018);
nor UO_159 (O_159,N_4216,N_4657);
and UO_160 (O_160,N_4272,N_4342);
nor UO_161 (O_161,N_4142,N_4088);
nor UO_162 (O_162,N_4591,N_4250);
and UO_163 (O_163,N_4597,N_4940);
xnor UO_164 (O_164,N_4723,N_4006);
nand UO_165 (O_165,N_4115,N_4247);
or UO_166 (O_166,N_4812,N_4136);
nand UO_167 (O_167,N_4344,N_4405);
nand UO_168 (O_168,N_4103,N_4106);
nand UO_169 (O_169,N_4549,N_4912);
nor UO_170 (O_170,N_4040,N_4495);
or UO_171 (O_171,N_4643,N_4644);
nor UO_172 (O_172,N_4128,N_4921);
or UO_173 (O_173,N_4379,N_4212);
nand UO_174 (O_174,N_4613,N_4338);
nand UO_175 (O_175,N_4655,N_4424);
nor UO_176 (O_176,N_4263,N_4627);
and UO_177 (O_177,N_4648,N_4325);
nor UO_178 (O_178,N_4104,N_4915);
nor UO_179 (O_179,N_4067,N_4278);
nand UO_180 (O_180,N_4797,N_4635);
nor UO_181 (O_181,N_4583,N_4187);
xor UO_182 (O_182,N_4513,N_4146);
or UO_183 (O_183,N_4210,N_4363);
nand UO_184 (O_184,N_4304,N_4596);
and UO_185 (O_185,N_4663,N_4640);
xor UO_186 (O_186,N_4083,N_4844);
nor UO_187 (O_187,N_4571,N_4710);
nor UO_188 (O_188,N_4188,N_4117);
nor UO_189 (O_189,N_4359,N_4863);
or UO_190 (O_190,N_4880,N_4748);
or UO_191 (O_191,N_4511,N_4897);
nor UO_192 (O_192,N_4682,N_4756);
nand UO_193 (O_193,N_4356,N_4875);
nand UO_194 (O_194,N_4244,N_4671);
or UO_195 (O_195,N_4747,N_4071);
nor UO_196 (O_196,N_4351,N_4725);
nand UO_197 (O_197,N_4110,N_4226);
or UO_198 (O_198,N_4786,N_4552);
nand UO_199 (O_199,N_4184,N_4539);
and UO_200 (O_200,N_4584,N_4874);
nor UO_201 (O_201,N_4052,N_4485);
and UO_202 (O_202,N_4678,N_4633);
or UO_203 (O_203,N_4126,N_4202);
and UO_204 (O_204,N_4063,N_4757);
and UO_205 (O_205,N_4819,N_4694);
nand UO_206 (O_206,N_4075,N_4380);
xor UO_207 (O_207,N_4836,N_4668);
or UO_208 (O_208,N_4955,N_4553);
and UO_209 (O_209,N_4487,N_4764);
and UO_210 (O_210,N_4167,N_4782);
and UO_211 (O_211,N_4616,N_4689);
and UO_212 (O_212,N_4855,N_4742);
nand UO_213 (O_213,N_4374,N_4034);
and UO_214 (O_214,N_4699,N_4409);
and UO_215 (O_215,N_4529,N_4980);
nand UO_216 (O_216,N_4559,N_4261);
nand UO_217 (O_217,N_4174,N_4258);
nand UO_218 (O_218,N_4364,N_4015);
and UO_219 (O_219,N_4249,N_4479);
nand UO_220 (O_220,N_4069,N_4528);
nor UO_221 (O_221,N_4223,N_4909);
and UO_222 (O_222,N_4802,N_4966);
and UO_223 (O_223,N_4521,N_4997);
and UO_224 (O_224,N_4219,N_4968);
and UO_225 (O_225,N_4675,N_4993);
nor UO_226 (O_226,N_4290,N_4264);
nand UO_227 (O_227,N_4585,N_4530);
nor UO_228 (O_228,N_4489,N_4677);
or UO_229 (O_229,N_4901,N_4220);
nor UO_230 (O_230,N_4831,N_4248);
nand UO_231 (O_231,N_4538,N_4758);
nand UO_232 (O_232,N_4014,N_4931);
nor UO_233 (O_233,N_4190,N_4566);
nand UO_234 (O_234,N_4406,N_4473);
or UO_235 (O_235,N_4729,N_4937);
nor UO_236 (O_236,N_4793,N_4568);
and UO_237 (O_237,N_4625,N_4316);
nand UO_238 (O_238,N_4512,N_4573);
or UO_239 (O_239,N_4975,N_4971);
nand UO_240 (O_240,N_4154,N_4331);
nor UO_241 (O_241,N_4158,N_4180);
nand UO_242 (O_242,N_4445,N_4932);
nor UO_243 (O_243,N_4701,N_4945);
xor UO_244 (O_244,N_4547,N_4038);
nor UO_245 (O_245,N_4369,N_4749);
nor UO_246 (O_246,N_4450,N_4676);
and UO_247 (O_247,N_4876,N_4131);
xor UO_248 (O_248,N_4673,N_4691);
nor UO_249 (O_249,N_4305,N_4818);
and UO_250 (O_250,N_4541,N_4506);
nand UO_251 (O_251,N_4957,N_4282);
and UO_252 (O_252,N_4230,N_4943);
or UO_253 (O_253,N_4926,N_4470);
or UO_254 (O_254,N_4619,N_4372);
and UO_255 (O_255,N_4232,N_4662);
and UO_256 (O_256,N_4520,N_4830);
nand UO_257 (O_257,N_4964,N_4442);
nand UO_258 (O_258,N_4478,N_4501);
and UO_259 (O_259,N_4806,N_4327);
or UO_260 (O_260,N_4389,N_4862);
and UO_261 (O_261,N_4215,N_4490);
and UO_262 (O_262,N_4630,N_4865);
and UO_263 (O_263,N_4581,N_4543);
xnor UO_264 (O_264,N_4022,N_4482);
xnor UO_265 (O_265,N_4070,N_4796);
nor UO_266 (O_266,N_4548,N_4496);
or UO_267 (O_267,N_4972,N_4550);
or UO_268 (O_268,N_4274,N_4760);
nor UO_269 (O_269,N_4554,N_4421);
xnor UO_270 (O_270,N_4270,N_4916);
nand UO_271 (O_271,N_4731,N_4822);
and UO_272 (O_272,N_4852,N_4843);
and UO_273 (O_273,N_4576,N_4012);
and UO_274 (O_274,N_4825,N_4693);
or UO_275 (O_275,N_4459,N_4618);
or UO_276 (O_276,N_4291,N_4408);
and UO_277 (O_277,N_4784,N_4878);
or UO_278 (O_278,N_4353,N_4498);
nor UO_279 (O_279,N_4848,N_4213);
nor UO_280 (O_280,N_4169,N_4095);
xnor UO_281 (O_281,N_4632,N_4265);
and UO_282 (O_282,N_4579,N_4096);
nor UO_283 (O_283,N_4612,N_4628);
or UO_284 (O_284,N_4833,N_4301);
and UO_285 (O_285,N_4835,N_4847);
xor UO_286 (O_286,N_4869,N_4780);
nor UO_287 (O_287,N_4224,N_4905);
nand UO_288 (O_288,N_4503,N_4638);
or UO_289 (O_289,N_4383,N_4911);
or UO_290 (O_290,N_4234,N_4908);
xor UO_291 (O_291,N_4650,N_4535);
nand UO_292 (O_292,N_4586,N_4133);
nor UO_293 (O_293,N_4277,N_4674);
nand UO_294 (O_294,N_4051,N_4564);
or UO_295 (O_295,N_4704,N_4703);
or UO_296 (O_296,N_4254,N_4194);
or UO_297 (O_297,N_4280,N_4228);
and UO_298 (O_298,N_4941,N_4658);
nand UO_299 (O_299,N_4033,N_4377);
or UO_300 (O_300,N_4609,N_4688);
nor UO_301 (O_301,N_4037,N_4339);
nor UO_302 (O_302,N_4524,N_4570);
nand UO_303 (O_303,N_4031,N_4161);
nand UO_304 (O_304,N_4563,N_4600);
and UO_305 (O_305,N_4685,N_4319);
nor UO_306 (O_306,N_4509,N_4864);
or UO_307 (O_307,N_4122,N_4533);
and UO_308 (O_308,N_4354,N_4292);
nand UO_309 (O_309,N_4745,N_4361);
and UO_310 (O_310,N_4773,N_4739);
or UO_311 (O_311,N_4269,N_4791);
xnor UO_312 (O_312,N_4626,N_4208);
or UO_313 (O_313,N_4141,N_4711);
nand UO_314 (O_314,N_4326,N_4615);
or UO_315 (O_315,N_4013,N_4741);
and UO_316 (O_316,N_4517,N_4058);
xnor UO_317 (O_317,N_4023,N_4266);
and UO_318 (O_318,N_4217,N_4598);
and UO_319 (O_319,N_4532,N_4330);
nand UO_320 (O_320,N_4065,N_4471);
nand UO_321 (O_321,N_4507,N_4854);
or UO_322 (O_322,N_4392,N_4059);
or UO_323 (O_323,N_4225,N_4944);
nand UO_324 (O_324,N_4881,N_4534);
xor UO_325 (O_325,N_4709,N_4838);
or UO_326 (O_326,N_4823,N_4771);
nor UO_327 (O_327,N_4516,N_4870);
nand UO_328 (O_328,N_4235,N_4114);
and UO_329 (O_329,N_4227,N_4365);
and UO_330 (O_330,N_4306,N_4716);
xnor UO_331 (O_331,N_4805,N_4645);
nor UO_332 (O_332,N_4949,N_4093);
nor UO_333 (O_333,N_4702,N_4191);
or UO_334 (O_334,N_4284,N_4454);
or UO_335 (O_335,N_4447,N_4956);
xnor UO_336 (O_336,N_4565,N_4717);
nor UO_337 (O_337,N_4428,N_4736);
xor UO_338 (O_338,N_4260,N_4954);
and UO_339 (O_339,N_4400,N_4713);
nor UO_340 (O_340,N_4346,N_4404);
nor UO_341 (O_341,N_4159,N_4525);
nor UO_342 (O_342,N_4724,N_4452);
or UO_343 (O_343,N_4774,N_4303);
nor UO_344 (O_344,N_4472,N_4950);
nand UO_345 (O_345,N_4121,N_4871);
xor UO_346 (O_346,N_4170,N_4770);
and UO_347 (O_347,N_4567,N_4253);
nor UO_348 (O_348,N_4750,N_4147);
and UO_349 (O_349,N_4016,N_4435);
or UO_350 (O_350,N_4336,N_4951);
nor UO_351 (O_351,N_4352,N_4575);
and UO_352 (O_352,N_4068,N_4969);
and UO_353 (O_353,N_4438,N_4456);
and UO_354 (O_354,N_4907,N_4201);
nor UO_355 (O_355,N_4712,N_4958);
and UO_356 (O_356,N_4105,N_4024);
and UO_357 (O_357,N_4540,N_4606);
and UO_358 (O_358,N_4120,N_4531);
and UO_359 (O_359,N_4680,N_4206);
nor UO_360 (O_360,N_4718,N_4378);
or UO_361 (O_361,N_4283,N_4500);
nor UO_362 (O_362,N_4233,N_4799);
nand UO_363 (O_363,N_4198,N_4172);
or UO_364 (O_364,N_4790,N_4842);
and UO_365 (O_365,N_4054,N_4965);
or UO_366 (O_366,N_4947,N_4515);
or UO_367 (O_367,N_4917,N_4340);
or UO_368 (O_368,N_4687,N_4281);
and UO_369 (O_369,N_4144,N_4021);
nor UO_370 (O_370,N_4286,N_4108);
and UO_371 (O_371,N_4125,N_4522);
nor UO_372 (O_372,N_4239,N_4608);
nor UO_373 (O_373,N_4508,N_4555);
nor UO_374 (O_374,N_4099,N_4307);
nor UO_375 (O_375,N_4197,N_4730);
nand UO_376 (O_376,N_4315,N_4076);
and UO_377 (O_377,N_4990,N_4588);
nand UO_378 (O_378,N_4294,N_4631);
and UO_379 (O_379,N_4236,N_4287);
or UO_380 (O_380,N_4868,N_4481);
nand UO_381 (O_381,N_4242,N_4107);
and UO_382 (O_382,N_4761,N_4610);
nor UO_383 (O_383,N_4946,N_4176);
nor UO_384 (O_384,N_4297,N_4082);
and UO_385 (O_385,N_4317,N_4518);
and UO_386 (O_386,N_4794,N_4998);
and UO_387 (O_387,N_4837,N_4629);
and UO_388 (O_388,N_4358,N_4207);
xnor UO_389 (O_389,N_4959,N_4480);
and UO_390 (O_390,N_4623,N_4475);
or UO_391 (O_391,N_4412,N_4890);
and UO_392 (O_392,N_4042,N_4150);
and UO_393 (O_393,N_4368,N_4776);
or UO_394 (O_394,N_4595,N_4321);
nor UO_395 (O_395,N_4367,N_4444);
nand UO_396 (O_396,N_4436,N_4417);
xor UO_397 (O_397,N_4410,N_4204);
and UO_398 (O_398,N_4753,N_4205);
or UO_399 (O_399,N_4705,N_4765);
nand UO_400 (O_400,N_4751,N_4324);
or UO_401 (O_401,N_4348,N_4259);
xor UO_402 (O_402,N_4928,N_4620);
or UO_403 (O_403,N_4913,N_4411);
nor UO_404 (O_404,N_4896,N_4433);
xnor UO_405 (O_405,N_4393,N_4523);
and UO_406 (O_406,N_4182,N_4816);
or UO_407 (O_407,N_4189,N_4341);
and UO_408 (O_408,N_4526,N_4094);
nor UO_409 (O_409,N_4004,N_4044);
nor UO_410 (O_410,N_4449,N_4853);
nand UO_411 (O_411,N_4569,N_4810);
or UO_412 (O_412,N_4920,N_4334);
nor UO_413 (O_413,N_4767,N_4382);
nor UO_414 (O_414,N_4241,N_4828);
nand UO_415 (O_415,N_4469,N_4113);
and UO_416 (O_416,N_4046,N_4192);
nor UO_417 (O_417,N_4746,N_4604);
nand UO_418 (O_418,N_4199,N_4960);
nand UO_419 (O_419,N_4592,N_4845);
and UO_420 (O_420,N_4394,N_4807);
xnor UO_421 (O_421,N_4856,N_4318);
nand UO_422 (O_422,N_4218,N_4601);
and UO_423 (O_423,N_4145,N_4298);
xor UO_424 (O_424,N_4989,N_4906);
or UO_425 (O_425,N_4935,N_4431);
nor UO_426 (O_426,N_4005,N_4743);
nor UO_427 (O_427,N_4246,N_4050);
and UO_428 (O_428,N_4492,N_4667);
and UO_429 (O_429,N_4849,N_4733);
nor UO_430 (O_430,N_4300,N_4337);
nor UO_431 (O_431,N_4275,N_4195);
xnor UO_432 (O_432,N_4308,N_4112);
or UO_433 (O_433,N_4766,N_4800);
and UO_434 (O_434,N_4451,N_4817);
and UO_435 (O_435,N_4310,N_4185);
xor UO_436 (O_436,N_4788,N_4988);
nor UO_437 (O_437,N_4978,N_4397);
or UO_438 (O_438,N_4462,N_4602);
nand UO_439 (O_439,N_4493,N_4887);
and UO_440 (O_440,N_4399,N_4461);
nand UO_441 (O_441,N_4162,N_4221);
or UO_442 (O_442,N_4706,N_4077);
nand UO_443 (O_443,N_4996,N_4979);
xor UO_444 (O_444,N_4323,N_4098);
nand UO_445 (O_445,N_4414,N_4755);
and UO_446 (O_446,N_4850,N_4320);
or UO_447 (O_447,N_4165,N_4017);
or UO_448 (O_448,N_4025,N_4078);
and UO_449 (O_449,N_4375,N_4737);
and UO_450 (O_450,N_4002,N_4056);
or UO_451 (O_451,N_4858,N_4582);
nor UO_452 (O_452,N_4652,N_4229);
or UO_453 (O_453,N_4045,N_4544);
nand UO_454 (O_454,N_4866,N_4804);
nand UO_455 (O_455,N_4314,N_4055);
nand UO_456 (O_456,N_4722,N_4064);
and UO_457 (O_457,N_4681,N_4429);
nor UO_458 (O_458,N_4684,N_4035);
nor UO_459 (O_459,N_4885,N_4081);
and UO_460 (O_460,N_4343,N_4922);
nor UO_461 (O_461,N_4129,N_4720);
and UO_462 (O_462,N_4659,N_4494);
nor UO_463 (O_463,N_4211,N_4402);
and UO_464 (O_464,N_4902,N_4127);
nor UO_465 (O_465,N_4925,N_4386);
or UO_466 (O_466,N_4859,N_4707);
nor UO_467 (O_467,N_4719,N_4546);
nand UO_468 (O_468,N_4072,N_4672);
nor UO_469 (O_469,N_4101,N_4256);
xor UO_470 (O_470,N_4740,N_4708);
nor UO_471 (O_471,N_4476,N_4036);
nand UO_472 (O_472,N_4443,N_4942);
and UO_473 (O_473,N_4387,N_4738);
or UO_474 (O_474,N_4446,N_4156);
nor UO_475 (O_475,N_4465,N_4641);
or UO_476 (O_476,N_4634,N_4692);
and UO_477 (O_477,N_4149,N_4970);
or UO_478 (O_478,N_4987,N_4697);
nand UO_479 (O_479,N_4637,N_4983);
nor UO_480 (O_480,N_4973,N_4962);
nor UO_481 (O_481,N_4815,N_4163);
or UO_482 (O_482,N_4043,N_4727);
nand UO_483 (O_483,N_4991,N_4578);
or UO_484 (O_484,N_4752,N_4097);
and UO_485 (O_485,N_4289,N_4974);
nor UO_486 (O_486,N_4086,N_4262);
nor UO_487 (O_487,N_4118,N_4279);
or UO_488 (O_488,N_4734,N_4007);
nor UO_489 (O_489,N_4542,N_4039);
nor UO_490 (O_490,N_4183,N_4079);
nand UO_491 (O_491,N_4060,N_4168);
nor UO_492 (O_492,N_4821,N_4639);
nor UO_493 (O_493,N_4934,N_4029);
nand UO_494 (O_494,N_4783,N_4066);
or UO_495 (O_495,N_4877,N_4510);
and UO_496 (O_496,N_4193,N_4271);
and UO_497 (O_497,N_4092,N_4660);
nand UO_498 (O_498,N_4698,N_4384);
nand UO_499 (O_499,N_4425,N_4840);
nor UO_500 (O_500,N_4803,N_4239);
or UO_501 (O_501,N_4288,N_4997);
nand UO_502 (O_502,N_4949,N_4821);
and UO_503 (O_503,N_4034,N_4163);
and UO_504 (O_504,N_4104,N_4539);
nor UO_505 (O_505,N_4160,N_4218);
xor UO_506 (O_506,N_4414,N_4551);
or UO_507 (O_507,N_4525,N_4089);
or UO_508 (O_508,N_4112,N_4244);
nand UO_509 (O_509,N_4972,N_4999);
or UO_510 (O_510,N_4519,N_4361);
nand UO_511 (O_511,N_4155,N_4044);
nor UO_512 (O_512,N_4033,N_4419);
nor UO_513 (O_513,N_4143,N_4752);
nand UO_514 (O_514,N_4670,N_4027);
nor UO_515 (O_515,N_4880,N_4972);
or UO_516 (O_516,N_4360,N_4172);
nor UO_517 (O_517,N_4028,N_4838);
or UO_518 (O_518,N_4946,N_4559);
xnor UO_519 (O_519,N_4948,N_4845);
and UO_520 (O_520,N_4920,N_4262);
xnor UO_521 (O_521,N_4350,N_4060);
and UO_522 (O_522,N_4568,N_4235);
and UO_523 (O_523,N_4870,N_4603);
nand UO_524 (O_524,N_4037,N_4502);
and UO_525 (O_525,N_4097,N_4256);
or UO_526 (O_526,N_4680,N_4548);
xor UO_527 (O_527,N_4348,N_4113);
or UO_528 (O_528,N_4982,N_4712);
nand UO_529 (O_529,N_4758,N_4038);
or UO_530 (O_530,N_4664,N_4399);
nor UO_531 (O_531,N_4675,N_4984);
nor UO_532 (O_532,N_4809,N_4701);
nor UO_533 (O_533,N_4499,N_4049);
and UO_534 (O_534,N_4292,N_4930);
nand UO_535 (O_535,N_4601,N_4110);
nor UO_536 (O_536,N_4609,N_4735);
and UO_537 (O_537,N_4150,N_4194);
nor UO_538 (O_538,N_4044,N_4768);
nor UO_539 (O_539,N_4655,N_4117);
or UO_540 (O_540,N_4048,N_4950);
nand UO_541 (O_541,N_4865,N_4895);
nor UO_542 (O_542,N_4841,N_4348);
and UO_543 (O_543,N_4876,N_4926);
nand UO_544 (O_544,N_4957,N_4325);
nor UO_545 (O_545,N_4042,N_4850);
nand UO_546 (O_546,N_4495,N_4801);
nand UO_547 (O_547,N_4204,N_4997);
nand UO_548 (O_548,N_4955,N_4031);
or UO_549 (O_549,N_4890,N_4609);
and UO_550 (O_550,N_4670,N_4521);
xnor UO_551 (O_551,N_4774,N_4223);
nor UO_552 (O_552,N_4210,N_4886);
or UO_553 (O_553,N_4495,N_4024);
nor UO_554 (O_554,N_4942,N_4972);
or UO_555 (O_555,N_4899,N_4275);
nand UO_556 (O_556,N_4884,N_4139);
and UO_557 (O_557,N_4777,N_4186);
and UO_558 (O_558,N_4172,N_4613);
nand UO_559 (O_559,N_4688,N_4130);
nor UO_560 (O_560,N_4100,N_4822);
nor UO_561 (O_561,N_4323,N_4727);
or UO_562 (O_562,N_4127,N_4017);
nand UO_563 (O_563,N_4749,N_4750);
nor UO_564 (O_564,N_4523,N_4003);
nand UO_565 (O_565,N_4897,N_4303);
xor UO_566 (O_566,N_4152,N_4690);
and UO_567 (O_567,N_4297,N_4322);
or UO_568 (O_568,N_4294,N_4042);
nand UO_569 (O_569,N_4088,N_4412);
nand UO_570 (O_570,N_4942,N_4786);
nand UO_571 (O_571,N_4386,N_4964);
or UO_572 (O_572,N_4700,N_4365);
or UO_573 (O_573,N_4615,N_4304);
xnor UO_574 (O_574,N_4327,N_4496);
or UO_575 (O_575,N_4183,N_4812);
nand UO_576 (O_576,N_4255,N_4205);
and UO_577 (O_577,N_4558,N_4884);
nand UO_578 (O_578,N_4988,N_4980);
nand UO_579 (O_579,N_4168,N_4354);
or UO_580 (O_580,N_4850,N_4649);
or UO_581 (O_581,N_4675,N_4706);
and UO_582 (O_582,N_4745,N_4377);
xnor UO_583 (O_583,N_4183,N_4323);
xor UO_584 (O_584,N_4588,N_4303);
nor UO_585 (O_585,N_4397,N_4383);
nand UO_586 (O_586,N_4048,N_4072);
or UO_587 (O_587,N_4097,N_4286);
nor UO_588 (O_588,N_4560,N_4506);
nor UO_589 (O_589,N_4009,N_4089);
or UO_590 (O_590,N_4467,N_4199);
or UO_591 (O_591,N_4080,N_4768);
nand UO_592 (O_592,N_4596,N_4169);
xor UO_593 (O_593,N_4832,N_4217);
xor UO_594 (O_594,N_4793,N_4144);
and UO_595 (O_595,N_4404,N_4355);
and UO_596 (O_596,N_4499,N_4292);
and UO_597 (O_597,N_4022,N_4331);
nor UO_598 (O_598,N_4680,N_4964);
nor UO_599 (O_599,N_4833,N_4954);
xnor UO_600 (O_600,N_4497,N_4505);
or UO_601 (O_601,N_4639,N_4520);
xnor UO_602 (O_602,N_4240,N_4695);
or UO_603 (O_603,N_4793,N_4835);
or UO_604 (O_604,N_4479,N_4888);
or UO_605 (O_605,N_4068,N_4582);
nor UO_606 (O_606,N_4706,N_4062);
and UO_607 (O_607,N_4746,N_4936);
nor UO_608 (O_608,N_4162,N_4425);
and UO_609 (O_609,N_4474,N_4833);
nand UO_610 (O_610,N_4891,N_4000);
xor UO_611 (O_611,N_4596,N_4520);
and UO_612 (O_612,N_4916,N_4626);
nand UO_613 (O_613,N_4964,N_4841);
nor UO_614 (O_614,N_4128,N_4613);
and UO_615 (O_615,N_4755,N_4061);
and UO_616 (O_616,N_4052,N_4676);
or UO_617 (O_617,N_4236,N_4881);
or UO_618 (O_618,N_4520,N_4628);
nand UO_619 (O_619,N_4415,N_4324);
and UO_620 (O_620,N_4510,N_4741);
or UO_621 (O_621,N_4743,N_4205);
or UO_622 (O_622,N_4730,N_4996);
nand UO_623 (O_623,N_4462,N_4905);
nand UO_624 (O_624,N_4436,N_4045);
nor UO_625 (O_625,N_4530,N_4932);
xor UO_626 (O_626,N_4477,N_4965);
xnor UO_627 (O_627,N_4182,N_4733);
and UO_628 (O_628,N_4254,N_4321);
and UO_629 (O_629,N_4023,N_4358);
and UO_630 (O_630,N_4552,N_4053);
and UO_631 (O_631,N_4202,N_4073);
nand UO_632 (O_632,N_4215,N_4728);
nor UO_633 (O_633,N_4699,N_4103);
nor UO_634 (O_634,N_4448,N_4140);
nor UO_635 (O_635,N_4004,N_4461);
and UO_636 (O_636,N_4371,N_4292);
or UO_637 (O_637,N_4301,N_4813);
or UO_638 (O_638,N_4875,N_4262);
xnor UO_639 (O_639,N_4597,N_4590);
nor UO_640 (O_640,N_4290,N_4324);
nor UO_641 (O_641,N_4471,N_4188);
or UO_642 (O_642,N_4541,N_4461);
and UO_643 (O_643,N_4331,N_4031);
or UO_644 (O_644,N_4095,N_4818);
nand UO_645 (O_645,N_4991,N_4312);
nor UO_646 (O_646,N_4632,N_4530);
nand UO_647 (O_647,N_4204,N_4999);
or UO_648 (O_648,N_4199,N_4983);
and UO_649 (O_649,N_4492,N_4372);
nor UO_650 (O_650,N_4176,N_4830);
or UO_651 (O_651,N_4564,N_4964);
nand UO_652 (O_652,N_4483,N_4960);
or UO_653 (O_653,N_4620,N_4432);
xor UO_654 (O_654,N_4836,N_4039);
or UO_655 (O_655,N_4253,N_4545);
or UO_656 (O_656,N_4877,N_4886);
and UO_657 (O_657,N_4846,N_4821);
nand UO_658 (O_658,N_4215,N_4821);
and UO_659 (O_659,N_4936,N_4818);
and UO_660 (O_660,N_4622,N_4925);
nor UO_661 (O_661,N_4587,N_4543);
nor UO_662 (O_662,N_4728,N_4691);
nor UO_663 (O_663,N_4965,N_4104);
nor UO_664 (O_664,N_4260,N_4498);
xor UO_665 (O_665,N_4316,N_4019);
and UO_666 (O_666,N_4016,N_4865);
and UO_667 (O_667,N_4882,N_4834);
xor UO_668 (O_668,N_4770,N_4216);
nand UO_669 (O_669,N_4716,N_4183);
and UO_670 (O_670,N_4544,N_4454);
nand UO_671 (O_671,N_4266,N_4507);
and UO_672 (O_672,N_4554,N_4247);
xor UO_673 (O_673,N_4895,N_4690);
nor UO_674 (O_674,N_4842,N_4720);
and UO_675 (O_675,N_4027,N_4845);
and UO_676 (O_676,N_4360,N_4442);
nor UO_677 (O_677,N_4806,N_4447);
nand UO_678 (O_678,N_4091,N_4451);
and UO_679 (O_679,N_4474,N_4830);
nor UO_680 (O_680,N_4934,N_4387);
or UO_681 (O_681,N_4662,N_4150);
or UO_682 (O_682,N_4911,N_4293);
nand UO_683 (O_683,N_4933,N_4445);
or UO_684 (O_684,N_4347,N_4578);
xnor UO_685 (O_685,N_4587,N_4663);
and UO_686 (O_686,N_4864,N_4504);
xor UO_687 (O_687,N_4839,N_4286);
or UO_688 (O_688,N_4463,N_4435);
nand UO_689 (O_689,N_4374,N_4503);
nor UO_690 (O_690,N_4313,N_4839);
nand UO_691 (O_691,N_4400,N_4079);
and UO_692 (O_692,N_4873,N_4153);
or UO_693 (O_693,N_4672,N_4812);
and UO_694 (O_694,N_4005,N_4728);
nor UO_695 (O_695,N_4695,N_4068);
and UO_696 (O_696,N_4182,N_4377);
nand UO_697 (O_697,N_4069,N_4922);
and UO_698 (O_698,N_4546,N_4782);
nand UO_699 (O_699,N_4839,N_4883);
nor UO_700 (O_700,N_4353,N_4084);
nor UO_701 (O_701,N_4419,N_4518);
nor UO_702 (O_702,N_4655,N_4758);
nor UO_703 (O_703,N_4111,N_4899);
and UO_704 (O_704,N_4164,N_4690);
nand UO_705 (O_705,N_4110,N_4744);
nor UO_706 (O_706,N_4405,N_4783);
and UO_707 (O_707,N_4376,N_4247);
or UO_708 (O_708,N_4212,N_4933);
or UO_709 (O_709,N_4082,N_4737);
or UO_710 (O_710,N_4389,N_4442);
xor UO_711 (O_711,N_4103,N_4624);
or UO_712 (O_712,N_4641,N_4070);
nor UO_713 (O_713,N_4967,N_4803);
and UO_714 (O_714,N_4789,N_4211);
nor UO_715 (O_715,N_4888,N_4372);
or UO_716 (O_716,N_4823,N_4095);
and UO_717 (O_717,N_4854,N_4747);
nand UO_718 (O_718,N_4283,N_4120);
nor UO_719 (O_719,N_4275,N_4464);
nor UO_720 (O_720,N_4500,N_4763);
nand UO_721 (O_721,N_4208,N_4288);
and UO_722 (O_722,N_4775,N_4141);
xor UO_723 (O_723,N_4938,N_4105);
nand UO_724 (O_724,N_4327,N_4392);
nand UO_725 (O_725,N_4977,N_4782);
nor UO_726 (O_726,N_4014,N_4611);
and UO_727 (O_727,N_4516,N_4601);
and UO_728 (O_728,N_4791,N_4575);
or UO_729 (O_729,N_4416,N_4060);
or UO_730 (O_730,N_4690,N_4641);
nor UO_731 (O_731,N_4760,N_4209);
nand UO_732 (O_732,N_4192,N_4397);
nor UO_733 (O_733,N_4740,N_4222);
or UO_734 (O_734,N_4460,N_4472);
nor UO_735 (O_735,N_4075,N_4216);
or UO_736 (O_736,N_4778,N_4114);
or UO_737 (O_737,N_4045,N_4047);
nand UO_738 (O_738,N_4048,N_4496);
and UO_739 (O_739,N_4856,N_4849);
or UO_740 (O_740,N_4554,N_4631);
nor UO_741 (O_741,N_4931,N_4981);
or UO_742 (O_742,N_4619,N_4702);
or UO_743 (O_743,N_4869,N_4737);
or UO_744 (O_744,N_4081,N_4371);
and UO_745 (O_745,N_4584,N_4709);
nor UO_746 (O_746,N_4632,N_4882);
nand UO_747 (O_747,N_4293,N_4930);
nand UO_748 (O_748,N_4565,N_4182);
nand UO_749 (O_749,N_4975,N_4234);
and UO_750 (O_750,N_4958,N_4083);
nand UO_751 (O_751,N_4286,N_4163);
nor UO_752 (O_752,N_4736,N_4432);
or UO_753 (O_753,N_4401,N_4925);
nand UO_754 (O_754,N_4711,N_4716);
or UO_755 (O_755,N_4512,N_4783);
nor UO_756 (O_756,N_4407,N_4915);
nor UO_757 (O_757,N_4575,N_4901);
nand UO_758 (O_758,N_4044,N_4421);
and UO_759 (O_759,N_4067,N_4047);
xor UO_760 (O_760,N_4167,N_4483);
nor UO_761 (O_761,N_4227,N_4326);
xnor UO_762 (O_762,N_4768,N_4991);
nor UO_763 (O_763,N_4933,N_4938);
and UO_764 (O_764,N_4581,N_4557);
nand UO_765 (O_765,N_4468,N_4515);
nor UO_766 (O_766,N_4339,N_4258);
and UO_767 (O_767,N_4208,N_4137);
and UO_768 (O_768,N_4955,N_4763);
nor UO_769 (O_769,N_4328,N_4035);
nor UO_770 (O_770,N_4360,N_4647);
nand UO_771 (O_771,N_4679,N_4153);
nor UO_772 (O_772,N_4786,N_4559);
nand UO_773 (O_773,N_4348,N_4000);
xor UO_774 (O_774,N_4220,N_4730);
nor UO_775 (O_775,N_4529,N_4869);
and UO_776 (O_776,N_4642,N_4659);
nand UO_777 (O_777,N_4767,N_4150);
nand UO_778 (O_778,N_4708,N_4654);
nand UO_779 (O_779,N_4944,N_4629);
and UO_780 (O_780,N_4783,N_4138);
xnor UO_781 (O_781,N_4040,N_4174);
and UO_782 (O_782,N_4359,N_4667);
and UO_783 (O_783,N_4465,N_4193);
nand UO_784 (O_784,N_4240,N_4707);
nor UO_785 (O_785,N_4165,N_4648);
and UO_786 (O_786,N_4360,N_4895);
or UO_787 (O_787,N_4906,N_4251);
and UO_788 (O_788,N_4261,N_4911);
nor UO_789 (O_789,N_4208,N_4226);
xor UO_790 (O_790,N_4214,N_4804);
or UO_791 (O_791,N_4692,N_4058);
nor UO_792 (O_792,N_4194,N_4393);
or UO_793 (O_793,N_4341,N_4380);
or UO_794 (O_794,N_4540,N_4112);
and UO_795 (O_795,N_4897,N_4938);
nand UO_796 (O_796,N_4981,N_4204);
and UO_797 (O_797,N_4830,N_4471);
nand UO_798 (O_798,N_4277,N_4958);
and UO_799 (O_799,N_4219,N_4474);
nand UO_800 (O_800,N_4696,N_4964);
nand UO_801 (O_801,N_4704,N_4070);
and UO_802 (O_802,N_4798,N_4998);
xnor UO_803 (O_803,N_4950,N_4432);
nand UO_804 (O_804,N_4746,N_4462);
nand UO_805 (O_805,N_4835,N_4415);
nor UO_806 (O_806,N_4616,N_4418);
and UO_807 (O_807,N_4631,N_4822);
xnor UO_808 (O_808,N_4033,N_4017);
or UO_809 (O_809,N_4487,N_4086);
nand UO_810 (O_810,N_4609,N_4467);
xor UO_811 (O_811,N_4440,N_4285);
nand UO_812 (O_812,N_4307,N_4854);
xor UO_813 (O_813,N_4777,N_4975);
nand UO_814 (O_814,N_4791,N_4934);
or UO_815 (O_815,N_4164,N_4552);
and UO_816 (O_816,N_4419,N_4098);
nand UO_817 (O_817,N_4800,N_4892);
and UO_818 (O_818,N_4537,N_4380);
nor UO_819 (O_819,N_4305,N_4608);
and UO_820 (O_820,N_4305,N_4946);
nand UO_821 (O_821,N_4624,N_4767);
or UO_822 (O_822,N_4045,N_4012);
nor UO_823 (O_823,N_4252,N_4685);
nand UO_824 (O_824,N_4784,N_4102);
or UO_825 (O_825,N_4231,N_4291);
nand UO_826 (O_826,N_4757,N_4990);
or UO_827 (O_827,N_4469,N_4401);
nand UO_828 (O_828,N_4641,N_4678);
nor UO_829 (O_829,N_4356,N_4380);
xnor UO_830 (O_830,N_4801,N_4435);
nand UO_831 (O_831,N_4322,N_4278);
nor UO_832 (O_832,N_4723,N_4843);
and UO_833 (O_833,N_4434,N_4976);
nand UO_834 (O_834,N_4433,N_4420);
nor UO_835 (O_835,N_4600,N_4395);
and UO_836 (O_836,N_4625,N_4064);
xnor UO_837 (O_837,N_4940,N_4640);
or UO_838 (O_838,N_4299,N_4972);
nand UO_839 (O_839,N_4301,N_4154);
nor UO_840 (O_840,N_4912,N_4591);
nand UO_841 (O_841,N_4018,N_4535);
and UO_842 (O_842,N_4999,N_4447);
nand UO_843 (O_843,N_4387,N_4743);
and UO_844 (O_844,N_4254,N_4549);
and UO_845 (O_845,N_4442,N_4986);
nor UO_846 (O_846,N_4758,N_4062);
and UO_847 (O_847,N_4814,N_4354);
and UO_848 (O_848,N_4418,N_4941);
xnor UO_849 (O_849,N_4483,N_4623);
or UO_850 (O_850,N_4935,N_4831);
nor UO_851 (O_851,N_4677,N_4863);
nor UO_852 (O_852,N_4692,N_4909);
xor UO_853 (O_853,N_4513,N_4556);
nor UO_854 (O_854,N_4041,N_4202);
nand UO_855 (O_855,N_4488,N_4957);
and UO_856 (O_856,N_4222,N_4283);
or UO_857 (O_857,N_4782,N_4273);
nand UO_858 (O_858,N_4283,N_4676);
or UO_859 (O_859,N_4809,N_4383);
nand UO_860 (O_860,N_4627,N_4777);
and UO_861 (O_861,N_4083,N_4652);
and UO_862 (O_862,N_4746,N_4301);
nor UO_863 (O_863,N_4201,N_4277);
nor UO_864 (O_864,N_4371,N_4435);
nand UO_865 (O_865,N_4273,N_4583);
nor UO_866 (O_866,N_4069,N_4717);
and UO_867 (O_867,N_4830,N_4390);
or UO_868 (O_868,N_4724,N_4271);
and UO_869 (O_869,N_4386,N_4044);
nor UO_870 (O_870,N_4317,N_4916);
or UO_871 (O_871,N_4205,N_4075);
nand UO_872 (O_872,N_4045,N_4989);
and UO_873 (O_873,N_4302,N_4119);
xor UO_874 (O_874,N_4709,N_4642);
nand UO_875 (O_875,N_4694,N_4871);
nand UO_876 (O_876,N_4963,N_4012);
or UO_877 (O_877,N_4304,N_4065);
nor UO_878 (O_878,N_4595,N_4072);
or UO_879 (O_879,N_4330,N_4441);
xnor UO_880 (O_880,N_4210,N_4697);
nor UO_881 (O_881,N_4707,N_4122);
and UO_882 (O_882,N_4363,N_4542);
nor UO_883 (O_883,N_4735,N_4401);
nand UO_884 (O_884,N_4952,N_4022);
or UO_885 (O_885,N_4810,N_4054);
nor UO_886 (O_886,N_4992,N_4731);
and UO_887 (O_887,N_4478,N_4632);
and UO_888 (O_888,N_4505,N_4648);
or UO_889 (O_889,N_4023,N_4481);
and UO_890 (O_890,N_4716,N_4723);
and UO_891 (O_891,N_4338,N_4692);
or UO_892 (O_892,N_4779,N_4980);
nand UO_893 (O_893,N_4901,N_4395);
nand UO_894 (O_894,N_4208,N_4123);
or UO_895 (O_895,N_4553,N_4035);
nor UO_896 (O_896,N_4473,N_4904);
or UO_897 (O_897,N_4783,N_4364);
and UO_898 (O_898,N_4942,N_4290);
and UO_899 (O_899,N_4993,N_4491);
nand UO_900 (O_900,N_4643,N_4471);
and UO_901 (O_901,N_4767,N_4187);
or UO_902 (O_902,N_4377,N_4415);
nand UO_903 (O_903,N_4928,N_4446);
nand UO_904 (O_904,N_4019,N_4540);
nand UO_905 (O_905,N_4743,N_4165);
xnor UO_906 (O_906,N_4455,N_4618);
nor UO_907 (O_907,N_4761,N_4696);
or UO_908 (O_908,N_4016,N_4534);
and UO_909 (O_909,N_4767,N_4925);
or UO_910 (O_910,N_4763,N_4707);
nor UO_911 (O_911,N_4718,N_4487);
or UO_912 (O_912,N_4161,N_4615);
nor UO_913 (O_913,N_4344,N_4023);
or UO_914 (O_914,N_4582,N_4388);
or UO_915 (O_915,N_4425,N_4220);
and UO_916 (O_916,N_4593,N_4600);
and UO_917 (O_917,N_4574,N_4474);
and UO_918 (O_918,N_4873,N_4052);
nor UO_919 (O_919,N_4280,N_4660);
nor UO_920 (O_920,N_4241,N_4886);
nor UO_921 (O_921,N_4227,N_4782);
nand UO_922 (O_922,N_4540,N_4221);
nand UO_923 (O_923,N_4816,N_4340);
xor UO_924 (O_924,N_4592,N_4705);
nand UO_925 (O_925,N_4738,N_4286);
xor UO_926 (O_926,N_4383,N_4498);
nand UO_927 (O_927,N_4155,N_4147);
and UO_928 (O_928,N_4291,N_4572);
xnor UO_929 (O_929,N_4895,N_4635);
xor UO_930 (O_930,N_4811,N_4683);
nand UO_931 (O_931,N_4701,N_4524);
nor UO_932 (O_932,N_4983,N_4504);
or UO_933 (O_933,N_4339,N_4657);
and UO_934 (O_934,N_4436,N_4504);
or UO_935 (O_935,N_4764,N_4486);
nor UO_936 (O_936,N_4296,N_4620);
nand UO_937 (O_937,N_4439,N_4013);
nor UO_938 (O_938,N_4431,N_4394);
xnor UO_939 (O_939,N_4148,N_4950);
nand UO_940 (O_940,N_4271,N_4154);
or UO_941 (O_941,N_4937,N_4250);
nor UO_942 (O_942,N_4381,N_4024);
nor UO_943 (O_943,N_4386,N_4899);
nand UO_944 (O_944,N_4565,N_4766);
xor UO_945 (O_945,N_4336,N_4231);
nand UO_946 (O_946,N_4868,N_4738);
nand UO_947 (O_947,N_4096,N_4376);
nand UO_948 (O_948,N_4814,N_4582);
nand UO_949 (O_949,N_4519,N_4134);
or UO_950 (O_950,N_4903,N_4104);
xor UO_951 (O_951,N_4725,N_4121);
xor UO_952 (O_952,N_4626,N_4694);
and UO_953 (O_953,N_4422,N_4250);
or UO_954 (O_954,N_4742,N_4096);
nor UO_955 (O_955,N_4070,N_4783);
or UO_956 (O_956,N_4478,N_4625);
and UO_957 (O_957,N_4867,N_4066);
or UO_958 (O_958,N_4567,N_4412);
or UO_959 (O_959,N_4237,N_4798);
and UO_960 (O_960,N_4084,N_4164);
nand UO_961 (O_961,N_4856,N_4669);
and UO_962 (O_962,N_4693,N_4522);
and UO_963 (O_963,N_4581,N_4996);
and UO_964 (O_964,N_4518,N_4014);
nand UO_965 (O_965,N_4386,N_4836);
nor UO_966 (O_966,N_4638,N_4931);
and UO_967 (O_967,N_4923,N_4731);
nor UO_968 (O_968,N_4084,N_4381);
nor UO_969 (O_969,N_4912,N_4887);
nor UO_970 (O_970,N_4452,N_4767);
or UO_971 (O_971,N_4050,N_4074);
or UO_972 (O_972,N_4030,N_4385);
xor UO_973 (O_973,N_4664,N_4188);
and UO_974 (O_974,N_4280,N_4301);
and UO_975 (O_975,N_4455,N_4897);
and UO_976 (O_976,N_4204,N_4457);
nand UO_977 (O_977,N_4171,N_4414);
or UO_978 (O_978,N_4855,N_4642);
or UO_979 (O_979,N_4628,N_4046);
nand UO_980 (O_980,N_4225,N_4197);
and UO_981 (O_981,N_4035,N_4881);
or UO_982 (O_982,N_4804,N_4046);
or UO_983 (O_983,N_4522,N_4379);
nor UO_984 (O_984,N_4081,N_4219);
nor UO_985 (O_985,N_4155,N_4935);
nand UO_986 (O_986,N_4256,N_4269);
and UO_987 (O_987,N_4416,N_4029);
nand UO_988 (O_988,N_4017,N_4849);
nand UO_989 (O_989,N_4159,N_4560);
and UO_990 (O_990,N_4674,N_4174);
or UO_991 (O_991,N_4658,N_4407);
and UO_992 (O_992,N_4091,N_4719);
nor UO_993 (O_993,N_4545,N_4223);
nand UO_994 (O_994,N_4184,N_4984);
nor UO_995 (O_995,N_4570,N_4150);
or UO_996 (O_996,N_4016,N_4267);
xor UO_997 (O_997,N_4264,N_4295);
nand UO_998 (O_998,N_4677,N_4460);
or UO_999 (O_999,N_4533,N_4390);
endmodule