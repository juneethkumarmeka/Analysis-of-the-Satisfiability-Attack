module basic_1000_10000_1500_2_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5009,N_5010,N_5011,N_5012,N_5015,N_5016,N_5017,N_5018,N_5019,N_5021,N_5023,N_5024,N_5028,N_5029,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5039,N_5040,N_5043,N_5045,N_5048,N_5050,N_5051,N_5052,N_5053,N_5055,N_5061,N_5062,N_5064,N_5068,N_5069,N_5070,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5082,N_5084,N_5087,N_5089,N_5090,N_5092,N_5093,N_5097,N_5098,N_5099,N_5101,N_5102,N_5104,N_5105,N_5107,N_5109,N_5110,N_5111,N_5112,N_5113,N_5115,N_5120,N_5121,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5130,N_5132,N_5134,N_5138,N_5139,N_5140,N_5141,N_5143,N_5144,N_5145,N_5152,N_5154,N_5155,N_5156,N_5157,N_5159,N_5161,N_5163,N_5168,N_5169,N_5170,N_5173,N_5174,N_5176,N_5177,N_5178,N_5179,N_5181,N_5182,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5194,N_5195,N_5196,N_5198,N_5202,N_5203,N_5204,N_5205,N_5207,N_5208,N_5209,N_5210,N_5211,N_5215,N_5218,N_5219,N_5220,N_5222,N_5223,N_5224,N_5225,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5236,N_5237,N_5240,N_5241,N_5242,N_5244,N_5245,N_5249,N_5250,N_5251,N_5252,N_5256,N_5257,N_5261,N_5262,N_5266,N_5267,N_5268,N_5272,N_5273,N_5274,N_5276,N_5280,N_5281,N_5286,N_5288,N_5290,N_5295,N_5296,N_5298,N_5299,N_5300,N_5301,N_5304,N_5306,N_5309,N_5310,N_5311,N_5312,N_5314,N_5315,N_5316,N_5317,N_5319,N_5320,N_5322,N_5324,N_5325,N_5326,N_5329,N_5332,N_5334,N_5335,N_5336,N_5338,N_5341,N_5342,N_5343,N_5346,N_5348,N_5351,N_5352,N_5353,N_5354,N_5355,N_5360,N_5362,N_5364,N_5365,N_5366,N_5367,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5390,N_5391,N_5394,N_5396,N_5398,N_5399,N_5401,N_5402,N_5405,N_5406,N_5408,N_5409,N_5412,N_5413,N_5414,N_5416,N_5417,N_5419,N_5421,N_5422,N_5424,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5443,N_5444,N_5445,N_5446,N_5447,N_5450,N_5453,N_5456,N_5457,N_5459,N_5460,N_5468,N_5470,N_5471,N_5474,N_5476,N_5477,N_5478,N_5479,N_5480,N_5482,N_5484,N_5486,N_5488,N_5489,N_5491,N_5492,N_5493,N_5495,N_5496,N_5497,N_5501,N_5503,N_5504,N_5505,N_5507,N_5508,N_5509,N_5510,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5519,N_5520,N_5521,N_5522,N_5523,N_5525,N_5526,N_5528,N_5529,N_5532,N_5534,N_5535,N_5536,N_5537,N_5538,N_5540,N_5542,N_5543,N_5544,N_5546,N_5547,N_5548,N_5549,N_5551,N_5554,N_5555,N_5557,N_5558,N_5559,N_5561,N_5564,N_5565,N_5567,N_5568,N_5570,N_5571,N_5572,N_5575,N_5576,N_5579,N_5580,N_5581,N_5582,N_5585,N_5586,N_5587,N_5589,N_5590,N_5592,N_5593,N_5594,N_5595,N_5600,N_5603,N_5606,N_5607,N_5608,N_5610,N_5612,N_5614,N_5616,N_5618,N_5619,N_5621,N_5622,N_5623,N_5625,N_5626,N_5627,N_5629,N_5631,N_5634,N_5635,N_5639,N_5641,N_5642,N_5643,N_5648,N_5649,N_5651,N_5653,N_5654,N_5656,N_5657,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5668,N_5670,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5681,N_5682,N_5684,N_5686,N_5687,N_5688,N_5689,N_5691,N_5692,N_5694,N_5697,N_5698,N_5699,N_5701,N_5702,N_5703,N_5707,N_5711,N_5712,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5721,N_5723,N_5724,N_5725,N_5729,N_5730,N_5731,N_5733,N_5734,N_5735,N_5736,N_5738,N_5740,N_5741,N_5743,N_5750,N_5751,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5762,N_5763,N_5765,N_5766,N_5767,N_5769,N_5771,N_5772,N_5774,N_5775,N_5777,N_5778,N_5780,N_5781,N_5782,N_5784,N_5785,N_5789,N_5790,N_5793,N_5796,N_5797,N_5799,N_5800,N_5802,N_5804,N_5805,N_5810,N_5811,N_5814,N_5816,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5825,N_5828,N_5829,N_5832,N_5833,N_5834,N_5837,N_5838,N_5840,N_5844,N_5845,N_5846,N_5848,N_5850,N_5854,N_5855,N_5856,N_5858,N_5859,N_5865,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5876,N_5877,N_5879,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5892,N_5893,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5903,N_5904,N_5909,N_5910,N_5911,N_5913,N_5917,N_5918,N_5919,N_5920,N_5921,N_5923,N_5924,N_5925,N_5926,N_5928,N_5929,N_5931,N_5933,N_5935,N_5938,N_5939,N_5942,N_5944,N_5946,N_5949,N_5952,N_5954,N_5955,N_5959,N_5960,N_5961,N_5962,N_5966,N_5967,N_5968,N_5970,N_5971,N_5973,N_5974,N_5975,N_5977,N_5978,N_5979,N_5980,N_5982,N_5983,N_5984,N_5986,N_5987,N_5988,N_5995,N_5996,N_5997,N_5999,N_6002,N_6003,N_6004,N_6006,N_6007,N_6009,N_6012,N_6013,N_6015,N_6019,N_6021,N_6022,N_6023,N_6024,N_6027,N_6030,N_6031,N_6032,N_6035,N_6037,N_6038,N_6039,N_6040,N_6041,N_6043,N_6044,N_6047,N_6048,N_6050,N_6051,N_6053,N_6056,N_6061,N_6064,N_6066,N_6067,N_6068,N_6070,N_6073,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6087,N_6088,N_6091,N_6093,N_6094,N_6095,N_6098,N_6099,N_6101,N_6103,N_6106,N_6110,N_6112,N_6113,N_6114,N_6115,N_6119,N_6120,N_6121,N_6122,N_6124,N_6125,N_6126,N_6127,N_6129,N_6130,N_6133,N_6136,N_6138,N_6139,N_6140,N_6142,N_6144,N_6145,N_6146,N_6148,N_6151,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6162,N_6164,N_6167,N_6169,N_6170,N_6171,N_6174,N_6175,N_6177,N_6179,N_6180,N_6181,N_6182,N_6185,N_6186,N_6187,N_6192,N_6194,N_6195,N_6196,N_6197,N_6201,N_6202,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6212,N_6214,N_6216,N_6219,N_6222,N_6223,N_6225,N_6226,N_6229,N_6230,N_6231,N_6232,N_6235,N_6236,N_6237,N_6241,N_6242,N_6243,N_6244,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6257,N_6265,N_6268,N_6269,N_6270,N_6272,N_6274,N_6276,N_6278,N_6279,N_6280,N_6281,N_6282,N_6285,N_6287,N_6288,N_6289,N_6293,N_6294,N_6295,N_6296,N_6297,N_6299,N_6303,N_6304,N_6305,N_6307,N_6313,N_6314,N_6315,N_6321,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6342,N_6343,N_6344,N_6346,N_6350,N_6351,N_6353,N_6355,N_6356,N_6357,N_6358,N_6360,N_6361,N_6362,N_6366,N_6367,N_6368,N_6371,N_6372,N_6373,N_6375,N_6377,N_6379,N_6381,N_6384,N_6385,N_6386,N_6387,N_6389,N_6390,N_6392,N_6393,N_6394,N_6395,N_6396,N_6398,N_6399,N_6400,N_6402,N_6405,N_6408,N_6409,N_6412,N_6414,N_6416,N_6418,N_6419,N_6420,N_6425,N_6430,N_6431,N_6433,N_6434,N_6435,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6449,N_6451,N_6452,N_6454,N_6455,N_6459,N_6462,N_6464,N_6465,N_6466,N_6469,N_6470,N_6472,N_6473,N_6477,N_6480,N_6481,N_6482,N_6484,N_6485,N_6487,N_6488,N_6489,N_6490,N_6492,N_6493,N_6494,N_6495,N_6497,N_6498,N_6499,N_6500,N_6503,N_6505,N_6506,N_6507,N_6511,N_6512,N_6514,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6530,N_6531,N_6532,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6541,N_6543,N_6544,N_6546,N_6548,N_6550,N_6552,N_6553,N_6554,N_6555,N_6557,N_6558,N_6560,N_6561,N_6562,N_6564,N_6565,N_6566,N_6567,N_6568,N_6570,N_6571,N_6572,N_6575,N_6577,N_6578,N_6584,N_6585,N_6586,N_6588,N_6589,N_6591,N_6592,N_6595,N_6596,N_6598,N_6601,N_6602,N_6604,N_6606,N_6607,N_6609,N_6611,N_6612,N_6613,N_6614,N_6617,N_6618,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6631,N_6634,N_6635,N_6638,N_6640,N_6641,N_6645,N_6646,N_6647,N_6655,N_6656,N_6657,N_6659,N_6664,N_6666,N_6667,N_6668,N_6670,N_6672,N_6674,N_6675,N_6677,N_6679,N_6681,N_6682,N_6684,N_6685,N_6687,N_6689,N_6690,N_6691,N_6692,N_6693,N_6696,N_6697,N_6698,N_6699,N_6701,N_6703,N_6704,N_6706,N_6709,N_6710,N_6711,N_6713,N_6714,N_6716,N_6717,N_6718,N_6720,N_6722,N_6723,N_6725,N_6726,N_6727,N_6728,N_6733,N_6734,N_6735,N_6736,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6752,N_6753,N_6754,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6768,N_6769,N_6771,N_6772,N_6773,N_6774,N_6778,N_6779,N_6784,N_6785,N_6789,N_6791,N_6792,N_6794,N_6795,N_6796,N_6797,N_6799,N_6801,N_6803,N_6804,N_6806,N_6808,N_6809,N_6810,N_6811,N_6813,N_6814,N_6821,N_6824,N_6825,N_6826,N_6827,N_6828,N_6831,N_6834,N_6835,N_6838,N_6840,N_6842,N_6843,N_6845,N_6849,N_6850,N_6851,N_6856,N_6857,N_6860,N_6862,N_6863,N_6864,N_6865,N_6867,N_6868,N_6870,N_6871,N_6873,N_6874,N_6876,N_6877,N_6879,N_6880,N_6882,N_6885,N_6886,N_6887,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6898,N_6899,N_6901,N_6902,N_6903,N_6904,N_6905,N_6907,N_6908,N_6909,N_6910,N_6912,N_6913,N_6914,N_6916,N_6918,N_6919,N_6920,N_6921,N_6925,N_6926,N_6927,N_6928,N_6929,N_6931,N_6932,N_6933,N_6934,N_6935,N_6937,N_6938,N_6939,N_6940,N_6941,N_6943,N_6945,N_6946,N_6947,N_6948,N_6949,N_6951,N_6952,N_6953,N_6954,N_6958,N_6959,N_6960,N_6961,N_6964,N_6966,N_6968,N_6971,N_6973,N_6974,N_6977,N_6978,N_6980,N_6982,N_6984,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6995,N_6997,N_6998,N_6999,N_7000,N_7001,N_7003,N_7005,N_7007,N_7008,N_7009,N_7011,N_7019,N_7020,N_7022,N_7025,N_7026,N_7027,N_7029,N_7030,N_7031,N_7032,N_7034,N_7036,N_7037,N_7040,N_7041,N_7042,N_7043,N_7045,N_7046,N_7050,N_7055,N_7059,N_7060,N_7061,N_7062,N_7064,N_7065,N_7073,N_7074,N_7075,N_7077,N_7078,N_7080,N_7081,N_7083,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7108,N_7109,N_7110,N_7112,N_7113,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7122,N_7124,N_7126,N_7127,N_7129,N_7133,N_7135,N_7136,N_7137,N_7138,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7149,N_7153,N_7157,N_7158,N_7159,N_7160,N_7162,N_7164,N_7165,N_7167,N_7172,N_7175,N_7176,N_7178,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7189,N_7190,N_7191,N_7193,N_7194,N_7195,N_7197,N_7198,N_7200,N_7202,N_7203,N_7205,N_7206,N_7207,N_7208,N_7209,N_7212,N_7213,N_7218,N_7220,N_7221,N_7224,N_7225,N_7226,N_7232,N_7235,N_7236,N_7237,N_7238,N_7239,N_7242,N_7245,N_7247,N_7249,N_7250,N_7251,N_7253,N_7254,N_7255,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7267,N_7268,N_7269,N_7270,N_7272,N_7274,N_7276,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7291,N_7292,N_7294,N_7295,N_7297,N_7299,N_7300,N_7301,N_7302,N_7303,N_7306,N_7308,N_7309,N_7311,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7320,N_7322,N_7323,N_7325,N_7326,N_7327,N_7328,N_7330,N_7336,N_7338,N_7339,N_7341,N_7342,N_7343,N_7344,N_7346,N_7348,N_7349,N_7351,N_7352,N_7353,N_7356,N_7357,N_7359,N_7361,N_7363,N_7364,N_7365,N_7367,N_7370,N_7373,N_7374,N_7375,N_7376,N_7377,N_7379,N_7380,N_7382,N_7384,N_7386,N_7387,N_7388,N_7391,N_7392,N_7394,N_7395,N_7397,N_7400,N_7401,N_7403,N_7404,N_7406,N_7407,N_7408,N_7410,N_7411,N_7416,N_7418,N_7420,N_7421,N_7423,N_7424,N_7425,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7435,N_7436,N_7438,N_7440,N_7446,N_7449,N_7450,N_7452,N_7453,N_7454,N_7455,N_7464,N_7466,N_7469,N_7470,N_7471,N_7473,N_7475,N_7476,N_7477,N_7478,N_7481,N_7482,N_7483,N_7485,N_7486,N_7489,N_7490,N_7491,N_7495,N_7496,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7508,N_7510,N_7512,N_7514,N_7515,N_7517,N_7518,N_7520,N_7521,N_7523,N_7524,N_7527,N_7528,N_7529,N_7530,N_7531,N_7534,N_7536,N_7538,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7548,N_7549,N_7554,N_7555,N_7557,N_7558,N_7559,N_7563,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7573,N_7574,N_7575,N_7576,N_7577,N_7580,N_7583,N_7584,N_7585,N_7587,N_7588,N_7590,N_7594,N_7596,N_7597,N_7598,N_7599,N_7600,N_7603,N_7604,N_7607,N_7608,N_7611,N_7612,N_7614,N_7615,N_7616,N_7618,N_7620,N_7622,N_7623,N_7626,N_7628,N_7629,N_7630,N_7631,N_7633,N_7635,N_7638,N_7639,N_7641,N_7642,N_7643,N_7644,N_7647,N_7649,N_7650,N_7651,N_7654,N_7655,N_7656,N_7657,N_7660,N_7661,N_7662,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7674,N_7675,N_7676,N_7678,N_7679,N_7680,N_7683,N_7684,N_7685,N_7686,N_7687,N_7689,N_7691,N_7695,N_7696,N_7697,N_7698,N_7703,N_7704,N_7706,N_7707,N_7708,N_7709,N_7710,N_7712,N_7713,N_7716,N_7717,N_7718,N_7720,N_7721,N_7722,N_7723,N_7725,N_7726,N_7728,N_7729,N_7730,N_7732,N_7733,N_7734,N_7735,N_7737,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7748,N_7750,N_7752,N_7753,N_7755,N_7756,N_7757,N_7759,N_7760,N_7761,N_7766,N_7767,N_7768,N_7769,N_7772,N_7773,N_7774,N_7776,N_7778,N_7779,N_7780,N_7783,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7794,N_7795,N_7796,N_7797,N_7801,N_7802,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7814,N_7815,N_7816,N_7817,N_7820,N_7821,N_7822,N_7823,N_7825,N_7828,N_7829,N_7834,N_7836,N_7839,N_7840,N_7843,N_7844,N_7845,N_7847,N_7852,N_7854,N_7855,N_7856,N_7857,N_7859,N_7862,N_7864,N_7869,N_7870,N_7873,N_7874,N_7876,N_7877,N_7879,N_7881,N_7882,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7891,N_7894,N_7895,N_7896,N_7900,N_7901,N_7902,N_7903,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7917,N_7919,N_7921,N_7922,N_7923,N_7924,N_7926,N_7927,N_7930,N_7933,N_7935,N_7937,N_7938,N_7940,N_7942,N_7943,N_7944,N_7946,N_7949,N_7950,N_7951,N_7952,N_7953,N_7955,N_7956,N_7957,N_7958,N_7961,N_7962,N_7963,N_7966,N_7968,N_7969,N_7971,N_7972,N_7973,N_7974,N_7975,N_7978,N_7981,N_7982,N_7985,N_7986,N_7987,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_8000,N_8002,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8016,N_8018,N_8019,N_8020,N_8024,N_8026,N_8027,N_8030,N_8032,N_8035,N_8036,N_8037,N_8038,N_8042,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8053,N_8057,N_8060,N_8062,N_8063,N_8064,N_8065,N_8069,N_8070,N_8073,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8083,N_8084,N_8086,N_8087,N_8089,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8100,N_8101,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8114,N_8116,N_8117,N_8118,N_8122,N_8123,N_8124,N_8127,N_8129,N_8132,N_8133,N_8134,N_8135,N_8137,N_8138,N_8140,N_8142,N_8144,N_8148,N_8149,N_8150,N_8151,N_8152,N_8154,N_8155,N_8157,N_8158,N_8159,N_8160,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8169,N_8171,N_8172,N_8174,N_8175,N_8176,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8191,N_8193,N_8194,N_8196,N_8197,N_8198,N_8199,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8224,N_8225,N_8226,N_8230,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8239,N_8241,N_8243,N_8244,N_8245,N_8247,N_8249,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8259,N_8260,N_8261,N_8262,N_8264,N_8266,N_8267,N_8269,N_8270,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8280,N_8283,N_8284,N_8290,N_8291,N_8292,N_8293,N_8294,N_8297,N_8299,N_8300,N_8301,N_8302,N_8303,N_8305,N_8306,N_8307,N_8312,N_8314,N_8315,N_8319,N_8320,N_8321,N_8326,N_8327,N_8329,N_8330,N_8331,N_8332,N_8333,N_8335,N_8336,N_8337,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8347,N_8348,N_8350,N_8351,N_8352,N_8354,N_8356,N_8358,N_8359,N_8360,N_8362,N_8364,N_8365,N_8366,N_8368,N_8369,N_8371,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8382,N_8383,N_8385,N_8387,N_8389,N_8390,N_8391,N_8392,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8403,N_8404,N_8409,N_8410,N_8413,N_8414,N_8415,N_8418,N_8420,N_8421,N_8423,N_8424,N_8427,N_8428,N_8431,N_8432,N_8433,N_8434,N_8437,N_8439,N_8440,N_8441,N_8442,N_8443,N_8445,N_8448,N_8451,N_8454,N_8458,N_8459,N_8460,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8474,N_8475,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8484,N_8487,N_8488,N_8489,N_8492,N_8493,N_8495,N_8498,N_8502,N_8503,N_8507,N_8508,N_8509,N_8511,N_8512,N_8513,N_8514,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8524,N_8529,N_8531,N_8532,N_8537,N_8538,N_8540,N_8541,N_8542,N_8543,N_8546,N_8547,N_8549,N_8550,N_8557,N_8558,N_8560,N_8563,N_8564,N_8566,N_8567,N_8568,N_8570,N_8571,N_8574,N_8575,N_8576,N_8577,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8594,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8603,N_8604,N_8607,N_8608,N_8609,N_8610,N_8611,N_8617,N_8622,N_8623,N_8624,N_8627,N_8628,N_8633,N_8635,N_8643,N_8644,N_8645,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8657,N_8658,N_8659,N_8660,N_8662,N_8663,N_8664,N_8667,N_8668,N_8669,N_8670,N_8673,N_8676,N_8678,N_8680,N_8681,N_8682,N_8683,N_8685,N_8687,N_8689,N_8692,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8701,N_8704,N_8707,N_8708,N_8710,N_8711,N_8713,N_8718,N_8721,N_8723,N_8725,N_8727,N_8728,N_8729,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8739,N_8741,N_8743,N_8746,N_8747,N_8749,N_8752,N_8753,N_8755,N_8756,N_8760,N_8762,N_8763,N_8764,N_8767,N_8770,N_8771,N_8774,N_8777,N_8778,N_8779,N_8780,N_8781,N_8784,N_8786,N_8789,N_8790,N_8794,N_8795,N_8796,N_8797,N_8802,N_8804,N_8805,N_8806,N_8808,N_8809,N_8811,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8821,N_8823,N_8824,N_8827,N_8829,N_8830,N_8834,N_8837,N_8839,N_8840,N_8841,N_8843,N_8846,N_8847,N_8849,N_8851,N_8853,N_8855,N_8856,N_8857,N_8860,N_8862,N_8863,N_8866,N_8868,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8879,N_8882,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8893,N_8897,N_8898,N_8904,N_8905,N_8907,N_8908,N_8910,N_8911,N_8912,N_8915,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8924,N_8927,N_8928,N_8931,N_8933,N_8936,N_8937,N_8938,N_8940,N_8941,N_8942,N_8945,N_8947,N_8948,N_8949,N_8951,N_8953,N_8954,N_8956,N_8960,N_8961,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8972,N_8973,N_8974,N_8975,N_8976,N_8987,N_8989,N_8994,N_8996,N_8997,N_9000,N_9002,N_9003,N_9005,N_9006,N_9007,N_9008,N_9009,N_9012,N_9016,N_9018,N_9019,N_9021,N_9025,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9037,N_9038,N_9039,N_9041,N_9042,N_9043,N_9045,N_9046,N_9048,N_9049,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9075,N_9076,N_9077,N_9078,N_9079,N_9081,N_9083,N_9084,N_9086,N_9087,N_9089,N_9090,N_9092,N_9093,N_9095,N_9097,N_9098,N_9100,N_9101,N_9102,N_9103,N_9105,N_9106,N_9108,N_9110,N_9111,N_9113,N_9114,N_9116,N_9117,N_9118,N_9119,N_9123,N_9125,N_9128,N_9130,N_9133,N_9134,N_9135,N_9136,N_9139,N_9140,N_9141,N_9142,N_9145,N_9146,N_9148,N_9149,N_9151,N_9152,N_9153,N_9156,N_9158,N_9161,N_9162,N_9163,N_9164,N_9166,N_9168,N_9169,N_9170,N_9172,N_9173,N_9176,N_9178,N_9180,N_9181,N_9183,N_9184,N_9186,N_9187,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9198,N_9200,N_9203,N_9204,N_9205,N_9208,N_9210,N_9211,N_9212,N_9218,N_9219,N_9221,N_9222,N_9223,N_9224,N_9225,N_9227,N_9228,N_9229,N_9230,N_9231,N_9233,N_9234,N_9236,N_9237,N_9238,N_9239,N_9241,N_9243,N_9245,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9259,N_9260,N_9261,N_9262,N_9264,N_9265,N_9266,N_9271,N_9272,N_9274,N_9276,N_9278,N_9279,N_9280,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9290,N_9291,N_9294,N_9295,N_9296,N_9300,N_9307,N_9309,N_9310,N_9312,N_9313,N_9315,N_9316,N_9318,N_9320,N_9321,N_9322,N_9323,N_9324,N_9326,N_9327,N_9328,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9338,N_9340,N_9342,N_9345,N_9347,N_9348,N_9350,N_9352,N_9353,N_9354,N_9355,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9370,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9379,N_9386,N_9393,N_9394,N_9395,N_9399,N_9400,N_9401,N_9403,N_9405,N_9407,N_9409,N_9411,N_9414,N_9415,N_9416,N_9420,N_9421,N_9422,N_9425,N_9426,N_9427,N_9428,N_9429,N_9432,N_9434,N_9435,N_9436,N_9439,N_9440,N_9441,N_9444,N_9445,N_9446,N_9447,N_9452,N_9453,N_9457,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9478,N_9479,N_9480,N_9481,N_9482,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9505,N_9506,N_9509,N_9510,N_9516,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9534,N_9535,N_9537,N_9538,N_9539,N_9542,N_9544,N_9546,N_9548,N_9550,N_9551,N_9552,N_9554,N_9557,N_9558,N_9559,N_9561,N_9562,N_9563,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9577,N_9578,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9587,N_9589,N_9591,N_9592,N_9597,N_9600,N_9601,N_9603,N_9604,N_9605,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9617,N_9619,N_9620,N_9621,N_9622,N_9623,N_9626,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9637,N_9639,N_9641,N_9642,N_9644,N_9645,N_9646,N_9647,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9659,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9669,N_9670,N_9672,N_9673,N_9674,N_9676,N_9677,N_9678,N_9679,N_9682,N_9685,N_9687,N_9688,N_9689,N_9692,N_9693,N_9694,N_9697,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9713,N_9714,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9732,N_9735,N_9737,N_9740,N_9742,N_9746,N_9754,N_9755,N_9760,N_9761,N_9764,N_9767,N_9769,N_9771,N_9772,N_9774,N_9776,N_9777,N_9778,N_9780,N_9781,N_9783,N_9786,N_9788,N_9789,N_9791,N_9792,N_9793,N_9794,N_9795,N_9799,N_9800,N_9802,N_9803,N_9805,N_9808,N_9809,N_9811,N_9813,N_9814,N_9815,N_9817,N_9819,N_9821,N_9822,N_9823,N_9825,N_9827,N_9828,N_9829,N_9830,N_9832,N_9833,N_9834,N_9837,N_9838,N_9839,N_9840,N_9841,N_9843,N_9844,N_9845,N_9847,N_9848,N_9849,N_9850,N_9852,N_9857,N_9858,N_9859,N_9860,N_9864,N_9865,N_9866,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9875,N_9877,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9888,N_9890,N_9891,N_9892,N_9893,N_9894,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9907,N_9910,N_9912,N_9914,N_9915,N_9920,N_9921,N_9924,N_9926,N_9927,N_9929,N_9931,N_9932,N_9933,N_9934,N_9936,N_9937,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9951,N_9952,N_9955,N_9956,N_9957,N_9959,N_9961,N_9962,N_9965,N_9966,N_9967,N_9968,N_9970,N_9973,N_9975,N_9979,N_9980,N_9981,N_9982,N_9984,N_9985,N_9987,N_9989,N_9990,N_9991,N_9993,N_9995,N_9997,N_9999;
xnor U0 (N_0,In_839,In_194);
xnor U1 (N_1,In_940,In_22);
xnor U2 (N_2,In_314,In_925);
or U3 (N_3,In_782,In_934);
or U4 (N_4,In_767,In_198);
and U5 (N_5,In_472,In_455);
xor U6 (N_6,In_571,In_698);
or U7 (N_7,In_538,In_360);
nand U8 (N_8,In_948,In_281);
nand U9 (N_9,In_971,In_844);
nand U10 (N_10,In_53,In_130);
nor U11 (N_11,In_846,In_123);
or U12 (N_12,In_81,In_254);
xnor U13 (N_13,In_329,In_45);
nand U14 (N_14,In_458,In_471);
xor U15 (N_15,In_299,In_745);
nor U16 (N_16,In_232,In_873);
xor U17 (N_17,In_319,In_418);
and U18 (N_18,In_772,In_167);
xor U19 (N_19,In_749,In_223);
xor U20 (N_20,In_808,In_568);
or U21 (N_21,In_677,In_193);
xor U22 (N_22,In_457,In_738);
nor U23 (N_23,In_180,In_32);
nand U24 (N_24,In_431,In_737);
nand U25 (N_25,In_57,In_803);
or U26 (N_26,In_91,In_220);
xor U27 (N_27,In_18,In_960);
nand U28 (N_28,In_906,In_185);
nand U29 (N_29,In_450,In_36);
xor U30 (N_30,In_136,In_325);
nand U31 (N_31,In_996,In_693);
and U32 (N_32,In_518,In_205);
nand U33 (N_33,In_357,In_736);
and U34 (N_34,In_424,In_597);
or U35 (N_35,In_927,In_886);
nor U36 (N_36,In_173,In_730);
or U37 (N_37,In_256,In_915);
xor U38 (N_38,In_134,In_499);
or U39 (N_39,In_346,In_747);
or U40 (N_40,In_542,In_689);
nor U41 (N_41,In_949,In_712);
xnor U42 (N_42,In_616,In_459);
xnor U43 (N_43,In_293,In_211);
and U44 (N_44,In_344,In_335);
or U45 (N_45,In_363,In_891);
and U46 (N_46,In_727,In_483);
or U47 (N_47,In_795,In_501);
and U48 (N_48,In_815,In_536);
or U49 (N_49,In_669,In_387);
nand U50 (N_50,In_74,In_48);
xnor U51 (N_51,In_365,In_402);
nor U52 (N_52,In_889,In_174);
xnor U53 (N_53,In_684,In_87);
or U54 (N_54,In_33,In_354);
or U55 (N_55,In_153,In_287);
or U56 (N_56,In_54,In_160);
or U57 (N_57,In_516,In_212);
xnor U58 (N_58,In_688,In_543);
or U59 (N_59,In_226,In_23);
nand U60 (N_60,In_559,In_961);
nand U61 (N_61,In_930,In_324);
nor U62 (N_62,In_312,In_3);
nand U63 (N_63,In_140,In_733);
nor U64 (N_64,In_389,In_526);
or U65 (N_65,In_98,In_842);
nor U66 (N_66,In_989,In_386);
and U67 (N_67,In_219,In_257);
nor U68 (N_68,In_676,In_432);
and U69 (N_69,In_61,In_297);
nor U70 (N_70,In_885,In_348);
xor U71 (N_71,In_711,In_638);
or U72 (N_72,In_14,In_233);
xnor U73 (N_73,In_908,In_548);
nand U74 (N_74,In_127,In_982);
and U75 (N_75,In_909,In_443);
xor U76 (N_76,In_343,In_63);
xor U77 (N_77,In_479,In_976);
nand U78 (N_78,In_739,In_979);
nor U79 (N_79,In_245,In_308);
nor U80 (N_80,In_300,In_251);
and U81 (N_81,In_465,In_784);
xor U82 (N_82,In_687,In_834);
nand U83 (N_83,In_30,In_635);
and U84 (N_84,In_980,In_657);
nand U85 (N_85,In_647,In_481);
nor U86 (N_86,In_392,In_436);
or U87 (N_87,In_316,In_261);
nand U88 (N_88,In_236,In_953);
and U89 (N_89,In_683,In_600);
xnor U90 (N_90,In_69,In_560);
xnor U91 (N_91,In_341,In_822);
or U92 (N_92,In_969,In_119);
and U93 (N_93,In_804,In_276);
nor U94 (N_94,In_285,In_120);
and U95 (N_95,In_611,In_983);
xnor U96 (N_96,In_621,In_932);
xor U97 (N_97,In_691,In_235);
and U98 (N_98,In_984,In_507);
and U99 (N_99,In_517,In_672);
nand U100 (N_100,In_385,In_661);
nand U101 (N_101,In_203,In_410);
nor U102 (N_102,In_905,In_441);
or U103 (N_103,In_463,In_615);
xnor U104 (N_104,In_567,In_572);
xnor U105 (N_105,In_487,In_322);
and U106 (N_106,In_475,In_556);
and U107 (N_107,In_342,In_665);
xnor U108 (N_108,In_337,In_714);
nor U109 (N_109,In_296,In_679);
xor U110 (N_110,In_188,In_849);
nor U111 (N_111,In_25,In_291);
nand U112 (N_112,In_345,In_10);
nand U113 (N_113,In_263,In_230);
xor U114 (N_114,In_710,In_419);
and U115 (N_115,In_29,In_309);
nor U116 (N_116,In_532,In_627);
nand U117 (N_117,In_580,In_164);
xor U118 (N_118,In_139,In_214);
or U119 (N_119,In_840,In_678);
or U120 (N_120,In_244,In_799);
or U121 (N_121,In_913,In_636);
xor U122 (N_122,In_366,In_90);
or U123 (N_123,In_525,In_398);
nand U124 (N_124,In_998,In_655);
or U125 (N_125,In_588,In_488);
nand U126 (N_126,In_495,In_978);
nand U127 (N_127,In_238,In_938);
nor U128 (N_128,In_225,In_381);
nor U129 (N_129,In_408,In_875);
and U130 (N_130,In_610,In_155);
nand U131 (N_131,In_768,In_492);
nand U132 (N_132,In_700,In_439);
nor U133 (N_133,In_202,In_821);
xor U134 (N_134,In_511,In_959);
nor U135 (N_135,In_453,In_673);
nor U136 (N_136,In_292,In_964);
nor U137 (N_137,In_863,In_777);
xor U138 (N_138,In_977,In_586);
or U139 (N_139,In_267,In_551);
nand U140 (N_140,In_310,In_447);
nor U141 (N_141,In_874,In_857);
nand U142 (N_142,In_259,In_380);
or U143 (N_143,In_390,In_550);
and U144 (N_144,In_731,In_861);
xnor U145 (N_145,In_829,In_544);
xnor U146 (N_146,In_21,In_192);
xor U147 (N_147,In_473,In_916);
xnor U148 (N_148,In_854,In_781);
nor U149 (N_149,In_651,In_968);
and U150 (N_150,In_106,In_869);
nand U151 (N_151,In_533,In_509);
nand U152 (N_152,In_872,In_255);
nand U153 (N_153,In_761,In_448);
or U154 (N_154,In_302,In_719);
nor U155 (N_155,In_89,In_537);
nand U156 (N_156,In_704,In_34);
or U157 (N_157,In_653,In_394);
nor U158 (N_158,In_288,In_512);
nand U159 (N_159,In_118,In_362);
nand U160 (N_160,In_248,In_209);
xor U161 (N_161,In_38,In_372);
nor U162 (N_162,In_933,In_7);
nand U163 (N_163,In_941,In_650);
or U164 (N_164,In_950,In_786);
and U165 (N_165,In_5,In_818);
nor U166 (N_166,In_125,In_830);
nor U167 (N_167,In_850,In_279);
nor U168 (N_168,In_298,In_612);
nand U169 (N_169,In_806,In_234);
and U170 (N_170,In_68,In_515);
and U171 (N_171,In_758,In_660);
or U172 (N_172,In_27,In_368);
nand U173 (N_173,In_218,In_652);
or U174 (N_174,In_617,In_801);
and U175 (N_175,In_67,In_184);
nand U176 (N_176,In_816,In_563);
and U177 (N_177,In_51,In_486);
and U178 (N_178,In_490,In_963);
and U179 (N_179,In_843,In_867);
xnor U180 (N_180,In_55,In_945);
xnor U181 (N_181,In_581,In_535);
or U182 (N_182,In_461,In_630);
nand U183 (N_183,In_485,In_78);
xnor U184 (N_184,In_216,In_413);
nor U185 (N_185,In_546,In_502);
nand U186 (N_186,In_491,In_370);
nor U187 (N_187,In_765,In_128);
or U188 (N_188,In_832,In_168);
xnor U189 (N_189,In_553,In_605);
or U190 (N_190,In_83,In_96);
nand U191 (N_191,In_587,In_24);
nor U192 (N_192,In_819,In_549);
or U193 (N_193,In_631,In_73);
and U194 (N_194,In_283,In_769);
or U195 (N_195,In_910,In_273);
xor U196 (N_196,In_468,In_975);
or U197 (N_197,In_703,In_265);
xnor U198 (N_198,In_250,In_303);
nor U199 (N_199,In_871,In_117);
xnor U200 (N_200,In_921,In_845);
nand U201 (N_201,In_80,In_156);
or U202 (N_202,In_620,In_506);
xor U203 (N_203,In_182,In_904);
nand U204 (N_204,In_753,In_760);
xor U205 (N_205,In_422,In_741);
and U206 (N_206,In_695,In_121);
nand U207 (N_207,In_56,In_562);
and U208 (N_208,In_498,In_624);
or U209 (N_209,In_353,In_809);
or U210 (N_210,In_877,In_527);
or U211 (N_211,In_375,In_124);
xnor U212 (N_212,In_951,In_242);
xnor U213 (N_213,In_409,In_897);
nor U214 (N_214,In_157,In_0);
and U215 (N_215,In_791,In_200);
xnor U216 (N_216,In_268,In_274);
nand U217 (N_217,In_939,In_505);
nor U218 (N_218,In_866,In_82);
nor U219 (N_219,In_755,In_813);
nor U220 (N_220,In_692,In_189);
and U221 (N_221,In_920,In_350);
nand U222 (N_222,In_247,In_898);
xnor U223 (N_223,In_187,In_606);
or U224 (N_224,In_847,In_545);
or U225 (N_225,In_271,In_554);
nand U226 (N_226,In_856,In_882);
and U227 (N_227,In_629,In_361);
xnor U228 (N_228,In_997,In_541);
or U229 (N_229,In_272,In_520);
nand U230 (N_230,In_162,In_446);
or U231 (N_231,In_955,In_331);
nand U232 (N_232,In_97,In_890);
nor U233 (N_233,In_681,In_379);
nand U234 (N_234,In_317,In_326);
or U235 (N_235,In_59,In_540);
xnor U236 (N_236,In_70,In_425);
xnor U237 (N_237,In_426,In_315);
nor U238 (N_238,In_417,In_6);
nor U239 (N_239,In_384,In_523);
nor U240 (N_240,In_65,In_812);
nor U241 (N_241,In_183,In_113);
xnor U242 (N_242,In_323,In_111);
or U243 (N_243,In_922,In_132);
nand U244 (N_244,In_107,In_43);
nor U245 (N_245,In_911,In_570);
nor U246 (N_246,In_790,In_510);
and U247 (N_247,In_598,In_601);
nand U248 (N_248,In_919,In_508);
xor U249 (N_249,In_207,In_148);
or U250 (N_250,In_364,In_286);
nor U251 (N_251,In_682,In_428);
or U252 (N_252,In_399,In_114);
and U253 (N_253,In_171,In_833);
or U254 (N_254,In_705,In_675);
nand U255 (N_255,In_775,In_237);
xnor U256 (N_256,In_870,In_987);
nand U257 (N_257,In_926,In_456);
or U258 (N_258,In_878,In_50);
or U259 (N_259,In_907,In_109);
or U260 (N_260,In_221,In_169);
xor U261 (N_261,In_720,In_264);
xnor U262 (N_262,In_99,In_590);
nand U263 (N_263,In_593,In_724);
xor U264 (N_264,In_599,In_800);
nor U265 (N_265,In_241,In_60);
nand U266 (N_266,In_307,In_92);
xor U267 (N_267,In_680,In_530);
xnor U268 (N_268,In_284,In_862);
nand U269 (N_269,In_912,In_622);
nor U270 (N_270,In_46,In_974);
xnor U271 (N_271,In_64,In_466);
nand U272 (N_272,In_88,In_573);
nor U273 (N_273,In_826,In_584);
or U274 (N_274,In_79,In_835);
xor U275 (N_275,In_914,In_947);
nor U276 (N_276,In_539,In_158);
and U277 (N_277,In_289,In_513);
xnor U278 (N_278,In_706,In_514);
and U279 (N_279,In_4,In_150);
nand U280 (N_280,In_376,In_792);
xnor U281 (N_281,In_894,In_699);
xor U282 (N_282,In_16,In_28);
xnor U283 (N_283,In_391,In_901);
xor U284 (N_284,In_58,In_336);
or U285 (N_285,In_715,In_957);
nand U286 (N_286,In_557,In_340);
nor U287 (N_287,In_49,In_41);
or U288 (N_288,In_531,In_306);
or U289 (N_289,In_269,In_744);
or U290 (N_290,In_602,In_865);
xor U291 (N_291,In_112,In_547);
and U292 (N_292,In_787,In_773);
nand U293 (N_293,In_824,In_435);
and U294 (N_294,In_240,In_311);
nor U295 (N_295,In_334,In_102);
or U296 (N_296,In_37,In_318);
xor U297 (N_297,In_433,In_469);
xor U298 (N_298,In_440,In_496);
nand U299 (N_299,In_94,In_565);
nor U300 (N_300,In_838,In_105);
nand U301 (N_301,In_243,In_659);
nor U302 (N_302,In_625,In_852);
xnor U303 (N_303,In_860,In_674);
and U304 (N_304,In_195,In_215);
xor U305 (N_305,In_393,In_766);
and U306 (N_306,In_880,In_258);
and U307 (N_307,In_990,In_848);
xor U308 (N_308,In_15,In_66);
xor U309 (N_309,In_742,In_163);
or U310 (N_310,In_789,In_131);
nor U311 (N_311,In_825,In_110);
nand U312 (N_312,In_640,In_966);
and U313 (N_313,In_999,In_476);
nand U314 (N_314,In_985,In_152);
and U315 (N_315,In_895,In_952);
and U316 (N_316,In_454,In_991);
nor U317 (N_317,In_764,In_864);
or U318 (N_318,In_759,In_278);
nor U319 (N_319,In_367,In_493);
nor U320 (N_320,In_396,In_589);
and U321 (N_321,In_115,In_266);
nor U322 (N_322,In_858,In_378);
nor U323 (N_323,In_579,In_355);
and U324 (N_324,In_702,In_841);
nor U325 (N_325,In_827,In_972);
and U326 (N_326,In_668,In_178);
nor U327 (N_327,In_592,In_726);
nand U328 (N_328,In_227,In_477);
and U329 (N_329,In_662,In_690);
or U330 (N_330,In_328,In_851);
xnor U331 (N_331,In_718,In_994);
or U332 (N_332,In_438,In_645);
xor U333 (N_333,In_137,In_262);
nand U334 (N_334,In_893,In_524);
xnor U335 (N_335,In_701,In_519);
nor U336 (N_336,In_321,In_100);
xnor U337 (N_337,In_144,In_552);
nor U338 (N_338,In_482,In_484);
or U339 (N_339,In_239,In_280);
nand U340 (N_340,In_903,In_754);
nor U341 (N_341,In_561,In_521);
and U342 (N_342,In_9,In_956);
and U343 (N_343,In_721,In_654);
xnor U344 (N_344,In_722,In_748);
or U345 (N_345,In_814,In_837);
xnor U346 (N_346,In_249,In_17);
nand U347 (N_347,In_222,In_805);
xnor U348 (N_348,In_534,In_667);
nand U349 (N_349,In_958,In_888);
nor U350 (N_350,In_569,In_883);
or U351 (N_351,In_937,In_147);
nand U352 (N_352,In_793,In_474);
nand U353 (N_353,In_771,In_836);
or U354 (N_354,In_725,In_811);
or U355 (N_355,In_802,In_172);
nor U356 (N_356,In_201,In_962);
or U357 (N_357,In_853,In_778);
nand U358 (N_358,In_750,In_176);
xnor U359 (N_359,In_252,In_896);
nand U360 (N_360,In_400,In_967);
and U361 (N_361,In_151,In_253);
xor U362 (N_362,In_728,In_859);
nand U363 (N_363,In_649,In_277);
and U364 (N_364,In_626,In_373);
nand U365 (N_365,In_327,In_820);
nand U366 (N_366,In_26,In_696);
and U367 (N_367,In_406,In_154);
nor U368 (N_368,In_713,In_663);
nand U369 (N_369,In_146,In_723);
nor U370 (N_370,In_191,In_648);
nor U371 (N_371,In_928,In_528);
nand U372 (N_372,In_887,In_72);
nor U373 (N_373,In_116,In_992);
nor U374 (N_374,In_47,In_217);
or U375 (N_375,In_434,In_179);
nand U376 (N_376,In_732,In_412);
nor U377 (N_377,In_141,In_986);
nor U378 (N_378,In_785,In_646);
nand U379 (N_379,In_388,In_213);
nand U380 (N_380,In_405,In_270);
nand U381 (N_381,In_103,In_19);
and U382 (N_382,In_632,In_159);
xor U383 (N_383,In_395,In_199);
xnor U384 (N_384,In_609,In_642);
and U385 (N_385,In_855,In_84);
or U386 (N_386,In_301,In_603);
and U387 (N_387,In_988,In_31);
nand U388 (N_388,In_884,In_429);
xnor U389 (N_389,In_196,In_145);
xnor U390 (N_390,In_282,In_946);
nor U391 (N_391,In_794,In_2);
or U392 (N_392,In_564,In_574);
and U393 (N_393,In_349,In_607);
xor U394 (N_394,In_42,In_451);
xnor U395 (N_395,In_104,In_170);
nor U396 (N_396,In_729,In_437);
or U397 (N_397,In_304,In_707);
and U398 (N_398,In_746,In_685);
and U399 (N_399,In_585,In_470);
or U400 (N_400,In_504,In_797);
nor U401 (N_401,In_467,In_210);
and U402 (N_402,In_313,In_807);
nand U403 (N_403,In_138,In_558);
xnor U404 (N_404,In_931,In_965);
nor U405 (N_405,In_973,In_555);
xor U406 (N_406,In_798,In_101);
xnor U407 (N_407,In_44,In_595);
xnor U408 (N_408,In_942,In_529);
nand U409 (N_409,In_407,In_817);
or U410 (N_410,In_810,In_197);
nor U411 (N_411,In_779,In_697);
xor U412 (N_412,In_421,In_780);
and U413 (N_413,In_382,In_397);
and U414 (N_414,In_166,In_416);
xnor U415 (N_415,In_566,In_623);
or U416 (N_416,In_671,In_757);
nor U417 (N_417,In_35,In_489);
and U418 (N_418,In_899,In_943);
xnor U419 (N_419,In_62,In_352);
nor U420 (N_420,In_954,In_756);
nand U421 (N_421,In_831,In_411);
or U422 (N_422,In_776,In_330);
nor U423 (N_423,In_204,In_20);
or U424 (N_424,In_305,In_497);
or U425 (N_425,In_135,In_604);
nand U426 (N_426,In_929,In_246);
or U427 (N_427,In_613,In_634);
nor U428 (N_428,In_442,In_93);
xor U429 (N_429,In_77,In_1);
nand U430 (N_430,In_369,In_414);
xor U431 (N_431,In_377,In_494);
nand U432 (N_432,In_639,In_177);
or U433 (N_433,In_161,In_462);
or U434 (N_434,In_39,In_637);
nand U435 (N_435,In_290,In_480);
nand U436 (N_436,In_347,In_332);
or U437 (N_437,In_401,In_75);
and U438 (N_438,In_619,In_923);
and U439 (N_439,In_892,In_614);
xor U440 (N_440,In_320,In_224);
and U441 (N_441,In_783,In_294);
nand U442 (N_442,In_464,In_774);
nor U443 (N_443,In_76,In_628);
nand U444 (N_444,In_694,In_181);
or U445 (N_445,In_734,In_770);
or U446 (N_446,In_333,In_752);
or U447 (N_447,In_709,In_666);
nand U448 (N_448,In_743,In_981);
xor U449 (N_449,In_175,In_763);
xnor U450 (N_450,In_993,In_576);
or U451 (N_451,In_740,In_275);
or U452 (N_452,In_478,In_460);
nand U453 (N_453,In_71,In_228);
and U454 (N_454,In_359,In_445);
or U455 (N_455,In_186,In_11);
nand U456 (N_456,In_944,In_85);
and U457 (N_457,In_40,In_995);
nand U458 (N_458,In_762,In_208);
nor U459 (N_459,In_633,In_356);
nor U460 (N_460,In_129,In_500);
xnor U461 (N_461,In_404,In_374);
and U462 (N_462,In_165,In_823);
xnor U463 (N_463,In_664,In_876);
or U464 (N_464,In_108,In_716);
xnor U465 (N_465,In_708,In_371);
and U466 (N_466,In_686,In_403);
or U467 (N_467,In_415,In_423);
or U468 (N_468,In_86,In_126);
nor U469 (N_469,In_917,In_522);
nand U470 (N_470,In_582,In_594);
nor U471 (N_471,In_260,In_751);
and U472 (N_472,In_583,In_190);
or U473 (N_473,In_142,In_881);
nand U474 (N_474,In_577,In_449);
nand U475 (N_475,In_13,In_828);
and U476 (N_476,In_643,In_591);
and U477 (N_477,In_936,In_575);
nand U478 (N_478,In_879,In_149);
and U479 (N_479,In_796,In_596);
nand U480 (N_480,In_52,In_206);
nor U481 (N_481,In_8,In_618);
and U482 (N_482,In_420,In_383);
and U483 (N_483,In_735,In_788);
xor U484 (N_484,In_644,In_918);
or U485 (N_485,In_295,In_452);
nor U486 (N_486,In_122,In_95);
nand U487 (N_487,In_868,In_444);
or U488 (N_488,In_351,In_503);
nor U489 (N_489,In_658,In_902);
nand U490 (N_490,In_970,In_229);
xor U491 (N_491,In_339,In_608);
nor U492 (N_492,In_231,In_578);
nor U493 (N_493,In_430,In_338);
nor U494 (N_494,In_143,In_427);
or U495 (N_495,In_641,In_900);
and U496 (N_496,In_717,In_935);
or U497 (N_497,In_656,In_133);
nand U498 (N_498,In_924,In_670);
or U499 (N_499,In_12,In_358);
xor U500 (N_500,In_70,In_934);
nand U501 (N_501,In_158,In_21);
or U502 (N_502,In_952,In_436);
nand U503 (N_503,In_619,In_385);
or U504 (N_504,In_285,In_441);
xnor U505 (N_505,In_214,In_839);
nand U506 (N_506,In_184,In_249);
and U507 (N_507,In_389,In_380);
and U508 (N_508,In_198,In_328);
or U509 (N_509,In_597,In_661);
or U510 (N_510,In_876,In_139);
nor U511 (N_511,In_126,In_24);
xnor U512 (N_512,In_292,In_530);
xor U513 (N_513,In_124,In_111);
xor U514 (N_514,In_379,In_407);
nand U515 (N_515,In_26,In_32);
xor U516 (N_516,In_295,In_835);
and U517 (N_517,In_296,In_665);
nor U518 (N_518,In_607,In_906);
nand U519 (N_519,In_431,In_484);
xnor U520 (N_520,In_217,In_415);
nor U521 (N_521,In_308,In_880);
and U522 (N_522,In_595,In_599);
xnor U523 (N_523,In_548,In_239);
or U524 (N_524,In_116,In_798);
nand U525 (N_525,In_29,In_48);
or U526 (N_526,In_69,In_890);
or U527 (N_527,In_107,In_569);
xnor U528 (N_528,In_138,In_41);
xnor U529 (N_529,In_745,In_256);
nor U530 (N_530,In_971,In_513);
xnor U531 (N_531,In_852,In_292);
nor U532 (N_532,In_459,In_57);
xor U533 (N_533,In_467,In_534);
or U534 (N_534,In_186,In_157);
nand U535 (N_535,In_439,In_762);
or U536 (N_536,In_635,In_892);
or U537 (N_537,In_598,In_142);
and U538 (N_538,In_126,In_930);
and U539 (N_539,In_599,In_704);
xor U540 (N_540,In_521,In_31);
or U541 (N_541,In_866,In_526);
xor U542 (N_542,In_807,In_332);
nor U543 (N_543,In_865,In_987);
nor U544 (N_544,In_40,In_816);
and U545 (N_545,In_100,In_833);
and U546 (N_546,In_309,In_492);
or U547 (N_547,In_876,In_147);
xnor U548 (N_548,In_588,In_584);
nor U549 (N_549,In_680,In_843);
and U550 (N_550,In_539,In_210);
nand U551 (N_551,In_810,In_566);
nor U552 (N_552,In_763,In_640);
nand U553 (N_553,In_831,In_19);
nor U554 (N_554,In_926,In_804);
and U555 (N_555,In_216,In_985);
xor U556 (N_556,In_30,In_918);
and U557 (N_557,In_373,In_394);
nor U558 (N_558,In_589,In_778);
xnor U559 (N_559,In_650,In_844);
or U560 (N_560,In_758,In_329);
and U561 (N_561,In_270,In_23);
or U562 (N_562,In_651,In_893);
nand U563 (N_563,In_286,In_821);
xor U564 (N_564,In_995,In_595);
or U565 (N_565,In_456,In_771);
xor U566 (N_566,In_491,In_990);
xor U567 (N_567,In_581,In_44);
or U568 (N_568,In_969,In_860);
xnor U569 (N_569,In_537,In_79);
and U570 (N_570,In_160,In_583);
nand U571 (N_571,In_338,In_582);
nor U572 (N_572,In_602,In_488);
and U573 (N_573,In_33,In_707);
xor U574 (N_574,In_503,In_670);
nor U575 (N_575,In_274,In_680);
xnor U576 (N_576,In_304,In_20);
and U577 (N_577,In_804,In_706);
and U578 (N_578,In_975,In_489);
xor U579 (N_579,In_131,In_205);
nor U580 (N_580,In_976,In_125);
nand U581 (N_581,In_350,In_892);
xor U582 (N_582,In_466,In_914);
nand U583 (N_583,In_876,In_840);
nor U584 (N_584,In_610,In_919);
nor U585 (N_585,In_371,In_250);
nand U586 (N_586,In_785,In_782);
nor U587 (N_587,In_262,In_780);
nor U588 (N_588,In_852,In_337);
nor U589 (N_589,In_362,In_580);
nor U590 (N_590,In_127,In_765);
xnor U591 (N_591,In_111,In_890);
nand U592 (N_592,In_114,In_28);
and U593 (N_593,In_975,In_86);
nor U594 (N_594,In_649,In_927);
or U595 (N_595,In_239,In_664);
nor U596 (N_596,In_118,In_270);
nand U597 (N_597,In_183,In_167);
nand U598 (N_598,In_286,In_731);
and U599 (N_599,In_119,In_900);
nor U600 (N_600,In_570,In_959);
and U601 (N_601,In_213,In_233);
and U602 (N_602,In_537,In_320);
or U603 (N_603,In_140,In_894);
and U604 (N_604,In_954,In_557);
xnor U605 (N_605,In_852,In_62);
or U606 (N_606,In_788,In_87);
nand U607 (N_607,In_512,In_455);
nand U608 (N_608,In_986,In_631);
xor U609 (N_609,In_524,In_25);
nand U610 (N_610,In_158,In_730);
xor U611 (N_611,In_953,In_323);
nor U612 (N_612,In_957,In_885);
or U613 (N_613,In_879,In_780);
xnor U614 (N_614,In_45,In_361);
and U615 (N_615,In_136,In_670);
nor U616 (N_616,In_110,In_788);
xor U617 (N_617,In_52,In_823);
nor U618 (N_618,In_122,In_315);
or U619 (N_619,In_587,In_179);
nand U620 (N_620,In_389,In_464);
or U621 (N_621,In_25,In_17);
xnor U622 (N_622,In_658,In_492);
and U623 (N_623,In_651,In_637);
nand U624 (N_624,In_502,In_984);
nand U625 (N_625,In_145,In_211);
nand U626 (N_626,In_768,In_506);
or U627 (N_627,In_560,In_754);
and U628 (N_628,In_566,In_367);
xor U629 (N_629,In_849,In_556);
nor U630 (N_630,In_852,In_416);
or U631 (N_631,In_477,In_174);
and U632 (N_632,In_837,In_473);
xnor U633 (N_633,In_294,In_848);
or U634 (N_634,In_782,In_249);
and U635 (N_635,In_436,In_479);
nor U636 (N_636,In_249,In_407);
xor U637 (N_637,In_909,In_750);
nor U638 (N_638,In_899,In_224);
xnor U639 (N_639,In_20,In_647);
nand U640 (N_640,In_420,In_109);
xor U641 (N_641,In_148,In_499);
nand U642 (N_642,In_559,In_597);
and U643 (N_643,In_65,In_639);
or U644 (N_644,In_526,In_832);
nand U645 (N_645,In_23,In_326);
xor U646 (N_646,In_9,In_302);
xnor U647 (N_647,In_238,In_509);
nor U648 (N_648,In_451,In_771);
and U649 (N_649,In_68,In_876);
xor U650 (N_650,In_558,In_497);
and U651 (N_651,In_489,In_907);
xor U652 (N_652,In_361,In_209);
xor U653 (N_653,In_843,In_702);
nand U654 (N_654,In_536,In_51);
nand U655 (N_655,In_107,In_115);
xor U656 (N_656,In_390,In_50);
nor U657 (N_657,In_495,In_190);
and U658 (N_658,In_645,In_906);
nor U659 (N_659,In_41,In_966);
xor U660 (N_660,In_427,In_821);
or U661 (N_661,In_829,In_709);
xor U662 (N_662,In_778,In_628);
nor U663 (N_663,In_571,In_664);
nor U664 (N_664,In_696,In_896);
nand U665 (N_665,In_972,In_494);
or U666 (N_666,In_3,In_144);
nand U667 (N_667,In_934,In_458);
or U668 (N_668,In_553,In_476);
nor U669 (N_669,In_577,In_793);
or U670 (N_670,In_412,In_590);
nor U671 (N_671,In_325,In_322);
nand U672 (N_672,In_253,In_612);
nand U673 (N_673,In_519,In_510);
xor U674 (N_674,In_357,In_682);
or U675 (N_675,In_848,In_167);
or U676 (N_676,In_887,In_845);
or U677 (N_677,In_444,In_93);
nor U678 (N_678,In_698,In_825);
xnor U679 (N_679,In_245,In_936);
nor U680 (N_680,In_440,In_447);
and U681 (N_681,In_879,In_109);
nor U682 (N_682,In_354,In_838);
nand U683 (N_683,In_587,In_108);
and U684 (N_684,In_271,In_548);
and U685 (N_685,In_794,In_623);
nand U686 (N_686,In_670,In_204);
xor U687 (N_687,In_817,In_25);
and U688 (N_688,In_769,In_411);
and U689 (N_689,In_541,In_331);
xor U690 (N_690,In_39,In_404);
and U691 (N_691,In_420,In_753);
xnor U692 (N_692,In_826,In_197);
nand U693 (N_693,In_253,In_872);
and U694 (N_694,In_445,In_199);
or U695 (N_695,In_661,In_751);
xnor U696 (N_696,In_56,In_328);
xnor U697 (N_697,In_649,In_164);
nor U698 (N_698,In_963,In_248);
nand U699 (N_699,In_85,In_848);
or U700 (N_700,In_795,In_493);
and U701 (N_701,In_584,In_62);
nand U702 (N_702,In_295,In_937);
nor U703 (N_703,In_719,In_585);
xor U704 (N_704,In_582,In_299);
xnor U705 (N_705,In_571,In_678);
and U706 (N_706,In_256,In_945);
or U707 (N_707,In_880,In_136);
nor U708 (N_708,In_754,In_410);
nand U709 (N_709,In_517,In_975);
and U710 (N_710,In_618,In_127);
nand U711 (N_711,In_106,In_617);
xor U712 (N_712,In_809,In_498);
nand U713 (N_713,In_455,In_490);
nor U714 (N_714,In_407,In_956);
or U715 (N_715,In_173,In_717);
and U716 (N_716,In_537,In_637);
nand U717 (N_717,In_902,In_545);
xor U718 (N_718,In_699,In_435);
xnor U719 (N_719,In_871,In_601);
or U720 (N_720,In_866,In_470);
nand U721 (N_721,In_185,In_189);
nor U722 (N_722,In_472,In_293);
xor U723 (N_723,In_530,In_53);
nand U724 (N_724,In_592,In_886);
and U725 (N_725,In_717,In_465);
nor U726 (N_726,In_610,In_715);
xor U727 (N_727,In_324,In_481);
nor U728 (N_728,In_557,In_465);
nand U729 (N_729,In_707,In_919);
and U730 (N_730,In_316,In_528);
xor U731 (N_731,In_899,In_440);
nor U732 (N_732,In_827,In_82);
and U733 (N_733,In_504,In_206);
and U734 (N_734,In_312,In_496);
nand U735 (N_735,In_955,In_686);
nand U736 (N_736,In_838,In_625);
or U737 (N_737,In_873,In_10);
nor U738 (N_738,In_846,In_532);
nand U739 (N_739,In_440,In_704);
xnor U740 (N_740,In_213,In_914);
xnor U741 (N_741,In_253,In_160);
nor U742 (N_742,In_838,In_20);
or U743 (N_743,In_203,In_619);
nand U744 (N_744,In_633,In_832);
nand U745 (N_745,In_221,In_859);
nand U746 (N_746,In_403,In_60);
or U747 (N_747,In_974,In_833);
xnor U748 (N_748,In_619,In_589);
xnor U749 (N_749,In_585,In_318);
xor U750 (N_750,In_98,In_543);
or U751 (N_751,In_185,In_910);
and U752 (N_752,In_644,In_621);
nand U753 (N_753,In_722,In_996);
nand U754 (N_754,In_892,In_938);
and U755 (N_755,In_451,In_423);
xnor U756 (N_756,In_3,In_799);
or U757 (N_757,In_82,In_906);
and U758 (N_758,In_706,In_395);
xnor U759 (N_759,In_301,In_711);
and U760 (N_760,In_260,In_841);
or U761 (N_761,In_701,In_461);
and U762 (N_762,In_835,In_131);
xnor U763 (N_763,In_355,In_60);
nor U764 (N_764,In_12,In_801);
xnor U765 (N_765,In_532,In_481);
nand U766 (N_766,In_358,In_532);
xor U767 (N_767,In_100,In_254);
nor U768 (N_768,In_445,In_785);
nand U769 (N_769,In_692,In_655);
xor U770 (N_770,In_568,In_81);
xor U771 (N_771,In_244,In_364);
xor U772 (N_772,In_922,In_300);
xor U773 (N_773,In_363,In_503);
nand U774 (N_774,In_702,In_720);
nand U775 (N_775,In_505,In_5);
xor U776 (N_776,In_137,In_843);
and U777 (N_777,In_605,In_942);
or U778 (N_778,In_698,In_813);
xnor U779 (N_779,In_366,In_551);
nor U780 (N_780,In_824,In_137);
nor U781 (N_781,In_377,In_933);
nor U782 (N_782,In_90,In_878);
and U783 (N_783,In_961,In_306);
nor U784 (N_784,In_732,In_617);
and U785 (N_785,In_412,In_118);
xnor U786 (N_786,In_160,In_682);
xnor U787 (N_787,In_757,In_500);
nand U788 (N_788,In_69,In_878);
and U789 (N_789,In_786,In_679);
and U790 (N_790,In_246,In_336);
nor U791 (N_791,In_692,In_378);
or U792 (N_792,In_290,In_113);
nand U793 (N_793,In_36,In_505);
and U794 (N_794,In_928,In_483);
xor U795 (N_795,In_194,In_101);
and U796 (N_796,In_645,In_889);
xnor U797 (N_797,In_895,In_553);
nand U798 (N_798,In_385,In_569);
xor U799 (N_799,In_876,In_588);
or U800 (N_800,In_745,In_486);
nand U801 (N_801,In_131,In_306);
xnor U802 (N_802,In_387,In_443);
or U803 (N_803,In_998,In_907);
nor U804 (N_804,In_906,In_106);
nor U805 (N_805,In_420,In_325);
nor U806 (N_806,In_695,In_148);
and U807 (N_807,In_315,In_23);
nand U808 (N_808,In_738,In_930);
and U809 (N_809,In_550,In_830);
nor U810 (N_810,In_118,In_827);
and U811 (N_811,In_107,In_518);
nor U812 (N_812,In_127,In_73);
nand U813 (N_813,In_301,In_700);
nand U814 (N_814,In_847,In_896);
and U815 (N_815,In_594,In_140);
or U816 (N_816,In_247,In_45);
nor U817 (N_817,In_308,In_135);
and U818 (N_818,In_201,In_972);
and U819 (N_819,In_53,In_815);
nand U820 (N_820,In_525,In_277);
and U821 (N_821,In_388,In_403);
and U822 (N_822,In_953,In_168);
or U823 (N_823,In_845,In_150);
and U824 (N_824,In_324,In_788);
and U825 (N_825,In_140,In_615);
or U826 (N_826,In_70,In_476);
nand U827 (N_827,In_837,In_147);
and U828 (N_828,In_22,In_749);
nand U829 (N_829,In_123,In_416);
and U830 (N_830,In_303,In_112);
nor U831 (N_831,In_237,In_907);
nand U832 (N_832,In_116,In_959);
or U833 (N_833,In_956,In_902);
nand U834 (N_834,In_266,In_501);
nor U835 (N_835,In_928,In_819);
or U836 (N_836,In_720,In_721);
xnor U837 (N_837,In_134,In_580);
nor U838 (N_838,In_489,In_567);
or U839 (N_839,In_651,In_588);
xnor U840 (N_840,In_294,In_403);
nor U841 (N_841,In_254,In_873);
xor U842 (N_842,In_980,In_778);
xor U843 (N_843,In_580,In_471);
or U844 (N_844,In_227,In_410);
xnor U845 (N_845,In_330,In_970);
xnor U846 (N_846,In_883,In_350);
nor U847 (N_847,In_651,In_897);
xnor U848 (N_848,In_732,In_869);
nand U849 (N_849,In_894,In_980);
nand U850 (N_850,In_566,In_96);
and U851 (N_851,In_854,In_391);
nor U852 (N_852,In_462,In_644);
xor U853 (N_853,In_425,In_826);
or U854 (N_854,In_11,In_912);
xnor U855 (N_855,In_85,In_5);
and U856 (N_856,In_322,In_389);
nor U857 (N_857,In_710,In_532);
nor U858 (N_858,In_565,In_612);
and U859 (N_859,In_13,In_9);
xnor U860 (N_860,In_875,In_490);
or U861 (N_861,In_214,In_851);
nor U862 (N_862,In_714,In_851);
and U863 (N_863,In_506,In_750);
xor U864 (N_864,In_987,In_251);
nor U865 (N_865,In_485,In_69);
or U866 (N_866,In_463,In_806);
or U867 (N_867,In_132,In_57);
xnor U868 (N_868,In_165,In_743);
xnor U869 (N_869,In_829,In_440);
and U870 (N_870,In_163,In_866);
and U871 (N_871,In_836,In_19);
nor U872 (N_872,In_501,In_63);
or U873 (N_873,In_111,In_481);
nand U874 (N_874,In_588,In_729);
or U875 (N_875,In_66,In_777);
or U876 (N_876,In_214,In_735);
nor U877 (N_877,In_97,In_138);
nor U878 (N_878,In_780,In_803);
and U879 (N_879,In_267,In_44);
xnor U880 (N_880,In_918,In_22);
or U881 (N_881,In_350,In_305);
or U882 (N_882,In_149,In_56);
or U883 (N_883,In_276,In_608);
or U884 (N_884,In_122,In_487);
nand U885 (N_885,In_267,In_588);
and U886 (N_886,In_981,In_27);
or U887 (N_887,In_23,In_535);
xor U888 (N_888,In_537,In_804);
xor U889 (N_889,In_236,In_433);
xnor U890 (N_890,In_664,In_812);
xor U891 (N_891,In_312,In_795);
xor U892 (N_892,In_486,In_427);
and U893 (N_893,In_691,In_564);
and U894 (N_894,In_498,In_603);
nor U895 (N_895,In_360,In_965);
nor U896 (N_896,In_44,In_858);
or U897 (N_897,In_294,In_600);
nor U898 (N_898,In_213,In_110);
xnor U899 (N_899,In_295,In_661);
or U900 (N_900,In_180,In_338);
nor U901 (N_901,In_481,In_380);
and U902 (N_902,In_359,In_189);
nand U903 (N_903,In_949,In_540);
or U904 (N_904,In_253,In_921);
xor U905 (N_905,In_477,In_808);
and U906 (N_906,In_903,In_676);
xor U907 (N_907,In_492,In_350);
and U908 (N_908,In_250,In_958);
xor U909 (N_909,In_616,In_879);
nor U910 (N_910,In_928,In_530);
or U911 (N_911,In_454,In_234);
nor U912 (N_912,In_190,In_213);
xor U913 (N_913,In_138,In_302);
or U914 (N_914,In_898,In_367);
xor U915 (N_915,In_131,In_794);
and U916 (N_916,In_179,In_868);
or U917 (N_917,In_21,In_879);
or U918 (N_918,In_44,In_257);
or U919 (N_919,In_841,In_898);
xor U920 (N_920,In_28,In_284);
nor U921 (N_921,In_415,In_341);
or U922 (N_922,In_747,In_101);
and U923 (N_923,In_724,In_99);
and U924 (N_924,In_138,In_159);
and U925 (N_925,In_344,In_656);
nand U926 (N_926,In_3,In_318);
and U927 (N_927,In_11,In_753);
nand U928 (N_928,In_300,In_983);
xor U929 (N_929,In_680,In_69);
xnor U930 (N_930,In_805,In_510);
xor U931 (N_931,In_973,In_683);
or U932 (N_932,In_486,In_336);
nor U933 (N_933,In_789,In_353);
nand U934 (N_934,In_82,In_212);
nand U935 (N_935,In_725,In_612);
nor U936 (N_936,In_76,In_254);
nand U937 (N_937,In_490,In_581);
xnor U938 (N_938,In_785,In_787);
and U939 (N_939,In_317,In_986);
xnor U940 (N_940,In_652,In_729);
and U941 (N_941,In_67,In_933);
or U942 (N_942,In_931,In_96);
nand U943 (N_943,In_181,In_142);
or U944 (N_944,In_432,In_821);
nand U945 (N_945,In_946,In_672);
and U946 (N_946,In_819,In_207);
nand U947 (N_947,In_527,In_600);
nand U948 (N_948,In_993,In_347);
nor U949 (N_949,In_682,In_784);
and U950 (N_950,In_849,In_298);
or U951 (N_951,In_859,In_997);
xor U952 (N_952,In_219,In_375);
and U953 (N_953,In_257,In_708);
nand U954 (N_954,In_673,In_749);
or U955 (N_955,In_46,In_5);
nor U956 (N_956,In_137,In_999);
xor U957 (N_957,In_574,In_236);
xor U958 (N_958,In_450,In_745);
and U959 (N_959,In_351,In_751);
and U960 (N_960,In_636,In_12);
or U961 (N_961,In_985,In_778);
xnor U962 (N_962,In_61,In_936);
nand U963 (N_963,In_882,In_408);
nand U964 (N_964,In_567,In_352);
and U965 (N_965,In_566,In_725);
or U966 (N_966,In_427,In_149);
xnor U967 (N_967,In_161,In_696);
xor U968 (N_968,In_152,In_652);
or U969 (N_969,In_746,In_717);
or U970 (N_970,In_827,In_848);
and U971 (N_971,In_97,In_907);
or U972 (N_972,In_283,In_323);
or U973 (N_973,In_428,In_710);
nor U974 (N_974,In_492,In_600);
xor U975 (N_975,In_573,In_773);
xor U976 (N_976,In_486,In_4);
and U977 (N_977,In_699,In_888);
and U978 (N_978,In_360,In_276);
nor U979 (N_979,In_429,In_901);
xor U980 (N_980,In_104,In_309);
nor U981 (N_981,In_626,In_172);
and U982 (N_982,In_339,In_422);
and U983 (N_983,In_664,In_953);
and U984 (N_984,In_934,In_464);
nor U985 (N_985,In_65,In_931);
xor U986 (N_986,In_520,In_283);
or U987 (N_987,In_316,In_43);
or U988 (N_988,In_146,In_775);
xor U989 (N_989,In_830,In_768);
and U990 (N_990,In_606,In_247);
nor U991 (N_991,In_462,In_163);
nand U992 (N_992,In_790,In_137);
nor U993 (N_993,In_104,In_143);
or U994 (N_994,In_630,In_671);
xnor U995 (N_995,In_508,In_80);
or U996 (N_996,In_147,In_404);
and U997 (N_997,In_291,In_780);
nor U998 (N_998,In_650,In_329);
or U999 (N_999,In_395,In_602);
and U1000 (N_1000,In_152,In_891);
xnor U1001 (N_1001,In_958,In_181);
or U1002 (N_1002,In_936,In_948);
or U1003 (N_1003,In_446,In_918);
nand U1004 (N_1004,In_359,In_795);
xor U1005 (N_1005,In_971,In_579);
nand U1006 (N_1006,In_858,In_161);
or U1007 (N_1007,In_851,In_341);
nand U1008 (N_1008,In_569,In_306);
and U1009 (N_1009,In_338,In_942);
or U1010 (N_1010,In_425,In_938);
xnor U1011 (N_1011,In_633,In_325);
or U1012 (N_1012,In_874,In_476);
nand U1013 (N_1013,In_856,In_626);
or U1014 (N_1014,In_819,In_583);
and U1015 (N_1015,In_404,In_477);
nand U1016 (N_1016,In_685,In_407);
and U1017 (N_1017,In_555,In_266);
and U1018 (N_1018,In_916,In_163);
nand U1019 (N_1019,In_417,In_681);
or U1020 (N_1020,In_322,In_171);
nand U1021 (N_1021,In_335,In_834);
and U1022 (N_1022,In_266,In_705);
and U1023 (N_1023,In_489,In_944);
xnor U1024 (N_1024,In_628,In_542);
nor U1025 (N_1025,In_723,In_444);
or U1026 (N_1026,In_356,In_151);
or U1027 (N_1027,In_795,In_562);
and U1028 (N_1028,In_428,In_558);
or U1029 (N_1029,In_120,In_643);
nand U1030 (N_1030,In_582,In_754);
and U1031 (N_1031,In_943,In_718);
or U1032 (N_1032,In_876,In_446);
or U1033 (N_1033,In_521,In_785);
xor U1034 (N_1034,In_279,In_127);
and U1035 (N_1035,In_25,In_104);
xnor U1036 (N_1036,In_296,In_920);
xor U1037 (N_1037,In_437,In_732);
or U1038 (N_1038,In_742,In_361);
nand U1039 (N_1039,In_339,In_666);
nand U1040 (N_1040,In_18,In_875);
nor U1041 (N_1041,In_159,In_477);
and U1042 (N_1042,In_217,In_389);
nor U1043 (N_1043,In_587,In_856);
or U1044 (N_1044,In_19,In_204);
and U1045 (N_1045,In_118,In_607);
nand U1046 (N_1046,In_367,In_287);
nand U1047 (N_1047,In_886,In_401);
nor U1048 (N_1048,In_536,In_21);
and U1049 (N_1049,In_871,In_899);
nor U1050 (N_1050,In_656,In_372);
or U1051 (N_1051,In_648,In_203);
nor U1052 (N_1052,In_477,In_397);
or U1053 (N_1053,In_940,In_593);
nor U1054 (N_1054,In_477,In_67);
nor U1055 (N_1055,In_805,In_367);
and U1056 (N_1056,In_241,In_493);
nor U1057 (N_1057,In_777,In_888);
xnor U1058 (N_1058,In_158,In_681);
nand U1059 (N_1059,In_785,In_761);
nor U1060 (N_1060,In_113,In_570);
or U1061 (N_1061,In_145,In_180);
or U1062 (N_1062,In_98,In_471);
and U1063 (N_1063,In_269,In_503);
xnor U1064 (N_1064,In_82,In_725);
and U1065 (N_1065,In_346,In_865);
or U1066 (N_1066,In_746,In_413);
nand U1067 (N_1067,In_980,In_813);
xor U1068 (N_1068,In_203,In_576);
and U1069 (N_1069,In_99,In_544);
nor U1070 (N_1070,In_10,In_379);
nand U1071 (N_1071,In_287,In_421);
nor U1072 (N_1072,In_52,In_924);
nand U1073 (N_1073,In_592,In_111);
and U1074 (N_1074,In_337,In_412);
xnor U1075 (N_1075,In_843,In_483);
or U1076 (N_1076,In_649,In_345);
nor U1077 (N_1077,In_202,In_645);
nor U1078 (N_1078,In_198,In_884);
nor U1079 (N_1079,In_642,In_935);
and U1080 (N_1080,In_268,In_7);
xor U1081 (N_1081,In_202,In_286);
or U1082 (N_1082,In_869,In_99);
or U1083 (N_1083,In_657,In_4);
or U1084 (N_1084,In_390,In_612);
xnor U1085 (N_1085,In_972,In_131);
or U1086 (N_1086,In_792,In_879);
nand U1087 (N_1087,In_394,In_513);
xnor U1088 (N_1088,In_301,In_113);
or U1089 (N_1089,In_165,In_438);
nor U1090 (N_1090,In_187,In_420);
or U1091 (N_1091,In_348,In_704);
nor U1092 (N_1092,In_384,In_729);
xor U1093 (N_1093,In_927,In_120);
and U1094 (N_1094,In_932,In_507);
xor U1095 (N_1095,In_144,In_966);
and U1096 (N_1096,In_844,In_161);
or U1097 (N_1097,In_239,In_789);
and U1098 (N_1098,In_411,In_711);
and U1099 (N_1099,In_402,In_980);
nand U1100 (N_1100,In_395,In_757);
xor U1101 (N_1101,In_169,In_166);
and U1102 (N_1102,In_292,In_711);
nor U1103 (N_1103,In_258,In_115);
nand U1104 (N_1104,In_607,In_247);
and U1105 (N_1105,In_908,In_124);
or U1106 (N_1106,In_749,In_774);
nand U1107 (N_1107,In_848,In_81);
and U1108 (N_1108,In_724,In_902);
xor U1109 (N_1109,In_653,In_571);
nor U1110 (N_1110,In_91,In_508);
xnor U1111 (N_1111,In_606,In_137);
nor U1112 (N_1112,In_6,In_748);
or U1113 (N_1113,In_304,In_245);
and U1114 (N_1114,In_734,In_890);
and U1115 (N_1115,In_893,In_36);
or U1116 (N_1116,In_579,In_883);
or U1117 (N_1117,In_667,In_747);
nor U1118 (N_1118,In_798,In_405);
xnor U1119 (N_1119,In_204,In_961);
nor U1120 (N_1120,In_922,In_563);
nand U1121 (N_1121,In_541,In_137);
and U1122 (N_1122,In_248,In_310);
and U1123 (N_1123,In_457,In_607);
and U1124 (N_1124,In_404,In_225);
or U1125 (N_1125,In_244,In_467);
and U1126 (N_1126,In_390,In_191);
nand U1127 (N_1127,In_468,In_863);
nand U1128 (N_1128,In_742,In_292);
or U1129 (N_1129,In_70,In_60);
or U1130 (N_1130,In_19,In_478);
and U1131 (N_1131,In_697,In_423);
nand U1132 (N_1132,In_149,In_159);
nand U1133 (N_1133,In_661,In_776);
or U1134 (N_1134,In_882,In_383);
nand U1135 (N_1135,In_281,In_769);
xnor U1136 (N_1136,In_235,In_560);
or U1137 (N_1137,In_88,In_519);
xor U1138 (N_1138,In_229,In_659);
nand U1139 (N_1139,In_147,In_30);
and U1140 (N_1140,In_122,In_546);
or U1141 (N_1141,In_931,In_936);
and U1142 (N_1142,In_689,In_746);
nor U1143 (N_1143,In_165,In_857);
and U1144 (N_1144,In_271,In_603);
nor U1145 (N_1145,In_974,In_202);
or U1146 (N_1146,In_50,In_689);
and U1147 (N_1147,In_161,In_578);
and U1148 (N_1148,In_992,In_770);
nor U1149 (N_1149,In_721,In_127);
xor U1150 (N_1150,In_345,In_426);
nand U1151 (N_1151,In_406,In_867);
nand U1152 (N_1152,In_817,In_348);
and U1153 (N_1153,In_706,In_709);
nor U1154 (N_1154,In_584,In_655);
xnor U1155 (N_1155,In_3,In_716);
xnor U1156 (N_1156,In_409,In_319);
nand U1157 (N_1157,In_996,In_298);
nor U1158 (N_1158,In_108,In_551);
nor U1159 (N_1159,In_70,In_394);
xnor U1160 (N_1160,In_677,In_928);
xor U1161 (N_1161,In_352,In_991);
and U1162 (N_1162,In_920,In_136);
nand U1163 (N_1163,In_719,In_315);
nand U1164 (N_1164,In_560,In_6);
or U1165 (N_1165,In_637,In_906);
xor U1166 (N_1166,In_844,In_920);
or U1167 (N_1167,In_478,In_231);
xnor U1168 (N_1168,In_855,In_374);
or U1169 (N_1169,In_319,In_59);
or U1170 (N_1170,In_127,In_739);
nor U1171 (N_1171,In_680,In_169);
nand U1172 (N_1172,In_528,In_526);
or U1173 (N_1173,In_414,In_617);
nand U1174 (N_1174,In_190,In_650);
and U1175 (N_1175,In_749,In_34);
and U1176 (N_1176,In_666,In_735);
nand U1177 (N_1177,In_814,In_828);
or U1178 (N_1178,In_255,In_523);
and U1179 (N_1179,In_880,In_678);
nand U1180 (N_1180,In_732,In_721);
xnor U1181 (N_1181,In_711,In_243);
nand U1182 (N_1182,In_701,In_741);
and U1183 (N_1183,In_433,In_449);
xnor U1184 (N_1184,In_931,In_698);
nand U1185 (N_1185,In_64,In_41);
xor U1186 (N_1186,In_941,In_395);
nand U1187 (N_1187,In_662,In_89);
nand U1188 (N_1188,In_516,In_54);
xor U1189 (N_1189,In_185,In_463);
nor U1190 (N_1190,In_717,In_607);
or U1191 (N_1191,In_578,In_977);
nor U1192 (N_1192,In_442,In_120);
or U1193 (N_1193,In_863,In_191);
and U1194 (N_1194,In_402,In_958);
nand U1195 (N_1195,In_481,In_183);
nor U1196 (N_1196,In_634,In_579);
xor U1197 (N_1197,In_760,In_841);
or U1198 (N_1198,In_886,In_449);
and U1199 (N_1199,In_213,In_82);
and U1200 (N_1200,In_214,In_874);
nand U1201 (N_1201,In_355,In_12);
or U1202 (N_1202,In_850,In_281);
nand U1203 (N_1203,In_117,In_105);
nor U1204 (N_1204,In_401,In_470);
nor U1205 (N_1205,In_685,In_594);
nand U1206 (N_1206,In_137,In_514);
and U1207 (N_1207,In_321,In_134);
and U1208 (N_1208,In_867,In_524);
and U1209 (N_1209,In_308,In_200);
or U1210 (N_1210,In_389,In_608);
or U1211 (N_1211,In_64,In_868);
or U1212 (N_1212,In_751,In_160);
xnor U1213 (N_1213,In_609,In_283);
nand U1214 (N_1214,In_997,In_108);
or U1215 (N_1215,In_197,In_419);
and U1216 (N_1216,In_695,In_838);
nand U1217 (N_1217,In_330,In_421);
nand U1218 (N_1218,In_228,In_822);
or U1219 (N_1219,In_830,In_385);
or U1220 (N_1220,In_705,In_616);
nor U1221 (N_1221,In_663,In_224);
nand U1222 (N_1222,In_508,In_632);
or U1223 (N_1223,In_265,In_856);
xor U1224 (N_1224,In_590,In_589);
and U1225 (N_1225,In_115,In_630);
nor U1226 (N_1226,In_404,In_772);
nor U1227 (N_1227,In_372,In_928);
and U1228 (N_1228,In_979,In_604);
nand U1229 (N_1229,In_418,In_397);
or U1230 (N_1230,In_881,In_616);
or U1231 (N_1231,In_271,In_4);
and U1232 (N_1232,In_410,In_748);
xor U1233 (N_1233,In_988,In_516);
and U1234 (N_1234,In_139,In_653);
or U1235 (N_1235,In_693,In_384);
and U1236 (N_1236,In_692,In_24);
nor U1237 (N_1237,In_842,In_66);
nand U1238 (N_1238,In_385,In_891);
xor U1239 (N_1239,In_912,In_648);
nor U1240 (N_1240,In_352,In_341);
nand U1241 (N_1241,In_921,In_920);
or U1242 (N_1242,In_35,In_610);
and U1243 (N_1243,In_246,In_346);
nor U1244 (N_1244,In_610,In_335);
nor U1245 (N_1245,In_937,In_749);
nand U1246 (N_1246,In_103,In_864);
nand U1247 (N_1247,In_41,In_728);
nand U1248 (N_1248,In_854,In_863);
or U1249 (N_1249,In_366,In_826);
xor U1250 (N_1250,In_241,In_683);
nand U1251 (N_1251,In_646,In_276);
or U1252 (N_1252,In_468,In_303);
nand U1253 (N_1253,In_574,In_159);
nand U1254 (N_1254,In_360,In_643);
and U1255 (N_1255,In_156,In_181);
xnor U1256 (N_1256,In_669,In_236);
or U1257 (N_1257,In_988,In_599);
nand U1258 (N_1258,In_121,In_792);
nor U1259 (N_1259,In_801,In_697);
nand U1260 (N_1260,In_509,In_663);
and U1261 (N_1261,In_530,In_398);
and U1262 (N_1262,In_56,In_696);
and U1263 (N_1263,In_809,In_703);
and U1264 (N_1264,In_33,In_360);
xor U1265 (N_1265,In_887,In_384);
xnor U1266 (N_1266,In_990,In_344);
nand U1267 (N_1267,In_813,In_269);
nand U1268 (N_1268,In_841,In_220);
xnor U1269 (N_1269,In_481,In_418);
nand U1270 (N_1270,In_148,In_732);
nor U1271 (N_1271,In_455,In_245);
xnor U1272 (N_1272,In_298,In_641);
nor U1273 (N_1273,In_601,In_931);
or U1274 (N_1274,In_347,In_991);
nand U1275 (N_1275,In_526,In_826);
or U1276 (N_1276,In_183,In_646);
or U1277 (N_1277,In_595,In_353);
nand U1278 (N_1278,In_940,In_224);
nand U1279 (N_1279,In_46,In_302);
and U1280 (N_1280,In_947,In_977);
and U1281 (N_1281,In_696,In_159);
xnor U1282 (N_1282,In_507,In_636);
and U1283 (N_1283,In_865,In_60);
nand U1284 (N_1284,In_152,In_881);
or U1285 (N_1285,In_59,In_316);
xnor U1286 (N_1286,In_385,In_360);
nor U1287 (N_1287,In_407,In_189);
or U1288 (N_1288,In_552,In_762);
nand U1289 (N_1289,In_563,In_152);
and U1290 (N_1290,In_312,In_637);
and U1291 (N_1291,In_389,In_802);
or U1292 (N_1292,In_969,In_9);
or U1293 (N_1293,In_208,In_817);
or U1294 (N_1294,In_419,In_445);
and U1295 (N_1295,In_832,In_573);
and U1296 (N_1296,In_656,In_809);
nor U1297 (N_1297,In_165,In_615);
or U1298 (N_1298,In_568,In_119);
nor U1299 (N_1299,In_642,In_704);
nand U1300 (N_1300,In_545,In_26);
or U1301 (N_1301,In_207,In_680);
and U1302 (N_1302,In_820,In_757);
or U1303 (N_1303,In_8,In_688);
and U1304 (N_1304,In_39,In_968);
and U1305 (N_1305,In_330,In_280);
and U1306 (N_1306,In_672,In_774);
nand U1307 (N_1307,In_191,In_213);
xnor U1308 (N_1308,In_91,In_544);
or U1309 (N_1309,In_857,In_228);
nand U1310 (N_1310,In_692,In_835);
nand U1311 (N_1311,In_144,In_636);
and U1312 (N_1312,In_156,In_297);
or U1313 (N_1313,In_916,In_937);
or U1314 (N_1314,In_526,In_231);
xnor U1315 (N_1315,In_224,In_712);
or U1316 (N_1316,In_532,In_14);
nor U1317 (N_1317,In_559,In_66);
nand U1318 (N_1318,In_3,In_112);
xnor U1319 (N_1319,In_585,In_539);
nor U1320 (N_1320,In_90,In_437);
nand U1321 (N_1321,In_598,In_18);
nor U1322 (N_1322,In_74,In_875);
nor U1323 (N_1323,In_698,In_883);
and U1324 (N_1324,In_319,In_131);
or U1325 (N_1325,In_828,In_482);
nand U1326 (N_1326,In_762,In_507);
nor U1327 (N_1327,In_276,In_11);
nor U1328 (N_1328,In_189,In_953);
xnor U1329 (N_1329,In_44,In_665);
and U1330 (N_1330,In_287,In_735);
nand U1331 (N_1331,In_223,In_162);
or U1332 (N_1332,In_467,In_490);
nand U1333 (N_1333,In_487,In_227);
or U1334 (N_1334,In_839,In_423);
nand U1335 (N_1335,In_632,In_850);
nor U1336 (N_1336,In_51,In_448);
nand U1337 (N_1337,In_319,In_555);
or U1338 (N_1338,In_664,In_544);
xor U1339 (N_1339,In_180,In_222);
or U1340 (N_1340,In_111,In_450);
nor U1341 (N_1341,In_679,In_612);
and U1342 (N_1342,In_265,In_602);
xor U1343 (N_1343,In_731,In_566);
xnor U1344 (N_1344,In_969,In_524);
nor U1345 (N_1345,In_344,In_978);
and U1346 (N_1346,In_676,In_968);
nand U1347 (N_1347,In_334,In_631);
xor U1348 (N_1348,In_305,In_597);
nor U1349 (N_1349,In_761,In_257);
nor U1350 (N_1350,In_732,In_164);
or U1351 (N_1351,In_180,In_236);
and U1352 (N_1352,In_961,In_104);
xor U1353 (N_1353,In_729,In_462);
nor U1354 (N_1354,In_850,In_489);
and U1355 (N_1355,In_313,In_52);
and U1356 (N_1356,In_315,In_366);
and U1357 (N_1357,In_547,In_773);
nor U1358 (N_1358,In_589,In_946);
or U1359 (N_1359,In_238,In_236);
and U1360 (N_1360,In_33,In_8);
or U1361 (N_1361,In_796,In_535);
nand U1362 (N_1362,In_851,In_335);
nor U1363 (N_1363,In_936,In_529);
nand U1364 (N_1364,In_314,In_96);
and U1365 (N_1365,In_203,In_49);
or U1366 (N_1366,In_134,In_337);
xor U1367 (N_1367,In_354,In_85);
and U1368 (N_1368,In_825,In_636);
and U1369 (N_1369,In_349,In_977);
and U1370 (N_1370,In_185,In_727);
xor U1371 (N_1371,In_101,In_411);
and U1372 (N_1372,In_277,In_489);
nor U1373 (N_1373,In_664,In_31);
nand U1374 (N_1374,In_175,In_861);
or U1375 (N_1375,In_380,In_587);
or U1376 (N_1376,In_622,In_712);
xnor U1377 (N_1377,In_228,In_148);
and U1378 (N_1378,In_306,In_544);
xnor U1379 (N_1379,In_118,In_742);
and U1380 (N_1380,In_836,In_232);
and U1381 (N_1381,In_850,In_420);
xor U1382 (N_1382,In_630,In_134);
nor U1383 (N_1383,In_572,In_733);
and U1384 (N_1384,In_762,In_153);
or U1385 (N_1385,In_911,In_699);
and U1386 (N_1386,In_932,In_95);
nand U1387 (N_1387,In_977,In_18);
nor U1388 (N_1388,In_830,In_123);
or U1389 (N_1389,In_301,In_942);
nor U1390 (N_1390,In_361,In_921);
or U1391 (N_1391,In_496,In_330);
and U1392 (N_1392,In_105,In_989);
nor U1393 (N_1393,In_15,In_692);
xnor U1394 (N_1394,In_588,In_665);
and U1395 (N_1395,In_862,In_322);
or U1396 (N_1396,In_298,In_526);
and U1397 (N_1397,In_168,In_320);
nand U1398 (N_1398,In_529,In_878);
nor U1399 (N_1399,In_66,In_120);
nand U1400 (N_1400,In_930,In_732);
xor U1401 (N_1401,In_323,In_523);
and U1402 (N_1402,In_67,In_614);
and U1403 (N_1403,In_257,In_987);
nand U1404 (N_1404,In_241,In_548);
nand U1405 (N_1405,In_537,In_779);
and U1406 (N_1406,In_513,In_423);
nor U1407 (N_1407,In_120,In_799);
or U1408 (N_1408,In_647,In_602);
or U1409 (N_1409,In_480,In_154);
nor U1410 (N_1410,In_279,In_343);
nand U1411 (N_1411,In_839,In_694);
xor U1412 (N_1412,In_217,In_20);
or U1413 (N_1413,In_498,In_622);
and U1414 (N_1414,In_546,In_132);
xnor U1415 (N_1415,In_302,In_862);
xor U1416 (N_1416,In_611,In_170);
and U1417 (N_1417,In_675,In_430);
and U1418 (N_1418,In_310,In_369);
xnor U1419 (N_1419,In_626,In_876);
nor U1420 (N_1420,In_295,In_722);
nor U1421 (N_1421,In_197,In_464);
nor U1422 (N_1422,In_433,In_597);
nand U1423 (N_1423,In_432,In_650);
and U1424 (N_1424,In_406,In_796);
nand U1425 (N_1425,In_91,In_786);
xnor U1426 (N_1426,In_318,In_265);
and U1427 (N_1427,In_972,In_359);
nand U1428 (N_1428,In_308,In_621);
nand U1429 (N_1429,In_887,In_876);
xnor U1430 (N_1430,In_605,In_99);
and U1431 (N_1431,In_104,In_830);
and U1432 (N_1432,In_161,In_612);
or U1433 (N_1433,In_361,In_182);
nor U1434 (N_1434,In_31,In_635);
xor U1435 (N_1435,In_342,In_629);
and U1436 (N_1436,In_358,In_624);
nor U1437 (N_1437,In_203,In_979);
or U1438 (N_1438,In_880,In_77);
xnor U1439 (N_1439,In_272,In_0);
and U1440 (N_1440,In_219,In_866);
nor U1441 (N_1441,In_702,In_231);
or U1442 (N_1442,In_796,In_914);
nor U1443 (N_1443,In_387,In_234);
and U1444 (N_1444,In_779,In_254);
and U1445 (N_1445,In_723,In_493);
or U1446 (N_1446,In_827,In_834);
and U1447 (N_1447,In_325,In_36);
or U1448 (N_1448,In_356,In_74);
xor U1449 (N_1449,In_280,In_885);
or U1450 (N_1450,In_942,In_306);
and U1451 (N_1451,In_634,In_671);
nand U1452 (N_1452,In_744,In_657);
or U1453 (N_1453,In_805,In_933);
xor U1454 (N_1454,In_273,In_73);
xor U1455 (N_1455,In_289,In_446);
nor U1456 (N_1456,In_251,In_323);
or U1457 (N_1457,In_360,In_5);
xor U1458 (N_1458,In_116,In_651);
and U1459 (N_1459,In_446,In_368);
or U1460 (N_1460,In_324,In_313);
nor U1461 (N_1461,In_837,In_414);
and U1462 (N_1462,In_17,In_628);
or U1463 (N_1463,In_739,In_310);
and U1464 (N_1464,In_270,In_958);
nor U1465 (N_1465,In_374,In_760);
nand U1466 (N_1466,In_644,In_875);
xnor U1467 (N_1467,In_545,In_255);
and U1468 (N_1468,In_780,In_698);
nor U1469 (N_1469,In_716,In_737);
or U1470 (N_1470,In_547,In_906);
xor U1471 (N_1471,In_375,In_535);
and U1472 (N_1472,In_907,In_672);
or U1473 (N_1473,In_935,In_639);
xnor U1474 (N_1474,In_183,In_960);
nor U1475 (N_1475,In_145,In_186);
or U1476 (N_1476,In_854,In_933);
and U1477 (N_1477,In_141,In_840);
and U1478 (N_1478,In_677,In_92);
nand U1479 (N_1479,In_772,In_398);
or U1480 (N_1480,In_602,In_515);
or U1481 (N_1481,In_50,In_565);
or U1482 (N_1482,In_20,In_779);
or U1483 (N_1483,In_844,In_712);
and U1484 (N_1484,In_917,In_334);
and U1485 (N_1485,In_608,In_9);
xor U1486 (N_1486,In_44,In_233);
nor U1487 (N_1487,In_170,In_483);
and U1488 (N_1488,In_723,In_383);
xnor U1489 (N_1489,In_106,In_889);
xor U1490 (N_1490,In_883,In_923);
or U1491 (N_1491,In_578,In_266);
nand U1492 (N_1492,In_428,In_358);
nand U1493 (N_1493,In_945,In_668);
or U1494 (N_1494,In_545,In_372);
xor U1495 (N_1495,In_708,In_111);
or U1496 (N_1496,In_780,In_351);
or U1497 (N_1497,In_656,In_551);
xor U1498 (N_1498,In_580,In_980);
nand U1499 (N_1499,In_191,In_552);
nand U1500 (N_1500,In_499,In_11);
and U1501 (N_1501,In_983,In_963);
and U1502 (N_1502,In_627,In_283);
and U1503 (N_1503,In_737,In_581);
nor U1504 (N_1504,In_264,In_790);
nand U1505 (N_1505,In_12,In_581);
xnor U1506 (N_1506,In_410,In_185);
xor U1507 (N_1507,In_369,In_53);
xor U1508 (N_1508,In_541,In_756);
nor U1509 (N_1509,In_552,In_77);
xor U1510 (N_1510,In_101,In_758);
nand U1511 (N_1511,In_727,In_681);
nor U1512 (N_1512,In_397,In_805);
or U1513 (N_1513,In_226,In_275);
and U1514 (N_1514,In_765,In_391);
or U1515 (N_1515,In_210,In_258);
nand U1516 (N_1516,In_57,In_9);
nor U1517 (N_1517,In_788,In_488);
and U1518 (N_1518,In_250,In_999);
nor U1519 (N_1519,In_104,In_218);
and U1520 (N_1520,In_94,In_526);
nor U1521 (N_1521,In_744,In_185);
xnor U1522 (N_1522,In_322,In_181);
nand U1523 (N_1523,In_550,In_260);
or U1524 (N_1524,In_121,In_326);
and U1525 (N_1525,In_705,In_422);
nor U1526 (N_1526,In_1,In_785);
and U1527 (N_1527,In_430,In_311);
or U1528 (N_1528,In_219,In_334);
nor U1529 (N_1529,In_393,In_899);
xnor U1530 (N_1530,In_113,In_231);
xnor U1531 (N_1531,In_760,In_819);
or U1532 (N_1532,In_953,In_923);
xnor U1533 (N_1533,In_38,In_889);
and U1534 (N_1534,In_994,In_704);
nand U1535 (N_1535,In_120,In_234);
and U1536 (N_1536,In_223,In_732);
and U1537 (N_1537,In_906,In_45);
or U1538 (N_1538,In_620,In_600);
xor U1539 (N_1539,In_752,In_699);
nand U1540 (N_1540,In_88,In_674);
nand U1541 (N_1541,In_138,In_503);
and U1542 (N_1542,In_0,In_993);
or U1543 (N_1543,In_118,In_379);
nand U1544 (N_1544,In_574,In_209);
or U1545 (N_1545,In_550,In_40);
and U1546 (N_1546,In_927,In_411);
or U1547 (N_1547,In_397,In_262);
nor U1548 (N_1548,In_228,In_526);
xnor U1549 (N_1549,In_604,In_591);
nor U1550 (N_1550,In_399,In_477);
nor U1551 (N_1551,In_757,In_910);
or U1552 (N_1552,In_529,In_263);
nor U1553 (N_1553,In_199,In_739);
nand U1554 (N_1554,In_477,In_48);
nor U1555 (N_1555,In_331,In_687);
or U1556 (N_1556,In_473,In_435);
nor U1557 (N_1557,In_412,In_18);
xnor U1558 (N_1558,In_188,In_688);
or U1559 (N_1559,In_870,In_12);
nand U1560 (N_1560,In_952,In_829);
xnor U1561 (N_1561,In_694,In_116);
and U1562 (N_1562,In_780,In_317);
nor U1563 (N_1563,In_606,In_852);
or U1564 (N_1564,In_664,In_995);
xnor U1565 (N_1565,In_102,In_202);
nor U1566 (N_1566,In_93,In_788);
and U1567 (N_1567,In_477,In_228);
nand U1568 (N_1568,In_485,In_668);
nor U1569 (N_1569,In_182,In_789);
or U1570 (N_1570,In_31,In_914);
or U1571 (N_1571,In_300,In_236);
and U1572 (N_1572,In_344,In_700);
xnor U1573 (N_1573,In_190,In_889);
and U1574 (N_1574,In_314,In_363);
nand U1575 (N_1575,In_703,In_540);
or U1576 (N_1576,In_350,In_616);
and U1577 (N_1577,In_580,In_107);
xnor U1578 (N_1578,In_624,In_866);
nand U1579 (N_1579,In_727,In_275);
or U1580 (N_1580,In_903,In_131);
nand U1581 (N_1581,In_180,In_451);
or U1582 (N_1582,In_480,In_296);
nor U1583 (N_1583,In_215,In_517);
nor U1584 (N_1584,In_556,In_570);
nand U1585 (N_1585,In_463,In_524);
nor U1586 (N_1586,In_401,In_108);
nand U1587 (N_1587,In_845,In_809);
nand U1588 (N_1588,In_785,In_139);
nor U1589 (N_1589,In_421,In_385);
nand U1590 (N_1590,In_369,In_945);
and U1591 (N_1591,In_907,In_385);
nand U1592 (N_1592,In_480,In_644);
or U1593 (N_1593,In_575,In_98);
nor U1594 (N_1594,In_366,In_188);
or U1595 (N_1595,In_475,In_403);
nor U1596 (N_1596,In_196,In_807);
or U1597 (N_1597,In_802,In_479);
nand U1598 (N_1598,In_452,In_75);
xnor U1599 (N_1599,In_397,In_373);
or U1600 (N_1600,In_360,In_959);
xnor U1601 (N_1601,In_945,In_923);
xnor U1602 (N_1602,In_503,In_60);
nand U1603 (N_1603,In_299,In_951);
or U1604 (N_1604,In_647,In_58);
nand U1605 (N_1605,In_207,In_85);
nor U1606 (N_1606,In_711,In_441);
nand U1607 (N_1607,In_292,In_995);
and U1608 (N_1608,In_517,In_144);
or U1609 (N_1609,In_379,In_111);
or U1610 (N_1610,In_677,In_355);
nand U1611 (N_1611,In_818,In_819);
and U1612 (N_1612,In_853,In_808);
nand U1613 (N_1613,In_687,In_99);
and U1614 (N_1614,In_967,In_0);
nor U1615 (N_1615,In_923,In_832);
and U1616 (N_1616,In_908,In_570);
xor U1617 (N_1617,In_553,In_96);
or U1618 (N_1618,In_23,In_786);
xor U1619 (N_1619,In_49,In_822);
nor U1620 (N_1620,In_128,In_260);
or U1621 (N_1621,In_829,In_981);
nor U1622 (N_1622,In_334,In_303);
xor U1623 (N_1623,In_423,In_419);
or U1624 (N_1624,In_343,In_820);
or U1625 (N_1625,In_728,In_589);
nand U1626 (N_1626,In_791,In_438);
and U1627 (N_1627,In_698,In_22);
or U1628 (N_1628,In_505,In_945);
and U1629 (N_1629,In_953,In_597);
or U1630 (N_1630,In_171,In_947);
nand U1631 (N_1631,In_159,In_590);
or U1632 (N_1632,In_41,In_285);
and U1633 (N_1633,In_40,In_314);
or U1634 (N_1634,In_905,In_362);
and U1635 (N_1635,In_542,In_209);
or U1636 (N_1636,In_355,In_161);
nand U1637 (N_1637,In_607,In_704);
xor U1638 (N_1638,In_153,In_714);
nand U1639 (N_1639,In_815,In_395);
xnor U1640 (N_1640,In_916,In_756);
or U1641 (N_1641,In_897,In_275);
xnor U1642 (N_1642,In_766,In_834);
nor U1643 (N_1643,In_408,In_338);
nand U1644 (N_1644,In_227,In_68);
and U1645 (N_1645,In_183,In_386);
or U1646 (N_1646,In_819,In_424);
nor U1647 (N_1647,In_179,In_16);
or U1648 (N_1648,In_79,In_85);
or U1649 (N_1649,In_769,In_117);
nand U1650 (N_1650,In_937,In_409);
xnor U1651 (N_1651,In_409,In_942);
xor U1652 (N_1652,In_318,In_763);
xnor U1653 (N_1653,In_261,In_57);
or U1654 (N_1654,In_895,In_648);
xor U1655 (N_1655,In_209,In_837);
nand U1656 (N_1656,In_899,In_632);
xor U1657 (N_1657,In_431,In_132);
and U1658 (N_1658,In_111,In_711);
and U1659 (N_1659,In_458,In_388);
xor U1660 (N_1660,In_163,In_720);
xnor U1661 (N_1661,In_0,In_588);
or U1662 (N_1662,In_982,In_647);
xor U1663 (N_1663,In_873,In_349);
nor U1664 (N_1664,In_63,In_729);
and U1665 (N_1665,In_301,In_112);
nor U1666 (N_1666,In_356,In_645);
and U1667 (N_1667,In_220,In_384);
or U1668 (N_1668,In_175,In_155);
or U1669 (N_1669,In_747,In_165);
nand U1670 (N_1670,In_700,In_261);
and U1671 (N_1671,In_182,In_120);
nor U1672 (N_1672,In_190,In_318);
or U1673 (N_1673,In_112,In_740);
and U1674 (N_1674,In_478,In_552);
and U1675 (N_1675,In_560,In_483);
or U1676 (N_1676,In_507,In_768);
xnor U1677 (N_1677,In_69,In_212);
and U1678 (N_1678,In_553,In_315);
nand U1679 (N_1679,In_957,In_571);
or U1680 (N_1680,In_103,In_95);
and U1681 (N_1681,In_455,In_586);
xnor U1682 (N_1682,In_62,In_196);
nand U1683 (N_1683,In_563,In_791);
xnor U1684 (N_1684,In_744,In_334);
and U1685 (N_1685,In_532,In_575);
xnor U1686 (N_1686,In_894,In_966);
or U1687 (N_1687,In_618,In_227);
nor U1688 (N_1688,In_50,In_701);
or U1689 (N_1689,In_709,In_927);
or U1690 (N_1690,In_531,In_910);
nor U1691 (N_1691,In_433,In_979);
nor U1692 (N_1692,In_106,In_667);
xor U1693 (N_1693,In_48,In_198);
or U1694 (N_1694,In_86,In_604);
nor U1695 (N_1695,In_685,In_445);
xor U1696 (N_1696,In_958,In_539);
or U1697 (N_1697,In_648,In_745);
nand U1698 (N_1698,In_74,In_617);
xnor U1699 (N_1699,In_2,In_981);
xor U1700 (N_1700,In_447,In_709);
and U1701 (N_1701,In_342,In_159);
and U1702 (N_1702,In_54,In_777);
xor U1703 (N_1703,In_250,In_515);
nor U1704 (N_1704,In_468,In_256);
or U1705 (N_1705,In_807,In_491);
nor U1706 (N_1706,In_366,In_464);
or U1707 (N_1707,In_301,In_745);
nor U1708 (N_1708,In_420,In_671);
xor U1709 (N_1709,In_815,In_887);
nor U1710 (N_1710,In_617,In_939);
and U1711 (N_1711,In_384,In_301);
nor U1712 (N_1712,In_526,In_23);
nand U1713 (N_1713,In_780,In_712);
xor U1714 (N_1714,In_603,In_871);
and U1715 (N_1715,In_514,In_808);
xnor U1716 (N_1716,In_964,In_129);
nand U1717 (N_1717,In_531,In_908);
nand U1718 (N_1718,In_842,In_726);
and U1719 (N_1719,In_486,In_22);
or U1720 (N_1720,In_332,In_232);
nand U1721 (N_1721,In_253,In_939);
nand U1722 (N_1722,In_60,In_841);
and U1723 (N_1723,In_580,In_146);
and U1724 (N_1724,In_836,In_343);
nand U1725 (N_1725,In_939,In_648);
nor U1726 (N_1726,In_493,In_561);
and U1727 (N_1727,In_632,In_947);
nand U1728 (N_1728,In_50,In_323);
xor U1729 (N_1729,In_199,In_279);
or U1730 (N_1730,In_605,In_610);
nand U1731 (N_1731,In_215,In_904);
xor U1732 (N_1732,In_236,In_487);
and U1733 (N_1733,In_60,In_609);
and U1734 (N_1734,In_988,In_608);
nand U1735 (N_1735,In_957,In_761);
nand U1736 (N_1736,In_909,In_21);
and U1737 (N_1737,In_432,In_17);
or U1738 (N_1738,In_502,In_145);
nand U1739 (N_1739,In_686,In_471);
nor U1740 (N_1740,In_116,In_124);
nand U1741 (N_1741,In_894,In_62);
and U1742 (N_1742,In_157,In_87);
nor U1743 (N_1743,In_176,In_664);
nor U1744 (N_1744,In_212,In_161);
and U1745 (N_1745,In_51,In_158);
nor U1746 (N_1746,In_22,In_406);
and U1747 (N_1747,In_562,In_312);
or U1748 (N_1748,In_857,In_518);
nand U1749 (N_1749,In_986,In_315);
nor U1750 (N_1750,In_56,In_510);
and U1751 (N_1751,In_959,In_626);
and U1752 (N_1752,In_254,In_80);
nor U1753 (N_1753,In_763,In_572);
or U1754 (N_1754,In_843,In_63);
nor U1755 (N_1755,In_87,In_480);
xnor U1756 (N_1756,In_967,In_977);
and U1757 (N_1757,In_766,In_560);
or U1758 (N_1758,In_843,In_837);
and U1759 (N_1759,In_916,In_824);
or U1760 (N_1760,In_468,In_914);
or U1761 (N_1761,In_115,In_743);
nor U1762 (N_1762,In_859,In_631);
or U1763 (N_1763,In_172,In_604);
xnor U1764 (N_1764,In_812,In_234);
xor U1765 (N_1765,In_342,In_471);
nand U1766 (N_1766,In_259,In_491);
xnor U1767 (N_1767,In_405,In_468);
nor U1768 (N_1768,In_369,In_244);
or U1769 (N_1769,In_861,In_785);
xor U1770 (N_1770,In_984,In_277);
nor U1771 (N_1771,In_564,In_754);
nor U1772 (N_1772,In_925,In_367);
nand U1773 (N_1773,In_55,In_297);
xor U1774 (N_1774,In_571,In_549);
nand U1775 (N_1775,In_138,In_739);
nand U1776 (N_1776,In_701,In_833);
and U1777 (N_1777,In_927,In_107);
xor U1778 (N_1778,In_859,In_273);
nor U1779 (N_1779,In_777,In_174);
or U1780 (N_1780,In_804,In_578);
nor U1781 (N_1781,In_993,In_33);
or U1782 (N_1782,In_876,In_151);
nand U1783 (N_1783,In_346,In_690);
nand U1784 (N_1784,In_439,In_807);
xnor U1785 (N_1785,In_769,In_878);
and U1786 (N_1786,In_335,In_410);
or U1787 (N_1787,In_57,In_817);
and U1788 (N_1788,In_865,In_345);
nand U1789 (N_1789,In_316,In_437);
nand U1790 (N_1790,In_934,In_693);
or U1791 (N_1791,In_467,In_288);
nor U1792 (N_1792,In_417,In_721);
nor U1793 (N_1793,In_497,In_288);
xnor U1794 (N_1794,In_977,In_612);
and U1795 (N_1795,In_790,In_964);
nor U1796 (N_1796,In_808,In_377);
nor U1797 (N_1797,In_535,In_355);
nor U1798 (N_1798,In_146,In_425);
xor U1799 (N_1799,In_1,In_620);
nand U1800 (N_1800,In_320,In_906);
xnor U1801 (N_1801,In_132,In_923);
xnor U1802 (N_1802,In_446,In_440);
xor U1803 (N_1803,In_428,In_380);
or U1804 (N_1804,In_611,In_567);
and U1805 (N_1805,In_202,In_21);
or U1806 (N_1806,In_1,In_115);
and U1807 (N_1807,In_955,In_387);
nand U1808 (N_1808,In_990,In_342);
xnor U1809 (N_1809,In_513,In_665);
nor U1810 (N_1810,In_576,In_18);
and U1811 (N_1811,In_56,In_26);
xnor U1812 (N_1812,In_106,In_188);
nand U1813 (N_1813,In_582,In_182);
or U1814 (N_1814,In_114,In_427);
or U1815 (N_1815,In_547,In_950);
or U1816 (N_1816,In_689,In_645);
nor U1817 (N_1817,In_383,In_55);
nand U1818 (N_1818,In_330,In_550);
nand U1819 (N_1819,In_380,In_402);
and U1820 (N_1820,In_404,In_507);
nor U1821 (N_1821,In_228,In_154);
and U1822 (N_1822,In_516,In_867);
xnor U1823 (N_1823,In_196,In_302);
or U1824 (N_1824,In_622,In_990);
nor U1825 (N_1825,In_12,In_534);
nor U1826 (N_1826,In_2,In_968);
or U1827 (N_1827,In_221,In_857);
nor U1828 (N_1828,In_914,In_266);
or U1829 (N_1829,In_770,In_123);
or U1830 (N_1830,In_713,In_1);
and U1831 (N_1831,In_225,In_908);
nand U1832 (N_1832,In_134,In_597);
and U1833 (N_1833,In_983,In_115);
and U1834 (N_1834,In_586,In_115);
or U1835 (N_1835,In_156,In_428);
xnor U1836 (N_1836,In_817,In_667);
xor U1837 (N_1837,In_555,In_947);
and U1838 (N_1838,In_525,In_353);
and U1839 (N_1839,In_103,In_433);
nor U1840 (N_1840,In_669,In_504);
nor U1841 (N_1841,In_780,In_133);
or U1842 (N_1842,In_834,In_174);
or U1843 (N_1843,In_351,In_864);
nor U1844 (N_1844,In_774,In_15);
and U1845 (N_1845,In_957,In_719);
and U1846 (N_1846,In_446,In_80);
and U1847 (N_1847,In_890,In_680);
xnor U1848 (N_1848,In_503,In_529);
nor U1849 (N_1849,In_195,In_795);
xnor U1850 (N_1850,In_226,In_970);
and U1851 (N_1851,In_226,In_331);
nor U1852 (N_1852,In_991,In_52);
nor U1853 (N_1853,In_796,In_414);
and U1854 (N_1854,In_994,In_661);
or U1855 (N_1855,In_101,In_8);
and U1856 (N_1856,In_573,In_392);
nand U1857 (N_1857,In_898,In_705);
or U1858 (N_1858,In_861,In_626);
xor U1859 (N_1859,In_105,In_52);
nand U1860 (N_1860,In_129,In_344);
or U1861 (N_1861,In_701,In_629);
nand U1862 (N_1862,In_172,In_907);
nand U1863 (N_1863,In_612,In_157);
nand U1864 (N_1864,In_865,In_925);
or U1865 (N_1865,In_538,In_209);
or U1866 (N_1866,In_746,In_613);
and U1867 (N_1867,In_692,In_478);
xnor U1868 (N_1868,In_800,In_988);
xnor U1869 (N_1869,In_813,In_589);
and U1870 (N_1870,In_872,In_196);
nand U1871 (N_1871,In_375,In_221);
and U1872 (N_1872,In_145,In_234);
nor U1873 (N_1873,In_799,In_952);
xor U1874 (N_1874,In_537,In_879);
or U1875 (N_1875,In_69,In_905);
and U1876 (N_1876,In_960,In_754);
or U1877 (N_1877,In_350,In_737);
nor U1878 (N_1878,In_289,In_514);
nor U1879 (N_1879,In_27,In_336);
xnor U1880 (N_1880,In_785,In_342);
nand U1881 (N_1881,In_352,In_722);
xor U1882 (N_1882,In_483,In_736);
or U1883 (N_1883,In_830,In_380);
nand U1884 (N_1884,In_802,In_983);
nor U1885 (N_1885,In_77,In_698);
nand U1886 (N_1886,In_112,In_598);
xnor U1887 (N_1887,In_789,In_600);
or U1888 (N_1888,In_61,In_348);
nor U1889 (N_1889,In_703,In_727);
xor U1890 (N_1890,In_794,In_556);
and U1891 (N_1891,In_100,In_342);
nand U1892 (N_1892,In_16,In_898);
and U1893 (N_1893,In_356,In_91);
xor U1894 (N_1894,In_629,In_240);
xnor U1895 (N_1895,In_484,In_995);
and U1896 (N_1896,In_155,In_228);
nand U1897 (N_1897,In_75,In_272);
nand U1898 (N_1898,In_351,In_11);
xor U1899 (N_1899,In_929,In_797);
and U1900 (N_1900,In_50,In_92);
xor U1901 (N_1901,In_55,In_673);
and U1902 (N_1902,In_428,In_678);
or U1903 (N_1903,In_395,In_605);
and U1904 (N_1904,In_24,In_689);
xnor U1905 (N_1905,In_90,In_257);
or U1906 (N_1906,In_970,In_185);
nand U1907 (N_1907,In_160,In_299);
and U1908 (N_1908,In_116,In_816);
xnor U1909 (N_1909,In_515,In_484);
and U1910 (N_1910,In_309,In_20);
nor U1911 (N_1911,In_546,In_660);
and U1912 (N_1912,In_284,In_63);
and U1913 (N_1913,In_589,In_125);
xor U1914 (N_1914,In_783,In_570);
xor U1915 (N_1915,In_273,In_660);
or U1916 (N_1916,In_87,In_70);
nand U1917 (N_1917,In_586,In_958);
xor U1918 (N_1918,In_934,In_475);
nor U1919 (N_1919,In_334,In_435);
nand U1920 (N_1920,In_537,In_970);
and U1921 (N_1921,In_239,In_966);
xor U1922 (N_1922,In_783,In_493);
and U1923 (N_1923,In_25,In_314);
nor U1924 (N_1924,In_252,In_879);
nand U1925 (N_1925,In_872,In_569);
and U1926 (N_1926,In_672,In_89);
or U1927 (N_1927,In_391,In_117);
or U1928 (N_1928,In_894,In_823);
or U1929 (N_1929,In_324,In_555);
and U1930 (N_1930,In_279,In_513);
nor U1931 (N_1931,In_165,In_274);
and U1932 (N_1932,In_788,In_355);
nor U1933 (N_1933,In_141,In_462);
or U1934 (N_1934,In_922,In_986);
xnor U1935 (N_1935,In_892,In_766);
xnor U1936 (N_1936,In_32,In_798);
nor U1937 (N_1937,In_588,In_461);
and U1938 (N_1938,In_927,In_707);
nand U1939 (N_1939,In_993,In_468);
or U1940 (N_1940,In_283,In_225);
nor U1941 (N_1941,In_156,In_625);
nand U1942 (N_1942,In_529,In_550);
nand U1943 (N_1943,In_639,In_159);
nor U1944 (N_1944,In_581,In_909);
nand U1945 (N_1945,In_61,In_201);
xnor U1946 (N_1946,In_221,In_144);
nand U1947 (N_1947,In_875,In_308);
xor U1948 (N_1948,In_186,In_918);
and U1949 (N_1949,In_726,In_685);
nor U1950 (N_1950,In_776,In_925);
nand U1951 (N_1951,In_841,In_940);
nor U1952 (N_1952,In_35,In_809);
and U1953 (N_1953,In_665,In_240);
or U1954 (N_1954,In_916,In_424);
nor U1955 (N_1955,In_665,In_809);
nand U1956 (N_1956,In_975,In_847);
nor U1957 (N_1957,In_56,In_656);
nand U1958 (N_1958,In_363,In_736);
and U1959 (N_1959,In_811,In_110);
nor U1960 (N_1960,In_150,In_412);
nand U1961 (N_1961,In_896,In_430);
and U1962 (N_1962,In_61,In_864);
xor U1963 (N_1963,In_237,In_585);
nor U1964 (N_1964,In_900,In_686);
or U1965 (N_1965,In_268,In_985);
nor U1966 (N_1966,In_333,In_823);
and U1967 (N_1967,In_860,In_48);
nor U1968 (N_1968,In_610,In_415);
nand U1969 (N_1969,In_789,In_843);
and U1970 (N_1970,In_472,In_483);
nand U1971 (N_1971,In_902,In_584);
xor U1972 (N_1972,In_137,In_993);
or U1973 (N_1973,In_486,In_917);
and U1974 (N_1974,In_667,In_840);
and U1975 (N_1975,In_937,In_628);
and U1976 (N_1976,In_858,In_231);
xnor U1977 (N_1977,In_253,In_431);
xor U1978 (N_1978,In_255,In_899);
xor U1979 (N_1979,In_366,In_425);
or U1980 (N_1980,In_221,In_692);
or U1981 (N_1981,In_193,In_920);
nand U1982 (N_1982,In_979,In_743);
nand U1983 (N_1983,In_51,In_793);
or U1984 (N_1984,In_941,In_811);
and U1985 (N_1985,In_601,In_690);
xor U1986 (N_1986,In_148,In_888);
nand U1987 (N_1987,In_837,In_310);
nand U1988 (N_1988,In_103,In_589);
and U1989 (N_1989,In_541,In_491);
or U1990 (N_1990,In_103,In_163);
and U1991 (N_1991,In_536,In_564);
nand U1992 (N_1992,In_649,In_650);
xor U1993 (N_1993,In_80,In_900);
xnor U1994 (N_1994,In_370,In_467);
or U1995 (N_1995,In_237,In_437);
nor U1996 (N_1996,In_245,In_380);
and U1997 (N_1997,In_62,In_830);
or U1998 (N_1998,In_774,In_333);
or U1999 (N_1999,In_456,In_138);
or U2000 (N_2000,In_53,In_618);
nand U2001 (N_2001,In_163,In_673);
xnor U2002 (N_2002,In_278,In_901);
and U2003 (N_2003,In_797,In_452);
nor U2004 (N_2004,In_505,In_187);
nand U2005 (N_2005,In_722,In_60);
or U2006 (N_2006,In_924,In_276);
or U2007 (N_2007,In_642,In_368);
or U2008 (N_2008,In_967,In_135);
or U2009 (N_2009,In_298,In_726);
nand U2010 (N_2010,In_52,In_230);
nor U2011 (N_2011,In_368,In_109);
xnor U2012 (N_2012,In_648,In_933);
nor U2013 (N_2013,In_147,In_465);
xnor U2014 (N_2014,In_784,In_515);
and U2015 (N_2015,In_150,In_23);
and U2016 (N_2016,In_262,In_687);
and U2017 (N_2017,In_357,In_185);
and U2018 (N_2018,In_329,In_780);
or U2019 (N_2019,In_645,In_849);
nand U2020 (N_2020,In_641,In_254);
xor U2021 (N_2021,In_977,In_674);
or U2022 (N_2022,In_988,In_486);
and U2023 (N_2023,In_611,In_98);
nor U2024 (N_2024,In_683,In_254);
nand U2025 (N_2025,In_175,In_285);
or U2026 (N_2026,In_745,In_468);
nor U2027 (N_2027,In_904,In_138);
nor U2028 (N_2028,In_167,In_811);
xnor U2029 (N_2029,In_320,In_232);
xnor U2030 (N_2030,In_991,In_418);
nor U2031 (N_2031,In_98,In_383);
nor U2032 (N_2032,In_819,In_290);
nor U2033 (N_2033,In_419,In_31);
and U2034 (N_2034,In_189,In_220);
nand U2035 (N_2035,In_316,In_201);
and U2036 (N_2036,In_396,In_993);
xor U2037 (N_2037,In_318,In_154);
xnor U2038 (N_2038,In_125,In_630);
xnor U2039 (N_2039,In_725,In_968);
and U2040 (N_2040,In_357,In_210);
xor U2041 (N_2041,In_414,In_263);
nor U2042 (N_2042,In_790,In_433);
nor U2043 (N_2043,In_131,In_419);
and U2044 (N_2044,In_104,In_873);
or U2045 (N_2045,In_986,In_144);
nor U2046 (N_2046,In_369,In_75);
nand U2047 (N_2047,In_400,In_808);
nand U2048 (N_2048,In_358,In_798);
nand U2049 (N_2049,In_960,In_752);
or U2050 (N_2050,In_423,In_969);
or U2051 (N_2051,In_275,In_403);
and U2052 (N_2052,In_219,In_441);
nor U2053 (N_2053,In_571,In_200);
nor U2054 (N_2054,In_566,In_74);
nor U2055 (N_2055,In_976,In_445);
or U2056 (N_2056,In_327,In_834);
and U2057 (N_2057,In_355,In_533);
xor U2058 (N_2058,In_581,In_880);
nand U2059 (N_2059,In_949,In_416);
xor U2060 (N_2060,In_48,In_952);
nand U2061 (N_2061,In_327,In_945);
and U2062 (N_2062,In_949,In_751);
and U2063 (N_2063,In_168,In_667);
or U2064 (N_2064,In_662,In_839);
nand U2065 (N_2065,In_728,In_717);
nand U2066 (N_2066,In_994,In_586);
and U2067 (N_2067,In_278,In_634);
and U2068 (N_2068,In_783,In_961);
and U2069 (N_2069,In_682,In_146);
xor U2070 (N_2070,In_347,In_564);
xnor U2071 (N_2071,In_762,In_161);
nor U2072 (N_2072,In_595,In_347);
nor U2073 (N_2073,In_140,In_130);
and U2074 (N_2074,In_570,In_59);
xnor U2075 (N_2075,In_183,In_178);
and U2076 (N_2076,In_580,In_419);
or U2077 (N_2077,In_112,In_326);
and U2078 (N_2078,In_430,In_904);
nand U2079 (N_2079,In_963,In_117);
xor U2080 (N_2080,In_181,In_7);
or U2081 (N_2081,In_772,In_136);
xnor U2082 (N_2082,In_340,In_738);
xor U2083 (N_2083,In_558,In_62);
and U2084 (N_2084,In_3,In_688);
xor U2085 (N_2085,In_423,In_977);
nand U2086 (N_2086,In_615,In_270);
xor U2087 (N_2087,In_31,In_332);
or U2088 (N_2088,In_700,In_92);
or U2089 (N_2089,In_665,In_54);
nor U2090 (N_2090,In_672,In_926);
xnor U2091 (N_2091,In_580,In_232);
nand U2092 (N_2092,In_685,In_978);
or U2093 (N_2093,In_406,In_348);
and U2094 (N_2094,In_49,In_318);
xnor U2095 (N_2095,In_877,In_499);
and U2096 (N_2096,In_925,In_127);
or U2097 (N_2097,In_358,In_671);
xor U2098 (N_2098,In_269,In_496);
xnor U2099 (N_2099,In_807,In_809);
nor U2100 (N_2100,In_757,In_89);
or U2101 (N_2101,In_614,In_980);
nor U2102 (N_2102,In_18,In_617);
and U2103 (N_2103,In_144,In_422);
nand U2104 (N_2104,In_745,In_871);
xor U2105 (N_2105,In_155,In_59);
nand U2106 (N_2106,In_579,In_256);
nand U2107 (N_2107,In_632,In_939);
xor U2108 (N_2108,In_764,In_684);
and U2109 (N_2109,In_696,In_657);
nand U2110 (N_2110,In_170,In_174);
nor U2111 (N_2111,In_58,In_626);
and U2112 (N_2112,In_982,In_739);
or U2113 (N_2113,In_366,In_87);
or U2114 (N_2114,In_766,In_549);
xnor U2115 (N_2115,In_113,In_832);
xnor U2116 (N_2116,In_653,In_647);
or U2117 (N_2117,In_86,In_660);
nor U2118 (N_2118,In_406,In_598);
nand U2119 (N_2119,In_589,In_803);
xor U2120 (N_2120,In_9,In_919);
xnor U2121 (N_2121,In_310,In_469);
xnor U2122 (N_2122,In_599,In_397);
or U2123 (N_2123,In_493,In_26);
nor U2124 (N_2124,In_291,In_779);
and U2125 (N_2125,In_224,In_33);
or U2126 (N_2126,In_765,In_670);
xor U2127 (N_2127,In_583,In_960);
nand U2128 (N_2128,In_701,In_403);
nand U2129 (N_2129,In_940,In_344);
nor U2130 (N_2130,In_611,In_75);
or U2131 (N_2131,In_578,In_467);
nor U2132 (N_2132,In_438,In_889);
nand U2133 (N_2133,In_44,In_60);
or U2134 (N_2134,In_131,In_469);
or U2135 (N_2135,In_603,In_869);
nand U2136 (N_2136,In_72,In_585);
or U2137 (N_2137,In_682,In_575);
nor U2138 (N_2138,In_99,In_17);
or U2139 (N_2139,In_223,In_918);
or U2140 (N_2140,In_387,In_4);
or U2141 (N_2141,In_138,In_379);
xor U2142 (N_2142,In_71,In_896);
nor U2143 (N_2143,In_578,In_696);
or U2144 (N_2144,In_575,In_862);
and U2145 (N_2145,In_258,In_616);
nor U2146 (N_2146,In_886,In_801);
nor U2147 (N_2147,In_742,In_818);
nor U2148 (N_2148,In_265,In_827);
nor U2149 (N_2149,In_307,In_450);
or U2150 (N_2150,In_515,In_175);
and U2151 (N_2151,In_785,In_175);
nor U2152 (N_2152,In_891,In_903);
xor U2153 (N_2153,In_35,In_181);
nor U2154 (N_2154,In_522,In_869);
nand U2155 (N_2155,In_838,In_430);
or U2156 (N_2156,In_755,In_551);
xor U2157 (N_2157,In_588,In_81);
nand U2158 (N_2158,In_680,In_847);
xnor U2159 (N_2159,In_216,In_920);
xnor U2160 (N_2160,In_44,In_173);
nor U2161 (N_2161,In_464,In_953);
xor U2162 (N_2162,In_478,In_215);
xor U2163 (N_2163,In_533,In_364);
and U2164 (N_2164,In_737,In_58);
nor U2165 (N_2165,In_849,In_520);
nand U2166 (N_2166,In_912,In_373);
nor U2167 (N_2167,In_112,In_876);
and U2168 (N_2168,In_418,In_631);
nand U2169 (N_2169,In_933,In_807);
xor U2170 (N_2170,In_823,In_292);
nand U2171 (N_2171,In_332,In_918);
or U2172 (N_2172,In_354,In_721);
nand U2173 (N_2173,In_503,In_408);
nor U2174 (N_2174,In_932,In_40);
or U2175 (N_2175,In_477,In_577);
xnor U2176 (N_2176,In_734,In_709);
nor U2177 (N_2177,In_82,In_941);
or U2178 (N_2178,In_664,In_587);
nand U2179 (N_2179,In_655,In_958);
nand U2180 (N_2180,In_289,In_283);
nand U2181 (N_2181,In_251,In_683);
xor U2182 (N_2182,In_716,In_531);
nor U2183 (N_2183,In_996,In_676);
nand U2184 (N_2184,In_537,In_995);
nor U2185 (N_2185,In_994,In_457);
or U2186 (N_2186,In_754,In_810);
nand U2187 (N_2187,In_217,In_449);
xor U2188 (N_2188,In_214,In_607);
or U2189 (N_2189,In_87,In_319);
xnor U2190 (N_2190,In_2,In_387);
xor U2191 (N_2191,In_166,In_638);
and U2192 (N_2192,In_361,In_140);
or U2193 (N_2193,In_585,In_764);
nand U2194 (N_2194,In_140,In_237);
nor U2195 (N_2195,In_505,In_934);
or U2196 (N_2196,In_146,In_577);
and U2197 (N_2197,In_424,In_716);
and U2198 (N_2198,In_829,In_56);
or U2199 (N_2199,In_117,In_435);
nand U2200 (N_2200,In_589,In_201);
and U2201 (N_2201,In_812,In_832);
or U2202 (N_2202,In_859,In_554);
xor U2203 (N_2203,In_432,In_993);
nor U2204 (N_2204,In_165,In_793);
and U2205 (N_2205,In_784,In_144);
nand U2206 (N_2206,In_294,In_265);
nor U2207 (N_2207,In_500,In_423);
xor U2208 (N_2208,In_218,In_582);
nor U2209 (N_2209,In_353,In_898);
and U2210 (N_2210,In_437,In_96);
xor U2211 (N_2211,In_226,In_919);
and U2212 (N_2212,In_326,In_515);
and U2213 (N_2213,In_909,In_402);
and U2214 (N_2214,In_591,In_731);
nand U2215 (N_2215,In_403,In_478);
and U2216 (N_2216,In_371,In_46);
or U2217 (N_2217,In_470,In_579);
or U2218 (N_2218,In_823,In_93);
and U2219 (N_2219,In_862,In_584);
nor U2220 (N_2220,In_537,In_845);
and U2221 (N_2221,In_425,In_40);
xor U2222 (N_2222,In_3,In_61);
nand U2223 (N_2223,In_480,In_663);
and U2224 (N_2224,In_477,In_743);
and U2225 (N_2225,In_429,In_360);
or U2226 (N_2226,In_389,In_866);
or U2227 (N_2227,In_103,In_631);
nand U2228 (N_2228,In_485,In_419);
and U2229 (N_2229,In_42,In_564);
nand U2230 (N_2230,In_409,In_678);
nor U2231 (N_2231,In_579,In_81);
nand U2232 (N_2232,In_914,In_974);
nor U2233 (N_2233,In_133,In_403);
nand U2234 (N_2234,In_384,In_739);
and U2235 (N_2235,In_117,In_626);
nor U2236 (N_2236,In_179,In_350);
xor U2237 (N_2237,In_174,In_533);
xnor U2238 (N_2238,In_27,In_969);
nor U2239 (N_2239,In_390,In_731);
xor U2240 (N_2240,In_127,In_871);
xor U2241 (N_2241,In_140,In_983);
nand U2242 (N_2242,In_655,In_2);
and U2243 (N_2243,In_308,In_50);
xor U2244 (N_2244,In_225,In_324);
xor U2245 (N_2245,In_616,In_547);
nor U2246 (N_2246,In_342,In_82);
or U2247 (N_2247,In_932,In_290);
nor U2248 (N_2248,In_618,In_694);
xnor U2249 (N_2249,In_315,In_885);
nor U2250 (N_2250,In_513,In_31);
xnor U2251 (N_2251,In_871,In_61);
or U2252 (N_2252,In_719,In_445);
nor U2253 (N_2253,In_578,In_249);
xnor U2254 (N_2254,In_896,In_279);
and U2255 (N_2255,In_701,In_974);
nor U2256 (N_2256,In_614,In_104);
nand U2257 (N_2257,In_376,In_259);
or U2258 (N_2258,In_86,In_136);
nor U2259 (N_2259,In_789,In_138);
and U2260 (N_2260,In_280,In_469);
and U2261 (N_2261,In_650,In_555);
xnor U2262 (N_2262,In_622,In_570);
nor U2263 (N_2263,In_431,In_650);
nand U2264 (N_2264,In_544,In_603);
nand U2265 (N_2265,In_14,In_24);
or U2266 (N_2266,In_684,In_1);
and U2267 (N_2267,In_484,In_881);
or U2268 (N_2268,In_788,In_426);
or U2269 (N_2269,In_355,In_132);
and U2270 (N_2270,In_767,In_83);
xor U2271 (N_2271,In_774,In_462);
xor U2272 (N_2272,In_44,In_102);
nand U2273 (N_2273,In_107,In_696);
or U2274 (N_2274,In_773,In_367);
nor U2275 (N_2275,In_148,In_929);
nand U2276 (N_2276,In_779,In_431);
or U2277 (N_2277,In_561,In_659);
xnor U2278 (N_2278,In_987,In_844);
nand U2279 (N_2279,In_580,In_530);
or U2280 (N_2280,In_261,In_128);
and U2281 (N_2281,In_248,In_169);
or U2282 (N_2282,In_585,In_290);
nand U2283 (N_2283,In_852,In_896);
xor U2284 (N_2284,In_306,In_630);
xnor U2285 (N_2285,In_604,In_885);
nand U2286 (N_2286,In_895,In_61);
and U2287 (N_2287,In_303,In_251);
or U2288 (N_2288,In_261,In_669);
or U2289 (N_2289,In_984,In_964);
nand U2290 (N_2290,In_34,In_166);
or U2291 (N_2291,In_860,In_395);
nor U2292 (N_2292,In_556,In_634);
nand U2293 (N_2293,In_542,In_796);
xnor U2294 (N_2294,In_217,In_987);
and U2295 (N_2295,In_855,In_867);
or U2296 (N_2296,In_727,In_473);
or U2297 (N_2297,In_290,In_607);
nor U2298 (N_2298,In_836,In_395);
or U2299 (N_2299,In_719,In_576);
or U2300 (N_2300,In_700,In_338);
xnor U2301 (N_2301,In_307,In_661);
nor U2302 (N_2302,In_968,In_434);
or U2303 (N_2303,In_559,In_841);
nand U2304 (N_2304,In_62,In_588);
or U2305 (N_2305,In_844,In_547);
and U2306 (N_2306,In_417,In_156);
and U2307 (N_2307,In_472,In_408);
nand U2308 (N_2308,In_305,In_833);
nor U2309 (N_2309,In_567,In_672);
nor U2310 (N_2310,In_194,In_960);
nand U2311 (N_2311,In_158,In_823);
nand U2312 (N_2312,In_790,In_449);
xnor U2313 (N_2313,In_49,In_437);
or U2314 (N_2314,In_380,In_237);
nand U2315 (N_2315,In_7,In_260);
nand U2316 (N_2316,In_966,In_411);
xnor U2317 (N_2317,In_866,In_698);
nor U2318 (N_2318,In_730,In_519);
or U2319 (N_2319,In_736,In_400);
and U2320 (N_2320,In_467,In_593);
xnor U2321 (N_2321,In_142,In_968);
or U2322 (N_2322,In_570,In_827);
and U2323 (N_2323,In_728,In_485);
xnor U2324 (N_2324,In_519,In_130);
or U2325 (N_2325,In_278,In_715);
xnor U2326 (N_2326,In_28,In_779);
or U2327 (N_2327,In_300,In_330);
or U2328 (N_2328,In_300,In_926);
and U2329 (N_2329,In_20,In_684);
xnor U2330 (N_2330,In_459,In_825);
and U2331 (N_2331,In_850,In_878);
nor U2332 (N_2332,In_232,In_328);
nand U2333 (N_2333,In_780,In_65);
nor U2334 (N_2334,In_961,In_487);
and U2335 (N_2335,In_43,In_643);
nand U2336 (N_2336,In_459,In_159);
xor U2337 (N_2337,In_943,In_937);
or U2338 (N_2338,In_130,In_889);
xnor U2339 (N_2339,In_536,In_409);
nand U2340 (N_2340,In_496,In_216);
or U2341 (N_2341,In_192,In_844);
or U2342 (N_2342,In_42,In_392);
and U2343 (N_2343,In_787,In_379);
nor U2344 (N_2344,In_91,In_440);
or U2345 (N_2345,In_532,In_441);
nand U2346 (N_2346,In_449,In_310);
or U2347 (N_2347,In_343,In_96);
and U2348 (N_2348,In_784,In_911);
xnor U2349 (N_2349,In_893,In_647);
or U2350 (N_2350,In_163,In_412);
xnor U2351 (N_2351,In_742,In_470);
xnor U2352 (N_2352,In_195,In_508);
nand U2353 (N_2353,In_41,In_548);
nand U2354 (N_2354,In_677,In_987);
or U2355 (N_2355,In_590,In_359);
or U2356 (N_2356,In_476,In_547);
nor U2357 (N_2357,In_162,In_83);
nor U2358 (N_2358,In_172,In_595);
nor U2359 (N_2359,In_815,In_254);
nand U2360 (N_2360,In_805,In_191);
xnor U2361 (N_2361,In_853,In_263);
or U2362 (N_2362,In_8,In_469);
xor U2363 (N_2363,In_692,In_377);
or U2364 (N_2364,In_833,In_900);
nor U2365 (N_2365,In_709,In_674);
or U2366 (N_2366,In_392,In_261);
or U2367 (N_2367,In_952,In_917);
xnor U2368 (N_2368,In_182,In_958);
xnor U2369 (N_2369,In_308,In_34);
nor U2370 (N_2370,In_108,In_403);
nor U2371 (N_2371,In_345,In_158);
xnor U2372 (N_2372,In_181,In_273);
or U2373 (N_2373,In_546,In_138);
nand U2374 (N_2374,In_742,In_594);
and U2375 (N_2375,In_320,In_525);
nor U2376 (N_2376,In_674,In_277);
or U2377 (N_2377,In_721,In_867);
nand U2378 (N_2378,In_653,In_99);
nand U2379 (N_2379,In_575,In_635);
xor U2380 (N_2380,In_240,In_509);
and U2381 (N_2381,In_111,In_174);
nor U2382 (N_2382,In_950,In_336);
nand U2383 (N_2383,In_464,In_396);
nor U2384 (N_2384,In_726,In_597);
nor U2385 (N_2385,In_246,In_388);
or U2386 (N_2386,In_480,In_717);
nand U2387 (N_2387,In_700,In_529);
and U2388 (N_2388,In_605,In_61);
nor U2389 (N_2389,In_638,In_230);
nor U2390 (N_2390,In_438,In_374);
xnor U2391 (N_2391,In_573,In_252);
nor U2392 (N_2392,In_657,In_87);
nor U2393 (N_2393,In_278,In_736);
xnor U2394 (N_2394,In_889,In_786);
nor U2395 (N_2395,In_395,In_405);
and U2396 (N_2396,In_518,In_686);
nor U2397 (N_2397,In_882,In_781);
nor U2398 (N_2398,In_780,In_983);
or U2399 (N_2399,In_916,In_395);
nor U2400 (N_2400,In_922,In_578);
and U2401 (N_2401,In_793,In_245);
nand U2402 (N_2402,In_935,In_415);
and U2403 (N_2403,In_976,In_692);
and U2404 (N_2404,In_451,In_713);
nand U2405 (N_2405,In_121,In_515);
nor U2406 (N_2406,In_214,In_341);
nor U2407 (N_2407,In_596,In_155);
nand U2408 (N_2408,In_88,In_760);
or U2409 (N_2409,In_481,In_902);
and U2410 (N_2410,In_578,In_474);
xnor U2411 (N_2411,In_23,In_407);
nor U2412 (N_2412,In_849,In_98);
xnor U2413 (N_2413,In_464,In_168);
or U2414 (N_2414,In_353,In_440);
and U2415 (N_2415,In_459,In_560);
nor U2416 (N_2416,In_377,In_125);
and U2417 (N_2417,In_604,In_37);
nand U2418 (N_2418,In_898,In_597);
and U2419 (N_2419,In_475,In_287);
nor U2420 (N_2420,In_472,In_428);
nor U2421 (N_2421,In_267,In_516);
and U2422 (N_2422,In_639,In_739);
xnor U2423 (N_2423,In_91,In_748);
or U2424 (N_2424,In_57,In_690);
nor U2425 (N_2425,In_933,In_628);
xor U2426 (N_2426,In_88,In_479);
xnor U2427 (N_2427,In_372,In_543);
nor U2428 (N_2428,In_208,In_616);
or U2429 (N_2429,In_935,In_725);
or U2430 (N_2430,In_532,In_454);
and U2431 (N_2431,In_20,In_984);
nand U2432 (N_2432,In_560,In_511);
or U2433 (N_2433,In_984,In_241);
or U2434 (N_2434,In_762,In_626);
or U2435 (N_2435,In_473,In_348);
and U2436 (N_2436,In_461,In_405);
or U2437 (N_2437,In_637,In_294);
xor U2438 (N_2438,In_953,In_166);
nand U2439 (N_2439,In_827,In_339);
or U2440 (N_2440,In_998,In_762);
nand U2441 (N_2441,In_953,In_105);
nand U2442 (N_2442,In_545,In_391);
and U2443 (N_2443,In_185,In_761);
nor U2444 (N_2444,In_718,In_910);
or U2445 (N_2445,In_132,In_20);
or U2446 (N_2446,In_39,In_575);
nand U2447 (N_2447,In_253,In_423);
or U2448 (N_2448,In_779,In_883);
xnor U2449 (N_2449,In_387,In_596);
nand U2450 (N_2450,In_99,In_973);
or U2451 (N_2451,In_352,In_363);
or U2452 (N_2452,In_100,In_725);
xor U2453 (N_2453,In_570,In_412);
and U2454 (N_2454,In_338,In_895);
nor U2455 (N_2455,In_668,In_124);
or U2456 (N_2456,In_737,In_47);
and U2457 (N_2457,In_0,In_126);
nand U2458 (N_2458,In_184,In_875);
nand U2459 (N_2459,In_989,In_817);
nand U2460 (N_2460,In_926,In_455);
nor U2461 (N_2461,In_379,In_611);
nand U2462 (N_2462,In_835,In_259);
nand U2463 (N_2463,In_731,In_304);
xnor U2464 (N_2464,In_289,In_968);
and U2465 (N_2465,In_410,In_955);
or U2466 (N_2466,In_785,In_864);
nor U2467 (N_2467,In_793,In_861);
xor U2468 (N_2468,In_77,In_390);
nand U2469 (N_2469,In_78,In_117);
or U2470 (N_2470,In_658,In_721);
and U2471 (N_2471,In_711,In_221);
and U2472 (N_2472,In_112,In_497);
nor U2473 (N_2473,In_949,In_302);
and U2474 (N_2474,In_984,In_762);
nor U2475 (N_2475,In_4,In_860);
xnor U2476 (N_2476,In_803,In_890);
nor U2477 (N_2477,In_576,In_860);
and U2478 (N_2478,In_445,In_230);
xor U2479 (N_2479,In_370,In_395);
nor U2480 (N_2480,In_839,In_618);
nor U2481 (N_2481,In_513,In_188);
nor U2482 (N_2482,In_868,In_633);
or U2483 (N_2483,In_424,In_465);
or U2484 (N_2484,In_573,In_949);
nand U2485 (N_2485,In_330,In_143);
nand U2486 (N_2486,In_233,In_25);
xor U2487 (N_2487,In_626,In_675);
or U2488 (N_2488,In_145,In_902);
nor U2489 (N_2489,In_675,In_414);
and U2490 (N_2490,In_413,In_708);
and U2491 (N_2491,In_596,In_416);
nor U2492 (N_2492,In_180,In_453);
or U2493 (N_2493,In_617,In_128);
nor U2494 (N_2494,In_188,In_811);
or U2495 (N_2495,In_361,In_896);
xor U2496 (N_2496,In_492,In_976);
nor U2497 (N_2497,In_976,In_377);
xor U2498 (N_2498,In_948,In_731);
xnor U2499 (N_2499,In_627,In_379);
nor U2500 (N_2500,In_810,In_604);
nor U2501 (N_2501,In_122,In_191);
or U2502 (N_2502,In_60,In_681);
nor U2503 (N_2503,In_47,In_585);
and U2504 (N_2504,In_781,In_292);
nand U2505 (N_2505,In_646,In_493);
nor U2506 (N_2506,In_73,In_601);
nand U2507 (N_2507,In_971,In_169);
or U2508 (N_2508,In_260,In_448);
nor U2509 (N_2509,In_544,In_665);
nand U2510 (N_2510,In_990,In_88);
xnor U2511 (N_2511,In_959,In_135);
nand U2512 (N_2512,In_764,In_874);
nand U2513 (N_2513,In_911,In_523);
and U2514 (N_2514,In_157,In_603);
xnor U2515 (N_2515,In_941,In_741);
or U2516 (N_2516,In_243,In_766);
xnor U2517 (N_2517,In_562,In_365);
or U2518 (N_2518,In_753,In_626);
nand U2519 (N_2519,In_858,In_227);
xnor U2520 (N_2520,In_109,In_207);
and U2521 (N_2521,In_87,In_347);
xor U2522 (N_2522,In_818,In_515);
nor U2523 (N_2523,In_791,In_178);
and U2524 (N_2524,In_82,In_234);
and U2525 (N_2525,In_599,In_504);
or U2526 (N_2526,In_992,In_533);
or U2527 (N_2527,In_503,In_40);
nand U2528 (N_2528,In_484,In_483);
xnor U2529 (N_2529,In_827,In_51);
or U2530 (N_2530,In_572,In_482);
nand U2531 (N_2531,In_119,In_191);
nand U2532 (N_2532,In_487,In_36);
xnor U2533 (N_2533,In_371,In_820);
nand U2534 (N_2534,In_331,In_344);
or U2535 (N_2535,In_726,In_65);
or U2536 (N_2536,In_434,In_265);
xnor U2537 (N_2537,In_313,In_236);
nand U2538 (N_2538,In_1,In_228);
nor U2539 (N_2539,In_156,In_290);
xor U2540 (N_2540,In_452,In_138);
or U2541 (N_2541,In_35,In_692);
nor U2542 (N_2542,In_582,In_827);
and U2543 (N_2543,In_291,In_879);
nand U2544 (N_2544,In_148,In_892);
xor U2545 (N_2545,In_39,In_400);
and U2546 (N_2546,In_87,In_521);
and U2547 (N_2547,In_553,In_743);
nor U2548 (N_2548,In_801,In_345);
nand U2549 (N_2549,In_888,In_99);
nor U2550 (N_2550,In_595,In_295);
nor U2551 (N_2551,In_229,In_720);
nand U2552 (N_2552,In_497,In_886);
nand U2553 (N_2553,In_127,In_639);
xnor U2554 (N_2554,In_241,In_42);
or U2555 (N_2555,In_762,In_212);
and U2556 (N_2556,In_636,In_285);
nor U2557 (N_2557,In_420,In_818);
nand U2558 (N_2558,In_850,In_890);
xnor U2559 (N_2559,In_713,In_712);
or U2560 (N_2560,In_599,In_503);
xnor U2561 (N_2561,In_223,In_818);
and U2562 (N_2562,In_644,In_909);
or U2563 (N_2563,In_633,In_792);
xor U2564 (N_2564,In_840,In_126);
nor U2565 (N_2565,In_27,In_745);
nor U2566 (N_2566,In_906,In_222);
and U2567 (N_2567,In_167,In_757);
nor U2568 (N_2568,In_222,In_121);
nand U2569 (N_2569,In_321,In_573);
and U2570 (N_2570,In_251,In_390);
and U2571 (N_2571,In_463,In_495);
xor U2572 (N_2572,In_990,In_842);
xnor U2573 (N_2573,In_356,In_698);
xnor U2574 (N_2574,In_505,In_504);
nor U2575 (N_2575,In_112,In_830);
and U2576 (N_2576,In_630,In_341);
and U2577 (N_2577,In_533,In_449);
xnor U2578 (N_2578,In_439,In_157);
or U2579 (N_2579,In_289,In_445);
or U2580 (N_2580,In_206,In_937);
and U2581 (N_2581,In_17,In_603);
or U2582 (N_2582,In_406,In_378);
or U2583 (N_2583,In_733,In_861);
and U2584 (N_2584,In_200,In_220);
nand U2585 (N_2585,In_960,In_918);
and U2586 (N_2586,In_674,In_474);
nand U2587 (N_2587,In_647,In_747);
or U2588 (N_2588,In_122,In_544);
nand U2589 (N_2589,In_800,In_344);
xnor U2590 (N_2590,In_408,In_934);
and U2591 (N_2591,In_699,In_945);
nand U2592 (N_2592,In_378,In_185);
or U2593 (N_2593,In_623,In_702);
nor U2594 (N_2594,In_712,In_2);
nor U2595 (N_2595,In_165,In_473);
and U2596 (N_2596,In_166,In_747);
nor U2597 (N_2597,In_391,In_905);
nor U2598 (N_2598,In_39,In_366);
xnor U2599 (N_2599,In_821,In_601);
and U2600 (N_2600,In_891,In_194);
nand U2601 (N_2601,In_61,In_580);
or U2602 (N_2602,In_838,In_480);
or U2603 (N_2603,In_883,In_385);
or U2604 (N_2604,In_776,In_908);
or U2605 (N_2605,In_329,In_944);
nand U2606 (N_2606,In_438,In_571);
and U2607 (N_2607,In_661,In_820);
and U2608 (N_2608,In_401,In_425);
xnor U2609 (N_2609,In_600,In_29);
or U2610 (N_2610,In_295,In_701);
and U2611 (N_2611,In_300,In_570);
and U2612 (N_2612,In_895,In_925);
xnor U2613 (N_2613,In_53,In_516);
nor U2614 (N_2614,In_851,In_502);
or U2615 (N_2615,In_309,In_153);
and U2616 (N_2616,In_286,In_385);
xor U2617 (N_2617,In_412,In_449);
nor U2618 (N_2618,In_351,In_501);
nand U2619 (N_2619,In_978,In_241);
or U2620 (N_2620,In_493,In_89);
xnor U2621 (N_2621,In_724,In_237);
nor U2622 (N_2622,In_101,In_998);
nor U2623 (N_2623,In_638,In_765);
nor U2624 (N_2624,In_863,In_380);
nand U2625 (N_2625,In_39,In_173);
nor U2626 (N_2626,In_255,In_734);
nand U2627 (N_2627,In_488,In_259);
xor U2628 (N_2628,In_497,In_417);
xor U2629 (N_2629,In_8,In_902);
and U2630 (N_2630,In_477,In_90);
or U2631 (N_2631,In_898,In_348);
nor U2632 (N_2632,In_44,In_472);
nand U2633 (N_2633,In_44,In_441);
and U2634 (N_2634,In_30,In_607);
or U2635 (N_2635,In_567,In_645);
nor U2636 (N_2636,In_419,In_409);
nor U2637 (N_2637,In_528,In_22);
nand U2638 (N_2638,In_614,In_190);
nand U2639 (N_2639,In_942,In_900);
nand U2640 (N_2640,In_503,In_65);
or U2641 (N_2641,In_607,In_464);
and U2642 (N_2642,In_84,In_497);
xnor U2643 (N_2643,In_449,In_538);
nor U2644 (N_2644,In_974,In_40);
and U2645 (N_2645,In_553,In_550);
nor U2646 (N_2646,In_580,In_771);
xnor U2647 (N_2647,In_287,In_561);
nand U2648 (N_2648,In_920,In_668);
or U2649 (N_2649,In_267,In_310);
and U2650 (N_2650,In_896,In_951);
nand U2651 (N_2651,In_821,In_332);
nand U2652 (N_2652,In_221,In_276);
and U2653 (N_2653,In_337,In_342);
xnor U2654 (N_2654,In_804,In_902);
xor U2655 (N_2655,In_10,In_874);
xnor U2656 (N_2656,In_386,In_339);
and U2657 (N_2657,In_38,In_314);
or U2658 (N_2658,In_200,In_319);
nand U2659 (N_2659,In_147,In_155);
and U2660 (N_2660,In_291,In_54);
nor U2661 (N_2661,In_947,In_92);
nor U2662 (N_2662,In_612,In_532);
nor U2663 (N_2663,In_791,In_407);
and U2664 (N_2664,In_101,In_129);
xor U2665 (N_2665,In_15,In_300);
or U2666 (N_2666,In_834,In_879);
nor U2667 (N_2667,In_852,In_832);
nand U2668 (N_2668,In_753,In_793);
and U2669 (N_2669,In_822,In_623);
and U2670 (N_2670,In_342,In_671);
nand U2671 (N_2671,In_778,In_248);
xor U2672 (N_2672,In_664,In_380);
nor U2673 (N_2673,In_663,In_803);
nand U2674 (N_2674,In_117,In_590);
or U2675 (N_2675,In_219,In_188);
and U2676 (N_2676,In_795,In_813);
nand U2677 (N_2677,In_79,In_684);
nor U2678 (N_2678,In_97,In_933);
or U2679 (N_2679,In_816,In_331);
xnor U2680 (N_2680,In_771,In_737);
nor U2681 (N_2681,In_200,In_467);
or U2682 (N_2682,In_762,In_508);
nand U2683 (N_2683,In_867,In_18);
nor U2684 (N_2684,In_50,In_381);
nor U2685 (N_2685,In_506,In_458);
nand U2686 (N_2686,In_435,In_770);
xnor U2687 (N_2687,In_959,In_923);
xor U2688 (N_2688,In_132,In_142);
nor U2689 (N_2689,In_684,In_458);
and U2690 (N_2690,In_129,In_173);
nor U2691 (N_2691,In_93,In_584);
nand U2692 (N_2692,In_514,In_830);
xnor U2693 (N_2693,In_291,In_711);
or U2694 (N_2694,In_542,In_534);
or U2695 (N_2695,In_715,In_475);
xor U2696 (N_2696,In_542,In_592);
nand U2697 (N_2697,In_929,In_987);
and U2698 (N_2698,In_618,In_296);
nor U2699 (N_2699,In_848,In_957);
nor U2700 (N_2700,In_685,In_417);
nor U2701 (N_2701,In_603,In_263);
xnor U2702 (N_2702,In_888,In_379);
nor U2703 (N_2703,In_562,In_781);
or U2704 (N_2704,In_335,In_848);
nand U2705 (N_2705,In_7,In_299);
and U2706 (N_2706,In_527,In_159);
xnor U2707 (N_2707,In_170,In_150);
and U2708 (N_2708,In_628,In_352);
or U2709 (N_2709,In_268,In_120);
or U2710 (N_2710,In_794,In_754);
or U2711 (N_2711,In_281,In_17);
and U2712 (N_2712,In_263,In_475);
nand U2713 (N_2713,In_924,In_231);
or U2714 (N_2714,In_6,In_961);
xnor U2715 (N_2715,In_534,In_811);
and U2716 (N_2716,In_723,In_597);
and U2717 (N_2717,In_439,In_435);
nand U2718 (N_2718,In_351,In_601);
nand U2719 (N_2719,In_741,In_736);
or U2720 (N_2720,In_413,In_373);
xor U2721 (N_2721,In_412,In_21);
or U2722 (N_2722,In_427,In_508);
nor U2723 (N_2723,In_170,In_729);
nor U2724 (N_2724,In_936,In_802);
nand U2725 (N_2725,In_769,In_613);
or U2726 (N_2726,In_720,In_900);
nor U2727 (N_2727,In_928,In_200);
or U2728 (N_2728,In_509,In_641);
nor U2729 (N_2729,In_875,In_143);
nand U2730 (N_2730,In_666,In_384);
xnor U2731 (N_2731,In_663,In_857);
nand U2732 (N_2732,In_208,In_934);
or U2733 (N_2733,In_15,In_320);
or U2734 (N_2734,In_511,In_752);
and U2735 (N_2735,In_780,In_393);
or U2736 (N_2736,In_519,In_702);
xnor U2737 (N_2737,In_933,In_965);
nand U2738 (N_2738,In_278,In_834);
xnor U2739 (N_2739,In_442,In_34);
nand U2740 (N_2740,In_301,In_358);
or U2741 (N_2741,In_797,In_822);
or U2742 (N_2742,In_711,In_157);
and U2743 (N_2743,In_30,In_23);
nand U2744 (N_2744,In_312,In_147);
nor U2745 (N_2745,In_846,In_616);
xnor U2746 (N_2746,In_586,In_572);
xor U2747 (N_2747,In_691,In_96);
nand U2748 (N_2748,In_915,In_44);
or U2749 (N_2749,In_118,In_527);
nor U2750 (N_2750,In_17,In_200);
xnor U2751 (N_2751,In_874,In_978);
xnor U2752 (N_2752,In_247,In_300);
nand U2753 (N_2753,In_376,In_874);
nor U2754 (N_2754,In_298,In_767);
xor U2755 (N_2755,In_807,In_771);
and U2756 (N_2756,In_341,In_569);
or U2757 (N_2757,In_995,In_957);
nand U2758 (N_2758,In_997,In_92);
xor U2759 (N_2759,In_66,In_470);
xor U2760 (N_2760,In_7,In_745);
and U2761 (N_2761,In_382,In_126);
nor U2762 (N_2762,In_821,In_65);
nor U2763 (N_2763,In_998,In_298);
or U2764 (N_2764,In_26,In_350);
nand U2765 (N_2765,In_948,In_836);
nand U2766 (N_2766,In_379,In_374);
nor U2767 (N_2767,In_815,In_275);
nor U2768 (N_2768,In_558,In_731);
nand U2769 (N_2769,In_367,In_198);
nor U2770 (N_2770,In_202,In_29);
and U2771 (N_2771,In_311,In_552);
nand U2772 (N_2772,In_585,In_576);
xor U2773 (N_2773,In_373,In_851);
xnor U2774 (N_2774,In_307,In_715);
and U2775 (N_2775,In_128,In_29);
nand U2776 (N_2776,In_97,In_682);
and U2777 (N_2777,In_753,In_534);
xor U2778 (N_2778,In_433,In_179);
nand U2779 (N_2779,In_889,In_913);
or U2780 (N_2780,In_695,In_158);
nor U2781 (N_2781,In_257,In_229);
nand U2782 (N_2782,In_935,In_950);
or U2783 (N_2783,In_804,In_717);
nor U2784 (N_2784,In_688,In_567);
nor U2785 (N_2785,In_326,In_685);
nand U2786 (N_2786,In_274,In_131);
or U2787 (N_2787,In_927,In_849);
or U2788 (N_2788,In_693,In_661);
and U2789 (N_2789,In_955,In_383);
nand U2790 (N_2790,In_411,In_715);
nand U2791 (N_2791,In_193,In_604);
xor U2792 (N_2792,In_637,In_115);
nand U2793 (N_2793,In_980,In_283);
and U2794 (N_2794,In_80,In_325);
xor U2795 (N_2795,In_470,In_813);
xor U2796 (N_2796,In_912,In_691);
nor U2797 (N_2797,In_530,In_157);
xor U2798 (N_2798,In_724,In_696);
and U2799 (N_2799,In_240,In_78);
or U2800 (N_2800,In_469,In_138);
and U2801 (N_2801,In_334,In_932);
and U2802 (N_2802,In_154,In_695);
and U2803 (N_2803,In_472,In_777);
nor U2804 (N_2804,In_386,In_791);
or U2805 (N_2805,In_904,In_66);
nand U2806 (N_2806,In_952,In_453);
xnor U2807 (N_2807,In_217,In_423);
xnor U2808 (N_2808,In_11,In_203);
xnor U2809 (N_2809,In_764,In_978);
or U2810 (N_2810,In_584,In_933);
nor U2811 (N_2811,In_681,In_716);
nor U2812 (N_2812,In_661,In_386);
nand U2813 (N_2813,In_719,In_130);
nand U2814 (N_2814,In_981,In_259);
nor U2815 (N_2815,In_86,In_357);
or U2816 (N_2816,In_569,In_720);
or U2817 (N_2817,In_951,In_199);
and U2818 (N_2818,In_137,In_637);
nor U2819 (N_2819,In_401,In_441);
or U2820 (N_2820,In_494,In_763);
nand U2821 (N_2821,In_213,In_155);
and U2822 (N_2822,In_449,In_653);
nand U2823 (N_2823,In_27,In_540);
and U2824 (N_2824,In_660,In_705);
or U2825 (N_2825,In_878,In_644);
nor U2826 (N_2826,In_716,In_939);
xnor U2827 (N_2827,In_254,In_668);
nand U2828 (N_2828,In_779,In_889);
or U2829 (N_2829,In_951,In_686);
xor U2830 (N_2830,In_123,In_926);
xor U2831 (N_2831,In_763,In_843);
nor U2832 (N_2832,In_674,In_404);
and U2833 (N_2833,In_609,In_845);
or U2834 (N_2834,In_982,In_128);
nand U2835 (N_2835,In_475,In_318);
or U2836 (N_2836,In_784,In_760);
and U2837 (N_2837,In_853,In_886);
or U2838 (N_2838,In_992,In_622);
and U2839 (N_2839,In_446,In_990);
nor U2840 (N_2840,In_472,In_31);
nand U2841 (N_2841,In_737,In_595);
or U2842 (N_2842,In_333,In_336);
xnor U2843 (N_2843,In_268,In_795);
nand U2844 (N_2844,In_817,In_553);
and U2845 (N_2845,In_766,In_333);
or U2846 (N_2846,In_115,In_446);
or U2847 (N_2847,In_257,In_592);
nor U2848 (N_2848,In_82,In_296);
or U2849 (N_2849,In_332,In_760);
nor U2850 (N_2850,In_233,In_279);
xnor U2851 (N_2851,In_355,In_104);
and U2852 (N_2852,In_596,In_390);
nand U2853 (N_2853,In_31,In_224);
xnor U2854 (N_2854,In_827,In_378);
and U2855 (N_2855,In_780,In_652);
xnor U2856 (N_2856,In_667,In_778);
or U2857 (N_2857,In_572,In_29);
and U2858 (N_2858,In_194,In_618);
xor U2859 (N_2859,In_561,In_408);
and U2860 (N_2860,In_797,In_621);
xor U2861 (N_2861,In_537,In_953);
nand U2862 (N_2862,In_100,In_754);
and U2863 (N_2863,In_592,In_210);
nor U2864 (N_2864,In_78,In_818);
nand U2865 (N_2865,In_533,In_740);
or U2866 (N_2866,In_31,In_417);
or U2867 (N_2867,In_303,In_853);
xor U2868 (N_2868,In_873,In_342);
xor U2869 (N_2869,In_23,In_980);
or U2870 (N_2870,In_515,In_341);
xnor U2871 (N_2871,In_636,In_64);
and U2872 (N_2872,In_818,In_970);
nand U2873 (N_2873,In_884,In_266);
and U2874 (N_2874,In_677,In_79);
xor U2875 (N_2875,In_381,In_80);
nand U2876 (N_2876,In_700,In_519);
xor U2877 (N_2877,In_20,In_229);
or U2878 (N_2878,In_253,In_731);
or U2879 (N_2879,In_732,In_938);
or U2880 (N_2880,In_724,In_374);
and U2881 (N_2881,In_13,In_619);
xor U2882 (N_2882,In_644,In_342);
and U2883 (N_2883,In_551,In_105);
nand U2884 (N_2884,In_72,In_817);
nand U2885 (N_2885,In_266,In_862);
nor U2886 (N_2886,In_34,In_912);
nand U2887 (N_2887,In_942,In_317);
or U2888 (N_2888,In_849,In_533);
nand U2889 (N_2889,In_954,In_266);
or U2890 (N_2890,In_820,In_663);
and U2891 (N_2891,In_837,In_520);
xnor U2892 (N_2892,In_70,In_121);
nand U2893 (N_2893,In_418,In_386);
xnor U2894 (N_2894,In_85,In_163);
xor U2895 (N_2895,In_176,In_995);
or U2896 (N_2896,In_764,In_490);
or U2897 (N_2897,In_798,In_980);
xor U2898 (N_2898,In_958,In_508);
xor U2899 (N_2899,In_779,In_467);
or U2900 (N_2900,In_362,In_183);
xor U2901 (N_2901,In_127,In_184);
xor U2902 (N_2902,In_578,In_14);
or U2903 (N_2903,In_613,In_288);
or U2904 (N_2904,In_918,In_219);
or U2905 (N_2905,In_492,In_520);
xnor U2906 (N_2906,In_264,In_756);
nand U2907 (N_2907,In_745,In_806);
xor U2908 (N_2908,In_604,In_84);
and U2909 (N_2909,In_161,In_50);
nand U2910 (N_2910,In_644,In_276);
nand U2911 (N_2911,In_967,In_66);
xnor U2912 (N_2912,In_189,In_474);
nor U2913 (N_2913,In_940,In_936);
nor U2914 (N_2914,In_315,In_189);
or U2915 (N_2915,In_911,In_794);
nand U2916 (N_2916,In_118,In_191);
and U2917 (N_2917,In_152,In_837);
xnor U2918 (N_2918,In_245,In_876);
or U2919 (N_2919,In_3,In_381);
or U2920 (N_2920,In_514,In_129);
nor U2921 (N_2921,In_38,In_713);
nor U2922 (N_2922,In_656,In_398);
xor U2923 (N_2923,In_736,In_839);
nor U2924 (N_2924,In_254,In_66);
and U2925 (N_2925,In_390,In_302);
or U2926 (N_2926,In_806,In_344);
and U2927 (N_2927,In_957,In_158);
and U2928 (N_2928,In_713,In_809);
or U2929 (N_2929,In_586,In_881);
or U2930 (N_2930,In_6,In_919);
nor U2931 (N_2931,In_880,In_98);
nand U2932 (N_2932,In_982,In_748);
and U2933 (N_2933,In_374,In_371);
nor U2934 (N_2934,In_867,In_436);
xor U2935 (N_2935,In_795,In_866);
xor U2936 (N_2936,In_329,In_115);
nand U2937 (N_2937,In_339,In_21);
nor U2938 (N_2938,In_244,In_171);
or U2939 (N_2939,In_813,In_134);
and U2940 (N_2940,In_45,In_511);
nor U2941 (N_2941,In_728,In_954);
or U2942 (N_2942,In_126,In_730);
or U2943 (N_2943,In_666,In_130);
nor U2944 (N_2944,In_536,In_849);
nand U2945 (N_2945,In_876,In_502);
nor U2946 (N_2946,In_617,In_130);
nand U2947 (N_2947,In_843,In_811);
or U2948 (N_2948,In_795,In_88);
nor U2949 (N_2949,In_881,In_724);
nor U2950 (N_2950,In_467,In_452);
nor U2951 (N_2951,In_489,In_236);
or U2952 (N_2952,In_409,In_382);
and U2953 (N_2953,In_393,In_351);
and U2954 (N_2954,In_689,In_417);
nand U2955 (N_2955,In_327,In_790);
and U2956 (N_2956,In_573,In_831);
or U2957 (N_2957,In_808,In_674);
xor U2958 (N_2958,In_311,In_184);
and U2959 (N_2959,In_460,In_266);
or U2960 (N_2960,In_446,In_553);
and U2961 (N_2961,In_807,In_490);
xor U2962 (N_2962,In_682,In_59);
nand U2963 (N_2963,In_398,In_923);
nor U2964 (N_2964,In_475,In_444);
or U2965 (N_2965,In_759,In_418);
nor U2966 (N_2966,In_245,In_724);
nand U2967 (N_2967,In_434,In_139);
nor U2968 (N_2968,In_273,In_842);
and U2969 (N_2969,In_938,In_131);
nand U2970 (N_2970,In_564,In_195);
or U2971 (N_2971,In_891,In_760);
nand U2972 (N_2972,In_333,In_943);
nand U2973 (N_2973,In_833,In_65);
nand U2974 (N_2974,In_198,In_547);
or U2975 (N_2975,In_121,In_772);
nand U2976 (N_2976,In_128,In_137);
or U2977 (N_2977,In_387,In_466);
xnor U2978 (N_2978,In_889,In_288);
nor U2979 (N_2979,In_501,In_133);
nand U2980 (N_2980,In_996,In_593);
nor U2981 (N_2981,In_93,In_486);
nor U2982 (N_2982,In_458,In_603);
nand U2983 (N_2983,In_697,In_363);
xor U2984 (N_2984,In_967,In_174);
xnor U2985 (N_2985,In_592,In_305);
xor U2986 (N_2986,In_974,In_150);
or U2987 (N_2987,In_123,In_199);
xnor U2988 (N_2988,In_470,In_558);
xnor U2989 (N_2989,In_38,In_678);
nor U2990 (N_2990,In_116,In_50);
nor U2991 (N_2991,In_443,In_766);
nor U2992 (N_2992,In_328,In_29);
nand U2993 (N_2993,In_430,In_603);
nor U2994 (N_2994,In_929,In_872);
xnor U2995 (N_2995,In_110,In_476);
or U2996 (N_2996,In_437,In_919);
nor U2997 (N_2997,In_732,In_569);
xnor U2998 (N_2998,In_575,In_679);
and U2999 (N_2999,In_235,In_414);
and U3000 (N_3000,In_782,In_963);
and U3001 (N_3001,In_811,In_476);
nor U3002 (N_3002,In_95,In_900);
nand U3003 (N_3003,In_898,In_140);
xnor U3004 (N_3004,In_100,In_504);
and U3005 (N_3005,In_376,In_843);
or U3006 (N_3006,In_607,In_890);
and U3007 (N_3007,In_87,In_566);
nand U3008 (N_3008,In_693,In_776);
xor U3009 (N_3009,In_63,In_552);
xor U3010 (N_3010,In_480,In_601);
or U3011 (N_3011,In_802,In_178);
or U3012 (N_3012,In_5,In_664);
nand U3013 (N_3013,In_699,In_838);
or U3014 (N_3014,In_533,In_293);
nor U3015 (N_3015,In_675,In_253);
and U3016 (N_3016,In_988,In_60);
xnor U3017 (N_3017,In_534,In_920);
and U3018 (N_3018,In_213,In_270);
nand U3019 (N_3019,In_630,In_195);
xor U3020 (N_3020,In_807,In_283);
xnor U3021 (N_3021,In_457,In_20);
nand U3022 (N_3022,In_488,In_990);
or U3023 (N_3023,In_286,In_920);
nor U3024 (N_3024,In_68,In_61);
nand U3025 (N_3025,In_864,In_168);
nor U3026 (N_3026,In_638,In_837);
or U3027 (N_3027,In_548,In_80);
and U3028 (N_3028,In_675,In_778);
nand U3029 (N_3029,In_849,In_609);
and U3030 (N_3030,In_847,In_945);
xnor U3031 (N_3031,In_567,In_207);
or U3032 (N_3032,In_22,In_95);
or U3033 (N_3033,In_378,In_850);
and U3034 (N_3034,In_413,In_991);
nor U3035 (N_3035,In_829,In_340);
nand U3036 (N_3036,In_7,In_931);
nand U3037 (N_3037,In_256,In_512);
nor U3038 (N_3038,In_77,In_593);
or U3039 (N_3039,In_454,In_79);
xnor U3040 (N_3040,In_945,In_471);
xnor U3041 (N_3041,In_579,In_900);
nor U3042 (N_3042,In_333,In_548);
xor U3043 (N_3043,In_995,In_0);
nor U3044 (N_3044,In_470,In_722);
or U3045 (N_3045,In_63,In_296);
or U3046 (N_3046,In_71,In_688);
nor U3047 (N_3047,In_375,In_861);
or U3048 (N_3048,In_129,In_631);
nor U3049 (N_3049,In_642,In_579);
nand U3050 (N_3050,In_72,In_125);
or U3051 (N_3051,In_951,In_144);
nand U3052 (N_3052,In_266,In_635);
or U3053 (N_3053,In_675,In_203);
nand U3054 (N_3054,In_771,In_127);
xnor U3055 (N_3055,In_683,In_95);
or U3056 (N_3056,In_441,In_371);
and U3057 (N_3057,In_198,In_28);
xor U3058 (N_3058,In_175,In_234);
nor U3059 (N_3059,In_977,In_442);
nor U3060 (N_3060,In_15,In_951);
nand U3061 (N_3061,In_111,In_300);
nor U3062 (N_3062,In_290,In_465);
and U3063 (N_3063,In_482,In_900);
xnor U3064 (N_3064,In_271,In_255);
and U3065 (N_3065,In_654,In_290);
nor U3066 (N_3066,In_538,In_144);
xor U3067 (N_3067,In_835,In_289);
nand U3068 (N_3068,In_97,In_296);
or U3069 (N_3069,In_335,In_806);
nand U3070 (N_3070,In_399,In_668);
xor U3071 (N_3071,In_451,In_248);
and U3072 (N_3072,In_933,In_169);
nor U3073 (N_3073,In_911,In_167);
nand U3074 (N_3074,In_431,In_727);
or U3075 (N_3075,In_709,In_929);
xnor U3076 (N_3076,In_404,In_767);
and U3077 (N_3077,In_641,In_464);
or U3078 (N_3078,In_209,In_166);
and U3079 (N_3079,In_893,In_126);
and U3080 (N_3080,In_84,In_304);
nand U3081 (N_3081,In_701,In_356);
xnor U3082 (N_3082,In_825,In_963);
xor U3083 (N_3083,In_765,In_279);
nor U3084 (N_3084,In_403,In_769);
xor U3085 (N_3085,In_342,In_498);
nor U3086 (N_3086,In_391,In_86);
or U3087 (N_3087,In_688,In_616);
xor U3088 (N_3088,In_803,In_182);
xor U3089 (N_3089,In_787,In_99);
nand U3090 (N_3090,In_87,In_563);
nor U3091 (N_3091,In_248,In_929);
xnor U3092 (N_3092,In_708,In_798);
and U3093 (N_3093,In_431,In_695);
or U3094 (N_3094,In_134,In_19);
or U3095 (N_3095,In_733,In_278);
nand U3096 (N_3096,In_210,In_203);
nor U3097 (N_3097,In_991,In_882);
nand U3098 (N_3098,In_115,In_287);
xnor U3099 (N_3099,In_398,In_62);
xnor U3100 (N_3100,In_191,In_393);
and U3101 (N_3101,In_147,In_339);
or U3102 (N_3102,In_102,In_994);
nor U3103 (N_3103,In_364,In_15);
or U3104 (N_3104,In_418,In_629);
nor U3105 (N_3105,In_394,In_293);
nand U3106 (N_3106,In_845,In_825);
nand U3107 (N_3107,In_137,In_956);
nor U3108 (N_3108,In_544,In_820);
nand U3109 (N_3109,In_951,In_546);
or U3110 (N_3110,In_144,In_529);
nand U3111 (N_3111,In_651,In_54);
xor U3112 (N_3112,In_991,In_836);
and U3113 (N_3113,In_30,In_762);
or U3114 (N_3114,In_977,In_105);
nand U3115 (N_3115,In_495,In_568);
and U3116 (N_3116,In_236,In_668);
xnor U3117 (N_3117,In_246,In_522);
xnor U3118 (N_3118,In_329,In_641);
nor U3119 (N_3119,In_460,In_514);
or U3120 (N_3120,In_880,In_320);
nand U3121 (N_3121,In_74,In_878);
nand U3122 (N_3122,In_271,In_908);
nor U3123 (N_3123,In_566,In_669);
or U3124 (N_3124,In_831,In_455);
or U3125 (N_3125,In_810,In_314);
nand U3126 (N_3126,In_61,In_130);
nand U3127 (N_3127,In_43,In_28);
nand U3128 (N_3128,In_525,In_645);
or U3129 (N_3129,In_908,In_334);
and U3130 (N_3130,In_105,In_192);
or U3131 (N_3131,In_737,In_677);
xnor U3132 (N_3132,In_978,In_399);
and U3133 (N_3133,In_708,In_968);
nand U3134 (N_3134,In_901,In_395);
nor U3135 (N_3135,In_787,In_955);
xor U3136 (N_3136,In_864,In_687);
xor U3137 (N_3137,In_787,In_746);
or U3138 (N_3138,In_454,In_383);
nor U3139 (N_3139,In_219,In_64);
and U3140 (N_3140,In_697,In_237);
nor U3141 (N_3141,In_169,In_947);
xnor U3142 (N_3142,In_943,In_658);
nand U3143 (N_3143,In_894,In_859);
and U3144 (N_3144,In_290,In_995);
nand U3145 (N_3145,In_517,In_629);
and U3146 (N_3146,In_22,In_113);
or U3147 (N_3147,In_526,In_115);
xnor U3148 (N_3148,In_778,In_758);
nor U3149 (N_3149,In_959,In_74);
nor U3150 (N_3150,In_843,In_494);
xor U3151 (N_3151,In_420,In_849);
nor U3152 (N_3152,In_403,In_615);
and U3153 (N_3153,In_213,In_120);
xor U3154 (N_3154,In_893,In_988);
and U3155 (N_3155,In_905,In_509);
and U3156 (N_3156,In_272,In_319);
xnor U3157 (N_3157,In_77,In_556);
nor U3158 (N_3158,In_905,In_883);
xor U3159 (N_3159,In_160,In_283);
and U3160 (N_3160,In_191,In_454);
xor U3161 (N_3161,In_725,In_663);
or U3162 (N_3162,In_534,In_836);
and U3163 (N_3163,In_619,In_63);
nor U3164 (N_3164,In_445,In_879);
and U3165 (N_3165,In_640,In_84);
nand U3166 (N_3166,In_551,In_797);
xor U3167 (N_3167,In_627,In_301);
or U3168 (N_3168,In_424,In_993);
nand U3169 (N_3169,In_209,In_755);
nand U3170 (N_3170,In_916,In_132);
nor U3171 (N_3171,In_920,In_902);
xor U3172 (N_3172,In_800,In_244);
and U3173 (N_3173,In_181,In_778);
or U3174 (N_3174,In_876,In_203);
nor U3175 (N_3175,In_66,In_241);
nand U3176 (N_3176,In_657,In_265);
xnor U3177 (N_3177,In_492,In_451);
nand U3178 (N_3178,In_753,In_740);
or U3179 (N_3179,In_645,In_775);
nor U3180 (N_3180,In_309,In_569);
and U3181 (N_3181,In_636,In_610);
nor U3182 (N_3182,In_632,In_422);
and U3183 (N_3183,In_597,In_834);
nand U3184 (N_3184,In_128,In_840);
nor U3185 (N_3185,In_180,In_998);
xnor U3186 (N_3186,In_506,In_972);
nand U3187 (N_3187,In_338,In_194);
or U3188 (N_3188,In_10,In_228);
nand U3189 (N_3189,In_496,In_93);
and U3190 (N_3190,In_970,In_747);
and U3191 (N_3191,In_212,In_927);
and U3192 (N_3192,In_297,In_774);
nand U3193 (N_3193,In_873,In_511);
or U3194 (N_3194,In_290,In_144);
nor U3195 (N_3195,In_384,In_95);
and U3196 (N_3196,In_486,In_834);
or U3197 (N_3197,In_149,In_861);
nor U3198 (N_3198,In_792,In_508);
nand U3199 (N_3199,In_115,In_335);
nor U3200 (N_3200,In_85,In_909);
or U3201 (N_3201,In_297,In_243);
nand U3202 (N_3202,In_546,In_17);
xor U3203 (N_3203,In_555,In_695);
and U3204 (N_3204,In_407,In_402);
and U3205 (N_3205,In_289,In_141);
and U3206 (N_3206,In_317,In_447);
nor U3207 (N_3207,In_959,In_180);
or U3208 (N_3208,In_367,In_878);
xnor U3209 (N_3209,In_689,In_266);
or U3210 (N_3210,In_835,In_873);
nand U3211 (N_3211,In_995,In_29);
or U3212 (N_3212,In_881,In_124);
or U3213 (N_3213,In_238,In_157);
or U3214 (N_3214,In_173,In_56);
or U3215 (N_3215,In_529,In_459);
nand U3216 (N_3216,In_828,In_679);
and U3217 (N_3217,In_193,In_923);
and U3218 (N_3218,In_401,In_649);
or U3219 (N_3219,In_59,In_124);
nor U3220 (N_3220,In_620,In_571);
nand U3221 (N_3221,In_828,In_630);
or U3222 (N_3222,In_803,In_382);
and U3223 (N_3223,In_439,In_300);
xnor U3224 (N_3224,In_707,In_833);
nor U3225 (N_3225,In_392,In_205);
nand U3226 (N_3226,In_165,In_210);
or U3227 (N_3227,In_314,In_129);
or U3228 (N_3228,In_998,In_727);
xor U3229 (N_3229,In_779,In_527);
or U3230 (N_3230,In_947,In_562);
nand U3231 (N_3231,In_840,In_931);
or U3232 (N_3232,In_238,In_392);
nor U3233 (N_3233,In_407,In_89);
nor U3234 (N_3234,In_244,In_396);
and U3235 (N_3235,In_859,In_488);
or U3236 (N_3236,In_383,In_797);
nand U3237 (N_3237,In_420,In_805);
nand U3238 (N_3238,In_471,In_824);
xnor U3239 (N_3239,In_631,In_536);
nor U3240 (N_3240,In_87,In_581);
xor U3241 (N_3241,In_635,In_179);
nand U3242 (N_3242,In_219,In_927);
and U3243 (N_3243,In_184,In_468);
nand U3244 (N_3244,In_920,In_566);
nor U3245 (N_3245,In_277,In_125);
or U3246 (N_3246,In_740,In_63);
and U3247 (N_3247,In_112,In_171);
nand U3248 (N_3248,In_323,In_441);
and U3249 (N_3249,In_209,In_386);
nor U3250 (N_3250,In_182,In_551);
or U3251 (N_3251,In_864,In_626);
xnor U3252 (N_3252,In_252,In_273);
nand U3253 (N_3253,In_935,In_714);
nor U3254 (N_3254,In_112,In_141);
and U3255 (N_3255,In_744,In_63);
nor U3256 (N_3256,In_106,In_546);
and U3257 (N_3257,In_711,In_701);
nand U3258 (N_3258,In_811,In_157);
nor U3259 (N_3259,In_857,In_266);
nor U3260 (N_3260,In_720,In_112);
and U3261 (N_3261,In_504,In_924);
and U3262 (N_3262,In_393,In_684);
and U3263 (N_3263,In_140,In_519);
nand U3264 (N_3264,In_328,In_92);
nor U3265 (N_3265,In_926,In_226);
xor U3266 (N_3266,In_154,In_250);
and U3267 (N_3267,In_44,In_450);
xor U3268 (N_3268,In_209,In_897);
and U3269 (N_3269,In_869,In_509);
or U3270 (N_3270,In_449,In_336);
nor U3271 (N_3271,In_542,In_175);
nand U3272 (N_3272,In_791,In_398);
nand U3273 (N_3273,In_892,In_406);
and U3274 (N_3274,In_710,In_445);
xor U3275 (N_3275,In_355,In_299);
nor U3276 (N_3276,In_751,In_832);
and U3277 (N_3277,In_488,In_179);
or U3278 (N_3278,In_241,In_575);
nor U3279 (N_3279,In_112,In_236);
and U3280 (N_3280,In_573,In_484);
or U3281 (N_3281,In_554,In_963);
xor U3282 (N_3282,In_609,In_655);
and U3283 (N_3283,In_722,In_762);
nor U3284 (N_3284,In_227,In_847);
and U3285 (N_3285,In_794,In_61);
nand U3286 (N_3286,In_28,In_771);
nor U3287 (N_3287,In_97,In_832);
xor U3288 (N_3288,In_943,In_556);
or U3289 (N_3289,In_653,In_500);
nor U3290 (N_3290,In_757,In_986);
nor U3291 (N_3291,In_633,In_641);
nor U3292 (N_3292,In_380,In_874);
nand U3293 (N_3293,In_755,In_165);
xnor U3294 (N_3294,In_224,In_439);
and U3295 (N_3295,In_406,In_647);
nand U3296 (N_3296,In_139,In_817);
nor U3297 (N_3297,In_793,In_481);
nand U3298 (N_3298,In_656,In_170);
and U3299 (N_3299,In_681,In_138);
nor U3300 (N_3300,In_762,In_390);
xnor U3301 (N_3301,In_162,In_936);
nor U3302 (N_3302,In_840,In_611);
nor U3303 (N_3303,In_32,In_683);
nand U3304 (N_3304,In_542,In_42);
and U3305 (N_3305,In_205,In_170);
or U3306 (N_3306,In_267,In_545);
nand U3307 (N_3307,In_203,In_552);
nor U3308 (N_3308,In_661,In_742);
nor U3309 (N_3309,In_57,In_467);
or U3310 (N_3310,In_203,In_789);
or U3311 (N_3311,In_531,In_643);
and U3312 (N_3312,In_194,In_142);
xor U3313 (N_3313,In_520,In_338);
nor U3314 (N_3314,In_559,In_236);
or U3315 (N_3315,In_449,In_855);
nand U3316 (N_3316,In_427,In_256);
xnor U3317 (N_3317,In_320,In_896);
or U3318 (N_3318,In_974,In_303);
and U3319 (N_3319,In_331,In_795);
nor U3320 (N_3320,In_961,In_522);
and U3321 (N_3321,In_663,In_332);
and U3322 (N_3322,In_865,In_633);
nand U3323 (N_3323,In_28,In_848);
nand U3324 (N_3324,In_715,In_486);
or U3325 (N_3325,In_24,In_3);
nor U3326 (N_3326,In_10,In_573);
or U3327 (N_3327,In_252,In_120);
nor U3328 (N_3328,In_893,In_318);
xnor U3329 (N_3329,In_450,In_455);
nand U3330 (N_3330,In_933,In_78);
xnor U3331 (N_3331,In_868,In_713);
nor U3332 (N_3332,In_990,In_521);
nand U3333 (N_3333,In_443,In_733);
nand U3334 (N_3334,In_202,In_359);
or U3335 (N_3335,In_626,In_992);
and U3336 (N_3336,In_782,In_613);
or U3337 (N_3337,In_862,In_288);
nor U3338 (N_3338,In_901,In_281);
nor U3339 (N_3339,In_261,In_126);
xnor U3340 (N_3340,In_166,In_363);
nand U3341 (N_3341,In_124,In_171);
xor U3342 (N_3342,In_548,In_673);
nand U3343 (N_3343,In_612,In_16);
nand U3344 (N_3344,In_312,In_650);
xnor U3345 (N_3345,In_180,In_614);
nor U3346 (N_3346,In_799,In_810);
and U3347 (N_3347,In_172,In_613);
nor U3348 (N_3348,In_156,In_249);
xor U3349 (N_3349,In_208,In_321);
nand U3350 (N_3350,In_603,In_698);
nor U3351 (N_3351,In_779,In_364);
or U3352 (N_3352,In_573,In_167);
and U3353 (N_3353,In_931,In_112);
nand U3354 (N_3354,In_806,In_182);
nor U3355 (N_3355,In_805,In_256);
nor U3356 (N_3356,In_869,In_35);
and U3357 (N_3357,In_85,In_51);
xor U3358 (N_3358,In_119,In_851);
and U3359 (N_3359,In_838,In_758);
nand U3360 (N_3360,In_449,In_502);
nor U3361 (N_3361,In_558,In_161);
nand U3362 (N_3362,In_27,In_58);
xor U3363 (N_3363,In_70,In_485);
or U3364 (N_3364,In_873,In_99);
nand U3365 (N_3365,In_868,In_24);
or U3366 (N_3366,In_131,In_910);
xnor U3367 (N_3367,In_179,In_481);
and U3368 (N_3368,In_762,In_566);
and U3369 (N_3369,In_695,In_493);
or U3370 (N_3370,In_417,In_80);
xor U3371 (N_3371,In_777,In_918);
nor U3372 (N_3372,In_466,In_541);
and U3373 (N_3373,In_979,In_915);
nand U3374 (N_3374,In_546,In_384);
and U3375 (N_3375,In_920,In_913);
nor U3376 (N_3376,In_304,In_208);
or U3377 (N_3377,In_768,In_46);
nor U3378 (N_3378,In_387,In_505);
or U3379 (N_3379,In_640,In_551);
and U3380 (N_3380,In_879,In_431);
and U3381 (N_3381,In_762,In_668);
nand U3382 (N_3382,In_258,In_756);
nand U3383 (N_3383,In_382,In_48);
and U3384 (N_3384,In_741,In_456);
and U3385 (N_3385,In_525,In_909);
or U3386 (N_3386,In_364,In_358);
nor U3387 (N_3387,In_454,In_611);
nand U3388 (N_3388,In_918,In_747);
or U3389 (N_3389,In_603,In_451);
nand U3390 (N_3390,In_313,In_639);
or U3391 (N_3391,In_480,In_220);
and U3392 (N_3392,In_389,In_92);
nand U3393 (N_3393,In_55,In_865);
nor U3394 (N_3394,In_3,In_14);
xnor U3395 (N_3395,In_563,In_978);
nor U3396 (N_3396,In_854,In_609);
nor U3397 (N_3397,In_820,In_94);
nor U3398 (N_3398,In_948,In_557);
nor U3399 (N_3399,In_16,In_224);
nand U3400 (N_3400,In_447,In_86);
nand U3401 (N_3401,In_276,In_756);
nand U3402 (N_3402,In_690,In_62);
nor U3403 (N_3403,In_888,In_22);
nor U3404 (N_3404,In_674,In_523);
and U3405 (N_3405,In_740,In_557);
and U3406 (N_3406,In_453,In_169);
nand U3407 (N_3407,In_657,In_786);
nor U3408 (N_3408,In_915,In_450);
nor U3409 (N_3409,In_702,In_559);
xor U3410 (N_3410,In_921,In_106);
and U3411 (N_3411,In_247,In_255);
and U3412 (N_3412,In_896,In_609);
xnor U3413 (N_3413,In_984,In_105);
nor U3414 (N_3414,In_708,In_876);
and U3415 (N_3415,In_204,In_281);
nand U3416 (N_3416,In_850,In_912);
xor U3417 (N_3417,In_470,In_388);
xor U3418 (N_3418,In_437,In_872);
and U3419 (N_3419,In_563,In_232);
xor U3420 (N_3420,In_462,In_783);
nand U3421 (N_3421,In_796,In_497);
xor U3422 (N_3422,In_622,In_441);
or U3423 (N_3423,In_968,In_690);
nand U3424 (N_3424,In_348,In_35);
or U3425 (N_3425,In_766,In_223);
nor U3426 (N_3426,In_143,In_224);
xnor U3427 (N_3427,In_758,In_694);
nand U3428 (N_3428,In_34,In_525);
and U3429 (N_3429,In_59,In_709);
nor U3430 (N_3430,In_812,In_410);
nand U3431 (N_3431,In_917,In_222);
and U3432 (N_3432,In_857,In_176);
or U3433 (N_3433,In_967,In_831);
nor U3434 (N_3434,In_191,In_692);
or U3435 (N_3435,In_29,In_807);
nand U3436 (N_3436,In_872,In_54);
nor U3437 (N_3437,In_126,In_436);
nor U3438 (N_3438,In_350,In_149);
and U3439 (N_3439,In_812,In_418);
nor U3440 (N_3440,In_931,In_510);
and U3441 (N_3441,In_895,In_180);
xor U3442 (N_3442,In_234,In_654);
nor U3443 (N_3443,In_440,In_256);
nor U3444 (N_3444,In_279,In_801);
xor U3445 (N_3445,In_557,In_108);
nor U3446 (N_3446,In_346,In_277);
xnor U3447 (N_3447,In_330,In_463);
and U3448 (N_3448,In_779,In_652);
xor U3449 (N_3449,In_999,In_978);
xnor U3450 (N_3450,In_348,In_326);
xnor U3451 (N_3451,In_111,In_173);
or U3452 (N_3452,In_80,In_991);
nor U3453 (N_3453,In_541,In_522);
and U3454 (N_3454,In_641,In_393);
and U3455 (N_3455,In_893,In_920);
xnor U3456 (N_3456,In_288,In_292);
nand U3457 (N_3457,In_636,In_906);
nand U3458 (N_3458,In_498,In_907);
or U3459 (N_3459,In_26,In_778);
or U3460 (N_3460,In_842,In_389);
nand U3461 (N_3461,In_979,In_129);
nand U3462 (N_3462,In_791,In_755);
and U3463 (N_3463,In_169,In_486);
xor U3464 (N_3464,In_938,In_939);
xor U3465 (N_3465,In_615,In_476);
and U3466 (N_3466,In_254,In_713);
nor U3467 (N_3467,In_893,In_175);
and U3468 (N_3468,In_26,In_651);
and U3469 (N_3469,In_886,In_344);
or U3470 (N_3470,In_648,In_944);
nand U3471 (N_3471,In_35,In_253);
nand U3472 (N_3472,In_735,In_816);
or U3473 (N_3473,In_197,In_517);
and U3474 (N_3474,In_229,In_301);
and U3475 (N_3475,In_165,In_307);
nand U3476 (N_3476,In_766,In_48);
nand U3477 (N_3477,In_776,In_240);
and U3478 (N_3478,In_90,In_321);
xnor U3479 (N_3479,In_81,In_861);
nand U3480 (N_3480,In_137,In_524);
nor U3481 (N_3481,In_781,In_269);
xor U3482 (N_3482,In_827,In_282);
or U3483 (N_3483,In_303,In_298);
nor U3484 (N_3484,In_713,In_835);
and U3485 (N_3485,In_924,In_849);
nor U3486 (N_3486,In_19,In_686);
nand U3487 (N_3487,In_59,In_698);
nor U3488 (N_3488,In_686,In_147);
or U3489 (N_3489,In_247,In_403);
nand U3490 (N_3490,In_427,In_659);
xnor U3491 (N_3491,In_433,In_230);
and U3492 (N_3492,In_370,In_909);
xnor U3493 (N_3493,In_589,In_527);
nand U3494 (N_3494,In_381,In_32);
or U3495 (N_3495,In_70,In_176);
nor U3496 (N_3496,In_502,In_669);
or U3497 (N_3497,In_757,In_191);
or U3498 (N_3498,In_250,In_288);
or U3499 (N_3499,In_517,In_118);
xnor U3500 (N_3500,In_602,In_143);
nand U3501 (N_3501,In_44,In_587);
nand U3502 (N_3502,In_132,In_703);
and U3503 (N_3503,In_970,In_205);
and U3504 (N_3504,In_564,In_874);
nor U3505 (N_3505,In_972,In_788);
nand U3506 (N_3506,In_276,In_381);
or U3507 (N_3507,In_133,In_856);
nand U3508 (N_3508,In_285,In_560);
nand U3509 (N_3509,In_786,In_71);
xnor U3510 (N_3510,In_221,In_522);
and U3511 (N_3511,In_839,In_381);
and U3512 (N_3512,In_900,In_385);
xor U3513 (N_3513,In_912,In_323);
xnor U3514 (N_3514,In_739,In_86);
xor U3515 (N_3515,In_366,In_323);
and U3516 (N_3516,In_565,In_625);
or U3517 (N_3517,In_617,In_344);
nor U3518 (N_3518,In_738,In_372);
nor U3519 (N_3519,In_953,In_363);
nand U3520 (N_3520,In_868,In_684);
nand U3521 (N_3521,In_904,In_968);
nor U3522 (N_3522,In_23,In_635);
nand U3523 (N_3523,In_207,In_22);
nand U3524 (N_3524,In_509,In_595);
nand U3525 (N_3525,In_271,In_948);
and U3526 (N_3526,In_454,In_936);
xor U3527 (N_3527,In_769,In_564);
or U3528 (N_3528,In_752,In_98);
or U3529 (N_3529,In_554,In_641);
or U3530 (N_3530,In_417,In_275);
nand U3531 (N_3531,In_14,In_942);
nor U3532 (N_3532,In_426,In_301);
and U3533 (N_3533,In_186,In_175);
nor U3534 (N_3534,In_263,In_374);
or U3535 (N_3535,In_888,In_910);
or U3536 (N_3536,In_596,In_350);
nand U3537 (N_3537,In_367,In_687);
nand U3538 (N_3538,In_898,In_703);
xor U3539 (N_3539,In_561,In_318);
nand U3540 (N_3540,In_366,In_929);
nand U3541 (N_3541,In_4,In_72);
xor U3542 (N_3542,In_121,In_417);
nand U3543 (N_3543,In_401,In_957);
and U3544 (N_3544,In_635,In_396);
nand U3545 (N_3545,In_823,In_187);
nor U3546 (N_3546,In_601,In_452);
xor U3547 (N_3547,In_981,In_525);
nand U3548 (N_3548,In_204,In_401);
and U3549 (N_3549,In_478,In_66);
nor U3550 (N_3550,In_220,In_359);
nor U3551 (N_3551,In_161,In_99);
or U3552 (N_3552,In_553,In_128);
xor U3553 (N_3553,In_980,In_303);
and U3554 (N_3554,In_484,In_802);
nand U3555 (N_3555,In_646,In_420);
nand U3556 (N_3556,In_880,In_630);
nand U3557 (N_3557,In_681,In_406);
and U3558 (N_3558,In_367,In_374);
nand U3559 (N_3559,In_796,In_345);
nand U3560 (N_3560,In_734,In_901);
or U3561 (N_3561,In_276,In_13);
and U3562 (N_3562,In_373,In_271);
xor U3563 (N_3563,In_311,In_880);
and U3564 (N_3564,In_991,In_23);
or U3565 (N_3565,In_843,In_213);
nand U3566 (N_3566,In_950,In_687);
nor U3567 (N_3567,In_790,In_72);
nor U3568 (N_3568,In_725,In_369);
nor U3569 (N_3569,In_960,In_340);
or U3570 (N_3570,In_445,In_123);
nand U3571 (N_3571,In_764,In_608);
or U3572 (N_3572,In_479,In_833);
and U3573 (N_3573,In_354,In_752);
nand U3574 (N_3574,In_142,In_801);
nand U3575 (N_3575,In_737,In_139);
nor U3576 (N_3576,In_277,In_584);
nand U3577 (N_3577,In_134,In_680);
or U3578 (N_3578,In_269,In_252);
nor U3579 (N_3579,In_91,In_482);
and U3580 (N_3580,In_465,In_471);
nand U3581 (N_3581,In_942,In_462);
nor U3582 (N_3582,In_437,In_682);
and U3583 (N_3583,In_978,In_464);
nor U3584 (N_3584,In_53,In_910);
or U3585 (N_3585,In_985,In_917);
nand U3586 (N_3586,In_949,In_279);
nand U3587 (N_3587,In_391,In_964);
nor U3588 (N_3588,In_841,In_973);
or U3589 (N_3589,In_584,In_440);
xnor U3590 (N_3590,In_858,In_773);
nand U3591 (N_3591,In_201,In_39);
nand U3592 (N_3592,In_843,In_808);
or U3593 (N_3593,In_611,In_579);
nand U3594 (N_3594,In_905,In_439);
xnor U3595 (N_3595,In_46,In_276);
and U3596 (N_3596,In_996,In_618);
nand U3597 (N_3597,In_490,In_761);
xnor U3598 (N_3598,In_58,In_17);
xnor U3599 (N_3599,In_95,In_349);
and U3600 (N_3600,In_687,In_386);
xnor U3601 (N_3601,In_374,In_669);
nand U3602 (N_3602,In_186,In_667);
xnor U3603 (N_3603,In_602,In_5);
or U3604 (N_3604,In_35,In_817);
and U3605 (N_3605,In_663,In_423);
nand U3606 (N_3606,In_402,In_890);
and U3607 (N_3607,In_595,In_14);
nand U3608 (N_3608,In_548,In_815);
and U3609 (N_3609,In_168,In_319);
or U3610 (N_3610,In_886,In_44);
nor U3611 (N_3611,In_119,In_332);
and U3612 (N_3612,In_546,In_30);
nor U3613 (N_3613,In_306,In_760);
nor U3614 (N_3614,In_620,In_726);
or U3615 (N_3615,In_572,In_159);
and U3616 (N_3616,In_934,In_392);
nor U3617 (N_3617,In_760,In_989);
xor U3618 (N_3618,In_761,In_209);
xor U3619 (N_3619,In_126,In_121);
and U3620 (N_3620,In_766,In_68);
nand U3621 (N_3621,In_3,In_802);
nand U3622 (N_3622,In_934,In_798);
and U3623 (N_3623,In_450,In_276);
nand U3624 (N_3624,In_306,In_651);
xnor U3625 (N_3625,In_421,In_487);
nor U3626 (N_3626,In_213,In_311);
xor U3627 (N_3627,In_484,In_608);
nand U3628 (N_3628,In_843,In_961);
or U3629 (N_3629,In_137,In_346);
or U3630 (N_3630,In_718,In_529);
nand U3631 (N_3631,In_868,In_527);
nand U3632 (N_3632,In_431,In_307);
or U3633 (N_3633,In_377,In_575);
nor U3634 (N_3634,In_405,In_956);
nand U3635 (N_3635,In_98,In_92);
xnor U3636 (N_3636,In_270,In_965);
xnor U3637 (N_3637,In_958,In_547);
and U3638 (N_3638,In_266,In_866);
nor U3639 (N_3639,In_764,In_297);
and U3640 (N_3640,In_195,In_720);
xnor U3641 (N_3641,In_225,In_235);
or U3642 (N_3642,In_841,In_798);
nor U3643 (N_3643,In_256,In_972);
and U3644 (N_3644,In_56,In_344);
xnor U3645 (N_3645,In_374,In_885);
nand U3646 (N_3646,In_143,In_97);
and U3647 (N_3647,In_772,In_526);
nor U3648 (N_3648,In_312,In_481);
nor U3649 (N_3649,In_392,In_408);
nor U3650 (N_3650,In_501,In_806);
nand U3651 (N_3651,In_254,In_835);
xor U3652 (N_3652,In_666,In_120);
nor U3653 (N_3653,In_62,In_693);
nand U3654 (N_3654,In_614,In_349);
nor U3655 (N_3655,In_32,In_405);
xnor U3656 (N_3656,In_40,In_188);
and U3657 (N_3657,In_445,In_790);
nor U3658 (N_3658,In_796,In_97);
or U3659 (N_3659,In_830,In_444);
xor U3660 (N_3660,In_662,In_608);
xor U3661 (N_3661,In_633,In_308);
nor U3662 (N_3662,In_932,In_399);
nand U3663 (N_3663,In_893,In_304);
nor U3664 (N_3664,In_239,In_357);
nor U3665 (N_3665,In_104,In_373);
nand U3666 (N_3666,In_92,In_155);
nor U3667 (N_3667,In_429,In_841);
and U3668 (N_3668,In_672,In_390);
and U3669 (N_3669,In_970,In_128);
and U3670 (N_3670,In_497,In_561);
nand U3671 (N_3671,In_283,In_115);
and U3672 (N_3672,In_135,In_647);
nor U3673 (N_3673,In_990,In_612);
nor U3674 (N_3674,In_81,In_574);
and U3675 (N_3675,In_252,In_66);
or U3676 (N_3676,In_536,In_546);
nor U3677 (N_3677,In_569,In_408);
and U3678 (N_3678,In_127,In_748);
nand U3679 (N_3679,In_880,In_730);
and U3680 (N_3680,In_408,In_88);
or U3681 (N_3681,In_954,In_708);
xor U3682 (N_3682,In_755,In_629);
xnor U3683 (N_3683,In_659,In_14);
xnor U3684 (N_3684,In_909,In_328);
nor U3685 (N_3685,In_616,In_305);
or U3686 (N_3686,In_343,In_590);
and U3687 (N_3687,In_846,In_296);
or U3688 (N_3688,In_436,In_184);
nand U3689 (N_3689,In_503,In_656);
xor U3690 (N_3690,In_777,In_374);
and U3691 (N_3691,In_17,In_120);
nand U3692 (N_3692,In_584,In_478);
and U3693 (N_3693,In_67,In_381);
and U3694 (N_3694,In_104,In_129);
or U3695 (N_3695,In_316,In_989);
and U3696 (N_3696,In_314,In_852);
nor U3697 (N_3697,In_270,In_332);
xnor U3698 (N_3698,In_167,In_830);
xor U3699 (N_3699,In_272,In_130);
nor U3700 (N_3700,In_548,In_972);
or U3701 (N_3701,In_966,In_289);
nor U3702 (N_3702,In_428,In_590);
xor U3703 (N_3703,In_490,In_821);
nand U3704 (N_3704,In_604,In_755);
xnor U3705 (N_3705,In_897,In_874);
nor U3706 (N_3706,In_105,In_647);
or U3707 (N_3707,In_285,In_779);
nor U3708 (N_3708,In_143,In_279);
nor U3709 (N_3709,In_342,In_362);
and U3710 (N_3710,In_200,In_650);
and U3711 (N_3711,In_770,In_585);
or U3712 (N_3712,In_923,In_171);
nand U3713 (N_3713,In_361,In_237);
nor U3714 (N_3714,In_595,In_103);
nor U3715 (N_3715,In_617,In_224);
nand U3716 (N_3716,In_652,In_384);
and U3717 (N_3717,In_727,In_832);
nand U3718 (N_3718,In_602,In_106);
or U3719 (N_3719,In_599,In_889);
or U3720 (N_3720,In_896,In_926);
nand U3721 (N_3721,In_470,In_492);
nor U3722 (N_3722,In_668,In_196);
and U3723 (N_3723,In_665,In_600);
and U3724 (N_3724,In_303,In_375);
or U3725 (N_3725,In_762,In_346);
and U3726 (N_3726,In_417,In_795);
and U3727 (N_3727,In_11,In_255);
or U3728 (N_3728,In_143,In_707);
or U3729 (N_3729,In_75,In_976);
nor U3730 (N_3730,In_83,In_732);
xnor U3731 (N_3731,In_195,In_663);
or U3732 (N_3732,In_597,In_197);
nand U3733 (N_3733,In_871,In_501);
and U3734 (N_3734,In_139,In_409);
nand U3735 (N_3735,In_631,In_91);
xnor U3736 (N_3736,In_305,In_96);
and U3737 (N_3737,In_697,In_906);
and U3738 (N_3738,In_629,In_490);
nor U3739 (N_3739,In_755,In_740);
or U3740 (N_3740,In_160,In_613);
xnor U3741 (N_3741,In_25,In_658);
nor U3742 (N_3742,In_708,In_548);
or U3743 (N_3743,In_256,In_437);
nand U3744 (N_3744,In_271,In_642);
or U3745 (N_3745,In_398,In_788);
nand U3746 (N_3746,In_17,In_251);
nand U3747 (N_3747,In_749,In_70);
or U3748 (N_3748,In_666,In_340);
and U3749 (N_3749,In_182,In_633);
xnor U3750 (N_3750,In_653,In_827);
or U3751 (N_3751,In_14,In_708);
nand U3752 (N_3752,In_324,In_599);
xnor U3753 (N_3753,In_956,In_309);
or U3754 (N_3754,In_273,In_688);
nand U3755 (N_3755,In_901,In_968);
nand U3756 (N_3756,In_525,In_321);
nand U3757 (N_3757,In_294,In_467);
or U3758 (N_3758,In_695,In_264);
or U3759 (N_3759,In_418,In_851);
xor U3760 (N_3760,In_773,In_455);
xor U3761 (N_3761,In_336,In_639);
xnor U3762 (N_3762,In_592,In_611);
or U3763 (N_3763,In_414,In_461);
nand U3764 (N_3764,In_28,In_711);
nor U3765 (N_3765,In_127,In_560);
and U3766 (N_3766,In_510,In_596);
and U3767 (N_3767,In_986,In_769);
nor U3768 (N_3768,In_508,In_263);
xor U3769 (N_3769,In_458,In_217);
and U3770 (N_3770,In_183,In_678);
or U3771 (N_3771,In_637,In_587);
nor U3772 (N_3772,In_268,In_324);
nand U3773 (N_3773,In_115,In_874);
or U3774 (N_3774,In_947,In_731);
nor U3775 (N_3775,In_413,In_183);
nor U3776 (N_3776,In_94,In_616);
xor U3777 (N_3777,In_274,In_827);
or U3778 (N_3778,In_407,In_312);
or U3779 (N_3779,In_0,In_699);
or U3780 (N_3780,In_622,In_402);
nor U3781 (N_3781,In_448,In_479);
or U3782 (N_3782,In_739,In_159);
nor U3783 (N_3783,In_136,In_200);
nor U3784 (N_3784,In_596,In_313);
xor U3785 (N_3785,In_304,In_485);
xnor U3786 (N_3786,In_267,In_413);
nand U3787 (N_3787,In_381,In_454);
xnor U3788 (N_3788,In_226,In_444);
nand U3789 (N_3789,In_435,In_679);
or U3790 (N_3790,In_152,In_431);
and U3791 (N_3791,In_228,In_218);
or U3792 (N_3792,In_795,In_55);
and U3793 (N_3793,In_66,In_200);
or U3794 (N_3794,In_488,In_151);
nor U3795 (N_3795,In_695,In_586);
xor U3796 (N_3796,In_451,In_255);
or U3797 (N_3797,In_243,In_357);
or U3798 (N_3798,In_16,In_641);
nor U3799 (N_3799,In_191,In_143);
xor U3800 (N_3800,In_683,In_101);
xor U3801 (N_3801,In_402,In_846);
nand U3802 (N_3802,In_289,In_711);
xor U3803 (N_3803,In_746,In_46);
nand U3804 (N_3804,In_874,In_937);
and U3805 (N_3805,In_244,In_964);
nand U3806 (N_3806,In_874,In_682);
or U3807 (N_3807,In_398,In_288);
nand U3808 (N_3808,In_719,In_116);
and U3809 (N_3809,In_872,In_470);
and U3810 (N_3810,In_515,In_24);
and U3811 (N_3811,In_227,In_462);
nand U3812 (N_3812,In_417,In_214);
and U3813 (N_3813,In_212,In_205);
nand U3814 (N_3814,In_568,In_334);
xnor U3815 (N_3815,In_342,In_622);
nor U3816 (N_3816,In_998,In_174);
nand U3817 (N_3817,In_523,In_656);
nand U3818 (N_3818,In_871,In_406);
and U3819 (N_3819,In_695,In_491);
or U3820 (N_3820,In_94,In_569);
nor U3821 (N_3821,In_425,In_842);
nor U3822 (N_3822,In_951,In_883);
and U3823 (N_3823,In_917,In_770);
and U3824 (N_3824,In_738,In_385);
xor U3825 (N_3825,In_694,In_183);
or U3826 (N_3826,In_474,In_30);
and U3827 (N_3827,In_503,In_900);
or U3828 (N_3828,In_422,In_831);
or U3829 (N_3829,In_534,In_411);
nor U3830 (N_3830,In_170,In_716);
nand U3831 (N_3831,In_322,In_379);
or U3832 (N_3832,In_793,In_566);
and U3833 (N_3833,In_715,In_785);
or U3834 (N_3834,In_815,In_843);
nor U3835 (N_3835,In_113,In_61);
and U3836 (N_3836,In_373,In_181);
nand U3837 (N_3837,In_958,In_410);
or U3838 (N_3838,In_705,In_561);
xor U3839 (N_3839,In_679,In_552);
nand U3840 (N_3840,In_321,In_934);
or U3841 (N_3841,In_584,In_330);
or U3842 (N_3842,In_314,In_650);
xnor U3843 (N_3843,In_771,In_151);
nand U3844 (N_3844,In_238,In_400);
xor U3845 (N_3845,In_279,In_618);
nand U3846 (N_3846,In_496,In_483);
nor U3847 (N_3847,In_928,In_982);
or U3848 (N_3848,In_685,In_30);
nand U3849 (N_3849,In_217,In_873);
nor U3850 (N_3850,In_682,In_765);
xor U3851 (N_3851,In_784,In_918);
and U3852 (N_3852,In_618,In_822);
nand U3853 (N_3853,In_469,In_109);
or U3854 (N_3854,In_419,In_803);
or U3855 (N_3855,In_208,In_226);
nor U3856 (N_3856,In_718,In_916);
nand U3857 (N_3857,In_178,In_560);
nor U3858 (N_3858,In_376,In_220);
nand U3859 (N_3859,In_379,In_383);
xnor U3860 (N_3860,In_248,In_264);
or U3861 (N_3861,In_448,In_617);
nor U3862 (N_3862,In_883,In_31);
or U3863 (N_3863,In_14,In_707);
or U3864 (N_3864,In_39,In_576);
nand U3865 (N_3865,In_298,In_130);
nor U3866 (N_3866,In_370,In_723);
and U3867 (N_3867,In_35,In_176);
and U3868 (N_3868,In_870,In_223);
or U3869 (N_3869,In_495,In_700);
or U3870 (N_3870,In_490,In_469);
nor U3871 (N_3871,In_654,In_933);
and U3872 (N_3872,In_637,In_311);
xnor U3873 (N_3873,In_543,In_54);
nor U3874 (N_3874,In_208,In_383);
xor U3875 (N_3875,In_258,In_242);
xor U3876 (N_3876,In_249,In_149);
nand U3877 (N_3877,In_6,In_763);
xor U3878 (N_3878,In_342,In_207);
and U3879 (N_3879,In_383,In_972);
xor U3880 (N_3880,In_453,In_175);
nor U3881 (N_3881,In_325,In_109);
xnor U3882 (N_3882,In_148,In_538);
nand U3883 (N_3883,In_16,In_589);
xor U3884 (N_3884,In_842,In_322);
nor U3885 (N_3885,In_955,In_629);
or U3886 (N_3886,In_564,In_94);
or U3887 (N_3887,In_911,In_825);
or U3888 (N_3888,In_223,In_694);
nand U3889 (N_3889,In_830,In_603);
and U3890 (N_3890,In_372,In_196);
nor U3891 (N_3891,In_426,In_341);
xor U3892 (N_3892,In_28,In_789);
and U3893 (N_3893,In_173,In_977);
nand U3894 (N_3894,In_474,In_25);
and U3895 (N_3895,In_258,In_309);
nor U3896 (N_3896,In_808,In_57);
or U3897 (N_3897,In_756,In_701);
nor U3898 (N_3898,In_207,In_498);
or U3899 (N_3899,In_592,In_392);
nand U3900 (N_3900,In_819,In_569);
nor U3901 (N_3901,In_151,In_63);
xor U3902 (N_3902,In_108,In_558);
xnor U3903 (N_3903,In_844,In_821);
nand U3904 (N_3904,In_930,In_95);
nor U3905 (N_3905,In_458,In_171);
or U3906 (N_3906,In_563,In_721);
nor U3907 (N_3907,In_144,In_980);
nand U3908 (N_3908,In_765,In_329);
nor U3909 (N_3909,In_45,In_466);
and U3910 (N_3910,In_15,In_347);
and U3911 (N_3911,In_105,In_230);
or U3912 (N_3912,In_188,In_62);
and U3913 (N_3913,In_12,In_877);
nand U3914 (N_3914,In_877,In_662);
nor U3915 (N_3915,In_828,In_538);
nand U3916 (N_3916,In_334,In_473);
xnor U3917 (N_3917,In_690,In_588);
nand U3918 (N_3918,In_878,In_845);
xnor U3919 (N_3919,In_502,In_522);
xor U3920 (N_3920,In_164,In_92);
xor U3921 (N_3921,In_359,In_419);
or U3922 (N_3922,In_710,In_565);
nand U3923 (N_3923,In_923,In_190);
nand U3924 (N_3924,In_746,In_710);
nor U3925 (N_3925,In_495,In_961);
and U3926 (N_3926,In_927,In_551);
or U3927 (N_3927,In_789,In_614);
and U3928 (N_3928,In_700,In_247);
and U3929 (N_3929,In_771,In_813);
nand U3930 (N_3930,In_960,In_520);
and U3931 (N_3931,In_83,In_51);
or U3932 (N_3932,In_453,In_445);
nand U3933 (N_3933,In_325,In_6);
nor U3934 (N_3934,In_37,In_296);
nand U3935 (N_3935,In_40,In_742);
nor U3936 (N_3936,In_121,In_472);
or U3937 (N_3937,In_970,In_962);
nand U3938 (N_3938,In_459,In_52);
or U3939 (N_3939,In_398,In_910);
nor U3940 (N_3940,In_549,In_725);
or U3941 (N_3941,In_857,In_627);
or U3942 (N_3942,In_969,In_714);
or U3943 (N_3943,In_571,In_66);
or U3944 (N_3944,In_874,In_869);
and U3945 (N_3945,In_776,In_124);
nor U3946 (N_3946,In_548,In_32);
xor U3947 (N_3947,In_70,In_915);
nor U3948 (N_3948,In_750,In_468);
and U3949 (N_3949,In_236,In_425);
or U3950 (N_3950,In_935,In_483);
nand U3951 (N_3951,In_547,In_190);
or U3952 (N_3952,In_788,In_397);
nor U3953 (N_3953,In_705,In_35);
nor U3954 (N_3954,In_610,In_619);
and U3955 (N_3955,In_564,In_732);
xor U3956 (N_3956,In_848,In_200);
xnor U3957 (N_3957,In_503,In_145);
nand U3958 (N_3958,In_657,In_716);
nand U3959 (N_3959,In_921,In_831);
nand U3960 (N_3960,In_563,In_691);
and U3961 (N_3961,In_237,In_44);
and U3962 (N_3962,In_69,In_67);
xor U3963 (N_3963,In_129,In_404);
nor U3964 (N_3964,In_131,In_937);
or U3965 (N_3965,In_485,In_918);
nand U3966 (N_3966,In_350,In_824);
xor U3967 (N_3967,In_238,In_346);
and U3968 (N_3968,In_168,In_962);
or U3969 (N_3969,In_325,In_706);
and U3970 (N_3970,In_950,In_205);
xnor U3971 (N_3971,In_456,In_498);
nand U3972 (N_3972,In_103,In_786);
or U3973 (N_3973,In_319,In_410);
and U3974 (N_3974,In_565,In_727);
and U3975 (N_3975,In_922,In_944);
and U3976 (N_3976,In_833,In_626);
and U3977 (N_3977,In_833,In_985);
nand U3978 (N_3978,In_480,In_362);
or U3979 (N_3979,In_970,In_264);
or U3980 (N_3980,In_173,In_420);
xnor U3981 (N_3981,In_707,In_177);
nand U3982 (N_3982,In_994,In_691);
or U3983 (N_3983,In_427,In_287);
nor U3984 (N_3984,In_907,In_685);
nor U3985 (N_3985,In_835,In_895);
xor U3986 (N_3986,In_828,In_486);
or U3987 (N_3987,In_377,In_302);
or U3988 (N_3988,In_264,In_241);
and U3989 (N_3989,In_712,In_245);
and U3990 (N_3990,In_102,In_258);
or U3991 (N_3991,In_337,In_62);
nor U3992 (N_3992,In_121,In_330);
xor U3993 (N_3993,In_241,In_612);
nor U3994 (N_3994,In_211,In_723);
xnor U3995 (N_3995,In_252,In_13);
nor U3996 (N_3996,In_575,In_641);
xor U3997 (N_3997,In_802,In_549);
xor U3998 (N_3998,In_749,In_848);
and U3999 (N_3999,In_547,In_315);
or U4000 (N_4000,In_924,In_877);
or U4001 (N_4001,In_245,In_228);
and U4002 (N_4002,In_497,In_317);
xor U4003 (N_4003,In_391,In_353);
xnor U4004 (N_4004,In_233,In_109);
nor U4005 (N_4005,In_754,In_868);
and U4006 (N_4006,In_249,In_183);
or U4007 (N_4007,In_738,In_854);
xor U4008 (N_4008,In_189,In_388);
and U4009 (N_4009,In_937,In_540);
xnor U4010 (N_4010,In_92,In_759);
nand U4011 (N_4011,In_716,In_242);
nor U4012 (N_4012,In_832,In_844);
nand U4013 (N_4013,In_926,In_872);
and U4014 (N_4014,In_271,In_361);
or U4015 (N_4015,In_145,In_929);
nand U4016 (N_4016,In_804,In_422);
nor U4017 (N_4017,In_511,In_884);
nor U4018 (N_4018,In_541,In_825);
and U4019 (N_4019,In_371,In_507);
nand U4020 (N_4020,In_547,In_698);
nand U4021 (N_4021,In_709,In_598);
or U4022 (N_4022,In_826,In_346);
nor U4023 (N_4023,In_422,In_953);
nor U4024 (N_4024,In_351,In_888);
nor U4025 (N_4025,In_467,In_971);
nand U4026 (N_4026,In_370,In_725);
and U4027 (N_4027,In_123,In_40);
or U4028 (N_4028,In_667,In_110);
nor U4029 (N_4029,In_940,In_780);
xnor U4030 (N_4030,In_67,In_369);
and U4031 (N_4031,In_356,In_655);
nor U4032 (N_4032,In_275,In_526);
or U4033 (N_4033,In_288,In_4);
xor U4034 (N_4034,In_12,In_605);
xor U4035 (N_4035,In_577,In_9);
xnor U4036 (N_4036,In_942,In_861);
xnor U4037 (N_4037,In_729,In_534);
nand U4038 (N_4038,In_967,In_329);
nor U4039 (N_4039,In_190,In_777);
nor U4040 (N_4040,In_19,In_748);
nand U4041 (N_4041,In_276,In_554);
nand U4042 (N_4042,In_263,In_557);
nor U4043 (N_4043,In_207,In_357);
nor U4044 (N_4044,In_870,In_752);
xor U4045 (N_4045,In_667,In_873);
xnor U4046 (N_4046,In_25,In_768);
nand U4047 (N_4047,In_765,In_30);
xor U4048 (N_4048,In_252,In_798);
xor U4049 (N_4049,In_910,In_934);
nand U4050 (N_4050,In_553,In_822);
or U4051 (N_4051,In_607,In_438);
or U4052 (N_4052,In_450,In_89);
xnor U4053 (N_4053,In_267,In_676);
nand U4054 (N_4054,In_749,In_428);
xor U4055 (N_4055,In_136,In_175);
and U4056 (N_4056,In_273,In_800);
xor U4057 (N_4057,In_669,In_631);
and U4058 (N_4058,In_278,In_176);
or U4059 (N_4059,In_196,In_857);
xor U4060 (N_4060,In_794,In_164);
nand U4061 (N_4061,In_733,In_244);
nor U4062 (N_4062,In_299,In_625);
xor U4063 (N_4063,In_307,In_881);
xor U4064 (N_4064,In_592,In_367);
nor U4065 (N_4065,In_219,In_634);
nor U4066 (N_4066,In_319,In_524);
xnor U4067 (N_4067,In_847,In_981);
or U4068 (N_4068,In_421,In_610);
nand U4069 (N_4069,In_904,In_164);
or U4070 (N_4070,In_32,In_133);
or U4071 (N_4071,In_346,In_175);
nand U4072 (N_4072,In_738,In_104);
nand U4073 (N_4073,In_269,In_734);
nor U4074 (N_4074,In_743,In_4);
nand U4075 (N_4075,In_5,In_580);
and U4076 (N_4076,In_423,In_368);
xor U4077 (N_4077,In_961,In_436);
xnor U4078 (N_4078,In_341,In_623);
xnor U4079 (N_4079,In_361,In_252);
and U4080 (N_4080,In_606,In_763);
or U4081 (N_4081,In_656,In_219);
nand U4082 (N_4082,In_971,In_22);
or U4083 (N_4083,In_511,In_368);
or U4084 (N_4084,In_446,In_621);
nor U4085 (N_4085,In_379,In_541);
xor U4086 (N_4086,In_927,In_74);
and U4087 (N_4087,In_657,In_670);
and U4088 (N_4088,In_793,In_69);
nor U4089 (N_4089,In_525,In_344);
nor U4090 (N_4090,In_844,In_849);
nor U4091 (N_4091,In_6,In_156);
nand U4092 (N_4092,In_68,In_729);
and U4093 (N_4093,In_265,In_782);
and U4094 (N_4094,In_169,In_916);
and U4095 (N_4095,In_612,In_506);
nand U4096 (N_4096,In_487,In_778);
and U4097 (N_4097,In_634,In_785);
nand U4098 (N_4098,In_859,In_466);
or U4099 (N_4099,In_52,In_543);
or U4100 (N_4100,In_469,In_609);
and U4101 (N_4101,In_720,In_64);
and U4102 (N_4102,In_399,In_275);
nand U4103 (N_4103,In_482,In_553);
or U4104 (N_4104,In_568,In_947);
or U4105 (N_4105,In_998,In_977);
or U4106 (N_4106,In_861,In_622);
xor U4107 (N_4107,In_330,In_879);
nor U4108 (N_4108,In_407,In_232);
nor U4109 (N_4109,In_564,In_723);
nand U4110 (N_4110,In_17,In_898);
or U4111 (N_4111,In_134,In_908);
xor U4112 (N_4112,In_222,In_976);
or U4113 (N_4113,In_49,In_975);
nand U4114 (N_4114,In_716,In_671);
nor U4115 (N_4115,In_458,In_490);
and U4116 (N_4116,In_821,In_137);
or U4117 (N_4117,In_374,In_139);
and U4118 (N_4118,In_649,In_658);
or U4119 (N_4119,In_480,In_159);
and U4120 (N_4120,In_156,In_532);
or U4121 (N_4121,In_853,In_484);
xor U4122 (N_4122,In_282,In_665);
nand U4123 (N_4123,In_972,In_82);
xnor U4124 (N_4124,In_0,In_906);
nand U4125 (N_4125,In_607,In_225);
and U4126 (N_4126,In_965,In_574);
or U4127 (N_4127,In_472,In_755);
xor U4128 (N_4128,In_1,In_19);
nor U4129 (N_4129,In_897,In_915);
xnor U4130 (N_4130,In_64,In_532);
nand U4131 (N_4131,In_475,In_538);
nand U4132 (N_4132,In_695,In_923);
nor U4133 (N_4133,In_924,In_556);
nor U4134 (N_4134,In_518,In_813);
nor U4135 (N_4135,In_353,In_476);
nand U4136 (N_4136,In_227,In_375);
nor U4137 (N_4137,In_847,In_63);
nand U4138 (N_4138,In_181,In_695);
xnor U4139 (N_4139,In_773,In_810);
and U4140 (N_4140,In_266,In_780);
or U4141 (N_4141,In_239,In_905);
nand U4142 (N_4142,In_697,In_796);
xnor U4143 (N_4143,In_396,In_877);
xnor U4144 (N_4144,In_534,In_613);
nand U4145 (N_4145,In_971,In_777);
xor U4146 (N_4146,In_667,In_59);
xor U4147 (N_4147,In_384,In_441);
xnor U4148 (N_4148,In_593,In_112);
nor U4149 (N_4149,In_774,In_23);
xnor U4150 (N_4150,In_802,In_173);
or U4151 (N_4151,In_192,In_640);
nor U4152 (N_4152,In_855,In_338);
and U4153 (N_4153,In_252,In_314);
or U4154 (N_4154,In_276,In_546);
or U4155 (N_4155,In_88,In_845);
nor U4156 (N_4156,In_368,In_450);
xor U4157 (N_4157,In_172,In_559);
xnor U4158 (N_4158,In_345,In_712);
nand U4159 (N_4159,In_645,In_785);
or U4160 (N_4160,In_260,In_484);
or U4161 (N_4161,In_728,In_537);
nor U4162 (N_4162,In_955,In_276);
xor U4163 (N_4163,In_274,In_774);
nand U4164 (N_4164,In_527,In_309);
nand U4165 (N_4165,In_516,In_617);
xor U4166 (N_4166,In_159,In_532);
or U4167 (N_4167,In_547,In_374);
xnor U4168 (N_4168,In_573,In_61);
or U4169 (N_4169,In_836,In_990);
nor U4170 (N_4170,In_167,In_189);
xnor U4171 (N_4171,In_442,In_203);
and U4172 (N_4172,In_179,In_502);
nor U4173 (N_4173,In_190,In_965);
nand U4174 (N_4174,In_677,In_176);
xor U4175 (N_4175,In_738,In_667);
nand U4176 (N_4176,In_649,In_54);
nand U4177 (N_4177,In_749,In_810);
nand U4178 (N_4178,In_992,In_96);
and U4179 (N_4179,In_573,In_72);
or U4180 (N_4180,In_535,In_664);
xnor U4181 (N_4181,In_542,In_805);
nand U4182 (N_4182,In_700,In_958);
and U4183 (N_4183,In_171,In_205);
and U4184 (N_4184,In_867,In_565);
nand U4185 (N_4185,In_725,In_21);
nor U4186 (N_4186,In_838,In_655);
nand U4187 (N_4187,In_732,In_954);
or U4188 (N_4188,In_154,In_637);
and U4189 (N_4189,In_302,In_794);
nor U4190 (N_4190,In_832,In_8);
nor U4191 (N_4191,In_540,In_953);
or U4192 (N_4192,In_443,In_459);
nand U4193 (N_4193,In_127,In_832);
nand U4194 (N_4194,In_774,In_952);
xnor U4195 (N_4195,In_14,In_402);
nor U4196 (N_4196,In_495,In_818);
xnor U4197 (N_4197,In_105,In_28);
nand U4198 (N_4198,In_0,In_933);
nor U4199 (N_4199,In_956,In_914);
and U4200 (N_4200,In_743,In_868);
and U4201 (N_4201,In_498,In_520);
xor U4202 (N_4202,In_805,In_391);
xor U4203 (N_4203,In_131,In_354);
xor U4204 (N_4204,In_136,In_977);
and U4205 (N_4205,In_242,In_741);
nor U4206 (N_4206,In_718,In_411);
xnor U4207 (N_4207,In_665,In_55);
xnor U4208 (N_4208,In_374,In_14);
and U4209 (N_4209,In_903,In_460);
or U4210 (N_4210,In_837,In_750);
xnor U4211 (N_4211,In_156,In_137);
xnor U4212 (N_4212,In_399,In_941);
or U4213 (N_4213,In_941,In_895);
xor U4214 (N_4214,In_34,In_768);
nor U4215 (N_4215,In_542,In_828);
nor U4216 (N_4216,In_465,In_889);
or U4217 (N_4217,In_832,In_651);
nand U4218 (N_4218,In_636,In_985);
xnor U4219 (N_4219,In_21,In_607);
nand U4220 (N_4220,In_30,In_444);
nand U4221 (N_4221,In_723,In_872);
or U4222 (N_4222,In_628,In_588);
nand U4223 (N_4223,In_0,In_836);
and U4224 (N_4224,In_331,In_869);
nor U4225 (N_4225,In_712,In_261);
nor U4226 (N_4226,In_605,In_780);
or U4227 (N_4227,In_667,In_470);
nand U4228 (N_4228,In_213,In_584);
xor U4229 (N_4229,In_425,In_364);
nor U4230 (N_4230,In_696,In_324);
or U4231 (N_4231,In_590,In_808);
or U4232 (N_4232,In_41,In_809);
xnor U4233 (N_4233,In_586,In_574);
nor U4234 (N_4234,In_622,In_802);
or U4235 (N_4235,In_868,In_397);
nand U4236 (N_4236,In_356,In_5);
or U4237 (N_4237,In_726,In_309);
nand U4238 (N_4238,In_343,In_558);
and U4239 (N_4239,In_64,In_368);
or U4240 (N_4240,In_344,In_702);
nor U4241 (N_4241,In_289,In_251);
or U4242 (N_4242,In_944,In_483);
nor U4243 (N_4243,In_477,In_447);
or U4244 (N_4244,In_620,In_327);
nor U4245 (N_4245,In_303,In_427);
nor U4246 (N_4246,In_695,In_597);
nand U4247 (N_4247,In_780,In_260);
xnor U4248 (N_4248,In_177,In_421);
nor U4249 (N_4249,In_231,In_338);
and U4250 (N_4250,In_904,In_688);
xor U4251 (N_4251,In_554,In_710);
or U4252 (N_4252,In_284,In_641);
nand U4253 (N_4253,In_382,In_540);
nand U4254 (N_4254,In_339,In_555);
nand U4255 (N_4255,In_628,In_508);
and U4256 (N_4256,In_271,In_533);
nor U4257 (N_4257,In_951,In_824);
and U4258 (N_4258,In_8,In_400);
nor U4259 (N_4259,In_652,In_34);
or U4260 (N_4260,In_329,In_757);
xnor U4261 (N_4261,In_897,In_809);
or U4262 (N_4262,In_992,In_772);
or U4263 (N_4263,In_408,In_565);
nand U4264 (N_4264,In_683,In_30);
xnor U4265 (N_4265,In_606,In_956);
and U4266 (N_4266,In_264,In_588);
xor U4267 (N_4267,In_819,In_897);
nor U4268 (N_4268,In_664,In_126);
xor U4269 (N_4269,In_404,In_638);
or U4270 (N_4270,In_210,In_166);
nand U4271 (N_4271,In_784,In_905);
or U4272 (N_4272,In_706,In_753);
nand U4273 (N_4273,In_426,In_68);
or U4274 (N_4274,In_805,In_712);
and U4275 (N_4275,In_725,In_288);
xor U4276 (N_4276,In_397,In_863);
or U4277 (N_4277,In_519,In_862);
nor U4278 (N_4278,In_223,In_482);
and U4279 (N_4279,In_938,In_309);
nor U4280 (N_4280,In_248,In_832);
xor U4281 (N_4281,In_432,In_507);
and U4282 (N_4282,In_428,In_542);
xnor U4283 (N_4283,In_134,In_817);
nor U4284 (N_4284,In_592,In_660);
nand U4285 (N_4285,In_786,In_535);
or U4286 (N_4286,In_622,In_575);
xnor U4287 (N_4287,In_741,In_229);
nand U4288 (N_4288,In_913,In_741);
nor U4289 (N_4289,In_306,In_823);
xor U4290 (N_4290,In_618,In_823);
nand U4291 (N_4291,In_525,In_762);
or U4292 (N_4292,In_597,In_128);
and U4293 (N_4293,In_53,In_806);
and U4294 (N_4294,In_983,In_487);
and U4295 (N_4295,In_749,In_152);
nor U4296 (N_4296,In_380,In_235);
nor U4297 (N_4297,In_468,In_856);
xnor U4298 (N_4298,In_883,In_648);
or U4299 (N_4299,In_501,In_974);
nand U4300 (N_4300,In_452,In_188);
or U4301 (N_4301,In_122,In_99);
nand U4302 (N_4302,In_665,In_608);
or U4303 (N_4303,In_504,In_613);
nand U4304 (N_4304,In_939,In_741);
xor U4305 (N_4305,In_646,In_199);
nand U4306 (N_4306,In_937,In_56);
and U4307 (N_4307,In_642,In_601);
or U4308 (N_4308,In_242,In_695);
nand U4309 (N_4309,In_47,In_719);
and U4310 (N_4310,In_917,In_337);
nor U4311 (N_4311,In_561,In_816);
nand U4312 (N_4312,In_366,In_720);
nand U4313 (N_4313,In_533,In_734);
nand U4314 (N_4314,In_619,In_587);
nor U4315 (N_4315,In_851,In_271);
or U4316 (N_4316,In_344,In_418);
nor U4317 (N_4317,In_95,In_611);
and U4318 (N_4318,In_329,In_215);
xor U4319 (N_4319,In_569,In_485);
nand U4320 (N_4320,In_369,In_68);
or U4321 (N_4321,In_63,In_787);
nor U4322 (N_4322,In_733,In_75);
nor U4323 (N_4323,In_697,In_448);
xnor U4324 (N_4324,In_431,In_12);
and U4325 (N_4325,In_759,In_515);
xor U4326 (N_4326,In_187,In_953);
nand U4327 (N_4327,In_808,In_594);
and U4328 (N_4328,In_309,In_583);
nor U4329 (N_4329,In_181,In_872);
xnor U4330 (N_4330,In_923,In_869);
and U4331 (N_4331,In_221,In_444);
and U4332 (N_4332,In_341,In_895);
nor U4333 (N_4333,In_735,In_695);
nor U4334 (N_4334,In_689,In_515);
nor U4335 (N_4335,In_831,In_764);
or U4336 (N_4336,In_455,In_496);
xnor U4337 (N_4337,In_402,In_369);
and U4338 (N_4338,In_728,In_314);
nor U4339 (N_4339,In_973,In_832);
and U4340 (N_4340,In_637,In_816);
and U4341 (N_4341,In_8,In_921);
nor U4342 (N_4342,In_427,In_662);
nand U4343 (N_4343,In_403,In_249);
nor U4344 (N_4344,In_746,In_552);
xnor U4345 (N_4345,In_474,In_928);
and U4346 (N_4346,In_273,In_210);
xor U4347 (N_4347,In_468,In_220);
or U4348 (N_4348,In_197,In_865);
or U4349 (N_4349,In_572,In_380);
nand U4350 (N_4350,In_514,In_386);
xor U4351 (N_4351,In_949,In_300);
xor U4352 (N_4352,In_691,In_518);
and U4353 (N_4353,In_946,In_626);
or U4354 (N_4354,In_731,In_196);
and U4355 (N_4355,In_505,In_688);
nand U4356 (N_4356,In_140,In_886);
nor U4357 (N_4357,In_435,In_874);
nor U4358 (N_4358,In_874,In_595);
or U4359 (N_4359,In_184,In_751);
and U4360 (N_4360,In_969,In_760);
xor U4361 (N_4361,In_56,In_958);
nand U4362 (N_4362,In_32,In_947);
or U4363 (N_4363,In_159,In_137);
xnor U4364 (N_4364,In_804,In_223);
xnor U4365 (N_4365,In_365,In_354);
nor U4366 (N_4366,In_425,In_852);
nand U4367 (N_4367,In_798,In_106);
or U4368 (N_4368,In_997,In_262);
nand U4369 (N_4369,In_238,In_686);
nand U4370 (N_4370,In_71,In_755);
or U4371 (N_4371,In_44,In_443);
nor U4372 (N_4372,In_624,In_619);
xnor U4373 (N_4373,In_447,In_476);
and U4374 (N_4374,In_937,In_922);
nor U4375 (N_4375,In_567,In_706);
and U4376 (N_4376,In_223,In_787);
nor U4377 (N_4377,In_177,In_847);
and U4378 (N_4378,In_161,In_147);
xnor U4379 (N_4379,In_760,In_385);
xor U4380 (N_4380,In_543,In_3);
and U4381 (N_4381,In_837,In_257);
or U4382 (N_4382,In_912,In_668);
nand U4383 (N_4383,In_102,In_870);
nand U4384 (N_4384,In_245,In_234);
xor U4385 (N_4385,In_666,In_670);
or U4386 (N_4386,In_942,In_647);
nor U4387 (N_4387,In_140,In_82);
nand U4388 (N_4388,In_67,In_506);
and U4389 (N_4389,In_135,In_872);
or U4390 (N_4390,In_724,In_255);
or U4391 (N_4391,In_488,In_849);
and U4392 (N_4392,In_900,In_628);
nor U4393 (N_4393,In_713,In_493);
nor U4394 (N_4394,In_157,In_353);
nand U4395 (N_4395,In_891,In_541);
xor U4396 (N_4396,In_662,In_177);
xnor U4397 (N_4397,In_675,In_647);
nor U4398 (N_4398,In_447,In_546);
xor U4399 (N_4399,In_609,In_210);
or U4400 (N_4400,In_645,In_464);
nand U4401 (N_4401,In_238,In_433);
and U4402 (N_4402,In_331,In_987);
and U4403 (N_4403,In_777,In_931);
nand U4404 (N_4404,In_27,In_211);
or U4405 (N_4405,In_69,In_895);
nand U4406 (N_4406,In_452,In_247);
nand U4407 (N_4407,In_906,In_186);
nand U4408 (N_4408,In_285,In_276);
nand U4409 (N_4409,In_144,In_807);
xor U4410 (N_4410,In_210,In_749);
xor U4411 (N_4411,In_658,In_826);
and U4412 (N_4412,In_51,In_268);
nand U4413 (N_4413,In_320,In_170);
and U4414 (N_4414,In_868,In_89);
nand U4415 (N_4415,In_35,In_476);
nand U4416 (N_4416,In_786,In_926);
nand U4417 (N_4417,In_976,In_196);
and U4418 (N_4418,In_225,In_664);
xor U4419 (N_4419,In_209,In_781);
xor U4420 (N_4420,In_277,In_332);
or U4421 (N_4421,In_437,In_62);
xnor U4422 (N_4422,In_510,In_433);
nor U4423 (N_4423,In_914,In_876);
nor U4424 (N_4424,In_636,In_910);
and U4425 (N_4425,In_209,In_725);
xor U4426 (N_4426,In_760,In_412);
and U4427 (N_4427,In_89,In_28);
nor U4428 (N_4428,In_893,In_328);
or U4429 (N_4429,In_210,In_701);
xnor U4430 (N_4430,In_460,In_566);
nor U4431 (N_4431,In_940,In_690);
nor U4432 (N_4432,In_867,In_307);
or U4433 (N_4433,In_90,In_882);
or U4434 (N_4434,In_505,In_339);
nor U4435 (N_4435,In_402,In_25);
or U4436 (N_4436,In_765,In_337);
nand U4437 (N_4437,In_184,In_192);
xor U4438 (N_4438,In_787,In_588);
nor U4439 (N_4439,In_721,In_935);
and U4440 (N_4440,In_272,In_647);
nand U4441 (N_4441,In_112,In_597);
xnor U4442 (N_4442,In_3,In_375);
or U4443 (N_4443,In_754,In_283);
nor U4444 (N_4444,In_488,In_682);
xor U4445 (N_4445,In_516,In_748);
or U4446 (N_4446,In_301,In_120);
nand U4447 (N_4447,In_371,In_625);
nand U4448 (N_4448,In_424,In_937);
xnor U4449 (N_4449,In_412,In_447);
nand U4450 (N_4450,In_126,In_842);
nor U4451 (N_4451,In_539,In_591);
and U4452 (N_4452,In_909,In_948);
xnor U4453 (N_4453,In_752,In_531);
or U4454 (N_4454,In_236,In_985);
or U4455 (N_4455,In_316,In_897);
and U4456 (N_4456,In_929,In_747);
nand U4457 (N_4457,In_84,In_302);
xnor U4458 (N_4458,In_701,In_768);
xor U4459 (N_4459,In_922,In_993);
xor U4460 (N_4460,In_937,In_884);
and U4461 (N_4461,In_674,In_983);
and U4462 (N_4462,In_279,In_806);
xor U4463 (N_4463,In_384,In_641);
xnor U4464 (N_4464,In_436,In_324);
and U4465 (N_4465,In_845,In_641);
or U4466 (N_4466,In_426,In_54);
xnor U4467 (N_4467,In_132,In_284);
nand U4468 (N_4468,In_671,In_565);
nor U4469 (N_4469,In_640,In_555);
xor U4470 (N_4470,In_88,In_895);
or U4471 (N_4471,In_373,In_571);
xnor U4472 (N_4472,In_773,In_94);
and U4473 (N_4473,In_173,In_493);
and U4474 (N_4474,In_698,In_566);
nand U4475 (N_4475,In_577,In_332);
nor U4476 (N_4476,In_469,In_19);
or U4477 (N_4477,In_315,In_773);
or U4478 (N_4478,In_278,In_945);
nor U4479 (N_4479,In_124,In_835);
xnor U4480 (N_4480,In_704,In_153);
and U4481 (N_4481,In_41,In_754);
xnor U4482 (N_4482,In_271,In_436);
or U4483 (N_4483,In_542,In_116);
xnor U4484 (N_4484,In_686,In_145);
nor U4485 (N_4485,In_753,In_501);
xnor U4486 (N_4486,In_591,In_70);
and U4487 (N_4487,In_711,In_273);
xnor U4488 (N_4488,In_42,In_226);
or U4489 (N_4489,In_609,In_697);
or U4490 (N_4490,In_49,In_319);
and U4491 (N_4491,In_125,In_703);
or U4492 (N_4492,In_342,In_419);
and U4493 (N_4493,In_123,In_134);
or U4494 (N_4494,In_408,In_908);
xnor U4495 (N_4495,In_707,In_552);
and U4496 (N_4496,In_769,In_939);
nand U4497 (N_4497,In_443,In_392);
or U4498 (N_4498,In_574,In_330);
nand U4499 (N_4499,In_596,In_909);
xnor U4500 (N_4500,In_410,In_517);
nand U4501 (N_4501,In_721,In_56);
nor U4502 (N_4502,In_446,In_400);
or U4503 (N_4503,In_487,In_601);
nor U4504 (N_4504,In_7,In_634);
xor U4505 (N_4505,In_65,In_456);
nand U4506 (N_4506,In_640,In_196);
xnor U4507 (N_4507,In_616,In_450);
and U4508 (N_4508,In_640,In_997);
xnor U4509 (N_4509,In_685,In_411);
nand U4510 (N_4510,In_969,In_108);
nand U4511 (N_4511,In_739,In_607);
nor U4512 (N_4512,In_841,In_777);
nor U4513 (N_4513,In_620,In_557);
nand U4514 (N_4514,In_848,In_670);
or U4515 (N_4515,In_713,In_863);
nand U4516 (N_4516,In_880,In_202);
and U4517 (N_4517,In_485,In_152);
nor U4518 (N_4518,In_556,In_725);
xor U4519 (N_4519,In_663,In_633);
or U4520 (N_4520,In_225,In_140);
xnor U4521 (N_4521,In_749,In_720);
and U4522 (N_4522,In_258,In_934);
or U4523 (N_4523,In_143,In_618);
nand U4524 (N_4524,In_218,In_132);
and U4525 (N_4525,In_139,In_402);
nand U4526 (N_4526,In_865,In_827);
nor U4527 (N_4527,In_146,In_613);
nand U4528 (N_4528,In_998,In_933);
xor U4529 (N_4529,In_510,In_937);
nand U4530 (N_4530,In_419,In_583);
xor U4531 (N_4531,In_754,In_619);
xor U4532 (N_4532,In_853,In_745);
nor U4533 (N_4533,In_118,In_552);
or U4534 (N_4534,In_493,In_746);
nand U4535 (N_4535,In_168,In_487);
nand U4536 (N_4536,In_576,In_108);
xnor U4537 (N_4537,In_958,In_737);
and U4538 (N_4538,In_13,In_505);
nor U4539 (N_4539,In_640,In_119);
and U4540 (N_4540,In_542,In_440);
and U4541 (N_4541,In_438,In_505);
and U4542 (N_4542,In_746,In_902);
and U4543 (N_4543,In_780,In_923);
xor U4544 (N_4544,In_498,In_324);
and U4545 (N_4545,In_298,In_943);
xnor U4546 (N_4546,In_249,In_474);
xnor U4547 (N_4547,In_507,In_176);
and U4548 (N_4548,In_125,In_79);
xor U4549 (N_4549,In_866,In_855);
or U4550 (N_4550,In_468,In_195);
nor U4551 (N_4551,In_388,In_1);
nor U4552 (N_4552,In_557,In_51);
nor U4553 (N_4553,In_116,In_643);
nand U4554 (N_4554,In_212,In_127);
or U4555 (N_4555,In_645,In_493);
or U4556 (N_4556,In_633,In_826);
nor U4557 (N_4557,In_505,In_140);
xnor U4558 (N_4558,In_945,In_750);
or U4559 (N_4559,In_907,In_563);
and U4560 (N_4560,In_713,In_394);
or U4561 (N_4561,In_894,In_482);
and U4562 (N_4562,In_860,In_864);
nand U4563 (N_4563,In_682,In_523);
xor U4564 (N_4564,In_738,In_207);
xor U4565 (N_4565,In_839,In_511);
nor U4566 (N_4566,In_802,In_381);
and U4567 (N_4567,In_471,In_34);
or U4568 (N_4568,In_19,In_635);
xor U4569 (N_4569,In_962,In_959);
nor U4570 (N_4570,In_474,In_478);
or U4571 (N_4571,In_662,In_782);
nand U4572 (N_4572,In_52,In_148);
xnor U4573 (N_4573,In_23,In_152);
nand U4574 (N_4574,In_401,In_456);
nor U4575 (N_4575,In_46,In_184);
or U4576 (N_4576,In_665,In_658);
nor U4577 (N_4577,In_414,In_819);
xnor U4578 (N_4578,In_745,In_506);
nor U4579 (N_4579,In_587,In_255);
xnor U4580 (N_4580,In_494,In_263);
nor U4581 (N_4581,In_292,In_609);
xnor U4582 (N_4582,In_30,In_872);
and U4583 (N_4583,In_114,In_200);
or U4584 (N_4584,In_669,In_766);
xnor U4585 (N_4585,In_919,In_720);
or U4586 (N_4586,In_498,In_600);
and U4587 (N_4587,In_991,In_433);
and U4588 (N_4588,In_495,In_276);
nor U4589 (N_4589,In_113,In_791);
xnor U4590 (N_4590,In_996,In_247);
or U4591 (N_4591,In_49,In_475);
nor U4592 (N_4592,In_935,In_20);
nor U4593 (N_4593,In_933,In_272);
or U4594 (N_4594,In_163,In_825);
or U4595 (N_4595,In_544,In_116);
nor U4596 (N_4596,In_374,In_138);
xor U4597 (N_4597,In_265,In_533);
nor U4598 (N_4598,In_217,In_528);
nand U4599 (N_4599,In_712,In_931);
nand U4600 (N_4600,In_432,In_611);
or U4601 (N_4601,In_671,In_383);
nand U4602 (N_4602,In_619,In_980);
and U4603 (N_4603,In_348,In_691);
xor U4604 (N_4604,In_134,In_698);
and U4605 (N_4605,In_434,In_534);
nor U4606 (N_4606,In_399,In_594);
nor U4607 (N_4607,In_735,In_499);
and U4608 (N_4608,In_223,In_748);
nor U4609 (N_4609,In_522,In_860);
nand U4610 (N_4610,In_343,In_639);
nor U4611 (N_4611,In_130,In_806);
nand U4612 (N_4612,In_95,In_588);
xnor U4613 (N_4613,In_86,In_653);
nor U4614 (N_4614,In_766,In_255);
or U4615 (N_4615,In_958,In_784);
or U4616 (N_4616,In_787,In_492);
xnor U4617 (N_4617,In_473,In_792);
or U4618 (N_4618,In_112,In_920);
and U4619 (N_4619,In_270,In_87);
or U4620 (N_4620,In_758,In_165);
or U4621 (N_4621,In_827,In_163);
xor U4622 (N_4622,In_559,In_491);
nand U4623 (N_4623,In_94,In_958);
nor U4624 (N_4624,In_618,In_76);
or U4625 (N_4625,In_929,In_640);
xor U4626 (N_4626,In_603,In_922);
nor U4627 (N_4627,In_479,In_664);
xnor U4628 (N_4628,In_196,In_774);
nor U4629 (N_4629,In_339,In_787);
or U4630 (N_4630,In_889,In_734);
and U4631 (N_4631,In_166,In_723);
nand U4632 (N_4632,In_512,In_945);
xor U4633 (N_4633,In_312,In_628);
and U4634 (N_4634,In_827,In_105);
or U4635 (N_4635,In_596,In_269);
and U4636 (N_4636,In_762,In_569);
or U4637 (N_4637,In_544,In_57);
nor U4638 (N_4638,In_124,In_447);
and U4639 (N_4639,In_885,In_670);
and U4640 (N_4640,In_352,In_113);
nand U4641 (N_4641,In_527,In_67);
xnor U4642 (N_4642,In_755,In_944);
or U4643 (N_4643,In_446,In_473);
xnor U4644 (N_4644,In_299,In_512);
nand U4645 (N_4645,In_759,In_247);
or U4646 (N_4646,In_335,In_527);
nor U4647 (N_4647,In_567,In_804);
xor U4648 (N_4648,In_252,In_171);
and U4649 (N_4649,In_294,In_950);
and U4650 (N_4650,In_709,In_845);
xnor U4651 (N_4651,In_212,In_919);
and U4652 (N_4652,In_426,In_995);
and U4653 (N_4653,In_307,In_240);
nor U4654 (N_4654,In_750,In_261);
nand U4655 (N_4655,In_460,In_879);
and U4656 (N_4656,In_705,In_520);
nor U4657 (N_4657,In_978,In_556);
and U4658 (N_4658,In_268,In_1);
or U4659 (N_4659,In_191,In_72);
and U4660 (N_4660,In_420,In_198);
or U4661 (N_4661,In_846,In_245);
or U4662 (N_4662,In_616,In_679);
nand U4663 (N_4663,In_665,In_392);
xor U4664 (N_4664,In_264,In_327);
and U4665 (N_4665,In_945,In_971);
or U4666 (N_4666,In_865,In_952);
nand U4667 (N_4667,In_815,In_593);
nand U4668 (N_4668,In_673,In_133);
xor U4669 (N_4669,In_637,In_246);
xnor U4670 (N_4670,In_783,In_502);
or U4671 (N_4671,In_447,In_608);
nor U4672 (N_4672,In_324,In_162);
nor U4673 (N_4673,In_657,In_747);
or U4674 (N_4674,In_462,In_23);
xnor U4675 (N_4675,In_387,In_236);
and U4676 (N_4676,In_200,In_777);
nand U4677 (N_4677,In_376,In_927);
or U4678 (N_4678,In_286,In_785);
nor U4679 (N_4679,In_629,In_527);
nand U4680 (N_4680,In_43,In_695);
xnor U4681 (N_4681,In_638,In_989);
or U4682 (N_4682,In_743,In_28);
or U4683 (N_4683,In_782,In_363);
and U4684 (N_4684,In_894,In_265);
nor U4685 (N_4685,In_565,In_815);
xnor U4686 (N_4686,In_845,In_245);
and U4687 (N_4687,In_323,In_354);
or U4688 (N_4688,In_146,In_181);
nand U4689 (N_4689,In_946,In_866);
or U4690 (N_4690,In_909,In_710);
nor U4691 (N_4691,In_807,In_58);
nand U4692 (N_4692,In_408,In_819);
xor U4693 (N_4693,In_417,In_364);
xnor U4694 (N_4694,In_711,In_394);
nor U4695 (N_4695,In_438,In_307);
nand U4696 (N_4696,In_598,In_146);
or U4697 (N_4697,In_902,In_284);
or U4698 (N_4698,In_562,In_124);
xor U4699 (N_4699,In_809,In_374);
and U4700 (N_4700,In_580,In_773);
nor U4701 (N_4701,In_363,In_43);
nand U4702 (N_4702,In_444,In_864);
or U4703 (N_4703,In_450,In_751);
or U4704 (N_4704,In_465,In_214);
xnor U4705 (N_4705,In_274,In_579);
nor U4706 (N_4706,In_914,In_570);
or U4707 (N_4707,In_858,In_607);
and U4708 (N_4708,In_349,In_355);
nor U4709 (N_4709,In_719,In_759);
nand U4710 (N_4710,In_171,In_594);
nor U4711 (N_4711,In_29,In_79);
or U4712 (N_4712,In_296,In_486);
or U4713 (N_4713,In_244,In_769);
nor U4714 (N_4714,In_920,In_16);
xnor U4715 (N_4715,In_600,In_934);
nand U4716 (N_4716,In_74,In_28);
nor U4717 (N_4717,In_171,In_492);
nand U4718 (N_4718,In_795,In_256);
or U4719 (N_4719,In_731,In_198);
nand U4720 (N_4720,In_766,In_295);
nand U4721 (N_4721,In_713,In_837);
and U4722 (N_4722,In_397,In_222);
xor U4723 (N_4723,In_829,In_545);
xor U4724 (N_4724,In_7,In_965);
and U4725 (N_4725,In_332,In_595);
nor U4726 (N_4726,In_123,In_404);
nor U4727 (N_4727,In_522,In_667);
and U4728 (N_4728,In_432,In_723);
nor U4729 (N_4729,In_519,In_719);
and U4730 (N_4730,In_850,In_891);
or U4731 (N_4731,In_685,In_428);
nor U4732 (N_4732,In_537,In_322);
nand U4733 (N_4733,In_735,In_751);
nor U4734 (N_4734,In_624,In_356);
and U4735 (N_4735,In_290,In_656);
xnor U4736 (N_4736,In_390,In_158);
xnor U4737 (N_4737,In_433,In_183);
xnor U4738 (N_4738,In_465,In_92);
nor U4739 (N_4739,In_233,In_65);
xnor U4740 (N_4740,In_269,In_2);
xnor U4741 (N_4741,In_221,In_440);
xor U4742 (N_4742,In_859,In_972);
nor U4743 (N_4743,In_617,In_456);
or U4744 (N_4744,In_241,In_598);
xor U4745 (N_4745,In_742,In_705);
xnor U4746 (N_4746,In_859,In_44);
xor U4747 (N_4747,In_129,In_30);
or U4748 (N_4748,In_424,In_20);
xnor U4749 (N_4749,In_119,In_579);
xnor U4750 (N_4750,In_671,In_89);
or U4751 (N_4751,In_638,In_313);
and U4752 (N_4752,In_822,In_548);
xnor U4753 (N_4753,In_512,In_946);
or U4754 (N_4754,In_923,In_993);
or U4755 (N_4755,In_287,In_247);
or U4756 (N_4756,In_28,In_885);
xor U4757 (N_4757,In_369,In_303);
nor U4758 (N_4758,In_137,In_988);
or U4759 (N_4759,In_807,In_953);
and U4760 (N_4760,In_354,In_531);
and U4761 (N_4761,In_549,In_75);
nor U4762 (N_4762,In_45,In_110);
and U4763 (N_4763,In_661,In_369);
nand U4764 (N_4764,In_306,In_649);
or U4765 (N_4765,In_264,In_413);
and U4766 (N_4766,In_917,In_978);
or U4767 (N_4767,In_824,In_594);
or U4768 (N_4768,In_151,In_322);
nor U4769 (N_4769,In_277,In_870);
xor U4770 (N_4770,In_39,In_391);
nor U4771 (N_4771,In_683,In_636);
or U4772 (N_4772,In_360,In_94);
or U4773 (N_4773,In_735,In_25);
xor U4774 (N_4774,In_275,In_587);
nand U4775 (N_4775,In_925,In_595);
xor U4776 (N_4776,In_40,In_297);
xnor U4777 (N_4777,In_961,In_375);
nand U4778 (N_4778,In_852,In_352);
or U4779 (N_4779,In_266,In_620);
nor U4780 (N_4780,In_181,In_174);
or U4781 (N_4781,In_859,In_620);
nand U4782 (N_4782,In_364,In_119);
and U4783 (N_4783,In_618,In_308);
xnor U4784 (N_4784,In_397,In_800);
nor U4785 (N_4785,In_265,In_951);
nand U4786 (N_4786,In_472,In_670);
nor U4787 (N_4787,In_591,In_189);
xor U4788 (N_4788,In_175,In_424);
and U4789 (N_4789,In_23,In_574);
and U4790 (N_4790,In_809,In_17);
or U4791 (N_4791,In_153,In_425);
and U4792 (N_4792,In_594,In_168);
or U4793 (N_4793,In_750,In_687);
nor U4794 (N_4794,In_797,In_854);
nor U4795 (N_4795,In_667,In_764);
and U4796 (N_4796,In_727,In_380);
xor U4797 (N_4797,In_744,In_797);
nand U4798 (N_4798,In_982,In_676);
and U4799 (N_4799,In_139,In_287);
and U4800 (N_4800,In_596,In_441);
nand U4801 (N_4801,In_829,In_200);
xnor U4802 (N_4802,In_411,In_763);
or U4803 (N_4803,In_727,In_30);
xor U4804 (N_4804,In_543,In_670);
and U4805 (N_4805,In_859,In_390);
nor U4806 (N_4806,In_10,In_146);
nor U4807 (N_4807,In_60,In_597);
nand U4808 (N_4808,In_802,In_304);
xor U4809 (N_4809,In_838,In_237);
xnor U4810 (N_4810,In_514,In_627);
or U4811 (N_4811,In_525,In_618);
nor U4812 (N_4812,In_984,In_556);
nor U4813 (N_4813,In_614,In_618);
nand U4814 (N_4814,In_160,In_972);
nand U4815 (N_4815,In_610,In_726);
xor U4816 (N_4816,In_239,In_95);
nand U4817 (N_4817,In_779,In_232);
nand U4818 (N_4818,In_442,In_950);
nor U4819 (N_4819,In_834,In_495);
nor U4820 (N_4820,In_937,In_532);
nor U4821 (N_4821,In_216,In_844);
nand U4822 (N_4822,In_388,In_715);
or U4823 (N_4823,In_298,In_512);
xor U4824 (N_4824,In_562,In_19);
or U4825 (N_4825,In_571,In_663);
nand U4826 (N_4826,In_235,In_105);
xor U4827 (N_4827,In_563,In_906);
or U4828 (N_4828,In_772,In_92);
or U4829 (N_4829,In_876,In_12);
nor U4830 (N_4830,In_953,In_328);
xnor U4831 (N_4831,In_93,In_241);
nor U4832 (N_4832,In_214,In_722);
nor U4833 (N_4833,In_563,In_754);
xor U4834 (N_4834,In_770,In_57);
nand U4835 (N_4835,In_148,In_215);
or U4836 (N_4836,In_246,In_113);
and U4837 (N_4837,In_449,In_501);
xor U4838 (N_4838,In_46,In_40);
and U4839 (N_4839,In_168,In_877);
nand U4840 (N_4840,In_113,In_228);
nand U4841 (N_4841,In_329,In_471);
or U4842 (N_4842,In_531,In_16);
and U4843 (N_4843,In_768,In_423);
nand U4844 (N_4844,In_702,In_642);
nand U4845 (N_4845,In_298,In_36);
nor U4846 (N_4846,In_699,In_660);
nor U4847 (N_4847,In_947,In_524);
nor U4848 (N_4848,In_69,In_280);
or U4849 (N_4849,In_656,In_218);
xor U4850 (N_4850,In_649,In_990);
xnor U4851 (N_4851,In_592,In_23);
nand U4852 (N_4852,In_452,In_724);
nand U4853 (N_4853,In_283,In_335);
xor U4854 (N_4854,In_737,In_833);
or U4855 (N_4855,In_288,In_33);
or U4856 (N_4856,In_276,In_114);
or U4857 (N_4857,In_14,In_446);
nand U4858 (N_4858,In_401,In_846);
nor U4859 (N_4859,In_202,In_932);
nand U4860 (N_4860,In_501,In_413);
xor U4861 (N_4861,In_980,In_349);
nor U4862 (N_4862,In_374,In_259);
xnor U4863 (N_4863,In_874,In_187);
nor U4864 (N_4864,In_951,In_120);
xor U4865 (N_4865,In_844,In_859);
or U4866 (N_4866,In_30,In_889);
xor U4867 (N_4867,In_141,In_85);
nand U4868 (N_4868,In_446,In_865);
or U4869 (N_4869,In_433,In_585);
and U4870 (N_4870,In_509,In_332);
nand U4871 (N_4871,In_962,In_73);
nor U4872 (N_4872,In_898,In_113);
nand U4873 (N_4873,In_380,In_654);
nor U4874 (N_4874,In_952,In_460);
and U4875 (N_4875,In_742,In_102);
nor U4876 (N_4876,In_117,In_668);
nand U4877 (N_4877,In_268,In_791);
nand U4878 (N_4878,In_895,In_558);
xor U4879 (N_4879,In_475,In_873);
nand U4880 (N_4880,In_801,In_439);
nor U4881 (N_4881,In_863,In_282);
nor U4882 (N_4882,In_535,In_445);
and U4883 (N_4883,In_584,In_444);
nand U4884 (N_4884,In_362,In_312);
or U4885 (N_4885,In_958,In_669);
and U4886 (N_4886,In_113,In_9);
nand U4887 (N_4887,In_873,In_62);
and U4888 (N_4888,In_809,In_411);
nor U4889 (N_4889,In_331,In_887);
nand U4890 (N_4890,In_118,In_833);
nor U4891 (N_4891,In_621,In_455);
nor U4892 (N_4892,In_343,In_240);
or U4893 (N_4893,In_373,In_749);
xnor U4894 (N_4894,In_420,In_115);
or U4895 (N_4895,In_675,In_984);
or U4896 (N_4896,In_298,In_257);
nor U4897 (N_4897,In_769,In_626);
nor U4898 (N_4898,In_614,In_959);
xor U4899 (N_4899,In_587,In_101);
and U4900 (N_4900,In_817,In_759);
and U4901 (N_4901,In_834,In_153);
nor U4902 (N_4902,In_367,In_359);
xor U4903 (N_4903,In_26,In_565);
and U4904 (N_4904,In_469,In_410);
xnor U4905 (N_4905,In_261,In_932);
xor U4906 (N_4906,In_554,In_651);
nand U4907 (N_4907,In_382,In_211);
and U4908 (N_4908,In_489,In_460);
nand U4909 (N_4909,In_543,In_641);
and U4910 (N_4910,In_999,In_715);
and U4911 (N_4911,In_643,In_925);
nor U4912 (N_4912,In_195,In_725);
and U4913 (N_4913,In_821,In_84);
and U4914 (N_4914,In_568,In_360);
nand U4915 (N_4915,In_759,In_438);
nor U4916 (N_4916,In_807,In_994);
and U4917 (N_4917,In_662,In_145);
nand U4918 (N_4918,In_534,In_254);
nand U4919 (N_4919,In_340,In_331);
nor U4920 (N_4920,In_905,In_246);
and U4921 (N_4921,In_514,In_78);
and U4922 (N_4922,In_497,In_857);
or U4923 (N_4923,In_248,In_231);
and U4924 (N_4924,In_267,In_268);
xor U4925 (N_4925,In_590,In_295);
nor U4926 (N_4926,In_504,In_810);
or U4927 (N_4927,In_601,In_126);
and U4928 (N_4928,In_37,In_127);
nand U4929 (N_4929,In_768,In_567);
xnor U4930 (N_4930,In_590,In_790);
nor U4931 (N_4931,In_951,In_443);
nor U4932 (N_4932,In_241,In_765);
or U4933 (N_4933,In_965,In_58);
xnor U4934 (N_4934,In_179,In_6);
nor U4935 (N_4935,In_517,In_332);
nand U4936 (N_4936,In_852,In_389);
nor U4937 (N_4937,In_587,In_580);
nand U4938 (N_4938,In_256,In_790);
and U4939 (N_4939,In_550,In_754);
and U4940 (N_4940,In_454,In_895);
nand U4941 (N_4941,In_959,In_835);
and U4942 (N_4942,In_396,In_615);
or U4943 (N_4943,In_195,In_602);
nand U4944 (N_4944,In_869,In_750);
and U4945 (N_4945,In_615,In_622);
nand U4946 (N_4946,In_948,In_327);
nor U4947 (N_4947,In_656,In_306);
xnor U4948 (N_4948,In_643,In_468);
nand U4949 (N_4949,In_756,In_456);
nand U4950 (N_4950,In_438,In_388);
and U4951 (N_4951,In_204,In_350);
and U4952 (N_4952,In_806,In_917);
nor U4953 (N_4953,In_664,In_376);
nand U4954 (N_4954,In_5,In_705);
or U4955 (N_4955,In_408,In_891);
xor U4956 (N_4956,In_965,In_106);
nor U4957 (N_4957,In_834,In_465);
nand U4958 (N_4958,In_978,In_673);
and U4959 (N_4959,In_747,In_752);
xor U4960 (N_4960,In_907,In_842);
xnor U4961 (N_4961,In_822,In_362);
nand U4962 (N_4962,In_491,In_352);
nor U4963 (N_4963,In_358,In_421);
xnor U4964 (N_4964,In_592,In_238);
nand U4965 (N_4965,In_923,In_196);
and U4966 (N_4966,In_62,In_700);
xnor U4967 (N_4967,In_18,In_466);
xor U4968 (N_4968,In_990,In_596);
or U4969 (N_4969,In_209,In_810);
or U4970 (N_4970,In_245,In_443);
nand U4971 (N_4971,In_490,In_415);
xnor U4972 (N_4972,In_55,In_861);
or U4973 (N_4973,In_61,In_561);
and U4974 (N_4974,In_26,In_437);
nor U4975 (N_4975,In_719,In_369);
nor U4976 (N_4976,In_200,In_540);
nand U4977 (N_4977,In_413,In_55);
or U4978 (N_4978,In_365,In_290);
nand U4979 (N_4979,In_743,In_605);
and U4980 (N_4980,In_437,In_41);
and U4981 (N_4981,In_194,In_446);
nor U4982 (N_4982,In_900,In_840);
nor U4983 (N_4983,In_520,In_119);
or U4984 (N_4984,In_927,In_610);
xnor U4985 (N_4985,In_698,In_955);
and U4986 (N_4986,In_169,In_250);
xnor U4987 (N_4987,In_775,In_895);
or U4988 (N_4988,In_61,In_507);
and U4989 (N_4989,In_831,In_955);
and U4990 (N_4990,In_9,In_612);
or U4991 (N_4991,In_852,In_154);
and U4992 (N_4992,In_793,In_14);
or U4993 (N_4993,In_638,In_579);
xor U4994 (N_4994,In_355,In_645);
and U4995 (N_4995,In_534,In_880);
and U4996 (N_4996,In_290,In_326);
and U4997 (N_4997,In_136,In_2);
and U4998 (N_4998,In_321,In_479);
or U4999 (N_4999,In_21,In_996);
nand U5000 (N_5000,N_1162,N_4706);
nand U5001 (N_5001,N_3376,N_1545);
nor U5002 (N_5002,N_1876,N_364);
and U5003 (N_5003,N_2199,N_85);
nand U5004 (N_5004,N_2223,N_3770);
and U5005 (N_5005,N_100,N_3517);
or U5006 (N_5006,N_2132,N_2275);
nand U5007 (N_5007,N_2078,N_2599);
and U5008 (N_5008,N_1078,N_1561);
nand U5009 (N_5009,N_4636,N_2147);
nand U5010 (N_5010,N_3,N_3858);
xnor U5011 (N_5011,N_2339,N_2084);
or U5012 (N_5012,N_3504,N_2806);
xnor U5013 (N_5013,N_4650,N_4056);
nor U5014 (N_5014,N_1409,N_353);
nand U5015 (N_5015,N_5,N_3387);
xnor U5016 (N_5016,N_3385,N_4285);
nand U5017 (N_5017,N_2650,N_4145);
nand U5018 (N_5018,N_4690,N_891);
nor U5019 (N_5019,N_3865,N_3221);
or U5020 (N_5020,N_4184,N_302);
xnor U5021 (N_5021,N_2971,N_649);
or U5022 (N_5022,N_1836,N_1222);
xnor U5023 (N_5023,N_633,N_1248);
xor U5024 (N_5024,N_3163,N_19);
nand U5025 (N_5025,N_4950,N_177);
and U5026 (N_5026,N_391,N_483);
xor U5027 (N_5027,N_3233,N_2855);
xor U5028 (N_5028,N_3894,N_624);
nand U5029 (N_5029,N_66,N_2757);
and U5030 (N_5030,N_308,N_2557);
nor U5031 (N_5031,N_966,N_716);
xnor U5032 (N_5032,N_3343,N_3723);
nor U5033 (N_5033,N_2949,N_407);
or U5034 (N_5034,N_3505,N_1103);
or U5035 (N_5035,N_3767,N_1124);
and U5036 (N_5036,N_3993,N_775);
xnor U5037 (N_5037,N_763,N_3256);
nand U5038 (N_5038,N_2658,N_882);
and U5039 (N_5039,N_176,N_2741);
or U5040 (N_5040,N_1421,N_3487);
and U5041 (N_5041,N_1475,N_414);
nand U5042 (N_5042,N_4613,N_4853);
or U5043 (N_5043,N_2433,N_693);
or U5044 (N_5044,N_2591,N_262);
xnor U5045 (N_5045,N_2884,N_1471);
nand U5046 (N_5046,N_637,N_3829);
nand U5047 (N_5047,N_1331,N_895);
nor U5048 (N_5048,N_3615,N_3442);
nor U5049 (N_5049,N_3599,N_1129);
nand U5050 (N_5050,N_546,N_2938);
nand U5051 (N_5051,N_3817,N_2897);
xor U5052 (N_5052,N_460,N_4361);
nand U5053 (N_5053,N_1377,N_1181);
xor U5054 (N_5054,N_4141,N_452);
nor U5055 (N_5055,N_4498,N_1369);
xnor U5056 (N_5056,N_2595,N_4235);
xnor U5057 (N_5057,N_872,N_3077);
nor U5058 (N_5058,N_509,N_3969);
and U5059 (N_5059,N_1108,N_33);
or U5060 (N_5060,N_2887,N_2969);
and U5061 (N_5061,N_588,N_4676);
nor U5062 (N_5062,N_1579,N_3763);
and U5063 (N_5063,N_1688,N_3853);
xnor U5064 (N_5064,N_2919,N_1821);
xnor U5065 (N_5065,N_4604,N_4571);
xnor U5066 (N_5066,N_4120,N_4480);
xnor U5067 (N_5067,N_1073,N_599);
and U5068 (N_5068,N_542,N_4575);
or U5069 (N_5069,N_2612,N_84);
or U5070 (N_5070,N_4257,N_3940);
xnor U5071 (N_5071,N_3590,N_1261);
xor U5072 (N_5072,N_1334,N_3701);
or U5073 (N_5073,N_1598,N_332);
nor U5074 (N_5074,N_754,N_3014);
xnor U5075 (N_5075,N_52,N_3951);
or U5076 (N_5076,N_3887,N_2305);
nor U5077 (N_5077,N_503,N_747);
nand U5078 (N_5078,N_1278,N_4703);
xnor U5079 (N_5079,N_2069,N_4905);
and U5080 (N_5080,N_4482,N_2614);
or U5081 (N_5081,N_2970,N_2226);
and U5082 (N_5082,N_1631,N_185);
and U5083 (N_5083,N_301,N_447);
nand U5084 (N_5084,N_4954,N_160);
or U5085 (N_5085,N_3276,N_3704);
and U5086 (N_5086,N_71,N_4733);
or U5087 (N_5087,N_3353,N_1931);
or U5088 (N_5088,N_1014,N_2169);
xor U5089 (N_5089,N_215,N_2935);
and U5090 (N_5090,N_4149,N_809);
and U5091 (N_5091,N_4555,N_2001);
xnor U5092 (N_5092,N_4956,N_1072);
nand U5093 (N_5093,N_1065,N_2415);
or U5094 (N_5094,N_903,N_4791);
nand U5095 (N_5095,N_2179,N_877);
nor U5096 (N_5096,N_4888,N_749);
nor U5097 (N_5097,N_2460,N_2847);
nor U5098 (N_5098,N_4828,N_1842);
or U5099 (N_5099,N_4046,N_505);
and U5100 (N_5100,N_4383,N_4894);
or U5101 (N_5101,N_717,N_2868);
xor U5102 (N_5102,N_3524,N_4692);
and U5103 (N_5103,N_2209,N_229);
and U5104 (N_5104,N_4583,N_1036);
xor U5105 (N_5105,N_3316,N_3898);
nand U5106 (N_5106,N_4123,N_1163);
nand U5107 (N_5107,N_1667,N_4887);
or U5108 (N_5108,N_516,N_2787);
and U5109 (N_5109,N_3844,N_2455);
nor U5110 (N_5110,N_626,N_3365);
nand U5111 (N_5111,N_3994,N_1279);
or U5112 (N_5112,N_2342,N_441);
nor U5113 (N_5113,N_4458,N_2880);
nor U5114 (N_5114,N_1998,N_2077);
and U5115 (N_5115,N_3296,N_550);
or U5116 (N_5116,N_2941,N_4927);
nor U5117 (N_5117,N_3691,N_2265);
nand U5118 (N_5118,N_1383,N_4724);
nand U5119 (N_5119,N_3210,N_2546);
xor U5120 (N_5120,N_4138,N_3067);
nand U5121 (N_5121,N_3911,N_3248);
nor U5122 (N_5122,N_673,N_2621);
and U5123 (N_5123,N_1634,N_662);
nand U5124 (N_5124,N_2268,N_4713);
and U5125 (N_5125,N_2921,N_4417);
or U5126 (N_5126,N_335,N_4239);
xnor U5127 (N_5127,N_4322,N_3892);
xnor U5128 (N_5128,N_4949,N_73);
and U5129 (N_5129,N_3293,N_2821);
and U5130 (N_5130,N_3058,N_3793);
nand U5131 (N_5131,N_1722,N_2665);
nor U5132 (N_5132,N_2845,N_3432);
nor U5133 (N_5133,N_4646,N_941);
xor U5134 (N_5134,N_405,N_4721);
nand U5135 (N_5135,N_379,N_1288);
xnor U5136 (N_5136,N_1760,N_2501);
xor U5137 (N_5137,N_4944,N_4060);
and U5138 (N_5138,N_2898,N_2058);
nand U5139 (N_5139,N_2710,N_2183);
nor U5140 (N_5140,N_1196,N_1179);
nand U5141 (N_5141,N_2146,N_1643);
xor U5142 (N_5142,N_67,N_1095);
xnor U5143 (N_5143,N_4456,N_2734);
and U5144 (N_5144,N_3882,N_1328);
and U5145 (N_5145,N_756,N_3947);
nand U5146 (N_5146,N_4674,N_1967);
nor U5147 (N_5147,N_777,N_1737);
xnor U5148 (N_5148,N_902,N_2812);
nor U5149 (N_5149,N_2200,N_2271);
nand U5150 (N_5150,N_4883,N_63);
xnor U5151 (N_5151,N_648,N_3870);
or U5152 (N_5152,N_1498,N_3259);
and U5153 (N_5153,N_3565,N_2831);
or U5154 (N_5154,N_1211,N_463);
or U5155 (N_5155,N_2815,N_2135);
xnor U5156 (N_5156,N_471,N_2028);
or U5157 (N_5157,N_1258,N_836);
nor U5158 (N_5158,N_1040,N_4521);
nand U5159 (N_5159,N_4971,N_1712);
or U5160 (N_5160,N_2804,N_3532);
or U5161 (N_5161,N_4275,N_962);
and U5162 (N_5162,N_277,N_4356);
or U5163 (N_5163,N_3946,N_4665);
nor U5164 (N_5164,N_219,N_2598);
and U5165 (N_5165,N_1742,N_4619);
or U5166 (N_5166,N_4207,N_4868);
nor U5167 (N_5167,N_3078,N_803);
xnor U5168 (N_5168,N_3582,N_689);
and U5169 (N_5169,N_597,N_1976);
nor U5170 (N_5170,N_3064,N_1188);
nor U5171 (N_5171,N_3936,N_26);
nand U5172 (N_5172,N_3754,N_1015);
or U5173 (N_5173,N_275,N_831);
and U5174 (N_5174,N_3627,N_3709);
xnor U5175 (N_5175,N_1618,N_4578);
or U5176 (N_5176,N_3978,N_1310);
or U5177 (N_5177,N_1984,N_1002);
and U5178 (N_5178,N_1201,N_1965);
nand U5179 (N_5179,N_1875,N_3018);
and U5180 (N_5180,N_3731,N_3373);
nor U5181 (N_5181,N_3589,N_25);
xor U5182 (N_5182,N_3133,N_4687);
or U5183 (N_5183,N_3162,N_1996);
and U5184 (N_5184,N_2326,N_867);
or U5185 (N_5185,N_1134,N_3099);
nand U5186 (N_5186,N_939,N_2492);
nand U5187 (N_5187,N_2645,N_2860);
and U5188 (N_5188,N_4847,N_745);
nand U5189 (N_5189,N_3366,N_2716);
and U5190 (N_5190,N_2116,N_4109);
and U5191 (N_5191,N_1653,N_4192);
xnor U5192 (N_5192,N_2027,N_3923);
or U5193 (N_5193,N_515,N_2863);
nand U5194 (N_5194,N_2382,N_1100);
nor U5195 (N_5195,N_4427,N_3838);
xor U5196 (N_5196,N_4700,N_4911);
or U5197 (N_5197,N_3242,N_1122);
and U5198 (N_5198,N_3631,N_1297);
nand U5199 (N_5199,N_2561,N_3328);
nand U5200 (N_5200,N_2467,N_2029);
xor U5201 (N_5201,N_4513,N_735);
nor U5202 (N_5202,N_4105,N_3305);
nand U5203 (N_5203,N_4463,N_2745);
xnor U5204 (N_5204,N_3482,N_1657);
nor U5205 (N_5205,N_3108,N_3737);
nand U5206 (N_5206,N_1338,N_548);
or U5207 (N_5207,N_3357,N_3997);
nor U5208 (N_5208,N_2487,N_315);
and U5209 (N_5209,N_761,N_932);
and U5210 (N_5210,N_4741,N_2365);
and U5211 (N_5211,N_2186,N_3840);
and U5212 (N_5212,N_3194,N_1128);
and U5213 (N_5213,N_788,N_3719);
nor U5214 (N_5214,N_684,N_4628);
and U5215 (N_5215,N_3780,N_4076);
and U5216 (N_5216,N_644,N_311);
and U5217 (N_5217,N_3687,N_427);
xor U5218 (N_5218,N_4761,N_2004);
xor U5219 (N_5219,N_3331,N_3681);
xor U5220 (N_5220,N_1479,N_4876);
nand U5221 (N_5221,N_3778,N_1774);
or U5222 (N_5222,N_1928,N_3106);
and U5223 (N_5223,N_1434,N_2024);
and U5224 (N_5224,N_2389,N_2089);
nand U5225 (N_5225,N_3313,N_3744);
nand U5226 (N_5226,N_1048,N_1696);
or U5227 (N_5227,N_778,N_4187);
nor U5228 (N_5228,N_1644,N_1704);
or U5229 (N_5229,N_4852,N_2442);
and U5230 (N_5230,N_2571,N_3121);
xnor U5231 (N_5231,N_4201,N_2222);
nand U5232 (N_5232,N_1028,N_382);
xor U5233 (N_5233,N_3741,N_1846);
and U5234 (N_5234,N_2411,N_1701);
nand U5235 (N_5235,N_2872,N_2021);
and U5236 (N_5236,N_1362,N_3799);
nor U5237 (N_5237,N_2309,N_303);
xnor U5238 (N_5238,N_3231,N_4952);
nand U5239 (N_5239,N_1245,N_1047);
nor U5240 (N_5240,N_729,N_4644);
nor U5241 (N_5241,N_3805,N_1);
xor U5242 (N_5242,N_1880,N_3007);
and U5243 (N_5243,N_4100,N_2177);
nor U5244 (N_5244,N_2870,N_1765);
xor U5245 (N_5245,N_2313,N_3956);
or U5246 (N_5246,N_1894,N_2759);
xor U5247 (N_5247,N_1370,N_196);
and U5248 (N_5248,N_604,N_2376);
nand U5249 (N_5249,N_1425,N_3932);
nand U5250 (N_5250,N_445,N_4842);
nand U5251 (N_5251,N_660,N_2681);
and U5252 (N_5252,N_1464,N_4566);
nand U5253 (N_5253,N_4374,N_3355);
or U5254 (N_5254,N_3608,N_3884);
xor U5255 (N_5255,N_2458,N_1626);
nor U5256 (N_5256,N_2842,N_4923);
or U5257 (N_5257,N_473,N_554);
nand U5258 (N_5258,N_2418,N_1799);
or U5259 (N_5259,N_141,N_4367);
xor U5260 (N_5260,N_2766,N_1625);
or U5261 (N_5261,N_2666,N_2481);
xor U5262 (N_5262,N_4357,N_3957);
and U5263 (N_5263,N_4068,N_1767);
xnor U5264 (N_5264,N_1980,N_4432);
xnor U5265 (N_5265,N_969,N_4772);
nor U5266 (N_5266,N_4892,N_2254);
xor U5267 (N_5267,N_2337,N_4328);
and U5268 (N_5268,N_107,N_2020);
or U5269 (N_5269,N_2422,N_3930);
and U5270 (N_5270,N_1729,N_883);
nor U5271 (N_5271,N_3413,N_4462);
xnor U5272 (N_5272,N_1609,N_2783);
nand U5273 (N_5273,N_4744,N_74);
xor U5274 (N_5274,N_502,N_2674);
xnor U5275 (N_5275,N_2857,N_4005);
nor U5276 (N_5276,N_694,N_96);
or U5277 (N_5277,N_134,N_3772);
xor U5278 (N_5278,N_1136,N_1446);
nand U5279 (N_5279,N_1818,N_3179);
nor U5280 (N_5280,N_2932,N_3555);
nand U5281 (N_5281,N_3502,N_2620);
nor U5282 (N_5282,N_2999,N_3283);
xor U5283 (N_5283,N_1091,N_2216);
xor U5284 (N_5284,N_4603,N_937);
and U5285 (N_5285,N_4580,N_4536);
nor U5286 (N_5286,N_3416,N_3753);
and U5287 (N_5287,N_2359,N_1466);
or U5288 (N_5288,N_2236,N_2565);
nand U5289 (N_5289,N_1178,N_2789);
nand U5290 (N_5290,N_866,N_1357);
nor U5291 (N_5291,N_791,N_2434);
xnor U5292 (N_5292,N_2228,N_1254);
or U5293 (N_5293,N_4034,N_4871);
and U5294 (N_5294,N_142,N_3860);
or U5295 (N_5295,N_171,N_1623);
nand U5296 (N_5296,N_3223,N_3617);
nor U5297 (N_5297,N_2749,N_2370);
xnor U5298 (N_5298,N_1403,N_580);
or U5299 (N_5299,N_704,N_3103);
and U5300 (N_5300,N_2279,N_4595);
nor U5301 (N_5301,N_4360,N_4183);
and U5302 (N_5302,N_1837,N_936);
nand U5303 (N_5303,N_2768,N_3815);
nor U5304 (N_5304,N_77,N_2986);
nor U5305 (N_5305,N_1796,N_2189);
nand U5306 (N_5306,N_3665,N_987);
or U5307 (N_5307,N_2597,N_1336);
or U5308 (N_5308,N_1534,N_3540);
nand U5309 (N_5309,N_3364,N_1067);
nand U5310 (N_5310,N_2841,N_1472);
and U5311 (N_5311,N_1795,N_2539);
or U5312 (N_5312,N_3302,N_4066);
or U5313 (N_5313,N_4838,N_3755);
xor U5314 (N_5314,N_3931,N_1683);
and U5315 (N_5315,N_3751,N_4256);
or U5316 (N_5316,N_4726,N_2774);
xnor U5317 (N_5317,N_2092,N_3303);
and U5318 (N_5318,N_1359,N_1728);
or U5319 (N_5319,N_3588,N_1456);
and U5320 (N_5320,N_2334,N_4786);
nand U5321 (N_5321,N_2231,N_4085);
or U5322 (N_5322,N_3843,N_2730);
nor U5323 (N_5323,N_2157,N_2378);
nor U5324 (N_5324,N_1097,N_1523);
nor U5325 (N_5325,N_166,N_2213);
nor U5326 (N_5326,N_4494,N_3928);
nor U5327 (N_5327,N_1037,N_462);
nand U5328 (N_5328,N_3325,N_1981);
or U5329 (N_5329,N_2979,N_1249);
and U5330 (N_5330,N_1919,N_4775);
nor U5331 (N_5331,N_2130,N_1467);
nor U5332 (N_5332,N_4220,N_4130);
or U5333 (N_5333,N_4258,N_2220);
and U5334 (N_5334,N_1244,N_2520);
or U5335 (N_5335,N_387,N_188);
and U5336 (N_5336,N_4885,N_4897);
xor U5337 (N_5337,N_1524,N_2534);
nor U5338 (N_5338,N_2685,N_4704);
nand U5339 (N_5339,N_538,N_3920);
nor U5340 (N_5340,N_1801,N_4902);
and U5341 (N_5341,N_338,N_3847);
nor U5342 (N_5342,N_1959,N_1542);
nand U5343 (N_5343,N_4439,N_2461);
nor U5344 (N_5344,N_3954,N_3145);
nand U5345 (N_5345,N_2448,N_3604);
nor U5346 (N_5346,N_1085,N_1603);
xnor U5347 (N_5347,N_3960,N_4880);
nor U5348 (N_5348,N_557,N_31);
and U5349 (N_5349,N_1418,N_3086);
xor U5350 (N_5350,N_1106,N_3529);
or U5351 (N_5351,N_4255,N_1590);
or U5352 (N_5352,N_833,N_24);
or U5353 (N_5353,N_2724,N_4379);
xor U5354 (N_5354,N_3310,N_2524);
nand U5355 (N_5355,N_1887,N_3542);
nor U5356 (N_5356,N_804,N_3149);
xnor U5357 (N_5357,N_751,N_880);
and U5358 (N_5358,N_3237,N_3886);
and U5359 (N_5359,N_3630,N_2703);
or U5360 (N_5360,N_4756,N_3094);
nor U5361 (N_5361,N_268,N_173);
nand U5362 (N_5362,N_430,N_1907);
nor U5363 (N_5363,N_1203,N_1373);
nand U5364 (N_5364,N_4754,N_708);
and U5365 (N_5365,N_1544,N_2102);
xor U5366 (N_5366,N_3267,N_3483);
nor U5367 (N_5367,N_625,N_3206);
or U5368 (N_5368,N_4233,N_4858);
or U5369 (N_5369,N_2090,N_3850);
or U5370 (N_5370,N_294,N_3809);
nor U5371 (N_5371,N_4174,N_2413);
xnor U5372 (N_5372,N_1253,N_207);
and U5373 (N_5373,N_1102,N_830);
nor U5374 (N_5374,N_2110,N_3459);
and U5375 (N_5375,N_155,N_1844);
xnor U5376 (N_5376,N_3675,N_1526);
xor U5377 (N_5377,N_2762,N_4631);
and U5378 (N_5378,N_3026,N_3451);
xor U5379 (N_5379,N_4999,N_1404);
xnor U5380 (N_5380,N_591,N_2782);
nand U5381 (N_5381,N_1933,N_4552);
nand U5382 (N_5382,N_2032,N_2755);
or U5383 (N_5383,N_1041,N_9);
and U5384 (N_5384,N_2450,N_2117);
nor U5385 (N_5385,N_93,N_832);
and U5386 (N_5386,N_4895,N_3804);
or U5387 (N_5387,N_965,N_2234);
nand U5388 (N_5388,N_3508,N_3560);
nand U5389 (N_5389,N_786,N_2549);
or U5390 (N_5390,N_3629,N_1259);
xnor U5391 (N_5391,N_2486,N_540);
and U5392 (N_5392,N_2316,N_1224);
xnor U5393 (N_5393,N_4525,N_4768);
or U5394 (N_5394,N_1034,N_4039);
nor U5395 (N_5395,N_1345,N_1615);
nand U5396 (N_5396,N_873,N_411);
nand U5397 (N_5397,N_4043,N_4242);
or U5398 (N_5398,N_4681,N_2444);
nor U5399 (N_5399,N_3258,N_2664);
nand U5400 (N_5400,N_4584,N_1930);
or U5401 (N_5401,N_3852,N_924);
xnor U5402 (N_5402,N_2975,N_2775);
xor U5403 (N_5403,N_598,N_4715);
and U5404 (N_5404,N_2012,N_4118);
or U5405 (N_5405,N_943,N_1871);
nor U5406 (N_5406,N_2158,N_2523);
xnor U5407 (N_5407,N_4198,N_2301);
nor U5408 (N_5408,N_4679,N_3453);
nor U5409 (N_5409,N_3776,N_2797);
xnor U5410 (N_5410,N_1327,N_223);
and U5411 (N_5411,N_116,N_641);
and U5412 (N_5412,N_340,N_3680);
nand U5413 (N_5413,N_741,N_4561);
and U5414 (N_5414,N_2925,N_1945);
nor U5415 (N_5415,N_3148,N_4764);
xor U5416 (N_5416,N_2005,N_222);
nand U5417 (N_5417,N_3834,N_1295);
nand U5418 (N_5418,N_3406,N_2803);
nor U5419 (N_5419,N_3452,N_4592);
and U5420 (N_5420,N_1063,N_620);
nand U5421 (N_5421,N_2283,N_495);
or U5422 (N_5422,N_4920,N_265);
or U5423 (N_5423,N_1068,N_1333);
or U5424 (N_5424,N_4453,N_3257);
nor U5425 (N_5425,N_4438,N_1789);
nand U5426 (N_5426,N_434,N_1448);
nand U5427 (N_5427,N_4342,N_612);
and U5428 (N_5428,N_4526,N_3401);
or U5429 (N_5429,N_1451,N_1496);
xor U5430 (N_5430,N_1740,N_3034);
nor U5431 (N_5431,N_2108,N_583);
or U5432 (N_5432,N_4994,N_1527);
nand U5433 (N_5433,N_3412,N_575);
and U5434 (N_5434,N_2773,N_4919);
nor U5435 (N_5435,N_4857,N_2300);
xor U5436 (N_5436,N_1482,N_3822);
xor U5437 (N_5437,N_4127,N_3122);
xnor U5438 (N_5438,N_1174,N_4618);
xor U5439 (N_5439,N_3929,N_4371);
nor U5440 (N_5440,N_2167,N_135);
nand U5441 (N_5441,N_287,N_4684);
or U5442 (N_5442,N_527,N_342);
nor U5443 (N_5443,N_2714,N_3176);
xnor U5444 (N_5444,N_1600,N_1671);
and U5445 (N_5445,N_935,N_333);
nand U5446 (N_5446,N_2864,N_3549);
nand U5447 (N_5447,N_4195,N_2208);
and U5448 (N_5448,N_545,N_4269);
nand U5449 (N_5449,N_2438,N_3374);
xnor U5450 (N_5450,N_4966,N_4098);
and U5451 (N_5451,N_1397,N_2103);
xnor U5452 (N_5452,N_4837,N_3501);
and U5453 (N_5453,N_4402,N_1676);
nand U5454 (N_5454,N_2000,N_726);
nand U5455 (N_5455,N_4222,N_2735);
nor U5456 (N_5456,N_489,N_233);
or U5457 (N_5457,N_2290,N_4496);
or U5458 (N_5458,N_3964,N_1551);
nand U5459 (N_5459,N_1512,N_1298);
or U5460 (N_5460,N_1828,N_728);
nand U5461 (N_5461,N_363,N_4353);
nor U5462 (N_5462,N_4182,N_4479);
nand U5463 (N_5463,N_2119,N_164);
xor U5464 (N_5464,N_950,N_1964);
and U5465 (N_5465,N_1845,N_1474);
and U5466 (N_5466,N_1738,N_2374);
xnor U5467 (N_5467,N_3247,N_4437);
xnor U5468 (N_5468,N_127,N_968);
or U5469 (N_5469,N_4623,N_2106);
nor U5470 (N_5470,N_4698,N_537);
nand U5471 (N_5471,N_3024,N_948);
xnor U5472 (N_5472,N_1923,N_3534);
nor U5473 (N_5473,N_587,N_3885);
nand U5474 (N_5474,N_4833,N_4866);
xnor U5475 (N_5475,N_696,N_4960);
nor U5476 (N_5476,N_2712,N_3942);
nand U5477 (N_5477,N_153,N_371);
nand U5478 (N_5478,N_2675,N_4405);
and U5479 (N_5479,N_191,N_3131);
nor U5480 (N_5480,N_2148,N_3298);
nor U5481 (N_5481,N_1390,N_3304);
and U5482 (N_5482,N_2902,N_306);
nor U5483 (N_5483,N_3747,N_4729);
and U5484 (N_5484,N_2498,N_2462);
xor U5485 (N_5485,N_1769,N_3378);
xor U5486 (N_5486,N_1239,N_3213);
and U5487 (N_5487,N_3117,N_1509);
nand U5488 (N_5488,N_766,N_748);
xor U5489 (N_5489,N_2865,N_3016);
nor U5490 (N_5490,N_1840,N_1568);
nor U5491 (N_5491,N_1974,N_999);
and U5492 (N_5492,N_4313,N_1552);
nor U5493 (N_5493,N_2335,N_4932);
and U5494 (N_5494,N_1198,N_3949);
nand U5495 (N_5495,N_3239,N_4722);
xnor U5496 (N_5496,N_440,N_2499);
xnor U5497 (N_5497,N_2348,N_319);
and U5498 (N_5498,N_4316,N_2488);
xnor U5499 (N_5499,N_1508,N_43);
xnor U5500 (N_5500,N_2982,N_1300);
nand U5501 (N_5501,N_1371,N_278);
xor U5502 (N_5502,N_953,N_4163);
nor U5503 (N_5503,N_1246,N_3246);
nand U5504 (N_5504,N_744,N_1673);
or U5505 (N_5505,N_1175,N_402);
and U5506 (N_5506,N_4226,N_1510);
nor U5507 (N_5507,N_4459,N_4125);
nand U5508 (N_5508,N_3377,N_642);
and U5509 (N_5509,N_4497,N_1231);
nand U5510 (N_5510,N_480,N_913);
nand U5511 (N_5511,N_3240,N_205);
xnor U5512 (N_5512,N_2943,N_768);
nor U5513 (N_5513,N_4097,N_1440);
or U5514 (N_5514,N_2,N_3685);
xnor U5515 (N_5515,N_3591,N_4305);
nand U5516 (N_5516,N_1050,N_61);
and U5517 (N_5517,N_280,N_1648);
nand U5518 (N_5518,N_124,N_3614);
nand U5519 (N_5519,N_4196,N_3663);
and U5520 (N_5520,N_2731,N_4042);
xor U5521 (N_5521,N_4160,N_1873);
or U5522 (N_5522,N_556,N_4412);
nand U5523 (N_5523,N_3201,N_1851);
or U5524 (N_5524,N_3988,N_2559);
or U5525 (N_5525,N_360,N_2683);
nor U5526 (N_5526,N_1127,N_4019);
or U5527 (N_5527,N_3825,N_1215);
and U5528 (N_5528,N_500,N_2071);
nor U5529 (N_5529,N_2023,N_1118);
xnor U5530 (N_5530,N_2728,N_1924);
and U5531 (N_5531,N_3289,N_712);
and U5532 (N_5532,N_3559,N_564);
and U5533 (N_5533,N_179,N_2306);
nand U5534 (N_5534,N_2204,N_2717);
or U5535 (N_5535,N_3393,N_231);
or U5536 (N_5536,N_286,N_4891);
xnor U5537 (N_5537,N_1316,N_4767);
nor U5538 (N_5538,N_2799,N_4889);
and U5539 (N_5539,N_1319,N_1937);
nor U5540 (N_5540,N_823,N_458);
and U5541 (N_5541,N_4906,N_4925);
xor U5542 (N_5542,N_3165,N_1082);
or U5543 (N_5543,N_3991,N_3666);
nor U5544 (N_5544,N_1536,N_1353);
nor U5545 (N_5545,N_4820,N_2330);
and U5546 (N_5546,N_451,N_1725);
or U5547 (N_5547,N_4645,N_798);
nor U5548 (N_5548,N_522,N_1164);
nor U5549 (N_5549,N_4219,N_609);
or U5550 (N_5550,N_4617,N_4616);
and U5551 (N_5551,N_1480,N_3877);
xor U5552 (N_5552,N_4745,N_3388);
nor U5553 (N_5553,N_89,N_4812);
and U5554 (N_5554,N_3538,N_2540);
xor U5555 (N_5555,N_2402,N_4648);
nand U5556 (N_5556,N_3174,N_3761);
nand U5557 (N_5557,N_4365,N_1433);
or U5558 (N_5558,N_2170,N_3679);
nor U5559 (N_5559,N_1192,N_4362);
nand U5560 (N_5560,N_1473,N_2361);
xnor U5561 (N_5561,N_1699,N_524);
nand U5562 (N_5562,N_4289,N_4212);
nor U5563 (N_5563,N_2464,N_2122);
nor U5564 (N_5564,N_1883,N_1199);
nand U5565 (N_5565,N_4587,N_3349);
and U5566 (N_5566,N_1839,N_565);
and U5567 (N_5567,N_3055,N_2750);
nor U5568 (N_5568,N_272,N_1872);
xnor U5569 (N_5569,N_2944,N_1172);
xnor U5570 (N_5570,N_1220,N_2793);
or U5571 (N_5571,N_133,N_3445);
and U5572 (N_5572,N_2277,N_2929);
nand U5573 (N_5573,N_1126,N_2667);
xor U5574 (N_5574,N_4489,N_3746);
nor U5575 (N_5575,N_1597,N_4122);
xnor U5576 (N_5576,N_2962,N_2767);
and U5577 (N_5577,N_4711,N_216);
nand U5578 (N_5578,N_4022,N_3199);
nor U5579 (N_5579,N_1807,N_3652);
nand U5580 (N_5580,N_1321,N_312);
or U5581 (N_5581,N_3536,N_4429);
or U5582 (N_5582,N_1637,N_3479);
and U5583 (N_5583,N_4079,N_281);
nor U5584 (N_5584,N_2178,N_1988);
or U5585 (N_5585,N_655,N_4544);
xor U5586 (N_5586,N_1555,N_1376);
nor U5587 (N_5587,N_3677,N_2551);
and U5588 (N_5588,N_2852,N_2663);
nand U5589 (N_5589,N_2893,N_4117);
or U5590 (N_5590,N_4961,N_4598);
nor U5591 (N_5591,N_4814,N_1189);
nor U5592 (N_5592,N_4253,N_531);
nor U5593 (N_5593,N_169,N_3136);
nor U5594 (N_5594,N_307,N_3288);
or U5595 (N_5595,N_988,N_3941);
xnor U5596 (N_5596,N_4176,N_3714);
nor U5597 (N_5597,N_3535,N_4037);
xor U5598 (N_5598,N_1366,N_2861);
xor U5599 (N_5599,N_843,N_4930);
or U5600 (N_5600,N_1578,N_3592);
or U5601 (N_5601,N_1602,N_3170);
and U5602 (N_5602,N_3004,N_2197);
nor U5603 (N_5603,N_4254,N_92);
nand U5604 (N_5604,N_978,N_3637);
nand U5605 (N_5605,N_3732,N_2631);
nand U5606 (N_5606,N_4302,N_841);
and U5607 (N_5607,N_3341,N_3730);
nand U5608 (N_5608,N_3193,N_3426);
nor U5609 (N_5609,N_2657,N_44);
nor U5610 (N_5610,N_3745,N_894);
xnor U5611 (N_5611,N_1481,N_4542);
or U5612 (N_5612,N_2287,N_4264);
nor U5613 (N_5613,N_3676,N_4779);
xor U5614 (N_5614,N_70,N_1329);
nor U5615 (N_5615,N_2052,N_4640);
nand U5616 (N_5616,N_1272,N_4593);
and U5617 (N_5617,N_1678,N_491);
nor U5618 (N_5618,N_2292,N_2280);
or U5619 (N_5619,N_4940,N_436);
or U5620 (N_5620,N_2740,N_3263);
nand U5621 (N_5621,N_1755,N_3602);
nor U5622 (N_5622,N_989,N_4044);
nand U5623 (N_5623,N_1219,N_1304);
nor U5624 (N_5624,N_2192,N_697);
nor U5625 (N_5625,N_395,N_4771);
xor U5626 (N_5626,N_1092,N_1702);
nor U5627 (N_5627,N_47,N_4394);
or U5628 (N_5628,N_566,N_2582);
nand U5629 (N_5629,N_3292,N_1372);
nor U5630 (N_5630,N_1431,N_3777);
nand U5631 (N_5631,N_95,N_2154);
or U5632 (N_5632,N_3757,N_2333);
nand U5633 (N_5633,N_2120,N_2639);
and U5634 (N_5634,N_4747,N_1121);
and U5635 (N_5635,N_348,N_3124);
and U5636 (N_5636,N_853,N_4935);
xor U5637 (N_5637,N_3419,N_3774);
or U5638 (N_5638,N_4271,N_3228);
nor U5639 (N_5639,N_4591,N_1863);
and U5640 (N_5640,N_3948,N_586);
xnor U5641 (N_5641,N_856,N_549);
and U5642 (N_5642,N_4996,N_1502);
or U5643 (N_5643,N_1721,N_4886);
xor U5644 (N_5644,N_1382,N_46);
nor U5645 (N_5645,N_459,N_808);
nand U5646 (N_5646,N_2794,N_1953);
nand U5647 (N_5647,N_1756,N_4985);
nand U5648 (N_5648,N_4028,N_2407);
or U5649 (N_5649,N_2161,N_475);
xor U5650 (N_5650,N_237,N_3661);
or U5651 (N_5651,N_1854,N_2668);
nor U5652 (N_5652,N_3656,N_3696);
nand U5653 (N_5653,N_2589,N_4803);
nand U5654 (N_5654,N_2629,N_3765);
and U5655 (N_5655,N_4126,N_3550);
nand U5656 (N_5656,N_971,N_1262);
xnor U5657 (N_5657,N_2726,N_1497);
nand U5658 (N_5658,N_3135,N_4942);
nand U5659 (N_5659,N_4528,N_397);
xnor U5660 (N_5660,N_1784,N_4510);
nor U5661 (N_5661,N_4844,N_1229);
xnor U5662 (N_5662,N_1350,N_2293);
nor U5663 (N_5663,N_4633,N_282);
nor U5664 (N_5664,N_2858,N_1180);
and U5665 (N_5665,N_4448,N_64);
or U5666 (N_5666,N_3903,N_2298);
xor U5667 (N_5667,N_3269,N_457);
and U5668 (N_5668,N_4227,N_2168);
or U5669 (N_5669,N_865,N_3114);
nor U5670 (N_5670,N_2874,N_3711);
nor U5671 (N_5671,N_1645,N_2965);
or U5672 (N_5672,N_2338,N_855);
nor U5673 (N_5673,N_3072,N_3647);
xor U5674 (N_5674,N_2329,N_3251);
and U5675 (N_5675,N_2695,N_3650);
nand U5676 (N_5676,N_668,N_862);
nor U5677 (N_5677,N_370,N_2319);
or U5678 (N_5678,N_4221,N_4333);
nor U5679 (N_5679,N_3274,N_283);
xnor U5680 (N_5680,N_1225,N_3689);
xor U5681 (N_5681,N_4045,N_4512);
and U5682 (N_5682,N_380,N_4727);
nand U5683 (N_5683,N_919,N_1968);
xor U5684 (N_5684,N_1485,N_1791);
and U5685 (N_5685,N_657,N_4947);
xor U5686 (N_5686,N_2472,N_4388);
nor U5687 (N_5687,N_3710,N_1823);
xnor U5688 (N_5688,N_3311,N_1247);
nand U5689 (N_5689,N_652,N_4080);
nand U5690 (N_5690,N_561,N_1879);
xnor U5691 (N_5691,N_3261,N_2661);
xor U5692 (N_5692,N_1173,N_1292);
nand U5693 (N_5693,N_4320,N_2790);
or U5694 (N_5694,N_1621,N_3161);
xor U5695 (N_5695,N_3545,N_944);
and U5696 (N_5696,N_98,N_4898);
nor U5697 (N_5697,N_1768,N_2410);
and U5698 (N_5698,N_3324,N_1956);
nor U5699 (N_5699,N_2611,N_2817);
and U5700 (N_5700,N_2939,N_1558);
or U5701 (N_5701,N_3628,N_431);
nor U5702 (N_5702,N_1891,N_4225);
or U5703 (N_5703,N_2654,N_3039);
nor U5704 (N_5704,N_2155,N_536);
xor U5705 (N_5705,N_812,N_1322);
nor U5706 (N_5706,N_4533,N_2074);
xor U5707 (N_5707,N_4259,N_1548);
and U5708 (N_5708,N_2255,N_2771);
nand U5709 (N_5709,N_3640,N_4652);
xnor U5710 (N_5710,N_1591,N_3514);
nor U5711 (N_5711,N_4504,N_1138);
nor U5712 (N_5712,N_3939,N_138);
or U5713 (N_5713,N_1238,N_2890);
or U5714 (N_5714,N_114,N_1094);
nand U5715 (N_5715,N_4801,N_2956);
xor U5716 (N_5716,N_3030,N_725);
or U5717 (N_5717,N_1672,N_4766);
nand U5718 (N_5718,N_187,N_4815);
or U5719 (N_5719,N_4554,N_4548);
xor U5720 (N_5720,N_3446,N_3196);
and U5721 (N_5721,N_3934,N_1158);
nand U5722 (N_5722,N_3224,N_1917);
nand U5723 (N_5723,N_1835,N_4641);
xor U5724 (N_5724,N_2476,N_1516);
nor U5725 (N_5725,N_3509,N_2452);
or U5726 (N_5726,N_4087,N_1986);
and U5727 (N_5727,N_3492,N_3579);
nand U5728 (N_5728,N_2791,N_826);
xor U5729 (N_5729,N_3626,N_3156);
xnor U5730 (N_5730,N_3112,N_520);
or U5731 (N_5731,N_1283,N_3003);
nand U5732 (N_5732,N_4487,N_259);
nand U5733 (N_5733,N_3972,N_1020);
and U5734 (N_5734,N_2953,N_3790);
nor U5735 (N_5735,N_2143,N_4987);
xor U5736 (N_5736,N_4446,N_3147);
xor U5737 (N_5737,N_2736,N_4629);
or U5738 (N_5738,N_1852,N_465);
nor U5739 (N_5739,N_1286,N_2034);
or U5740 (N_5740,N_2588,N_1488);
xor U5741 (N_5741,N_4535,N_4071);
and U5742 (N_5742,N_3725,N_2584);
nand U5743 (N_5743,N_2867,N_690);
nand U5744 (N_5744,N_3874,N_2136);
xnor U5745 (N_5745,N_316,N_4849);
or U5746 (N_5746,N_139,N_3164);
nand U5747 (N_5747,N_4164,N_2826);
nor U5748 (N_5748,N_1104,N_4596);
or U5749 (N_5749,N_4472,N_922);
and U5750 (N_5750,N_1908,N_314);
nand U5751 (N_5751,N_3391,N_3139);
nor U5752 (N_5752,N_2545,N_4813);
and U5753 (N_5753,N_2428,N_1393);
nand U5754 (N_5754,N_3557,N_3967);
xnor U5755 (N_5755,N_7,N_3520);
xor U5756 (N_5756,N_787,N_917);
and U5757 (N_5757,N_3610,N_241);
nor U5758 (N_5758,N_2015,N_1778);
and U5759 (N_5759,N_1572,N_2350);
and U5760 (N_5760,N_1133,N_4778);
and U5761 (N_5761,N_1194,N_428);
xor U5762 (N_5762,N_2607,N_4345);
xnor U5763 (N_5763,N_1652,N_2763);
nand U5764 (N_5764,N_874,N_1414);
nor U5765 (N_5765,N_1026,N_3861);
xnor U5766 (N_5766,N_2276,N_2241);
or U5767 (N_5767,N_3919,N_3115);
xor U5768 (N_5768,N_1083,N_3278);
xnor U5769 (N_5769,N_3081,N_4491);
or U5770 (N_5770,N_4055,N_647);
nand U5771 (N_5771,N_636,N_2356);
or U5772 (N_5772,N_2572,N_376);
nand U5773 (N_5773,N_250,N_3782);
nor U5774 (N_5774,N_3983,N_1006);
and U5775 (N_5775,N_4769,N_4840);
nor U5776 (N_5776,N_1003,N_829);
or U5777 (N_5777,N_4082,N_1825);
nor U5778 (N_5778,N_1817,N_1834);
and U5779 (N_5779,N_4829,N_1200);
nor U5780 (N_5780,N_1870,N_3367);
or U5781 (N_5781,N_1999,N_4441);
nor U5782 (N_5782,N_2918,N_3370);
xor U5783 (N_5783,N_1882,N_2219);
and U5784 (N_5784,N_2676,N_2249);
nand U5785 (N_5785,N_2947,N_1087);
or U5786 (N_5786,N_2784,N_337);
nor U5787 (N_5787,N_645,N_3718);
xnor U5788 (N_5788,N_329,N_1950);
or U5789 (N_5789,N_2412,N_1131);
nor U5790 (N_5790,N_2095,N_486);
or U5791 (N_5791,N_4011,N_3396);
nand U5792 (N_5792,N_3315,N_3380);
nand U5793 (N_5793,N_2958,N_870);
nor U5794 (N_5794,N_4001,N_709);
or U5795 (N_5795,N_3970,N_674);
or U5796 (N_5796,N_426,N_4798);
xor U5797 (N_5797,N_4057,N_4998);
and U5798 (N_5798,N_2733,N_816);
and U5799 (N_5799,N_3285,N_810);
nor U5800 (N_5800,N_4414,N_168);
nand U5801 (N_5801,N_4824,N_4211);
and U5802 (N_5802,N_4624,N_3091);
and U5803 (N_5803,N_3749,N_779);
nor U5804 (N_5804,N_1115,N_1909);
nor U5805 (N_5805,N_2358,N_603);
xnor U5806 (N_5806,N_2818,N_523);
or U5807 (N_5807,N_322,N_1918);
or U5808 (N_5808,N_701,N_2619);
nand U5809 (N_5809,N_3119,N_1468);
or U5810 (N_5810,N_1110,N_2430);
nand U5811 (N_5811,N_3169,N_581);
or U5812 (N_5812,N_3280,N_1154);
xnor U5813 (N_5813,N_3580,N_3795);
or U5814 (N_5814,N_570,N_2655);
or U5815 (N_5815,N_800,N_120);
or U5816 (N_5816,N_423,N_2404);
or U5817 (N_5817,N_2033,N_2651);
nand U5818 (N_5818,N_3598,N_576);
xor U5819 (N_5819,N_3097,N_2528);
xor U5820 (N_5820,N_3662,N_4229);
nor U5821 (N_5821,N_4175,N_4827);
and U5822 (N_5822,N_2180,N_3528);
nand U5823 (N_5823,N_3301,N_1962);
nand U5824 (N_5824,N_1029,N_3976);
nor U5825 (N_5825,N_1443,N_1938);
or U5826 (N_5826,N_4004,N_3218);
or U5827 (N_5827,N_3109,N_2839);
or U5828 (N_5828,N_1169,N_3049);
nand U5829 (N_5829,N_518,N_4486);
or U5830 (N_5830,N_324,N_1783);
xnor U5831 (N_5831,N_958,N_2371);
xnor U5832 (N_5832,N_4358,N_2062);
nand U5833 (N_5833,N_2543,N_3657);
nand U5834 (N_5834,N_3820,N_2053);
xor U5835 (N_5835,N_3600,N_4475);
xnor U5836 (N_5836,N_682,N_991);
or U5837 (N_5837,N_3061,N_3668);
and U5838 (N_5838,N_104,N_163);
xor U5839 (N_5839,N_2202,N_720);
or U5840 (N_5840,N_3699,N_3633);
nand U5841 (N_5841,N_2087,N_4026);
nand U5842 (N_5842,N_130,N_4549);
nor U5843 (N_5843,N_4830,N_2896);
and U5844 (N_5844,N_4467,N_3390);
xnor U5845 (N_5845,N_1687,N_1385);
nor U5846 (N_5846,N_2396,N_1663);
nand U5847 (N_5847,N_4817,N_3713);
or U5848 (N_5848,N_3428,N_3358);
nor U5849 (N_5849,N_1217,N_2706);
xor U5850 (N_5850,N_1798,N_2085);
xnor U5851 (N_5851,N_3466,N_1822);
xnor U5852 (N_5852,N_961,N_3005);
and U5853 (N_5853,N_3845,N_1709);
nand U5854 (N_5854,N_4714,N_562);
nor U5855 (N_5855,N_2233,N_4989);
xor U5856 (N_5856,N_1586,N_3674);
nand U5857 (N_5857,N_1537,N_327);
nand U5858 (N_5858,N_1264,N_1715);
or U5859 (N_5859,N_3862,N_4569);
and U5860 (N_5860,N_3712,N_2862);
xnor U5861 (N_5861,N_4424,N_4567);
or U5862 (N_5862,N_432,N_3695);
nand U5863 (N_5863,N_782,N_2384);
or U5864 (N_5864,N_1989,N_4755);
and U5865 (N_5865,N_4341,N_4983);
nor U5866 (N_5866,N_4329,N_3322);
xor U5867 (N_5867,N_2099,N_3986);
and U5868 (N_5868,N_1308,N_3572);
and U5869 (N_5869,N_4081,N_1237);
nand U5870 (N_5870,N_534,N_1664);
and U5871 (N_5871,N_3915,N_4216);
nand U5872 (N_5872,N_1903,N_2905);
nand U5873 (N_5873,N_2240,N_476);
and U5874 (N_5874,N_3352,N_1465);
xnor U5875 (N_5875,N_3891,N_404);
and U5876 (N_5876,N_1406,N_3485);
and U5877 (N_5877,N_110,N_3998);
nand U5878 (N_5878,N_2454,N_2278);
nor U5879 (N_5879,N_2984,N_330);
xor U5880 (N_5880,N_2575,N_1939);
nand U5881 (N_5881,N_3806,N_90);
nand U5882 (N_5882,N_3044,N_1086);
or U5883 (N_5883,N_2538,N_1992);
and U5884 (N_5884,N_1629,N_3499);
xor U5885 (N_5885,N_3060,N_8);
and U5886 (N_5886,N_3118,N_1833);
xor U5887 (N_5887,N_4084,N_1780);
or U5888 (N_5888,N_236,N_3551);
xor U5889 (N_5889,N_3904,N_3070);
and U5890 (N_5890,N_1389,N_496);
xnor U5891 (N_5891,N_2594,N_771);
xnor U5892 (N_5892,N_3192,N_621);
nand U5893 (N_5893,N_2048,N_3036);
or U5894 (N_5894,N_4964,N_4301);
nor U5895 (N_5895,N_521,N_4283);
and U5896 (N_5896,N_925,N_4708);
and U5897 (N_5897,N_2282,N_4121);
xor U5898 (N_5898,N_4962,N_3329);
or U5899 (N_5899,N_654,N_4995);
nand U5900 (N_5900,N_4608,N_106);
xnor U5901 (N_5901,N_2883,N_1265);
and U5902 (N_5902,N_3211,N_938);
nor U5903 (N_5903,N_349,N_532);
and U5904 (N_5904,N_906,N_3319);
and U5905 (N_5905,N_1042,N_757);
xor U5906 (N_5906,N_450,N_2570);
xor U5907 (N_5907,N_4155,N_3129);
nor U5908 (N_5908,N_4520,N_4795);
nor U5909 (N_5909,N_3241,N_2525);
or U5910 (N_5910,N_3262,N_4419);
nor U5911 (N_5911,N_197,N_3048);
nor U5912 (N_5912,N_3339,N_700);
nand U5913 (N_5913,N_755,N_3461);
nand U5914 (N_5914,N_1521,N_1141);
and U5915 (N_5915,N_907,N_3340);
or U5916 (N_5916,N_3063,N_4565);
or U5917 (N_5917,N_3641,N_4319);
or U5918 (N_5918,N_2618,N_1611);
xnor U5919 (N_5919,N_2801,N_2973);
nor U5920 (N_5920,N_1518,N_4324);
nor U5921 (N_5921,N_4941,N_2964);
xor U5922 (N_5922,N_1391,N_3634);
nand U5923 (N_5923,N_4601,N_526);
xnor U5924 (N_5924,N_3596,N_2972);
nor U5925 (N_5925,N_639,N_470);
and U5926 (N_5926,N_699,N_3144);
xor U5927 (N_5927,N_1075,N_3739);
nand U5928 (N_5928,N_257,N_3826);
nor U5929 (N_5929,N_2195,N_149);
nand U5930 (N_5930,N_157,N_2187);
xnor U5931 (N_5931,N_4425,N_4738);
xnor U5932 (N_5932,N_1785,N_2420);
or U5933 (N_5933,N_3337,N_1592);
nand U5934 (N_5934,N_663,N_1375);
nor U5935 (N_5935,N_4705,N_4112);
nor U5936 (N_5936,N_4531,N_4540);
and U5937 (N_5937,N_263,N_4089);
nor U5938 (N_5938,N_2586,N_3012);
nor U5939 (N_5939,N_634,N_4236);
or U5940 (N_5940,N_4279,N_485);
or U5941 (N_5941,N_1519,N_1604);
and U5942 (N_5942,N_4352,N_3575);
nand U5943 (N_5943,N_4428,N_1595);
nand U5944 (N_5944,N_3512,N_1243);
xor U5945 (N_5945,N_1478,N_4718);
nand U5946 (N_5946,N_507,N_3833);
and U5947 (N_5947,N_4481,N_2347);
or U5948 (N_5948,N_4774,N_1214);
xnor U5949 (N_5949,N_4202,N_2563);
and U5950 (N_5950,N_4465,N_838);
xnor U5951 (N_5951,N_3859,N_494);
nor U5952 (N_5952,N_2463,N_3486);
xnor U5953 (N_5953,N_1395,N_1010);
or U5954 (N_5954,N_1585,N_1940);
xnor U5955 (N_5955,N_2746,N_1384);
or U5956 (N_5956,N_1904,N_2907);
xor U5957 (N_5957,N_1686,N_253);
xnor U5958 (N_5958,N_1815,N_2043);
and U5959 (N_5959,N_4108,N_1727);
and U5960 (N_5960,N_2416,N_136);
and U5961 (N_5961,N_1013,N_50);
or U5962 (N_5962,N_3720,N_3281);
and U5963 (N_5963,N_814,N_758);
nand U5964 (N_5964,N_1570,N_1948);
nand U5965 (N_5965,N_326,N_3856);
nand U5966 (N_5966,N_1236,N_4929);
xnor U5967 (N_5967,N_1954,N_4506);
xor U5968 (N_5968,N_3474,N_4789);
nand U5969 (N_5969,N_4061,N_2640);
xnor U5970 (N_5970,N_3198,N_2700);
nand U5971 (N_5971,N_355,N_638);
xnor U5972 (N_5972,N_1553,N_1556);
nor U5973 (N_5973,N_4938,N_4731);
nand U5974 (N_5974,N_4083,N_4020);
nor U5975 (N_5975,N_1985,N_653);
nor U5976 (N_5976,N_723,N_4214);
xnor U5977 (N_5977,N_2889,N_3214);
or U5978 (N_5978,N_3900,N_4102);
xor U5979 (N_5979,N_1461,N_4389);
nor U5980 (N_5980,N_2656,N_4832);
or U5981 (N_5981,N_119,N_3697);
or U5982 (N_5982,N_2694,N_2625);
nand U5983 (N_5983,N_1787,N_1654);
and U5984 (N_5984,N_2687,N_1906);
xnor U5985 (N_5985,N_3227,N_1540);
xnor U5986 (N_5986,N_3980,N_1946);
and U5987 (N_5987,N_1005,N_1935);
and U5988 (N_5988,N_847,N_2604);
or U5989 (N_5989,N_1056,N_2081);
nor U5990 (N_5990,N_4490,N_3544);
and U5991 (N_5991,N_1970,N_1594);
nor U5992 (N_5992,N_1506,N_1921);
nor U5993 (N_5993,N_4238,N_4545);
or U5994 (N_5994,N_3219,N_3275);
or U5995 (N_5995,N_2141,N_1043);
and U5996 (N_5996,N_211,N_2747);
nand U5997 (N_5997,N_2159,N_2564);
nor U5998 (N_5998,N_517,N_4511);
and U5999 (N_5999,N_2814,N_1779);
nor U6000 (N_6000,N_3792,N_30);
nor U6001 (N_6001,N_878,N_1811);
nor U6002 (N_6002,N_4366,N_4368);
nor U6003 (N_6003,N_1662,N_1661);
xor U6004 (N_6004,N_746,N_3624);
nor U6005 (N_6005,N_1584,N_4582);
nor U6006 (N_6006,N_889,N_3120);
nor U6007 (N_6007,N_1949,N_3693);
or U6008 (N_6008,N_2094,N_3738);
xnor U6009 (N_6009,N_58,N_2312);
xnor U6010 (N_6010,N_1032,N_2340);
and U6011 (N_6011,N_1276,N_1387);
xor U6012 (N_6012,N_2960,N_4208);
and U6013 (N_6013,N_4694,N_69);
nor U6014 (N_6014,N_3125,N_1208);
xor U6015 (N_6015,N_3468,N_1266);
and U6016 (N_6016,N_664,N_2210);
nor U6017 (N_6017,N_1332,N_2459);
or U6018 (N_6018,N_4893,N_4758);
nor U6019 (N_6019,N_1079,N_4823);
or U6020 (N_6020,N_1330,N_2581);
nor U6021 (N_6021,N_4110,N_584);
nor U6022 (N_6022,N_2653,N_3541);
and U6023 (N_6023,N_4074,N_4945);
nand U6024 (N_6024,N_159,N_4901);
or U6025 (N_6025,N_4077,N_343);
xor U6026 (N_6026,N_656,N_3022);
xor U6027 (N_6027,N_818,N_1071);
or U6028 (N_6028,N_390,N_2377);
or U6029 (N_6029,N_3047,N_4303);
nor U6030 (N_6030,N_1700,N_1771);
or U6031 (N_6031,N_4686,N_1400);
or U6032 (N_6032,N_1751,N_232);
nor U6033 (N_6033,N_1748,N_3605);
or U6034 (N_6034,N_1335,N_4449);
nor U6035 (N_6035,N_4062,N_3824);
nor U6036 (N_6036,N_4147,N_1402);
or U6037 (N_6037,N_2489,N_3828);
or U6038 (N_6038,N_1640,N_2696);
or U6039 (N_6039,N_2165,N_4291);
nand U6040 (N_6040,N_1444,N_2429);
nor U6041 (N_6041,N_3484,N_2922);
nand U6042 (N_6042,N_1274,N_4716);
nor U6043 (N_6043,N_3955,N_2936);
or U6044 (N_6044,N_2137,N_2050);
xnor U6045 (N_6045,N_4922,N_271);
and U6046 (N_6046,N_3642,N_4484);
and U6047 (N_6047,N_904,N_3107);
xnor U6048 (N_6048,N_182,N_3606);
and U6049 (N_6049,N_4244,N_1099);
nor U6050 (N_6050,N_3925,N_4017);
xnor U6051 (N_6051,N_210,N_805);
and U6052 (N_6052,N_834,N_707);
or U6053 (N_6053,N_3140,N_2114);
nand U6054 (N_6054,N_4218,N_406);
or U6055 (N_6055,N_2441,N_2603);
nor U6056 (N_6056,N_220,N_4637);
nand U6057 (N_6057,N_2010,N_2691);
nand U6058 (N_6058,N_2267,N_1743);
nor U6059 (N_6059,N_2205,N_848);
nand U6060 (N_6060,N_2991,N_1982);
or U6061 (N_6061,N_102,N_2553);
nor U6062 (N_6062,N_1877,N_3664);
nand U6063 (N_6063,N_4132,N_3134);
xnor U6064 (N_6064,N_959,N_2928);
and U6065 (N_6065,N_1983,N_2190);
or U6066 (N_6066,N_296,N_3173);
and U6067 (N_6067,N_2723,N_1853);
or U6068 (N_6068,N_4859,N_3209);
xnor U6069 (N_6069,N_2203,N_289);
nand U6070 (N_6070,N_1392,N_3568);
nand U6071 (N_6071,N_1492,N_3327);
or U6072 (N_6072,N_1240,N_3052);
nor U6073 (N_6073,N_3386,N_3425);
xor U6074 (N_6074,N_722,N_1899);
nand U6075 (N_6075,N_2304,N_4890);
nor U6076 (N_6076,N_2809,N_3405);
xor U6077 (N_6077,N_3456,N_3454);
or U6078 (N_6078,N_940,N_1352);
nor U6079 (N_6079,N_615,N_1731);
and U6080 (N_6080,N_849,N_4793);
nor U6081 (N_6081,N_4967,N_703);
nor U6082 (N_6082,N_4171,N_2013);
and U6083 (N_6083,N_4142,N_1197);
nor U6084 (N_6084,N_1802,N_4749);
or U6085 (N_6085,N_3950,N_4806);
nand U6086 (N_6086,N_1449,N_377);
and U6087 (N_6087,N_4734,N_2917);
nand U6088 (N_6088,N_243,N_2440);
xor U6089 (N_6089,N_2624,N_3875);
nor U6090 (N_6090,N_1412,N_1567);
nand U6091 (N_6091,N_1212,N_3607);
nor U6092 (N_6092,N_4398,N_4024);
or U6093 (N_6093,N_806,N_3230);
and U6094 (N_6094,N_3924,N_2526);
xor U6095 (N_6095,N_1881,N_632);
and U6096 (N_6096,N_4470,N_1430);
nor U6097 (N_6097,N_3071,N_3764);
nor U6098 (N_6098,N_2704,N_331);
or U6099 (N_6099,N_2509,N_3851);
and U6100 (N_6100,N_378,N_4457);
or U6101 (N_6101,N_1241,N_573);
nand U6102 (N_6102,N_3457,N_4390);
nor U6103 (N_6103,N_4915,N_923);
or U6104 (N_6104,N_4471,N_4104);
and U6105 (N_6105,N_4790,N_2967);
nand U6106 (N_6106,N_2218,N_4811);
xnor U6107 (N_6107,N_1675,N_4991);
nand U6108 (N_6108,N_2049,N_1139);
nand U6109 (N_6109,N_893,N_3435);
and U6110 (N_6110,N_2484,N_1257);
xnor U6111 (N_6111,N_3333,N_3392);
nor U6112 (N_6112,N_175,N_736);
xnor U6113 (N_6113,N_2066,N_4508);
nor U6114 (N_6114,N_3977,N_4753);
xor U6115 (N_6115,N_1064,N_1587);
nand U6116 (N_6116,N_4570,N_4800);
and U6117 (N_6117,N_1744,N_1358);
nor U6118 (N_6118,N_4907,N_4407);
xnor U6119 (N_6119,N_3611,N_3441);
and U6120 (N_6120,N_3644,N_3126);
nor U6121 (N_6121,N_2041,N_3756);
nor U6122 (N_6122,N_4206,N_1786);
nor U6123 (N_6123,N_2164,N_1024);
or U6124 (N_6124,N_239,N_508);
xnor U6125 (N_6125,N_3424,N_3558);
xor U6126 (N_6126,N_3041,N_2808);
and U6127 (N_6127,N_3821,N_248);
xnor U6128 (N_6128,N_2022,N_796);
or U6129 (N_6129,N_295,N_1991);
and U6130 (N_6130,N_2576,N_3268);
or U6131 (N_6131,N_3491,N_702);
xor U6132 (N_6132,N_2230,N_1800);
xor U6133 (N_6133,N_1829,N_97);
xnor U6134 (N_6134,N_4180,N_1011);
nand U6135 (N_6135,N_4036,N_392);
and U6136 (N_6136,N_881,N_4607);
nor U6137 (N_6137,N_2777,N_4739);
xnor U6138 (N_6138,N_4194,N_2567);
or U6139 (N_6139,N_4403,N_3684);
xnor U6140 (N_6140,N_2061,N_2709);
nand U6141 (N_6141,N_2485,N_2910);
xnor U6142 (N_6142,N_4969,N_1273);
nand U6143 (N_6143,N_1405,N_2495);
or U6144 (N_6144,N_4992,N_448);
or U6145 (N_6145,N_1550,N_437);
xor U6146 (N_6146,N_3272,N_3318);
and U6147 (N_6147,N_1008,N_1624);
and U6148 (N_6148,N_1997,N_2878);
and U6149 (N_6149,N_1583,N_438);
or U6150 (N_6150,N_1943,N_3800);
or U6151 (N_6151,N_4916,N_3105);
xnor U6152 (N_6152,N_3092,N_3181);
and U6153 (N_6153,N_3574,N_4488);
or U6154 (N_6154,N_3154,N_1520);
xor U6155 (N_6155,N_3507,N_1315);
and U6156 (N_6156,N_563,N_2800);
nor U6157 (N_6157,N_2995,N_4205);
or U6158 (N_6158,N_3095,N_4191);
or U6159 (N_6159,N_4167,N_156);
xnor U6160 (N_6160,N_743,N_582);
nand U6161 (N_6161,N_661,N_3914);
and U6162 (N_6162,N_1776,N_2036);
nor U6163 (N_6163,N_4970,N_2453);
and U6164 (N_6164,N_2719,N_996);
or U6165 (N_6165,N_132,N_3455);
or U6166 (N_6166,N_2992,N_4247);
or U6167 (N_6167,N_4263,N_1693);
and U6168 (N_6168,N_2556,N_942);
nor U6169 (N_6169,N_1437,N_528);
and U6170 (N_6170,N_1947,N_4839);
nand U6171 (N_6171,N_1915,N_4307);
nor U6172 (N_6172,N_4553,N_3819);
and U6173 (N_6173,N_957,N_714);
and U6174 (N_6174,N_1320,N_137);
nand U6175 (N_6175,N_2142,N_172);
or U6176 (N_6176,N_4327,N_62);
xnor U6177 (N_6177,N_3781,N_3813);
xor U6178 (N_6178,N_4131,N_4736);
xor U6179 (N_6179,N_36,N_4973);
and U6180 (N_6180,N_4381,N_2437);
nor U6181 (N_6181,N_1896,N_4499);
nor U6182 (N_6182,N_3045,N_1420);
nand U6183 (N_6183,N_2707,N_1547);
and U6184 (N_6184,N_23,N_734);
nor U6185 (N_6185,N_2660,N_1733);
and U6186 (N_6186,N_764,N_4444);
or U6187 (N_6187,N_2977,N_2067);
nand U6188 (N_6188,N_3658,N_2446);
and U6189 (N_6189,N_1232,N_762);
nor U6190 (N_6190,N_2352,N_618);
xor U6191 (N_6191,N_1459,N_3447);
xnor U6192 (N_6192,N_57,N_1832);
and U6193 (N_6193,N_2802,N_3649);
nand U6194 (N_6194,N_2648,N_3185);
nor U6195 (N_6195,N_658,N_3394);
and U6196 (N_6196,N_3518,N_2807);
or U6197 (N_6197,N_686,N_113);
xnor U6198 (N_6198,N_4776,N_2214);
or U6199 (N_6199,N_3769,N_1182);
nor U6200 (N_6200,N_1902,N_2045);
and U6201 (N_6201,N_2388,N_1435);
and U6202 (N_6202,N_415,N_3621);
nor U6203 (N_6203,N_4534,N_1306);
nor U6204 (N_6204,N_54,N_101);
xnor U6205 (N_6205,N_578,N_799);
nand U6206 (N_6206,N_4173,N_4717);
or U6207 (N_6207,N_567,N_695);
xnor U6208 (N_6208,N_1772,N_478);
nor U6209 (N_6209,N_1337,N_2318);
and U6210 (N_6210,N_2270,N_4826);
and U6211 (N_6211,N_1569,N_2642);
and U6212 (N_6212,N_4300,N_1588);
nor U6213 (N_6213,N_4651,N_1764);
or U6214 (N_6214,N_4349,N_2617);
nand U6215 (N_6215,N_3075,N_710);
or U6216 (N_6216,N_2310,N_369);
xnor U6217 (N_6217,N_2840,N_2876);
and U6218 (N_6218,N_3748,N_3354);
xor U6219 (N_6219,N_4720,N_973);
or U6220 (N_6220,N_4957,N_1869);
nand U6221 (N_6221,N_3279,N_2981);
xnor U6222 (N_6222,N_3581,N_4958);
and U6223 (N_6223,N_3336,N_3516);
nor U6224 (N_6224,N_2632,N_202);
nand U6225 (N_6225,N_1500,N_2468);
and U6226 (N_6226,N_3132,N_590);
nor U6227 (N_6227,N_4030,N_1655);
nor U6228 (N_6228,N_4666,N_1573);
and U6229 (N_6229,N_2264,N_75);
nand U6230 (N_6230,N_1515,N_4610);
or U6231 (N_6231,N_2544,N_1256);
nand U6232 (N_6232,N_2637,N_425);
nand U6233 (N_6233,N_4150,N_947);
xor U6234 (N_6234,N_375,N_4626);
or U6235 (N_6235,N_266,N_2963);
nand U6236 (N_6236,N_3750,N_4059);
and U6237 (N_6237,N_2035,N_4455);
nor U6238 (N_6238,N_2307,N_4541);
and U6239 (N_6239,N_706,N_1864);
and U6240 (N_6240,N_1271,N_3526);
and U6241 (N_6241,N_1714,N_2083);
xor U6242 (N_6242,N_4308,N_1098);
and U6243 (N_6243,N_2682,N_3908);
nor U6244 (N_6244,N_2211,N_2829);
and U6245 (N_6245,N_4144,N_4050);
and U6246 (N_6246,N_2251,N_1758);
nand U6247 (N_6247,N_2026,N_1424);
nor U6248 (N_6248,N_2424,N_926);
or U6249 (N_6249,N_3473,N_1221);
or U6250 (N_6250,N_4392,N_1088);
nor U6251 (N_6251,N_4975,N_2284);
or U6252 (N_6252,N_984,N_4474);
and U6253 (N_6253,N_4272,N_1081);
or U6254 (N_6254,N_1759,N_1190);
or U6255 (N_6255,N_111,N_1838);
xor U6256 (N_6256,N_3926,N_4804);
or U6257 (N_6257,N_2098,N_2515);
nand U6258 (N_6258,N_718,N_3724);
and U6259 (N_6259,N_1401,N_2901);
xnor U6260 (N_6260,N_2239,N_2299);
nand U6261 (N_6261,N_2988,N_3742);
nor U6262 (N_6262,N_4997,N_3597);
nor U6263 (N_6263,N_4464,N_2046);
xor U6264 (N_6264,N_3420,N_1302);
or U6265 (N_6265,N_4468,N_4434);
or U6266 (N_6266,N_3195,N_4159);
xor U6267 (N_6267,N_1499,N_2003);
or U6268 (N_6268,N_2297,N_2367);
nor U6269 (N_6269,N_3217,N_2670);
and U6270 (N_6270,N_79,N_801);
and U6271 (N_6271,N_650,N_1599);
nand U6272 (N_6272,N_2987,N_1364);
or U6273 (N_6273,N_2899,N_1454);
and U6274 (N_6274,N_3651,N_2832);
nor U6275 (N_6275,N_3478,N_2605);
and U6276 (N_6276,N_3849,N_821);
nor U6277 (N_6277,N_2647,N_3382);
xor U6278 (N_6278,N_2281,N_665);
nor U6279 (N_6279,N_3481,N_2671);
and U6280 (N_6280,N_4581,N_3038);
and U6281 (N_6281,N_1165,N_1886);
or U6282 (N_6282,N_3480,N_2980);
xor U6283 (N_6283,N_770,N_1285);
xnor U6284 (N_6284,N_819,N_3053);
or U6285 (N_6285,N_4311,N_2127);
nand U6286 (N_6286,N_1270,N_339);
xnor U6287 (N_6287,N_837,N_1975);
or U6288 (N_6288,N_4620,N_905);
nand U6289 (N_6289,N_1684,N_204);
nor U6290 (N_6290,N_1130,N_2126);
nor U6291 (N_6291,N_1410,N_374);
nand U6292 (N_6292,N_3175,N_2606);
and U6293 (N_6293,N_2974,N_4702);
and U6294 (N_6294,N_4128,N_3421);
nand U6295 (N_6295,N_1090,N_2060);
xor U6296 (N_6296,N_1827,N_4835);
xor U6297 (N_6297,N_117,N_2400);
and U6298 (N_6298,N_2521,N_409);
nand U6299 (N_6299,N_2480,N_2892);
nand U6300 (N_6300,N_4473,N_4404);
or U6301 (N_6301,N_3905,N_511);
and U6302 (N_6302,N_1560,N_742);
nor U6303 (N_6303,N_4267,N_1911);
xor U6304 (N_6304,N_2247,N_490);
and U6305 (N_6305,N_2121,N_2353);
nor U6306 (N_6306,N_1455,N_1647);
and U6307 (N_6307,N_3671,N_1135);
and U6308 (N_6308,N_4794,N_38);
xor U6309 (N_6309,N_4306,N_4699);
nand U6310 (N_6310,N_2837,N_3212);
nand U6311 (N_6311,N_4007,N_2006);
and U6312 (N_6312,N_4568,N_398);
nand U6313 (N_6313,N_4124,N_817);
xnor U6314 (N_6314,N_4093,N_3308);
nand U6315 (N_6315,N_2751,N_276);
nor U6316 (N_6316,N_1415,N_692);
and U6317 (N_6317,N_218,N_4040);
nor U6318 (N_6318,N_1143,N_13);
nand U6319 (N_6319,N_4334,N_1525);
nor U6320 (N_6320,N_2592,N_3968);
or U6321 (N_6321,N_2810,N_3153);
nor U6322 (N_6322,N_2105,N_4659);
nor U6323 (N_6323,N_3102,N_997);
nand U6324 (N_6324,N_1290,N_4065);
nand U6325 (N_6325,N_442,N_519);
nand U6326 (N_6326,N_4270,N_1922);
nor U6327 (N_6327,N_3638,N_2162);
nor U6328 (N_6328,N_1325,N_679);
xnor U6329 (N_6329,N_1408,N_2153);
xnor U6330 (N_6330,N_759,N_3966);
nand U6331 (N_6331,N_1501,N_1291);
and U6332 (N_6332,N_2737,N_4450);
xor U6333 (N_6333,N_2457,N_3791);
nand U6334 (N_6334,N_1341,N_4304);
and U6335 (N_6335,N_1788,N_3810);
xor U6336 (N_6336,N_2693,N_3220);
xor U6337 (N_6337,N_3273,N_3830);
nor U6338 (N_6338,N_492,N_920);
xnor U6339 (N_6339,N_1074,N_1027);
and U6340 (N_6340,N_2291,N_4558);
nand U6341 (N_6341,N_3513,N_4594);
or U6342 (N_6342,N_2449,N_1388);
or U6343 (N_6343,N_4476,N_3880);
and U6344 (N_6344,N_1650,N_4393);
nand U6345 (N_6345,N_2866,N_2518);
xor U6346 (N_6346,N_2732,N_4347);
nor U6347 (N_6347,N_3255,N_760);
or U6348 (N_6348,N_4177,N_245);
nor U6349 (N_6349,N_4153,N_765);
nand U6350 (N_6350,N_140,N_1460);
or U6351 (N_6351,N_3577,N_1206);
nand U6352 (N_6352,N_4415,N_506);
nor U6353 (N_6353,N_4677,N_2877);
nand U6354 (N_6354,N_78,N_357);
and U6355 (N_6355,N_2079,N_795);
xor U6356 (N_6356,N_0,N_2630);
and U6357 (N_6357,N_2820,N_2643);
xnor U6358 (N_6358,N_180,N_186);
xor U6359 (N_6359,N_2391,N_3758);
nand U6360 (N_6360,N_1149,N_2101);
or U6361 (N_6361,N_4658,N_4675);
or U6362 (N_6362,N_2662,N_1226);
nor U6363 (N_6363,N_2188,N_2451);
xor U6364 (N_6364,N_3076,N_4517);
nand U6365 (N_6365,N_4355,N_3775);
and U6366 (N_6366,N_3152,N_3440);
or U6367 (N_6367,N_2252,N_2764);
xor U6368 (N_6368,N_2144,N_4430);
xnor U6369 (N_6369,N_1062,N_525);
nor U6370 (N_6370,N_2445,N_4466);
nand U6371 (N_6371,N_2916,N_780);
or U6372 (N_6372,N_3216,N_1004);
nor U6373 (N_6373,N_4924,N_4431);
and U6374 (N_6374,N_896,N_3672);
nor U6375 (N_6375,N_4363,N_2830);
or U6376 (N_6376,N_1897,N_225);
and U6377 (N_6377,N_4373,N_2957);
or U6378 (N_6378,N_3655,N_4148);
and U6379 (N_6379,N_128,N_4728);
and U6380 (N_6380,N_3913,N_4516);
and U6381 (N_6381,N_2224,N_666);
and U6382 (N_6382,N_3836,N_3653);
nor U6383 (N_6383,N_1114,N_1535);
nand U6384 (N_6384,N_3085,N_2431);
or U6385 (N_6385,N_1794,N_3619);
nand U6386 (N_6386,N_1689,N_4926);
nor U6387 (N_6387,N_4725,N_1734);
or U6388 (N_6388,N_4426,N_1176);
and U6389 (N_6389,N_2976,N_2123);
nor U6390 (N_6390,N_4501,N_2244);
nand U6391 (N_6391,N_4914,N_4621);
nand U6392 (N_6392,N_3562,N_424);
xnor U6393 (N_6393,N_928,N_3783);
nand U6394 (N_6394,N_433,N_439);
nand U6395 (N_6395,N_2482,N_261);
and U6396 (N_6396,N_195,N_2920);
nand U6397 (N_6397,N_3417,N_3110);
nand U6398 (N_6398,N_3338,N_539);
or U6399 (N_6399,N_2931,N_3043);
nor U6400 (N_6400,N_4606,N_1605);
and U6401 (N_6401,N_3146,N_3788);
nor U6402 (N_6402,N_3837,N_981);
or U6403 (N_6403,N_2983,N_1137);
or U6404 (N_6404,N_37,N_4781);
nor U6405 (N_6405,N_1207,N_3506);
nand U6406 (N_6406,N_4154,N_4331);
nand U6407 (N_6407,N_2635,N_559);
or U6408 (N_6408,N_68,N_1720);
and U6409 (N_6409,N_2533,N_1925);
and U6410 (N_6410,N_3471,N_3789);
nand U6411 (N_6411,N_2952,N_4518);
xor U6412 (N_6412,N_481,N_345);
nand U6413 (N_6413,N_2346,N_11);
or U6414 (N_6414,N_1713,N_955);
or U6415 (N_6415,N_1749,N_807);
nand U6416 (N_6416,N_3389,N_4136);
nand U6417 (N_6417,N_671,N_4865);
xor U6418 (N_6418,N_4443,N_285);
xor U6419 (N_6419,N_3694,N_3187);
nor U6420 (N_6420,N_2702,N_2532);
or U6421 (N_6421,N_974,N_4653);
nor U6422 (N_6422,N_4156,N_162);
and U6423 (N_6423,N_863,N_2259);
or U6424 (N_6424,N_3089,N_1790);
or U6425 (N_6425,N_4086,N_2258);
nand U6426 (N_6426,N_334,N_1416);
nand U6427 (N_6427,N_354,N_3381);
nand U6428 (N_6428,N_2679,N_850);
nor U6429 (N_6429,N_949,N_3051);
and U6430 (N_6430,N_3660,N_3876);
nand U6431 (N_6431,N_4977,N_2888);
and U6432 (N_6432,N_1717,N_3743);
and U6433 (N_6433,N_675,N_1612);
nor U6434 (N_6434,N_267,N_121);
nor U6435 (N_6435,N_876,N_1972);
xor U6436 (N_6436,N_3360,N_4937);
or U6437 (N_6437,N_3616,N_1177);
or U6438 (N_6438,N_4189,N_273);
nand U6439 (N_6439,N_2659,N_1379);
xnor U6440 (N_6440,N_4413,N_1927);
nor U6441 (N_6441,N_151,N_1752);
nand U6442 (N_6442,N_2331,N_3654);
or U6443 (N_6443,N_1514,N_2229);
xor U6444 (N_6444,N_4409,N_356);
xnor U6445 (N_6445,N_1166,N_32);
or U6446 (N_6446,N_2360,N_1680);
nand U6447 (N_6447,N_630,N_3084);
or U6448 (N_6448,N_3530,N_3893);
and U6449 (N_6449,N_2002,N_1589);
or U6450 (N_6450,N_3205,N_174);
nor U6451 (N_6451,N_857,N_264);
or U6452 (N_6452,N_900,N_4685);
xor U6453 (N_6453,N_918,N_2930);
and U6454 (N_6454,N_3869,N_3973);
nand U6455 (N_6455,N_4759,N_1490);
xnor U6456 (N_6456,N_2725,N_1228);
nor U6457 (N_6457,N_1955,N_4237);
nand U6458 (N_6458,N_212,N_3229);
nor U6459 (N_6459,N_4197,N_2473);
nand U6460 (N_6460,N_4029,N_1719);
nor U6461 (N_6461,N_3368,N_2881);
and U6462 (N_6462,N_4843,N_1209);
nand U6463 (N_6463,N_1546,N_977);
nand U6464 (N_6464,N_553,N_1462);
nor U6465 (N_6465,N_3066,N_4369);
xnor U6466 (N_6466,N_4538,N_1021);
and U6467 (N_6467,N_4784,N_249);
or U6468 (N_6468,N_1347,N_1269);
nor U6469 (N_6469,N_192,N_227);
and U6470 (N_6470,N_341,N_3028);
or U6471 (N_6471,N_1503,N_4730);
nand U6472 (N_6472,N_3307,N_3418);
nor U6473 (N_6473,N_1349,N_2708);
or U6474 (N_6474,N_3158,N_4288);
nor U6475 (N_6475,N_346,N_4408);
or U6476 (N_6476,N_3907,N_2175);
nand U6477 (N_6477,N_711,N_3143);
nor U6478 (N_6478,N_846,N_4557);
or U6479 (N_6479,N_4612,N_1035);
nand U6480 (N_6480,N_1355,N_4090);
xor U6481 (N_6481,N_2343,N_4013);
and U6482 (N_6482,N_1117,N_2753);
xor U6483 (N_6483,N_2398,N_1413);
nand U6484 (N_6484,N_4052,N_2344);
xnor U6485 (N_6485,N_1849,N_1531);
xor U6486 (N_6486,N_3404,N_336);
xnor U6487 (N_6487,N_4252,N_3245);
and U6488 (N_6488,N_4103,N_4281);
and U6489 (N_6489,N_2978,N_2181);
xnor U6490 (N_6490,N_4860,N_396);
nand U6491 (N_6491,N_4818,N_2891);
or U6492 (N_6492,N_290,N_1898);
or U6493 (N_6493,N_3707,N_2368);
xnor U6494 (N_6494,N_4477,N_3899);
nor U6495 (N_6495,N_1187,N_3796);
xnor U6496 (N_6496,N_2633,N_3040);
nor U6497 (N_6497,N_3079,N_3659);
nand U6498 (N_6498,N_2133,N_1533);
or U6499 (N_6499,N_2173,N_3846);
nand U6500 (N_6500,N_2672,N_4634);
and U6501 (N_6501,N_3042,N_1750);
nand U6502 (N_6502,N_2320,N_2075);
and U6503 (N_6503,N_1511,N_3729);
or U6504 (N_6504,N_513,N_533);
and U6505 (N_6505,N_934,N_3963);
and U6506 (N_6506,N_1718,N_879);
nand U6507 (N_6507,N_4078,N_769);
or U6508 (N_6508,N_386,N_1484);
nand U6509 (N_6509,N_4332,N_871);
or U6510 (N_6510,N_401,N_3771);
nand U6511 (N_6511,N_2836,N_4682);
xor U6512 (N_6512,N_4401,N_1309);
nor U6513 (N_6513,N_2399,N_2517);
nor U6514 (N_6514,N_194,N_3087);
nor U6515 (N_6515,N_1305,N_4014);
or U6516 (N_6516,N_1808,N_3431);
and U6517 (N_6517,N_613,N_1168);
xnor U6518 (N_6518,N_4025,N_4106);
or U6519 (N_6519,N_724,N_3369);
and U6520 (N_6520,N_4968,N_3400);
and U6521 (N_6521,N_3309,N_2176);
or U6522 (N_6522,N_951,N_2578);
and U6523 (N_6523,N_954,N_688);
and U6524 (N_6524,N_4872,N_1307);
xor U6525 (N_6525,N_2721,N_2541);
nor U6526 (N_6526,N_366,N_21);
nand U6527 (N_6527,N_4298,N_1342);
nand U6528 (N_6528,N_558,N_91);
nor U6529 (N_6529,N_3971,N_4875);
xnor U6530 (N_6530,N_3935,N_4848);
nand U6531 (N_6531,N_3794,N_2994);
or U6532 (N_6532,N_1910,N_49);
xor U6533 (N_6533,N_3571,N_3069);
and U6534 (N_6534,N_1111,N_4530);
or U6535 (N_6535,N_1263,N_4577);
and U6536 (N_6536,N_1830,N_2269);
xnor U6537 (N_6537,N_2819,N_3264);
nor U6538 (N_6538,N_4933,N_4143);
or U6539 (N_6539,N_2886,N_1892);
or U6540 (N_6540,N_3835,N_1848);
xnor U6541 (N_6541,N_479,N_3027);
xnor U6542 (N_6542,N_3918,N_577);
or U6543 (N_6543,N_1952,N_3909);
xnor U6544 (N_6544,N_4884,N_86);
and U6545 (N_6545,N_3816,N_4485);
and U6546 (N_6546,N_3138,N_2503);
or U6547 (N_6547,N_2780,N_4667);
nand U6548 (N_6548,N_4777,N_2626);
and U6549 (N_6549,N_4519,N_1522);
nand U6550 (N_6550,N_3944,N_3722);
nand U6551 (N_6551,N_224,N_2478);
nand U6552 (N_6552,N_551,N_3226);
nand U6553 (N_6553,N_34,N_3467);
xor U6554 (N_6554,N_2166,N_3728);
and U6555 (N_6555,N_3100,N_4680);
and U6556 (N_6556,N_3083,N_4151);
or U6557 (N_6557,N_1639,N_4546);
nor U6558 (N_6558,N_4493,N_2403);
nor U6559 (N_6559,N_2838,N_3434);
or U6560 (N_6560,N_2869,N_3189);
nand U6561 (N_6561,N_2387,N_1781);
nand U6562 (N_6562,N_1723,N_1770);
nor U6563 (N_6563,N_3525,N_4514);
xor U6564 (N_6564,N_1532,N_784);
or U6565 (N_6565,N_3232,N_560);
and U6566 (N_6566,N_1803,N_3031);
nor U6567 (N_6567,N_2998,N_2409);
nand U6568 (N_6568,N_3706,N_3916);
nand U6569 (N_6569,N_3645,N_3708);
nand U6570 (N_6570,N_1901,N_4284);
nand U6571 (N_6571,N_4831,N_1724);
or U6572 (N_6572,N_131,N_3814);
and U6573 (N_6573,N_4041,N_170);
and U6574 (N_6574,N_552,N_3249);
nor U6575 (N_6575,N_299,N_4693);
nand U6576 (N_6576,N_1439,N_2007);
nor U6577 (N_6577,N_4799,N_1299);
nor U6578 (N_6578,N_381,N_4101);
nand U6579 (N_6579,N_389,N_2823);
nand U6580 (N_6580,N_1757,N_2788);
and U6581 (N_6581,N_3465,N_3056);
nand U6582 (N_6582,N_2742,N_631);
nor U6583 (N_6583,N_87,N_781);
and U6584 (N_6584,N_1476,N_1294);
and U6585 (N_6585,N_828,N_4873);
nor U6586 (N_6586,N_4963,N_4224);
and U6587 (N_6587,N_669,N_4695);
xnor U6588 (N_6588,N_4782,N_3768);
nor U6589 (N_6589,N_3300,N_568);
nor U6590 (N_6590,N_4315,N_794);
xor U6591 (N_6591,N_3430,N_4669);
and U6592 (N_6592,N_4819,N_1889);
xnor U6593 (N_6593,N_3458,N_1159);
and U6594 (N_6594,N_3495,N_4846);
nor U6595 (N_6595,N_4335,N_1089);
or U6596 (N_6596,N_2196,N_555);
xnor U6597 (N_6597,N_1691,N_3766);
or U6598 (N_6598,N_1185,N_1538);
and U6599 (N_6599,N_2761,N_1566);
nor U6600 (N_6600,N_3570,N_3059);
or U6601 (N_6601,N_2286,N_1819);
or U6602 (N_6602,N_3797,N_2380);
xor U6603 (N_6603,N_1052,N_2068);
or U6604 (N_6604,N_3818,N_1407);
nor U6605 (N_6605,N_3449,N_3902);
xnor U6606 (N_6606,N_3323,N_3726);
or U6607 (N_6607,N_574,N_3578);
xor U6608 (N_6608,N_854,N_2414);
xor U6609 (N_6609,N_3802,N_4965);
and U6610 (N_6610,N_4032,N_1365);
nand U6611 (N_6611,N_852,N_3155);
nand U6612 (N_6612,N_3552,N_4070);
or U6613 (N_6613,N_4016,N_4241);
and U6614 (N_6614,N_2752,N_1017);
and U6615 (N_6615,N_1289,N_4354);
nand U6616 (N_6616,N_2738,N_1381);
or U6617 (N_6617,N_4643,N_3648);
and U6618 (N_6618,N_4719,N_2940);
and U6619 (N_6619,N_4344,N_235);
nor U6620 (N_6620,N_2989,N_3586);
or U6621 (N_6621,N_4047,N_2554);
nor U6622 (N_6622,N_887,N_3409);
nor U6623 (N_6623,N_228,N_1161);
or U6624 (N_6624,N_1140,N_3912);
or U6625 (N_6625,N_2390,N_2688);
and U6626 (N_6626,N_3808,N_3984);
or U6627 (N_6627,N_2225,N_3035);
xnor U6628 (N_6628,N_1171,N_48);
nand U6629 (N_6629,N_946,N_4296);
and U6630 (N_6630,N_1378,N_963);
and U6631 (N_6631,N_2113,N_4321);
nor U6632 (N_6632,N_3803,N_579);
xnor U6633 (N_6633,N_3609,N_2698);
xor U6634 (N_6634,N_3603,N_1023);
nand U6635 (N_6635,N_269,N_3593);
xor U6636 (N_6636,N_4573,N_3244);
and U6637 (N_6637,N_2317,N_1862);
xor U6638 (N_6638,N_3786,N_3623);
nor U6639 (N_6639,N_3716,N_4012);
or U6640 (N_6640,N_979,N_3141);
and U6641 (N_6641,N_72,N_585);
xnor U6642 (N_6642,N_3583,N_1018);
or U6643 (N_6643,N_4003,N_3533);
and U6644 (N_6644,N_4796,N_4746);
xnor U6645 (N_6645,N_189,N_2959);
xor U6646 (N_6646,N_2542,N_1971);
and U6647 (N_6647,N_2057,N_2321);
or U6648 (N_6648,N_3411,N_569);
nand U6649 (N_6649,N_3987,N_4186);
nor U6650 (N_6650,N_298,N_493);
and U6651 (N_6651,N_2727,N_3601);
and U6652 (N_6652,N_4787,N_916);
nand U6653 (N_6653,N_990,N_4751);
nand U6654 (N_6654,N_2047,N_3362);
nor U6655 (N_6655,N_2243,N_1549);
and U6656 (N_6656,N_1399,N_417);
or U6657 (N_6657,N_4881,N_2622);
and U6658 (N_6658,N_4397,N_3238);
or U6659 (N_6659,N_1227,N_297);
nor U6660 (N_6660,N_1267,N_122);
or U6661 (N_6661,N_3889,N_2684);
and U6662 (N_6662,N_2294,N_3104);
nand U6663 (N_6663,N_1374,N_1505);
nand U6664 (N_6664,N_4158,N_783);
xor U6665 (N_6665,N_3975,N_3020);
xnor U6666 (N_6666,N_4825,N_1153);
nand U6667 (N_6667,N_1705,N_325);
and U6668 (N_6668,N_4091,N_4689);
or U6669 (N_6669,N_178,N_3490);
xnor U6670 (N_6670,N_1470,N_3299);
xnor U6671 (N_6671,N_651,N_2516);
and U6672 (N_6672,N_4855,N_4265);
or U6673 (N_6673,N_2748,N_2822);
xor U6674 (N_6674,N_2990,N_2364);
nand U6675 (N_6675,N_1564,N_1268);
xnor U6676 (N_6676,N_1831,N_2996);
nand U6677 (N_6677,N_2408,N_184);
nor U6678 (N_6678,N_858,N_4422);
and U6679 (N_6679,N_4878,N_2491);
or U6680 (N_6680,N_4075,N_1951);
or U6681 (N_6681,N_3933,N_4783);
xnor U6682 (N_6682,N_4166,N_2882);
or U6683 (N_6683,N_4276,N_504);
nor U6684 (N_6684,N_4451,N_3314);
or U6685 (N_6685,N_4625,N_2770);
nand U6686 (N_6686,N_822,N_3312);
xor U6687 (N_6687,N_1574,N_1314);
nor U6688 (N_6688,N_1033,N_1994);
nand U6689 (N_6689,N_4317,N_2602);
xnor U6690 (N_6690,N_152,N_4877);
and U6691 (N_6691,N_1346,N_2846);
nand U6692 (N_6692,N_1147,N_1860);
xnor U6693 (N_6693,N_274,N_1916);
and U6694 (N_6694,N_4370,N_1920);
or U6695 (N_6695,N_208,N_4051);
or U6696 (N_6696,N_986,N_811);
nor U6697 (N_6697,N_4092,N_472);
nand U6698 (N_6698,N_3350,N_4856);
xor U6699 (N_6699,N_1284,N_4979);
xnor U6700 (N_6700,N_2873,N_3402);
xnor U6701 (N_6701,N_20,N_2853);
or U6702 (N_6702,N_1495,N_2471);
nand U6703 (N_6703,N_3733,N_4179);
or U6704 (N_6704,N_4200,N_4399);
or U6705 (N_6705,N_4792,N_2435);
and U6706 (N_6706,N_4190,N_4454);
or U6707 (N_6707,N_3287,N_3669);
xor U6708 (N_6708,N_4378,N_309);
and U6709 (N_6709,N_672,N_3408);
xnor U6710 (N_6710,N_2713,N_115);
and U6711 (N_6711,N_3265,N_2616);
and U6712 (N_6712,N_1051,N_4921);
or U6713 (N_6713,N_3320,N_3372);
xnor U6714 (N_6714,N_2923,N_3321);
or U6715 (N_6715,N_2373,N_1156);
xnor U6716 (N_6716,N_929,N_3160);
or U6717 (N_6717,N_931,N_3519);
nand U6718 (N_6718,N_640,N_1747);
nor U6719 (N_6719,N_3439,N_2811);
xor U6720 (N_6720,N_616,N_1613);
and U6721 (N_6721,N_3253,N_2332);
nor U6722 (N_6722,N_2198,N_2207);
nand U6723 (N_6723,N_385,N_252);
xnor U6724 (N_6724,N_4348,N_1096);
or U6725 (N_6725,N_2406,N_1995);
nand U6726 (N_6726,N_3564,N_4615);
and U6727 (N_6727,N_3576,N_2369);
or U6728 (N_6728,N_4867,N_2322);
xnor U6729 (N_6729,N_3010,N_1120);
nor U6730 (N_6730,N_3811,N_3945);
and U6731 (N_6731,N_1044,N_1046);
and U6732 (N_6732,N_2568,N_3937);
nand U6733 (N_6733,N_4119,N_4309);
xor U6734 (N_6734,N_1255,N_4982);
nand U6735 (N_6735,N_3866,N_2037);
nor U6736 (N_6736,N_1210,N_824);
nand U6737 (N_6737,N_4622,N_1233);
nand U6738 (N_6738,N_3897,N_4822);
nand U6739 (N_6739,N_995,N_2423);
xnor U6740 (N_6740,N_1963,N_4854);
or U6741 (N_6741,N_607,N_4834);
nor U6742 (N_6742,N_4008,N_909);
nor U6743 (N_6743,N_2851,N_2593);
nor U6744 (N_6744,N_2772,N_2500);
xnor U6745 (N_6745,N_3347,N_4912);
xnor U6746 (N_6746,N_501,N_2397);
and U6747 (N_6747,N_4904,N_3171);
and U6748 (N_6748,N_2547,N_1494);
or U6749 (N_6749,N_2042,N_2421);
or U6750 (N_6750,N_2221,N_4805);
and U6751 (N_6751,N_3901,N_2039);
xnor U6752 (N_6752,N_1754,N_1773);
and U6753 (N_6753,N_970,N_2913);
nor U6754 (N_6754,N_1324,N_3703);
and U6755 (N_6755,N_1151,N_1941);
and U6756 (N_6756,N_4021,N_3008);
nand U6757 (N_6757,N_3332,N_16);
xnor U6758 (N_6758,N_1356,N_2856);
or U6759 (N_6759,N_1601,N_687);
and U6760 (N_6760,N_146,N_317);
xor U6761 (N_6761,N_3622,N_2895);
xor U6762 (N_6762,N_80,N_785);
nor U6763 (N_6763,N_1493,N_4524);
nand U6764 (N_6764,N_1739,N_2961);
nor U6765 (N_6765,N_3476,N_1557);
and U6766 (N_6766,N_1160,N_1251);
nand U6767 (N_6767,N_2885,N_4033);
or U6768 (N_6768,N_2535,N_2504);
nor U6769 (N_6769,N_4785,N_1367);
and U6770 (N_6770,N_4550,N_1642);
nand U6771 (N_6771,N_2064,N_1632);
nor U6772 (N_6772,N_3167,N_2150);
or U6773 (N_6773,N_3235,N_2927);
nor U6774 (N_6774,N_4009,N_2954);
or U6775 (N_6775,N_3736,N_3510);
nand U6776 (N_6776,N_885,N_2336);
nand U6777 (N_6777,N_1856,N_3922);
and U6778 (N_6778,N_2017,N_898);
xnor U6779 (N_6779,N_1183,N_4140);
xnor U6780 (N_6780,N_256,N_3686);
or U6781 (N_6781,N_1427,N_3342);
or U6782 (N_6782,N_1055,N_2785);
nor U6783 (N_6783,N_1857,N_2848);
or U6784 (N_6784,N_4656,N_4168);
and U6785 (N_6785,N_3854,N_4605);
and U6786 (N_6786,N_1698,N_4765);
nand U6787 (N_6787,N_2426,N_35);
and U6788 (N_6788,N_2149,N_2531);
xnor U6789 (N_6789,N_2507,N_1458);
nor U6790 (N_6790,N_4243,N_3345);
or U6791 (N_6791,N_3497,N_429);
nor U6792 (N_6792,N_2754,N_1890);
nor U6793 (N_6793,N_3317,N_3306);
nand U6794 (N_6794,N_2673,N_2261);
nor U6795 (N_6795,N_3543,N_3215);
nor U6796 (N_6796,N_1627,N_244);
or U6797 (N_6797,N_2608,N_4069);
or U6798 (N_6798,N_416,N_4299);
xnor U6799 (N_6799,N_3282,N_474);
and U6800 (N_6800,N_2756,N_4869);
nand U6801 (N_6801,N_1053,N_2519);
and U6802 (N_6802,N_4172,N_910);
and U6803 (N_6803,N_4002,N_1084);
and U6804 (N_6804,N_3734,N_4228);
nand U6805 (N_6805,N_3667,N_4662);
or U6806 (N_6806,N_4063,N_2131);
or U6807 (N_6807,N_466,N_3397);
xnor U6808 (N_6808,N_4318,N_1205);
nand U6809 (N_6809,N_455,N_3643);
xnor U6810 (N_6810,N_3398,N_4436);
and U6811 (N_6811,N_1394,N_1732);
or U6812 (N_6812,N_2152,N_2527);
or U6813 (N_6813,N_1577,N_4111);
nor U6814 (N_6814,N_4586,N_2677);
nor U6815 (N_6815,N_2560,N_4287);
nand U6816 (N_6816,N_3995,N_1543);
or U6817 (N_6817,N_3286,N_1900);
nor U6818 (N_6818,N_3068,N_983);
and U6819 (N_6819,N_3297,N_2926);
xnor U6820 (N_6820,N_2097,N_3959);
or U6821 (N_6821,N_2341,N_1944);
nand U6822 (N_6822,N_4948,N_4752);
xnor U6823 (N_6823,N_2835,N_4290);
xnor U6824 (N_6824,N_1610,N_3190);
nor U6825 (N_6825,N_2263,N_789);
nor U6826 (N_6826,N_1223,N_753);
and U6827 (N_6827,N_617,N_1144);
nand U6828 (N_6828,N_4170,N_12);
nand U6829 (N_6829,N_2610,N_927);
xnor U6830 (N_6830,N_964,N_543);
and U6831 (N_6831,N_1979,N_1866);
xor U6832 (N_6832,N_1805,N_3832);
nor U6833 (N_6833,N_3831,N_945);
and U6834 (N_6834,N_1730,N_4274);
nand U6835 (N_6835,N_3142,N_3554);
and U6836 (N_6836,N_4523,N_3873);
xnor U6837 (N_6837,N_1685,N_2827);
xor U6838 (N_6838,N_1507,N_461);
and U6839 (N_6839,N_1874,N_1000);
nor U6840 (N_6840,N_2072,N_1855);
and U6841 (N_6841,N_4735,N_2718);
and U6842 (N_6842,N_2510,N_4053);
nand U6843 (N_6843,N_2937,N_993);
and U6844 (N_6844,N_667,N_2109);
xnor U6845 (N_6845,N_4423,N_4447);
xor U6846 (N_6846,N_2381,N_4232);
xor U6847 (N_6847,N_2112,N_292);
nor U6848 (N_6848,N_4277,N_3183);
nor U6849 (N_6849,N_1396,N_4146);
xor U6850 (N_6850,N_3383,N_1929);
xor U6851 (N_6851,N_4978,N_2134);
nor U6852 (N_6852,N_4913,N_4723);
nor U6853 (N_6853,N_2951,N_2385);
nand U6854 (N_6854,N_3363,N_541);
nand U6855 (N_6855,N_3595,N_469);
xor U6856 (N_6856,N_4742,N_1157);
nand U6857 (N_6857,N_1562,N_2652);
nand U6858 (N_6858,N_975,N_3965);
xnor U6859 (N_6859,N_1841,N_352);
nor U6860 (N_6860,N_960,N_3415);
nand U6861 (N_6861,N_2118,N_1607);
nand U6862 (N_6862,N_1656,N_4500);
nand U6863 (N_6863,N_3773,N_1638);
xnor U6864 (N_6864,N_1487,N_2395);
xor U6865 (N_6865,N_2354,N_2722);
nand U6866 (N_6866,N_4152,N_1242);
xnor U6867 (N_6867,N_2583,N_845);
and U6868 (N_6868,N_2934,N_4788);
nand U6869 (N_6869,N_2601,N_3872);
nor U6870 (N_6870,N_2363,N_2419);
nand U6871 (N_6871,N_2760,N_4245);
xnor U6872 (N_6872,N_1735,N_514);
and U6873 (N_6873,N_4435,N_3974);
and U6874 (N_6874,N_1109,N_4851);
or U6875 (N_6875,N_76,N_3625);
nor U6876 (N_6876,N_2615,N_1530);
xor U6877 (N_6877,N_1942,N_305);
nor U6878 (N_6878,N_510,N_792);
nand U6879 (N_6879,N_3127,N_199);
xor U6880 (N_6880,N_4576,N_410);
nand U6881 (N_6881,N_4712,N_1080);
nand U6882 (N_6882,N_1312,N_10);
or U6883 (N_6883,N_1195,N_3202);
and U6884 (N_6884,N_3137,N_246);
and U6885 (N_6885,N_2115,N_3760);
nand U6886 (N_6886,N_320,N_3001);
and U6887 (N_6887,N_3943,N_482);
or U6888 (N_6888,N_3620,N_1007);
or U6889 (N_6889,N_3025,N_4340);
nand U6890 (N_6890,N_1354,N_3539);
and U6891 (N_6891,N_1692,N_1066);
and U6892 (N_6892,N_393,N_3348);
or U6893 (N_6893,N_2701,N_4203);
nor U6894 (N_6894,N_739,N_1934);
xnor U6895 (N_6895,N_60,N_2900);
or U6896 (N_6896,N_4899,N_3384);
nor U6897 (N_6897,N_2697,N_2494);
nand U6898 (N_6898,N_4387,N_4903);
nor U6899 (N_6899,N_4574,N_4809);
nand U6900 (N_6900,N_4709,N_2914);
and U6901 (N_6901,N_2946,N_512);
nor U6902 (N_6902,N_4527,N_1614);
nand U6903 (N_6903,N_4585,N_3088);
and U6904 (N_6904,N_1677,N_2834);
xor U6905 (N_6905,N_4492,N_2357);
and U6906 (N_6906,N_4336,N_42);
or U6907 (N_6907,N_2477,N_3673);
xor U6908 (N_6908,N_1489,N_2871);
nor U6909 (N_6909,N_1746,N_2235);
nand U6910 (N_6910,N_51,N_3291);
xor U6911 (N_6911,N_2795,N_738);
nand U6912 (N_6912,N_3450,N_730);
xor U6913 (N_6913,N_2600,N_4058);
and U6914 (N_6914,N_1193,N_4181);
or U6915 (N_6915,N_4210,N_1706);
nor U6916 (N_6916,N_1669,N_2073);
xor U6917 (N_6917,N_4807,N_1641);
xnor U6918 (N_6918,N_994,N_1463);
and U6919 (N_6919,N_2392,N_572);
xnor U6920 (N_6920,N_1884,N_1363);
or U6921 (N_6921,N_53,N_2911);
nand U6922 (N_6922,N_498,N_3172);
or U6923 (N_6923,N_17,N_3883);
nor U6924 (N_6924,N_998,N_820);
or U6925 (N_6925,N_2427,N_2505);
xnor U6926 (N_6926,N_4337,N_4597);
or U6927 (N_6927,N_3335,N_1281);
nand U6928 (N_6928,N_230,N_1777);
or U6929 (N_6929,N_4951,N_2351);
nand U6930 (N_6930,N_2111,N_3678);
and U6931 (N_6931,N_3002,N_4678);
nor U6932 (N_6932,N_1152,N_4808);
xnor U6933 (N_6933,N_4273,N_2100);
nor U6934 (N_6934,N_3587,N_2056);
or U6935 (N_6935,N_3438,N_1445);
nor U6936 (N_6936,N_1303,N_368);
and U6937 (N_6937,N_446,N_4323);
and U6938 (N_6938,N_2849,N_1417);
nand U6939 (N_6939,N_3361,N_2729);
xor U6940 (N_6940,N_3429,N_4260);
xor U6941 (N_6941,N_254,N_547);
or U6942 (N_6942,N_2744,N_3503);
nand U6943 (N_6943,N_773,N_3927);
nor U6944 (N_6944,N_992,N_844);
nand U6945 (N_6945,N_3128,N_3632);
nor U6946 (N_6946,N_125,N_1711);
and U6947 (N_6947,N_4917,N_318);
nand U6948 (N_6948,N_1977,N_4647);
xor U6949 (N_6949,N_4133,N_3990);
and U6950 (N_6950,N_2699,N_544);
nor U6951 (N_6951,N_3798,N_732);
nand U6952 (N_6952,N_3326,N_4976);
nand U6953 (N_6953,N_4375,N_3700);
and U6954 (N_6954,N_4841,N_2638);
xor U6955 (N_6955,N_2328,N_1596);
nand U6956 (N_6956,N_3197,N_3952);
or U6957 (N_6957,N_4116,N_1716);
and U6958 (N_6958,N_14,N_365);
nand U6959 (N_6959,N_1861,N_3636);
nor U6960 (N_6960,N_260,N_2088);
and U6961 (N_6961,N_3500,N_1031);
and U6962 (N_6962,N_1030,N_1125);
xor U6963 (N_6963,N_614,N_88);
nand U6964 (N_6964,N_3823,N_4981);
xnor U6965 (N_6965,N_825,N_1554);
and U6966 (N_6966,N_3527,N_864);
nand U6967 (N_6967,N_4278,N_1386);
nand U6968 (N_6968,N_1076,N_4993);
or U6969 (N_6969,N_1260,N_3895);
and U6970 (N_6970,N_238,N_1155);
and U6971 (N_6971,N_1682,N_2906);
nor U6972 (N_6972,N_1361,N_1707);
nand U6973 (N_6973,N_608,N_3029);
or U6974 (N_6974,N_2649,N_1660);
or U6975 (N_6975,N_2128,N_972);
or U6976 (N_6976,N_82,N_3252);
nand U6977 (N_6977,N_1635,N_4114);
nor U6978 (N_6978,N_2140,N_3785);
nand U6979 (N_6979,N_2227,N_1670);
nand U6980 (N_6980,N_715,N_4262);
nor U6981 (N_6981,N_4420,N_4188);
nand U6982 (N_6982,N_4562,N_1296);
nand U6983 (N_6983,N_1736,N_1658);
xnor U6984 (N_6984,N_2833,N_2669);
and U6985 (N_6985,N_3841,N_3399);
xnor U6986 (N_6986,N_4380,N_4115);
and U6987 (N_6987,N_4673,N_2915);
xor U6988 (N_6988,N_165,N_251);
nor U6989 (N_6989,N_623,N_3346);
or U6990 (N_6990,N_4483,N_4959);
and U6991 (N_6991,N_2942,N_2627);
or U6992 (N_6992,N_912,N_1093);
or U6993 (N_6993,N_4701,N_4551);
and U6994 (N_6994,N_2522,N_2038);
xnor U6995 (N_6995,N_2466,N_497);
nand U6996 (N_6996,N_2145,N_2217);
or U6997 (N_6997,N_2912,N_2432);
xnor U6998 (N_6998,N_449,N_1216);
and U6999 (N_6999,N_2366,N_4939);
nor U7000 (N_7000,N_3437,N_3801);
nand U7001 (N_7001,N_698,N_1905);
or U7002 (N_7002,N_4359,N_956);
xor U7003 (N_7003,N_4564,N_4135);
nor U7004 (N_7004,N_2993,N_4230);
nor U7005 (N_7005,N_2051,N_4268);
and U7006 (N_7006,N_3981,N_1636);
xnor U7007 (N_7007,N_1101,N_2798);
xor U7008 (N_7008,N_3531,N_1659);
xnor U7009 (N_7009,N_4372,N_1617);
and U7010 (N_7010,N_1703,N_1447);
xor U7011 (N_7011,N_2933,N_1633);
xor U7012 (N_7012,N_1593,N_3698);
or U7013 (N_7013,N_4445,N_1608);
or U7014 (N_7014,N_56,N_2025);
nor U7015 (N_7015,N_3989,N_3150);
nand U7016 (N_7016,N_2262,N_1824);
or U7017 (N_7017,N_3982,N_1398);
or U7018 (N_7018,N_240,N_2393);
or U7019 (N_7019,N_2014,N_610);
and U7020 (N_7020,N_221,N_2859);
nor U7021 (N_7021,N_3881,N_2908);
nor U7022 (N_7022,N_3563,N_4410);
or U7023 (N_7023,N_1012,N_2394);
xnor U7024 (N_7024,N_4740,N_2490);
nand U7025 (N_7025,N_835,N_1646);
and U7026 (N_7026,N_713,N_2479);
nor U7027 (N_7027,N_3207,N_2256);
and U7028 (N_7028,N_897,N_4543);
xnor U7029 (N_7029,N_3863,N_3537);
xnor U7030 (N_7030,N_4178,N_2182);
xor U7031 (N_7031,N_2436,N_3715);
or U7032 (N_7032,N_4129,N_300);
or U7033 (N_7033,N_350,N_148);
or U7034 (N_7034,N_4249,N_1888);
nor U7035 (N_7035,N_4350,N_1146);
and U7036 (N_7036,N_4421,N_4614);
nand U7037 (N_7037,N_4107,N_3521);
or U7038 (N_7038,N_4588,N_3938);
and U7039 (N_7039,N_3006,N_2044);
nand U7040 (N_7040,N_4896,N_1912);
nand U7041 (N_7041,N_627,N_123);
nor U7042 (N_7042,N_1009,N_3752);
xnor U7043 (N_7043,N_1804,N_1426);
nand U7044 (N_7044,N_1762,N_4015);
or U7045 (N_7045,N_361,N_982);
and U7046 (N_7046,N_802,N_4185);
or U7047 (N_7047,N_1753,N_453);
xnor U7048 (N_7048,N_2242,N_1116);
and U7049 (N_7049,N_635,N_3896);
nor U7050 (N_7050,N_3054,N_3979);
xor U7051 (N_7051,N_1775,N_2273);
xor U7052 (N_7052,N_875,N_869);
xnor U7053 (N_7053,N_4773,N_4215);
and U7054 (N_7054,N_4955,N_206);
nor U7055 (N_7055,N_2289,N_1360);
and U7056 (N_7056,N_2138,N_2758);
nand U7057 (N_7057,N_1745,N_4251);
nor U7058 (N_7058,N_4099,N_3498);
xor U7059 (N_7059,N_2511,N_3567);
xnor U7060 (N_7060,N_790,N_3842);
and U7061 (N_7061,N_2508,N_3496);
xnor U7062 (N_7062,N_2246,N_1318);
and U7063 (N_7063,N_2308,N_3344);
nor U7064 (N_7064,N_2082,N_2585);
and U7065 (N_7065,N_1529,N_1112);
nor U7066 (N_7066,N_4762,N_1202);
nand U7067 (N_7067,N_915,N_2628);
nor U7068 (N_7068,N_2513,N_1429);
nor U7069 (N_7069,N_4294,N_1878);
or U7070 (N_7070,N_2302,N_2966);
or U7071 (N_7071,N_2260,N_1766);
or U7072 (N_7072,N_40,N_1761);
nor U7073 (N_7073,N_3168,N_4295);
nand U7074 (N_7074,N_4440,N_4338);
nor U7075 (N_7075,N_4266,N_2590);
xor U7076 (N_7076,N_4697,N_1213);
or U7077 (N_7077,N_4314,N_980);
or U7078 (N_7078,N_1275,N_2474);
or U7079 (N_7079,N_112,N_2125);
nand U7080 (N_7080,N_3612,N_147);
and U7081 (N_7081,N_161,N_4386);
or U7082 (N_7082,N_1668,N_4770);
nor U7083 (N_7083,N_4900,N_767);
nor U7084 (N_7084,N_1958,N_4246);
xnor U7085 (N_7085,N_4529,N_193);
nor U7086 (N_7086,N_2776,N_1679);
and U7087 (N_7087,N_3584,N_3407);
nor U7088 (N_7088,N_2345,N_3180);
nor U7089 (N_7089,N_4250,N_1914);
xnor U7090 (N_7090,N_737,N_595);
nand U7091 (N_7091,N_1486,N_3462);
xor U7092 (N_7092,N_258,N_4088);
and U7093 (N_7093,N_3033,N_3573);
xnor U7094 (N_7094,N_1477,N_4282);
nand U7095 (N_7095,N_288,N_4630);
nor U7096 (N_7096,N_4213,N_4049);
and U7097 (N_7097,N_4217,N_2272);
nand U7098 (N_7098,N_1186,N_2055);
or U7099 (N_7099,N_1343,N_3921);
and U7100 (N_7100,N_1340,N_2828);
or U7101 (N_7101,N_3443,N_4655);
or U7102 (N_7102,N_733,N_2562);
nor U7103 (N_7103,N_1070,N_1313);
nand U7104 (N_7104,N_1234,N_1441);
xnor U7105 (N_7105,N_2285,N_1978);
nand U7106 (N_7106,N_3444,N_2894);
or U7107 (N_7107,N_399,N_4836);
and U7108 (N_7108,N_2443,N_4537);
nor U7109 (N_7109,N_592,N_3494);
nor U7110 (N_7110,N_4821,N_3735);
nor U7111 (N_7111,N_721,N_3023);
nand U7112 (N_7112,N_4199,N_1113);
nor U7113 (N_7113,N_3878,N_18);
nor U7114 (N_7114,N_774,N_1571);
nand U7115 (N_7115,N_2854,N_2813);
nor U7116 (N_7116,N_605,N_1167);
xnor U7117 (N_7117,N_3166,N_2566);
nor U7118 (N_7118,N_3290,N_1666);
and U7119 (N_7119,N_2193,N_868);
nor U7120 (N_7120,N_3561,N_2646);
and U7121 (N_7121,N_3705,N_3266);
nor U7122 (N_7122,N_3098,N_487);
xor U7123 (N_7123,N_118,N_4635);
nor U7124 (N_7124,N_181,N_3688);
nand U7125 (N_7125,N_1868,N_2470);
or U7126 (N_7126,N_3702,N_899);
nor U7127 (N_7127,N_1850,N_4661);
xnor U7128 (N_7128,N_1287,N_3057);
nor U7129 (N_7129,N_4990,N_2201);
nor U7130 (N_7130,N_840,N_1797);
and U7131 (N_7131,N_367,N_1695);
or U7132 (N_7132,N_3260,N_150);
nor U7133 (N_7133,N_596,N_4326);
xor U7134 (N_7134,N_2163,N_2475);
xnor U7135 (N_7135,N_2171,N_2018);
and U7136 (N_7136,N_4433,N_4972);
xor U7137 (N_7137,N_619,N_4064);
and U7138 (N_7138,N_571,N_154);
xnor U7139 (N_7139,N_4710,N_1348);
xnor U7140 (N_7140,N_594,N_1969);
and U7141 (N_7141,N_1809,N_3807);
nand U7142 (N_7142,N_2909,N_530);
nand U7143 (N_7143,N_3594,N_4157);
and U7144 (N_7144,N_2232,N_1961);
nor U7145 (N_7145,N_3236,N_4986);
or U7146 (N_7146,N_3433,N_1150);
or U7147 (N_7147,N_4073,N_1867);
xnor U7148 (N_7148,N_421,N_1932);
or U7149 (N_7149,N_750,N_2040);
nand U7150 (N_7150,N_4816,N_2160);
xnor U7151 (N_7151,N_4980,N_420);
nand U7152 (N_7152,N_183,N_4928);
nor U7153 (N_7153,N_3522,N_2238);
nor U7154 (N_7154,N_1816,N_1606);
nand U7155 (N_7155,N_255,N_3015);
nand U7156 (N_7156,N_313,N_4169);
nand U7157 (N_7157,N_2955,N_3046);
and U7158 (N_7158,N_2206,N_4);
xnor U7159 (N_7159,N_1528,N_226);
xor U7160 (N_7160,N_2641,N_351);
or U7161 (N_7161,N_158,N_4627);
xor U7162 (N_7162,N_4054,N_2502);
nand U7163 (N_7163,N_65,N_3548);
nor U7164 (N_7164,N_3613,N_2875);
xor U7165 (N_7165,N_3090,N_1039);
or U7166 (N_7166,N_2824,N_3065);
and U7167 (N_7167,N_468,N_3270);
xor U7168 (N_7168,N_3864,N_1368);
nor U7169 (N_7169,N_4067,N_4953);
and U7170 (N_7170,N_3177,N_4522);
nor U7171 (N_7171,N_3868,N_1069);
xor U7172 (N_7172,N_908,N_930);
and U7173 (N_7173,N_2191,N_1810);
and U7174 (N_7174,N_167,N_4672);
or U7175 (N_7175,N_4609,N_3379);
nor U7176 (N_7176,N_109,N_198);
or U7177 (N_7177,N_3635,N_4031);
or U7178 (N_7178,N_2825,N_1380);
xnor U7179 (N_7179,N_1694,N_731);
xnor U7180 (N_7180,N_1812,N_2065);
xnor U7181 (N_7181,N_4649,N_1847);
nand U7182 (N_7182,N_1973,N_143);
nand U7183 (N_7183,N_727,N_2030);
or U7184 (N_7184,N_3436,N_1541);
or U7185 (N_7185,N_413,N_1060);
and U7186 (N_7186,N_22,N_2579);
nor U7187 (N_7187,N_2623,N_2580);
xor U7188 (N_7188,N_601,N_3395);
xnor U7189 (N_7189,N_388,N_4478);
or U7190 (N_7190,N_4863,N_4639);
and U7191 (N_7191,N_4113,N_418);
or U7192 (N_7192,N_403,N_4870);
or U7193 (N_7193,N_3463,N_3334);
and U7194 (N_7194,N_4671,N_3827);
nand U7195 (N_7195,N_1491,N_4292);
and U7196 (N_7196,N_4802,N_2779);
xnor U7197 (N_7197,N_4590,N_3184);
nand U7198 (N_7198,N_1191,N_4240);
nand U7199 (N_7199,N_1697,N_3032);
xnor U7200 (N_7200,N_2379,N_3011);
nor U7201 (N_7201,N_3159,N_291);
nor U7202 (N_7202,N_2879,N_2596);
nor U7203 (N_7203,N_1057,N_681);
and U7204 (N_7204,N_454,N_2129);
xnor U7205 (N_7205,N_2070,N_4909);
xnor U7206 (N_7206,N_2174,N_3855);
xnor U7207 (N_7207,N_3019,N_4559);
nor U7208 (N_7208,N_2372,N_4502);
nand U7209 (N_7209,N_860,N_2469);
xor U7210 (N_7210,N_3113,N_1438);
and U7211 (N_7211,N_1504,N_2417);
nor U7212 (N_7212,N_3116,N_1517);
xor U7213 (N_7213,N_3692,N_4023);
nand U7214 (N_7214,N_3996,N_685);
or U7215 (N_7215,N_3489,N_4732);
or U7216 (N_7216,N_3867,N_105);
nor U7217 (N_7217,N_1559,N_4910);
or U7218 (N_7218,N_1457,N_1651);
and U7219 (N_7219,N_372,N_2156);
nor U7220 (N_7220,N_201,N_2080);
or U7221 (N_7221,N_772,N_2059);
and U7222 (N_7222,N_933,N_1148);
xor U7223 (N_7223,N_2439,N_83);
nand U7224 (N_7224,N_3784,N_94);
nand U7225 (N_7225,N_1170,N_911);
and U7226 (N_7226,N_2456,N_347);
xnor U7227 (N_7227,N_1580,N_4696);
or U7228 (N_7228,N_1726,N_1960);
and U7229 (N_7229,N_1674,N_129);
nor U7230 (N_7230,N_400,N_914);
nand U7231 (N_7231,N_3727,N_1132);
nand U7232 (N_7232,N_1649,N_190);
nor U7233 (N_7233,N_683,N_4547);
nand U7234 (N_7234,N_4072,N_293);
xnor U7235 (N_7235,N_2743,N_1741);
nand U7236 (N_7236,N_677,N_443);
nand U7237 (N_7237,N_4737,N_108);
xor U7238 (N_7238,N_680,N_2315);
and U7239 (N_7239,N_4988,N_1058);
nand U7240 (N_7240,N_4000,N_815);
or U7241 (N_7241,N_3857,N_247);
or U7242 (N_7242,N_3556,N_1565);
and U7243 (N_7243,N_3469,N_1311);
and U7244 (N_7244,N_1049,N_3888);
and U7245 (N_7245,N_4507,N_422);
or U7246 (N_7246,N_952,N_600);
nor U7247 (N_7247,N_3958,N_4027);
and U7248 (N_7248,N_1630,N_4760);
nor U7249 (N_7249,N_4048,N_1025);
xor U7250 (N_7250,N_3787,N_1826);
and U7251 (N_7251,N_488,N_2248);
xnor U7252 (N_7252,N_3013,N_4165);
nor U7253 (N_7253,N_1581,N_4757);
nor U7254 (N_7254,N_1843,N_28);
nor U7255 (N_7255,N_144,N_793);
and U7256 (N_7256,N_1045,N_4010);
xnor U7257 (N_7257,N_1858,N_2383);
or U7258 (N_7258,N_691,N_4563);
xnor U7259 (N_7259,N_4442,N_1616);
nor U7260 (N_7260,N_2425,N_1250);
xor U7261 (N_7261,N_1204,N_2016);
or U7262 (N_7262,N_4515,N_4396);
or U7263 (N_7263,N_321,N_589);
nand U7264 (N_7264,N_976,N_3682);
xor U7265 (N_7265,N_1665,N_1681);
or U7266 (N_7266,N_2796,N_217);
and U7267 (N_7267,N_4094,N_4918);
xor U7268 (N_7268,N_1038,N_622);
nor U7269 (N_7269,N_467,N_1105);
or U7270 (N_7270,N_670,N_2405);
or U7271 (N_7271,N_3009,N_3203);
or U7272 (N_7272,N_4416,N_3243);
and U7273 (N_7273,N_4984,N_3178);
or U7274 (N_7274,N_3812,N_2558);
nand U7275 (N_7275,N_2692,N_4461);
nor U7276 (N_7276,N_499,N_362);
or U7277 (N_7277,N_606,N_2019);
and U7278 (N_7278,N_2573,N_3410);
or U7279 (N_7279,N_103,N_2493);
nand U7280 (N_7280,N_1450,N_4293);
nand U7281 (N_7281,N_4096,N_4688);
nor U7282 (N_7282,N_1142,N_4638);
and U7283 (N_7283,N_4572,N_1453);
and U7284 (N_7284,N_1054,N_4351);
nand U7285 (N_7285,N_2609,N_629);
nor U7286 (N_7286,N_328,N_214);
nor U7287 (N_7287,N_1022,N_2634);
and U7288 (N_7288,N_1293,N_2924);
and U7289 (N_7289,N_3917,N_2237);
nand U7290 (N_7290,N_3191,N_2031);
and U7291 (N_7291,N_4261,N_2245);
and U7292 (N_7292,N_2253,N_2086);
xnor U7293 (N_7293,N_3200,N_3000);
or U7294 (N_7294,N_3250,N_1077);
nor U7295 (N_7295,N_3547,N_2349);
or U7296 (N_7296,N_419,N_827);
xnor U7297 (N_7297,N_3096,N_3050);
or U7298 (N_7298,N_886,N_705);
or U7299 (N_7299,N_3021,N_1575);
and U7300 (N_7300,N_2945,N_2613);
or U7301 (N_7301,N_3569,N_3448);
or U7302 (N_7302,N_4382,N_719);
nor U7303 (N_7303,N_4509,N_2816);
xnor U7304 (N_7304,N_2569,N_628);
or U7305 (N_7305,N_4346,N_921);
xnor U7306 (N_7306,N_4193,N_3553);
and U7307 (N_7307,N_678,N_3204);
and U7308 (N_7308,N_3460,N_1442);
nand U7309 (N_7309,N_4668,N_209);
xnor U7310 (N_7310,N_2530,N_4312);
nor U7311 (N_7311,N_4469,N_2636);
or U7312 (N_7312,N_2303,N_1690);
or U7313 (N_7313,N_3182,N_3839);
and U7314 (N_7314,N_4861,N_2705);
nor U7315 (N_7315,N_1913,N_535);
nor U7316 (N_7316,N_4589,N_242);
and U7317 (N_7317,N_1483,N_2577);
and U7318 (N_7318,N_2274,N_384);
and U7319 (N_7319,N_310,N_1282);
xor U7320 (N_7320,N_3082,N_2555);
or U7321 (N_7321,N_2288,N_4654);
nand U7322 (N_7322,N_2151,N_3254);
or U7323 (N_7323,N_1280,N_1539);
nand U7324 (N_7324,N_4600,N_3670);
or U7325 (N_7325,N_2172,N_4161);
nand U7326 (N_7326,N_2786,N_4874);
xor U7327 (N_7327,N_2574,N_2107);
or U7328 (N_7328,N_2096,N_1230);
nand U7329 (N_7329,N_3157,N_59);
and U7330 (N_7330,N_435,N_55);
xor U7331 (N_7331,N_4384,N_4286);
nor U7332 (N_7332,N_1619,N_1620);
or U7333 (N_7333,N_4280,N_4495);
xnor U7334 (N_7334,N_2011,N_2076);
or U7335 (N_7335,N_859,N_4707);
nand U7336 (N_7336,N_3618,N_6);
xor U7337 (N_7337,N_3423,N_2739);
xor U7338 (N_7338,N_3511,N_3111);
nand U7339 (N_7339,N_3871,N_408);
and U7340 (N_7340,N_4943,N_2536);
nand U7341 (N_7341,N_4579,N_2904);
nor U7342 (N_7342,N_4209,N_3080);
and U7343 (N_7343,N_2552,N_1582);
nand U7344 (N_7344,N_890,N_4377);
nand U7345 (N_7345,N_1895,N_2314);
or U7346 (N_7346,N_2537,N_1865);
and U7347 (N_7347,N_1710,N_126);
xor U7348 (N_7348,N_3294,N_4095);
nor U7349 (N_7349,N_676,N_529);
nor U7350 (N_7350,N_1452,N_3284);
nand U7351 (N_7351,N_3566,N_344);
and U7352 (N_7352,N_1966,N_2215);
or U7353 (N_7353,N_4539,N_323);
nor U7354 (N_7354,N_1059,N_2250);
or U7355 (N_7355,N_1622,N_3523);
xor U7356 (N_7356,N_2781,N_484);
and U7357 (N_7357,N_4339,N_1422);
and U7358 (N_7358,N_3295,N_2063);
and U7359 (N_7359,N_1419,N_3234);
or U7360 (N_7360,N_3879,N_1563);
nor U7361 (N_7361,N_4204,N_3037);
nand U7362 (N_7362,N_4660,N_1859);
nand U7363 (N_7363,N_2497,N_3493);
or U7364 (N_7364,N_3470,N_2587);
nand U7365 (N_7365,N_3683,N_2985);
or U7366 (N_7366,N_839,N_1351);
or U7367 (N_7367,N_2844,N_4850);
or U7368 (N_7368,N_3740,N_4503);
nand U7369 (N_7369,N_81,N_1428);
nor U7370 (N_7370,N_4343,N_4134);
xor U7371 (N_7371,N_2401,N_4664);
xor U7372 (N_7372,N_284,N_412);
nor U7373 (N_7373,N_2465,N_3779);
or U7374 (N_7374,N_2903,N_2362);
xnor U7375 (N_7375,N_3359,N_1926);
xor U7376 (N_7376,N_4325,N_3961);
nand U7377 (N_7377,N_2091,N_2375);
xor U7378 (N_7378,N_4364,N_3464);
or U7379 (N_7379,N_776,N_1317);
or U7380 (N_7380,N_1019,N_1628);
or U7381 (N_7381,N_4642,N_2514);
nand U7382 (N_7382,N_1993,N_3222);
and U7383 (N_7383,N_4936,N_3414);
nand U7384 (N_7384,N_2948,N_2506);
nand U7385 (N_7385,N_1235,N_813);
nor U7386 (N_7386,N_2139,N_3721);
nand U7387 (N_7387,N_3123,N_611);
nor U7388 (N_7388,N_41,N_2778);
or U7389 (N_7389,N_270,N_2447);
or U7390 (N_7390,N_2295,N_1990);
xnor U7391 (N_7391,N_304,N_444);
and U7392 (N_7392,N_4223,N_4946);
and U7393 (N_7393,N_3151,N_4864);
or U7394 (N_7394,N_3188,N_3375);
or U7395 (N_7395,N_3762,N_2257);
nor U7396 (N_7396,N_1016,N_4750);
nor U7397 (N_7397,N_4035,N_4632);
nor U7398 (N_7398,N_1432,N_1806);
nand U7399 (N_7399,N_3910,N_797);
or U7400 (N_7400,N_3351,N_2296);
xnor U7401 (N_7401,N_4810,N_4400);
xnor U7402 (N_7402,N_3890,N_3356);
or U7403 (N_7403,N_2769,N_477);
or U7404 (N_7404,N_3546,N_213);
and U7405 (N_7405,N_2512,N_394);
nor U7406 (N_7406,N_3639,N_1436);
nand U7407 (N_7407,N_1423,N_4406);
nor U7408 (N_7408,N_145,N_4908);
nand U7409 (N_7409,N_464,N_1119);
or U7410 (N_7410,N_3403,N_4385);
nor U7411 (N_7411,N_1145,N_2212);
nand U7412 (N_7412,N_3992,N_2009);
or U7413 (N_7413,N_2194,N_3759);
or U7414 (N_7414,N_4611,N_4310);
and U7415 (N_7415,N_1813,N_3962);
nor U7416 (N_7416,N_3130,N_3330);
xnor U7417 (N_7417,N_1123,N_2266);
nand U7418 (N_7418,N_1782,N_4139);
or U7419 (N_7419,N_659,N_602);
and U7420 (N_7420,N_1957,N_1987);
and U7421 (N_7421,N_2968,N_646);
xor U7422 (N_7422,N_99,N_2008);
and U7423 (N_7423,N_842,N_1576);
nand U7424 (N_7424,N_200,N_2093);
or U7425 (N_7425,N_383,N_3277);
and U7426 (N_7426,N_2311,N_1218);
and U7427 (N_7427,N_3690,N_359);
nor U7428 (N_7428,N_861,N_1326);
nor U7429 (N_7429,N_2327,N_27);
or U7430 (N_7430,N_2185,N_2686);
xnor U7431 (N_7431,N_373,N_1301);
and U7432 (N_7432,N_967,N_2483);
or U7433 (N_7433,N_2496,N_4560);
and U7434 (N_7434,N_4452,N_740);
nand U7435 (N_7435,N_3472,N_3515);
xor U7436 (N_7436,N_4797,N_884);
and U7437 (N_7437,N_4763,N_3475);
xnor U7438 (N_7438,N_3074,N_4743);
nor U7439 (N_7439,N_851,N_4748);
xor U7440 (N_7440,N_4780,N_2690);
nand U7441 (N_7441,N_2715,N_4657);
nand U7442 (N_7442,N_1469,N_4845);
or U7443 (N_7443,N_4556,N_4411);
nand U7444 (N_7444,N_2997,N_4670);
nor U7445 (N_7445,N_2184,N_1885);
or U7446 (N_7446,N_643,N_1763);
nand U7447 (N_7447,N_1820,N_3717);
nor U7448 (N_7448,N_2355,N_15);
nand U7449 (N_7449,N_1793,N_4460);
and U7450 (N_7450,N_2644,N_3186);
xnor U7451 (N_7451,N_3585,N_2323);
xor U7452 (N_7452,N_4018,N_3225);
nand U7453 (N_7453,N_4505,N_29);
xnor U7454 (N_7454,N_203,N_3062);
nand U7455 (N_7455,N_4248,N_3488);
nand U7456 (N_7456,N_3906,N_4599);
and U7457 (N_7457,N_279,N_3093);
and U7458 (N_7458,N_1411,N_4391);
xnor U7459 (N_7459,N_456,N_1277);
nor U7460 (N_7460,N_3427,N_4532);
xor U7461 (N_7461,N_2843,N_4376);
or U7462 (N_7462,N_3208,N_3953);
or U7463 (N_7463,N_1061,N_1708);
nand U7464 (N_7464,N_3371,N_2386);
or U7465 (N_7465,N_3101,N_1792);
nand U7466 (N_7466,N_2711,N_4691);
or U7467 (N_7467,N_4330,N_4297);
xor U7468 (N_7468,N_2680,N_1936);
nand U7469 (N_7469,N_1323,N_4683);
xnor U7470 (N_7470,N_1107,N_2550);
nor U7471 (N_7471,N_3271,N_888);
xnor U7472 (N_7472,N_1814,N_1513);
xnor U7473 (N_7473,N_2689,N_1252);
nand U7474 (N_7474,N_4418,N_2850);
xor U7475 (N_7475,N_358,N_4234);
nand U7476 (N_7476,N_4862,N_3985);
and U7477 (N_7477,N_2720,N_2792);
and U7478 (N_7478,N_2805,N_4974);
or U7479 (N_7479,N_2054,N_4602);
xor U7480 (N_7480,N_1001,N_3073);
nor U7481 (N_7481,N_2950,N_4038);
nand U7482 (N_7482,N_1344,N_901);
nand U7483 (N_7483,N_1184,N_4006);
nor U7484 (N_7484,N_752,N_2678);
nand U7485 (N_7485,N_3646,N_593);
xnor U7486 (N_7486,N_2104,N_1893);
nand U7487 (N_7487,N_4231,N_3017);
xnor U7488 (N_7488,N_4879,N_3422);
nor U7489 (N_7489,N_4162,N_3999);
xor U7490 (N_7490,N_2765,N_4934);
nor U7491 (N_7491,N_2548,N_39);
nand U7492 (N_7492,N_3848,N_985);
nand U7493 (N_7493,N_4882,N_4931);
or U7494 (N_7494,N_892,N_1339);
xnor U7495 (N_7495,N_2124,N_4395);
xnor U7496 (N_7496,N_3477,N_2529);
or U7497 (N_7497,N_234,N_4137);
xnor U7498 (N_7498,N_2324,N_45);
nor U7499 (N_7499,N_4663,N_2325);
or U7500 (N_7500,N_366,N_433);
or U7501 (N_7501,N_143,N_3433);
nor U7502 (N_7502,N_4649,N_1768);
xor U7503 (N_7503,N_359,N_36);
nand U7504 (N_7504,N_2289,N_2480);
nor U7505 (N_7505,N_4209,N_265);
nor U7506 (N_7506,N_3891,N_1976);
or U7507 (N_7507,N_3529,N_4303);
xnor U7508 (N_7508,N_1070,N_2540);
xor U7509 (N_7509,N_4670,N_4843);
xnor U7510 (N_7510,N_3759,N_3193);
and U7511 (N_7511,N_2005,N_2239);
nor U7512 (N_7512,N_340,N_2279);
nor U7513 (N_7513,N_4257,N_2491);
nand U7514 (N_7514,N_3235,N_1769);
xor U7515 (N_7515,N_4995,N_1274);
and U7516 (N_7516,N_4831,N_4079);
nor U7517 (N_7517,N_2638,N_2585);
xor U7518 (N_7518,N_2756,N_1746);
xnor U7519 (N_7519,N_4225,N_4046);
and U7520 (N_7520,N_509,N_1341);
nand U7521 (N_7521,N_3771,N_1520);
and U7522 (N_7522,N_1508,N_791);
nand U7523 (N_7523,N_6,N_3778);
nor U7524 (N_7524,N_2188,N_3434);
or U7525 (N_7525,N_2878,N_322);
and U7526 (N_7526,N_1519,N_4906);
or U7527 (N_7527,N_1580,N_4731);
nand U7528 (N_7528,N_4083,N_4117);
nand U7529 (N_7529,N_4741,N_72);
xnor U7530 (N_7530,N_1818,N_3362);
or U7531 (N_7531,N_2897,N_2110);
nor U7532 (N_7532,N_75,N_1029);
and U7533 (N_7533,N_1877,N_2521);
xnor U7534 (N_7534,N_3811,N_3270);
nand U7535 (N_7535,N_3784,N_4835);
nor U7536 (N_7536,N_2659,N_1681);
nor U7537 (N_7537,N_4287,N_3258);
or U7538 (N_7538,N_4709,N_3040);
and U7539 (N_7539,N_1873,N_2864);
or U7540 (N_7540,N_1957,N_4830);
nor U7541 (N_7541,N_1214,N_3472);
nand U7542 (N_7542,N_3108,N_3824);
or U7543 (N_7543,N_3382,N_1441);
and U7544 (N_7544,N_3747,N_1663);
xor U7545 (N_7545,N_3831,N_1012);
nor U7546 (N_7546,N_3997,N_905);
or U7547 (N_7547,N_2905,N_1638);
or U7548 (N_7548,N_2239,N_2316);
and U7549 (N_7549,N_3347,N_1044);
or U7550 (N_7550,N_2846,N_4009);
nand U7551 (N_7551,N_1900,N_3786);
xnor U7552 (N_7552,N_1587,N_4750);
and U7553 (N_7553,N_2734,N_3923);
nand U7554 (N_7554,N_2880,N_4830);
nand U7555 (N_7555,N_1552,N_1489);
nor U7556 (N_7556,N_1130,N_1497);
xor U7557 (N_7557,N_3369,N_3765);
nand U7558 (N_7558,N_1710,N_1661);
and U7559 (N_7559,N_800,N_2703);
or U7560 (N_7560,N_1799,N_2818);
nand U7561 (N_7561,N_2457,N_1134);
nor U7562 (N_7562,N_3348,N_4301);
and U7563 (N_7563,N_635,N_1851);
nor U7564 (N_7564,N_2553,N_4009);
nand U7565 (N_7565,N_402,N_4484);
xnor U7566 (N_7566,N_3917,N_2416);
nand U7567 (N_7567,N_2948,N_2390);
nor U7568 (N_7568,N_1535,N_3768);
or U7569 (N_7569,N_4528,N_2250);
nor U7570 (N_7570,N_1171,N_4906);
or U7571 (N_7571,N_2851,N_567);
nand U7572 (N_7572,N_4900,N_4260);
or U7573 (N_7573,N_1921,N_3013);
or U7574 (N_7574,N_2108,N_4473);
nor U7575 (N_7575,N_4242,N_3325);
or U7576 (N_7576,N_521,N_3573);
nand U7577 (N_7577,N_2481,N_2966);
xnor U7578 (N_7578,N_786,N_3050);
or U7579 (N_7579,N_3942,N_2027);
xnor U7580 (N_7580,N_850,N_2716);
nand U7581 (N_7581,N_1854,N_1913);
and U7582 (N_7582,N_1149,N_1979);
or U7583 (N_7583,N_501,N_113);
or U7584 (N_7584,N_1649,N_4907);
xor U7585 (N_7585,N_4124,N_3419);
or U7586 (N_7586,N_1663,N_2902);
nor U7587 (N_7587,N_109,N_1854);
nor U7588 (N_7588,N_4583,N_2689);
xnor U7589 (N_7589,N_1484,N_4516);
and U7590 (N_7590,N_848,N_4176);
or U7591 (N_7591,N_3076,N_3467);
xor U7592 (N_7592,N_649,N_3705);
or U7593 (N_7593,N_3509,N_3385);
xor U7594 (N_7594,N_4176,N_3145);
nor U7595 (N_7595,N_2045,N_9);
nor U7596 (N_7596,N_1064,N_1628);
xnor U7597 (N_7597,N_1437,N_3419);
nand U7598 (N_7598,N_3250,N_3778);
and U7599 (N_7599,N_2572,N_3102);
nor U7600 (N_7600,N_2563,N_3270);
nor U7601 (N_7601,N_1473,N_4205);
nor U7602 (N_7602,N_884,N_3457);
nand U7603 (N_7603,N_1114,N_2993);
or U7604 (N_7604,N_2942,N_2036);
nor U7605 (N_7605,N_4341,N_4407);
or U7606 (N_7606,N_749,N_4014);
xor U7607 (N_7607,N_4856,N_4611);
or U7608 (N_7608,N_3339,N_4953);
nand U7609 (N_7609,N_3498,N_402);
xnor U7610 (N_7610,N_3600,N_3465);
nand U7611 (N_7611,N_509,N_4209);
or U7612 (N_7612,N_3893,N_2521);
or U7613 (N_7613,N_4969,N_2838);
or U7614 (N_7614,N_118,N_182);
xnor U7615 (N_7615,N_1437,N_4926);
nor U7616 (N_7616,N_1620,N_1246);
nand U7617 (N_7617,N_3186,N_4213);
xnor U7618 (N_7618,N_4483,N_4530);
or U7619 (N_7619,N_961,N_4804);
and U7620 (N_7620,N_1732,N_2915);
nand U7621 (N_7621,N_754,N_3676);
nand U7622 (N_7622,N_3437,N_1535);
nand U7623 (N_7623,N_2147,N_1755);
nand U7624 (N_7624,N_3657,N_4363);
nor U7625 (N_7625,N_1769,N_3986);
or U7626 (N_7626,N_4921,N_2926);
nor U7627 (N_7627,N_887,N_3628);
and U7628 (N_7628,N_768,N_73);
and U7629 (N_7629,N_4395,N_270);
or U7630 (N_7630,N_2682,N_2698);
nand U7631 (N_7631,N_3280,N_985);
or U7632 (N_7632,N_4152,N_3273);
or U7633 (N_7633,N_4768,N_3265);
xor U7634 (N_7634,N_3188,N_1501);
xnor U7635 (N_7635,N_2388,N_4844);
nand U7636 (N_7636,N_1756,N_619);
nand U7637 (N_7637,N_2179,N_1506);
and U7638 (N_7638,N_2980,N_3646);
or U7639 (N_7639,N_3023,N_3661);
and U7640 (N_7640,N_1065,N_3231);
xor U7641 (N_7641,N_1494,N_1217);
nor U7642 (N_7642,N_41,N_1221);
nor U7643 (N_7643,N_1653,N_1654);
xor U7644 (N_7644,N_3069,N_3753);
or U7645 (N_7645,N_204,N_3164);
xnor U7646 (N_7646,N_4723,N_1217);
nand U7647 (N_7647,N_1035,N_1911);
nand U7648 (N_7648,N_1555,N_935);
and U7649 (N_7649,N_1441,N_3378);
nor U7650 (N_7650,N_4616,N_2827);
or U7651 (N_7651,N_1983,N_2912);
nand U7652 (N_7652,N_3821,N_3621);
nand U7653 (N_7653,N_159,N_2522);
nand U7654 (N_7654,N_2404,N_3196);
nand U7655 (N_7655,N_4855,N_620);
xor U7656 (N_7656,N_3628,N_1901);
or U7657 (N_7657,N_990,N_4972);
nand U7658 (N_7658,N_1051,N_2740);
xor U7659 (N_7659,N_4354,N_165);
and U7660 (N_7660,N_2180,N_791);
xor U7661 (N_7661,N_2673,N_3893);
and U7662 (N_7662,N_4274,N_4717);
nor U7663 (N_7663,N_1594,N_41);
and U7664 (N_7664,N_1189,N_467);
xor U7665 (N_7665,N_602,N_631);
nor U7666 (N_7666,N_4540,N_2262);
or U7667 (N_7667,N_3497,N_280);
nand U7668 (N_7668,N_4326,N_1714);
and U7669 (N_7669,N_307,N_691);
nor U7670 (N_7670,N_2327,N_1986);
nand U7671 (N_7671,N_841,N_3917);
and U7672 (N_7672,N_216,N_1102);
or U7673 (N_7673,N_993,N_3767);
nor U7674 (N_7674,N_4002,N_493);
or U7675 (N_7675,N_2365,N_1014);
and U7676 (N_7676,N_3165,N_2127);
or U7677 (N_7677,N_4609,N_2963);
and U7678 (N_7678,N_2308,N_276);
nand U7679 (N_7679,N_4684,N_399);
nand U7680 (N_7680,N_2487,N_1474);
and U7681 (N_7681,N_134,N_924);
xor U7682 (N_7682,N_135,N_4680);
xor U7683 (N_7683,N_4955,N_2311);
and U7684 (N_7684,N_2190,N_1842);
nand U7685 (N_7685,N_1712,N_425);
xnor U7686 (N_7686,N_1225,N_3505);
xor U7687 (N_7687,N_4292,N_3215);
xor U7688 (N_7688,N_2011,N_2708);
and U7689 (N_7689,N_3447,N_67);
nand U7690 (N_7690,N_4713,N_2383);
nand U7691 (N_7691,N_213,N_2949);
xnor U7692 (N_7692,N_3073,N_1862);
xnor U7693 (N_7693,N_4778,N_4049);
or U7694 (N_7694,N_2856,N_2397);
or U7695 (N_7695,N_3808,N_2932);
xnor U7696 (N_7696,N_1242,N_4562);
xnor U7697 (N_7697,N_1839,N_3159);
nor U7698 (N_7698,N_8,N_3808);
nor U7699 (N_7699,N_2756,N_1118);
nor U7700 (N_7700,N_403,N_2677);
xor U7701 (N_7701,N_3255,N_798);
or U7702 (N_7702,N_2697,N_1482);
or U7703 (N_7703,N_3982,N_314);
and U7704 (N_7704,N_617,N_3852);
nor U7705 (N_7705,N_115,N_3931);
and U7706 (N_7706,N_384,N_1815);
xnor U7707 (N_7707,N_510,N_135);
and U7708 (N_7708,N_3772,N_3433);
xor U7709 (N_7709,N_4317,N_2808);
and U7710 (N_7710,N_3013,N_862);
nand U7711 (N_7711,N_1557,N_2753);
and U7712 (N_7712,N_4367,N_3430);
and U7713 (N_7713,N_3326,N_2177);
nor U7714 (N_7714,N_3272,N_4642);
nor U7715 (N_7715,N_3701,N_481);
nor U7716 (N_7716,N_3450,N_1923);
nor U7717 (N_7717,N_283,N_3919);
nand U7718 (N_7718,N_3824,N_2948);
nor U7719 (N_7719,N_4516,N_1637);
xor U7720 (N_7720,N_292,N_2771);
or U7721 (N_7721,N_3878,N_4858);
nand U7722 (N_7722,N_3325,N_4222);
xor U7723 (N_7723,N_3278,N_1555);
nand U7724 (N_7724,N_2199,N_4042);
xnor U7725 (N_7725,N_3892,N_4433);
nor U7726 (N_7726,N_3692,N_1354);
nand U7727 (N_7727,N_4810,N_65);
and U7728 (N_7728,N_2920,N_3798);
xnor U7729 (N_7729,N_3875,N_4738);
and U7730 (N_7730,N_1364,N_1089);
nor U7731 (N_7731,N_820,N_3472);
or U7732 (N_7732,N_1603,N_3751);
nand U7733 (N_7733,N_3638,N_4390);
nor U7734 (N_7734,N_2794,N_254);
or U7735 (N_7735,N_2624,N_1242);
or U7736 (N_7736,N_3098,N_2626);
nand U7737 (N_7737,N_607,N_196);
or U7738 (N_7738,N_4333,N_1251);
and U7739 (N_7739,N_1361,N_1302);
nand U7740 (N_7740,N_1070,N_559);
nand U7741 (N_7741,N_2397,N_4723);
nand U7742 (N_7742,N_903,N_1782);
nor U7743 (N_7743,N_4031,N_2682);
nand U7744 (N_7744,N_1947,N_2629);
or U7745 (N_7745,N_4830,N_2017);
or U7746 (N_7746,N_676,N_4070);
xnor U7747 (N_7747,N_2748,N_2557);
and U7748 (N_7748,N_3956,N_1672);
xor U7749 (N_7749,N_3330,N_578);
and U7750 (N_7750,N_615,N_3428);
or U7751 (N_7751,N_522,N_3213);
or U7752 (N_7752,N_2513,N_2065);
nand U7753 (N_7753,N_2876,N_4849);
or U7754 (N_7754,N_66,N_2942);
nor U7755 (N_7755,N_851,N_2831);
or U7756 (N_7756,N_4407,N_814);
or U7757 (N_7757,N_2019,N_888);
nand U7758 (N_7758,N_2494,N_2282);
or U7759 (N_7759,N_2364,N_1765);
or U7760 (N_7760,N_2953,N_3387);
nor U7761 (N_7761,N_4179,N_3667);
or U7762 (N_7762,N_1648,N_3582);
nor U7763 (N_7763,N_895,N_1634);
and U7764 (N_7764,N_3975,N_2954);
xnor U7765 (N_7765,N_4141,N_1184);
nor U7766 (N_7766,N_1247,N_786);
xnor U7767 (N_7767,N_4877,N_1316);
xor U7768 (N_7768,N_998,N_4839);
or U7769 (N_7769,N_3608,N_3959);
and U7770 (N_7770,N_4540,N_3564);
xor U7771 (N_7771,N_1434,N_4272);
or U7772 (N_7772,N_3909,N_4149);
and U7773 (N_7773,N_4664,N_3048);
nor U7774 (N_7774,N_666,N_2684);
nor U7775 (N_7775,N_3126,N_258);
nor U7776 (N_7776,N_1867,N_1680);
or U7777 (N_7777,N_4557,N_1268);
nand U7778 (N_7778,N_1834,N_4080);
and U7779 (N_7779,N_75,N_608);
nand U7780 (N_7780,N_896,N_3491);
and U7781 (N_7781,N_4822,N_3192);
nor U7782 (N_7782,N_420,N_3727);
xor U7783 (N_7783,N_587,N_276);
or U7784 (N_7784,N_3609,N_3589);
nor U7785 (N_7785,N_4296,N_4265);
or U7786 (N_7786,N_4811,N_4465);
and U7787 (N_7787,N_2285,N_649);
and U7788 (N_7788,N_1226,N_2010);
or U7789 (N_7789,N_956,N_3488);
or U7790 (N_7790,N_53,N_4360);
xor U7791 (N_7791,N_3359,N_1469);
and U7792 (N_7792,N_1119,N_454);
nand U7793 (N_7793,N_347,N_2214);
nand U7794 (N_7794,N_4987,N_4338);
or U7795 (N_7795,N_1396,N_2925);
xor U7796 (N_7796,N_1807,N_4179);
and U7797 (N_7797,N_3132,N_2568);
or U7798 (N_7798,N_122,N_964);
nor U7799 (N_7799,N_3783,N_4211);
xor U7800 (N_7800,N_807,N_2462);
or U7801 (N_7801,N_4949,N_4194);
xor U7802 (N_7802,N_1818,N_1971);
or U7803 (N_7803,N_4269,N_2521);
xnor U7804 (N_7804,N_1135,N_2385);
xor U7805 (N_7805,N_4144,N_799);
and U7806 (N_7806,N_2742,N_2303);
or U7807 (N_7807,N_2420,N_4972);
xor U7808 (N_7808,N_2397,N_1127);
nand U7809 (N_7809,N_2283,N_984);
or U7810 (N_7810,N_1977,N_2434);
or U7811 (N_7811,N_4464,N_363);
and U7812 (N_7812,N_4943,N_3110);
nand U7813 (N_7813,N_511,N_4363);
nand U7814 (N_7814,N_3543,N_2534);
nor U7815 (N_7815,N_1786,N_3054);
and U7816 (N_7816,N_3327,N_2664);
nand U7817 (N_7817,N_4718,N_2362);
xnor U7818 (N_7818,N_2861,N_2486);
and U7819 (N_7819,N_751,N_1055);
xnor U7820 (N_7820,N_969,N_717);
xnor U7821 (N_7821,N_4759,N_3802);
and U7822 (N_7822,N_1812,N_3043);
or U7823 (N_7823,N_4519,N_95);
and U7824 (N_7824,N_4433,N_4233);
xnor U7825 (N_7825,N_646,N_349);
or U7826 (N_7826,N_2892,N_3921);
nand U7827 (N_7827,N_2819,N_4785);
xnor U7828 (N_7828,N_309,N_4036);
xnor U7829 (N_7829,N_631,N_510);
and U7830 (N_7830,N_1106,N_1327);
or U7831 (N_7831,N_834,N_558);
or U7832 (N_7832,N_4185,N_3765);
xnor U7833 (N_7833,N_2270,N_1076);
xor U7834 (N_7834,N_4180,N_2924);
and U7835 (N_7835,N_1699,N_4911);
or U7836 (N_7836,N_854,N_1998);
xor U7837 (N_7837,N_4597,N_679);
nor U7838 (N_7838,N_325,N_1546);
or U7839 (N_7839,N_1466,N_2299);
nor U7840 (N_7840,N_3151,N_373);
nand U7841 (N_7841,N_1605,N_4060);
and U7842 (N_7842,N_3973,N_2005);
and U7843 (N_7843,N_1478,N_3107);
or U7844 (N_7844,N_702,N_1730);
and U7845 (N_7845,N_3445,N_2971);
and U7846 (N_7846,N_2263,N_1578);
xor U7847 (N_7847,N_4026,N_1070);
xnor U7848 (N_7848,N_4149,N_4452);
nand U7849 (N_7849,N_4106,N_4690);
nor U7850 (N_7850,N_500,N_4782);
xor U7851 (N_7851,N_4643,N_1250);
or U7852 (N_7852,N_16,N_3700);
and U7853 (N_7853,N_2987,N_979);
nor U7854 (N_7854,N_2139,N_790);
nor U7855 (N_7855,N_554,N_601);
xnor U7856 (N_7856,N_2923,N_1812);
or U7857 (N_7857,N_836,N_4184);
and U7858 (N_7858,N_625,N_3057);
nand U7859 (N_7859,N_2348,N_2238);
xor U7860 (N_7860,N_4215,N_1541);
and U7861 (N_7861,N_958,N_240);
and U7862 (N_7862,N_568,N_4042);
nor U7863 (N_7863,N_4939,N_915);
nor U7864 (N_7864,N_4911,N_3515);
and U7865 (N_7865,N_4150,N_579);
nor U7866 (N_7866,N_3486,N_184);
or U7867 (N_7867,N_4495,N_1124);
nand U7868 (N_7868,N_4705,N_3449);
or U7869 (N_7869,N_4973,N_3608);
nand U7870 (N_7870,N_1929,N_3657);
nand U7871 (N_7871,N_1203,N_2598);
and U7872 (N_7872,N_2449,N_4676);
nor U7873 (N_7873,N_3930,N_1063);
nor U7874 (N_7874,N_3892,N_2536);
nand U7875 (N_7875,N_1569,N_722);
or U7876 (N_7876,N_1292,N_2532);
nand U7877 (N_7877,N_4836,N_483);
nand U7878 (N_7878,N_1947,N_1258);
nand U7879 (N_7879,N_4478,N_2511);
xnor U7880 (N_7880,N_2758,N_4886);
xor U7881 (N_7881,N_2259,N_4652);
nor U7882 (N_7882,N_284,N_1596);
or U7883 (N_7883,N_2004,N_1998);
nand U7884 (N_7884,N_3718,N_2745);
or U7885 (N_7885,N_499,N_3174);
or U7886 (N_7886,N_3724,N_4273);
nand U7887 (N_7887,N_3052,N_4830);
xor U7888 (N_7888,N_552,N_3445);
nor U7889 (N_7889,N_2453,N_2046);
nor U7890 (N_7890,N_2443,N_2071);
xnor U7891 (N_7891,N_2461,N_3263);
and U7892 (N_7892,N_4692,N_4073);
and U7893 (N_7893,N_4874,N_3952);
or U7894 (N_7894,N_1994,N_2057);
nor U7895 (N_7895,N_4469,N_475);
nand U7896 (N_7896,N_920,N_4730);
or U7897 (N_7897,N_2927,N_4449);
or U7898 (N_7898,N_3852,N_1648);
xor U7899 (N_7899,N_2448,N_1075);
nor U7900 (N_7900,N_4180,N_3521);
xnor U7901 (N_7901,N_465,N_1976);
nor U7902 (N_7902,N_963,N_1881);
nand U7903 (N_7903,N_2030,N_4935);
nand U7904 (N_7904,N_700,N_2415);
nand U7905 (N_7905,N_3736,N_4579);
nor U7906 (N_7906,N_2690,N_143);
nor U7907 (N_7907,N_4420,N_3335);
nor U7908 (N_7908,N_2674,N_4596);
nor U7909 (N_7909,N_2729,N_3546);
xnor U7910 (N_7910,N_2877,N_412);
nand U7911 (N_7911,N_982,N_3016);
and U7912 (N_7912,N_1913,N_4085);
xor U7913 (N_7913,N_2990,N_1767);
nand U7914 (N_7914,N_3096,N_1520);
nand U7915 (N_7915,N_2370,N_4111);
or U7916 (N_7916,N_1387,N_3530);
and U7917 (N_7917,N_3211,N_3475);
nor U7918 (N_7918,N_3293,N_4472);
nor U7919 (N_7919,N_1135,N_1480);
nor U7920 (N_7920,N_2786,N_3162);
and U7921 (N_7921,N_3312,N_1388);
or U7922 (N_7922,N_1884,N_2668);
xnor U7923 (N_7923,N_4797,N_3563);
nor U7924 (N_7924,N_2524,N_4347);
xor U7925 (N_7925,N_1846,N_3479);
xnor U7926 (N_7926,N_4566,N_3968);
nand U7927 (N_7927,N_132,N_1919);
nor U7928 (N_7928,N_3144,N_3973);
nand U7929 (N_7929,N_4090,N_1836);
or U7930 (N_7930,N_499,N_3184);
xor U7931 (N_7931,N_1504,N_1733);
or U7932 (N_7932,N_2378,N_206);
nand U7933 (N_7933,N_4597,N_3510);
nand U7934 (N_7934,N_3408,N_3970);
nand U7935 (N_7935,N_2583,N_2845);
xnor U7936 (N_7936,N_3781,N_2779);
nor U7937 (N_7937,N_4912,N_4285);
or U7938 (N_7938,N_2613,N_2052);
and U7939 (N_7939,N_3633,N_1112);
and U7940 (N_7940,N_4663,N_925);
or U7941 (N_7941,N_307,N_3237);
nor U7942 (N_7942,N_2143,N_2554);
or U7943 (N_7943,N_809,N_1804);
nand U7944 (N_7944,N_1451,N_4607);
nand U7945 (N_7945,N_581,N_4780);
nand U7946 (N_7946,N_297,N_1890);
and U7947 (N_7947,N_4980,N_2106);
nor U7948 (N_7948,N_2191,N_183);
nand U7949 (N_7949,N_3220,N_2786);
xor U7950 (N_7950,N_39,N_4268);
nor U7951 (N_7951,N_4296,N_672);
nand U7952 (N_7952,N_365,N_3703);
and U7953 (N_7953,N_15,N_3470);
or U7954 (N_7954,N_4807,N_3241);
xnor U7955 (N_7955,N_2807,N_2279);
and U7956 (N_7956,N_1677,N_830);
xnor U7957 (N_7957,N_3973,N_3553);
and U7958 (N_7958,N_3161,N_3355);
xnor U7959 (N_7959,N_2962,N_4845);
nand U7960 (N_7960,N_793,N_1233);
or U7961 (N_7961,N_3303,N_2195);
xor U7962 (N_7962,N_1359,N_1095);
nor U7963 (N_7963,N_3240,N_1423);
xnor U7964 (N_7964,N_4015,N_66);
xor U7965 (N_7965,N_144,N_3843);
or U7966 (N_7966,N_968,N_1293);
nor U7967 (N_7967,N_83,N_3288);
nor U7968 (N_7968,N_326,N_1606);
nor U7969 (N_7969,N_1157,N_331);
or U7970 (N_7970,N_2009,N_2674);
xor U7971 (N_7971,N_2348,N_1588);
or U7972 (N_7972,N_3346,N_2607);
nor U7973 (N_7973,N_746,N_94);
nand U7974 (N_7974,N_136,N_3669);
nand U7975 (N_7975,N_3436,N_4539);
nand U7976 (N_7976,N_3842,N_4249);
and U7977 (N_7977,N_4675,N_3118);
and U7978 (N_7978,N_1319,N_510);
xnor U7979 (N_7979,N_4929,N_2064);
nand U7980 (N_7980,N_4889,N_4431);
and U7981 (N_7981,N_725,N_1189);
and U7982 (N_7982,N_1135,N_3470);
nor U7983 (N_7983,N_1237,N_769);
nor U7984 (N_7984,N_2522,N_2947);
xnor U7985 (N_7985,N_2426,N_1034);
nor U7986 (N_7986,N_4769,N_4624);
or U7987 (N_7987,N_4988,N_4782);
xor U7988 (N_7988,N_900,N_199);
or U7989 (N_7989,N_490,N_1349);
nor U7990 (N_7990,N_602,N_2065);
and U7991 (N_7991,N_1300,N_3460);
and U7992 (N_7992,N_2983,N_3447);
nor U7993 (N_7993,N_1670,N_4959);
and U7994 (N_7994,N_2971,N_427);
and U7995 (N_7995,N_4873,N_3574);
xor U7996 (N_7996,N_3291,N_3801);
and U7997 (N_7997,N_2225,N_3468);
xor U7998 (N_7998,N_2685,N_206);
or U7999 (N_7999,N_4243,N_675);
xor U8000 (N_8000,N_3322,N_4175);
and U8001 (N_8001,N_206,N_4190);
xnor U8002 (N_8002,N_3410,N_3558);
nand U8003 (N_8003,N_2194,N_1156);
nor U8004 (N_8004,N_4550,N_463);
and U8005 (N_8005,N_2286,N_4640);
nand U8006 (N_8006,N_4049,N_4294);
nor U8007 (N_8007,N_3922,N_4780);
and U8008 (N_8008,N_953,N_1806);
xor U8009 (N_8009,N_1259,N_3861);
nand U8010 (N_8010,N_3869,N_1033);
and U8011 (N_8011,N_2040,N_531);
and U8012 (N_8012,N_4220,N_2750);
and U8013 (N_8013,N_4253,N_3029);
nand U8014 (N_8014,N_1904,N_3713);
and U8015 (N_8015,N_2273,N_453);
xnor U8016 (N_8016,N_69,N_2963);
and U8017 (N_8017,N_2871,N_2938);
nor U8018 (N_8018,N_587,N_1168);
nor U8019 (N_8019,N_62,N_472);
or U8020 (N_8020,N_3024,N_1763);
nor U8021 (N_8021,N_4243,N_1691);
nand U8022 (N_8022,N_1283,N_316);
and U8023 (N_8023,N_949,N_3165);
nor U8024 (N_8024,N_1175,N_2986);
or U8025 (N_8025,N_4399,N_1948);
and U8026 (N_8026,N_3312,N_2377);
nand U8027 (N_8027,N_2374,N_351);
xor U8028 (N_8028,N_1644,N_396);
and U8029 (N_8029,N_3597,N_1326);
nand U8030 (N_8030,N_4061,N_4767);
or U8031 (N_8031,N_4851,N_2198);
xnor U8032 (N_8032,N_3348,N_1159);
and U8033 (N_8033,N_3021,N_144);
or U8034 (N_8034,N_30,N_4708);
or U8035 (N_8035,N_4488,N_4407);
nand U8036 (N_8036,N_1260,N_137);
nor U8037 (N_8037,N_2477,N_3674);
or U8038 (N_8038,N_1788,N_2312);
and U8039 (N_8039,N_4269,N_294);
nand U8040 (N_8040,N_3814,N_272);
nand U8041 (N_8041,N_4628,N_166);
and U8042 (N_8042,N_296,N_3319);
or U8043 (N_8043,N_1080,N_4327);
or U8044 (N_8044,N_3727,N_199);
nand U8045 (N_8045,N_1267,N_1201);
or U8046 (N_8046,N_403,N_2129);
nand U8047 (N_8047,N_4049,N_2085);
or U8048 (N_8048,N_1180,N_1545);
nor U8049 (N_8049,N_2875,N_3537);
nor U8050 (N_8050,N_3920,N_1832);
nor U8051 (N_8051,N_1811,N_2415);
or U8052 (N_8052,N_1997,N_2784);
or U8053 (N_8053,N_3827,N_314);
xnor U8054 (N_8054,N_2490,N_1193);
xor U8055 (N_8055,N_4355,N_684);
xnor U8056 (N_8056,N_221,N_3533);
and U8057 (N_8057,N_3068,N_3933);
or U8058 (N_8058,N_1896,N_4345);
and U8059 (N_8059,N_4492,N_4778);
nor U8060 (N_8060,N_3519,N_1678);
nand U8061 (N_8061,N_924,N_112);
xnor U8062 (N_8062,N_1258,N_1166);
or U8063 (N_8063,N_3503,N_1493);
or U8064 (N_8064,N_3552,N_4862);
and U8065 (N_8065,N_1898,N_825);
nand U8066 (N_8066,N_2374,N_3236);
and U8067 (N_8067,N_1180,N_159);
nor U8068 (N_8068,N_3028,N_168);
and U8069 (N_8069,N_2702,N_3800);
and U8070 (N_8070,N_4467,N_4455);
nor U8071 (N_8071,N_4827,N_33);
or U8072 (N_8072,N_4480,N_2571);
nor U8073 (N_8073,N_1683,N_1141);
nor U8074 (N_8074,N_1258,N_1716);
and U8075 (N_8075,N_3302,N_1524);
and U8076 (N_8076,N_233,N_528);
nor U8077 (N_8077,N_1270,N_2003);
nand U8078 (N_8078,N_2376,N_3488);
xnor U8079 (N_8079,N_110,N_4347);
and U8080 (N_8080,N_4223,N_2129);
xor U8081 (N_8081,N_122,N_4296);
and U8082 (N_8082,N_1138,N_1627);
nand U8083 (N_8083,N_732,N_3096);
xor U8084 (N_8084,N_2774,N_2685);
nor U8085 (N_8085,N_564,N_3137);
and U8086 (N_8086,N_832,N_2345);
and U8087 (N_8087,N_2159,N_3799);
nor U8088 (N_8088,N_534,N_1939);
or U8089 (N_8089,N_3289,N_2701);
and U8090 (N_8090,N_2206,N_839);
and U8091 (N_8091,N_3364,N_4980);
nand U8092 (N_8092,N_103,N_2438);
and U8093 (N_8093,N_2034,N_4611);
nand U8094 (N_8094,N_2146,N_2840);
xnor U8095 (N_8095,N_4282,N_535);
nor U8096 (N_8096,N_2385,N_3878);
nand U8097 (N_8097,N_4184,N_803);
nor U8098 (N_8098,N_2957,N_1620);
nand U8099 (N_8099,N_0,N_4225);
and U8100 (N_8100,N_1712,N_957);
and U8101 (N_8101,N_1289,N_2050);
xor U8102 (N_8102,N_784,N_4801);
nand U8103 (N_8103,N_3415,N_247);
and U8104 (N_8104,N_2411,N_2068);
xor U8105 (N_8105,N_4737,N_4854);
and U8106 (N_8106,N_2158,N_4301);
nor U8107 (N_8107,N_4193,N_4413);
nor U8108 (N_8108,N_1250,N_548);
and U8109 (N_8109,N_2220,N_1103);
nand U8110 (N_8110,N_4636,N_842);
nor U8111 (N_8111,N_2810,N_1878);
nand U8112 (N_8112,N_4930,N_4005);
and U8113 (N_8113,N_2381,N_3339);
or U8114 (N_8114,N_4533,N_2407);
and U8115 (N_8115,N_500,N_670);
nand U8116 (N_8116,N_1551,N_3057);
xnor U8117 (N_8117,N_3581,N_3654);
and U8118 (N_8118,N_1518,N_2283);
or U8119 (N_8119,N_2262,N_1418);
xnor U8120 (N_8120,N_3592,N_3812);
and U8121 (N_8121,N_571,N_3288);
nand U8122 (N_8122,N_2207,N_4264);
nor U8123 (N_8123,N_1044,N_2711);
xor U8124 (N_8124,N_1369,N_3949);
xnor U8125 (N_8125,N_470,N_4401);
nor U8126 (N_8126,N_4517,N_87);
or U8127 (N_8127,N_162,N_2874);
xnor U8128 (N_8128,N_4560,N_3829);
nor U8129 (N_8129,N_3752,N_2311);
nor U8130 (N_8130,N_4645,N_659);
nand U8131 (N_8131,N_255,N_2875);
nand U8132 (N_8132,N_4021,N_4900);
or U8133 (N_8133,N_508,N_2731);
nand U8134 (N_8134,N_2092,N_747);
xnor U8135 (N_8135,N_3099,N_1859);
nor U8136 (N_8136,N_2386,N_2988);
or U8137 (N_8137,N_918,N_2274);
nand U8138 (N_8138,N_3808,N_1219);
and U8139 (N_8139,N_4238,N_3162);
xor U8140 (N_8140,N_3422,N_1874);
or U8141 (N_8141,N_3917,N_4357);
nor U8142 (N_8142,N_2273,N_607);
and U8143 (N_8143,N_3506,N_1168);
or U8144 (N_8144,N_4930,N_4068);
or U8145 (N_8145,N_1488,N_381);
or U8146 (N_8146,N_2202,N_1948);
xor U8147 (N_8147,N_4940,N_1458);
xor U8148 (N_8148,N_2529,N_4427);
nor U8149 (N_8149,N_3446,N_2805);
and U8150 (N_8150,N_4669,N_1678);
and U8151 (N_8151,N_155,N_692);
xnor U8152 (N_8152,N_1514,N_3770);
or U8153 (N_8153,N_1020,N_3085);
or U8154 (N_8154,N_3709,N_2611);
xor U8155 (N_8155,N_4786,N_156);
and U8156 (N_8156,N_3625,N_732);
nor U8157 (N_8157,N_2612,N_3517);
xnor U8158 (N_8158,N_2044,N_2411);
or U8159 (N_8159,N_1079,N_1929);
nand U8160 (N_8160,N_4421,N_1562);
nand U8161 (N_8161,N_4414,N_601);
or U8162 (N_8162,N_4155,N_366);
nand U8163 (N_8163,N_1449,N_2130);
nor U8164 (N_8164,N_1529,N_1603);
xnor U8165 (N_8165,N_2859,N_1686);
nor U8166 (N_8166,N_1417,N_2659);
and U8167 (N_8167,N_4700,N_1906);
nand U8168 (N_8168,N_4005,N_1882);
or U8169 (N_8169,N_4570,N_4329);
nor U8170 (N_8170,N_363,N_3372);
nor U8171 (N_8171,N_3237,N_4918);
or U8172 (N_8172,N_365,N_4095);
nor U8173 (N_8173,N_1619,N_2596);
nand U8174 (N_8174,N_2820,N_4805);
or U8175 (N_8175,N_695,N_4663);
nand U8176 (N_8176,N_2543,N_3597);
nor U8177 (N_8177,N_3085,N_4934);
and U8178 (N_8178,N_1086,N_2217);
and U8179 (N_8179,N_3,N_2686);
nor U8180 (N_8180,N_1906,N_2842);
nand U8181 (N_8181,N_2263,N_3849);
and U8182 (N_8182,N_366,N_3333);
or U8183 (N_8183,N_3194,N_2094);
nor U8184 (N_8184,N_2011,N_4933);
or U8185 (N_8185,N_4924,N_4501);
nor U8186 (N_8186,N_2419,N_2368);
and U8187 (N_8187,N_2125,N_3705);
nand U8188 (N_8188,N_1982,N_2414);
nor U8189 (N_8189,N_2538,N_4241);
xor U8190 (N_8190,N_4205,N_3088);
nor U8191 (N_8191,N_3432,N_2556);
nor U8192 (N_8192,N_3038,N_554);
and U8193 (N_8193,N_2333,N_3758);
xor U8194 (N_8194,N_1851,N_4004);
or U8195 (N_8195,N_1037,N_1454);
or U8196 (N_8196,N_72,N_3696);
or U8197 (N_8197,N_3833,N_129);
nor U8198 (N_8198,N_4460,N_4481);
nand U8199 (N_8199,N_449,N_1948);
and U8200 (N_8200,N_3338,N_4111);
or U8201 (N_8201,N_4595,N_2082);
nor U8202 (N_8202,N_184,N_2760);
nand U8203 (N_8203,N_4412,N_3006);
nor U8204 (N_8204,N_2315,N_1553);
and U8205 (N_8205,N_2364,N_4566);
xnor U8206 (N_8206,N_1616,N_2268);
xnor U8207 (N_8207,N_1675,N_1079);
xnor U8208 (N_8208,N_3233,N_3824);
nor U8209 (N_8209,N_3874,N_753);
and U8210 (N_8210,N_200,N_3951);
or U8211 (N_8211,N_2983,N_3204);
nor U8212 (N_8212,N_3692,N_4807);
and U8213 (N_8213,N_3866,N_1613);
nand U8214 (N_8214,N_16,N_899);
and U8215 (N_8215,N_1388,N_1964);
nand U8216 (N_8216,N_4603,N_1662);
nor U8217 (N_8217,N_2891,N_3112);
nand U8218 (N_8218,N_3689,N_1871);
xnor U8219 (N_8219,N_1074,N_1200);
nor U8220 (N_8220,N_1878,N_2498);
xnor U8221 (N_8221,N_2682,N_2275);
or U8222 (N_8222,N_4717,N_3206);
nor U8223 (N_8223,N_2650,N_1968);
or U8224 (N_8224,N_4747,N_804);
nand U8225 (N_8225,N_1615,N_2666);
nand U8226 (N_8226,N_1427,N_2214);
nand U8227 (N_8227,N_4982,N_191);
or U8228 (N_8228,N_1065,N_1039);
nor U8229 (N_8229,N_1225,N_2251);
or U8230 (N_8230,N_2556,N_4028);
or U8231 (N_8231,N_2573,N_3145);
and U8232 (N_8232,N_1944,N_3592);
nor U8233 (N_8233,N_1676,N_1626);
nand U8234 (N_8234,N_4365,N_4751);
or U8235 (N_8235,N_47,N_955);
or U8236 (N_8236,N_927,N_2228);
and U8237 (N_8237,N_4449,N_3551);
nand U8238 (N_8238,N_543,N_3022);
and U8239 (N_8239,N_938,N_963);
nand U8240 (N_8240,N_2338,N_4877);
nand U8241 (N_8241,N_471,N_3451);
nor U8242 (N_8242,N_4657,N_880);
xnor U8243 (N_8243,N_1356,N_3650);
nor U8244 (N_8244,N_2767,N_266);
nor U8245 (N_8245,N_3767,N_66);
or U8246 (N_8246,N_3103,N_2793);
or U8247 (N_8247,N_502,N_2293);
and U8248 (N_8248,N_967,N_4382);
nand U8249 (N_8249,N_3501,N_4945);
nor U8250 (N_8250,N_575,N_1859);
xnor U8251 (N_8251,N_4916,N_327);
nand U8252 (N_8252,N_2596,N_4362);
or U8253 (N_8253,N_586,N_2175);
nor U8254 (N_8254,N_3743,N_4388);
or U8255 (N_8255,N_534,N_2428);
nor U8256 (N_8256,N_2091,N_2697);
nand U8257 (N_8257,N_760,N_4666);
or U8258 (N_8258,N_2481,N_2483);
or U8259 (N_8259,N_3181,N_4564);
xor U8260 (N_8260,N_3991,N_3039);
xor U8261 (N_8261,N_2848,N_2043);
or U8262 (N_8262,N_1888,N_651);
or U8263 (N_8263,N_1843,N_4527);
xnor U8264 (N_8264,N_1719,N_1800);
or U8265 (N_8265,N_1999,N_3195);
or U8266 (N_8266,N_3004,N_1688);
or U8267 (N_8267,N_1075,N_4430);
or U8268 (N_8268,N_4079,N_94);
and U8269 (N_8269,N_3527,N_1765);
nand U8270 (N_8270,N_4687,N_4904);
nor U8271 (N_8271,N_4660,N_3320);
and U8272 (N_8272,N_1030,N_583);
xor U8273 (N_8273,N_3764,N_2564);
or U8274 (N_8274,N_426,N_2065);
nor U8275 (N_8275,N_3400,N_1101);
nor U8276 (N_8276,N_4301,N_3722);
or U8277 (N_8277,N_3615,N_540);
xor U8278 (N_8278,N_510,N_2420);
and U8279 (N_8279,N_737,N_4295);
nor U8280 (N_8280,N_615,N_2722);
xor U8281 (N_8281,N_3599,N_244);
xnor U8282 (N_8282,N_3497,N_4873);
nand U8283 (N_8283,N_2892,N_4230);
or U8284 (N_8284,N_4201,N_2565);
or U8285 (N_8285,N_3891,N_715);
and U8286 (N_8286,N_3904,N_1546);
nand U8287 (N_8287,N_1241,N_2583);
and U8288 (N_8288,N_3447,N_825);
nor U8289 (N_8289,N_622,N_1775);
and U8290 (N_8290,N_403,N_4459);
nand U8291 (N_8291,N_855,N_3451);
or U8292 (N_8292,N_3800,N_1807);
nor U8293 (N_8293,N_767,N_2985);
xnor U8294 (N_8294,N_3512,N_3426);
and U8295 (N_8295,N_657,N_2118);
or U8296 (N_8296,N_1812,N_2500);
or U8297 (N_8297,N_4852,N_3012);
or U8298 (N_8298,N_2313,N_2673);
nand U8299 (N_8299,N_2006,N_1802);
and U8300 (N_8300,N_1180,N_3871);
nor U8301 (N_8301,N_2864,N_4320);
or U8302 (N_8302,N_3658,N_4454);
or U8303 (N_8303,N_4257,N_490);
nor U8304 (N_8304,N_1704,N_2041);
or U8305 (N_8305,N_2760,N_4340);
xor U8306 (N_8306,N_2769,N_851);
nand U8307 (N_8307,N_1865,N_655);
or U8308 (N_8308,N_2737,N_330);
or U8309 (N_8309,N_3477,N_2599);
or U8310 (N_8310,N_3759,N_1573);
nor U8311 (N_8311,N_4061,N_448);
nand U8312 (N_8312,N_2183,N_3565);
and U8313 (N_8313,N_1854,N_4860);
and U8314 (N_8314,N_2764,N_4480);
nor U8315 (N_8315,N_2947,N_1157);
nand U8316 (N_8316,N_2663,N_452);
nand U8317 (N_8317,N_3897,N_2436);
or U8318 (N_8318,N_2583,N_4280);
nand U8319 (N_8319,N_3812,N_3637);
xnor U8320 (N_8320,N_4334,N_3587);
or U8321 (N_8321,N_4690,N_4395);
and U8322 (N_8322,N_2618,N_1359);
nand U8323 (N_8323,N_4997,N_1239);
nand U8324 (N_8324,N_3430,N_2445);
and U8325 (N_8325,N_4828,N_2817);
xnor U8326 (N_8326,N_2318,N_2065);
or U8327 (N_8327,N_970,N_1101);
or U8328 (N_8328,N_33,N_321);
or U8329 (N_8329,N_2635,N_1857);
or U8330 (N_8330,N_634,N_4047);
nor U8331 (N_8331,N_1773,N_1649);
nor U8332 (N_8332,N_22,N_1965);
nor U8333 (N_8333,N_2086,N_1668);
nand U8334 (N_8334,N_4043,N_791);
xor U8335 (N_8335,N_3118,N_4988);
xnor U8336 (N_8336,N_3333,N_160);
nand U8337 (N_8337,N_4759,N_1520);
nor U8338 (N_8338,N_4697,N_2147);
nand U8339 (N_8339,N_576,N_1580);
nand U8340 (N_8340,N_3966,N_4149);
and U8341 (N_8341,N_1538,N_3300);
xor U8342 (N_8342,N_3498,N_3221);
and U8343 (N_8343,N_2930,N_4578);
nand U8344 (N_8344,N_3000,N_4216);
nor U8345 (N_8345,N_4105,N_1172);
or U8346 (N_8346,N_4673,N_3327);
xnor U8347 (N_8347,N_3731,N_1603);
xor U8348 (N_8348,N_4432,N_3587);
and U8349 (N_8349,N_2945,N_35);
and U8350 (N_8350,N_747,N_4527);
nor U8351 (N_8351,N_1131,N_2817);
xor U8352 (N_8352,N_221,N_1972);
xor U8353 (N_8353,N_463,N_1916);
or U8354 (N_8354,N_4956,N_4768);
nand U8355 (N_8355,N_2304,N_3936);
and U8356 (N_8356,N_3974,N_1989);
and U8357 (N_8357,N_4281,N_763);
xor U8358 (N_8358,N_4008,N_549);
nor U8359 (N_8359,N_1845,N_282);
xnor U8360 (N_8360,N_4893,N_1827);
xnor U8361 (N_8361,N_2047,N_1161);
nand U8362 (N_8362,N_4401,N_163);
or U8363 (N_8363,N_1014,N_3259);
xnor U8364 (N_8364,N_4514,N_3247);
and U8365 (N_8365,N_3620,N_800);
nor U8366 (N_8366,N_1041,N_2240);
xnor U8367 (N_8367,N_4897,N_1790);
and U8368 (N_8368,N_3317,N_1089);
nor U8369 (N_8369,N_4192,N_1865);
or U8370 (N_8370,N_4158,N_2801);
nand U8371 (N_8371,N_4903,N_4557);
and U8372 (N_8372,N_918,N_1570);
or U8373 (N_8373,N_3347,N_3111);
or U8374 (N_8374,N_793,N_2105);
nor U8375 (N_8375,N_1830,N_3667);
and U8376 (N_8376,N_4522,N_4261);
and U8377 (N_8377,N_181,N_4682);
and U8378 (N_8378,N_3402,N_1701);
xnor U8379 (N_8379,N_202,N_3177);
nand U8380 (N_8380,N_1266,N_693);
xor U8381 (N_8381,N_513,N_3476);
nand U8382 (N_8382,N_584,N_4361);
nand U8383 (N_8383,N_4966,N_540);
or U8384 (N_8384,N_2152,N_2167);
nand U8385 (N_8385,N_2670,N_1336);
xor U8386 (N_8386,N_3459,N_3759);
nand U8387 (N_8387,N_766,N_3071);
and U8388 (N_8388,N_3485,N_471);
nor U8389 (N_8389,N_230,N_1414);
and U8390 (N_8390,N_1938,N_1469);
and U8391 (N_8391,N_2117,N_699);
xor U8392 (N_8392,N_4115,N_2898);
nor U8393 (N_8393,N_2504,N_2157);
or U8394 (N_8394,N_259,N_300);
and U8395 (N_8395,N_308,N_2284);
and U8396 (N_8396,N_2823,N_231);
nor U8397 (N_8397,N_750,N_2985);
or U8398 (N_8398,N_2229,N_522);
nand U8399 (N_8399,N_3524,N_1006);
nor U8400 (N_8400,N_1303,N_3334);
or U8401 (N_8401,N_4230,N_3221);
or U8402 (N_8402,N_4082,N_3343);
nor U8403 (N_8403,N_297,N_1493);
xor U8404 (N_8404,N_730,N_2410);
nor U8405 (N_8405,N_843,N_1294);
and U8406 (N_8406,N_1108,N_4153);
xnor U8407 (N_8407,N_2786,N_4734);
or U8408 (N_8408,N_4583,N_669);
xnor U8409 (N_8409,N_615,N_4391);
xnor U8410 (N_8410,N_3243,N_1814);
and U8411 (N_8411,N_1954,N_2514);
and U8412 (N_8412,N_3133,N_693);
nand U8413 (N_8413,N_4170,N_3371);
xor U8414 (N_8414,N_1559,N_2237);
or U8415 (N_8415,N_1643,N_3806);
xor U8416 (N_8416,N_2484,N_578);
nand U8417 (N_8417,N_2483,N_2099);
nand U8418 (N_8418,N_4664,N_2906);
nor U8419 (N_8419,N_2314,N_1289);
xor U8420 (N_8420,N_3675,N_1382);
xor U8421 (N_8421,N_363,N_12);
or U8422 (N_8422,N_537,N_1199);
or U8423 (N_8423,N_3949,N_934);
and U8424 (N_8424,N_1842,N_4222);
nand U8425 (N_8425,N_3315,N_3811);
and U8426 (N_8426,N_620,N_3162);
or U8427 (N_8427,N_1717,N_4900);
nand U8428 (N_8428,N_1038,N_3030);
nor U8429 (N_8429,N_3504,N_1975);
or U8430 (N_8430,N_2757,N_4979);
nand U8431 (N_8431,N_1589,N_1789);
xor U8432 (N_8432,N_1928,N_4197);
nor U8433 (N_8433,N_254,N_2466);
and U8434 (N_8434,N_3310,N_670);
xor U8435 (N_8435,N_2552,N_2581);
xor U8436 (N_8436,N_2737,N_3960);
xor U8437 (N_8437,N_191,N_4845);
nand U8438 (N_8438,N_2479,N_3984);
xor U8439 (N_8439,N_1440,N_3319);
xor U8440 (N_8440,N_1537,N_2735);
and U8441 (N_8441,N_2171,N_831);
or U8442 (N_8442,N_843,N_1150);
nand U8443 (N_8443,N_2460,N_761);
nand U8444 (N_8444,N_3594,N_4357);
xor U8445 (N_8445,N_1756,N_1411);
nor U8446 (N_8446,N_3561,N_3714);
nor U8447 (N_8447,N_2265,N_1122);
nor U8448 (N_8448,N_1262,N_519);
nand U8449 (N_8449,N_2207,N_1196);
xnor U8450 (N_8450,N_3635,N_4420);
xnor U8451 (N_8451,N_2888,N_3200);
nor U8452 (N_8452,N_4267,N_2398);
and U8453 (N_8453,N_1331,N_2902);
or U8454 (N_8454,N_1460,N_1209);
xnor U8455 (N_8455,N_4010,N_4784);
nor U8456 (N_8456,N_3722,N_2762);
xor U8457 (N_8457,N_1152,N_22);
and U8458 (N_8458,N_3052,N_4916);
and U8459 (N_8459,N_171,N_2860);
or U8460 (N_8460,N_138,N_718);
nor U8461 (N_8461,N_1894,N_1339);
nand U8462 (N_8462,N_230,N_4566);
or U8463 (N_8463,N_3480,N_2445);
xnor U8464 (N_8464,N_4427,N_1882);
nand U8465 (N_8465,N_3002,N_321);
nor U8466 (N_8466,N_1339,N_2309);
nor U8467 (N_8467,N_618,N_3218);
and U8468 (N_8468,N_1533,N_1879);
xor U8469 (N_8469,N_698,N_281);
xnor U8470 (N_8470,N_4524,N_3131);
or U8471 (N_8471,N_4473,N_4381);
and U8472 (N_8472,N_2489,N_2825);
nand U8473 (N_8473,N_3220,N_3120);
or U8474 (N_8474,N_3528,N_1185);
nand U8475 (N_8475,N_2725,N_4123);
nor U8476 (N_8476,N_3073,N_4278);
and U8477 (N_8477,N_1723,N_575);
nand U8478 (N_8478,N_2711,N_1585);
nor U8479 (N_8479,N_3114,N_4739);
nand U8480 (N_8480,N_1997,N_2243);
or U8481 (N_8481,N_3995,N_743);
and U8482 (N_8482,N_3199,N_2294);
or U8483 (N_8483,N_4104,N_3887);
or U8484 (N_8484,N_4276,N_934);
xnor U8485 (N_8485,N_160,N_1628);
or U8486 (N_8486,N_4240,N_4825);
nand U8487 (N_8487,N_3783,N_1792);
nor U8488 (N_8488,N_4787,N_1609);
nor U8489 (N_8489,N_3076,N_3325);
nand U8490 (N_8490,N_1007,N_1809);
nand U8491 (N_8491,N_657,N_4769);
xor U8492 (N_8492,N_4172,N_1126);
xor U8493 (N_8493,N_814,N_2235);
nand U8494 (N_8494,N_4768,N_2857);
xnor U8495 (N_8495,N_731,N_146);
nor U8496 (N_8496,N_3946,N_782);
or U8497 (N_8497,N_1139,N_4156);
and U8498 (N_8498,N_508,N_2528);
xnor U8499 (N_8499,N_2704,N_1422);
xnor U8500 (N_8500,N_1457,N_669);
xnor U8501 (N_8501,N_2967,N_872);
nor U8502 (N_8502,N_1268,N_4841);
nand U8503 (N_8503,N_1999,N_4253);
xor U8504 (N_8504,N_2479,N_588);
nor U8505 (N_8505,N_2242,N_87);
nor U8506 (N_8506,N_3530,N_664);
or U8507 (N_8507,N_3482,N_1642);
or U8508 (N_8508,N_268,N_4634);
nor U8509 (N_8509,N_3635,N_3044);
nand U8510 (N_8510,N_4969,N_643);
and U8511 (N_8511,N_845,N_4570);
and U8512 (N_8512,N_167,N_4239);
or U8513 (N_8513,N_1741,N_3006);
nand U8514 (N_8514,N_885,N_2363);
nand U8515 (N_8515,N_2677,N_1740);
and U8516 (N_8516,N_78,N_2732);
xnor U8517 (N_8517,N_1055,N_1843);
or U8518 (N_8518,N_2772,N_3144);
and U8519 (N_8519,N_1418,N_482);
nor U8520 (N_8520,N_1224,N_161);
nor U8521 (N_8521,N_627,N_2148);
xnor U8522 (N_8522,N_4796,N_956);
nor U8523 (N_8523,N_4330,N_113);
or U8524 (N_8524,N_1540,N_1951);
xnor U8525 (N_8525,N_861,N_1082);
and U8526 (N_8526,N_39,N_1924);
or U8527 (N_8527,N_1477,N_1302);
or U8528 (N_8528,N_3827,N_1370);
or U8529 (N_8529,N_201,N_474);
and U8530 (N_8530,N_3571,N_940);
and U8531 (N_8531,N_1105,N_4015);
and U8532 (N_8532,N_1913,N_2198);
nor U8533 (N_8533,N_3877,N_2650);
and U8534 (N_8534,N_2390,N_3037);
xnor U8535 (N_8535,N_2061,N_3821);
nand U8536 (N_8536,N_3470,N_500);
nor U8537 (N_8537,N_2207,N_2940);
nor U8538 (N_8538,N_4915,N_316);
or U8539 (N_8539,N_2367,N_3595);
xnor U8540 (N_8540,N_1280,N_1892);
and U8541 (N_8541,N_102,N_1397);
nor U8542 (N_8542,N_2840,N_1563);
xor U8543 (N_8543,N_2168,N_1910);
or U8544 (N_8544,N_3032,N_4085);
nand U8545 (N_8545,N_4718,N_352);
and U8546 (N_8546,N_610,N_1204);
or U8547 (N_8547,N_1544,N_2356);
or U8548 (N_8548,N_1220,N_2145);
or U8549 (N_8549,N_3621,N_4166);
or U8550 (N_8550,N_2432,N_577);
xor U8551 (N_8551,N_891,N_1797);
nand U8552 (N_8552,N_165,N_4691);
nor U8553 (N_8553,N_3815,N_2538);
or U8554 (N_8554,N_2252,N_265);
or U8555 (N_8555,N_336,N_4984);
nand U8556 (N_8556,N_4973,N_2663);
nand U8557 (N_8557,N_3759,N_2686);
or U8558 (N_8558,N_4417,N_3401);
nand U8559 (N_8559,N_625,N_75);
nor U8560 (N_8560,N_4743,N_349);
nor U8561 (N_8561,N_3037,N_4660);
and U8562 (N_8562,N_4684,N_4719);
or U8563 (N_8563,N_2911,N_2727);
or U8564 (N_8564,N_1168,N_3354);
xor U8565 (N_8565,N_1995,N_2437);
nor U8566 (N_8566,N_233,N_2232);
or U8567 (N_8567,N_1660,N_2915);
or U8568 (N_8568,N_4679,N_4293);
nand U8569 (N_8569,N_2547,N_126);
nor U8570 (N_8570,N_3309,N_3848);
or U8571 (N_8571,N_2659,N_4457);
and U8572 (N_8572,N_605,N_1916);
or U8573 (N_8573,N_4385,N_3750);
and U8574 (N_8574,N_2193,N_2663);
and U8575 (N_8575,N_728,N_3809);
nand U8576 (N_8576,N_372,N_4080);
or U8577 (N_8577,N_308,N_798);
nand U8578 (N_8578,N_4700,N_1850);
nand U8579 (N_8579,N_4158,N_3807);
nand U8580 (N_8580,N_2324,N_4272);
and U8581 (N_8581,N_2702,N_3007);
xnor U8582 (N_8582,N_2975,N_4678);
or U8583 (N_8583,N_2954,N_2609);
or U8584 (N_8584,N_3647,N_4220);
nor U8585 (N_8585,N_2914,N_4393);
or U8586 (N_8586,N_4548,N_2720);
nand U8587 (N_8587,N_3409,N_3760);
xnor U8588 (N_8588,N_469,N_1267);
and U8589 (N_8589,N_2035,N_638);
xor U8590 (N_8590,N_3439,N_2970);
nor U8591 (N_8591,N_4052,N_2701);
and U8592 (N_8592,N_4843,N_3311);
nor U8593 (N_8593,N_3679,N_836);
nor U8594 (N_8594,N_2771,N_619);
and U8595 (N_8595,N_3755,N_2567);
xor U8596 (N_8596,N_780,N_984);
nor U8597 (N_8597,N_1535,N_2170);
nor U8598 (N_8598,N_3700,N_615);
nand U8599 (N_8599,N_1046,N_4437);
and U8600 (N_8600,N_4563,N_4833);
nand U8601 (N_8601,N_4493,N_1911);
or U8602 (N_8602,N_2885,N_2514);
xnor U8603 (N_8603,N_2445,N_2547);
nand U8604 (N_8604,N_448,N_3743);
or U8605 (N_8605,N_2884,N_4633);
nand U8606 (N_8606,N_3165,N_129);
and U8607 (N_8607,N_963,N_1902);
or U8608 (N_8608,N_710,N_421);
nand U8609 (N_8609,N_1576,N_4954);
and U8610 (N_8610,N_1774,N_3087);
and U8611 (N_8611,N_4073,N_4992);
nand U8612 (N_8612,N_731,N_3917);
nand U8613 (N_8613,N_2778,N_4702);
nor U8614 (N_8614,N_1945,N_3970);
or U8615 (N_8615,N_4036,N_2673);
xor U8616 (N_8616,N_1125,N_596);
nand U8617 (N_8617,N_424,N_4552);
nand U8618 (N_8618,N_308,N_472);
nor U8619 (N_8619,N_2600,N_928);
and U8620 (N_8620,N_1875,N_4317);
nand U8621 (N_8621,N_3468,N_1182);
or U8622 (N_8622,N_2168,N_3836);
nand U8623 (N_8623,N_2496,N_2240);
or U8624 (N_8624,N_3560,N_3180);
nand U8625 (N_8625,N_851,N_4085);
nor U8626 (N_8626,N_3509,N_3913);
nor U8627 (N_8627,N_4997,N_4835);
and U8628 (N_8628,N_4585,N_2679);
nor U8629 (N_8629,N_4810,N_3509);
nand U8630 (N_8630,N_598,N_2587);
nand U8631 (N_8631,N_1335,N_950);
nand U8632 (N_8632,N_1167,N_4173);
or U8633 (N_8633,N_2840,N_3149);
nor U8634 (N_8634,N_1719,N_408);
or U8635 (N_8635,N_1677,N_4334);
xnor U8636 (N_8636,N_1387,N_1918);
xor U8637 (N_8637,N_2279,N_145);
or U8638 (N_8638,N_685,N_304);
nand U8639 (N_8639,N_3943,N_843);
or U8640 (N_8640,N_1650,N_2587);
nand U8641 (N_8641,N_1031,N_1742);
and U8642 (N_8642,N_2394,N_946);
nand U8643 (N_8643,N_1204,N_1696);
nand U8644 (N_8644,N_23,N_4249);
xnor U8645 (N_8645,N_2123,N_1223);
nor U8646 (N_8646,N_78,N_3518);
nand U8647 (N_8647,N_149,N_4308);
nand U8648 (N_8648,N_4017,N_2110);
or U8649 (N_8649,N_2339,N_788);
or U8650 (N_8650,N_2933,N_2071);
xor U8651 (N_8651,N_858,N_3190);
and U8652 (N_8652,N_1209,N_495);
nand U8653 (N_8653,N_2943,N_1290);
xor U8654 (N_8654,N_2914,N_2890);
nor U8655 (N_8655,N_4064,N_567);
xor U8656 (N_8656,N_2741,N_3684);
xor U8657 (N_8657,N_4064,N_3651);
or U8658 (N_8658,N_1824,N_4853);
nor U8659 (N_8659,N_1755,N_4663);
nor U8660 (N_8660,N_4903,N_4592);
or U8661 (N_8661,N_918,N_171);
or U8662 (N_8662,N_889,N_814);
or U8663 (N_8663,N_1683,N_4164);
or U8664 (N_8664,N_1215,N_2492);
nand U8665 (N_8665,N_3383,N_2594);
or U8666 (N_8666,N_1473,N_4072);
nor U8667 (N_8667,N_2199,N_1053);
xnor U8668 (N_8668,N_1601,N_2018);
or U8669 (N_8669,N_968,N_1504);
and U8670 (N_8670,N_2995,N_1078);
xnor U8671 (N_8671,N_2838,N_3355);
and U8672 (N_8672,N_3270,N_2732);
or U8673 (N_8673,N_171,N_3808);
nand U8674 (N_8674,N_1783,N_3405);
or U8675 (N_8675,N_3496,N_3909);
nand U8676 (N_8676,N_839,N_4097);
nor U8677 (N_8677,N_4834,N_2569);
and U8678 (N_8678,N_1449,N_804);
xor U8679 (N_8679,N_2021,N_3483);
xor U8680 (N_8680,N_1083,N_2430);
or U8681 (N_8681,N_231,N_4752);
or U8682 (N_8682,N_1643,N_2728);
and U8683 (N_8683,N_2467,N_1952);
and U8684 (N_8684,N_725,N_4786);
xnor U8685 (N_8685,N_4496,N_4745);
nor U8686 (N_8686,N_3191,N_890);
and U8687 (N_8687,N_542,N_4304);
and U8688 (N_8688,N_1726,N_3533);
and U8689 (N_8689,N_2966,N_4949);
and U8690 (N_8690,N_3094,N_1383);
nor U8691 (N_8691,N_1392,N_2629);
xor U8692 (N_8692,N_3809,N_2977);
xor U8693 (N_8693,N_1333,N_900);
xor U8694 (N_8694,N_1156,N_1032);
nor U8695 (N_8695,N_1902,N_4246);
nor U8696 (N_8696,N_3971,N_1638);
and U8697 (N_8697,N_1512,N_2989);
and U8698 (N_8698,N_1464,N_4279);
xnor U8699 (N_8699,N_3438,N_4407);
nand U8700 (N_8700,N_3992,N_4913);
and U8701 (N_8701,N_2159,N_2137);
and U8702 (N_8702,N_1196,N_3620);
nand U8703 (N_8703,N_3771,N_3185);
or U8704 (N_8704,N_1077,N_4487);
xnor U8705 (N_8705,N_362,N_3384);
xor U8706 (N_8706,N_1533,N_460);
xor U8707 (N_8707,N_4958,N_1710);
or U8708 (N_8708,N_2672,N_3613);
or U8709 (N_8709,N_1026,N_2807);
xor U8710 (N_8710,N_229,N_1033);
xnor U8711 (N_8711,N_2511,N_2497);
and U8712 (N_8712,N_4858,N_218);
nor U8713 (N_8713,N_3488,N_3141);
and U8714 (N_8714,N_2033,N_542);
or U8715 (N_8715,N_3337,N_1234);
and U8716 (N_8716,N_1629,N_4105);
or U8717 (N_8717,N_1689,N_1124);
nor U8718 (N_8718,N_4105,N_4328);
xor U8719 (N_8719,N_4372,N_248);
nor U8720 (N_8720,N_147,N_4250);
or U8721 (N_8721,N_1616,N_155);
xor U8722 (N_8722,N_298,N_1476);
nand U8723 (N_8723,N_4891,N_1647);
nand U8724 (N_8724,N_2787,N_1969);
or U8725 (N_8725,N_210,N_3165);
xor U8726 (N_8726,N_1555,N_2725);
nand U8727 (N_8727,N_1222,N_177);
or U8728 (N_8728,N_1759,N_4145);
or U8729 (N_8729,N_2670,N_4595);
xnor U8730 (N_8730,N_4631,N_944);
or U8731 (N_8731,N_4274,N_945);
xnor U8732 (N_8732,N_2498,N_3595);
or U8733 (N_8733,N_701,N_551);
nor U8734 (N_8734,N_892,N_4750);
nor U8735 (N_8735,N_519,N_237);
nor U8736 (N_8736,N_3694,N_1293);
xnor U8737 (N_8737,N_3938,N_2602);
or U8738 (N_8738,N_425,N_3117);
or U8739 (N_8739,N_1489,N_622);
and U8740 (N_8740,N_2962,N_1751);
nor U8741 (N_8741,N_2906,N_4176);
xnor U8742 (N_8742,N_404,N_4662);
nand U8743 (N_8743,N_4404,N_1946);
xor U8744 (N_8744,N_865,N_42);
nand U8745 (N_8745,N_1981,N_621);
nor U8746 (N_8746,N_3428,N_1013);
nand U8747 (N_8747,N_4884,N_203);
nand U8748 (N_8748,N_929,N_4875);
xnor U8749 (N_8749,N_1591,N_2415);
nor U8750 (N_8750,N_1913,N_2650);
nor U8751 (N_8751,N_3876,N_2444);
xor U8752 (N_8752,N_1515,N_927);
nand U8753 (N_8753,N_4019,N_4811);
or U8754 (N_8754,N_4736,N_4119);
xor U8755 (N_8755,N_3212,N_1231);
nor U8756 (N_8756,N_2943,N_4856);
and U8757 (N_8757,N_4668,N_191);
nor U8758 (N_8758,N_1955,N_2806);
and U8759 (N_8759,N_4837,N_170);
nor U8760 (N_8760,N_1007,N_2114);
or U8761 (N_8761,N_4683,N_2925);
or U8762 (N_8762,N_3544,N_1350);
xor U8763 (N_8763,N_4032,N_3711);
xor U8764 (N_8764,N_2890,N_62);
nand U8765 (N_8765,N_1703,N_918);
xnor U8766 (N_8766,N_4926,N_3374);
and U8767 (N_8767,N_4250,N_2293);
or U8768 (N_8768,N_3782,N_2036);
and U8769 (N_8769,N_1153,N_4942);
xor U8770 (N_8770,N_4369,N_3716);
or U8771 (N_8771,N_3760,N_1741);
nand U8772 (N_8772,N_2016,N_3345);
xnor U8773 (N_8773,N_415,N_2088);
nor U8774 (N_8774,N_3406,N_1882);
nand U8775 (N_8775,N_4526,N_2187);
nor U8776 (N_8776,N_1106,N_4267);
nor U8777 (N_8777,N_3366,N_205);
nor U8778 (N_8778,N_4046,N_3503);
xor U8779 (N_8779,N_398,N_295);
xor U8780 (N_8780,N_4905,N_1080);
nor U8781 (N_8781,N_4623,N_4829);
and U8782 (N_8782,N_3063,N_66);
xnor U8783 (N_8783,N_1535,N_2998);
and U8784 (N_8784,N_1713,N_1833);
nor U8785 (N_8785,N_671,N_2140);
nor U8786 (N_8786,N_3119,N_382);
xor U8787 (N_8787,N_1484,N_1141);
or U8788 (N_8788,N_3995,N_4318);
xnor U8789 (N_8789,N_1128,N_332);
nand U8790 (N_8790,N_4766,N_4412);
nand U8791 (N_8791,N_1780,N_3291);
nand U8792 (N_8792,N_2369,N_3074);
nand U8793 (N_8793,N_423,N_4594);
nand U8794 (N_8794,N_2707,N_3976);
xnor U8795 (N_8795,N_3312,N_4596);
or U8796 (N_8796,N_2216,N_1808);
xor U8797 (N_8797,N_171,N_3288);
nor U8798 (N_8798,N_1632,N_707);
and U8799 (N_8799,N_2828,N_4373);
nand U8800 (N_8800,N_3727,N_1460);
xnor U8801 (N_8801,N_2648,N_415);
or U8802 (N_8802,N_3416,N_2297);
xor U8803 (N_8803,N_2550,N_3964);
and U8804 (N_8804,N_1488,N_2393);
xor U8805 (N_8805,N_2705,N_2769);
nor U8806 (N_8806,N_2557,N_4515);
nand U8807 (N_8807,N_2329,N_1529);
and U8808 (N_8808,N_2874,N_894);
xnor U8809 (N_8809,N_3941,N_1877);
xnor U8810 (N_8810,N_617,N_3592);
nor U8811 (N_8811,N_2207,N_2814);
or U8812 (N_8812,N_3291,N_2270);
and U8813 (N_8813,N_3669,N_2419);
or U8814 (N_8814,N_3517,N_4228);
nor U8815 (N_8815,N_1559,N_2805);
and U8816 (N_8816,N_2323,N_4000);
nand U8817 (N_8817,N_4821,N_3974);
xnor U8818 (N_8818,N_3247,N_2019);
or U8819 (N_8819,N_1481,N_4459);
or U8820 (N_8820,N_806,N_1324);
or U8821 (N_8821,N_936,N_4821);
xor U8822 (N_8822,N_4148,N_4192);
nor U8823 (N_8823,N_2000,N_4599);
or U8824 (N_8824,N_979,N_3483);
xor U8825 (N_8825,N_4443,N_3984);
nor U8826 (N_8826,N_1983,N_2039);
xor U8827 (N_8827,N_21,N_1919);
nor U8828 (N_8828,N_971,N_3995);
nor U8829 (N_8829,N_4644,N_1242);
nand U8830 (N_8830,N_1648,N_4168);
xor U8831 (N_8831,N_1727,N_163);
nand U8832 (N_8832,N_2479,N_2285);
nor U8833 (N_8833,N_4703,N_4104);
or U8834 (N_8834,N_2780,N_4964);
xor U8835 (N_8835,N_4878,N_1908);
xnor U8836 (N_8836,N_919,N_2825);
and U8837 (N_8837,N_4146,N_2647);
xnor U8838 (N_8838,N_189,N_3399);
or U8839 (N_8839,N_1598,N_1005);
or U8840 (N_8840,N_3843,N_585);
nor U8841 (N_8841,N_413,N_556);
nand U8842 (N_8842,N_502,N_1189);
nor U8843 (N_8843,N_4863,N_388);
nor U8844 (N_8844,N_1935,N_278);
xor U8845 (N_8845,N_1665,N_2635);
or U8846 (N_8846,N_4571,N_1833);
nand U8847 (N_8847,N_1660,N_3914);
and U8848 (N_8848,N_874,N_4775);
xnor U8849 (N_8849,N_1310,N_1471);
or U8850 (N_8850,N_1450,N_3488);
nand U8851 (N_8851,N_3679,N_4834);
or U8852 (N_8852,N_1575,N_1230);
xnor U8853 (N_8853,N_4761,N_60);
nor U8854 (N_8854,N_4206,N_827);
nor U8855 (N_8855,N_4077,N_1435);
or U8856 (N_8856,N_3896,N_3217);
nand U8857 (N_8857,N_2004,N_1974);
xnor U8858 (N_8858,N_3671,N_4685);
nand U8859 (N_8859,N_1177,N_633);
nor U8860 (N_8860,N_4116,N_4903);
or U8861 (N_8861,N_1913,N_714);
and U8862 (N_8862,N_4102,N_4190);
nor U8863 (N_8863,N_2323,N_1025);
nand U8864 (N_8864,N_4894,N_2657);
and U8865 (N_8865,N_872,N_4595);
or U8866 (N_8866,N_4714,N_544);
xnor U8867 (N_8867,N_1958,N_4379);
nor U8868 (N_8868,N_1119,N_2218);
nand U8869 (N_8869,N_3623,N_1709);
and U8870 (N_8870,N_2308,N_1945);
or U8871 (N_8871,N_2067,N_4588);
nor U8872 (N_8872,N_2105,N_3062);
or U8873 (N_8873,N_343,N_3791);
and U8874 (N_8874,N_2414,N_2257);
and U8875 (N_8875,N_2243,N_1505);
nand U8876 (N_8876,N_3526,N_1909);
nand U8877 (N_8877,N_2932,N_3141);
nor U8878 (N_8878,N_2597,N_3483);
and U8879 (N_8879,N_2490,N_2883);
and U8880 (N_8880,N_701,N_2008);
or U8881 (N_8881,N_1910,N_230);
and U8882 (N_8882,N_389,N_4546);
xnor U8883 (N_8883,N_2490,N_1026);
nor U8884 (N_8884,N_2617,N_1933);
and U8885 (N_8885,N_1715,N_4355);
and U8886 (N_8886,N_2322,N_2577);
and U8887 (N_8887,N_35,N_2771);
xnor U8888 (N_8888,N_1331,N_3710);
or U8889 (N_8889,N_815,N_4012);
or U8890 (N_8890,N_3791,N_4467);
and U8891 (N_8891,N_2771,N_1238);
and U8892 (N_8892,N_1146,N_3969);
or U8893 (N_8893,N_279,N_4265);
xor U8894 (N_8894,N_1802,N_4753);
nor U8895 (N_8895,N_3467,N_3446);
and U8896 (N_8896,N_2256,N_2310);
xnor U8897 (N_8897,N_4899,N_2768);
xnor U8898 (N_8898,N_2416,N_3627);
xnor U8899 (N_8899,N_509,N_3039);
xnor U8900 (N_8900,N_4735,N_3105);
xor U8901 (N_8901,N_3918,N_495);
or U8902 (N_8902,N_1994,N_2380);
xor U8903 (N_8903,N_1750,N_4135);
and U8904 (N_8904,N_157,N_4109);
xor U8905 (N_8905,N_2568,N_2088);
xnor U8906 (N_8906,N_333,N_3417);
and U8907 (N_8907,N_1890,N_2416);
nand U8908 (N_8908,N_4730,N_2094);
nand U8909 (N_8909,N_4398,N_3679);
nand U8910 (N_8910,N_4707,N_4582);
and U8911 (N_8911,N_1829,N_2578);
nand U8912 (N_8912,N_3632,N_983);
nand U8913 (N_8913,N_696,N_4019);
nor U8914 (N_8914,N_1688,N_482);
nor U8915 (N_8915,N_2675,N_2497);
or U8916 (N_8916,N_825,N_949);
or U8917 (N_8917,N_3590,N_3352);
or U8918 (N_8918,N_2297,N_625);
and U8919 (N_8919,N_3607,N_4831);
and U8920 (N_8920,N_894,N_587);
nor U8921 (N_8921,N_4064,N_1596);
nor U8922 (N_8922,N_2963,N_4643);
or U8923 (N_8923,N_2529,N_4571);
xor U8924 (N_8924,N_1405,N_425);
or U8925 (N_8925,N_4973,N_4318);
nand U8926 (N_8926,N_2651,N_2579);
nand U8927 (N_8927,N_2471,N_4397);
nand U8928 (N_8928,N_3423,N_3072);
nor U8929 (N_8929,N_2775,N_3783);
nor U8930 (N_8930,N_1572,N_4081);
and U8931 (N_8931,N_4908,N_4439);
nor U8932 (N_8932,N_3872,N_4451);
and U8933 (N_8933,N_3319,N_4810);
nor U8934 (N_8934,N_1538,N_289);
nand U8935 (N_8935,N_4207,N_773);
or U8936 (N_8936,N_82,N_844);
and U8937 (N_8937,N_4305,N_921);
nor U8938 (N_8938,N_2093,N_615);
or U8939 (N_8939,N_846,N_552);
nor U8940 (N_8940,N_1998,N_4467);
xnor U8941 (N_8941,N_729,N_1846);
xor U8942 (N_8942,N_3685,N_1700);
nor U8943 (N_8943,N_1553,N_4423);
xnor U8944 (N_8944,N_4469,N_1053);
or U8945 (N_8945,N_2206,N_4631);
nand U8946 (N_8946,N_3705,N_2503);
nand U8947 (N_8947,N_927,N_2943);
nor U8948 (N_8948,N_1019,N_4109);
nand U8949 (N_8949,N_3372,N_4543);
or U8950 (N_8950,N_4393,N_2723);
nor U8951 (N_8951,N_2926,N_2453);
or U8952 (N_8952,N_506,N_3618);
and U8953 (N_8953,N_3315,N_488);
nand U8954 (N_8954,N_3556,N_3832);
and U8955 (N_8955,N_2574,N_1216);
and U8956 (N_8956,N_2335,N_132);
nand U8957 (N_8957,N_1285,N_3256);
nor U8958 (N_8958,N_814,N_1861);
or U8959 (N_8959,N_2370,N_4092);
nor U8960 (N_8960,N_1041,N_4058);
nor U8961 (N_8961,N_1971,N_4536);
nand U8962 (N_8962,N_2591,N_208);
xnor U8963 (N_8963,N_3643,N_2675);
nor U8964 (N_8964,N_3969,N_591);
or U8965 (N_8965,N_969,N_1371);
and U8966 (N_8966,N_4863,N_4475);
or U8967 (N_8967,N_2821,N_4313);
nand U8968 (N_8968,N_2020,N_4950);
xor U8969 (N_8969,N_2453,N_0);
and U8970 (N_8970,N_4896,N_1461);
and U8971 (N_8971,N_834,N_1179);
and U8972 (N_8972,N_3317,N_507);
nand U8973 (N_8973,N_549,N_1407);
nor U8974 (N_8974,N_4891,N_4238);
and U8975 (N_8975,N_926,N_2725);
and U8976 (N_8976,N_1766,N_1904);
nand U8977 (N_8977,N_3069,N_3959);
and U8978 (N_8978,N_4671,N_4024);
xnor U8979 (N_8979,N_3865,N_2256);
or U8980 (N_8980,N_2086,N_3304);
nand U8981 (N_8981,N_3940,N_2537);
xnor U8982 (N_8982,N_4766,N_2213);
or U8983 (N_8983,N_4423,N_4976);
nand U8984 (N_8984,N_3002,N_933);
xor U8985 (N_8985,N_1376,N_1467);
or U8986 (N_8986,N_2218,N_3054);
nor U8987 (N_8987,N_1916,N_2978);
nor U8988 (N_8988,N_1966,N_2658);
nand U8989 (N_8989,N_2259,N_1259);
nor U8990 (N_8990,N_32,N_156);
xor U8991 (N_8991,N_1292,N_2327);
and U8992 (N_8992,N_938,N_1964);
xor U8993 (N_8993,N_319,N_1359);
and U8994 (N_8994,N_594,N_4079);
nor U8995 (N_8995,N_1008,N_4110);
nand U8996 (N_8996,N_1006,N_2752);
and U8997 (N_8997,N_4248,N_4892);
nor U8998 (N_8998,N_480,N_522);
and U8999 (N_8999,N_4933,N_3829);
nor U9000 (N_9000,N_2409,N_2052);
nand U9001 (N_9001,N_4303,N_2026);
and U9002 (N_9002,N_1360,N_234);
and U9003 (N_9003,N_4446,N_552);
or U9004 (N_9004,N_3418,N_3958);
xnor U9005 (N_9005,N_3632,N_3355);
nand U9006 (N_9006,N_3478,N_4164);
nand U9007 (N_9007,N_2469,N_3603);
xor U9008 (N_9008,N_1131,N_4649);
and U9009 (N_9009,N_1726,N_1350);
or U9010 (N_9010,N_3925,N_2850);
nand U9011 (N_9011,N_3888,N_1270);
nor U9012 (N_9012,N_278,N_1846);
xnor U9013 (N_9013,N_274,N_3663);
and U9014 (N_9014,N_1217,N_176);
nor U9015 (N_9015,N_3659,N_2090);
or U9016 (N_9016,N_834,N_2591);
nor U9017 (N_9017,N_4242,N_3066);
or U9018 (N_9018,N_3782,N_3508);
and U9019 (N_9019,N_2182,N_574);
or U9020 (N_9020,N_75,N_1017);
or U9021 (N_9021,N_4643,N_3508);
or U9022 (N_9022,N_913,N_4118);
and U9023 (N_9023,N_1385,N_468);
nand U9024 (N_9024,N_1505,N_2275);
nor U9025 (N_9025,N_2075,N_350);
nor U9026 (N_9026,N_3481,N_850);
xor U9027 (N_9027,N_862,N_503);
xor U9028 (N_9028,N_3644,N_1298);
nor U9029 (N_9029,N_3393,N_756);
nand U9030 (N_9030,N_3842,N_2124);
and U9031 (N_9031,N_4609,N_3258);
xnor U9032 (N_9032,N_4834,N_3339);
and U9033 (N_9033,N_2051,N_4218);
nand U9034 (N_9034,N_226,N_207);
nand U9035 (N_9035,N_3697,N_4988);
and U9036 (N_9036,N_4604,N_2969);
or U9037 (N_9037,N_4432,N_4272);
and U9038 (N_9038,N_4223,N_3440);
nand U9039 (N_9039,N_3770,N_3758);
nor U9040 (N_9040,N_3270,N_3367);
nand U9041 (N_9041,N_4796,N_2827);
or U9042 (N_9042,N_3552,N_146);
nor U9043 (N_9043,N_4981,N_353);
xor U9044 (N_9044,N_4502,N_3581);
and U9045 (N_9045,N_3442,N_761);
xor U9046 (N_9046,N_4105,N_1776);
and U9047 (N_9047,N_2807,N_1175);
nor U9048 (N_9048,N_4439,N_4592);
nand U9049 (N_9049,N_1400,N_2734);
and U9050 (N_9050,N_1751,N_2404);
or U9051 (N_9051,N_3298,N_706);
or U9052 (N_9052,N_301,N_1183);
nor U9053 (N_9053,N_4331,N_23);
nand U9054 (N_9054,N_1164,N_3387);
nand U9055 (N_9055,N_2610,N_1569);
and U9056 (N_9056,N_4705,N_340);
and U9057 (N_9057,N_3118,N_4962);
nor U9058 (N_9058,N_678,N_961);
nand U9059 (N_9059,N_1705,N_3955);
xnor U9060 (N_9060,N_1105,N_3147);
nor U9061 (N_9061,N_1976,N_4090);
nor U9062 (N_9062,N_3892,N_3376);
or U9063 (N_9063,N_156,N_1865);
or U9064 (N_9064,N_1541,N_1843);
or U9065 (N_9065,N_2097,N_444);
and U9066 (N_9066,N_35,N_2005);
nor U9067 (N_9067,N_2029,N_1357);
nor U9068 (N_9068,N_1963,N_1263);
and U9069 (N_9069,N_3757,N_3545);
or U9070 (N_9070,N_3024,N_1592);
nor U9071 (N_9071,N_2484,N_2828);
or U9072 (N_9072,N_4373,N_1228);
nand U9073 (N_9073,N_1983,N_4890);
xor U9074 (N_9074,N_620,N_2037);
and U9075 (N_9075,N_834,N_4024);
nand U9076 (N_9076,N_562,N_279);
nand U9077 (N_9077,N_1167,N_3380);
or U9078 (N_9078,N_2770,N_3438);
or U9079 (N_9079,N_2624,N_68);
and U9080 (N_9080,N_682,N_2106);
xnor U9081 (N_9081,N_3933,N_449);
and U9082 (N_9082,N_2697,N_4303);
or U9083 (N_9083,N_880,N_2931);
nor U9084 (N_9084,N_4743,N_3097);
or U9085 (N_9085,N_192,N_441);
and U9086 (N_9086,N_1923,N_353);
xnor U9087 (N_9087,N_4008,N_3952);
nand U9088 (N_9088,N_3512,N_4087);
and U9089 (N_9089,N_3684,N_4190);
or U9090 (N_9090,N_1622,N_2996);
nand U9091 (N_9091,N_3039,N_4038);
xnor U9092 (N_9092,N_4470,N_4664);
nor U9093 (N_9093,N_3820,N_383);
nand U9094 (N_9094,N_418,N_2038);
nand U9095 (N_9095,N_1316,N_2717);
nor U9096 (N_9096,N_1644,N_1769);
nand U9097 (N_9097,N_1575,N_3765);
and U9098 (N_9098,N_2882,N_4844);
or U9099 (N_9099,N_2832,N_4733);
nor U9100 (N_9100,N_2760,N_1370);
and U9101 (N_9101,N_3657,N_1599);
and U9102 (N_9102,N_197,N_759);
xnor U9103 (N_9103,N_492,N_3200);
and U9104 (N_9104,N_2695,N_4433);
or U9105 (N_9105,N_4508,N_3283);
nand U9106 (N_9106,N_4285,N_2489);
and U9107 (N_9107,N_4559,N_4687);
and U9108 (N_9108,N_1528,N_2445);
nand U9109 (N_9109,N_3383,N_2098);
xor U9110 (N_9110,N_4057,N_360);
or U9111 (N_9111,N_2004,N_4123);
and U9112 (N_9112,N_283,N_4790);
and U9113 (N_9113,N_2891,N_4682);
nand U9114 (N_9114,N_2715,N_4858);
nand U9115 (N_9115,N_1670,N_861);
or U9116 (N_9116,N_4664,N_3541);
nand U9117 (N_9117,N_4883,N_791);
nor U9118 (N_9118,N_4123,N_845);
nor U9119 (N_9119,N_2584,N_1596);
or U9120 (N_9120,N_2590,N_3389);
xor U9121 (N_9121,N_14,N_4810);
and U9122 (N_9122,N_3211,N_2965);
and U9123 (N_9123,N_4373,N_4314);
and U9124 (N_9124,N_900,N_3147);
and U9125 (N_9125,N_1298,N_2096);
and U9126 (N_9126,N_387,N_3512);
nor U9127 (N_9127,N_3181,N_1472);
nor U9128 (N_9128,N_4024,N_2019);
xor U9129 (N_9129,N_1833,N_2272);
xnor U9130 (N_9130,N_3857,N_4933);
and U9131 (N_9131,N_4582,N_1716);
nand U9132 (N_9132,N_2496,N_269);
nand U9133 (N_9133,N_4020,N_3819);
and U9134 (N_9134,N_3439,N_3822);
xnor U9135 (N_9135,N_1362,N_1887);
nand U9136 (N_9136,N_630,N_1312);
or U9137 (N_9137,N_3030,N_2248);
or U9138 (N_9138,N_784,N_4033);
nor U9139 (N_9139,N_117,N_1398);
xnor U9140 (N_9140,N_2038,N_1028);
nand U9141 (N_9141,N_772,N_1163);
xnor U9142 (N_9142,N_4749,N_198);
xnor U9143 (N_9143,N_2429,N_4877);
xnor U9144 (N_9144,N_338,N_2165);
nor U9145 (N_9145,N_99,N_2832);
nor U9146 (N_9146,N_331,N_2251);
nor U9147 (N_9147,N_4232,N_2076);
nand U9148 (N_9148,N_2425,N_1700);
or U9149 (N_9149,N_2762,N_2784);
and U9150 (N_9150,N_3998,N_3538);
nand U9151 (N_9151,N_3641,N_4999);
nand U9152 (N_9152,N_3344,N_3422);
nand U9153 (N_9153,N_3285,N_1295);
and U9154 (N_9154,N_652,N_1224);
or U9155 (N_9155,N_4603,N_889);
nand U9156 (N_9156,N_3607,N_224);
and U9157 (N_9157,N_3738,N_2778);
or U9158 (N_9158,N_2435,N_1351);
nand U9159 (N_9159,N_1938,N_3957);
nand U9160 (N_9160,N_3086,N_1410);
nor U9161 (N_9161,N_1212,N_4156);
xnor U9162 (N_9162,N_3413,N_4337);
nand U9163 (N_9163,N_3875,N_2067);
or U9164 (N_9164,N_971,N_4812);
xnor U9165 (N_9165,N_3052,N_2602);
and U9166 (N_9166,N_285,N_946);
or U9167 (N_9167,N_769,N_695);
nor U9168 (N_9168,N_2226,N_2696);
or U9169 (N_9169,N_1520,N_1996);
and U9170 (N_9170,N_3611,N_4739);
and U9171 (N_9171,N_3214,N_2448);
and U9172 (N_9172,N_896,N_4087);
nand U9173 (N_9173,N_3546,N_821);
nor U9174 (N_9174,N_4380,N_4946);
or U9175 (N_9175,N_4070,N_3276);
xnor U9176 (N_9176,N_1741,N_2681);
xnor U9177 (N_9177,N_961,N_3842);
xor U9178 (N_9178,N_4041,N_4894);
xnor U9179 (N_9179,N_756,N_1358);
or U9180 (N_9180,N_1381,N_4130);
or U9181 (N_9181,N_162,N_2033);
xnor U9182 (N_9182,N_4444,N_2317);
or U9183 (N_9183,N_314,N_838);
nor U9184 (N_9184,N_1277,N_2824);
nand U9185 (N_9185,N_4471,N_359);
nand U9186 (N_9186,N_3230,N_3001);
nor U9187 (N_9187,N_2541,N_1716);
or U9188 (N_9188,N_2504,N_240);
or U9189 (N_9189,N_1373,N_1417);
xor U9190 (N_9190,N_4695,N_1953);
xnor U9191 (N_9191,N_2666,N_3270);
nand U9192 (N_9192,N_198,N_1230);
and U9193 (N_9193,N_2953,N_1032);
or U9194 (N_9194,N_1632,N_3705);
nand U9195 (N_9195,N_3598,N_1361);
or U9196 (N_9196,N_3863,N_3434);
and U9197 (N_9197,N_1319,N_2243);
nand U9198 (N_9198,N_1389,N_1549);
nand U9199 (N_9199,N_4246,N_3210);
and U9200 (N_9200,N_1663,N_3134);
or U9201 (N_9201,N_433,N_4498);
and U9202 (N_9202,N_667,N_1330);
nor U9203 (N_9203,N_2965,N_1282);
and U9204 (N_9204,N_4718,N_1294);
or U9205 (N_9205,N_1768,N_2183);
nand U9206 (N_9206,N_2489,N_3749);
or U9207 (N_9207,N_810,N_3886);
xor U9208 (N_9208,N_882,N_3636);
xnor U9209 (N_9209,N_1195,N_2379);
and U9210 (N_9210,N_3590,N_4014);
and U9211 (N_9211,N_594,N_3898);
and U9212 (N_9212,N_416,N_607);
xnor U9213 (N_9213,N_2601,N_106);
nor U9214 (N_9214,N_1658,N_2038);
nand U9215 (N_9215,N_1602,N_1054);
xor U9216 (N_9216,N_1737,N_1095);
and U9217 (N_9217,N_1985,N_31);
and U9218 (N_9218,N_186,N_1084);
xnor U9219 (N_9219,N_1283,N_305);
or U9220 (N_9220,N_4401,N_1613);
or U9221 (N_9221,N_3691,N_4858);
or U9222 (N_9222,N_2269,N_3453);
nand U9223 (N_9223,N_2852,N_4969);
and U9224 (N_9224,N_3116,N_1427);
xor U9225 (N_9225,N_1777,N_658);
nor U9226 (N_9226,N_3969,N_2081);
and U9227 (N_9227,N_3065,N_2541);
xnor U9228 (N_9228,N_2953,N_3590);
nor U9229 (N_9229,N_1204,N_4678);
and U9230 (N_9230,N_286,N_2389);
and U9231 (N_9231,N_4223,N_682);
nor U9232 (N_9232,N_818,N_780);
and U9233 (N_9233,N_207,N_676);
or U9234 (N_9234,N_1533,N_18);
nor U9235 (N_9235,N_3275,N_3267);
and U9236 (N_9236,N_3154,N_4384);
nand U9237 (N_9237,N_4836,N_2187);
or U9238 (N_9238,N_4330,N_1134);
nand U9239 (N_9239,N_4366,N_4580);
or U9240 (N_9240,N_4383,N_2487);
nand U9241 (N_9241,N_1663,N_3763);
or U9242 (N_9242,N_2250,N_3863);
nand U9243 (N_9243,N_933,N_1402);
nor U9244 (N_9244,N_1845,N_2250);
nand U9245 (N_9245,N_4645,N_3857);
nand U9246 (N_9246,N_3672,N_2014);
and U9247 (N_9247,N_720,N_4026);
xor U9248 (N_9248,N_2106,N_1669);
nand U9249 (N_9249,N_1450,N_1838);
and U9250 (N_9250,N_3909,N_3162);
and U9251 (N_9251,N_3419,N_4165);
nand U9252 (N_9252,N_3264,N_2592);
xnor U9253 (N_9253,N_2088,N_3915);
nor U9254 (N_9254,N_381,N_1495);
nor U9255 (N_9255,N_3127,N_1543);
or U9256 (N_9256,N_1307,N_3722);
xor U9257 (N_9257,N_235,N_756);
or U9258 (N_9258,N_4879,N_180);
xnor U9259 (N_9259,N_1776,N_75);
xor U9260 (N_9260,N_614,N_916);
nand U9261 (N_9261,N_217,N_2744);
nor U9262 (N_9262,N_262,N_385);
xor U9263 (N_9263,N_3519,N_240);
and U9264 (N_9264,N_392,N_634);
and U9265 (N_9265,N_4246,N_1945);
or U9266 (N_9266,N_2867,N_4041);
nor U9267 (N_9267,N_36,N_1069);
and U9268 (N_9268,N_4686,N_457);
nor U9269 (N_9269,N_2577,N_1406);
and U9270 (N_9270,N_4877,N_363);
and U9271 (N_9271,N_4071,N_1825);
and U9272 (N_9272,N_495,N_3656);
nand U9273 (N_9273,N_3930,N_3433);
or U9274 (N_9274,N_3477,N_2129);
xor U9275 (N_9275,N_2065,N_923);
nor U9276 (N_9276,N_243,N_4312);
nor U9277 (N_9277,N_851,N_122);
nand U9278 (N_9278,N_3594,N_4128);
xnor U9279 (N_9279,N_3202,N_600);
and U9280 (N_9280,N_2215,N_539);
and U9281 (N_9281,N_188,N_4416);
nand U9282 (N_9282,N_1465,N_2449);
xor U9283 (N_9283,N_1549,N_3577);
or U9284 (N_9284,N_851,N_3638);
nor U9285 (N_9285,N_4164,N_2584);
and U9286 (N_9286,N_1392,N_1318);
nor U9287 (N_9287,N_2455,N_4962);
and U9288 (N_9288,N_4160,N_1650);
nand U9289 (N_9289,N_673,N_3504);
or U9290 (N_9290,N_1232,N_1844);
or U9291 (N_9291,N_3771,N_4921);
or U9292 (N_9292,N_4310,N_281);
and U9293 (N_9293,N_4893,N_1447);
xor U9294 (N_9294,N_3019,N_4117);
nor U9295 (N_9295,N_4820,N_3785);
xor U9296 (N_9296,N_3534,N_4267);
nand U9297 (N_9297,N_1214,N_3519);
or U9298 (N_9298,N_598,N_4600);
nor U9299 (N_9299,N_4981,N_4843);
and U9300 (N_9300,N_2575,N_802);
or U9301 (N_9301,N_1077,N_1884);
xor U9302 (N_9302,N_3833,N_1409);
or U9303 (N_9303,N_4370,N_2263);
nor U9304 (N_9304,N_729,N_2734);
nand U9305 (N_9305,N_1694,N_4580);
or U9306 (N_9306,N_2466,N_1562);
or U9307 (N_9307,N_780,N_934);
xnor U9308 (N_9308,N_4870,N_1570);
nand U9309 (N_9309,N_4372,N_3441);
or U9310 (N_9310,N_1527,N_482);
xnor U9311 (N_9311,N_1771,N_4784);
nand U9312 (N_9312,N_4304,N_9);
nor U9313 (N_9313,N_754,N_1091);
nor U9314 (N_9314,N_1039,N_2939);
nor U9315 (N_9315,N_584,N_2881);
or U9316 (N_9316,N_1578,N_4795);
or U9317 (N_9317,N_1504,N_2784);
and U9318 (N_9318,N_3237,N_2283);
nor U9319 (N_9319,N_521,N_2238);
nand U9320 (N_9320,N_1317,N_4423);
nor U9321 (N_9321,N_4824,N_3431);
nor U9322 (N_9322,N_1514,N_3467);
or U9323 (N_9323,N_3420,N_1208);
nor U9324 (N_9324,N_3469,N_4085);
and U9325 (N_9325,N_1517,N_693);
nor U9326 (N_9326,N_1505,N_657);
and U9327 (N_9327,N_3816,N_1993);
or U9328 (N_9328,N_1809,N_836);
xor U9329 (N_9329,N_967,N_1783);
nand U9330 (N_9330,N_224,N_380);
xor U9331 (N_9331,N_455,N_4248);
and U9332 (N_9332,N_4145,N_1602);
nand U9333 (N_9333,N_3724,N_1489);
nor U9334 (N_9334,N_2984,N_596);
xor U9335 (N_9335,N_664,N_3830);
nand U9336 (N_9336,N_1689,N_1494);
and U9337 (N_9337,N_1232,N_3338);
or U9338 (N_9338,N_2288,N_2111);
nand U9339 (N_9339,N_537,N_1858);
nand U9340 (N_9340,N_977,N_1455);
or U9341 (N_9341,N_99,N_3013);
or U9342 (N_9342,N_4686,N_30);
nand U9343 (N_9343,N_2943,N_1311);
nand U9344 (N_9344,N_1019,N_2003);
and U9345 (N_9345,N_2700,N_4177);
or U9346 (N_9346,N_3940,N_3314);
or U9347 (N_9347,N_4888,N_2506);
xnor U9348 (N_9348,N_1597,N_1796);
nand U9349 (N_9349,N_505,N_4601);
and U9350 (N_9350,N_2252,N_4162);
nor U9351 (N_9351,N_609,N_3447);
nand U9352 (N_9352,N_3081,N_795);
nand U9353 (N_9353,N_4613,N_2975);
and U9354 (N_9354,N_1838,N_737);
xor U9355 (N_9355,N_2492,N_2477);
nor U9356 (N_9356,N_3265,N_915);
and U9357 (N_9357,N_500,N_2299);
and U9358 (N_9358,N_455,N_4328);
or U9359 (N_9359,N_2236,N_4582);
and U9360 (N_9360,N_1666,N_3051);
or U9361 (N_9361,N_1083,N_4042);
xor U9362 (N_9362,N_3478,N_2021);
nor U9363 (N_9363,N_1909,N_998);
and U9364 (N_9364,N_4002,N_2065);
nand U9365 (N_9365,N_2463,N_1608);
xor U9366 (N_9366,N_1999,N_1264);
xnor U9367 (N_9367,N_1260,N_1248);
or U9368 (N_9368,N_2224,N_87);
xnor U9369 (N_9369,N_2818,N_3266);
and U9370 (N_9370,N_598,N_2204);
nand U9371 (N_9371,N_215,N_3210);
nand U9372 (N_9372,N_2969,N_1204);
nor U9373 (N_9373,N_1016,N_1067);
nor U9374 (N_9374,N_890,N_174);
or U9375 (N_9375,N_3508,N_4699);
or U9376 (N_9376,N_1596,N_2612);
xnor U9377 (N_9377,N_4068,N_3704);
and U9378 (N_9378,N_897,N_336);
or U9379 (N_9379,N_2303,N_1170);
nor U9380 (N_9380,N_3983,N_2748);
nand U9381 (N_9381,N_1621,N_2677);
and U9382 (N_9382,N_2820,N_4955);
and U9383 (N_9383,N_70,N_3274);
and U9384 (N_9384,N_4398,N_4842);
or U9385 (N_9385,N_4951,N_2854);
or U9386 (N_9386,N_2727,N_1294);
nand U9387 (N_9387,N_1413,N_1234);
or U9388 (N_9388,N_4728,N_1086);
or U9389 (N_9389,N_895,N_2494);
and U9390 (N_9390,N_4160,N_3355);
xnor U9391 (N_9391,N_4494,N_3579);
xnor U9392 (N_9392,N_3872,N_2744);
nor U9393 (N_9393,N_1587,N_2202);
nand U9394 (N_9394,N_2588,N_296);
and U9395 (N_9395,N_4502,N_1904);
xnor U9396 (N_9396,N_4445,N_4171);
or U9397 (N_9397,N_3890,N_1073);
or U9398 (N_9398,N_3517,N_3900);
nor U9399 (N_9399,N_1822,N_290);
and U9400 (N_9400,N_2679,N_933);
and U9401 (N_9401,N_1774,N_3540);
nor U9402 (N_9402,N_681,N_2225);
xnor U9403 (N_9403,N_4649,N_2293);
and U9404 (N_9404,N_4687,N_971);
xor U9405 (N_9405,N_3784,N_4934);
nand U9406 (N_9406,N_2246,N_4260);
nand U9407 (N_9407,N_4763,N_644);
nor U9408 (N_9408,N_1215,N_2297);
and U9409 (N_9409,N_4273,N_1004);
nand U9410 (N_9410,N_3462,N_2478);
nand U9411 (N_9411,N_517,N_95);
or U9412 (N_9412,N_2127,N_4203);
nor U9413 (N_9413,N_1083,N_2356);
nor U9414 (N_9414,N_2592,N_3523);
or U9415 (N_9415,N_1459,N_4697);
or U9416 (N_9416,N_2450,N_1717);
xor U9417 (N_9417,N_4625,N_1315);
or U9418 (N_9418,N_3959,N_3208);
and U9419 (N_9419,N_3105,N_4949);
or U9420 (N_9420,N_2240,N_2818);
and U9421 (N_9421,N_990,N_2639);
xnor U9422 (N_9422,N_2804,N_1659);
nor U9423 (N_9423,N_4243,N_2482);
and U9424 (N_9424,N_2025,N_403);
or U9425 (N_9425,N_4702,N_417);
and U9426 (N_9426,N_1028,N_2893);
nor U9427 (N_9427,N_1366,N_3333);
or U9428 (N_9428,N_4767,N_3564);
and U9429 (N_9429,N_4873,N_322);
nor U9430 (N_9430,N_582,N_198);
nor U9431 (N_9431,N_444,N_415);
and U9432 (N_9432,N_1022,N_4390);
xor U9433 (N_9433,N_4092,N_4493);
and U9434 (N_9434,N_2366,N_3310);
xnor U9435 (N_9435,N_4594,N_1092);
or U9436 (N_9436,N_2318,N_4305);
nor U9437 (N_9437,N_536,N_4764);
and U9438 (N_9438,N_4210,N_1209);
and U9439 (N_9439,N_4261,N_581);
nor U9440 (N_9440,N_4504,N_2623);
or U9441 (N_9441,N_4263,N_3015);
and U9442 (N_9442,N_1211,N_2640);
and U9443 (N_9443,N_1121,N_494);
xnor U9444 (N_9444,N_1613,N_2471);
nand U9445 (N_9445,N_4238,N_2079);
and U9446 (N_9446,N_523,N_4217);
or U9447 (N_9447,N_4459,N_4371);
xnor U9448 (N_9448,N_1396,N_1646);
or U9449 (N_9449,N_1752,N_684);
nor U9450 (N_9450,N_3704,N_1355);
nor U9451 (N_9451,N_1603,N_3779);
nand U9452 (N_9452,N_186,N_994);
nand U9453 (N_9453,N_592,N_3542);
xor U9454 (N_9454,N_89,N_2632);
xor U9455 (N_9455,N_4032,N_1350);
or U9456 (N_9456,N_1925,N_3114);
xnor U9457 (N_9457,N_475,N_578);
or U9458 (N_9458,N_3248,N_2426);
nor U9459 (N_9459,N_4627,N_2588);
xor U9460 (N_9460,N_2225,N_1775);
xnor U9461 (N_9461,N_321,N_1567);
nand U9462 (N_9462,N_513,N_1609);
or U9463 (N_9463,N_2449,N_4400);
xor U9464 (N_9464,N_378,N_2468);
xnor U9465 (N_9465,N_3369,N_3024);
or U9466 (N_9466,N_4978,N_3131);
nor U9467 (N_9467,N_1487,N_794);
nand U9468 (N_9468,N_1744,N_1572);
or U9469 (N_9469,N_1195,N_192);
and U9470 (N_9470,N_877,N_3856);
and U9471 (N_9471,N_2883,N_3965);
xor U9472 (N_9472,N_252,N_1681);
or U9473 (N_9473,N_849,N_2268);
and U9474 (N_9474,N_2123,N_2798);
nor U9475 (N_9475,N_3047,N_2176);
or U9476 (N_9476,N_1094,N_4281);
nor U9477 (N_9477,N_3002,N_987);
xnor U9478 (N_9478,N_1874,N_508);
nor U9479 (N_9479,N_4940,N_780);
or U9480 (N_9480,N_1015,N_1950);
and U9481 (N_9481,N_4431,N_4937);
nor U9482 (N_9482,N_3770,N_3997);
nor U9483 (N_9483,N_3257,N_1695);
or U9484 (N_9484,N_1092,N_1589);
nor U9485 (N_9485,N_130,N_4375);
and U9486 (N_9486,N_885,N_2035);
nor U9487 (N_9487,N_1288,N_3348);
or U9488 (N_9488,N_1154,N_4136);
nor U9489 (N_9489,N_3147,N_1463);
and U9490 (N_9490,N_4603,N_3507);
and U9491 (N_9491,N_2757,N_1169);
and U9492 (N_9492,N_3282,N_16);
nand U9493 (N_9493,N_2959,N_4646);
nand U9494 (N_9494,N_3207,N_1933);
nor U9495 (N_9495,N_1996,N_1367);
xnor U9496 (N_9496,N_3964,N_900);
and U9497 (N_9497,N_3282,N_1321);
nor U9498 (N_9498,N_2652,N_1106);
xor U9499 (N_9499,N_2379,N_4893);
xnor U9500 (N_9500,N_4889,N_1748);
nand U9501 (N_9501,N_1115,N_3039);
xnor U9502 (N_9502,N_492,N_4610);
nor U9503 (N_9503,N_1080,N_815);
and U9504 (N_9504,N_4433,N_296);
xnor U9505 (N_9505,N_3364,N_4667);
xnor U9506 (N_9506,N_4659,N_2274);
or U9507 (N_9507,N_3858,N_1515);
xnor U9508 (N_9508,N_941,N_1193);
nor U9509 (N_9509,N_4942,N_4668);
or U9510 (N_9510,N_3454,N_1709);
and U9511 (N_9511,N_3238,N_4499);
nand U9512 (N_9512,N_807,N_4502);
nand U9513 (N_9513,N_3062,N_706);
and U9514 (N_9514,N_894,N_3763);
xor U9515 (N_9515,N_4199,N_394);
or U9516 (N_9516,N_4898,N_1582);
and U9517 (N_9517,N_1202,N_346);
xnor U9518 (N_9518,N_885,N_1465);
and U9519 (N_9519,N_874,N_2011);
xor U9520 (N_9520,N_4008,N_3367);
nand U9521 (N_9521,N_2046,N_610);
nor U9522 (N_9522,N_4177,N_713);
nor U9523 (N_9523,N_3985,N_742);
or U9524 (N_9524,N_685,N_275);
and U9525 (N_9525,N_1152,N_3711);
nor U9526 (N_9526,N_1237,N_4372);
or U9527 (N_9527,N_960,N_2829);
xor U9528 (N_9528,N_2250,N_738);
or U9529 (N_9529,N_799,N_4359);
and U9530 (N_9530,N_1174,N_1924);
nor U9531 (N_9531,N_3965,N_104);
nor U9532 (N_9532,N_3682,N_1506);
xnor U9533 (N_9533,N_2663,N_1544);
or U9534 (N_9534,N_995,N_4287);
and U9535 (N_9535,N_375,N_3902);
nand U9536 (N_9536,N_476,N_3955);
or U9537 (N_9537,N_3133,N_714);
and U9538 (N_9538,N_3362,N_3327);
nor U9539 (N_9539,N_1435,N_4237);
xor U9540 (N_9540,N_4815,N_4295);
nand U9541 (N_9541,N_876,N_4876);
nand U9542 (N_9542,N_2046,N_2000);
nand U9543 (N_9543,N_3132,N_3979);
and U9544 (N_9544,N_679,N_3742);
xor U9545 (N_9545,N_3505,N_3458);
nand U9546 (N_9546,N_3154,N_399);
nand U9547 (N_9547,N_1688,N_2792);
or U9548 (N_9548,N_222,N_2137);
nand U9549 (N_9549,N_2432,N_4229);
xor U9550 (N_9550,N_448,N_480);
nand U9551 (N_9551,N_3439,N_3135);
or U9552 (N_9552,N_2283,N_4650);
or U9553 (N_9553,N_78,N_1685);
and U9554 (N_9554,N_1257,N_4812);
nand U9555 (N_9555,N_2022,N_4881);
or U9556 (N_9556,N_137,N_1654);
nor U9557 (N_9557,N_1139,N_2721);
or U9558 (N_9558,N_473,N_1270);
and U9559 (N_9559,N_3717,N_2330);
and U9560 (N_9560,N_4304,N_460);
and U9561 (N_9561,N_798,N_4709);
and U9562 (N_9562,N_1713,N_1393);
nor U9563 (N_9563,N_4333,N_2734);
and U9564 (N_9564,N_752,N_2896);
nor U9565 (N_9565,N_1569,N_3625);
or U9566 (N_9566,N_1845,N_3348);
nor U9567 (N_9567,N_1234,N_4460);
or U9568 (N_9568,N_1037,N_229);
and U9569 (N_9569,N_91,N_4834);
and U9570 (N_9570,N_44,N_4183);
nand U9571 (N_9571,N_1566,N_1820);
nor U9572 (N_9572,N_3117,N_777);
nand U9573 (N_9573,N_882,N_2927);
nor U9574 (N_9574,N_2710,N_2167);
and U9575 (N_9575,N_1342,N_2191);
nor U9576 (N_9576,N_4558,N_2390);
and U9577 (N_9577,N_861,N_4261);
xnor U9578 (N_9578,N_92,N_1805);
nor U9579 (N_9579,N_3282,N_4754);
xor U9580 (N_9580,N_3415,N_4828);
nand U9581 (N_9581,N_2650,N_2048);
nor U9582 (N_9582,N_452,N_3252);
nand U9583 (N_9583,N_992,N_1942);
or U9584 (N_9584,N_163,N_2395);
nor U9585 (N_9585,N_672,N_1772);
and U9586 (N_9586,N_3959,N_3716);
nor U9587 (N_9587,N_3716,N_4807);
xnor U9588 (N_9588,N_1400,N_187);
and U9589 (N_9589,N_3467,N_3663);
nor U9590 (N_9590,N_2496,N_3658);
or U9591 (N_9591,N_57,N_3505);
nor U9592 (N_9592,N_1350,N_4090);
nand U9593 (N_9593,N_1340,N_1068);
nor U9594 (N_9594,N_4572,N_4287);
nand U9595 (N_9595,N_4123,N_4910);
xnor U9596 (N_9596,N_1183,N_2546);
and U9597 (N_9597,N_4845,N_3581);
nand U9598 (N_9598,N_4923,N_2211);
xor U9599 (N_9599,N_3156,N_3555);
xor U9600 (N_9600,N_4817,N_400);
nor U9601 (N_9601,N_3098,N_4449);
or U9602 (N_9602,N_1544,N_2743);
xnor U9603 (N_9603,N_3284,N_1118);
and U9604 (N_9604,N_709,N_2159);
nor U9605 (N_9605,N_2170,N_3702);
nor U9606 (N_9606,N_4769,N_3928);
nand U9607 (N_9607,N_804,N_3794);
nand U9608 (N_9608,N_3464,N_2322);
xnor U9609 (N_9609,N_3371,N_96);
and U9610 (N_9610,N_2786,N_2365);
xor U9611 (N_9611,N_2034,N_1237);
nor U9612 (N_9612,N_1427,N_2267);
nand U9613 (N_9613,N_366,N_506);
nand U9614 (N_9614,N_55,N_319);
nor U9615 (N_9615,N_134,N_2948);
and U9616 (N_9616,N_4851,N_4495);
nor U9617 (N_9617,N_868,N_2954);
nand U9618 (N_9618,N_1768,N_4971);
nor U9619 (N_9619,N_2710,N_2197);
nor U9620 (N_9620,N_4693,N_2759);
nor U9621 (N_9621,N_2484,N_1595);
nand U9622 (N_9622,N_2334,N_3191);
nand U9623 (N_9623,N_2064,N_4941);
nor U9624 (N_9624,N_2401,N_3596);
or U9625 (N_9625,N_4254,N_4804);
nand U9626 (N_9626,N_1734,N_4226);
and U9627 (N_9627,N_1182,N_4104);
or U9628 (N_9628,N_4873,N_1002);
nand U9629 (N_9629,N_1312,N_895);
and U9630 (N_9630,N_790,N_4136);
nor U9631 (N_9631,N_4473,N_4666);
or U9632 (N_9632,N_1905,N_1934);
xor U9633 (N_9633,N_3102,N_4763);
nor U9634 (N_9634,N_3024,N_1603);
nor U9635 (N_9635,N_2362,N_3175);
and U9636 (N_9636,N_1308,N_3190);
nand U9637 (N_9637,N_1082,N_3642);
nor U9638 (N_9638,N_996,N_3366);
nor U9639 (N_9639,N_4507,N_1541);
xor U9640 (N_9640,N_2188,N_2444);
and U9641 (N_9641,N_3886,N_2585);
nand U9642 (N_9642,N_4013,N_2023);
xor U9643 (N_9643,N_3696,N_2877);
nor U9644 (N_9644,N_4002,N_2142);
xor U9645 (N_9645,N_2414,N_4061);
nand U9646 (N_9646,N_4574,N_4840);
nand U9647 (N_9647,N_1721,N_3663);
xor U9648 (N_9648,N_503,N_3942);
and U9649 (N_9649,N_790,N_3015);
or U9650 (N_9650,N_756,N_103);
nand U9651 (N_9651,N_2694,N_126);
and U9652 (N_9652,N_4274,N_4054);
or U9653 (N_9653,N_1778,N_4210);
and U9654 (N_9654,N_3672,N_2287);
or U9655 (N_9655,N_2906,N_3087);
nand U9656 (N_9656,N_1833,N_4338);
or U9657 (N_9657,N_1674,N_147);
and U9658 (N_9658,N_433,N_2058);
or U9659 (N_9659,N_28,N_1429);
and U9660 (N_9660,N_2636,N_3863);
nor U9661 (N_9661,N_1118,N_1516);
nor U9662 (N_9662,N_2310,N_722);
and U9663 (N_9663,N_481,N_4092);
or U9664 (N_9664,N_3831,N_4640);
or U9665 (N_9665,N_1553,N_704);
xnor U9666 (N_9666,N_2498,N_564);
and U9667 (N_9667,N_360,N_453);
and U9668 (N_9668,N_4439,N_965);
nor U9669 (N_9669,N_2506,N_1241);
nor U9670 (N_9670,N_559,N_3166);
or U9671 (N_9671,N_1568,N_612);
nand U9672 (N_9672,N_1838,N_628);
nand U9673 (N_9673,N_4037,N_370);
or U9674 (N_9674,N_2956,N_4181);
xor U9675 (N_9675,N_2721,N_3071);
nand U9676 (N_9676,N_245,N_697);
or U9677 (N_9677,N_4677,N_974);
or U9678 (N_9678,N_3427,N_947);
nand U9679 (N_9679,N_983,N_300);
nor U9680 (N_9680,N_3886,N_2695);
or U9681 (N_9681,N_4881,N_247);
and U9682 (N_9682,N_1856,N_2385);
and U9683 (N_9683,N_2034,N_1892);
nor U9684 (N_9684,N_2744,N_684);
nor U9685 (N_9685,N_177,N_1254);
xnor U9686 (N_9686,N_3839,N_2384);
and U9687 (N_9687,N_4783,N_1542);
nor U9688 (N_9688,N_550,N_4296);
nand U9689 (N_9689,N_1817,N_48);
xor U9690 (N_9690,N_382,N_4587);
or U9691 (N_9691,N_65,N_2548);
nor U9692 (N_9692,N_2062,N_4653);
and U9693 (N_9693,N_1951,N_128);
and U9694 (N_9694,N_2103,N_4026);
xnor U9695 (N_9695,N_4944,N_1870);
nand U9696 (N_9696,N_441,N_1237);
or U9697 (N_9697,N_1155,N_1032);
and U9698 (N_9698,N_304,N_4123);
or U9699 (N_9699,N_683,N_987);
or U9700 (N_9700,N_998,N_2025);
or U9701 (N_9701,N_3071,N_4505);
nand U9702 (N_9702,N_3224,N_1941);
or U9703 (N_9703,N_977,N_1574);
and U9704 (N_9704,N_4655,N_2483);
and U9705 (N_9705,N_4877,N_3867);
nor U9706 (N_9706,N_4085,N_1373);
or U9707 (N_9707,N_4975,N_2837);
or U9708 (N_9708,N_1629,N_350);
and U9709 (N_9709,N_1176,N_4075);
nand U9710 (N_9710,N_4459,N_2777);
xor U9711 (N_9711,N_3757,N_2328);
nor U9712 (N_9712,N_4486,N_4633);
xor U9713 (N_9713,N_3026,N_4449);
or U9714 (N_9714,N_3284,N_3612);
nand U9715 (N_9715,N_467,N_694);
or U9716 (N_9716,N_1655,N_2759);
or U9717 (N_9717,N_71,N_1688);
or U9718 (N_9718,N_2917,N_3793);
nand U9719 (N_9719,N_1974,N_2986);
or U9720 (N_9720,N_1393,N_999);
or U9721 (N_9721,N_112,N_565);
nand U9722 (N_9722,N_314,N_3696);
nor U9723 (N_9723,N_3159,N_3915);
xor U9724 (N_9724,N_2429,N_4928);
or U9725 (N_9725,N_2182,N_187);
nand U9726 (N_9726,N_4092,N_1389);
or U9727 (N_9727,N_1054,N_4237);
and U9728 (N_9728,N_2713,N_4964);
and U9729 (N_9729,N_781,N_3686);
xnor U9730 (N_9730,N_1239,N_3501);
nand U9731 (N_9731,N_3268,N_1068);
xor U9732 (N_9732,N_423,N_2951);
and U9733 (N_9733,N_4247,N_3869);
nor U9734 (N_9734,N_2090,N_2248);
nor U9735 (N_9735,N_546,N_3738);
xnor U9736 (N_9736,N_2754,N_3659);
xor U9737 (N_9737,N_3727,N_1976);
and U9738 (N_9738,N_3347,N_877);
xnor U9739 (N_9739,N_3793,N_4724);
and U9740 (N_9740,N_2227,N_2058);
nor U9741 (N_9741,N_369,N_4210);
nor U9742 (N_9742,N_50,N_4225);
and U9743 (N_9743,N_843,N_3416);
and U9744 (N_9744,N_808,N_1073);
nor U9745 (N_9745,N_1905,N_3645);
or U9746 (N_9746,N_1875,N_4857);
nand U9747 (N_9747,N_4398,N_2149);
xnor U9748 (N_9748,N_1575,N_2836);
nor U9749 (N_9749,N_1731,N_1127);
or U9750 (N_9750,N_1392,N_790);
nor U9751 (N_9751,N_4865,N_2883);
nor U9752 (N_9752,N_343,N_2983);
and U9753 (N_9753,N_1770,N_561);
and U9754 (N_9754,N_193,N_280);
or U9755 (N_9755,N_647,N_3058);
or U9756 (N_9756,N_657,N_3153);
xnor U9757 (N_9757,N_4161,N_169);
and U9758 (N_9758,N_2621,N_4101);
nor U9759 (N_9759,N_1156,N_876);
xor U9760 (N_9760,N_3049,N_2344);
and U9761 (N_9761,N_585,N_728);
nand U9762 (N_9762,N_433,N_2955);
nor U9763 (N_9763,N_416,N_2889);
nor U9764 (N_9764,N_4250,N_595);
or U9765 (N_9765,N_3392,N_1647);
xor U9766 (N_9766,N_1649,N_4314);
or U9767 (N_9767,N_3437,N_4461);
xor U9768 (N_9768,N_1967,N_4923);
and U9769 (N_9769,N_1760,N_2859);
and U9770 (N_9770,N_3855,N_2393);
and U9771 (N_9771,N_4070,N_3478);
xnor U9772 (N_9772,N_4536,N_2844);
or U9773 (N_9773,N_3921,N_476);
xnor U9774 (N_9774,N_4114,N_153);
or U9775 (N_9775,N_4423,N_7);
and U9776 (N_9776,N_2533,N_4177);
and U9777 (N_9777,N_1836,N_753);
nor U9778 (N_9778,N_1492,N_1215);
xnor U9779 (N_9779,N_2967,N_1205);
nor U9780 (N_9780,N_768,N_245);
or U9781 (N_9781,N_2532,N_1315);
nand U9782 (N_9782,N_1313,N_1430);
or U9783 (N_9783,N_2722,N_4149);
xor U9784 (N_9784,N_158,N_2410);
and U9785 (N_9785,N_439,N_3309);
xor U9786 (N_9786,N_443,N_543);
xnor U9787 (N_9787,N_948,N_2096);
and U9788 (N_9788,N_758,N_1061);
and U9789 (N_9789,N_4089,N_1508);
nor U9790 (N_9790,N_3559,N_234);
or U9791 (N_9791,N_1728,N_116);
or U9792 (N_9792,N_4656,N_874);
nor U9793 (N_9793,N_119,N_4087);
nor U9794 (N_9794,N_3020,N_1216);
nand U9795 (N_9795,N_4518,N_335);
xnor U9796 (N_9796,N_3121,N_3360);
or U9797 (N_9797,N_2015,N_1053);
xor U9798 (N_9798,N_3675,N_2717);
and U9799 (N_9799,N_3829,N_2935);
xnor U9800 (N_9800,N_1155,N_4839);
xnor U9801 (N_9801,N_1189,N_4528);
and U9802 (N_9802,N_850,N_4341);
nor U9803 (N_9803,N_4782,N_3911);
nor U9804 (N_9804,N_2867,N_3793);
nor U9805 (N_9805,N_4895,N_3417);
or U9806 (N_9806,N_1612,N_4806);
nand U9807 (N_9807,N_3740,N_4275);
nor U9808 (N_9808,N_2139,N_32);
or U9809 (N_9809,N_1608,N_107);
and U9810 (N_9810,N_559,N_4632);
nor U9811 (N_9811,N_2211,N_332);
or U9812 (N_9812,N_252,N_410);
and U9813 (N_9813,N_621,N_1948);
nor U9814 (N_9814,N_77,N_2980);
nor U9815 (N_9815,N_4770,N_2307);
xor U9816 (N_9816,N_2105,N_698);
or U9817 (N_9817,N_1279,N_581);
or U9818 (N_9818,N_4167,N_1674);
nand U9819 (N_9819,N_367,N_4255);
nor U9820 (N_9820,N_64,N_623);
nand U9821 (N_9821,N_3792,N_4713);
xor U9822 (N_9822,N_4386,N_2296);
or U9823 (N_9823,N_4331,N_695);
or U9824 (N_9824,N_2488,N_813);
and U9825 (N_9825,N_90,N_1842);
nand U9826 (N_9826,N_3321,N_1168);
nand U9827 (N_9827,N_4440,N_2335);
and U9828 (N_9828,N_2725,N_2728);
nand U9829 (N_9829,N_3864,N_1761);
or U9830 (N_9830,N_2554,N_2781);
xor U9831 (N_9831,N_723,N_2199);
or U9832 (N_9832,N_2329,N_3694);
nor U9833 (N_9833,N_652,N_2510);
and U9834 (N_9834,N_1043,N_690);
or U9835 (N_9835,N_694,N_1212);
nand U9836 (N_9836,N_2249,N_1082);
xor U9837 (N_9837,N_4034,N_4043);
nor U9838 (N_9838,N_2204,N_3317);
nand U9839 (N_9839,N_2689,N_808);
nand U9840 (N_9840,N_4078,N_48);
or U9841 (N_9841,N_4847,N_4084);
and U9842 (N_9842,N_4243,N_4162);
nor U9843 (N_9843,N_1201,N_3529);
nor U9844 (N_9844,N_3750,N_4103);
and U9845 (N_9845,N_4450,N_4979);
nor U9846 (N_9846,N_973,N_4745);
or U9847 (N_9847,N_2954,N_2264);
nor U9848 (N_9848,N_168,N_2558);
and U9849 (N_9849,N_4410,N_3457);
xnor U9850 (N_9850,N_105,N_4496);
and U9851 (N_9851,N_1730,N_584);
or U9852 (N_9852,N_2470,N_4700);
nand U9853 (N_9853,N_2999,N_2887);
nand U9854 (N_9854,N_335,N_4696);
nand U9855 (N_9855,N_3207,N_1225);
nor U9856 (N_9856,N_4480,N_151);
nor U9857 (N_9857,N_1820,N_6);
xnor U9858 (N_9858,N_1904,N_3022);
and U9859 (N_9859,N_1051,N_2949);
nand U9860 (N_9860,N_606,N_317);
and U9861 (N_9861,N_4208,N_4314);
xnor U9862 (N_9862,N_4761,N_866);
and U9863 (N_9863,N_4395,N_1184);
xor U9864 (N_9864,N_1596,N_998);
nor U9865 (N_9865,N_2660,N_1254);
or U9866 (N_9866,N_2150,N_1692);
nand U9867 (N_9867,N_2429,N_2742);
or U9868 (N_9868,N_4502,N_2631);
or U9869 (N_9869,N_4890,N_3545);
nor U9870 (N_9870,N_1164,N_310);
xor U9871 (N_9871,N_3162,N_3384);
nand U9872 (N_9872,N_3964,N_567);
xor U9873 (N_9873,N_4874,N_2679);
or U9874 (N_9874,N_3689,N_2898);
nor U9875 (N_9875,N_4072,N_2787);
xor U9876 (N_9876,N_4344,N_2430);
and U9877 (N_9877,N_2219,N_1953);
nor U9878 (N_9878,N_4327,N_3355);
xor U9879 (N_9879,N_4916,N_3578);
and U9880 (N_9880,N_3020,N_1308);
or U9881 (N_9881,N_2223,N_1046);
or U9882 (N_9882,N_2079,N_3817);
nor U9883 (N_9883,N_10,N_4296);
nand U9884 (N_9884,N_1639,N_1449);
and U9885 (N_9885,N_366,N_49);
and U9886 (N_9886,N_3853,N_4756);
nand U9887 (N_9887,N_1318,N_666);
or U9888 (N_9888,N_2948,N_95);
xnor U9889 (N_9889,N_3313,N_4891);
and U9890 (N_9890,N_4112,N_3724);
or U9891 (N_9891,N_3359,N_3569);
or U9892 (N_9892,N_3038,N_4955);
nor U9893 (N_9893,N_2041,N_3463);
or U9894 (N_9894,N_4572,N_4376);
and U9895 (N_9895,N_4840,N_3232);
and U9896 (N_9896,N_2628,N_4251);
nor U9897 (N_9897,N_4666,N_1017);
or U9898 (N_9898,N_773,N_1265);
nand U9899 (N_9899,N_4973,N_997);
nor U9900 (N_9900,N_3950,N_4308);
nand U9901 (N_9901,N_2624,N_2870);
and U9902 (N_9902,N_2836,N_3703);
nor U9903 (N_9903,N_3930,N_141);
or U9904 (N_9904,N_3704,N_962);
or U9905 (N_9905,N_3004,N_2854);
nand U9906 (N_9906,N_4993,N_3983);
and U9907 (N_9907,N_2306,N_3543);
and U9908 (N_9908,N_3289,N_268);
or U9909 (N_9909,N_1784,N_1941);
and U9910 (N_9910,N_1750,N_2494);
xor U9911 (N_9911,N_2219,N_1937);
or U9912 (N_9912,N_2448,N_1660);
xnor U9913 (N_9913,N_1069,N_831);
xnor U9914 (N_9914,N_3207,N_2362);
and U9915 (N_9915,N_3175,N_1761);
nand U9916 (N_9916,N_1145,N_2457);
nand U9917 (N_9917,N_4826,N_84);
and U9918 (N_9918,N_671,N_1454);
nand U9919 (N_9919,N_4489,N_2187);
or U9920 (N_9920,N_2231,N_117);
and U9921 (N_9921,N_757,N_3751);
nand U9922 (N_9922,N_3419,N_2249);
or U9923 (N_9923,N_4445,N_2811);
xor U9924 (N_9924,N_292,N_2073);
xor U9925 (N_9925,N_1392,N_987);
and U9926 (N_9926,N_4507,N_3718);
or U9927 (N_9927,N_4988,N_3336);
nor U9928 (N_9928,N_2321,N_2816);
nand U9929 (N_9929,N_2029,N_2893);
xnor U9930 (N_9930,N_4668,N_1089);
xor U9931 (N_9931,N_3517,N_631);
nand U9932 (N_9932,N_3126,N_3969);
nor U9933 (N_9933,N_3474,N_2640);
nor U9934 (N_9934,N_657,N_562);
nor U9935 (N_9935,N_2881,N_1827);
and U9936 (N_9936,N_1829,N_2788);
or U9937 (N_9937,N_3596,N_2308);
and U9938 (N_9938,N_4403,N_3917);
nand U9939 (N_9939,N_983,N_1459);
nor U9940 (N_9940,N_1943,N_401);
nor U9941 (N_9941,N_4502,N_3933);
nor U9942 (N_9942,N_1762,N_3639);
nor U9943 (N_9943,N_3886,N_2231);
xor U9944 (N_9944,N_3419,N_749);
xor U9945 (N_9945,N_1939,N_1036);
and U9946 (N_9946,N_2701,N_1242);
and U9947 (N_9947,N_586,N_1260);
and U9948 (N_9948,N_422,N_410);
and U9949 (N_9949,N_1111,N_4740);
nand U9950 (N_9950,N_4785,N_2138);
nand U9951 (N_9951,N_487,N_3694);
and U9952 (N_9952,N_1820,N_3264);
and U9953 (N_9953,N_1281,N_2177);
and U9954 (N_9954,N_4115,N_211);
nor U9955 (N_9955,N_625,N_3365);
nand U9956 (N_9956,N_3177,N_1946);
nor U9957 (N_9957,N_3191,N_3873);
and U9958 (N_9958,N_4941,N_623);
xor U9959 (N_9959,N_1141,N_1725);
nor U9960 (N_9960,N_1187,N_4811);
or U9961 (N_9961,N_3945,N_2544);
nand U9962 (N_9962,N_2604,N_672);
and U9963 (N_9963,N_1506,N_90);
nor U9964 (N_9964,N_4019,N_399);
xor U9965 (N_9965,N_2112,N_35);
or U9966 (N_9966,N_832,N_72);
or U9967 (N_9967,N_3791,N_3487);
xnor U9968 (N_9968,N_552,N_4993);
nand U9969 (N_9969,N_798,N_539);
nand U9970 (N_9970,N_2400,N_2199);
or U9971 (N_9971,N_3979,N_1548);
nand U9972 (N_9972,N_1361,N_3855);
nand U9973 (N_9973,N_2929,N_4673);
nand U9974 (N_9974,N_1260,N_3341);
xor U9975 (N_9975,N_2542,N_2781);
nand U9976 (N_9976,N_2747,N_3062);
and U9977 (N_9977,N_2628,N_547);
and U9978 (N_9978,N_2954,N_597);
xnor U9979 (N_9979,N_1363,N_4319);
nor U9980 (N_9980,N_4121,N_2157);
nor U9981 (N_9981,N_4028,N_161);
xnor U9982 (N_9982,N_3441,N_1941);
nand U9983 (N_9983,N_850,N_299);
and U9984 (N_9984,N_53,N_4674);
or U9985 (N_9985,N_4259,N_3862);
nand U9986 (N_9986,N_2779,N_2961);
xor U9987 (N_9987,N_908,N_2263);
nand U9988 (N_9988,N_3453,N_4794);
and U9989 (N_9989,N_3031,N_86);
nand U9990 (N_9990,N_2412,N_3714);
xnor U9991 (N_9991,N_1144,N_2103);
nor U9992 (N_9992,N_4827,N_2005);
nand U9993 (N_9993,N_796,N_2447);
and U9994 (N_9994,N_4269,N_1227);
and U9995 (N_9995,N_3813,N_706);
xor U9996 (N_9996,N_2432,N_3315);
or U9997 (N_9997,N_3469,N_2207);
xor U9998 (N_9998,N_2232,N_370);
nand U9999 (N_9999,N_2959,N_1497);
xor UO_0 (O_0,N_8872,N_9041);
xnor UO_1 (O_1,N_5332,N_7981);
or UO_2 (O_2,N_5493,N_5051);
and UO_3 (O_3,N_8741,N_7141);
and UO_4 (O_4,N_5845,N_7505);
nand UO_5 (O_5,N_6953,N_7062);
nor UO_6 (O_6,N_8284,N_9870);
and UO_7 (O_7,N_8300,N_9840);
or UO_8 (O_8,N_7352,N_7559);
xor UO_9 (O_9,N_6430,N_7449);
or UO_10 (O_10,N_9705,N_8243);
nor UO_11 (O_11,N_7703,N_9101);
nor UO_12 (O_12,N_9559,N_7870);
and UO_13 (O_13,N_8818,N_8645);
xor UO_14 (O_14,N_6353,N_9118);
and UO_15 (O_15,N_8537,N_6591);
or UO_16 (O_16,N_6960,N_8718);
xnor UO_17 (O_17,N_8516,N_8364);
and UO_18 (O_18,N_8654,N_9716);
and UO_19 (O_19,N_6753,N_8274);
nor UO_20 (O_20,N_5000,N_7450);
or UO_21 (O_21,N_6051,N_6338);
nor UO_22 (O_22,N_8360,N_8174);
nand UO_23 (O_23,N_5892,N_6948);
xor UO_24 (O_24,N_7109,N_8673);
nor UO_25 (O_25,N_9941,N_8351);
xnor UO_26 (O_26,N_7691,N_5895);
nand UO_27 (O_27,N_5141,N_6598);
xor UO_28 (O_28,N_5581,N_7902);
nand UO_29 (O_29,N_9526,N_7958);
nor UO_30 (O_30,N_6909,N_5157);
or UO_31 (O_31,N_8948,N_9042);
nand UO_32 (O_32,N_5774,N_5398);
and UO_33 (O_33,N_6366,N_6167);
nor UO_34 (O_34,N_8512,N_7353);
xor UO_35 (O_35,N_5223,N_9321);
nand UO_36 (O_36,N_9318,N_8368);
or UO_37 (O_37,N_8681,N_8834);
xor UO_38 (O_38,N_7735,N_5971);
nor UO_39 (O_39,N_6821,N_6696);
and UO_40 (O_40,N_6826,N_8011);
nand UO_41 (O_41,N_5497,N_8137);
nand UO_42 (O_42,N_6933,N_9914);
xor UO_43 (O_43,N_6265,N_9725);
nor UO_44 (O_44,N_5804,N_6813);
or UO_45 (O_45,N_9287,N_9558);
nand UO_46 (O_46,N_6585,N_9432);
or UO_47 (O_47,N_7162,N_6394);
nor UO_48 (O_48,N_5919,N_7395);
nor UO_49 (O_49,N_9803,N_7009);
and UO_50 (O_50,N_8877,N_8520);
and UO_51 (O_51,N_7834,N_5382);
or UO_52 (O_52,N_7388,N_9012);
or UO_53 (O_53,N_6466,N_7836);
and UO_54 (O_54,N_5828,N_6640);
and UO_55 (O_55,N_7265,N_6929);
nand UO_56 (O_56,N_6409,N_6856);
nand UO_57 (O_57,N_8194,N_6657);
nor UO_58 (O_58,N_9336,N_5612);
nand UO_59 (O_59,N_5353,N_6679);
nor UO_60 (O_60,N_7294,N_7864);
and UO_61 (O_61,N_9907,N_7187);
or UO_62 (O_62,N_9173,N_7452);
nor UO_63 (O_63,N_5268,N_6385);
or UO_64 (O_64,N_9875,N_5504);
nor UO_65 (O_65,N_5379,N_8016);
nor UO_66 (O_66,N_5717,N_7862);
and UO_67 (O_67,N_8968,N_9530);
nor UO_68 (O_68,N_8752,N_9873);
or UO_69 (O_69,N_7926,N_5756);
xor UO_70 (O_70,N_5621,N_7618);
nand UO_71 (O_71,N_7175,N_7485);
xor UO_72 (O_72,N_9839,N_7055);
and UO_73 (O_73,N_8603,N_9663);
or UO_74 (O_74,N_6281,N_5301);
or UO_75 (O_75,N_6305,N_6279);
and UO_76 (O_76,N_8433,N_6002);
nor UO_77 (O_77,N_5300,N_5743);
and UO_78 (O_78,N_9834,N_6882);
and UO_79 (O_79,N_5189,N_7940);
nand UO_80 (O_80,N_9029,N_5754);
xor UO_81 (O_81,N_6481,N_8847);
nor UO_82 (O_82,N_8611,N_6898);
nand UO_83 (O_83,N_8070,N_7603);
and UO_84 (O_84,N_5435,N_6984);
or UO_85 (O_85,N_8777,N_8348);
nor UO_86 (O_86,N_9373,N_6631);
and UO_87 (O_87,N_8568,N_9621);
or UO_88 (O_88,N_9847,N_5968);
or UO_89 (O_89,N_7122,N_9735);
and UO_90 (O_90,N_7668,N_6516);
xnor UO_91 (O_91,N_8189,N_8019);
nor UO_92 (O_92,N_8305,N_8538);
xor UO_93 (O_93,N_8134,N_5984);
or UO_94 (O_94,N_9521,N_5833);
xor UO_95 (O_95,N_6534,N_8669);
nor UO_96 (O_96,N_8811,N_7146);
nand UO_97 (O_97,N_8098,N_6901);
and UO_98 (O_98,N_9825,N_5762);
and UO_99 (O_99,N_8254,N_7558);
and UO_100 (O_100,N_9689,N_7569);
nor UO_101 (O_101,N_5168,N_7847);
or UO_102 (O_102,N_6612,N_6857);
xnor UO_103 (O_103,N_6088,N_7761);
nand UO_104 (O_104,N_9229,N_8375);
nand UO_105 (O_105,N_5933,N_9929);
nand UO_106 (O_106,N_5288,N_5535);
or UO_107 (O_107,N_8276,N_7276);
and UO_108 (O_108,N_6511,N_6920);
or UO_109 (O_109,N_5371,N_9676);
nor UO_110 (O_110,N_9113,N_6698);
xor UO_111 (O_111,N_9255,N_6442);
nand UO_112 (O_112,N_9257,N_6503);
nand UO_113 (O_113,N_8269,N_7978);
xnor UO_114 (O_114,N_6810,N_6398);
and UO_115 (O_115,N_9322,N_7059);
and UO_116 (O_116,N_5196,N_5935);
xor UO_117 (O_117,N_8108,N_6151);
xnor UO_118 (O_118,N_5983,N_5097);
xor UO_119 (O_119,N_5145,N_8094);
nand UO_120 (O_120,N_6614,N_5564);
nand UO_121 (O_121,N_9482,N_7104);
xor UO_122 (O_122,N_9271,N_8451);
or UO_123 (O_123,N_5394,N_7514);
nand UO_124 (O_124,N_8885,N_9655);
nand UO_125 (O_125,N_9926,N_8292);
and UO_126 (O_126,N_7218,N_5069);
nor UO_127 (O_127,N_8020,N_5486);
or UO_128 (O_128,N_8365,N_9078);
or UO_129 (O_129,N_8936,N_9228);
nand UO_130 (O_130,N_7822,N_7046);
nand UO_131 (O_131,N_5405,N_7616);
nor UO_132 (O_132,N_6333,N_7742);
or UO_133 (O_133,N_5973,N_9999);
or UO_134 (O_134,N_8805,N_7628);
and UO_135 (O_135,N_6356,N_9256);
and UO_136 (O_136,N_7597,N_6850);
or UO_137 (O_137,N_7089,N_8107);
or UO_138 (O_138,N_8106,N_9066);
xnor UO_139 (O_139,N_8882,N_6015);
and UO_140 (O_140,N_7184,N_9612);
or UO_141 (O_141,N_7120,N_6144);
xor UO_142 (O_142,N_6874,N_6368);
or UO_143 (O_143,N_8198,N_5309);
nor UO_144 (O_144,N_9584,N_5215);
or UO_145 (O_145,N_6758,N_9623);
nand UO_146 (O_146,N_9714,N_9234);
or UO_147 (O_147,N_5859,N_6606);
or UO_148 (O_148,N_6433,N_8181);
nand UO_149 (O_149,N_7729,N_8997);
xnor UO_150 (O_150,N_8756,N_8283);
nor UO_151 (O_151,N_5496,N_7239);
nand UO_152 (O_152,N_8856,N_9848);
xor UO_153 (O_153,N_6910,N_9062);
or UO_154 (O_154,N_6532,N_6507);
or UO_155 (O_155,N_9231,N_8418);
xnor UO_156 (O_156,N_9615,N_6455);
xor UO_157 (O_157,N_6304,N_5838);
and UO_158 (O_158,N_7806,N_9224);
nor UO_159 (O_159,N_9046,N_6623);
nand UO_160 (O_160,N_5520,N_9103);
and UO_161 (O_161,N_5034,N_5618);
nor UO_162 (O_162,N_9493,N_5074);
nand UO_163 (O_163,N_5738,N_7855);
nor UO_164 (O_164,N_6334,N_9161);
and UO_165 (O_165,N_9815,N_8509);
nor UO_166 (O_166,N_7888,N_5622);
or UO_167 (O_167,N_7759,N_6472);
and UO_168 (O_168,N_8007,N_9279);
xor UO_169 (O_169,N_7531,N_5256);
or UO_170 (O_170,N_7433,N_7684);
xor UO_171 (O_171,N_6538,N_9828);
or UO_172 (O_172,N_5124,N_5163);
and UO_173 (O_173,N_5821,N_6505);
xor UO_174 (O_174,N_9542,N_7687);
nand UO_175 (O_175,N_7748,N_5355);
nand UO_176 (O_176,N_7805,N_7828);
or UO_177 (O_177,N_7882,N_8518);
and UO_178 (O_178,N_6794,N_8924);
and UO_179 (O_179,N_5408,N_7901);
xnor UO_180 (O_180,N_6219,N_7722);
nor UO_181 (O_181,N_7432,N_6425);
or UO_182 (O_182,N_5729,N_6718);
xnor UO_183 (O_183,N_9470,N_5996);
nand UO_184 (O_184,N_5154,N_9672);
nor UO_185 (O_185,N_7985,N_7650);
xnor UO_186 (O_186,N_9110,N_9019);
or UO_187 (O_187,N_9393,N_7491);
or UO_188 (O_188,N_5188,N_5447);
nor UO_189 (O_189,N_9358,N_6935);
xnor UO_190 (O_190,N_8374,N_8657);
or UO_191 (O_191,N_9697,N_8089);
nor UO_192 (O_192,N_9933,N_7428);
nor UO_193 (O_193,N_5575,N_5579);
xor UO_194 (O_194,N_5440,N_9665);
or UO_195 (O_195,N_6487,N_8564);
and UO_196 (O_196,N_9491,N_8692);
or UO_197 (O_197,N_9794,N_7671);
xor UO_198 (O_198,N_8479,N_8468);
or UO_199 (O_199,N_9375,N_7253);
or UO_200 (O_200,N_7642,N_5707);
and UO_201 (O_201,N_6441,N_9561);
nor UO_202 (O_202,N_7065,N_9890);
nor UO_203 (O_203,N_6645,N_5468);
and UO_204 (O_204,N_8315,N_9645);
or UO_205 (O_205,N_9984,N_8140);
xor UO_206 (O_206,N_5600,N_9600);
xor UO_207 (O_207,N_8275,N_8012);
or UO_208 (O_208,N_9902,N_6918);
nor UO_209 (O_209,N_6655,N_5898);
and UO_210 (O_210,N_6525,N_7744);
or UO_211 (O_211,N_8400,N_9755);
or UO_212 (O_212,N_5075,N_8027);
nand UO_213 (O_213,N_7105,N_8169);
or UO_214 (O_214,N_9463,N_9364);
nand UO_215 (O_215,N_6814,N_9883);
or UO_216 (O_216,N_9340,N_7922);
and UO_217 (O_217,N_5873,N_9076);
nor UO_218 (O_218,N_5219,N_8122);
and UO_219 (O_219,N_5286,N_8336);
nand UO_220 (O_220,N_9720,N_7669);
nand UO_221 (O_221,N_5592,N_6521);
and UO_222 (O_222,N_9376,N_8332);
or UO_223 (O_223,N_7466,N_7568);
nand UO_224 (O_224,N_9326,N_6785);
nand UO_225 (O_225,N_7886,N_5503);
and UO_226 (O_226,N_5663,N_9291);
and UO_227 (O_227,N_8735,N_9464);
or UO_228 (O_228,N_6119,N_9614);
nand UO_229 (O_229,N_8695,N_6772);
nor UO_230 (O_230,N_7580,N_5312);
nor UO_231 (O_231,N_5923,N_8949);
nor UO_232 (O_232,N_5176,N_6030);
nand UO_233 (O_233,N_8710,N_5885);
xnor UO_234 (O_234,N_7318,N_7145);
xnor UO_235 (O_235,N_8172,N_7357);
xnor UO_236 (O_236,N_7136,N_5884);
nand UO_237 (O_237,N_5987,N_8585);
and UO_238 (O_238,N_5876,N_5820);
xnor UO_239 (O_239,N_9479,N_5546);
and UO_240 (O_240,N_6709,N_5766);
nand UO_241 (O_241,N_9251,N_7753);
xnor UO_242 (O_242,N_6225,N_5513);
nor UO_243 (O_243,N_5413,N_6945);
and UO_244 (O_244,N_6469,N_8101);
and UO_245 (O_245,N_7817,N_5457);
xor UO_246 (O_246,N_5537,N_8321);
and UO_247 (O_247,N_6667,N_7129);
xor UO_248 (O_248,N_9637,N_6527);
xnor UO_249 (O_249,N_8260,N_7946);
and UO_250 (O_250,N_5775,N_5002);
xor UO_251 (O_251,N_6313,N_5220);
or UO_252 (O_252,N_5536,N_7328);
or UO_253 (O_253,N_7356,N_8245);
nand UO_254 (O_254,N_7571,N_9009);
and UO_255 (O_255,N_6907,N_9669);
nand UO_256 (O_256,N_6687,N_6351);
or UO_257 (O_257,N_9888,N_7030);
nor UO_258 (O_258,N_6023,N_8668);
or UO_259 (O_259,N_9630,N_8566);
nor UO_260 (O_260,N_6031,N_9932);
xor UO_261 (O_261,N_7386,N_9539);
nand UO_262 (O_262,N_9075,N_9721);
nand UO_263 (O_263,N_5001,N_8591);
xor UO_264 (O_264,N_9746,N_6617);
or UO_265 (O_265,N_5336,N_6293);
xor UO_266 (O_266,N_6159,N_7225);
and UO_267 (O_267,N_8737,N_5205);
or UO_268 (O_268,N_5173,N_7283);
and UO_269 (O_269,N_6210,N_9116);
xor UO_270 (O_270,N_9860,N_9253);
nand UO_271 (O_271,N_7102,N_5589);
and UO_272 (O_272,N_6870,N_5169);
nor UO_273 (O_273,N_6746,N_7942);
nor UO_274 (O_274,N_7630,N_6893);
and UO_275 (O_275,N_6685,N_8829);
nor UO_276 (O_276,N_6835,N_6021);
or UO_277 (O_277,N_5068,N_7477);
or UO_278 (O_278,N_7431,N_7191);
and UO_279 (O_279,N_9499,N_7809);
or UO_280 (O_280,N_8781,N_9719);
nand UO_281 (O_281,N_9701,N_8648);
xnor UO_282 (O_282,N_5144,N_5225);
nand UO_283 (O_283,N_9710,N_6926);
nand UO_284 (O_284,N_5675,N_7308);
or UO_285 (O_285,N_8947,N_8633);
nand UO_286 (O_286,N_5211,N_7411);
nor UO_287 (O_287,N_6384,N_7407);
nand UO_288 (O_288,N_8644,N_7099);
or UO_289 (O_289,N_8076,N_8397);
and UO_290 (O_290,N_5921,N_9591);
xnor UO_291 (O_291,N_8623,N_5796);
nand UO_292 (O_292,N_9903,N_5209);
or UO_293 (O_293,N_6247,N_8047);
or UO_294 (O_294,N_5416,N_6588);
nor UO_295 (O_295,N_5011,N_7521);
or UO_296 (O_296,N_9944,N_7220);
or UO_297 (O_297,N_7440,N_7137);
nand UO_298 (O_298,N_5610,N_9693);
or UO_299 (O_299,N_5508,N_5802);
xor UO_300 (O_300,N_5351,N_5896);
nand UO_301 (O_301,N_5037,N_9064);
and UO_302 (O_302,N_5102,N_8459);
xor UO_303 (O_303,N_7314,N_6541);
nor UO_304 (O_304,N_5132,N_5869);
xnor UO_305 (O_305,N_8294,N_6971);
nor UO_306 (O_306,N_6187,N_9570);
nor UO_307 (O_307,N_6289,N_7042);
and UO_308 (O_308,N_5814,N_6462);
nand UO_309 (O_309,N_5893,N_9682);
xor UO_310 (O_310,N_6492,N_6526);
xor UO_311 (O_311,N_7877,N_5450);
xnor UO_312 (O_312,N_7588,N_5396);
nand UO_313 (O_313,N_7649,N_5510);
nand UO_314 (O_314,N_5822,N_6083);
and UO_315 (O_315,N_8840,N_9218);
nor UO_316 (O_316,N_6004,N_7598);
xnor UO_317 (O_317,N_8000,N_8767);
and UO_318 (O_318,N_5800,N_6235);
or UO_319 (O_319,N_7453,N_5322);
nand UO_320 (O_320,N_8144,N_9105);
nand UO_321 (O_321,N_6714,N_9332);
nand UO_322 (O_322,N_9760,N_5961);
xnor UO_323 (O_323,N_9038,N_7664);
or UO_324 (O_324,N_8330,N_6892);
nand UO_325 (O_325,N_9245,N_6244);
nor UO_326 (O_326,N_6039,N_6997);
or UO_327 (O_327,N_8335,N_5784);
and UO_328 (O_328,N_9045,N_6127);
or UO_329 (O_329,N_9192,N_9538);
or UO_330 (O_330,N_7778,N_8839);
and UO_331 (O_331,N_5326,N_9195);
or UO_332 (O_332,N_8086,N_6554);
nor UO_333 (O_333,N_7857,N_5039);
or UO_334 (O_334,N_6885,N_5179);
xnor UO_335 (O_335,N_8138,N_5390);
or UO_336 (O_336,N_9777,N_5701);
and UO_337 (O_337,N_5544,N_9492);
nor UO_338 (O_338,N_6958,N_6138);
xor UO_339 (O_339,N_8721,N_8129);
xor UO_340 (O_340,N_5453,N_6952);
nand UO_341 (O_341,N_9951,N_6443);
or UO_342 (O_342,N_7773,N_9363);
and UO_343 (O_343,N_8409,N_8358);
xor UO_344 (O_344,N_8466,N_8945);
or UO_345 (O_345,N_9718,N_6765);
xnor UO_346 (O_346,N_9061,N_5651);
and UO_347 (O_347,N_7181,N_9833);
nor UO_348 (O_348,N_9982,N_6435);
nand UO_349 (O_349,N_6343,N_6125);
and UO_350 (O_350,N_5829,N_7299);
xor UO_351 (O_351,N_8257,N_5978);
xor UO_352 (O_352,N_8080,N_6209);
nand UO_353 (O_353,N_5538,N_7288);
xnor UO_354 (O_354,N_6158,N_8376);
xor UO_355 (O_355,N_7845,N_7320);
xnor UO_356 (O_356,N_7106,N_5501);
or UO_357 (O_357,N_8480,N_8975);
nand UO_358 (O_358,N_7032,N_7697);
nor UO_359 (O_359,N_9310,N_7844);
nor UO_360 (O_360,N_8427,N_5623);
nor UO_361 (O_361,N_9737,N_8211);
xnor UO_362 (O_362,N_9901,N_9990);
xor UO_363 (O_363,N_8532,N_6195);
nor UO_364 (O_364,N_7992,N_6402);
nor UO_365 (O_365,N_9985,N_9799);
nand UO_366 (O_366,N_9086,N_6741);
and UO_367 (O_367,N_8083,N_7952);
and UO_368 (O_368,N_7380,N_7950);
and UO_369 (O_369,N_9441,N_6939);
xor UO_370 (O_370,N_5988,N_8837);
and UO_371 (O_371,N_9181,N_5422);
xnor UO_372 (O_372,N_7090,N_9415);
xor UO_373 (O_373,N_7843,N_8697);
nand UO_374 (O_374,N_7473,N_8915);
nor UO_375 (O_375,N_7909,N_6180);
and UO_376 (O_376,N_5276,N_8327);
nand UO_377 (O_377,N_5625,N_9677);
nor UO_378 (O_378,N_6387,N_9102);
nor UO_379 (O_379,N_5128,N_5409);
nand UO_380 (O_380,N_7295,N_5035);
nand UO_381 (O_381,N_7726,N_5816);
nor UO_382 (O_382,N_9771,N_5582);
nor UO_383 (O_383,N_5719,N_9140);
xor UO_384 (O_384,N_6727,N_7127);
nand UO_385 (O_385,N_6236,N_5492);
or UO_386 (O_386,N_6294,N_6517);
xor UO_387 (O_387,N_5725,N_9077);
and UO_388 (O_388,N_5227,N_7119);
and UO_389 (O_389,N_7418,N_8860);
or UO_390 (O_390,N_8157,N_9858);
nand UO_391 (O_391,N_5594,N_5755);
or UO_392 (O_392,N_7036,N_8378);
nand UO_393 (O_393,N_7250,N_7768);
nand UO_394 (O_394,N_7410,N_6038);
nand UO_395 (O_395,N_8164,N_8683);
and UO_396 (O_396,N_5364,N_7767);
or UO_397 (O_397,N_6624,N_5648);
nand UO_398 (O_398,N_9829,N_7501);
nor UO_399 (O_399,N_6396,N_5653);
or UO_400 (O_400,N_5509,N_8326);
xnor UO_401 (O_401,N_8290,N_8116);
or UO_402 (O_402,N_6733,N_5608);
and UO_403 (O_403,N_6327,N_5439);
or UO_404 (O_404,N_9184,N_8222);
xor UO_405 (O_405,N_6171,N_6690);
nor UO_406 (O_406,N_9359,N_6493);
nand UO_407 (O_407,N_6246,N_9172);
nand UO_408 (O_408,N_6362,N_5152);
xnor UO_409 (O_409,N_5529,N_7894);
xnor UO_410 (O_410,N_8857,N_6328);
nand UO_411 (O_411,N_5819,N_7416);
xnor UO_412 (O_412,N_7756,N_6194);
and UO_413 (O_413,N_9347,N_9704);
and UO_414 (O_414,N_7995,N_9031);
and UO_415 (O_415,N_7245,N_5926);
nand UO_416 (O_416,N_6987,N_7096);
and UO_417 (O_417,N_9210,N_8478);
xnor UO_418 (O_418,N_5028,N_6796);
and UO_419 (O_419,N_8897,N_5055);
nor UO_420 (O_420,N_5789,N_9395);
and UO_421 (O_421,N_8236,N_8794);
nor UO_422 (O_422,N_8075,N_6990);
and UO_423 (O_423,N_7790,N_7391);
nor UO_424 (O_424,N_5723,N_9717);
and UO_425 (O_425,N_7178,N_6186);
or UO_426 (O_426,N_5681,N_7011);
or UO_427 (O_427,N_8320,N_7093);
or UO_428 (O_428,N_6752,N_5338);
nor UO_429 (O_429,N_9662,N_5178);
xnor UO_430 (O_430,N_8180,N_9243);
or UO_431 (O_431,N_8185,N_8004);
and UO_432 (O_432,N_5299,N_9647);
nor UO_433 (O_433,N_8660,N_6734);
xor UO_434 (O_434,N_7376,N_7213);
nand UO_435 (O_435,N_8853,N_6913);
or UO_436 (O_436,N_7587,N_6009);
xnor UO_437 (O_437,N_7638,N_7060);
nor UO_438 (O_438,N_6991,N_6827);
or UO_439 (O_439,N_9355,N_7541);
or UO_440 (O_440,N_9793,N_5391);
xnor UO_441 (O_441,N_7476,N_8599);
and UO_442 (O_442,N_7153,N_6416);
nor UO_443 (O_443,N_7755,N_5187);
or UO_444 (O_444,N_7975,N_8749);
or UO_445 (O_445,N_6622,N_7944);
xnor UO_446 (O_446,N_6112,N_8392);
nand UO_447 (O_447,N_8064,N_8733);
or UO_448 (O_448,N_5319,N_5848);
or UO_449 (O_449,N_7115,N_5429);
xnor UO_450 (O_450,N_5105,N_6681);
xnor UO_451 (O_451,N_9548,N_9633);
xnor UO_452 (O_452,N_5938,N_5314);
nor UO_453 (O_453,N_6592,N_5772);
and UO_454 (O_454,N_8583,N_5882);
nor UO_455 (O_455,N_6040,N_5750);
and UO_456 (O_456,N_9652,N_6488);
and UO_457 (O_457,N_8928,N_8344);
xnor UO_458 (O_458,N_5092,N_6214);
xnor UO_459 (O_459,N_8736,N_7034);
and UO_460 (O_460,N_6562,N_5712);
or UO_461 (O_461,N_8341,N_6431);
xor UO_462 (O_462,N_8790,N_8974);
and UO_463 (O_463,N_5021,N_6565);
or UO_464 (O_464,N_5619,N_5682);
or UO_465 (O_465,N_7287,N_9502);
and UO_466 (O_466,N_5399,N_7164);
nand UO_467 (O_467,N_6181,N_7117);
nor UO_468 (O_468,N_5274,N_8824);
nor UO_469 (O_469,N_6400,N_7791);
and UO_470 (O_470,N_7683,N_9817);
nor UO_471 (O_471,N_6296,N_9457);
xnor UO_472 (O_472,N_9572,N_5082);
xnor UO_473 (O_473,N_8987,N_9169);
nand UO_474 (O_474,N_8343,N_7919);
nand UO_475 (O_475,N_9506,N_8604);
nand UO_476 (O_476,N_9190,N_9320);
or UO_477 (O_477,N_9480,N_8707);
xnor UO_478 (O_478,N_9469,N_6899);
nand UO_479 (O_479,N_7923,N_8149);
xnor UO_480 (O_480,N_8018,N_8815);
or UO_481 (O_481,N_5315,N_9178);
and UO_482 (O_482,N_6231,N_9128);
nor UO_483 (O_483,N_9562,N_8937);
and UO_484 (O_484,N_5568,N_9130);
and UO_485 (O_485,N_5009,N_9943);
nor UO_486 (O_486,N_9955,N_7050);
xnor UO_487 (O_487,N_9176,N_6692);
nand UO_488 (O_488,N_7567,N_6331);
or UO_489 (O_489,N_6684,N_6405);
nand UO_490 (O_490,N_7856,N_5677);
or UO_491 (O_491,N_7272,N_7656);
nor UO_492 (O_492,N_5664,N_6230);
or UO_493 (O_493,N_9481,N_9205);
nand UO_494 (O_494,N_6216,N_7949);
or UO_495 (O_495,N_9139,N_9087);
and UO_496 (O_496,N_5385,N_8395);
xor UO_497 (O_497,N_9892,N_9808);
xor UO_498 (O_498,N_8879,N_9642);
xor UO_499 (O_499,N_5052,N_6921);
or UO_500 (O_500,N_9421,N_8655);
or UO_501 (O_501,N_9574,N_7745);
and UO_502 (O_502,N_9357,N_9910);
xor UO_503 (O_503,N_7540,N_9617);
xnor UO_504 (O_504,N_8784,N_6735);
xor UO_505 (O_505,N_5785,N_8884);
or UO_506 (O_506,N_7518,N_6082);
xnor UO_507 (O_507,N_6050,N_8747);
nand UO_508 (O_508,N_5686,N_9476);
and UO_509 (O_509,N_9800,N_7769);
nand UO_510 (O_510,N_8301,N_5298);
nor UO_511 (O_511,N_6868,N_8942);
nand UO_512 (O_512,N_9227,N_7594);
or UO_513 (O_513,N_7757,N_9043);
and UO_514 (O_514,N_8610,N_8676);
nor UO_515 (O_515,N_9072,N_9189);
and UO_516 (O_516,N_7182,N_7086);
nor UO_517 (O_517,N_5375,N_7972);
or UO_518 (O_518,N_6743,N_6555);
and UO_519 (O_519,N_8780,N_7599);
or UO_520 (O_520,N_7291,N_5428);
xnor UO_521 (O_521,N_6196,N_9822);
or UO_522 (O_522,N_6392,N_6949);
xnor UO_523 (O_523,N_9567,N_5657);
nand UO_524 (O_524,N_7576,N_5140);
xnor UO_525 (O_525,N_6041,N_6804);
nor UO_526 (O_526,N_6867,N_6891);
or UO_527 (O_527,N_7274,N_9995);
or UO_528 (O_528,N_5202,N_6270);
or UO_529 (O_529,N_9965,N_7359);
xor UO_530 (O_530,N_8622,N_6084);
nand UO_531 (O_531,N_8133,N_6122);
or UO_532 (O_532,N_9583,N_7135);
xnor UO_533 (O_533,N_7400,N_6113);
nand UO_534 (O_534,N_5159,N_6070);
and UO_535 (O_535,N_7794,N_5139);
nand UO_536 (O_536,N_8340,N_8577);
or UO_537 (O_537,N_7674,N_5778);
nand UO_538 (O_538,N_7825,N_6459);
xor UO_539 (O_539,N_7061,N_8337);
or UO_540 (O_540,N_9027,N_6386);
or UO_541 (O_541,N_7517,N_5767);
and UO_542 (O_542,N_6053,N_6375);
nand UO_543 (O_543,N_6197,N_5555);
nor UO_544 (O_544,N_7373,N_9987);
xnor UO_545 (O_545,N_9809,N_6484);
nor UO_546 (O_546,N_9294,N_6243);
and UO_547 (O_547,N_7506,N_6774);
nand UO_548 (O_548,N_7375,N_9708);
or UO_549 (O_549,N_9148,N_8732);
nor UO_550 (O_550,N_6121,N_6420);
xor UO_551 (O_551,N_7647,N_5547);
nand UO_552 (O_552,N_7471,N_8394);
xor UO_553 (O_553,N_5901,N_7342);
nor UO_554 (O_554,N_8241,N_5954);
and UO_555 (O_555,N_8331,N_7365);
and UO_556 (O_556,N_6146,N_8291);
nor UO_557 (O_557,N_9611,N_8196);
nand UO_558 (O_558,N_9168,N_7895);
nor UO_559 (O_559,N_6572,N_6656);
and UO_560 (O_560,N_7924,N_8220);
xnor UO_561 (O_561,N_5649,N_8024);
nand UO_562 (O_562,N_6495,N_5203);
xnor UO_563 (O_563,N_8524,N_9571);
xnor UO_564 (O_564,N_6584,N_6295);
xor UO_565 (O_565,N_9767,N_6789);
or UO_566 (O_566,N_8445,N_5295);
or UO_567 (O_567,N_9475,N_5526);
or UO_568 (O_568,N_5015,N_6252);
and UO_569 (O_569,N_5525,N_7596);
nand UO_570 (O_570,N_9092,N_9125);
nor UO_571 (O_571,N_5488,N_6522);
and UO_572 (O_572,N_7750,N_9880);
or UO_573 (O_573,N_8350,N_7091);
nor UO_574 (O_574,N_6621,N_9980);
nor UO_575 (O_575,N_5656,N_6806);
or UO_576 (O_576,N_9654,N_9278);
and UO_577 (O_577,N_8960,N_5229);
or UO_578 (O_578,N_8297,N_9290);
or UO_579 (O_579,N_8213,N_5459);
xnor UO_580 (O_580,N_5691,N_9772);
or UO_581 (O_581,N_5019,N_6988);
and UO_582 (O_582,N_9444,N_6845);
nor UO_583 (O_583,N_6206,N_7193);
and UO_584 (O_584,N_7704,N_7557);
xnor UO_585 (O_585,N_5290,N_9813);
or UO_586 (O_586,N_9774,N_9864);
or UO_587 (O_587,N_5191,N_8218);
xnor UO_588 (O_588,N_5780,N_5210);
xnor UO_589 (O_589,N_9814,N_7377);
or UO_590 (O_590,N_6093,N_7730);
and UO_591 (O_591,N_9518,N_5740);
and UO_592 (O_592,N_6799,N_9795);
or UO_593 (O_593,N_5757,N_9465);
xor UO_594 (O_594,N_5155,N_6871);
xor UO_595 (O_595,N_9723,N_5585);
nand UO_596 (O_596,N_7873,N_9535);
nor UO_597 (O_597,N_7631,N_8100);
or UO_598 (O_598,N_8233,N_5437);
and UO_599 (O_599,N_5073,N_5017);
nand UO_600 (O_600,N_6344,N_6768);
nor UO_601 (O_601,N_5558,N_9924);
xor UO_602 (O_602,N_7885,N_7675);
xnor UO_603 (O_603,N_8084,N_5104);
or UO_604 (O_604,N_9284,N_6880);
xor UO_605 (O_605,N_7670,N_6863);
nor UO_606 (O_606,N_5317,N_5557);
nand UO_607 (O_607,N_7300,N_8148);
or UO_608 (O_608,N_7689,N_7074);
nor UO_609 (O_609,N_5484,N_6155);
nand UO_610 (O_610,N_5078,N_5662);
or UO_611 (O_611,N_5942,N_8651);
nand UO_612 (O_612,N_6464,N_5523);
and UO_613 (O_613,N_8132,N_8186);
nand UO_614 (O_614,N_8789,N_6160);
nor UO_615 (O_615,N_7370,N_5242);
nor UO_616 (O_616,N_6762,N_7133);
or UO_617 (O_617,N_7080,N_5402);
nand UO_618 (O_618,N_6887,N_7716);
or UO_619 (O_619,N_6558,N_7167);
nand UO_620 (O_620,N_9471,N_5631);
xnor UO_621 (O_621,N_6797,N_9659);
or UO_622 (O_622,N_5182,N_5903);
nor UO_623 (O_623,N_9968,N_9656);
xor UO_624 (O_624,N_6745,N_6498);
and UO_625 (O_625,N_8663,N_7481);
xnor UO_626 (O_626,N_5974,N_6831);
nor UO_627 (O_627,N_5634,N_7911);
xor UO_628 (O_628,N_7026,N_9724);
xor UO_629 (O_629,N_9252,N_5698);
nor UO_630 (O_630,N_5540,N_7935);
xor UO_631 (O_631,N_7269,N_9117);
and UO_632 (O_632,N_5703,N_5161);
nor UO_633 (O_633,N_9208,N_8771);
nor UO_634 (O_634,N_5883,N_5670);
nor UO_635 (O_635,N_9032,N_9706);
and UO_636 (O_636,N_7292,N_5790);
and UO_637 (O_637,N_5639,N_9629);
nor UO_638 (O_638,N_6940,N_8010);
nor UO_639 (O_639,N_8264,N_7190);
and UO_640 (O_640,N_7205,N_9626);
and UO_641 (O_641,N_6157,N_9628);
xnor UO_642 (O_642,N_8907,N_8594);
nor UO_643 (O_643,N_5230,N_9300);
nand UO_644 (O_644,N_6148,N_6760);
xnor UO_645 (O_645,N_7820,N_5380);
xor UO_646 (O_646,N_9857,N_7971);
nand UO_647 (O_647,N_8410,N_9592);
or UO_648 (O_648,N_6641,N_6519);
nand UO_649 (O_649,N_8576,N_9791);
nor UO_650 (O_650,N_6757,N_5997);
xor UO_651 (O_651,N_7887,N_7615);
or UO_652 (O_652,N_6736,N_5512);
nor UO_653 (O_653,N_8307,N_9769);
nor UO_654 (O_654,N_8382,N_8624);
xnor UO_655 (O_655,N_5348,N_8489);
xnor UO_656 (O_656,N_7991,N_6169);
xor UO_657 (O_657,N_5419,N_9578);
xnor UO_658 (O_658,N_6618,N_5204);
nand UO_659 (O_659,N_7027,N_8543);
and UO_660 (O_660,N_8216,N_9632);
nor UO_661 (O_661,N_5093,N_7500);
and UO_662 (O_662,N_7538,N_7363);
nand UO_663 (O_663,N_8911,N_9945);
nand UO_664 (O_664,N_8708,N_8588);
or UO_665 (O_665,N_5414,N_7737);
or UO_666 (O_666,N_8467,N_6784);
nor UO_667 (O_667,N_9348,N_7235);
and UO_668 (O_668,N_9016,N_7302);
nand UO_669 (O_669,N_5665,N_7760);
xor UO_670 (O_670,N_6346,N_6840);
or UO_671 (O_671,N_9250,N_5949);
nor UO_672 (O_672,N_9651,N_6756);
nand UO_673 (O_673,N_6372,N_7112);
nor UO_674 (O_674,N_6489,N_8215);
xnor UO_675 (O_675,N_9037,N_7486);
or UO_676 (O_676,N_7325,N_5121);
or UO_677 (O_677,N_6250,N_8927);
or UO_678 (O_678,N_8495,N_9619);
xor UO_679 (O_679,N_9528,N_5910);
and UO_680 (O_680,N_5194,N_8855);
nor UO_681 (O_681,N_7189,N_7678);
and UO_682 (O_682,N_7326,N_9802);
nand UO_683 (O_683,N_5240,N_9937);
and UO_684 (O_684,N_9899,N_7921);
xor UO_685 (O_685,N_7262,N_5018);
or UO_686 (O_686,N_6803,N_7343);
xnor UO_687 (O_687,N_5195,N_8764);
nand UO_688 (O_688,N_9732,N_8414);
nor UO_689 (O_689,N_8154,N_9033);
nand UO_690 (O_690,N_9030,N_6027);
and UO_691 (O_691,N_6208,N_6139);
or UO_692 (O_692,N_7612,N_5050);
xor UO_693 (O_693,N_9183,N_8217);
nand UO_694 (O_694,N_8966,N_8972);
nor UO_695 (O_695,N_6130,N_7475);
or UO_696 (O_696,N_9573,N_9309);
nor UO_697 (O_697,N_5040,N_6675);
nand UO_698 (O_698,N_7641,N_5952);
or UO_699 (O_699,N_5920,N_6321);
or UO_700 (O_700,N_7268,N_7384);
nor UO_701 (O_701,N_9966,N_6682);
xnor UO_702 (O_702,N_9859,N_8994);
or UO_703 (O_703,N_9764,N_6035);
or UO_704 (O_704,N_9285,N_5925);
and UO_705 (O_705,N_7542,N_8609);
and UO_706 (O_706,N_5899,N_9563);
xor UO_707 (O_707,N_9973,N_9523);
xnor UO_708 (O_708,N_9365,N_6977);
and UO_709 (O_709,N_6602,N_8689);
nor UO_710 (O_710,N_7159,N_9145);
nor UO_711 (O_711,N_5823,N_7022);
or UO_712 (O_712,N_9707,N_8760);
xnor UO_713 (O_713,N_7313,N_9409);
or UO_714 (O_714,N_7197,N_5304);
xnor UO_715 (O_715,N_9141,N_6314);
nor UO_716 (O_716,N_8303,N_8237);
nand UO_717 (O_717,N_7364,N_7963);
xor UO_718 (O_718,N_9018,N_5311);
and UO_719 (O_719,N_5228,N_6626);
or UO_720 (O_720,N_8731,N_8051);
xor UO_721 (O_721,N_9505,N_6693);
xnor UO_722 (O_722,N_9089,N_6672);
nand UO_723 (O_723,N_9534,N_9453);
nand UO_724 (O_724,N_9936,N_9156);
and UO_725 (O_725,N_5445,N_7176);
xor UO_726 (O_726,N_5872,N_9000);
or UO_727 (O_727,N_9370,N_7548);
xnor UO_728 (O_728,N_6499,N_5342);
and UO_729 (O_729,N_5281,N_7927);
and UO_730 (O_730,N_5716,N_8439);
nor UO_731 (O_731,N_7408,N_7577);
and UO_732 (O_732,N_9070,N_5495);
and UO_733 (O_733,N_6120,N_9604);
or UO_734 (O_734,N_6237,N_9366);
and UO_735 (O_735,N_5565,N_5635);
nor UO_736 (O_736,N_9426,N_8191);
xor UO_737 (O_737,N_9610,N_8540);
nor UO_738 (O_738,N_7008,N_7323);
xor UO_739 (O_739,N_9108,N_8694);
and UO_740 (O_740,N_6544,N_7854);
and UO_741 (O_741,N_6916,N_7338);
nand UO_742 (O_742,N_9186,N_8255);
and UO_743 (O_743,N_8464,N_5250);
nand UO_744 (O_744,N_8465,N_5174);
xor UO_745 (O_745,N_6638,N_8687);
or UO_746 (O_746,N_5109,N_9589);
xnor UO_747 (O_747,N_6824,N_5946);
or UO_748 (O_748,N_6860,N_7427);
and UO_749 (O_749,N_9422,N_7429);
xnor UO_750 (O_750,N_9472,N_7994);
and UO_751 (O_751,N_8440,N_5237);
nor UO_752 (O_752,N_9551,N_5837);
xor UO_753 (O_753,N_7254,N_5931);
nor UO_754 (O_754,N_6722,N_6931);
and UO_755 (O_755,N_5661,N_5079);
or UO_756 (O_756,N_6142,N_7483);
nand UO_757 (O_757,N_5687,N_6494);
xor UO_758 (O_758,N_7698,N_6808);
nand UO_759 (O_759,N_9272,N_5543);
or UO_760 (O_760,N_7160,N_7686);
or UO_761 (O_761,N_5517,N_5062);
or UO_762 (O_762,N_8617,N_9569);
nor UO_763 (O_763,N_7943,N_9219);
xnor UO_764 (O_764,N_7695,N_8529);
and UO_765 (O_765,N_7140,N_6635);
nor UO_766 (O_766,N_9852,N_9362);
nor UO_767 (O_767,N_8150,N_9484);
nand UO_768 (O_768,N_8888,N_8770);
nand UO_769 (O_769,N_9048,N_6578);
nand UO_770 (O_770,N_9687,N_9265);
nor UO_771 (O_771,N_7969,N_5016);
and UO_772 (O_772,N_6843,N_5982);
and UO_773 (O_773,N_8964,N_7423);
nand UO_774 (O_774,N_9352,N_6500);
and UO_775 (O_775,N_8057,N_7665);
nor UO_776 (O_776,N_5257,N_7088);
and UO_777 (O_777,N_9670,N_6332);
and UO_778 (O_778,N_7772,N_6518);
nor UO_779 (O_779,N_8940,N_6864);
nor UO_780 (O_780,N_6337,N_9407);
xor UO_781 (O_781,N_5889,N_5005);
nand UO_782 (O_782,N_8077,N_6613);
xnor UO_783 (O_783,N_8698,N_6890);
xor UO_784 (O_784,N_9920,N_7020);
nand UO_785 (O_785,N_8658,N_8184);
or UO_786 (O_786,N_6223,N_9898);
and UO_787 (O_787,N_5198,N_8199);
nor UO_788 (O_788,N_7814,N_5113);
and UO_789 (O_789,N_6066,N_9552);
or UO_790 (O_790,N_8114,N_5120);
nor UO_791 (O_791,N_6454,N_5280);
nor UO_792 (O_792,N_9106,N_9531);
or UO_793 (O_793,N_9374,N_7092);
nor UO_794 (O_794,N_7261,N_6465);
or UO_795 (O_795,N_6257,N_7394);
nand UO_796 (O_796,N_7604,N_7563);
nand UO_797 (O_797,N_6202,N_7263);
and UO_798 (O_798,N_5854,N_9927);
and UO_799 (O_799,N_6659,N_9237);
nor UO_800 (O_800,N_7108,N_5799);
or UO_801 (O_801,N_8557,N_9993);
xor UO_802 (O_802,N_8590,N_9931);
nand UO_803 (O_803,N_6434,N_6315);
nand UO_804 (O_804,N_6064,N_7574);
nor UO_805 (O_805,N_8171,N_7707);
nor UO_806 (O_806,N_9372,N_8008);
and UO_807 (O_807,N_7528,N_5273);
or UO_808 (O_808,N_6201,N_5818);
and UO_809 (O_809,N_6523,N_5781);
and UO_810 (O_810,N_9071,N_7987);
or UO_811 (O_811,N_8050,N_7712);
and UO_812 (O_812,N_5521,N_8862);
nor UO_813 (O_813,N_9211,N_6274);
nor UO_814 (O_814,N_9646,N_6056);
and UO_815 (O_815,N_7654,N_8598);
nor UO_816 (O_816,N_9942,N_7212);
or UO_817 (O_817,N_7267,N_8032);
nor UO_818 (O_818,N_9674,N_6357);
and UO_819 (O_819,N_8182,N_6711);
nand UO_820 (O_820,N_6085,N_9991);
and UO_821 (O_821,N_9603,N_7264);
or UO_822 (O_822,N_6251,N_8475);
and UO_823 (O_823,N_6037,N_8558);
and UO_824 (O_824,N_9095,N_6668);
or UO_825 (O_825,N_7786,N_8379);
or UO_826 (O_826,N_7382,N_7713);
nand UO_827 (O_827,N_9158,N_8244);
xor UO_828 (O_828,N_5856,N_6838);
nor UO_829 (O_829,N_6754,N_9975);
nor UO_830 (O_830,N_5477,N_8723);
xnor UO_831 (O_831,N_9241,N_5654);
or UO_832 (O_832,N_7570,N_6068);
or UO_833 (O_833,N_9702,N_5810);
or UO_834 (O_834,N_8234,N_9180);
and UO_835 (O_835,N_7774,N_6530);
nor UO_836 (O_836,N_8167,N_5735);
nor UO_837 (O_837,N_6528,N_5367);
nor UO_838 (O_838,N_5955,N_7907);
or UO_839 (O_839,N_6470,N_8841);
and UO_840 (O_840,N_6222,N_7661);
xnor UO_841 (O_841,N_7077,N_6999);
nand UO_842 (O_842,N_9221,N_9338);
or UO_843 (O_843,N_7172,N_6170);
or UO_844 (O_844,N_8755,N_5966);
xor UO_845 (O_845,N_9164,N_7508);
or UO_846 (O_846,N_9097,N_6205);
xor UO_847 (O_847,N_8843,N_5676);
and UO_848 (O_848,N_6081,N_6568);
nor UO_849 (O_849,N_6801,N_6399);
or UO_850 (O_850,N_9053,N_8659);
xor UO_851 (O_851,N_8253,N_9959);
nand UO_852 (O_852,N_9754,N_5699);
nand UO_853 (O_853,N_7910,N_9057);
and UO_854 (O_854,N_6013,N_9891);
xnor UO_855 (O_855,N_8587,N_8542);
nand UO_856 (O_856,N_7260,N_9850);
nand UO_857 (O_857,N_8487,N_5674);
xor UO_858 (O_858,N_7696,N_9079);
nor UO_859 (O_859,N_8575,N_9866);
nor UO_860 (O_860,N_6932,N_9641);
xnor UO_861 (O_861,N_5470,N_6706);
nor UO_862 (O_862,N_7406,N_5406);
nand UO_863 (O_863,N_6951,N_5576);
or UO_864 (O_864,N_7498,N_8938);
xnor UO_865 (O_865,N_7124,N_9494);
nor UO_866 (O_866,N_5549,N_9354);
nand UO_867 (O_867,N_8069,N_5222);
nand UO_868 (O_868,N_9473,N_6288);
xnor UO_869 (O_869,N_8898,N_9830);
and UO_870 (O_870,N_8502,N_5177);
xnor UO_871 (O_871,N_7435,N_7635);
nor UO_872 (O_872,N_6242,N_7025);
nand UO_873 (O_873,N_6003,N_7706);
or UO_874 (O_874,N_5960,N_8713);
xnor UO_875 (O_875,N_7776,N_9843);
nand UO_876 (O_876,N_6982,N_5053);
and UO_877 (O_877,N_8212,N_5231);
and UO_878 (O_878,N_9386,N_9679);
and UO_879 (O_879,N_8398,N_8649);
nand UO_880 (O_880,N_8104,N_9377);
nor UO_881 (O_881,N_8210,N_6894);
nor UO_882 (O_882,N_6697,N_7144);
nor UO_883 (O_883,N_9805,N_7374);
xnor UO_884 (O_884,N_5939,N_7341);
nor UO_885 (O_885,N_9323,N_9328);
or UO_886 (O_886,N_5607,N_8415);
nand UO_887 (O_887,N_8404,N_8463);
and UO_888 (O_888,N_6412,N_5913);
nand UO_889 (O_889,N_6282,N_7546);
xor UO_890 (O_890,N_5143,N_7397);
xor UO_891 (O_891,N_7802,N_9440);
and UO_892 (O_892,N_5586,N_7344);
or UO_893 (O_893,N_7989,N_5692);
nor UO_894 (O_894,N_5252,N_7029);
nand UO_895 (O_895,N_8165,N_9827);
or UO_896 (O_896,N_8314,N_7708);
nand UO_897 (O_897,N_5373,N_8729);
and UO_898 (O_898,N_7869,N_8571);
nand UO_899 (O_899,N_8482,N_5758);
nor UO_900 (O_900,N_5559,N_6024);
and UO_901 (O_901,N_8823,N_7741);
xnor UO_902 (O_902,N_8813,N_7142);
nand UO_903 (O_903,N_7286,N_9496);
xor UO_904 (O_904,N_8912,N_8390);
xor UO_905 (O_905,N_8763,N_6779);
and UO_906 (O_906,N_7322,N_8247);
or UO_907 (O_907,N_7200,N_6717);
nand UO_908 (O_908,N_7889,N_9871);
nand UO_909 (O_909,N_6452,N_9093);
nand UO_910 (O_910,N_7657,N_6689);
or UO_911 (O_911,N_6177,N_7808);
or UO_912 (O_912,N_6566,N_8711);
xnor UO_913 (O_913,N_6873,N_5335);
nand UO_914 (O_914,N_6514,N_8293);
nand UO_915 (O_915,N_5376,N_8597);
or UO_916 (O_916,N_8280,N_5616);
nor UO_917 (O_917,N_8685,N_8431);
and UO_918 (O_918,N_8214,N_5424);
xor UO_919 (O_919,N_9664,N_7933);
xnor UO_920 (O_920,N_5441,N_6928);
xnor UO_921 (O_921,N_8142,N_7208);
and UO_922 (O_922,N_6825,N_8919);
nand UO_923 (O_923,N_6809,N_6625);
nor UO_924 (O_924,N_9119,N_8549);
xnor UO_925 (O_925,N_6876,N_7720);
or UO_926 (O_926,N_8256,N_9879);
xnor UO_927 (O_927,N_9781,N_6611);
nor UO_928 (O_928,N_8809,N_7728);
nor UO_929 (O_929,N_5446,N_8155);
or UO_930 (O_930,N_9520,N_6179);
or UO_931 (O_931,N_8728,N_6524);
or UO_932 (O_932,N_7666,N_7037);
and UO_933 (O_933,N_8224,N_8887);
and UO_934 (O_934,N_6192,N_5567);
nor UO_935 (O_935,N_6414,N_7180);
nand UO_936 (O_936,N_9490,N_8110);
nor UO_937 (O_937,N_6674,N_6303);
nor UO_938 (O_938,N_7351,N_7249);
nor UO_939 (O_939,N_6520,N_7811);
xor UO_940 (O_940,N_8302,N_5642);
or UO_941 (O_941,N_8060,N_8420);
xor UO_942 (O_942,N_5868,N_9259);
and UO_943 (O_943,N_6232,N_8221);
or UO_944 (O_944,N_6249,N_9204);
and UO_945 (O_945,N_8391,N_8873);
or UO_946 (O_946,N_6974,N_6927);
or UO_947 (O_947,N_7183,N_9059);
xnor UO_948 (O_948,N_9884,N_8124);
and UO_949 (O_949,N_5427,N_8312);
nand UO_950 (O_950,N_6601,N_6634);
nand UO_951 (O_951,N_9905,N_8739);
and UO_952 (O_952,N_8802,N_8087);
or UO_953 (O_953,N_6728,N_8354);
nand UO_954 (O_954,N_8550,N_6548);
xor UO_955 (O_955,N_9550,N_8062);
xor UO_956 (O_956,N_5360,N_6535);
and UO_957 (O_957,N_5421,N_9519);
xnor UO_958 (O_958,N_9661,N_6080);
nor UO_959 (O_959,N_8827,N_5929);
nand UO_960 (O_960,N_5329,N_6325);
xor UO_961 (O_961,N_6278,N_5769);
nand UO_962 (O_962,N_8922,N_6989);
or UO_963 (O_963,N_9345,N_5045);
or UO_964 (O_964,N_8207,N_7953);
xor UO_965 (O_965,N_7361,N_5548);
xor UO_966 (O_966,N_7138,N_9844);
nor UO_967 (O_967,N_7957,N_9367);
nand UO_968 (O_968,N_8574,N_5551);
xnor UO_969 (O_969,N_5730,N_5310);
or UO_970 (O_970,N_9487,N_5924);
or UO_971 (O_971,N_6964,N_6140);
xnor UO_972 (O_972,N_7534,N_6912);
xor UO_973 (O_973,N_8209,N_8797);
or UO_974 (O_974,N_6851,N_7912);
nand UO_975 (O_975,N_7379,N_8424);
nand UO_976 (O_976,N_5267,N_9940);
and UO_977 (O_977,N_9315,N_9934);
nor UO_978 (O_978,N_8319,N_8272);
nand UO_979 (O_979,N_5572,N_9083);
and UO_980 (O_980,N_8474,N_8904);
xnor UO_981 (O_981,N_7430,N_6091);
and UO_982 (O_982,N_9510,N_5668);
or UO_983 (O_983,N_5689,N_9727);
nor UO_984 (O_984,N_9100,N_5688);
nor UO_985 (O_985,N_8918,N_8377);
or UO_986 (O_986,N_9286,N_6371);
xor UO_987 (O_987,N_7007,N_6747);
nand UO_988 (O_988,N_6154,N_5694);
xor UO_989 (O_989,N_5272,N_8814);
nand UO_990 (O_990,N_5061,N_6350);
nand UO_991 (O_991,N_9447,N_5724);
nor UO_992 (O_992,N_6701,N_9266);
and UO_993 (O_993,N_7040,N_8514);
nand UO_994 (O_994,N_6367,N_8225);
and UO_995 (O_995,N_9811,N_7633);
xnor UO_996 (O_996,N_7348,N_9961);
or UO_997 (O_997,N_7387,N_5825);
and UO_998 (O_998,N_7607,N_8009);
nand UO_999 (O_999,N_9868,N_8454);
or UO_1000 (O_1000,N_8517,N_9872);
or UO_1001 (O_1001,N_9435,N_5587);
or UO_1002 (O_1002,N_5138,N_9445);
or UO_1003 (O_1003,N_5316,N_5249);
nor UO_1004 (O_1004,N_9002,N_5793);
or UO_1005 (O_1005,N_8795,N_7993);
and UO_1006 (O_1006,N_6726,N_5352);
xnor UO_1007 (O_1007,N_7779,N_9728);
nand UO_1008 (O_1008,N_5979,N_6145);
nor UO_1009 (O_1009,N_8356,N_6596);
or UO_1010 (O_1010,N_6886,N_9249);
nor UO_1011 (O_1011,N_8601,N_9056);
or UO_1012 (O_1012,N_8458,N_5346);
and UO_1013 (O_1013,N_7608,N_7644);
nand UO_1014 (O_1014,N_8704,N_9452);
or UO_1015 (O_1015,N_9613,N_5343);
nand UO_1016 (O_1016,N_7336,N_9264);
or UO_1017 (O_1017,N_7425,N_7401);
and UO_1018 (O_1018,N_7392,N_5383);
and UO_1019 (O_1019,N_5036,N_7549);
nand UO_1020 (O_1020,N_5554,N_6577);
nand UO_1021 (O_1021,N_7740,N_7499);
and UO_1022 (O_1022,N_8306,N_6162);
or UO_1023 (O_1023,N_7840,N_7198);
nand UO_1024 (O_1024,N_5386,N_9997);
and UO_1025 (O_1025,N_6677,N_5944);
and UO_1026 (O_1026,N_6115,N_7743);
xnor UO_1027 (O_1027,N_5805,N_8175);
nand UO_1028 (O_1028,N_8266,N_9331);
or UO_1029 (O_1029,N_7504,N_9709);
or UO_1030 (O_1030,N_6947,N_7495);
nor UO_1031 (O_1031,N_8863,N_9688);
xnor UO_1032 (O_1032,N_8806,N_7510);
nand UO_1033 (O_1033,N_5911,N_8038);
and UO_1034 (O_1034,N_8586,N_6664);
or UO_1035 (O_1035,N_5900,N_5033);
nand UO_1036 (O_1036,N_8969,N_5534);
nor UO_1037 (O_1037,N_8699,N_6925);
or UO_1038 (O_1038,N_8910,N_7284);
xnor UO_1039 (O_1039,N_7710,N_5101);
xnor UO_1040 (O_1040,N_8680,N_7496);
or UO_1041 (O_1041,N_6390,N_9631);
nor UO_1042 (O_1042,N_9639,N_9350);
nor UO_1043 (O_1043,N_7639,N_8821);
nor UO_1044 (O_1044,N_9230,N_8734);
and UO_1045 (O_1045,N_7789,N_6713);
xor UO_1046 (O_1046,N_8874,N_9685);
nand UO_1047 (O_1047,N_6941,N_5507);
nor UO_1048 (O_1048,N_7938,N_5614);
or UO_1049 (O_1049,N_9152,N_9203);
nor UO_1050 (O_1050,N_9461,N_5334);
xnor UO_1051 (O_1051,N_6153,N_5266);
xor UO_1052 (O_1052,N_5888,N_7367);
nand UO_1053 (O_1053,N_5185,N_9198);
xor UO_1054 (O_1054,N_8753,N_8931);
or UO_1055 (O_1055,N_7226,N_9233);
and UO_1056 (O_1056,N_9052,N_5731);
or UO_1057 (O_1057,N_5515,N_7891);
nor UO_1058 (O_1058,N_9554,N_7852);
xor UO_1059 (O_1059,N_7420,N_5306);
xnor UO_1060 (O_1060,N_8096,N_7078);
nand UO_1061 (O_1061,N_6773,N_8329);
nand UO_1062 (O_1062,N_9488,N_9436);
xor UO_1063 (O_1063,N_9400,N_7839);
or UO_1064 (O_1064,N_9865,N_6006);
nand UO_1065 (O_1065,N_6106,N_7490);
xor UO_1066 (O_1066,N_5130,N_8434);
nor UO_1067 (O_1067,N_6061,N_7611);
nand UO_1068 (O_1068,N_8049,N_6849);
nor UO_1069 (O_1069,N_5846,N_6101);
nand UO_1070 (O_1070,N_9111,N_7810);
nand UO_1071 (O_1071,N_7041,N_8423);
or UO_1072 (O_1072,N_8193,N_5763);
nand UO_1073 (O_1073,N_5733,N_9849);
xnor UO_1074 (O_1074,N_8299,N_7544);
or UO_1075 (O_1075,N_8383,N_8277);
nand UO_1076 (O_1076,N_8403,N_8488);
and UO_1077 (O_1077,N_5023,N_5855);
or UO_1078 (O_1078,N_5366,N_8030);
nor UO_1079 (O_1079,N_5134,N_6272);
or UO_1080 (O_1080,N_8432,N_9090);
xor UO_1081 (O_1081,N_7583,N_9581);
nand UO_1082 (O_1082,N_8389,N_9334);
or UO_1083 (O_1083,N_6473,N_9420);
nand UO_1084 (O_1084,N_9361,N_9274);
or UO_1085 (O_1085,N_7101,N_5870);
nor UO_1086 (O_1086,N_7896,N_7962);
and UO_1087 (O_1087,N_9740,N_7973);
nand UO_1088 (O_1088,N_5471,N_6326);
xor UO_1089 (O_1089,N_9254,N_6241);
nand UO_1090 (O_1090,N_7404,N_7585);
or UO_1091 (O_1091,N_6828,N_9236);
nand UO_1092 (O_1092,N_7968,N_9039);
or UO_1093 (O_1093,N_6269,N_7879);
nand UO_1094 (O_1094,N_7660,N_8002);
and UO_1095 (O_1095,N_8046,N_7000);
nor UO_1096 (O_1096,N_9821,N_8048);
and UO_1097 (O_1097,N_7306,N_6919);
or UO_1098 (O_1098,N_9557,N_7206);
nand UO_1099 (O_1099,N_6114,N_5032);
and UO_1100 (O_1100,N_9403,N_7285);
and UO_1101 (O_1101,N_9501,N_6905);
or UO_1102 (O_1102,N_9780,N_8097);
or UO_1103 (O_1103,N_5871,N_5076);
and UO_1104 (O_1104,N_7232,N_7997);
nand UO_1105 (O_1105,N_7237,N_8273);
or UO_1106 (O_1106,N_8152,N_7780);
or UO_1107 (O_1107,N_8876,N_6408);
xnor UO_1108 (O_1108,N_6902,N_7796);
nand UO_1109 (O_1109,N_5012,N_7876);
nand UO_1110 (O_1110,N_7469,N_5232);
nand UO_1111 (O_1111,N_6552,N_9915);
nand UO_1112 (O_1112,N_5561,N_8063);
and UO_1113 (O_1113,N_5962,N_7309);
and UO_1114 (O_1114,N_8352,N_8628);
nand UO_1115 (O_1115,N_8643,N_5029);
nand UO_1116 (O_1116,N_6586,N_7081);
xnor UO_1117 (O_1117,N_7804,N_6791);
nand UO_1118 (O_1118,N_5917,N_8026);
or UO_1119 (O_1119,N_7512,N_6759);
nor UO_1120 (O_1120,N_8584,N_7143);
nand UO_1121 (O_1121,N_5218,N_9509);
or UO_1122 (O_1122,N_6761,N_7797);
xnor UO_1123 (O_1123,N_5977,N_7455);
nor UO_1124 (O_1124,N_9282,N_9427);
nand UO_1125 (O_1125,N_9260,N_9006);
and UO_1126 (O_1126,N_7575,N_8235);
and UO_1127 (O_1127,N_7315,N_8095);
nor UO_1128 (O_1128,N_6543,N_9881);
and UO_1129 (O_1129,N_6445,N_7996);
nand UO_1130 (O_1130,N_8188,N_7543);
nor UO_1131 (O_1131,N_7829,N_5031);
and UO_1132 (O_1132,N_6553,N_5354);
nand UO_1133 (O_1133,N_5734,N_5190);
or UO_1134 (O_1134,N_8078,N_7317);
xnor UO_1135 (O_1135,N_6212,N_7807);
nand UO_1136 (O_1136,N_7626,N_8163);
or UO_1137 (O_1137,N_7723,N_5084);
and UO_1138 (O_1138,N_9055,N_6087);
xnor UO_1139 (O_1139,N_9904,N_7990);
and UO_1140 (O_1140,N_9474,N_7584);
nor UO_1141 (O_1141,N_9489,N_9170);
nand UO_1142 (O_1142,N_9789,N_5251);
nand UO_1143 (O_1143,N_9967,N_6792);
nand UO_1144 (O_1144,N_9446,N_6007);
or UO_1145 (O_1145,N_5741,N_5384);
and UO_1146 (O_1146,N_5460,N_6943);
nand UO_1147 (O_1147,N_6485,N_6110);
and UO_1148 (O_1148,N_7801,N_7194);
xnor UO_1149 (O_1149,N_7874,N_8037);
nand UO_1150 (O_1150,N_5170,N_6723);
xor UO_1151 (O_1151,N_7186,N_5324);
nand UO_1152 (O_1152,N_5024,N_9068);
xnor UO_1153 (O_1153,N_5678,N_8093);
or UO_1154 (O_1154,N_9585,N_6451);
or UO_1155 (O_1155,N_5684,N_5072);
and UO_1156 (O_1156,N_5480,N_5850);
xnor UO_1157 (O_1157,N_6903,N_9837);
nand UO_1158 (O_1158,N_7524,N_9114);
nand UO_1159 (O_1159,N_6073,N_5528);
xnor UO_1160 (O_1160,N_7464,N_8261);
or UO_1161 (O_1161,N_7974,N_8580);
nand UO_1162 (O_1162,N_9295,N_8151);
or UO_1163 (O_1163,N_6744,N_8849);
nand UO_1164 (O_1164,N_6725,N_9912);
nor UO_1165 (O_1165,N_7986,N_9952);
nor UO_1166 (O_1166,N_6771,N_8109);
nand UO_1167 (O_1167,N_7795,N_6691);
xnor UO_1168 (O_1168,N_5010,N_5241);
xor UO_1169 (O_1169,N_7003,N_9049);
nand UO_1170 (O_1170,N_8437,N_9666);
nor UO_1171 (O_1171,N_9414,N_9673);
xnor UO_1172 (O_1172,N_7655,N_8600);
and UO_1173 (O_1173,N_5482,N_9425);
and UO_1174 (O_1174,N_8036,N_8664);
nor UO_1175 (O_1175,N_6834,N_9428);
nor UO_1176 (O_1176,N_6879,N_5438);
and UO_1177 (O_1177,N_5999,N_5262);
xor UO_1178 (O_1178,N_5928,N_8816);
nand UO_1179 (O_1179,N_9819,N_6393);
or UO_1180 (O_1180,N_5505,N_7718);
and UO_1181 (O_1181,N_6647,N_7242);
and UO_1182 (O_1182,N_5897,N_5867);
or UO_1183 (O_1183,N_9778,N_6720);
nand UO_1184 (O_1184,N_8342,N_6126);
xor UO_1185 (O_1185,N_5986,N_5456);
nand UO_1186 (O_1186,N_5374,N_8830);
xnor UO_1187 (O_1187,N_7238,N_9529);
and UO_1188 (O_1188,N_8127,N_5970);
nor UO_1189 (O_1189,N_6966,N_8230);
xnor UO_1190 (O_1190,N_5126,N_5417);
or UO_1191 (O_1191,N_7110,N_5571);
nor UO_1192 (O_1192,N_9212,N_5244);
or UO_1193 (O_1193,N_9149,N_8443);
nor UO_1194 (O_1194,N_7679,N_8045);
or UO_1195 (O_1195,N_5834,N_7185);
or UO_1196 (O_1196,N_7126,N_9069);
nand UO_1197 (O_1197,N_9694,N_8387);
nor UO_1198 (O_1198,N_9544,N_7503);
nand UO_1199 (O_1199,N_8158,N_8073);
xor UO_1200 (O_1200,N_8567,N_9605);
xor UO_1201 (O_1201,N_9313,N_9054);
or UO_1202 (O_1202,N_5004,N_9568);
nand UO_1203 (O_1203,N_9478,N_6358);
or UO_1204 (O_1204,N_9845,N_5629);
and UO_1205 (O_1205,N_9956,N_9416);
and UO_1206 (O_1206,N_9970,N_6098);
and UO_1207 (O_1207,N_6536,N_6570);
nor UO_1208 (O_1208,N_9894,N_6908);
and UO_1209 (O_1209,N_7573,N_9008);
xnor UO_1210 (O_1210,N_5320,N_8973);
xnor UO_1211 (O_1211,N_8105,N_8804);
nand UO_1212 (O_1212,N_8239,N_8541);
xnor UO_1213 (O_1213,N_6986,N_7001);
nand UO_1214 (O_1214,N_6094,N_5516);
or UO_1215 (O_1215,N_7478,N_9466);
xor UO_1216 (O_1216,N_5064,N_7236);
and UO_1217 (O_1217,N_8249,N_6666);
nor UO_1218 (O_1218,N_8953,N_8635);
nand UO_1219 (O_1219,N_8941,N_8252);
or UO_1220 (O_1220,N_7158,N_5918);
xor UO_1221 (O_1221,N_8362,N_8006);
or UO_1222 (O_1222,N_5112,N_6156);
nand UO_1223 (O_1223,N_9503,N_7620);
nor UO_1224 (O_1224,N_9462,N_7961);
xor UO_1225 (O_1225,N_8817,N_9335);
nand UO_1226 (O_1226,N_6419,N_6512);
and UO_1227 (O_1227,N_7725,N_6136);
nor UO_1228 (O_1228,N_7788,N_8570);
nand UO_1229 (O_1229,N_5627,N_9123);
nor UO_1230 (O_1230,N_9136,N_8871);
or UO_1231 (O_1231,N_8889,N_7955);
nand UO_1232 (O_1232,N_6185,N_5443);
nand UO_1233 (O_1233,N_6537,N_5797);
xnor UO_1234 (O_1234,N_6567,N_6978);
xor UO_1235 (O_1235,N_6182,N_6287);
nand UO_1236 (O_1236,N_8262,N_7247);
xnor UO_1237 (O_1237,N_5542,N_9239);
xnor UO_1238 (O_1238,N_9921,N_7005);
or UO_1239 (O_1239,N_6377,N_9379);
xor UO_1240 (O_1240,N_6299,N_9516);
nor UO_1241 (O_1241,N_7651,N_7157);
nor UO_1242 (O_1242,N_9957,N_8967);
and UO_1243 (O_1243,N_5098,N_6276);
or UO_1244 (O_1244,N_5886,N_5261);
nand UO_1245 (O_1245,N_9196,N_9163);
xnor UO_1246 (O_1246,N_6561,N_8448);
or UO_1247 (O_1247,N_9327,N_5090);
xnor UO_1248 (O_1248,N_6253,N_5522);
or UO_1249 (O_1249,N_6564,N_5714);
or UO_1250 (O_1250,N_6571,N_5715);
nor UO_1251 (O_1251,N_5207,N_5673);
or UO_1252 (O_1252,N_7083,N_6048);
nor UO_1253 (O_1253,N_9162,N_6995);
nor UO_1254 (O_1254,N_8608,N_9405);
nor UO_1255 (O_1255,N_6980,N_7303);
nand UO_1256 (O_1256,N_6670,N_7075);
nand UO_1257 (O_1257,N_6133,N_6946);
and UO_1258 (O_1258,N_8875,N_7421);
nor UO_1259 (O_1259,N_6811,N_7667);
nor UO_1260 (O_1260,N_5641,N_8396);
xor UO_1261 (O_1261,N_6604,N_7930);
nor UO_1262 (O_1262,N_5660,N_5967);
nand UO_1263 (O_1263,N_9577,N_8746);
xnor UO_1264 (O_1264,N_7203,N_7031);
nand UO_1265 (O_1265,N_9296,N_6324);
or UO_1266 (O_1266,N_6099,N_8725);
xnor UO_1267 (O_1267,N_5381,N_5721);
xnor UO_1268 (O_1268,N_6248,N_8786);
nor UO_1269 (O_1269,N_9312,N_7103);
xnor UO_1270 (O_1270,N_9522,N_9060);
and UO_1271 (O_1271,N_9897,N_8560);
or UO_1272 (O_1272,N_8696,N_9597);
nand UO_1273 (O_1273,N_7812,N_8596);
or UO_1274 (O_1274,N_9193,N_5341);
nand UO_1275 (O_1275,N_9587,N_6012);
or UO_1276 (O_1276,N_7732,N_9166);
or UO_1277 (O_1277,N_7529,N_6954);
nor UO_1278 (O_1278,N_8123,N_5476);
xnor UO_1279 (O_1279,N_8079,N_6904);
nand UO_1280 (O_1280,N_9622,N_5123);
xor UO_1281 (O_1281,N_9316,N_8118);
nor UO_1282 (O_1282,N_9276,N_5909);
nor UO_1283 (O_1283,N_6395,N_8399);
and UO_1284 (O_1284,N_6742,N_7502);
or UO_1285 (O_1285,N_7816,N_5580);
nand UO_1286 (O_1286,N_9411,N_5877);
or UO_1287 (O_1287,N_7717,N_8359);
nor UO_1288 (O_1288,N_6716,N_8851);
nor UO_1289 (O_1289,N_6207,N_8498);
nand UO_1290 (O_1290,N_7821,N_9726);
nor UO_1291 (O_1291,N_5003,N_6865);
and UO_1292 (O_1292,N_6307,N_8589);
or UO_1293 (O_1293,N_8727,N_7149);
nor UO_1294 (O_1294,N_7752,N_6704);
xnor UO_1295 (O_1295,N_8868,N_5840);
xor UO_1296 (O_1296,N_6550,N_9084);
and UO_1297 (O_1297,N_8166,N_5759);
nor UO_1298 (O_1298,N_9222,N_8954);
nor UO_1299 (O_1299,N_9333,N_5233);
xor UO_1300 (O_1300,N_7900,N_7436);
nor UO_1301 (O_1301,N_5431,N_6329);
xor UO_1302 (O_1302,N_6449,N_5115);
and UO_1303 (O_1303,N_7446,N_8627);
xor UO_1304 (O_1304,N_8366,N_7998);
or UO_1305 (O_1305,N_9989,N_5811);
nor UO_1306 (O_1306,N_5089,N_8380);
nand UO_1307 (O_1307,N_6710,N_9742);
nand UO_1308 (O_1308,N_7515,N_8976);
or UO_1309 (O_1309,N_8469,N_6506);
or UO_1310 (O_1310,N_6342,N_5865);
xor UO_1311 (O_1311,N_9223,N_9776);
xor UO_1312 (O_1312,N_5590,N_6842);
nand UO_1313 (O_1313,N_8232,N_9601);
nand UO_1314 (O_1314,N_5995,N_5593);
nor UO_1315 (O_1315,N_6914,N_9283);
and UO_1316 (O_1316,N_8259,N_5370);
nand UO_1317 (O_1317,N_9893,N_7903);
and UO_1318 (O_1318,N_7064,N_7823);
nor UO_1319 (O_1319,N_9838,N_5532);
and UO_1320 (O_1320,N_7680,N_7590);
and UO_1321 (O_1321,N_6360,N_5603);
or UO_1322 (O_1322,N_9262,N_5702);
nand UO_1323 (O_1323,N_6766,N_9869);
nor UO_1324 (O_1324,N_9434,N_6877);
xnor UO_1325 (O_1325,N_5236,N_6575);
xor UO_1326 (O_1326,N_7349,N_7815);
nand UO_1327 (O_1327,N_8492,N_8653);
and UO_1328 (O_1328,N_8905,N_5765);
or UO_1329 (O_1329,N_9194,N_7555);
and UO_1330 (O_1330,N_8762,N_5519);
or UO_1331 (O_1331,N_9342,N_8162);
xnor UO_1332 (O_1332,N_9644,N_5111);
and UO_1333 (O_1333,N_9429,N_6204);
xor UO_1334 (O_1334,N_6067,N_8951);
or UO_1335 (O_1335,N_8219,N_8933);
and UO_1336 (O_1336,N_8670,N_7327);
nor UO_1337 (O_1337,N_9620,N_6968);
or UO_1338 (O_1338,N_8385,N_7454);
or UO_1339 (O_1339,N_7165,N_7523);
nor UO_1340 (O_1340,N_7259,N_5697);
nor UO_1341 (O_1341,N_8547,N_8650);
xor UO_1342 (O_1342,N_5489,N_9498);
nor UO_1343 (O_1343,N_7956,N_8893);
nor UO_1344 (O_1344,N_6019,N_5711);
and UO_1345 (O_1345,N_9225,N_8183);
nor UO_1346 (O_1346,N_7913,N_5980);
xor UO_1347 (O_1347,N_7951,N_6961);
or UO_1348 (O_1348,N_5478,N_5444);
nor UO_1349 (O_1349,N_8519,N_5887);
nor UO_1350 (O_1350,N_8961,N_5372);
nor UO_1351 (O_1351,N_7043,N_6373);
and UO_1352 (O_1352,N_8965,N_6763);
and UO_1353 (O_1353,N_6124,N_7733);
nor UO_1354 (O_1354,N_6446,N_7881);
nand UO_1355 (O_1355,N_6703,N_6129);
nor UO_1356 (O_1356,N_7676,N_7251);
xor UO_1357 (O_1357,N_5879,N_9394);
nand UO_1358 (O_1358,N_9098,N_8176);
or UO_1359 (O_1359,N_9832,N_9761);
xor UO_1360 (O_1360,N_5771,N_9786);
nor UO_1361 (O_1361,N_6497,N_7643);
or UO_1362 (O_1362,N_7566,N_5844);
or UO_1363 (O_1363,N_7966,N_9134);
nand UO_1364 (O_1364,N_7438,N_5181);
nand UO_1365 (O_1365,N_7520,N_9081);
and UO_1366 (O_1366,N_5362,N_6938);
or UO_1367 (O_1367,N_8513,N_8484);
and UO_1368 (O_1368,N_6973,N_9191);
nand UO_1369 (O_1369,N_8796,N_5107);
xor UO_1370 (O_1370,N_8507,N_5156);
or UO_1371 (O_1371,N_9005,N_8347);
nor UO_1372 (O_1372,N_7207,N_5208);
nor UO_1373 (O_1373,N_9527,N_6889);
nand UO_1374 (O_1374,N_7113,N_8563);
and UO_1375 (O_1375,N_5077,N_8701);
and UO_1376 (O_1376,N_9133,N_8333);
nor UO_1377 (O_1377,N_7623,N_6764);
xor UO_1378 (O_1378,N_7087,N_8808);
xnor UO_1379 (O_1379,N_9028,N_6032);
xnor UO_1380 (O_1380,N_9979,N_5904);
and UO_1381 (O_1381,N_8159,N_5751);
nand UO_1382 (O_1382,N_9703,N_5401);
and UO_1383 (O_1383,N_9792,N_7209);
xor UO_1384 (O_1384,N_6379,N_6539);
or UO_1385 (O_1385,N_5087,N_6482);
xnor UO_1386 (O_1386,N_6285,N_7527);
nand UO_1387 (O_1387,N_7330,N_6335);
or UO_1388 (O_1388,N_5643,N_9486);
nand UO_1389 (O_1389,N_9353,N_9546);
and UO_1390 (O_1390,N_7721,N_7982);
xnor UO_1391 (O_1391,N_6381,N_8920);
and UO_1392 (O_1392,N_5975,N_8477);
nor UO_1393 (O_1393,N_7536,N_6229);
or UO_1394 (O_1394,N_5595,N_5048);
or UO_1395 (O_1395,N_9500,N_6280);
nor UO_1396 (O_1396,N_5782,N_7255);
or UO_1397 (O_1397,N_8135,N_6769);
or UO_1398 (O_1398,N_5125,N_8774);
nand UO_1399 (O_1399,N_9788,N_5491);
nor UO_1400 (O_1400,N_6418,N_7094);
and UO_1401 (O_1401,N_7908,N_6444);
xor UO_1402 (O_1402,N_8503,N_8371);
or UO_1403 (O_1403,N_6043,N_6490);
nor UO_1404 (O_1404,N_7489,N_8035);
nand UO_1405 (O_1405,N_7734,N_6355);
nand UO_1406 (O_1406,N_6557,N_7095);
nand UO_1407 (O_1407,N_7859,N_9153);
or UO_1408 (O_1408,N_5365,N_9823);
nand UO_1409 (O_1409,N_7709,N_9280);
and UO_1410 (O_1410,N_5514,N_8531);
or UO_1411 (O_1411,N_7783,N_8270);
nor UO_1412 (O_1412,N_7424,N_5430);
and UO_1413 (O_1413,N_9021,N_8678);
and UO_1414 (O_1414,N_8908,N_9067);
or UO_1415 (O_1415,N_5626,N_7118);
nor UO_1416 (O_1416,N_9007,N_9877);
xor UO_1417 (O_1417,N_8117,N_5186);
and UO_1418 (O_1418,N_9151,N_6795);
nand UO_1419 (O_1419,N_5479,N_6175);
nand UO_1420 (O_1420,N_7316,N_7297);
or UO_1421 (O_1421,N_8989,N_5777);
xor UO_1422 (O_1422,N_8652,N_7339);
nand UO_1423 (O_1423,N_7346,N_8667);
and UO_1424 (O_1424,N_9025,N_6609);
xnor UO_1425 (O_1425,N_5296,N_7100);
and UO_1426 (O_1426,N_7116,N_8042);
or UO_1427 (O_1427,N_7019,N_8160);
and UO_1428 (O_1428,N_8005,N_5570);
or UO_1429 (O_1429,N_9058,N_6268);
and UO_1430 (O_1430,N_6560,N_9439);
or UO_1431 (O_1431,N_7662,N_7787);
xor UO_1432 (O_1432,N_7482,N_8369);
or UO_1433 (O_1433,N_5245,N_7622);
nand UO_1434 (O_1434,N_8460,N_7554);
and UO_1435 (O_1435,N_8607,N_6959);
nor UO_1436 (O_1436,N_9678,N_7224);
xnor UO_1437 (O_1437,N_8682,N_6022);
nand UO_1438 (O_1438,N_8413,N_5474);
and UO_1439 (O_1439,N_9580,N_9537);
or UO_1440 (O_1440,N_5378,N_5224);
and UO_1441 (O_1441,N_7884,N_7470);
xnor UO_1442 (O_1442,N_9238,N_7685);
and UO_1443 (O_1443,N_8493,N_5736);
and UO_1444 (O_1444,N_8996,N_8208);
nand UO_1445 (O_1445,N_9063,N_6336);
or UO_1446 (O_1446,N_7937,N_8582);
xnor UO_1447 (O_1447,N_5099,N_8428);
nor UO_1448 (O_1448,N_6164,N_6226);
xor UO_1449 (O_1449,N_9146,N_9485);
nand UO_1450 (O_1450,N_6044,N_7614);
nand UO_1451 (O_1451,N_6477,N_6546);
xor UO_1452 (O_1452,N_9003,N_9142);
nand UO_1453 (O_1453,N_9900,N_5718);
or UO_1454 (O_1454,N_6480,N_8226);
nor UO_1455 (O_1455,N_8866,N_5832);
nor UO_1456 (O_1456,N_8441,N_5070);
and UO_1457 (O_1457,N_7629,N_8065);
or UO_1458 (O_1458,N_9713,N_9187);
xnor UO_1459 (O_1459,N_8846,N_6047);
nor UO_1460 (O_1460,N_7221,N_5606);
nor UO_1461 (O_1461,N_6778,N_9962);
nand UO_1462 (O_1462,N_5959,N_9981);
nor UO_1463 (O_1463,N_6297,N_9073);
xor UO_1464 (O_1464,N_6646,N_8917);
xor UO_1465 (O_1465,N_8442,N_7917);
nand UO_1466 (O_1466,N_8921,N_7311);
or UO_1467 (O_1467,N_6595,N_6998);
or UO_1468 (O_1468,N_9200,N_6361);
nor UO_1469 (O_1469,N_7766,N_7270);
and UO_1470 (O_1470,N_5127,N_8743);
nor UO_1471 (O_1471,N_5858,N_6589);
nor UO_1472 (O_1472,N_7600,N_8511);
xor UO_1473 (O_1473,N_7073,N_8546);
nand UO_1474 (O_1474,N_6862,N_8778);
nand UO_1475 (O_1475,N_8521,N_8662);
xor UO_1476 (O_1476,N_9783,N_6095);
or UO_1477 (O_1477,N_8886,N_6937);
and UO_1478 (O_1478,N_9653,N_8197);
xnor UO_1479 (O_1479,N_8187,N_7403);
or UO_1480 (O_1480,N_5110,N_7045);
nand UO_1481 (O_1481,N_7545,N_9360);
nor UO_1482 (O_1482,N_5426,N_9399);
nand UO_1483 (O_1483,N_7195,N_8339);
nor UO_1484 (O_1484,N_6607,N_6699);
and UO_1485 (O_1485,N_8779,N_6174);
xnor UO_1486 (O_1486,N_8421,N_6389);
or UO_1487 (O_1487,N_9135,N_9841);
and UO_1488 (O_1488,N_9261,N_9307);
and UO_1489 (O_1489,N_6934,N_5436);
or UO_1490 (O_1490,N_7530,N_6103);
nor UO_1491 (O_1491,N_8267,N_9324);
and UO_1492 (O_1492,N_9582,N_9497);
nand UO_1493 (O_1493,N_9692,N_8956);
nand UO_1494 (O_1494,N_9401,N_7301);
and UO_1495 (O_1495,N_8508,N_9882);
nand UO_1496 (O_1496,N_8053,N_8481);
nor UO_1497 (O_1497,N_5412,N_5325);
and UO_1498 (O_1498,N_5043,N_6531);
nand UO_1499 (O_1499,N_7202,N_8581);
endmodule